magic
tech sky130A
magscale 1 2
timestamp 1717201555
<< metal1 >>
rect 21110 9160 21506 9190
rect 12884 8850 12890 9150
rect 13190 8850 13196 9150
rect 21110 8860 21140 9160
rect 21440 8860 21506 9160
rect 12890 8650 13190 8850
rect 12890 8344 13190 8350
rect 21110 8660 21506 8860
rect 21110 8360 21140 8660
rect 21440 8360 21506 8660
rect 21110 7520 21506 8360
rect 12884 7210 12890 7510
rect 13190 7210 13196 7510
rect 21110 7220 21140 7520
rect 21440 7220 21506 7520
rect 21110 6810 21506 7220
rect 12884 6500 12890 6800
rect 13190 6500 13196 6800
rect 21110 6510 21140 6810
rect 21440 6510 21506 6810
rect 21110 6130 21506 6510
rect 12884 5820 12890 6120
rect 13190 5820 13196 6120
rect 21110 5830 21140 6130
rect 21440 5830 21506 6130
rect 21110 5270 21506 5830
rect 12890 5260 13190 5266
rect 12884 4960 12890 5260
rect 13190 4960 13196 5260
rect 21110 4970 21140 5270
rect 21440 4970 21506 5270
rect 12890 4954 13190 4960
rect 21110 4390 21506 4970
rect 12884 4080 12890 4380
rect 13190 4080 13196 4380
rect 21110 4090 21140 4390
rect 21440 4090 21506 4390
rect 21110 3410 21506 4090
rect 12884 3100 12890 3400
rect 13190 3100 13196 3400
rect 21110 3110 21140 3410
rect 21440 3110 21506 3410
rect 12890 2690 13190 3100
rect 12890 2384 13190 2390
rect 21110 2700 21506 3110
rect 21110 2400 21140 2700
rect 21440 2400 21506 2700
rect 21110 2170 21506 2400
rect 29100 9150 29480 9170
rect 29100 8850 29130 9150
rect 29430 8850 29480 9150
rect 29100 8650 29480 8850
rect 29100 8350 29130 8650
rect 29430 8350 29480 8650
rect 29100 7510 29480 8350
rect 29100 7210 29130 7510
rect 29430 7210 29480 7510
rect 29100 6800 29480 7210
rect 29100 6500 29130 6800
rect 29430 6500 29480 6800
rect 29100 6120 29480 6500
rect 29100 5820 29130 6120
rect 29430 5820 29480 6120
rect 29100 5260 29480 5820
rect 29100 4960 29130 5260
rect 29430 4960 29480 5260
rect 29100 4380 29480 4960
rect 29100 4080 29130 4380
rect 29430 4080 29480 4380
rect 29100 3400 29480 4080
rect 29100 3100 29130 3400
rect 29430 3100 29480 3400
rect 29100 2690 29480 3100
rect 29100 2390 29130 2690
rect 29430 2390 29480 2690
rect 29100 2180 29480 2390
rect 24831 1319 25249 1325
rect 16208 1103 16740 1123
rect 16878 1103 17343 1109
rect 8328 901 8772 907
rect 7648 457 8328 901
rect 16208 658 16878 1103
rect 16740 638 16878 658
rect 24071 901 24831 1319
rect 24831 895 25249 901
rect 16878 632 17343 638
rect 8328 451 8772 457
<< via1 >>
rect 12890 8850 13190 9150
rect 21140 8860 21440 9160
rect 12890 8350 13190 8650
rect 21140 8360 21440 8660
rect 12890 7210 13190 7510
rect 21140 7220 21440 7520
rect 12890 6500 13190 6800
rect 21140 6510 21440 6810
rect 12890 5820 13190 6120
rect 21140 5830 21440 6130
rect 12890 4960 13190 5260
rect 21140 4970 21440 5270
rect 12890 4080 13190 4380
rect 21140 4090 21440 4390
rect 12890 3100 13190 3400
rect 21140 3110 21440 3410
rect 12890 2390 13190 2690
rect 21140 2400 21440 2700
rect 29130 8850 29430 9150
rect 29130 8350 29430 8650
rect 29130 7210 29430 7510
rect 29130 6500 29430 6800
rect 29130 5820 29430 6120
rect 29130 4960 29430 5260
rect 29130 4080 29430 4380
rect 29130 3100 29430 3400
rect 29130 2390 29430 2690
rect 8328 457 8772 901
rect 16878 638 17343 1103
rect 24831 901 25249 1319
<< metal2 >>
rect 15692 44180 15748 44187
rect 15690 44178 15750 44180
rect 15690 44122 15692 44178
rect 15748 44122 15750 44178
rect 5390 43588 5450 43590
rect 5383 43532 5392 43588
rect 5448 43532 5457 43588
rect 5390 43138 5450 43532
rect 6860 43448 6920 43450
rect 6853 43392 6862 43448
rect 6918 43392 6927 43448
rect 5386 43020 5450 43138
rect 6860 43058 6920 43392
rect 8330 43308 8390 43310
rect 8323 43252 8332 43308
rect 8388 43252 8397 43308
rect 5386 42752 5442 43020
rect 6858 42930 6920 43058
rect 8330 42940 8390 43252
rect 12740 42988 12800 42990
rect 9802 42980 9858 42987
rect 9800 42978 9860 42980
rect 11270 42978 11330 42980
rect 6858 42672 6914 42930
rect 8330 42702 8386 42940
rect 9800 42922 9802 42978
rect 9858 42922 9860 42978
rect 11263 42922 11272 42978
rect 11328 42922 11337 42978
rect 12733 42932 12742 42988
rect 12798 42932 12807 42988
rect 14210 42978 14270 42980
rect 9800 42740 9860 42922
rect 11270 42740 11330 42922
rect 12740 42818 12800 42932
rect 14203 42922 14212 42978
rect 14268 42922 14277 42978
rect 12740 42760 12802 42818
rect 12746 42740 12802 42760
rect 14210 42808 14270 42922
rect 15690 42920 15750 44122
rect 17160 44038 17220 44040
rect 17153 43982 17162 44038
rect 17218 43982 17227 44038
rect 14210 42740 14274 42808
rect 15690 42740 15746 42920
rect 17160 42740 17220 43982
rect 18632 43910 18688 43917
rect 18630 43908 18690 43910
rect 18630 43852 18632 43908
rect 18688 43852 18690 43908
rect 18630 42740 18690 43852
rect 20112 43770 20168 43777
rect 20110 43768 20170 43770
rect 20110 43712 20112 43768
rect 20168 43712 20170 43768
rect 20110 42768 20170 43712
rect 21582 43630 21638 43637
rect 21580 43628 21640 43630
rect 21580 43572 21582 43628
rect 21638 43572 21640 43628
rect 21580 42778 21640 43572
rect 23052 43480 23108 43487
rect 20106 42740 20170 42768
rect 21578 42740 21640 42778
rect 23050 43478 23110 43480
rect 23050 43422 23052 43478
rect 23108 43422 23110 43478
rect 23050 42740 23110 43422
rect 24522 43350 24578 43357
rect 24520 43348 24580 43350
rect 24520 43292 24522 43348
rect 24578 43292 24580 43348
rect 24520 42740 24580 43292
rect 25990 43218 26050 43220
rect 25983 43162 25992 43218
rect 26048 43162 26057 43218
rect 25990 42740 26050 43162
rect 27460 43092 27516 43099
rect 27458 43090 27518 43092
rect 27458 43034 27460 43090
rect 27516 43034 27518 43090
rect 27458 42740 27518 43034
rect 28938 42958 28994 42965
rect 28936 42956 28996 42958
rect 28936 42900 28938 42956
rect 28994 42900 28996 42956
rect 28936 42740 28996 42900
rect 30514 42828 30570 42835
rect 30408 42826 30572 42828
rect 30408 42770 30514 42826
rect 30570 42770 30572 42826
rect 30408 42768 30572 42770
rect 30408 42740 30468 42768
rect 30514 42761 30570 42768
rect 24522 42722 24578 42740
rect 5754 9948 5810 10940
rect 6306 10358 6362 10974
rect 6858 10478 6914 10922
rect 7410 10578 7466 10940
rect 7962 10688 8018 10952
rect 8514 10798 8570 10956
rect 8514 10742 8768 10798
rect 7962 10632 8248 10688
rect 7410 10522 7848 10578
rect 6858 10422 7528 10478
rect 6306 10302 7228 10358
rect 5754 9892 6948 9948
rect 7172 9782 7228 10302
rect 7472 9782 7528 10422
rect 7792 9792 7848 10522
rect 8192 9782 8248 10632
rect 8712 9812 8768 10742
rect 9066 9848 9122 10996
rect 9066 9792 9308 9848
rect 9618 9792 9674 11014
rect 10170 9848 10226 10966
rect 10722 10068 10778 11000
rect 11274 10398 11330 10962
rect 9962 9792 10226 9848
rect 10432 10012 10778 10068
rect 10842 10342 11330 10398
rect 10432 9802 10488 10012
rect 10842 9802 10898 10342
rect 11826 10298 11882 10970
rect 11232 10242 11882 10298
rect 11232 9812 11288 10242
rect 12378 10188 12434 10942
rect 11602 10132 12434 10188
rect 11602 9802 11658 10132
rect 12930 10078 12986 10940
rect 12040 10022 12986 10078
rect 12040 9786 12096 10022
rect 13482 9956 13538 10900
rect 14034 10438 14090 10932
rect 14586 10558 14642 10980
rect 15138 10688 15194 10946
rect 15690 10788 15746 10980
rect 15690 10732 16098 10788
rect 15138 10632 15768 10688
rect 14586 10502 15468 10558
rect 14034 10382 15078 10438
rect 12294 9900 13538 9956
rect 15022 9952 15078 10382
rect 15412 9952 15468 10502
rect 15712 9952 15768 10632
rect 16042 9952 16098 10732
rect 16242 10548 16298 10940
rect 16242 10492 16488 10548
rect 16432 9962 16488 10492
rect 16794 10028 16850 10990
rect 17346 10388 17402 10962
rect 17346 10332 17468 10388
rect 16794 9972 17118 10028
rect 17412 9952 17468 10332
rect 17898 9962 17954 10966
rect 18450 10498 18506 10972
rect 19002 10628 19058 10956
rect 18312 10442 18506 10498
rect 18672 10572 19058 10628
rect 18312 9962 18368 10442
rect 18672 9962 18728 10572
rect 19554 10518 19610 10956
rect 19082 10462 19610 10518
rect 19082 9962 19138 10462
rect 20106 10418 20162 10966
rect 19472 10362 20162 10418
rect 19472 9972 19528 10362
rect 20658 10314 20714 10946
rect 19852 10258 20714 10314
rect 19852 9972 19908 10258
rect 21210 10222 21266 10932
rect 20280 10166 21266 10222
rect 20280 9958 20336 10166
rect 21762 10092 21818 10912
rect 22314 10578 22370 10900
rect 22866 10668 22922 10900
rect 23418 10668 23474 10900
rect 23970 10678 24026 10900
rect 22866 10612 23348 10668
rect 23418 10612 23858 10668
rect 23970 10622 24168 10678
rect 22314 10522 23048 10578
rect 22992 10288 23048 10522
rect 23292 10288 23348 10612
rect 22992 10232 23148 10288
rect 23292 10232 23568 10288
rect 23802 10242 23858 10612
rect 24112 10242 24168 10622
rect 24522 10298 24578 10900
rect 25074 10318 25130 10938
rect 25626 10518 25682 10928
rect 26178 10518 26234 10928
rect 26730 10608 26786 10908
rect 27282 10688 27338 10938
rect 27834 10798 27890 10918
rect 25022 10308 25130 10318
rect 24412 10242 24578 10298
rect 24962 10252 25130 10308
rect 25482 10462 25682 10518
rect 25912 10462 26234 10518
rect 26282 10552 26786 10608
rect 26922 10632 27338 10688
rect 27622 10742 27890 10798
rect 25482 10242 25538 10462
rect 25912 10232 25968 10462
rect 26282 10252 26338 10552
rect 26922 10518 26978 10632
rect 27622 10598 27678 10742
rect 28386 10698 28442 10908
rect 26632 10462 26978 10518
rect 27042 10542 27678 10598
rect 27782 10642 28442 10698
rect 26632 10272 26688 10462
rect 27042 10252 27098 10542
rect 27782 10498 27838 10642
rect 28938 10598 28994 10938
rect 27442 10442 27838 10498
rect 27942 10542 28994 10598
rect 27442 10312 27498 10442
rect 27942 10388 27998 10542
rect 29490 10498 29546 10900
rect 27792 10332 27998 10388
rect 28262 10442 29546 10498
rect 28262 10262 28318 10442
rect 30042 10298 30098 10928
rect 28522 10242 30098 10298
rect 20556 10036 21818 10092
rect 22325 9730 22615 9734
rect 22320 9725 22620 9730
rect 22320 9435 22325 9725
rect 22615 9435 22620 9725
rect 14375 9420 14665 9424
rect 14370 9415 14670 9420
rect 6125 9280 6415 9284
rect 6120 9275 6420 9280
rect 6120 8985 6125 9275
rect 6415 8985 6420 9275
rect 6120 8380 6420 8985
rect 12890 9150 13190 9156
rect 12890 8650 13190 8850
rect 14370 9125 14375 9415
rect 14665 9125 14670 9415
rect 14370 8730 14670 9125
rect 21140 9160 21440 9166
rect 22320 8950 22620 9435
rect 29130 9150 29430 9156
rect 21140 8660 21440 8860
rect 12884 8350 12890 8650
rect 13190 8350 13196 8650
rect 21134 8360 21140 8660
rect 21440 8360 21446 8660
rect 29130 8650 29430 8850
rect 12890 8075 13190 8350
rect 12890 7785 12895 8075
rect 13185 7785 13190 8075
rect 12890 7510 13190 7785
rect 12890 6800 13190 7210
rect 12890 6120 13190 6500
rect 12890 5260 13190 5820
rect 21140 8085 21440 8360
rect 29124 8350 29130 8650
rect 29430 8350 29436 8650
rect 21140 7795 21145 8085
rect 21435 7795 21440 8085
rect 21140 7520 21440 7795
rect 21140 6810 21440 7220
rect 21140 6130 21440 6510
rect 21140 5270 21440 5830
rect 29130 8075 29430 8350
rect 29130 7785 29135 8075
rect 29425 7785 29430 8075
rect 29130 7510 29430 7785
rect 29130 6800 29430 7210
rect 29130 6120 29430 6500
rect 12884 4960 12890 5260
rect 13190 4960 13196 5260
rect 21134 4970 21140 5270
rect 21440 4970 21446 5270
rect 29130 5260 29430 5820
rect 12890 4380 13190 4960
rect 12890 3400 13190 4080
rect 12890 2690 13190 3100
rect 21140 4390 21440 4970
rect 29124 4960 29130 5260
rect 29430 4960 29436 5260
rect 21140 3410 21440 4090
rect 21140 2700 21440 3110
rect 29130 4380 29430 4960
rect 29130 3400 29430 4080
rect 12884 2390 12890 2690
rect 13190 2390 13196 2690
rect 21134 2400 21140 2700
rect 21440 2400 21446 2700
rect 29130 2690 29430 3100
rect 12890 2200 13190 2390
rect 21140 2210 21440 2400
rect 29124 2390 29130 2690
rect 29430 2390 29436 2690
rect 29130 2200 29430 2390
rect 25566 1319 25974 1323
rect 17493 1103 17948 1107
rect 8883 901 9317 905
rect 8322 457 8328 901
rect 8772 896 9322 901
rect 8772 462 8883 896
rect 9317 462 9322 896
rect 16872 638 16878 1103
rect 17343 1098 17953 1103
rect 17343 643 17493 1098
rect 17948 643 17953 1098
rect 24825 901 24831 1319
rect 25249 1314 25979 1319
rect 25249 906 25566 1314
rect 25974 906 25979 1314
rect 25249 901 25979 906
rect 25566 897 25974 901
rect 17343 638 17953 643
rect 17493 634 17948 638
rect 8772 457 9322 462
rect 8883 453 9317 457
<< via2 >>
rect 15692 44122 15748 44178
rect 5392 43532 5448 43588
rect 6862 43392 6918 43448
rect 8332 43252 8388 43308
rect 9802 42922 9858 42978
rect 11272 42922 11328 42978
rect 12742 42932 12798 42988
rect 14212 42922 14268 42978
rect 17162 43982 17218 44038
rect 18632 43852 18688 43908
rect 20112 43712 20168 43768
rect 21582 43572 21638 43628
rect 23052 43422 23108 43478
rect 24522 43292 24578 43348
rect 25992 43162 26048 43218
rect 27460 43034 27516 43090
rect 28938 42900 28994 42956
rect 30514 42770 30570 42826
rect 22325 9435 22615 9725
rect 6125 8985 6415 9275
rect 14375 9125 14665 9415
rect 12895 7785 13185 8075
rect 21145 7795 21435 8085
rect 29135 7785 29425 8075
rect 8883 462 9317 896
rect 17493 643 17948 1098
rect 25566 906 25974 1314
<< metal3 >>
rect 16246 44778 16252 44842
rect 16316 44778 16322 44842
rect 16982 44778 16988 44842
rect 17052 44778 17058 44842
rect 17718 44778 17724 44842
rect 17788 44778 17794 44842
rect 15687 44180 15753 44183
rect 15838 44182 15902 44188
rect 15687 44178 15838 44180
rect 15687 44122 15692 44178
rect 15748 44122 15838 44178
rect 15687 44120 15838 44122
rect 15687 44117 15753 44120
rect 15838 44112 15902 44118
rect 5387 43590 5453 43593
rect 16254 43590 16314 44778
rect 5387 43588 16314 43590
rect 5387 43532 5392 43588
rect 5448 43532 16314 43588
rect 5387 43530 16314 43532
rect 5387 43527 5453 43530
rect 6857 43450 6923 43453
rect 16990 43450 17050 44778
rect 17157 44040 17223 44043
rect 17318 44042 17382 44048
rect 17157 44038 17318 44040
rect 17157 43982 17162 44038
rect 17218 43982 17318 44038
rect 17157 43980 17318 43982
rect 17157 43977 17223 43980
rect 17318 43972 17382 43978
rect 6857 43448 17050 43450
rect 6857 43392 6862 43448
rect 6918 43392 17050 43448
rect 6857 43390 17050 43392
rect 6857 43387 6923 43390
rect 8327 43310 8393 43313
rect 17726 43310 17786 44778
rect 18627 43910 18693 43913
rect 18808 43912 18872 43918
rect 18627 43908 18808 43910
rect 18627 43852 18632 43908
rect 18688 43852 18808 43908
rect 18627 43850 18808 43852
rect 18627 43847 18693 43850
rect 18808 43842 18872 43848
rect 20107 43770 20173 43773
rect 20298 43772 20362 43778
rect 20107 43768 20298 43770
rect 20107 43712 20112 43768
rect 20168 43712 20298 43768
rect 20107 43710 20298 43712
rect 20107 43707 20173 43710
rect 20298 43702 20362 43708
rect 21577 43630 21643 43633
rect 21738 43632 21802 43638
rect 21577 43628 21738 43630
rect 21577 43572 21582 43628
rect 21638 43572 21738 43628
rect 21577 43570 21738 43572
rect 21577 43567 21643 43570
rect 21738 43562 21802 43568
rect 23047 43480 23113 43483
rect 23208 43482 23272 43488
rect 23047 43478 23208 43480
rect 23047 43422 23052 43478
rect 23108 43422 23208 43478
rect 23047 43420 23208 43422
rect 23047 43417 23113 43420
rect 23208 43412 23272 43418
rect 8327 43308 17786 43310
rect 8327 43252 8332 43308
rect 8388 43252 17786 43308
rect 24517 43350 24583 43353
rect 24678 43352 24742 43358
rect 24517 43348 24678 43350
rect 24517 43292 24522 43348
rect 24578 43292 24678 43348
rect 24517 43290 24678 43292
rect 24517 43287 24583 43290
rect 24678 43282 24742 43288
rect 8327 43250 17786 43252
rect 8327 43247 8393 43250
rect 25987 43220 26053 43223
rect 26168 43222 26232 43228
rect 25987 43218 26168 43220
rect 11268 43172 11332 43178
rect 9792 43108 9798 43172
rect 9862 43108 9868 43172
rect 9800 42983 9860 43108
rect 11268 43102 11332 43108
rect 12738 43172 12802 43178
rect 25987 43162 25992 43218
rect 26048 43162 26168 43218
rect 25987 43160 26168 43162
rect 25987 43157 26053 43160
rect 26168 43152 26232 43158
rect 12738 43102 12802 43108
rect 11270 42983 11330 43102
rect 12740 42993 12800 43102
rect 27455 43092 27521 43095
rect 27712 43094 27776 43100
rect 27455 43090 27712 43092
rect 27455 43034 27460 43090
rect 27516 43034 27712 43090
rect 27455 43032 27712 43034
rect 27455 43029 27521 43032
rect 27712 43024 27776 43030
rect 12737 42988 12803 42993
rect 9797 42978 9863 42983
rect 9797 42922 9802 42978
rect 9858 42922 9863 42978
rect 9797 42917 9863 42922
rect 11267 42978 11333 42983
rect 11267 42922 11272 42978
rect 11328 42922 11333 42978
rect 12737 42932 12742 42988
rect 12798 42932 12803 42988
rect 14210 42983 14270 42990
rect 12737 42927 12803 42932
rect 14207 42980 14273 42983
rect 14388 42982 14452 42988
rect 14207 42978 14388 42980
rect 11267 42917 11333 42922
rect 14207 42922 14212 42978
rect 14268 42922 14388 42978
rect 14207 42920 14388 42922
rect 14207 42917 14273 42920
rect 14388 42912 14452 42918
rect 28933 42958 28999 42961
rect 29174 42960 29238 42966
rect 28933 42956 29174 42958
rect 28933 42900 28938 42956
rect 28994 42900 29174 42956
rect 28933 42898 29174 42900
rect 28933 42895 28999 42898
rect 29174 42890 29238 42896
rect 30509 42828 30575 42831
rect 30700 42830 30764 42836
rect 30509 42826 30700 42828
rect 30509 42770 30514 42826
rect 30570 42770 30700 42826
rect 30509 42768 30700 42770
rect 30509 42765 30575 42768
rect 30700 42760 30764 42766
rect 7750 10796 8050 10802
rect 21196 10782 21496 10788
rect 5391 9280 5689 9285
rect 5390 9279 6420 9280
rect 5390 8981 5391 9279
rect 5689 9275 6420 9279
rect 5689 8985 6125 9275
rect 6415 8985 6420 9275
rect 5689 8981 6420 8985
rect 5390 8980 6420 8981
rect 5391 8975 5689 8980
rect 1001 8080 1299 8085
rect 7750 8080 8050 10496
rect 14456 10482 14462 10782
rect 14762 10482 15594 10782
rect 13660 9419 14670 9420
rect 13655 9121 13661 9419
rect 13959 9415 14670 9419
rect 13959 9125 14375 9415
rect 14665 9125 14670 9415
rect 13959 9121 14670 9125
rect 13660 9120 14670 9121
rect 15294 8080 15594 10482
rect 21196 8090 21496 10482
rect 27896 10782 28196 10788
rect 21831 9730 22129 9735
rect 21830 9729 22620 9730
rect 21830 9431 21831 9729
rect 22129 9725 22620 9729
rect 22129 9435 22325 9725
rect 22615 9435 22620 9725
rect 22129 9431 22620 9435
rect 21830 9430 22620 9431
rect 21831 9425 22129 9430
rect 21110 8085 21510 8090
rect 21110 8080 21145 8085
rect 1000 8079 21145 8080
rect 1000 7781 1001 8079
rect 1299 8075 21145 8079
rect 1299 7785 12895 8075
rect 13185 7795 21145 8075
rect 21435 8080 21510 8085
rect 27896 8080 28196 10482
rect 21435 8075 29480 8080
rect 21435 7795 29135 8075
rect 13185 7785 29135 7795
rect 29425 7785 29480 8075
rect 1299 7781 29480 7785
rect 1000 7780 29480 7781
rect 1001 7775 1299 7780
rect 25561 1314 26689 1319
rect 17488 1098 18733 1103
rect 8878 896 10302 901
rect 8878 462 8883 896
rect 9317 834 10302 896
rect 10447 834 10754 839
rect 9317 833 10755 834
rect 9317 526 10447 833
rect 10754 526 10755 833
rect 17488 643 17493 1098
rect 17948 1019 18733 1098
rect 20542 1019 20838 1024
rect 17948 1018 20839 1019
rect 17948 722 20542 1018
rect 20838 722 20839 1018
rect 25561 906 25566 1314
rect 25974 1261 26689 1314
rect 29890 1261 30190 1266
rect 25974 1260 30191 1261
rect 25974 960 29890 1260
rect 30190 960 30191 1260
rect 25974 959 30191 960
rect 25974 906 26689 959
rect 29890 954 30190 959
rect 25561 901 26689 906
rect 17948 721 20839 722
rect 17948 643 18733 721
rect 20542 716 20838 721
rect 17488 638 18733 643
rect 9317 525 10755 526
rect 9317 462 10302 525
rect 10447 520 10754 525
rect 8878 457 10302 462
<< via3 >>
rect 16252 44778 16316 44842
rect 16988 44778 17052 44842
rect 17724 44778 17788 44842
rect 15838 44118 15902 44182
rect 17318 43978 17382 44042
rect 18808 43848 18872 43912
rect 20298 43708 20362 43772
rect 21738 43568 21802 43632
rect 23208 43418 23272 43482
rect 24678 43288 24742 43352
rect 9798 43108 9862 43172
rect 11268 43108 11332 43172
rect 12738 43108 12802 43172
rect 26168 43158 26232 43222
rect 27712 43030 27776 43094
rect 14388 42918 14452 42982
rect 29174 42896 29238 42960
rect 30700 42766 30764 42830
rect 7750 10496 8050 10796
rect 5391 8981 5689 9279
rect 14462 10482 14762 10782
rect 13661 9121 13959 9419
rect 21196 10482 21496 10782
rect 27896 10482 28196 10782
rect 21831 9431 22129 9729
rect 1001 7781 1299 8079
rect 10447 526 10754 833
rect 20542 722 20838 1018
rect 29890 960 30190 1260
<< metal4 >>
rect 798 44900 858 45152
rect 790 44800 870 44900
rect 1534 44800 1594 45152
rect 2270 44800 2330 45152
rect 3006 44800 3066 45152
rect 3742 44800 3802 45152
rect 4478 44800 4538 45152
rect 5214 44800 5274 45152
rect 5950 44800 6010 45152
rect 6686 44800 6746 45152
rect 7422 44800 7482 45152
rect 8158 44800 8218 45152
rect 8894 44800 8954 45152
rect 9630 44800 9690 45152
rect 10366 44800 10426 45152
rect 11102 44800 11162 45152
rect 11838 44800 11898 45152
rect 12574 44800 12634 45152
rect 13310 44800 13370 45152
rect 14046 44800 14106 45152
rect 14782 44800 14842 45152
rect 15518 44800 15578 45152
rect 16254 44843 16314 45152
rect 16990 44843 17050 45152
rect 17726 44843 17786 45152
rect 18462 44860 18522 45152
rect 19198 44860 19258 45152
rect 19934 44860 19994 45152
rect 20670 44860 20730 45152
rect 790 44740 15578 44800
rect 16251 44842 16317 44843
rect 16251 44778 16252 44842
rect 16316 44778 16317 44842
rect 16251 44777 16317 44778
rect 16987 44842 17053 44843
rect 16987 44778 16988 44842
rect 17052 44778 17053 44842
rect 16987 44777 17053 44778
rect 17723 44842 17789 44843
rect 17723 44778 17724 44842
rect 17788 44778 17789 44842
rect 17723 44777 17789 44778
rect 790 44720 14840 44740
rect 1530 44500 14840 44720
rect 21406 44680 21466 45152
rect 15030 44620 21466 44680
rect 200 8080 500 44152
rect 1800 9730 2100 44500
rect 15030 43840 15090 44620
rect 22142 44560 22202 45152
rect 9800 43780 15090 43840
rect 15190 44500 22202 44560
rect 9800 43173 9860 43780
rect 15190 43710 15250 44500
rect 22878 44440 22938 45152
rect 11270 43650 15250 43710
rect 15350 44380 22938 44440
rect 11270 43173 11330 43650
rect 12740 43173 12800 43180
rect 9797 43172 9863 43173
rect 9797 43108 9798 43172
rect 9862 43108 9863 43172
rect 9797 43107 9863 43108
rect 11267 43172 11333 43173
rect 11267 43108 11268 43172
rect 11332 43108 11333 43172
rect 11267 43107 11333 43108
rect 12737 43172 12803 43173
rect 12737 43108 12738 43172
rect 12802 43170 12803 43172
rect 14050 43170 14110 43180
rect 15350 43170 15410 44380
rect 23614 44310 23674 45152
rect 15520 44250 23674 44310
rect 15520 43170 15580 44250
rect 15837 44182 15903 44183
rect 15837 44118 15838 44182
rect 15902 44180 15903 44182
rect 24350 44180 24410 45152
rect 15902 44120 24410 44180
rect 15902 44118 15903 44120
rect 15837 44117 15903 44118
rect 17317 44042 17383 44043
rect 17317 43978 17318 44042
rect 17382 44040 17383 44042
rect 25086 44040 25146 45152
rect 17382 43980 25146 44040
rect 17382 43978 17383 43980
rect 17317 43977 17383 43978
rect 18807 43912 18873 43913
rect 18807 43848 18808 43912
rect 18872 43910 18873 43912
rect 25822 43910 25882 45152
rect 18872 43850 25882 43910
rect 18872 43848 18873 43850
rect 18807 43847 18873 43848
rect 20297 43772 20363 43773
rect 20297 43708 20298 43772
rect 20362 43770 20363 43772
rect 26558 43770 26618 45152
rect 20362 43710 26618 43770
rect 20362 43708 20363 43710
rect 20297 43707 20363 43708
rect 21737 43632 21803 43633
rect 21737 43568 21738 43632
rect 21802 43630 21803 43632
rect 27294 43630 27354 45152
rect 21802 43570 27354 43630
rect 21802 43568 21803 43570
rect 21737 43567 21803 43568
rect 23207 43482 23273 43483
rect 23207 43418 23208 43482
rect 23272 43480 23273 43482
rect 28030 43480 28090 45152
rect 23272 43420 28090 43480
rect 23272 43418 23273 43420
rect 23207 43417 23273 43418
rect 24677 43352 24743 43353
rect 24677 43288 24678 43352
rect 24742 43350 24743 43352
rect 28766 43350 28826 45152
rect 24742 43290 28826 43350
rect 24742 43288 24743 43290
rect 24677 43287 24743 43288
rect 12802 43110 15410 43170
rect 15510 43110 15580 43170
rect 26167 43222 26233 43223
rect 26167 43158 26168 43222
rect 26232 43220 26233 43222
rect 29502 43220 29562 45152
rect 26232 43160 29562 43220
rect 26232 43158 26233 43160
rect 26167 43157 26233 43158
rect 12802 43108 12803 43110
rect 12737 43107 12803 43108
rect 14387 42982 14453 42983
rect 14387 42918 14388 42982
rect 14452 42980 14453 42982
rect 15520 42980 15580 43110
rect 27711 43094 27777 43095
rect 27711 43030 27712 43094
rect 27776 43092 27777 43094
rect 30238 43092 30298 45152
rect 27776 43032 30298 43092
rect 27776 43030 27777 43032
rect 27711 43029 27777 43030
rect 14452 42920 15580 42980
rect 29173 42960 29239 42961
rect 14452 42918 14453 42920
rect 14387 42917 14453 42918
rect 29173 42896 29174 42960
rect 29238 42958 29239 42960
rect 30974 42958 31034 45152
rect 29238 42898 31034 42958
rect 29238 42896 29239 42898
rect 29173 42895 29239 42896
rect 30699 42830 30765 42831
rect 30699 42766 30700 42830
rect 30764 42828 30765 42830
rect 31710 42828 31770 45152
rect 30764 42768 31770 42828
rect 30764 42766 30765 42768
rect 30699 42765 30765 42766
rect 7750 10797 8050 41900
rect 7749 10796 8051 10797
rect 7749 10496 7750 10796
rect 8050 10496 8051 10796
rect 7749 10495 8051 10496
rect 11098 9730 11398 41878
rect 14462 10783 14762 41822
rect 14461 10782 14763 10783
rect 14461 10482 14462 10782
rect 14762 10482 14763 10782
rect 14461 10481 14763 10482
rect 17826 9730 18126 41900
rect 21196 10783 21496 41850
rect 21195 10782 21497 10783
rect 21195 10482 21196 10782
rect 21496 10482 21497 10782
rect 21195 10481 21497 10482
rect 24554 9730 24854 41894
rect 27896 10783 28196 41906
rect 27895 10782 28197 10783
rect 27895 10482 27896 10782
rect 28196 10482 28197 10782
rect 27895 10481 28197 10482
rect 31250 9730 31550 41888
rect 1800 9729 31550 9730
rect 1800 9431 21831 9729
rect 22129 9431 31550 9729
rect 1800 9430 31550 9431
rect 200 8079 1300 8080
rect 200 7781 1001 8079
rect 1299 7781 1300 8079
rect 200 7780 1300 7781
rect 200 1000 500 7780
rect 1800 1000 2100 9430
rect 5390 9279 5690 9430
rect 5390 8981 5391 9279
rect 5689 8981 5690 9279
rect 13660 9419 13960 9430
rect 13660 9121 13661 9419
rect 13959 9121 13960 9419
rect 13660 9120 13960 9121
rect 5390 8980 5690 8981
rect 29889 1260 31460 1261
rect 21630 1019 21970 1020
rect 20541 1018 21970 1019
rect 12176 834 12894 835
rect 10446 833 12894 834
rect 10446 526 10447 833
rect 10754 526 12894 833
rect 20541 722 20542 1018
rect 20838 780 21970 1018
rect 29889 960 29890 1260
rect 30190 960 31462 1260
rect 29889 959 31462 960
rect 20838 722 27046 780
rect 20541 721 27046 722
rect 21620 600 27046 721
rect 10446 525 12894 526
rect 12585 456 12894 525
rect 12585 286 22630 456
rect 12640 276 22630 286
rect 370 0 550 200
rect 4786 0 4966 200
rect 9202 0 9382 200
rect 13618 0 13798 200
rect 18034 0 18214 200
rect 22450 0 22630 276
rect 26866 0 27046 600
rect 31282 0 31462 959
use ay8913  ay8913_0
timestamp 1717176801
transform 1 0 3988 0 1 10844
box 514 0 27576 32000
use dac_16nfet  dac_16nfet_0
timestamp 1716419193
transform 0 -1 22676 -1 0 10400
box -11 -6800 9500 406
use dac_16nfet  dac_16nfet_1
timestamp 1716419193
transform 0 -1 14700 -1 0 10120
box -11 -6800 9500 406
use dac_16nfet  dac_16nfet_2
timestamp 1716419193
transform 0 -1 6456 -1 0 9952
box -11 -6800 9500 406
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31282 0 31462 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26866 0 27046 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22450 0 22630 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18034 0 18214 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13618 0 13798 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9202 0 9382 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4786 0 4966 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 370 0 550 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 4800 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 1800 1000 2100 44152 1 FreeSans 4800 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
