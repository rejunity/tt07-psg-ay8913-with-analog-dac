VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_rejunity_ay8913
  CLASS BLOCK ;
  FOREIGN tt_um_rejunity_ay8913 ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 13.148600 ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 13.148600 ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 13.148600 ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1172.472900 ;
    ANTENNADIFFAREA 999.351990 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1172.472900 ;
    ANTENNADIFFAREA 999.351990 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1172.472900 ;
    ANTENNADIFFAREA 999.351990 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1172.472900 ;
    ANTENNADIFFAREA 999.351990 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1172.472900 ;
    ANTENNADIFFAREA 999.351990 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1172.472900 ;
    ANTENNADIFFAREA 999.351990 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1172.472900 ;
    ANTENNADIFFAREA 999.351990 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1172.472900 ;
    ANTENNADIFFAREA 999.351990 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1172.472900 ;
    ANTENNADIFFAREA 999.351990 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1172.472900 ;
    ANTENNADIFFAREA 999.351990 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1172.472900 ;
    ANTENNADIFFAREA 999.351990 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1172.472900 ;
    ANTENNADIFFAREA 999.351990 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1172.472900 ;
    ANTENNADIFFAREA 999.351990 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1172.472900 ;
    ANTENNADIFFAREA 999.351990 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1172.472900 ;
    ANTENNADIFFAREA 999.351990 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1172.472900 ;
    ANTENNADIFFAREA 999.351990 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1172.472900 ;
    ANTENNADIFFAREA 999.351990 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1172.472900 ;
    ANTENNADIFFAREA 999.351990 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1172.472900 ;
    ANTENNADIFFAREA 999.351990 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1172.472900 ;
    ANTENNADIFFAREA 999.351990 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1172.472900 ;
    ANTENNADIFFAREA 999.351990 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 9.000 5.000 10.500 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 22.845 209.155 23.015 209.345 ;
        RECT 24.225 209.155 24.395 209.345 ;
        RECT 29.745 209.155 29.915 209.345 ;
        RECT 35.260 209.205 35.380 209.315 ;
        RECT 36.185 209.155 36.355 209.345 ;
        RECT 41.705 209.155 41.875 209.345 ;
        RECT 47.225 209.155 47.395 209.345 ;
        RECT 22.705 208.345 24.075 209.155 ;
        RECT 24.085 208.345 29.595 209.155 ;
        RECT 29.605 208.345 35.115 209.155 ;
        RECT 35.595 208.285 36.025 209.070 ;
        RECT 36.045 208.345 41.555 209.155 ;
        RECT 41.565 208.345 47.075 209.155 ;
        RECT 47.085 208.345 48.455 209.155 ;
        RECT 49.070 209.125 49.240 209.345 ;
        RECT 51.820 209.155 51.990 209.345 ;
        RECT 55.965 209.155 56.135 209.345 ;
        RECT 56.435 209.200 56.595 209.310 ;
        RECT 60.565 209.155 60.735 209.345 ;
        RECT 61.020 209.205 61.140 209.315 ;
        RECT 62.865 209.155 63.035 209.345 ;
        RECT 63.335 209.200 63.495 209.310 ;
        RECT 64.245 209.155 64.415 209.345 ;
        RECT 65.625 209.155 65.795 209.345 ;
        RECT 69.300 209.205 69.420 209.315 ;
        RECT 71.605 209.155 71.775 209.345 ;
        RECT 72.065 209.155 72.235 209.345 ;
        RECT 73.455 209.200 73.615 209.310 ;
        RECT 74.825 209.155 74.995 209.345 ;
        RECT 78.500 209.205 78.620 209.315 ;
        RECT 78.965 209.155 79.135 209.345 ;
        RECT 80.800 209.155 80.970 209.345 ;
        RECT 82.180 209.205 82.300 209.315 ;
        RECT 85.865 209.155 86.035 209.345 ;
        RECT 86.335 209.200 86.495 209.310 ;
        RECT 91.390 209.155 91.560 209.345 ;
        RECT 91.845 209.155 92.015 209.345 ;
        RECT 93.685 209.155 93.855 209.345 ;
        RECT 95.525 209.155 95.695 209.345 ;
        RECT 99.215 209.200 99.375 209.310 ;
        RECT 50.730 209.125 51.675 209.155 ;
        RECT 48.475 208.285 48.905 209.070 ;
        RECT 48.925 208.445 51.675 209.125 ;
        RECT 50.730 208.245 51.675 208.445 ;
        RECT 51.705 208.245 53.055 209.155 ;
        RECT 53.065 208.245 56.175 209.155 ;
        RECT 57.300 208.475 60.765 209.155 ;
        RECT 57.300 208.245 58.220 208.475 ;
        RECT 61.355 208.285 61.785 209.070 ;
        RECT 61.805 208.375 63.175 209.155 ;
        RECT 64.105 208.375 65.475 209.155 ;
        RECT 65.485 208.345 69.155 209.155 ;
        RECT 69.625 208.475 71.915 209.155 ;
        RECT 69.625 208.245 70.545 208.475 ;
        RECT 71.925 208.375 73.295 209.155 ;
        RECT 74.235 208.285 74.665 209.070 ;
        RECT 74.685 208.345 78.355 209.155 ;
        RECT 78.825 208.475 80.655 209.155 ;
        RECT 79.310 208.245 80.655 208.475 ;
        RECT 80.685 208.245 82.035 209.155 ;
        RECT 82.600 208.475 86.065 209.155 ;
        RECT 82.600 208.245 83.520 208.475 ;
        RECT 87.115 208.285 87.545 209.070 ;
        RECT 87.565 208.245 91.670 209.155 ;
        RECT 91.705 208.345 93.535 209.155 ;
        RECT 93.545 208.475 95.375 209.155 ;
        RECT 94.030 208.245 95.375 208.475 ;
        RECT 95.385 208.345 99.055 209.155 ;
        RECT 100.445 209.125 101.390 209.155 ;
        RECT 103.345 209.125 103.515 209.345 ;
        RECT 103.805 209.155 103.975 209.345 ;
        RECT 105.185 209.155 105.355 209.345 ;
        RECT 107.020 209.205 107.140 209.315 ;
        RECT 110.245 209.155 110.415 209.345 ;
        RECT 112.085 209.155 112.255 209.345 ;
        RECT 112.540 209.205 112.660 209.315 ;
        RECT 113.465 209.155 113.635 209.345 ;
        RECT 116.695 209.200 116.855 209.310 ;
        RECT 120.825 209.155 120.995 209.345 ;
        RECT 122.665 209.155 122.835 209.345 ;
        RECT 124.505 209.155 124.675 209.345 ;
        RECT 124.975 209.200 125.135 209.310 ;
        RECT 126.345 209.155 126.515 209.345 ;
        RECT 130.020 209.205 130.140 209.315 ;
        RECT 131.865 209.155 132.035 209.345 ;
        RECT 132.325 209.155 132.495 209.345 ;
        RECT 134.625 209.155 134.795 209.345 ;
        RECT 135.085 209.155 135.255 209.345 ;
        RECT 139.200 209.175 139.370 209.345 ;
        RECT 139.260 209.155 139.370 209.175 ;
        RECT 143.825 209.155 143.995 209.345 ;
        RECT 149.345 209.155 149.515 209.345 ;
        RECT 151.180 209.205 151.300 209.315 ;
        RECT 152.100 209.205 152.220 209.315 ;
        RECT 153.485 209.155 153.655 209.345 ;
        RECT 153.945 209.155 154.115 209.345 ;
        RECT 156.705 209.155 156.875 209.345 ;
        RECT 99.995 208.285 100.425 209.070 ;
        RECT 100.445 208.925 103.515 209.125 ;
        RECT 100.445 208.445 103.655 208.925 ;
        RECT 100.445 208.245 101.390 208.445 ;
        RECT 102.725 208.245 103.655 208.445 ;
        RECT 103.665 208.375 105.035 209.155 ;
        RECT 105.045 208.345 106.875 209.155 ;
        RECT 107.345 208.245 110.555 209.155 ;
        RECT 110.565 208.475 112.395 209.155 ;
        RECT 112.875 208.285 113.305 209.070 ;
        RECT 113.325 208.245 116.535 209.155 ;
        RECT 117.560 208.475 121.025 209.155 ;
        RECT 121.145 208.475 122.975 209.155 ;
        RECT 122.985 208.475 124.815 209.155 ;
        RECT 117.560 208.245 118.480 208.475 ;
        RECT 125.755 208.285 126.185 209.070 ;
        RECT 126.205 208.345 129.875 209.155 ;
        RECT 130.345 208.475 132.175 209.155 ;
        RECT 132.185 208.345 133.555 209.155 ;
        RECT 133.565 208.375 134.935 209.155 ;
        RECT 134.945 208.345 138.615 209.155 ;
        RECT 138.635 208.285 139.065 209.070 ;
        RECT 139.260 208.475 143.675 209.155 ;
        RECT 139.745 208.245 143.675 208.475 ;
        RECT 143.685 208.345 149.195 209.155 ;
        RECT 149.205 208.345 151.035 209.155 ;
        RECT 151.515 208.285 151.945 209.070 ;
        RECT 152.425 208.375 153.795 209.155 ;
        RECT 153.805 208.345 155.635 209.155 ;
        RECT 155.645 208.345 157.015 209.155 ;
      LAYER nwell ;
        RECT 22.510 205.125 157.210 207.955 ;
      LAYER pwell ;
        RECT 22.705 203.925 24.075 204.735 ;
        RECT 24.085 203.925 27.755 204.735 ;
        RECT 27.845 204.605 29.615 204.835 ;
        RECT 31.150 204.605 32.060 204.825 ;
        RECT 27.845 203.925 35.575 204.605 ;
        RECT 35.595 204.010 36.025 204.795 ;
        RECT 39.560 204.605 40.470 204.825 ;
        RECT 42.005 204.605 43.775 204.835 ;
        RECT 47.380 204.605 48.290 204.825 ;
        RECT 49.825 204.605 51.175 204.835 ;
        RECT 36.045 203.925 43.775 204.605 ;
        RECT 43.865 203.925 51.175 204.605 ;
        RECT 51.685 203.925 53.055 204.705 ;
        RECT 56.580 204.605 57.490 204.825 ;
        RECT 59.025 204.605 60.375 204.835 ;
        RECT 53.065 203.925 60.375 204.605 ;
        RECT 61.355 204.010 61.785 204.795 ;
        RECT 61.825 203.925 63.175 204.835 ;
        RECT 63.185 203.925 64.555 204.705 ;
        RECT 64.575 203.925 65.925 204.835 ;
        RECT 65.945 203.925 67.315 204.705 ;
        RECT 70.840 204.605 71.750 204.825 ;
        RECT 73.285 204.605 74.635 204.835 ;
        RECT 67.325 203.925 74.635 204.605 ;
        RECT 75.165 203.925 76.515 204.835 ;
        RECT 80.040 204.605 80.950 204.825 ;
        RECT 82.485 204.605 83.835 204.835 ;
        RECT 76.525 203.925 83.835 204.605 ;
        RECT 83.885 203.925 85.255 204.735 ;
        RECT 85.750 204.605 87.095 204.835 ;
        RECT 85.265 203.925 87.095 204.605 ;
        RECT 87.115 204.010 87.545 204.795 ;
        RECT 87.565 203.925 88.935 204.705 ;
        RECT 89.445 204.605 90.795 204.835 ;
        RECT 92.330 204.605 93.240 204.825 ;
        RECT 89.445 203.925 96.755 204.605 ;
        RECT 96.765 203.925 98.135 204.705 ;
        RECT 98.605 203.925 99.975 204.705 ;
        RECT 100.025 204.605 101.375 204.835 ;
        RECT 102.910 204.605 103.820 204.825 ;
        RECT 100.025 203.925 107.335 204.605 ;
        RECT 107.345 203.925 109.175 204.735 ;
        RECT 109.280 204.605 110.200 204.835 ;
        RECT 109.280 203.925 112.745 204.605 ;
        RECT 112.875 204.010 113.305 204.795 ;
        RECT 117.760 204.605 118.670 204.825 ;
        RECT 120.205 204.605 121.555 204.835 ;
        RECT 114.245 203.925 121.555 204.605 ;
        RECT 121.645 203.925 124.815 204.835 ;
        RECT 124.825 204.605 125.755 204.835 ;
        RECT 129.405 204.605 130.335 204.835 ;
        RECT 134.780 204.605 135.690 204.825 ;
        RECT 137.225 204.605 138.575 204.835 ;
        RECT 124.825 203.925 127.575 204.605 ;
        RECT 127.585 203.925 130.335 204.605 ;
        RECT 131.265 203.925 138.575 204.605 ;
        RECT 138.635 204.010 139.065 204.795 ;
        RECT 139.085 203.925 140.455 204.705 ;
        RECT 140.505 204.605 141.855 204.835 ;
        RECT 143.390 204.605 144.300 204.825 ;
        RECT 140.505 203.925 147.815 204.605 ;
        RECT 147.825 203.925 153.335 204.735 ;
        RECT 153.345 203.925 155.175 204.735 ;
        RECT 155.645 203.925 157.015 204.735 ;
        RECT 22.845 203.715 23.015 203.925 ;
        RECT 24.225 203.735 24.395 203.925 ;
        RECT 31.585 203.715 31.755 203.905 ;
        RECT 32.055 203.760 32.215 203.870 ;
        RECT 32.965 203.755 33.135 203.905 ;
        RECT 22.705 202.905 24.075 203.715 ;
        RECT 24.165 203.035 31.895 203.715 ;
        RECT 24.165 202.805 25.935 203.035 ;
        RECT 27.470 202.815 28.380 203.035 ;
        RECT 32.845 202.805 33.735 203.755 ;
        RECT 33.885 203.715 34.055 203.905 ;
        RECT 35.265 203.735 35.435 203.925 ;
        RECT 36.185 203.735 36.355 203.925 ;
        RECT 37.565 203.715 37.735 203.905 ;
        RECT 39.870 203.715 40.040 203.905 ;
        RECT 40.320 203.765 40.440 203.875 ;
        RECT 40.785 203.715 40.955 203.905 ;
        RECT 44.005 203.735 44.175 203.925 ;
        RECT 46.765 203.715 46.935 203.905 ;
        RECT 47.225 203.715 47.395 203.905 ;
        RECT 51.360 203.765 51.480 203.875 ;
        RECT 52.745 203.735 52.915 203.925 ;
        RECT 53.205 203.735 53.375 203.925 ;
        RECT 56.420 203.715 56.590 203.905 ;
        RECT 56.885 203.715 57.055 203.905 ;
        RECT 59.640 203.765 59.760 203.875 ;
        RECT 60.105 203.715 60.275 203.905 ;
        RECT 60.575 203.770 60.735 203.880 ;
        RECT 61.940 203.735 62.110 203.925 ;
        RECT 64.245 203.735 64.415 203.925 ;
        RECT 65.625 203.735 65.795 203.925 ;
        RECT 66.085 203.735 66.255 203.925 ;
        RECT 67.465 203.715 67.635 203.925 ;
        RECT 70.220 203.765 70.340 203.875 ;
        RECT 72.525 203.735 72.695 203.905 ;
        RECT 72.525 203.715 72.690 203.735 ;
        RECT 73.910 203.715 74.080 203.905 ;
        RECT 74.825 203.875 74.995 203.905 ;
        RECT 74.820 203.765 74.995 203.875 ;
        RECT 74.825 203.715 74.995 203.765 ;
        RECT 75.280 203.735 75.450 203.925 ;
        RECT 76.665 203.755 76.835 203.925 ;
        RECT 77.135 203.760 77.295 203.870 ;
        RECT 33.745 202.905 37.415 203.715 ;
        RECT 37.425 202.905 38.795 203.715 ;
        RECT 38.805 202.805 40.155 203.715 ;
        RECT 40.645 202.935 42.015 203.715 ;
        RECT 42.260 203.035 47.075 203.715 ;
        RECT 47.085 202.905 48.455 203.715 ;
        RECT 48.475 202.845 48.905 203.630 ;
        RECT 48.985 202.805 56.735 203.715 ;
        RECT 56.745 202.905 59.495 203.715 ;
        RECT 59.965 203.035 67.275 203.715 ;
        RECT 63.480 202.815 64.390 203.035 ;
        RECT 65.925 202.805 67.275 203.035 ;
        RECT 67.325 202.905 70.075 203.715 ;
        RECT 70.855 203.035 72.690 203.715 ;
        RECT 70.855 202.805 71.785 203.035 ;
        RECT 72.845 202.805 74.195 203.715 ;
        RECT 74.235 202.845 74.665 203.630 ;
        RECT 74.685 202.905 76.055 203.715 ;
        RECT 76.065 202.805 76.955 203.755 ;
        RECT 78.050 203.715 78.220 203.905 ;
        RECT 82.185 203.715 82.355 203.905 ;
        RECT 83.565 203.715 83.735 203.905 ;
        RECT 84.025 203.735 84.195 203.925 ;
        RECT 85.405 203.735 85.575 203.925 ;
        RECT 88.625 203.735 88.795 203.925 ;
        RECT 89.080 203.765 89.200 203.875 ;
        RECT 90.935 203.760 91.095 203.870 ;
        RECT 91.845 203.735 92.015 203.905 ;
        RECT 91.850 203.715 92.015 203.735 ;
        RECT 77.905 203.035 82.035 203.715 ;
        RECT 80.645 202.805 82.035 203.035 ;
        RECT 82.045 202.905 83.415 203.715 ;
        RECT 83.425 203.035 90.735 203.715 ;
        RECT 91.850 203.035 93.685 203.715 ;
        RECT 94.150 203.685 94.320 203.905 ;
        RECT 96.445 203.735 96.615 203.925 ;
        RECT 97.825 203.735 97.995 203.925 ;
        RECT 98.280 203.765 98.400 203.875 ;
        RECT 98.745 203.735 98.915 203.925 ;
        RECT 99.205 203.735 99.375 203.905 ;
        RECT 99.660 203.765 99.780 203.875 ;
        RECT 99.205 203.715 99.355 203.735 ;
        RECT 96.280 203.685 97.215 203.715 ;
        RECT 94.150 203.485 97.215 203.685 ;
        RECT 86.940 202.815 87.850 203.035 ;
        RECT 89.385 202.805 90.735 203.035 ;
        RECT 92.755 202.805 93.685 203.035 ;
        RECT 94.005 203.005 97.215 203.485 ;
        RECT 94.005 202.805 94.935 203.005 ;
        RECT 96.265 202.805 97.215 203.005 ;
        RECT 97.425 202.895 99.355 203.715 ;
        RECT 100.445 203.685 101.380 203.715 ;
        RECT 103.340 203.685 103.510 203.905 ;
        RECT 103.805 203.715 103.975 203.905 ;
        RECT 106.565 203.715 106.735 203.905 ;
        RECT 107.025 203.735 107.195 203.925 ;
        RECT 107.485 203.735 107.655 203.925 ;
        RECT 112.545 203.735 112.715 203.925 ;
        RECT 113.475 203.770 113.635 203.880 ;
        RECT 113.925 203.715 114.095 203.905 ;
        RECT 114.385 203.735 114.555 203.925 ;
        RECT 121.745 203.735 121.915 203.925 ;
        RECT 124.505 203.715 124.675 203.905 ;
        RECT 124.975 203.760 125.135 203.870 ;
        RECT 127.265 203.735 127.435 203.925 ;
        RECT 127.725 203.735 127.895 203.925 ;
        RECT 128.645 203.735 128.815 203.905 ;
        RECT 128.645 203.715 128.775 203.735 ;
        RECT 97.425 202.805 98.375 202.895 ;
        RECT 99.995 202.845 100.425 203.630 ;
        RECT 100.445 203.485 103.510 203.685 ;
        RECT 100.445 203.005 103.655 203.485 ;
        RECT 103.665 203.035 106.405 203.715 ;
        RECT 106.425 203.035 113.735 203.715 ;
        RECT 113.785 203.035 121.095 203.715 ;
        RECT 100.445 202.805 101.395 203.005 ;
        RECT 102.725 202.805 103.655 203.005 ;
        RECT 109.940 202.815 110.850 203.035 ;
        RECT 112.385 202.805 113.735 203.035 ;
        RECT 117.300 202.815 118.210 203.035 ;
        RECT 119.745 202.805 121.095 203.035 ;
        RECT 121.240 203.035 124.705 203.715 ;
        RECT 121.240 202.805 122.160 203.035 ;
        RECT 125.755 202.845 126.185 203.630 ;
        RECT 126.925 203.485 128.775 203.715 ;
        RECT 129.100 203.685 129.270 203.905 ;
        RECT 130.495 203.770 130.655 203.880 ;
        RECT 131.405 203.715 131.575 203.925 ;
        RECT 130.300 203.685 131.255 203.715 ;
        RECT 126.440 202.805 128.775 203.485 ;
        RECT 128.975 203.005 131.255 203.685 ;
        RECT 131.265 203.035 134.475 203.715 ;
        RECT 130.300 202.805 131.255 203.005 ;
        RECT 133.340 202.805 134.475 203.035 ;
        RECT 134.485 203.685 135.420 203.715 ;
        RECT 137.380 203.685 137.550 203.905 ;
        RECT 134.485 203.485 137.550 203.685 ;
        RECT 137.850 203.685 138.020 203.905 ;
        RECT 139.225 203.735 139.395 203.925 ;
        RECT 141.065 203.715 141.235 203.905 ;
        RECT 142.905 203.715 143.075 203.905 ;
        RECT 146.125 203.715 146.295 203.905 ;
        RECT 147.505 203.735 147.675 203.925 ;
        RECT 147.965 203.735 148.135 203.925 ;
        RECT 153.485 203.735 153.655 203.925 ;
        RECT 155.325 203.875 155.495 203.905 ;
        RECT 155.320 203.765 155.495 203.875 ;
        RECT 155.325 203.715 155.495 203.765 ;
        RECT 156.705 203.715 156.875 203.925 ;
        RECT 139.980 203.685 140.915 203.715 ;
        RECT 137.850 203.485 140.915 203.685 ;
        RECT 134.485 203.005 137.695 203.485 ;
        RECT 134.485 202.805 135.435 203.005 ;
        RECT 136.765 202.805 137.695 203.005 ;
        RECT 137.705 203.005 140.915 203.485 ;
        RECT 137.705 202.805 138.635 203.005 ;
        RECT 139.965 202.805 140.915 203.005 ;
        RECT 140.925 202.905 142.755 203.715 ;
        RECT 142.865 202.805 145.975 203.715 ;
        RECT 145.985 202.905 151.495 203.715 ;
        RECT 151.515 202.845 151.945 203.630 ;
        RECT 152.060 203.035 155.525 203.715 ;
        RECT 152.060 202.805 152.980 203.035 ;
        RECT 155.645 202.905 157.015 203.715 ;
      LAYER nwell ;
        RECT 22.510 199.685 157.210 202.515 ;
      LAYER pwell ;
        RECT 22.705 198.485 24.075 199.295 ;
        RECT 24.085 198.485 29.595 199.295 ;
        RECT 29.605 198.485 35.115 199.295 ;
        RECT 35.595 198.570 36.025 199.355 ;
        RECT 36.045 198.485 37.415 199.295 ;
        RECT 40.940 199.165 41.850 199.385 ;
        RECT 43.385 199.165 44.735 199.395 ;
        RECT 37.425 198.485 44.735 199.165 ;
        RECT 44.795 198.485 47.525 199.395 ;
        RECT 49.365 199.165 50.295 199.395 ;
        RECT 47.545 198.485 50.295 199.165 ;
        RECT 50.305 198.485 52.135 199.395 ;
        RECT 52.145 198.485 57.655 199.295 ;
        RECT 57.665 198.485 61.335 199.295 ;
        RECT 61.355 198.570 61.785 199.355 ;
        RECT 61.805 199.195 62.755 199.395 ;
        RECT 64.085 199.195 65.015 199.395 ;
        RECT 61.805 198.715 65.015 199.195 ;
        RECT 61.805 198.515 64.870 198.715 ;
        RECT 61.805 198.485 62.740 198.515 ;
        RECT 22.845 198.275 23.015 198.485 ;
        RECT 24.225 198.275 24.395 198.485 ;
        RECT 29.745 198.275 29.915 198.485 ;
        RECT 35.260 198.325 35.380 198.435 ;
        RECT 36.185 198.295 36.355 198.485 ;
        RECT 37.565 198.295 37.735 198.485 ;
        RECT 39.405 198.275 39.575 198.465 ;
        RECT 39.865 198.275 40.035 198.465 ;
        RECT 41.700 198.325 41.820 198.435 ;
        RECT 44.005 198.275 44.175 198.465 ;
        RECT 44.465 198.275 44.635 198.465 ;
        RECT 44.925 198.295 45.095 198.485 ;
        RECT 47.685 198.295 47.855 198.485 ;
        RECT 51.820 198.465 51.990 198.485 ;
        RECT 48.140 198.325 48.260 198.435 ;
        RECT 51.820 198.295 51.995 198.465 ;
        RECT 51.825 198.275 51.995 198.295 ;
        RECT 52.285 198.275 52.455 198.485 ;
        RECT 57.805 198.295 57.975 198.485 ;
        RECT 64.700 198.465 64.870 198.515 ;
        RECT 65.025 198.485 66.375 199.395 ;
        RECT 66.865 198.485 68.235 199.265 ;
        RECT 68.245 198.485 70.075 199.295 ;
        RECT 70.105 198.485 71.455 199.395 ;
        RECT 71.465 198.485 74.215 199.295 ;
        RECT 75.735 199.165 76.665 199.395 ;
        RECT 74.830 198.485 76.665 199.165 ;
        RECT 77.000 198.485 78.815 199.395 ;
        RECT 78.825 198.485 84.335 199.295 ;
        RECT 85.855 199.165 86.785 199.395 ;
        RECT 84.950 198.485 86.785 199.165 ;
        RECT 87.115 198.570 87.545 199.355 ;
        RECT 87.565 198.485 93.075 199.295 ;
        RECT 93.085 198.485 95.835 199.295 ;
        RECT 97.355 199.165 98.285 199.395 ;
        RECT 96.450 198.485 98.285 199.165 ;
        RECT 98.605 198.485 100.435 199.295 ;
        RECT 101.815 199.165 102.735 199.395 ;
        RECT 100.445 198.485 102.735 199.165 ;
        RECT 102.765 198.485 104.115 199.395 ;
        RECT 104.125 198.485 105.495 199.265 ;
        RECT 105.505 198.485 111.015 199.295 ;
        RECT 111.025 198.485 112.855 199.295 ;
        RECT 112.875 198.570 113.305 199.355 ;
        RECT 113.325 198.485 116.535 199.395 ;
        RECT 116.545 198.485 120.215 199.295 ;
        RECT 122.030 199.195 122.975 199.395 ;
        RECT 120.225 198.515 122.975 199.195 ;
        RECT 61.485 198.275 61.655 198.465 ;
        RECT 63.320 198.275 63.490 198.465 ;
        RECT 63.795 198.320 63.955 198.430 ;
        RECT 64.700 198.295 64.875 198.465 ;
        RECT 65.170 198.295 65.340 198.485 ;
        RECT 66.540 198.325 66.660 198.435 ;
        RECT 67.925 198.295 68.095 198.485 ;
        RECT 68.385 198.295 68.555 198.485 ;
        RECT 70.220 198.295 70.390 198.485 ;
        RECT 71.605 198.295 71.775 198.485 ;
        RECT 74.830 198.465 74.995 198.485 ;
        RECT 64.705 198.275 64.875 198.295 ;
        RECT 72.980 198.275 73.150 198.465 ;
        RECT 73.455 198.320 73.615 198.430 ;
        RECT 74.360 198.325 74.480 198.435 ;
        RECT 74.825 198.275 74.995 198.465 ;
        RECT 22.705 197.465 24.075 198.275 ;
        RECT 24.085 197.465 29.595 198.275 ;
        RECT 29.605 197.465 32.355 198.275 ;
        RECT 32.405 197.595 39.715 198.275 ;
        RECT 32.405 197.365 33.755 197.595 ;
        RECT 35.290 197.375 36.200 197.595 ;
        RECT 39.725 197.465 41.555 198.275 ;
        RECT 42.025 197.595 44.315 198.275 ;
        RECT 42.025 197.365 42.945 197.595 ;
        RECT 44.325 197.465 47.995 198.275 ;
        RECT 48.475 197.405 48.905 198.190 ;
        RECT 48.925 197.365 52.035 198.275 ;
        RECT 52.145 197.595 59.455 198.275 ;
        RECT 55.660 197.375 56.570 197.595 ;
        RECT 58.105 197.365 59.455 197.595 ;
        RECT 59.505 197.595 61.795 198.275 ;
        RECT 59.505 197.365 60.425 197.595 ;
        RECT 61.805 197.365 63.635 198.275 ;
        RECT 64.565 197.595 71.875 198.275 ;
        RECT 68.080 197.375 68.990 197.595 ;
        RECT 70.525 197.365 71.875 197.595 ;
        RECT 71.945 197.365 73.295 198.275 ;
        RECT 74.235 197.405 74.665 198.190 ;
        RECT 74.695 197.365 76.045 198.275 ;
        RECT 76.210 198.245 76.380 198.465 ;
        RECT 77.125 198.295 77.295 198.485 ;
        RECT 78.965 198.295 79.135 198.485 ;
        RECT 84.950 198.465 85.115 198.485 ;
        RECT 79.425 198.275 79.595 198.465 ;
        RECT 83.105 198.275 83.275 198.465 ;
        RECT 84.490 198.435 84.660 198.465 ;
        RECT 84.480 198.325 84.660 198.435 ;
        RECT 78.340 198.245 79.275 198.275 ;
        RECT 76.210 198.045 79.275 198.245 ;
        RECT 76.065 197.565 79.275 198.045 ;
        RECT 76.065 197.365 76.995 197.565 ;
        RECT 78.325 197.365 79.275 197.565 ;
        RECT 79.285 197.465 82.955 198.275 ;
        RECT 82.965 197.465 84.335 198.275 ;
        RECT 84.490 198.245 84.660 198.325 ;
        RECT 84.945 198.295 85.115 198.465 ;
        RECT 87.705 198.275 87.875 198.485 ;
        RECT 86.620 198.245 87.555 198.275 ;
        RECT 84.490 198.045 87.555 198.245 ;
        RECT 84.345 197.565 87.555 198.045 ;
        RECT 84.345 197.365 85.275 197.565 ;
        RECT 86.605 197.365 87.555 197.565 ;
        RECT 87.565 197.465 88.935 198.275 ;
        RECT 89.090 198.245 89.260 198.465 ;
        RECT 92.305 198.295 92.475 198.465 ;
        RECT 93.225 198.295 93.395 198.485 ;
        RECT 96.450 198.465 96.615 198.485 ;
        RECT 94.600 198.325 94.720 198.435 ;
        RECT 92.310 198.275 92.475 198.295 ;
        RECT 95.065 198.275 95.235 198.465 ;
        RECT 95.980 198.325 96.100 198.435 ;
        RECT 96.445 198.295 96.615 198.465 ;
        RECT 97.365 198.275 97.535 198.465 ;
        RECT 98.745 198.295 98.915 198.485 ;
        RECT 99.215 198.320 99.375 198.430 ;
        RECT 100.585 198.295 100.755 198.485 ;
        RECT 102.880 198.430 103.050 198.485 ;
        RECT 102.880 198.320 103.055 198.430 ;
        RECT 102.880 198.295 103.050 198.320 ;
        RECT 100.590 198.275 100.755 198.295 ;
        RECT 103.805 198.275 103.975 198.465 ;
        RECT 104.265 198.295 104.435 198.485 ;
        RECT 105.645 198.295 105.815 198.485 ;
        RECT 111.165 198.295 111.335 198.485 ;
        RECT 112.085 198.275 112.255 198.465 ;
        RECT 112.555 198.320 112.715 198.430 ;
        RECT 113.465 198.275 113.635 198.465 ;
        RECT 116.225 198.295 116.395 198.485 ;
        RECT 116.685 198.295 116.855 198.485 ;
        RECT 120.370 198.295 120.540 198.515 ;
        RECT 122.030 198.485 122.975 198.515 ;
        RECT 122.985 198.485 125.735 199.295 ;
        RECT 127.540 199.195 128.495 199.395 ;
        RECT 126.215 198.515 128.495 199.195 ;
        RECT 123.125 198.295 123.295 198.485 ;
        RECT 124.045 198.275 124.215 198.465 ;
        RECT 124.505 198.275 124.675 198.465 ;
        RECT 125.880 198.325 126.000 198.435 ;
        RECT 126.340 198.295 126.510 198.515 ;
        RECT 127.540 198.485 128.495 198.515 ;
        RECT 128.505 198.485 131.255 199.295 ;
        RECT 133.095 199.165 134.015 199.395 ;
        RECT 131.725 198.485 134.015 199.165 ;
        RECT 134.035 198.485 135.385 199.395 ;
        RECT 135.415 198.485 138.145 199.395 ;
        RECT 138.635 198.570 139.065 199.355 ;
        RECT 143.520 199.165 144.430 199.385 ;
        RECT 145.965 199.165 147.315 199.395 ;
        RECT 150.880 199.165 151.790 199.385 ;
        RECT 153.325 199.165 154.675 199.395 ;
        RECT 140.005 198.485 147.315 199.165 ;
        RECT 147.365 198.485 154.675 199.165 ;
        RECT 155.645 198.485 157.015 199.295 ;
        RECT 128.645 198.295 128.815 198.485 ;
        RECT 130.945 198.275 131.115 198.465 ;
        RECT 131.400 198.325 131.520 198.435 ;
        RECT 131.865 198.295 132.035 198.485 ;
        RECT 133.245 198.295 133.415 198.465 ;
        RECT 133.245 198.275 133.395 198.295 ;
        RECT 133.705 198.275 133.875 198.465 ;
        RECT 135.085 198.295 135.255 198.485 ;
        RECT 135.545 198.295 135.715 198.485 ;
        RECT 136.460 198.325 136.580 198.435 ;
        RECT 136.925 198.295 137.095 198.465 ;
        RECT 138.300 198.325 138.420 198.435 ;
        RECT 139.235 198.320 139.395 198.440 ;
        RECT 136.930 198.275 137.095 198.295 ;
        RECT 140.145 198.275 140.315 198.485 ;
        RECT 141.525 198.275 141.695 198.465 ;
        RECT 147.040 198.275 147.210 198.465 ;
        RECT 147.505 198.295 147.675 198.485 ;
        RECT 148.425 198.275 148.595 198.465 ;
        RECT 151.180 198.325 151.300 198.435 ;
        RECT 152.105 198.275 152.275 198.465 ;
        RECT 154.875 198.330 155.035 198.440 ;
        RECT 156.705 198.275 156.875 198.485 ;
        RECT 91.220 198.245 92.155 198.275 ;
        RECT 89.090 198.045 92.155 198.245 ;
        RECT 88.945 197.565 92.155 198.045 ;
        RECT 92.310 197.595 94.145 198.275 ;
        RECT 94.925 197.595 97.215 198.275 ;
        RECT 97.225 197.595 99.055 198.275 ;
        RECT 88.945 197.365 89.875 197.565 ;
        RECT 91.205 197.365 92.155 197.565 ;
        RECT 93.215 197.365 94.145 197.595 ;
        RECT 96.295 197.365 97.215 197.595 ;
        RECT 99.995 197.405 100.425 198.190 ;
        RECT 100.590 197.595 102.425 198.275 ;
        RECT 103.665 197.595 110.975 198.275 ;
        RECT 101.495 197.365 102.425 197.595 ;
        RECT 107.180 197.375 108.090 197.595 ;
        RECT 109.625 197.365 110.975 197.595 ;
        RECT 111.035 197.365 112.385 198.275 ;
        RECT 113.325 197.595 120.635 198.275 ;
        RECT 116.840 197.375 117.750 197.595 ;
        RECT 119.285 197.365 120.635 197.595 ;
        RECT 120.780 197.595 124.245 198.275 ;
        RECT 120.780 197.365 121.700 197.595 ;
        RECT 124.365 197.465 125.735 198.275 ;
        RECT 125.755 197.405 126.185 198.190 ;
        RECT 126.440 197.595 131.255 198.275 ;
        RECT 131.465 197.455 133.395 198.275 ;
        RECT 133.565 197.465 136.315 198.275 ;
        RECT 136.930 197.595 138.765 198.275 ;
        RECT 131.465 197.365 132.415 197.455 ;
        RECT 137.835 197.365 138.765 197.595 ;
        RECT 140.005 197.495 141.375 198.275 ;
        RECT 141.385 197.465 146.895 198.275 ;
        RECT 146.925 197.365 148.275 198.275 ;
        RECT 148.285 197.465 151.035 198.275 ;
        RECT 151.515 197.405 151.945 198.190 ;
        RECT 151.965 197.465 155.635 198.275 ;
        RECT 155.645 197.465 157.015 198.275 ;
      LAYER nwell ;
        RECT 22.510 194.245 157.210 197.075 ;
      LAYER pwell ;
        RECT 22.705 193.045 24.075 193.855 ;
        RECT 24.085 193.045 29.595 193.855 ;
        RECT 29.605 193.045 32.355 193.855 ;
        RECT 33.135 193.725 34.065 193.955 ;
        RECT 33.135 193.045 34.970 193.725 ;
        RECT 35.595 193.130 36.025 193.915 ;
        RECT 36.045 193.045 37.415 193.825 ;
        RECT 37.425 193.045 39.255 193.855 ;
        RECT 39.265 193.045 40.635 193.825 ;
        RECT 40.645 193.045 46.155 193.855 ;
        RECT 46.165 193.045 47.535 193.855 ;
        RECT 47.555 193.045 48.905 193.955 ;
        RECT 50.730 193.755 51.675 193.955 ;
        RECT 48.925 193.075 51.675 193.755 ;
        RECT 22.845 192.835 23.015 193.045 ;
        RECT 24.225 192.835 24.395 193.045 ;
        RECT 27.915 192.880 28.075 192.990 ;
        RECT 28.825 192.835 28.995 193.025 ;
        RECT 29.745 192.855 29.915 193.045 ;
        RECT 34.805 193.025 34.970 193.045 ;
        RECT 30.675 192.880 30.835 192.990 ;
        RECT 22.705 192.025 24.075 192.835 ;
        RECT 24.085 192.025 27.755 192.835 ;
        RECT 28.685 192.155 30.515 192.835 ;
        RECT 31.590 192.805 31.760 193.025 ;
        RECT 32.500 192.885 32.620 192.995 ;
        RECT 34.805 192.855 34.975 193.025 ;
        RECT 35.260 192.885 35.380 192.995 ;
        RECT 36.185 192.855 36.355 193.045 ;
        RECT 36.645 192.855 36.815 193.025 ;
        RECT 37.100 192.885 37.220 192.995 ;
        RECT 36.645 192.835 36.795 192.855 ;
        RECT 37.565 192.835 37.735 193.045 ;
        RECT 40.325 192.855 40.495 193.045 ;
        RECT 40.785 192.855 40.955 193.045 ;
        RECT 44.920 192.885 45.040 192.995 ;
        RECT 45.385 192.835 45.555 193.025 ;
        RECT 46.305 192.855 46.475 193.045 ;
        RECT 47.685 192.855 47.855 193.045 ;
        RECT 49.070 192.855 49.240 193.075 ;
        RECT 50.730 193.045 51.675 193.075 ;
        RECT 51.685 193.045 54.425 193.725 ;
        RECT 54.445 193.045 55.815 193.825 ;
        RECT 55.825 193.045 57.655 193.855 ;
        RECT 58.135 193.045 60.865 193.955 ;
        RECT 61.355 193.130 61.785 193.915 ;
        RECT 61.805 193.045 64.555 193.855 ;
        RECT 69.625 193.755 70.575 193.955 ;
        RECT 71.905 193.755 72.835 193.955 ;
        RECT 64.565 193.045 69.380 193.725 ;
        RECT 69.625 193.275 72.835 193.755 ;
        RECT 72.845 193.725 73.980 193.955 ;
        RECT 80.040 193.725 80.950 193.945 ;
        RECT 82.485 193.725 83.835 193.955 ;
        RECT 69.625 193.075 72.690 193.275 ;
        RECT 69.625 193.045 70.560 193.075 ;
        RECT 51.365 192.835 51.535 193.025 ;
        RECT 51.825 192.855 51.995 193.045 ;
        RECT 55.505 192.855 55.675 193.045 ;
        RECT 55.965 192.855 56.135 193.045 ;
        RECT 57.800 192.885 57.920 192.995 ;
        RECT 58.725 192.835 58.895 193.025 ;
        RECT 59.185 192.835 59.355 193.025 ;
        RECT 60.565 192.855 60.735 193.045 ;
        RECT 61.020 192.885 61.140 192.995 ;
        RECT 61.945 192.855 62.115 193.045 ;
        RECT 62.865 192.835 63.035 193.025 ;
        RECT 64.705 192.855 64.875 193.045 ;
        RECT 67.925 192.835 68.095 193.025 ;
        RECT 68.385 192.835 68.555 193.025 ;
        RECT 72.060 192.885 72.180 192.995 ;
        RECT 72.520 192.855 72.690 193.075 ;
        RECT 72.845 193.045 76.055 193.725 ;
        RECT 76.525 193.045 83.835 193.725 ;
        RECT 85.005 193.865 85.955 193.955 ;
        RECT 85.005 193.045 86.935 193.865 ;
        RECT 87.115 193.130 87.545 193.915 ;
        RECT 88.935 193.725 89.855 193.955 ;
        RECT 87.565 193.045 89.855 193.725 ;
        RECT 89.905 193.725 91.255 193.955 ;
        RECT 92.790 193.725 93.700 193.945 ;
        RECT 100.340 193.725 101.260 193.955 ;
        RECT 104.880 193.725 105.790 193.945 ;
        RECT 107.325 193.725 108.675 193.955 ;
        RECT 111.380 193.725 112.300 193.955 ;
        RECT 89.905 193.045 97.215 193.725 ;
        RECT 97.795 193.045 101.260 193.725 ;
        RECT 101.365 193.045 108.675 193.725 ;
        RECT 108.835 193.045 112.300 193.725 ;
        RECT 112.875 193.130 113.305 193.915 ;
        RECT 113.325 193.045 116.535 193.955 ;
        RECT 116.545 193.045 120.215 193.855 ;
        RECT 122.490 193.755 123.435 193.955 ;
        RECT 120.685 193.075 123.435 193.755 ;
        RECT 73.445 192.835 73.615 193.025 ;
        RECT 73.900 192.885 74.020 192.995 ;
        RECT 74.825 192.835 74.995 193.025 ;
        RECT 75.745 192.855 75.915 193.045 ;
        RECT 76.200 192.885 76.320 192.995 ;
        RECT 76.665 192.855 76.835 193.045 ;
        RECT 86.785 193.025 86.935 193.045 ;
        RECT 77.580 192.885 77.700 192.995 ;
        RECT 78.965 192.835 79.135 193.025 ;
        RECT 80.345 192.835 80.515 193.025 ;
        RECT 80.805 192.835 80.975 193.025 ;
        RECT 84.035 192.890 84.195 193.000 ;
        RECT 84.480 192.885 84.600 192.995 ;
        RECT 85.865 192.835 86.035 193.025 ;
        RECT 86.325 192.835 86.495 193.025 ;
        RECT 86.785 192.855 86.955 193.025 ;
        RECT 87.705 192.855 87.875 193.045 ;
        RECT 88.625 192.835 88.795 193.025 ;
        RECT 89.085 192.835 89.255 193.025 ;
        RECT 90.920 192.885 91.040 192.995 ;
        RECT 91.385 192.835 91.555 193.025 ;
        RECT 92.775 192.880 92.935 192.990 ;
        RECT 94.605 192.835 94.775 193.025 ;
        RECT 95.065 192.835 95.235 193.025 ;
        RECT 96.905 192.995 97.075 193.045 ;
        RECT 96.900 192.885 97.075 192.995 ;
        RECT 97.360 192.885 97.480 192.995 ;
        RECT 96.905 192.855 97.075 192.885 ;
        RECT 97.825 192.855 97.995 193.045 ;
        RECT 98.285 192.835 98.455 193.025 ;
        RECT 98.745 192.835 98.915 193.025 ;
        RECT 100.585 192.855 100.755 193.025 ;
        RECT 101.505 192.855 101.675 193.045 ;
        RECT 103.355 192.880 103.515 192.990 ;
        RECT 100.735 192.835 100.755 192.855 ;
        RECT 108.865 192.835 109.035 193.045 ;
        RECT 109.325 192.835 109.495 193.025 ;
        RECT 112.540 192.885 112.660 192.995 ;
        RECT 116.225 192.855 116.395 193.045 ;
        RECT 116.685 192.835 116.855 193.045 ;
        RECT 120.360 192.885 120.480 192.995 ;
        RECT 120.830 192.855 121.000 193.075 ;
        RECT 122.490 193.045 123.435 193.075 ;
        RECT 123.905 193.045 125.720 193.955 ;
        RECT 126.235 193.045 128.955 193.955 ;
        RECT 128.965 193.045 130.795 193.855 ;
        RECT 130.805 193.045 132.155 193.955 ;
        RECT 132.185 193.045 134.935 193.855 ;
        RECT 134.945 193.045 136.295 193.955 ;
        RECT 137.375 193.725 138.305 193.955 ;
        RECT 136.470 193.045 138.305 193.725 ;
        RECT 138.635 193.130 139.065 193.915 ;
        RECT 139.085 193.725 140.005 193.955 ;
        RECT 141.385 193.725 142.305 193.955 ;
        RECT 139.085 193.045 141.375 193.725 ;
        RECT 141.385 193.045 143.675 193.725 ;
        RECT 143.685 193.045 145.515 193.855 ;
        RECT 145.525 193.045 146.895 193.825 ;
        RECT 146.905 193.045 152.415 193.855 ;
        RECT 152.425 193.045 155.175 193.855 ;
        RECT 155.645 193.045 157.015 193.855 ;
        RECT 123.580 192.885 123.700 192.995 ;
        RECT 124.045 192.835 124.215 193.025 ;
        RECT 125.425 192.855 125.595 193.045 ;
        RECT 125.880 192.885 126.000 192.995 ;
        RECT 126.340 192.885 126.460 192.995 ;
        RECT 128.185 192.835 128.355 193.025 ;
        RECT 128.645 192.855 128.815 193.045 ;
        RECT 129.105 192.855 129.275 193.045 ;
        RECT 130.950 192.855 131.120 193.045 ;
        RECT 33.720 192.805 34.655 192.835 ;
        RECT 31.590 192.605 34.655 192.805 ;
        RECT 31.445 192.125 34.655 192.605 ;
        RECT 31.445 191.925 32.375 192.125 ;
        RECT 33.705 191.925 34.655 192.125 ;
        RECT 34.865 192.015 36.795 192.835 ;
        RECT 37.425 192.155 44.735 192.835 ;
        RECT 45.245 192.155 48.455 192.835 ;
        RECT 34.865 191.925 35.815 192.015 ;
        RECT 40.940 191.935 41.850 192.155 ;
        RECT 43.385 191.925 44.735 192.155 ;
        RECT 47.320 191.925 48.455 192.155 ;
        RECT 48.475 191.965 48.905 192.750 ;
        RECT 48.955 191.925 51.675 192.835 ;
        RECT 51.725 192.155 59.035 192.835 ;
        RECT 51.725 191.925 53.075 192.155 ;
        RECT 54.610 191.935 55.520 192.155 ;
        RECT 59.045 192.025 62.715 192.835 ;
        RECT 62.725 192.155 65.475 192.835 ;
        RECT 64.545 191.925 65.475 192.155 ;
        RECT 65.485 192.155 68.235 192.835 ;
        RECT 65.485 191.925 66.415 192.155 ;
        RECT 68.245 192.025 71.915 192.835 ;
        RECT 72.395 191.925 73.745 192.835 ;
        RECT 74.235 191.965 74.665 192.750 ;
        RECT 74.685 192.025 77.435 192.835 ;
        RECT 77.905 192.055 79.275 192.835 ;
        RECT 79.295 191.925 80.645 192.835 ;
        RECT 80.665 192.025 84.335 192.835 ;
        RECT 84.815 191.925 86.165 192.835 ;
        RECT 86.185 192.025 87.555 192.835 ;
        RECT 87.575 191.925 88.925 192.835 ;
        RECT 88.945 192.025 90.775 192.835 ;
        RECT 91.245 192.055 92.615 192.835 ;
        RECT 93.555 191.925 94.905 192.835 ;
        RECT 94.925 192.025 96.755 192.835 ;
        RECT 97.235 191.925 98.585 192.835 ;
        RECT 98.605 192.025 99.975 192.835 ;
        RECT 99.995 191.965 100.425 192.750 ;
        RECT 100.735 192.155 103.185 192.835 ;
        RECT 104.360 192.155 109.175 192.835 ;
        RECT 109.185 192.155 116.495 192.835 ;
        RECT 116.545 192.155 123.855 192.835 ;
        RECT 101.225 191.925 103.185 192.155 ;
        RECT 112.700 191.935 113.610 192.155 ;
        RECT 115.145 191.925 116.495 192.155 ;
        RECT 120.060 191.935 120.970 192.155 ;
        RECT 122.505 191.925 123.855 192.155 ;
        RECT 123.905 192.025 125.735 192.835 ;
        RECT 125.755 191.965 126.185 192.750 ;
        RECT 126.665 191.925 128.480 192.835 ;
        RECT 128.505 192.805 129.455 192.835 ;
        RECT 131.860 192.805 132.030 193.025 ;
        RECT 132.325 192.855 132.495 193.045 ;
        RECT 135.085 192.835 135.255 193.025 ;
        RECT 135.545 192.835 135.715 193.025 ;
        RECT 136.010 192.855 136.180 193.045 ;
        RECT 136.470 193.025 136.635 193.045 ;
        RECT 141.065 193.025 141.235 193.045 ;
        RECT 136.465 192.855 136.635 193.025 ;
        RECT 137.850 192.835 138.020 193.025 ;
        RECT 139.225 192.835 139.395 193.025 ;
        RECT 139.685 192.835 139.855 193.025 ;
        RECT 141.065 192.855 141.240 193.025 ;
        RECT 143.365 192.855 143.535 193.045 ;
        RECT 143.825 192.855 143.995 193.045 ;
        RECT 145.665 192.855 145.835 193.045 ;
        RECT 147.045 192.855 147.215 193.045 ;
        RECT 128.505 192.125 132.175 192.805 ;
        RECT 128.505 191.925 129.455 192.125 ;
        RECT 132.185 191.925 135.395 192.835 ;
        RECT 135.405 192.025 136.775 192.835 ;
        RECT 136.785 191.925 138.135 192.835 ;
        RECT 138.175 191.925 139.525 192.835 ;
        RECT 139.545 192.025 140.915 192.835 ;
        RECT 141.070 192.805 141.240 192.855 ;
        RECT 151.185 192.835 151.355 193.025 ;
        RECT 152.105 192.835 152.275 193.025 ;
        RECT 152.565 192.855 152.735 193.045 ;
        RECT 155.320 192.885 155.440 192.995 ;
        RECT 156.705 192.835 156.875 193.045 ;
        RECT 143.200 192.805 144.135 192.835 ;
        RECT 141.070 192.605 144.135 192.805 ;
        RECT 140.925 192.125 144.135 192.605 ;
        RECT 140.925 191.925 141.855 192.125 ;
        RECT 143.185 191.925 144.135 192.125 ;
        RECT 144.185 192.155 151.495 192.835 ;
        RECT 144.185 191.925 145.535 192.155 ;
        RECT 147.070 191.935 147.980 192.155 ;
        RECT 151.515 191.965 151.945 192.750 ;
        RECT 151.965 192.025 155.635 192.835 ;
        RECT 155.645 192.025 157.015 192.835 ;
      LAYER nwell ;
        RECT 22.510 188.805 157.210 191.635 ;
      LAYER pwell ;
        RECT 22.705 187.605 24.075 188.415 ;
        RECT 27.600 188.285 28.510 188.505 ;
        RECT 30.045 188.285 31.395 188.515 ;
        RECT 24.085 187.605 31.395 188.285 ;
        RECT 31.445 188.315 32.395 188.515 ;
        RECT 33.725 188.315 34.655 188.515 ;
        RECT 31.445 187.835 34.655 188.315 ;
        RECT 31.445 187.635 34.510 187.835 ;
        RECT 35.595 187.690 36.025 188.475 ;
        RECT 31.445 187.605 32.380 187.635 ;
        RECT 22.845 187.395 23.015 187.605 ;
        RECT 24.225 187.395 24.395 187.605 ;
        RECT 26.525 187.395 26.695 187.585 ;
        RECT 26.985 187.395 27.155 187.585 ;
        RECT 30.675 187.440 30.835 187.550 ;
        RECT 33.425 187.395 33.595 187.585 ;
        RECT 34.340 187.415 34.510 187.635 ;
        RECT 36.045 187.605 37.875 188.415 ;
        RECT 37.885 188.315 38.815 188.515 ;
        RECT 40.145 188.315 41.095 188.515 ;
        RECT 37.885 187.835 41.095 188.315 ;
        RECT 38.030 187.635 41.095 187.835 ;
        RECT 34.815 187.450 34.975 187.560 ;
        RECT 35.725 187.415 35.895 187.585 ;
        RECT 35.725 187.395 35.890 187.415 ;
        RECT 36.185 187.395 36.355 187.605 ;
        RECT 37.565 187.395 37.735 187.585 ;
        RECT 38.030 187.415 38.200 187.635 ;
        RECT 40.160 187.605 41.095 187.635 ;
        RECT 41.105 187.605 42.475 188.415 ;
        RECT 42.485 187.605 45.405 188.515 ;
        RECT 45.705 187.605 47.535 188.415 ;
        RECT 48.005 188.315 48.950 188.515 ;
        RECT 48.005 187.635 50.755 188.315 ;
        RECT 48.005 187.605 48.950 187.635 ;
        RECT 39.400 187.445 39.520 187.555 ;
        RECT 39.865 187.395 40.035 187.585 ;
        RECT 41.245 187.415 41.415 187.605 ;
        RECT 42.630 187.585 42.800 187.605 ;
        RECT 42.625 187.415 42.800 187.585 ;
        RECT 45.380 187.445 45.500 187.555 ;
        RECT 42.625 187.395 42.795 187.415 ;
        RECT 45.845 187.395 46.015 187.605 ;
        RECT 47.680 187.445 47.800 187.555 ;
        RECT 50.440 187.415 50.610 187.635 ;
        RECT 50.765 187.605 53.975 188.515 ;
        RECT 56.640 188.285 57.560 188.515 ;
        RECT 54.095 187.605 57.560 188.285 ;
        RECT 57.760 188.285 58.680 188.515 ;
        RECT 57.760 187.605 61.225 188.285 ;
        RECT 61.355 187.690 61.785 188.475 ;
        RECT 64.070 188.315 65.015 188.515 ;
        RECT 62.265 187.635 65.015 188.315 ;
        RECT 50.905 187.415 51.075 187.605 ;
        RECT 51.835 187.395 52.005 187.585 ;
        RECT 52.295 187.440 52.455 187.550 ;
        RECT 53.205 187.395 53.375 187.585 ;
        RECT 54.125 187.415 54.295 187.605 ;
        RECT 60.565 187.395 60.735 187.585 ;
        RECT 61.025 187.415 61.195 187.605 ;
        RECT 61.945 187.555 62.115 187.585 ;
        RECT 61.940 187.445 62.115 187.555 ;
        RECT 61.945 187.395 62.115 187.445 ;
        RECT 62.410 187.415 62.580 187.635 ;
        RECT 64.070 187.605 65.015 187.635 ;
        RECT 65.025 187.605 68.680 188.515 ;
        RECT 68.715 187.605 71.445 188.515 ;
        RECT 71.465 187.605 74.675 188.515 ;
        RECT 74.685 187.605 76.055 188.415 ;
        RECT 76.065 187.605 79.275 188.515 ;
        RECT 79.745 187.605 82.955 188.515 ;
        RECT 83.425 187.605 86.635 188.515 ;
        RECT 87.115 187.690 87.545 188.475 ;
        RECT 87.565 187.605 90.775 188.515 ;
        RECT 91.245 187.605 93.060 188.515 ;
        RECT 93.085 187.605 96.295 188.515 ;
        RECT 96.765 187.605 99.975 188.515 ;
        RECT 99.985 187.605 105.495 188.415 ;
        RECT 105.965 187.605 109.175 188.515 ;
        RECT 109.645 187.605 112.855 188.515 ;
        RECT 112.875 187.690 113.305 188.475 ;
        RECT 113.420 188.285 114.340 188.515 ;
        RECT 113.420 187.605 116.885 188.285 ;
        RECT 117.005 187.605 118.835 188.415 ;
        RECT 118.940 188.285 119.860 188.515 ;
        RECT 118.940 187.605 122.405 188.285 ;
        RECT 122.525 187.605 124.355 188.415 ;
        RECT 124.385 187.605 125.735 188.515 ;
        RECT 127.550 188.315 128.495 188.515 ;
        RECT 125.745 187.635 128.495 188.315 ;
        RECT 64.245 187.395 64.415 187.585 ;
        RECT 65.170 187.415 65.340 187.605 ;
        RECT 67.015 187.440 67.175 187.550 ;
        RECT 71.145 187.395 71.315 187.605 ;
        RECT 71.600 187.445 71.720 187.555 ;
        RECT 73.905 187.395 74.075 187.585 ;
        RECT 74.365 187.415 74.535 187.605 ;
        RECT 74.825 187.395 74.995 187.605 ;
        RECT 76.205 187.415 76.375 187.605 ;
        RECT 78.965 187.395 79.135 187.585 ;
        RECT 79.425 187.555 79.595 187.585 ;
        RECT 79.420 187.445 79.595 187.555 ;
        RECT 79.425 187.395 79.595 187.445 ;
        RECT 79.885 187.415 80.055 187.605 ;
        RECT 82.185 187.395 82.355 187.585 ;
        RECT 83.100 187.445 83.220 187.555 ;
        RECT 83.565 187.415 83.735 187.605 ;
        RECT 85.865 187.395 86.035 187.585 ;
        RECT 86.325 187.395 86.495 187.585 ;
        RECT 86.780 187.445 86.900 187.555 ;
        RECT 90.465 187.415 90.635 187.605 ;
        RECT 90.920 187.445 91.040 187.555 ;
        RECT 91.845 187.395 92.015 187.585 ;
        RECT 92.765 187.415 92.935 187.605 ;
        RECT 93.225 187.415 93.395 187.605 ;
        RECT 96.440 187.445 96.560 187.555 ;
        RECT 96.895 187.415 97.065 187.605 ;
        RECT 97.375 187.440 97.535 187.550 ;
        RECT 98.290 187.395 98.460 187.585 ;
        RECT 100.125 187.415 100.295 187.605 ;
        RECT 100.580 187.395 100.750 187.585 ;
        RECT 105.640 187.445 105.760 187.555 ;
        RECT 106.105 187.415 106.275 187.605 ;
        RECT 22.705 186.585 24.075 187.395 ;
        RECT 24.085 186.585 25.455 187.395 ;
        RECT 25.465 186.615 26.835 187.395 ;
        RECT 26.845 186.585 30.515 187.395 ;
        RECT 31.445 186.715 33.735 187.395 ;
        RECT 34.055 186.715 35.890 187.395 ;
        RECT 31.445 186.485 32.365 186.715 ;
        RECT 34.055 186.485 34.985 186.715 ;
        RECT 36.055 186.485 37.405 187.395 ;
        RECT 37.425 186.585 39.255 187.395 ;
        RECT 39.725 186.715 42.475 187.395 ;
        RECT 41.545 186.485 42.475 186.715 ;
        RECT 42.485 186.585 45.235 187.395 ;
        RECT 45.715 186.485 48.445 187.395 ;
        RECT 48.475 186.525 48.905 187.310 ;
        RECT 48.925 186.485 52.135 187.395 ;
        RECT 53.065 186.715 60.375 187.395 ;
        RECT 56.580 186.495 57.490 186.715 ;
        RECT 59.025 186.485 60.375 186.715 ;
        RECT 60.425 186.585 61.795 187.395 ;
        RECT 61.805 186.715 64.095 187.395 ;
        RECT 63.175 186.485 64.095 186.715 ;
        RECT 64.115 186.485 66.845 187.395 ;
        RECT 67.880 186.715 71.345 187.395 ;
        RECT 71.925 186.715 74.215 187.395 ;
        RECT 67.880 186.485 68.800 186.715 ;
        RECT 71.925 186.485 72.845 186.715 ;
        RECT 74.235 186.525 74.665 187.310 ;
        RECT 74.685 186.585 76.515 187.395 ;
        RECT 76.535 186.485 79.265 187.395 ;
        RECT 79.295 186.485 82.025 187.395 ;
        RECT 82.045 186.585 83.415 187.395 ;
        RECT 83.435 186.485 86.165 187.395 ;
        RECT 86.185 186.585 91.695 187.395 ;
        RECT 91.705 186.585 97.215 187.395 ;
        RECT 98.145 186.485 99.975 187.395 ;
        RECT 99.995 186.525 100.425 187.310 ;
        RECT 100.455 186.485 103.655 187.395 ;
        RECT 103.665 187.365 104.610 187.395 ;
        RECT 106.565 187.365 106.735 187.585 ;
        RECT 109.320 187.445 109.440 187.555 ;
        RECT 109.785 187.395 109.955 187.605 ;
        RECT 110.245 187.395 110.415 187.585 ;
        RECT 116.685 187.395 116.855 187.605 ;
        RECT 117.145 187.415 117.315 187.605 ;
        RECT 121.285 187.395 121.455 187.585 ;
        RECT 121.740 187.445 121.860 187.555 ;
        RECT 122.205 187.395 122.375 187.605 ;
        RECT 122.665 187.415 122.835 187.605 ;
        RECT 124.500 187.415 124.670 187.605 ;
        RECT 125.420 187.445 125.540 187.555 ;
        RECT 125.890 187.415 126.060 187.635 ;
        RECT 127.550 187.605 128.495 187.635 ;
        RECT 129.275 188.285 130.205 188.515 ;
        RECT 129.275 187.605 131.110 188.285 ;
        RECT 131.265 187.605 134.935 188.415 ;
        RECT 135.415 187.605 136.765 188.515 ;
        RECT 136.785 187.605 138.615 188.415 ;
        RECT 138.635 187.690 139.065 188.475 ;
        RECT 140.135 188.285 141.065 188.515 ;
        RECT 142.525 188.425 143.475 188.515 ;
        RECT 139.230 187.605 141.065 188.285 ;
        RECT 141.545 187.605 143.475 188.425 ;
        RECT 143.685 188.315 144.615 188.515 ;
        RECT 145.945 188.315 146.895 188.515 ;
        RECT 143.685 187.835 146.895 188.315 ;
        RECT 151.340 188.285 152.250 188.505 ;
        RECT 153.785 188.285 155.135 188.515 ;
        RECT 143.830 187.635 146.895 187.835 ;
        RECT 130.945 187.585 131.110 187.605 ;
        RECT 126.350 187.395 126.520 187.585 ;
        RECT 128.640 187.445 128.760 187.555 ;
        RECT 129.565 187.395 129.735 187.585 ;
        RECT 130.945 187.415 131.115 187.585 ;
        RECT 131.405 187.415 131.575 187.605 ;
        RECT 135.080 187.445 135.200 187.555 ;
        RECT 135.545 187.395 135.715 187.585 ;
        RECT 136.465 187.415 136.635 187.605 ;
        RECT 136.925 187.395 137.095 187.605 ;
        RECT 139.230 187.585 139.395 187.605 ;
        RECT 141.545 187.585 141.695 187.605 ;
        RECT 138.760 187.445 138.880 187.555 ;
        RECT 139.225 187.415 139.395 187.585 ;
        RECT 141.065 187.395 141.235 187.585 ;
        RECT 141.525 187.395 141.695 187.585 ;
        RECT 143.830 187.415 144.000 187.635 ;
        RECT 145.960 187.605 146.895 187.635 ;
        RECT 147.825 187.605 155.135 188.285 ;
        RECT 155.645 187.605 157.015 188.415 ;
        RECT 145.205 187.415 145.375 187.585 ;
        RECT 145.205 187.395 145.370 187.415 ;
        RECT 145.665 187.395 145.835 187.585 ;
        RECT 147.055 187.450 147.215 187.560 ;
        RECT 147.500 187.445 147.620 187.555 ;
        RECT 147.965 187.395 148.135 187.605 ;
        RECT 149.345 187.395 149.515 187.585 ;
        RECT 151.180 187.445 151.300 187.555 ;
        RECT 152.105 187.395 152.275 187.585 ;
        RECT 155.320 187.445 155.440 187.555 ;
        RECT 156.705 187.395 156.875 187.605 ;
        RECT 103.665 187.165 106.735 187.365 ;
        RECT 103.665 186.685 106.875 187.165 ;
        RECT 103.665 186.485 104.610 186.685 ;
        RECT 105.945 186.485 106.875 186.685 ;
        RECT 106.885 186.485 110.055 187.395 ;
        RECT 110.105 186.485 113.315 187.395 ;
        RECT 113.420 186.715 116.885 187.395 ;
        RECT 118.020 186.715 121.485 187.395 ;
        RECT 113.420 186.485 114.340 186.715 ;
        RECT 118.020 186.485 118.940 186.715 ;
        RECT 122.065 186.485 125.275 187.395 ;
        RECT 125.755 186.525 126.185 187.310 ;
        RECT 126.205 186.485 129.415 187.395 ;
        RECT 129.425 186.585 134.935 187.395 ;
        RECT 135.405 186.615 136.775 187.395 ;
        RECT 136.785 186.585 138.615 187.395 ;
        RECT 139.085 186.715 141.375 187.395 ;
        RECT 139.085 186.485 140.005 186.715 ;
        RECT 141.385 186.585 143.215 187.395 ;
        RECT 143.535 186.715 145.370 187.395 ;
        RECT 143.535 186.485 144.465 186.715 ;
        RECT 145.525 186.585 147.355 187.395 ;
        RECT 147.825 186.615 149.195 187.395 ;
        RECT 149.205 186.585 151.035 187.395 ;
        RECT 151.515 186.525 151.945 187.310 ;
        RECT 151.965 186.585 155.635 187.395 ;
        RECT 155.645 186.585 157.015 187.395 ;
      LAYER nwell ;
        RECT 22.510 183.365 157.210 186.195 ;
      LAYER pwell ;
        RECT 22.705 182.165 24.075 182.975 ;
        RECT 24.085 182.165 29.595 182.975 ;
        RECT 29.605 182.165 31.435 182.975 ;
        RECT 31.445 182.165 32.795 183.075 ;
        RECT 32.845 182.165 34.195 183.075 ;
        RECT 34.205 182.165 35.575 182.945 ;
        RECT 35.595 182.250 36.025 183.035 ;
        RECT 36.045 182.165 40.860 182.845 ;
        RECT 41.105 182.165 42.935 182.975 ;
        RECT 43.405 182.165 46.325 183.075 ;
        RECT 46.625 182.165 52.135 182.975 ;
        RECT 52.145 182.165 54.895 182.975 ;
        RECT 54.905 182.165 58.115 183.075 ;
        RECT 60.415 182.845 61.335 183.075 ;
        RECT 59.045 182.165 61.335 182.845 ;
        RECT 61.355 182.250 61.785 183.035 ;
        RECT 65.320 182.845 66.230 183.065 ;
        RECT 67.765 182.845 69.115 183.075 ;
        RECT 61.805 182.165 69.115 182.845 ;
        RECT 69.625 182.165 72.835 183.075 ;
        RECT 72.845 182.165 74.215 182.975 ;
        RECT 79.380 182.845 80.300 183.075 ;
        RECT 86.080 182.845 87.000 183.075 ;
        RECT 74.225 182.165 79.040 182.845 ;
        RECT 79.380 182.165 82.845 182.845 ;
        RECT 83.535 182.165 87.000 182.845 ;
        RECT 87.115 182.250 87.545 183.035 ;
        RECT 91.080 182.845 91.990 183.065 ;
        RECT 93.525 182.845 94.875 183.075 ;
        RECT 87.565 182.165 94.875 182.845 ;
        RECT 95.125 182.985 96.075 183.075 ;
        RECT 98.365 182.985 99.315 183.075 ;
        RECT 95.125 182.165 97.055 182.985 ;
        RECT 22.845 181.955 23.015 182.165 ;
        RECT 24.225 181.955 24.395 182.165 ;
        RECT 29.745 181.975 29.915 182.165 ;
        RECT 31.585 181.975 31.755 182.145 ;
        RECT 32.510 181.975 32.680 182.165 ;
        RECT 32.960 181.975 33.130 182.165 ;
        RECT 31.590 181.955 31.755 181.975 ;
        RECT 33.885 181.955 34.055 182.145 ;
        RECT 34.345 181.975 34.515 182.165 ;
        RECT 36.185 181.975 36.355 182.165 ;
        RECT 41.245 181.975 41.415 182.165 ;
        RECT 43.080 182.005 43.200 182.115 ;
        RECT 43.550 181.975 43.720 182.165 ;
        RECT 22.705 181.145 24.075 181.955 ;
        RECT 24.085 181.275 31.395 181.955 ;
        RECT 31.590 181.275 33.425 181.955 ;
        RECT 33.745 181.275 41.055 181.955 ;
        RECT 27.600 181.055 28.510 181.275 ;
        RECT 30.045 181.045 31.395 181.275 ;
        RECT 32.495 181.045 33.425 181.275 ;
        RECT 37.260 181.055 38.170 181.275 ;
        RECT 39.705 181.045 41.055 181.275 ;
        RECT 42.025 181.925 42.970 181.955 ;
        RECT 44.925 181.925 45.095 182.145 ;
        RECT 42.025 181.725 45.095 181.925 ;
        RECT 45.385 181.925 45.555 182.145 ;
        RECT 46.765 181.975 46.935 182.165 ;
        RECT 49.065 181.955 49.235 182.145 ;
        RECT 52.285 181.975 52.455 182.165 ;
        RECT 56.420 181.955 56.590 182.145 ;
        RECT 56.895 182.000 57.055 182.110 ;
        RECT 57.805 181.975 57.975 182.165 ;
        RECT 58.275 182.010 58.435 182.120 ;
        RECT 59.185 181.975 59.355 182.165 ;
        RECT 60.565 181.955 60.735 182.145 ;
        RECT 61.025 181.955 61.195 182.145 ;
        RECT 61.945 181.975 62.115 182.165 ;
        RECT 65.625 181.955 65.795 182.145 ;
        RECT 69.305 182.115 69.475 182.145 ;
        RECT 66.095 182.000 66.255 182.110 ;
        RECT 69.300 182.005 69.475 182.115 ;
        RECT 69.305 181.955 69.475 182.005 ;
        RECT 69.765 181.975 69.935 182.165 ;
        RECT 72.985 181.955 73.155 182.165 ;
        RECT 73.455 182.000 73.615 182.110 ;
        RECT 74.365 181.975 74.535 182.165 ;
        RECT 74.835 182.000 74.995 182.110 ;
        RECT 75.745 181.955 75.915 182.145 ;
        RECT 82.645 181.975 82.815 182.165 ;
        RECT 83.100 182.005 83.220 182.115 ;
        RECT 83.565 181.975 83.735 182.165 ;
        RECT 84.945 181.955 85.115 182.145 ;
        RECT 85.405 181.955 85.575 182.145 ;
        RECT 87.705 181.975 87.875 182.165 ;
        RECT 96.905 182.145 97.055 182.165 ;
        RECT 97.385 182.165 99.315 182.985 ;
        RECT 102.025 182.985 102.975 183.075 ;
        RECT 99.525 182.165 101.355 182.975 ;
        RECT 102.025 182.165 103.955 182.985 ;
        RECT 104.125 182.165 107.795 182.975 ;
        RECT 108.265 182.165 111.475 183.075 ;
        RECT 111.485 182.165 112.855 182.975 ;
        RECT 112.875 182.250 113.305 183.035 ;
        RECT 116.840 182.845 117.750 183.065 ;
        RECT 119.285 182.845 120.635 183.075 ;
        RECT 113.325 182.165 120.635 182.845 ;
        RECT 120.685 182.165 122.500 183.075 ;
        RECT 123.645 182.985 124.595 183.075 ;
        RECT 123.645 182.165 125.575 182.985 ;
        RECT 125.755 182.165 127.105 183.075 ;
        RECT 127.125 182.165 130.795 182.975 ;
        RECT 131.305 182.845 132.655 183.075 ;
        RECT 134.190 182.845 135.100 183.065 ;
        RECT 131.305 182.165 138.615 182.845 ;
        RECT 138.635 182.250 139.065 183.035 ;
        RECT 139.085 182.845 140.005 183.075 ;
        RECT 141.385 182.875 142.315 183.075 ;
        RECT 143.645 182.875 144.595 183.075 ;
        RECT 139.085 182.165 141.375 182.845 ;
        RECT 141.385 182.395 144.595 182.875 ;
        RECT 141.530 182.195 144.595 182.395 ;
        RECT 97.385 182.145 97.535 182.165 ;
        RECT 89.080 182.005 89.200 182.115 ;
        RECT 90.465 181.955 90.635 182.145 ;
        RECT 90.935 182.000 91.095 182.110 ;
        RECT 92.120 181.955 92.290 182.145 ;
        RECT 95.985 181.955 96.155 182.145 ;
        RECT 96.905 181.975 97.075 182.145 ;
        RECT 97.365 181.975 97.535 182.145 ;
        RECT 99.665 182.115 99.835 182.165 ;
        RECT 103.805 182.145 103.955 182.165 ;
        RECT 99.660 182.005 99.835 182.115 ;
        RECT 99.665 181.975 99.835 182.005 ;
        RECT 100.585 181.955 100.755 182.145 ;
        RECT 101.500 182.005 101.620 182.115 ;
        RECT 103.805 181.975 103.975 182.145 ;
        RECT 104.265 181.975 104.435 182.165 ;
        RECT 106.105 181.955 106.275 182.145 ;
        RECT 107.940 182.005 108.060 182.115 ;
        RECT 108.865 181.955 109.035 182.145 ;
        RECT 111.165 181.975 111.335 182.165 ;
        RECT 111.625 181.975 111.795 182.165 ;
        RECT 113.465 181.975 113.635 182.165 ;
        RECT 116.225 181.955 116.395 182.145 ;
        RECT 119.915 182.000 120.075 182.110 ;
        RECT 120.825 181.955 120.995 182.145 ;
        RECT 122.205 181.955 122.375 182.165 ;
        RECT 125.425 182.145 125.575 182.165 ;
        RECT 122.675 182.010 122.835 182.120 ;
        RECT 125.425 181.975 125.595 182.145 ;
        RECT 125.885 181.975 126.055 182.165 ;
        RECT 126.340 182.005 126.460 182.115 ;
        RECT 126.805 181.975 126.975 182.145 ;
        RECT 127.265 181.975 127.435 182.165 ;
        RECT 130.940 182.005 131.060 182.115 ;
        RECT 126.805 181.955 127.005 181.975 ;
        RECT 133.240 181.955 133.410 182.145 ;
        RECT 133.705 181.975 133.875 182.145 ;
        RECT 136.015 182.000 136.175 182.110 ;
        RECT 138.305 181.975 138.475 182.165 ;
        RECT 138.765 181.975 138.935 182.145 ;
        RECT 133.725 181.955 133.875 181.975 ;
        RECT 138.765 181.955 138.930 181.975 ;
        RECT 140.150 181.955 140.320 182.145 ;
        RECT 140.605 181.955 140.775 182.145 ;
        RECT 141.065 181.975 141.235 182.165 ;
        RECT 141.530 181.975 141.700 182.195 ;
        RECT 143.660 182.165 144.595 182.195 ;
        RECT 144.645 182.845 145.995 183.075 ;
        RECT 147.530 182.845 148.440 183.065 ;
        RECT 144.645 182.165 151.955 182.845 ;
        RECT 151.965 182.165 155.635 182.975 ;
        RECT 155.645 182.165 157.015 182.975 ;
        RECT 142.440 182.005 142.560 182.115 ;
        RECT 142.905 181.955 143.075 182.145 ;
        RECT 144.740 182.005 144.860 182.115 ;
        RECT 145.205 181.955 145.375 182.145 ;
        RECT 146.585 181.955 146.755 182.145 ;
        RECT 151.645 181.975 151.815 182.165 ;
        RECT 152.105 181.955 152.275 182.165 ;
        RECT 156.705 181.955 156.875 182.165 ;
        RECT 47.510 181.925 48.455 181.955 ;
        RECT 45.385 181.725 48.455 181.925 ;
        RECT 42.025 181.245 45.235 181.725 ;
        RECT 42.025 181.045 42.970 181.245 ;
        RECT 44.305 181.045 45.235 181.245 ;
        RECT 45.245 181.245 48.455 181.725 ;
        RECT 45.245 181.045 46.175 181.245 ;
        RECT 47.510 181.045 48.455 181.245 ;
        RECT 48.475 181.085 48.905 181.870 ;
        RECT 48.925 181.145 54.435 181.955 ;
        RECT 54.525 181.045 56.735 181.955 ;
        RECT 57.665 181.045 60.875 181.955 ;
        RECT 60.885 181.145 62.255 181.955 ;
        RECT 62.360 181.275 65.825 181.955 ;
        RECT 62.360 181.045 63.280 181.275 ;
        RECT 66.875 181.045 69.605 181.955 ;
        RECT 69.720 181.275 73.185 181.955 ;
        RECT 69.720 181.045 70.640 181.275 ;
        RECT 74.235 181.085 74.665 181.870 ;
        RECT 75.605 181.275 82.915 181.955 ;
        RECT 79.120 181.055 80.030 181.275 ;
        RECT 81.565 181.045 82.915 181.275 ;
        RECT 82.965 181.275 85.255 181.955 ;
        RECT 82.965 181.045 83.885 181.275 ;
        RECT 85.265 181.145 88.935 181.955 ;
        RECT 89.405 181.175 90.775 181.955 ;
        RECT 91.705 181.275 95.605 181.955 ;
        RECT 91.705 181.045 92.635 181.275 ;
        RECT 95.845 181.145 99.515 181.955 ;
        RECT 99.995 181.085 100.425 181.870 ;
        RECT 100.445 181.145 105.955 181.955 ;
        RECT 105.965 181.145 108.715 181.955 ;
        RECT 108.725 181.275 116.035 181.955 ;
        RECT 112.240 181.055 113.150 181.275 ;
        RECT 114.685 181.045 116.035 181.275 ;
        RECT 116.085 181.145 119.755 181.955 ;
        RECT 120.695 181.045 122.045 181.955 ;
        RECT 122.065 181.145 125.735 181.955 ;
        RECT 125.755 181.085 126.185 181.870 ;
        RECT 126.805 181.275 130.335 181.955 ;
        RECT 127.510 181.045 130.335 181.275 ;
        RECT 130.635 181.045 133.555 181.955 ;
        RECT 133.725 181.135 135.655 181.955 ;
        RECT 134.705 181.045 135.655 181.135 ;
        RECT 137.095 181.275 138.930 181.955 ;
        RECT 137.095 181.045 138.025 181.275 ;
        RECT 139.085 181.045 140.435 181.955 ;
        RECT 140.465 181.145 142.295 181.955 ;
        RECT 142.765 181.275 144.595 181.955 ;
        RECT 145.065 181.175 146.435 181.955 ;
        RECT 146.445 181.275 151.260 181.955 ;
        RECT 151.515 181.085 151.945 181.870 ;
        RECT 151.965 181.145 155.635 181.955 ;
        RECT 155.645 181.145 157.015 181.955 ;
      LAYER nwell ;
        RECT 22.510 177.925 157.210 180.755 ;
      LAYER pwell ;
        RECT 22.705 176.725 24.075 177.535 ;
        RECT 25.005 176.725 26.375 177.505 ;
        RECT 26.385 176.725 28.215 177.535 ;
        RECT 28.225 177.405 29.145 177.635 ;
        RECT 28.225 176.725 30.515 177.405 ;
        RECT 30.525 176.725 31.895 177.535 ;
        RECT 33.275 177.405 34.195 177.635 ;
        RECT 31.905 176.725 34.195 177.405 ;
        RECT 34.215 176.725 35.565 177.635 ;
        RECT 35.595 176.810 36.025 177.595 ;
        RECT 36.045 176.725 39.715 177.535 ;
        RECT 41.990 177.435 42.935 177.635 ;
        RECT 40.185 176.755 42.935 177.435 ;
        RECT 22.845 176.515 23.015 176.725 ;
        RECT 24.225 176.515 24.395 176.705 ;
        RECT 26.065 176.535 26.235 176.725 ;
        RECT 26.525 176.535 26.695 176.725 ;
        RECT 27.915 176.560 28.075 176.670 ;
        RECT 29.750 176.515 29.920 176.705 ;
        RECT 30.205 176.535 30.375 176.725 ;
        RECT 30.665 176.535 30.835 176.725 ;
        RECT 32.045 176.535 32.215 176.725 ;
        RECT 32.515 176.560 32.675 176.670 ;
        RECT 32.045 176.515 32.195 176.535 ;
        RECT 34.345 176.515 34.515 176.725 ;
        RECT 34.805 176.515 34.975 176.705 ;
        RECT 36.185 176.535 36.355 176.725 ;
        RECT 40.330 176.705 40.500 176.755 ;
        RECT 41.990 176.725 42.935 176.755 ;
        RECT 43.445 176.725 46.615 177.635 ;
        RECT 46.625 176.725 48.455 177.535 ;
        RECT 48.505 177.405 49.855 177.635 ;
        RECT 51.390 177.405 52.300 177.625 ;
        RECT 55.920 177.405 56.840 177.635 ;
        RECT 48.505 176.725 55.815 177.405 ;
        RECT 55.920 176.725 59.385 177.405 ;
        RECT 59.505 176.725 61.335 177.535 ;
        RECT 61.355 176.810 61.785 177.595 ;
        RECT 61.805 176.725 63.175 177.535 ;
        RECT 66.700 177.405 67.610 177.625 ;
        RECT 69.145 177.405 70.495 177.635 ;
        RECT 74.060 177.405 74.970 177.625 ;
        RECT 76.505 177.405 77.855 177.635 ;
        RECT 63.185 176.725 70.495 177.405 ;
        RECT 70.545 176.725 77.855 177.405 ;
        RECT 77.905 176.725 79.735 177.535 ;
        RECT 83.260 177.405 84.170 177.625 ;
        RECT 85.705 177.405 87.055 177.635 ;
        RECT 79.745 176.725 87.055 177.405 ;
        RECT 87.115 176.810 87.545 177.595 ;
        RECT 90.680 177.405 91.600 177.635 ;
        RECT 88.135 176.725 91.600 177.405 ;
        RECT 91.705 177.405 92.625 177.635 ;
        RECT 95.585 177.545 96.535 177.635 ;
        RECT 91.705 176.725 93.995 177.405 ;
        RECT 94.005 176.725 95.375 177.505 ;
        RECT 95.585 176.725 97.515 177.545 ;
        RECT 98.145 176.725 99.515 177.505 ;
        RECT 103.040 177.405 103.950 177.625 ;
        RECT 105.485 177.405 106.835 177.635 ;
        RECT 99.525 176.725 106.835 177.405 ;
        RECT 107.085 177.545 108.035 177.635 ;
        RECT 107.085 176.725 109.015 177.545 ;
        RECT 109.725 176.725 111.935 177.635 ;
        RECT 112.875 176.810 113.305 177.595 ;
        RECT 113.325 176.725 115.155 177.535 ;
        RECT 115.165 176.725 116.535 177.505 ;
        RECT 120.060 177.405 120.970 177.625 ;
        RECT 122.505 177.405 123.855 177.635 ;
        RECT 116.545 176.725 123.855 177.405 ;
        RECT 123.905 176.725 127.575 177.535 ;
        RECT 129.865 177.405 130.795 177.635 ;
        RECT 128.045 176.725 130.795 177.405 ;
        RECT 130.805 176.725 134.475 177.535 ;
        RECT 134.945 177.435 135.875 177.635 ;
        RECT 137.210 177.435 138.155 177.635 ;
        RECT 134.945 176.955 138.155 177.435 ;
        RECT 135.085 176.755 138.155 176.955 ;
        RECT 138.635 176.810 139.065 177.595 ;
        RECT 140.455 177.405 141.375 177.635 ;
        RECT 39.860 176.565 39.980 176.675 ;
        RECT 40.325 176.535 40.500 176.705 ;
        RECT 43.080 176.565 43.200 176.675 ;
        RECT 43.545 176.535 43.715 176.725 ;
        RECT 40.325 176.515 40.495 176.535 ;
        RECT 22.705 175.705 24.075 176.515 ;
        RECT 24.085 175.705 27.755 176.515 ;
        RECT 28.685 175.605 30.035 176.515 ;
        RECT 30.265 175.695 32.195 176.515 ;
        RECT 30.265 175.605 31.215 175.695 ;
        RECT 33.295 175.605 34.645 176.515 ;
        RECT 34.665 175.705 40.175 176.515 ;
        RECT 40.185 175.705 41.555 176.515 ;
        RECT 41.565 176.485 42.510 176.515 ;
        RECT 44.000 176.485 44.170 176.705 ;
        RECT 44.465 176.515 44.635 176.705 ;
        RECT 46.765 176.535 46.935 176.725 ;
        RECT 48.140 176.565 48.260 176.675 ;
        RECT 49.065 176.515 49.235 176.705 ;
        RECT 53.665 176.515 53.835 176.705 ;
        RECT 54.125 176.515 54.295 176.705 ;
        RECT 55.505 176.535 55.675 176.725 ;
        RECT 57.345 176.515 57.515 176.705 ;
        RECT 59.185 176.535 59.355 176.725 ;
        RECT 59.645 176.535 59.815 176.725 ;
        RECT 61.945 176.535 62.115 176.725 ;
        RECT 63.325 176.535 63.495 176.725 ;
        RECT 64.705 176.515 64.875 176.705 ;
        RECT 66.545 176.515 66.715 176.705 ;
        RECT 69.305 176.515 69.475 176.705 ;
        RECT 70.685 176.535 70.855 176.725 ;
        RECT 72.525 176.515 72.695 176.705 ;
        RECT 72.985 176.515 73.155 176.705 ;
        RECT 78.045 176.515 78.215 176.725 ;
        RECT 79.885 176.515 80.055 176.725 ;
        RECT 80.345 176.515 80.515 176.705 ;
        RECT 83.105 176.515 83.275 176.705 ;
        RECT 85.865 176.515 86.035 176.705 ;
        RECT 87.700 176.565 87.820 176.675 ;
        RECT 88.165 176.535 88.335 176.725 ;
        RECT 89.545 176.515 89.715 176.705 ;
        RECT 90.925 176.515 91.095 176.705 ;
        RECT 93.685 176.535 93.855 176.725 ;
        RECT 95.065 176.535 95.235 176.725 ;
        RECT 97.365 176.705 97.515 176.725 ;
        RECT 97.365 176.535 97.535 176.705 ;
        RECT 97.820 176.565 97.940 176.675 ;
        RECT 98.285 176.515 98.455 176.725 ;
        RECT 99.665 176.535 99.835 176.725 ;
        RECT 108.865 176.705 109.015 176.725 ;
        RECT 100.860 176.515 101.030 176.705 ;
        RECT 104.725 176.515 104.895 176.705 ;
        RECT 107.480 176.565 107.600 176.675 ;
        RECT 108.865 176.535 109.035 176.705 ;
        RECT 109.320 176.565 109.440 176.675 ;
        RECT 109.785 176.535 109.955 176.705 ;
        RECT 109.785 176.515 109.935 176.535 ;
        RECT 110.245 176.515 110.415 176.705 ;
        RECT 111.620 176.535 111.790 176.725 ;
        RECT 112.095 176.570 112.255 176.680 ;
        RECT 113.465 176.535 113.635 176.725 ;
        RECT 113.920 176.565 114.040 176.675 ;
        RECT 115.305 176.535 115.475 176.725 ;
        RECT 116.225 176.535 116.395 176.705 ;
        RECT 116.685 176.535 116.855 176.725 ;
        RECT 116.225 176.515 116.375 176.535 ;
        RECT 117.880 176.515 118.050 176.705 ;
        RECT 123.585 176.535 123.755 176.705 ;
        RECT 123.585 176.515 123.735 176.535 ;
        RECT 124.045 176.515 124.215 176.725 ;
        RECT 126.340 176.565 126.460 176.675 ;
        RECT 126.805 176.535 126.975 176.705 ;
        RECT 127.720 176.565 127.840 176.675 ;
        RECT 128.185 176.535 128.355 176.725 ;
        RECT 126.815 176.515 126.975 176.535 ;
        RECT 130.945 176.515 131.115 176.725 ;
        RECT 132.780 176.565 132.900 176.675 ;
        RECT 134.620 176.565 134.740 176.675 ;
        RECT 135.085 176.535 135.255 176.755 ;
        RECT 137.210 176.725 138.155 176.755 ;
        RECT 139.085 176.725 141.375 177.405 ;
        RECT 141.395 176.725 142.745 177.635 ;
        RECT 142.765 176.725 144.135 177.505 ;
        RECT 144.165 176.725 145.515 177.635 ;
        RECT 145.545 176.725 146.895 177.635 ;
        RECT 146.905 176.725 148.275 177.535 ;
        RECT 151.800 177.405 152.710 177.625 ;
        RECT 154.245 177.405 155.595 177.635 ;
        RECT 148.285 176.725 155.595 177.405 ;
        RECT 155.645 176.725 157.015 177.535 ;
        RECT 136.465 176.515 136.635 176.705 ;
        RECT 136.925 176.515 137.095 176.705 ;
        RECT 138.300 176.565 138.420 176.675 ;
        RECT 138.765 176.515 138.935 176.705 ;
        RECT 139.225 176.535 139.395 176.725 ;
        RECT 141.525 176.535 141.695 176.725 ;
        RECT 142.905 176.535 143.075 176.725 ;
        RECT 144.280 176.705 144.450 176.725 ;
        RECT 145.660 176.705 145.830 176.725 ;
        RECT 144.280 176.535 144.455 176.705 ;
        RECT 144.755 176.560 144.915 176.670 ;
        RECT 145.660 176.535 145.835 176.705 ;
        RECT 147.045 176.535 147.215 176.725 ;
        RECT 144.285 176.515 144.450 176.535 ;
        RECT 41.565 175.805 44.315 176.485 ;
        RECT 41.565 175.605 42.510 175.805 ;
        RECT 44.325 175.705 47.995 176.515 ;
        RECT 48.475 175.645 48.905 176.430 ;
        RECT 48.925 175.705 50.755 176.515 ;
        RECT 50.765 175.605 53.975 176.515 ;
        RECT 53.985 175.605 57.195 176.515 ;
        RECT 57.205 175.835 64.515 176.515 ;
        RECT 60.720 175.615 61.630 175.835 ;
        RECT 63.165 175.605 64.515 175.835 ;
        RECT 64.565 175.705 66.395 176.515 ;
        RECT 66.415 175.605 69.145 176.515 ;
        RECT 69.165 175.705 70.535 176.515 ;
        RECT 70.545 175.835 72.835 176.515 ;
        RECT 70.545 175.605 71.465 175.835 ;
        RECT 72.845 175.705 74.215 176.515 ;
        RECT 74.235 175.645 74.665 176.430 ;
        RECT 74.780 175.835 78.245 176.515 ;
        RECT 78.365 175.835 80.195 176.515 ;
        RECT 74.780 175.605 75.700 175.835 ;
        RECT 80.205 175.705 82.955 176.515 ;
        RECT 82.975 175.605 85.705 176.515 ;
        RECT 85.725 175.705 89.395 176.515 ;
        RECT 89.405 175.705 90.775 176.515 ;
        RECT 90.785 175.835 98.095 176.515 ;
        RECT 94.300 175.615 95.210 175.835 ;
        RECT 96.745 175.605 98.095 175.835 ;
        RECT 98.145 175.705 99.975 176.515 ;
        RECT 99.995 175.645 100.425 176.430 ;
        RECT 100.445 175.835 104.345 176.515 ;
        RECT 100.445 175.605 101.375 175.835 ;
        RECT 104.585 175.705 107.335 176.515 ;
        RECT 108.005 175.695 109.935 176.515 ;
        RECT 110.105 175.705 113.775 176.515 ;
        RECT 114.445 175.695 116.375 176.515 ;
        RECT 117.465 175.835 121.365 176.515 ;
        RECT 108.005 175.605 108.955 175.695 ;
        RECT 114.445 175.605 115.395 175.695 ;
        RECT 117.465 175.605 118.395 175.835 ;
        RECT 121.805 175.695 123.735 176.515 ;
        RECT 123.905 175.705 125.735 176.515 ;
        RECT 121.805 175.605 122.755 175.695 ;
        RECT 125.755 175.645 126.185 176.430 ;
        RECT 126.815 175.605 130.470 176.515 ;
        RECT 130.805 175.705 132.635 176.515 ;
        RECT 133.200 175.835 136.665 176.515 ;
        RECT 133.200 175.605 134.120 175.835 ;
        RECT 136.800 175.605 138.615 176.515 ;
        RECT 138.735 175.835 142.200 176.515 ;
        RECT 141.280 175.605 142.200 175.835 ;
        RECT 142.615 175.835 144.450 176.515 ;
        RECT 145.670 176.515 145.835 176.535 ;
        RECT 147.965 176.515 148.135 176.705 ;
        RECT 148.425 176.535 148.595 176.725 ;
        RECT 151.185 176.515 151.355 176.705 ;
        RECT 152.105 176.515 152.275 176.705 ;
        RECT 154.405 176.515 154.575 176.705 ;
        RECT 154.875 176.560 155.035 176.670 ;
        RECT 156.705 176.515 156.875 176.725 ;
        RECT 145.670 175.835 147.505 176.515 ;
        RECT 147.825 175.835 150.115 176.515 ;
        RECT 142.615 175.605 143.545 175.835 ;
        RECT 146.575 175.605 147.505 175.835 ;
        RECT 149.195 175.605 150.115 175.835 ;
        RECT 150.125 175.735 151.495 176.515 ;
        RECT 151.515 175.645 151.945 176.430 ;
        RECT 151.965 175.705 153.335 176.515 ;
        RECT 153.355 175.605 154.705 176.515 ;
        RECT 155.645 175.705 157.015 176.515 ;
      LAYER nwell ;
        RECT 22.510 172.485 157.210 175.315 ;
      LAYER pwell ;
        RECT 22.705 171.285 24.075 172.095 ;
        RECT 24.085 171.285 25.455 172.065 ;
        RECT 25.485 171.285 26.835 172.195 ;
        RECT 26.845 171.995 27.795 172.195 ;
        RECT 29.125 171.995 30.055 172.195 ;
        RECT 26.845 171.515 30.055 171.995 ;
        RECT 31.895 171.965 32.815 172.195 ;
        RECT 26.845 171.315 29.910 171.515 ;
        RECT 26.845 171.285 27.780 171.315 ;
        RECT 22.845 171.075 23.015 171.285 ;
        RECT 24.225 171.075 24.395 171.285 ;
        RECT 25.600 171.095 25.770 171.285 ;
        RECT 29.740 171.095 29.910 171.315 ;
        RECT 30.525 171.285 32.815 171.965 ;
        RECT 32.825 171.965 33.745 172.195 ;
        RECT 32.825 171.285 35.115 171.965 ;
        RECT 35.595 171.370 36.025 172.155 ;
        RECT 36.975 171.285 38.325 172.195 ;
        RECT 38.635 171.285 41.555 172.195 ;
        RECT 41.565 171.285 44.775 172.195 ;
        RECT 46.120 171.995 47.075 172.195 ;
        RECT 44.795 171.315 47.075 171.995 ;
        RECT 50.600 171.965 51.510 172.185 ;
        RECT 53.045 171.965 54.395 172.195 ;
        RECT 30.200 171.125 30.320 171.235 ;
        RECT 30.665 171.095 30.835 171.285 ;
        RECT 31.595 171.120 31.755 171.230 ;
        RECT 22.705 170.265 24.075 171.075 ;
        RECT 24.085 170.395 31.395 171.075 ;
        RECT 32.510 171.045 32.680 171.265 ;
        RECT 34.805 171.095 34.975 171.285 ;
        RECT 35.265 171.235 35.435 171.265 ;
        RECT 35.260 171.125 35.435 171.235 ;
        RECT 36.195 171.130 36.355 171.240 ;
        RECT 35.265 171.075 35.435 171.125 ;
        RECT 37.105 171.095 37.275 171.285 ;
        RECT 38.485 171.075 38.655 171.265 ;
        RECT 39.865 171.095 40.035 171.265 ;
        RECT 41.240 171.095 41.410 171.285 ;
        RECT 41.705 171.095 41.875 171.285 ;
        RECT 39.990 171.075 40.035 171.095 ;
        RECT 44.010 171.075 44.180 171.265 ;
        RECT 44.465 171.075 44.635 171.265 ;
        RECT 44.920 171.095 45.090 171.315 ;
        RECT 46.120 171.285 47.075 171.315 ;
        RECT 47.085 171.285 54.395 171.965 ;
        RECT 54.445 171.285 55.815 172.095 ;
        RECT 55.920 171.965 56.840 172.195 ;
        RECT 55.920 171.285 59.385 171.965 ;
        RECT 59.505 171.285 61.335 172.095 ;
        RECT 61.355 171.370 61.785 172.155 ;
        RECT 61.900 171.965 62.820 172.195 ;
        RECT 61.900 171.285 65.365 171.965 ;
        RECT 65.485 171.285 67.315 172.095 ;
        RECT 70.840 171.965 71.750 172.185 ;
        RECT 73.285 171.965 74.635 172.195 ;
        RECT 80.040 171.965 80.950 172.185 ;
        RECT 82.485 171.965 83.835 172.195 ;
        RECT 67.325 171.285 74.635 171.965 ;
        RECT 74.685 171.285 76.515 171.965 ;
        RECT 76.525 171.285 83.835 171.965 ;
        RECT 83.885 171.285 86.095 172.195 ;
        RECT 87.115 171.370 87.545 172.155 ;
        RECT 87.565 171.965 88.485 172.195 ;
        RECT 87.565 171.285 89.855 171.965 ;
        RECT 89.865 171.285 91.235 172.065 ;
        RECT 91.245 171.285 93.075 172.095 ;
        RECT 93.085 171.965 94.015 172.195 ;
        RECT 93.085 171.285 96.985 171.965 ;
        RECT 97.225 171.285 99.055 172.095 ;
        RECT 99.525 171.285 102.265 171.965 ;
        RECT 102.285 171.285 103.655 172.065 ;
        RECT 107.180 171.965 108.090 172.185 ;
        RECT 109.625 171.965 110.975 172.195 ;
        RECT 103.665 171.285 110.975 171.965 ;
        RECT 111.485 171.285 112.855 172.065 ;
        RECT 112.875 171.370 113.305 172.155 ;
        RECT 116.840 171.965 117.750 172.185 ;
        RECT 119.285 171.965 120.635 172.195 ;
        RECT 113.325 171.285 120.635 171.965 ;
        RECT 120.885 172.105 121.835 172.195 ;
        RECT 120.885 171.285 122.815 172.105 ;
        RECT 123.445 171.285 126.655 172.195 ;
        RECT 126.680 171.285 130.335 172.195 ;
        RECT 134.780 171.965 135.690 172.185 ;
        RECT 137.225 171.965 138.575 172.195 ;
        RECT 131.265 171.285 138.575 171.965 ;
        RECT 138.635 171.370 139.065 172.155 ;
        RECT 140.045 171.965 141.395 172.195 ;
        RECT 142.930 171.965 143.840 172.185 ;
        RECT 148.145 171.965 150.105 172.195 ;
        RECT 140.045 171.285 147.355 171.965 ;
        RECT 147.655 171.285 150.105 171.965 ;
        RECT 150.125 171.285 151.955 172.095 ;
        RECT 152.435 171.285 153.785 172.195 ;
        RECT 153.805 171.285 155.635 172.095 ;
        RECT 155.645 171.285 157.015 172.095 ;
        RECT 47.225 171.095 47.395 171.285 ;
        RECT 48.140 171.125 48.260 171.235 ;
        RECT 49.060 171.125 49.180 171.235 ;
        RECT 49.530 171.075 49.700 171.265 ;
        RECT 54.585 171.095 54.755 171.285 ;
        RECT 55.045 171.075 55.215 171.265 ;
        RECT 55.505 171.075 55.675 171.265 ;
        RECT 59.185 171.095 59.355 171.285 ;
        RECT 59.645 171.095 59.815 171.285 ;
        RECT 65.165 171.095 65.335 171.285 ;
        RECT 65.625 171.075 65.795 171.285 ;
        RECT 66.085 171.075 66.255 171.265 ;
        RECT 67.465 171.095 67.635 171.285 ;
        RECT 69.765 171.075 69.935 171.265 ;
        RECT 72.525 171.075 72.695 171.265 ;
        RECT 74.825 171.075 74.995 171.265 ;
        RECT 76.205 171.095 76.375 171.285 ;
        RECT 76.665 171.095 76.835 171.285 ;
        RECT 78.500 171.125 78.620 171.235 ;
        RECT 78.965 171.075 79.135 171.265 ;
        RECT 81.735 171.120 81.895 171.230 ;
        RECT 84.030 171.095 84.200 171.285 ;
        RECT 86.050 171.075 86.220 171.265 ;
        RECT 86.335 171.130 86.495 171.240 ;
        RECT 86.785 171.075 86.955 171.265 ;
        RECT 89.545 171.095 89.715 171.285 ;
        RECT 90.925 171.095 91.095 171.285 ;
        RECT 91.385 171.095 91.555 171.285 ;
        RECT 93.500 171.095 93.670 171.285 ;
        RECT 94.145 171.075 94.315 171.265 ;
        RECT 95.980 171.125 96.100 171.235 ;
        RECT 97.365 171.075 97.535 171.285 ;
        RECT 97.825 171.095 97.995 171.265 ;
        RECT 99.200 171.125 99.320 171.235 ;
        RECT 99.665 171.095 99.835 171.285 ;
        RECT 97.845 171.075 97.995 171.095 ;
        RECT 100.860 171.075 101.030 171.265 ;
        RECT 102.425 171.095 102.595 171.285 ;
        RECT 103.805 171.095 103.975 171.285 ;
        RECT 104.720 171.125 104.840 171.235 ;
        RECT 105.460 171.075 105.630 171.265 ;
        RECT 109.325 171.075 109.495 171.265 ;
        RECT 111.160 171.125 111.280 171.235 ;
        RECT 111.625 171.095 111.795 171.285 ;
        RECT 112.360 171.075 112.530 171.265 ;
        RECT 113.465 171.095 113.635 171.285 ;
        RECT 122.665 171.265 122.815 171.285 ;
        RECT 116.235 171.120 116.395 171.230 ;
        RECT 117.145 171.075 117.315 171.265 ;
        RECT 118.525 171.075 118.695 171.265 ;
        RECT 122.665 171.095 122.835 171.265 ;
        RECT 123.120 171.125 123.240 171.235 ;
        RECT 126.345 171.075 126.515 171.285 ;
        RECT 130.020 171.095 130.190 171.285 ;
        RECT 130.495 171.130 130.655 171.240 ;
        RECT 131.405 171.095 131.575 171.285 ;
        RECT 132.325 171.075 132.495 171.265 ;
        RECT 132.785 171.075 132.955 171.265 ;
        RECT 139.225 171.075 139.395 171.265 ;
        RECT 139.685 171.075 139.855 171.265 ;
        RECT 141.525 171.075 141.695 171.265 ;
        RECT 143.825 171.075 143.995 171.265 ;
        RECT 147.045 171.095 147.215 171.285 ;
        RECT 147.655 171.265 147.675 171.285 ;
        RECT 147.505 171.095 147.675 171.265 ;
        RECT 149.345 171.075 149.515 171.265 ;
        RECT 150.265 171.095 150.435 171.285 ;
        RECT 151.180 171.125 151.300 171.235 ;
        RECT 152.100 171.125 152.220 171.235 ;
        RECT 153.485 171.095 153.655 171.285 ;
        RECT 153.945 171.095 154.115 171.285 ;
        RECT 155.325 171.075 155.495 171.265 ;
        RECT 156.705 171.075 156.875 171.285 ;
        RECT 34.170 171.045 35.115 171.075 ;
        RECT 27.600 170.175 28.510 170.395 ;
        RECT 30.045 170.165 31.395 170.395 ;
        RECT 32.365 170.365 35.115 171.045 ;
        RECT 34.170 170.165 35.115 170.365 ;
        RECT 35.125 170.165 38.335 171.075 ;
        RECT 38.345 170.265 39.715 171.075 ;
        RECT 39.990 170.165 42.925 171.075 ;
        RECT 42.945 170.165 44.295 171.075 ;
        RECT 44.325 170.265 47.995 171.075 ;
        RECT 48.475 170.205 48.905 170.990 ;
        RECT 49.385 170.165 51.995 171.075 ;
        RECT 52.145 170.165 55.355 171.075 ;
        RECT 55.365 170.165 58.575 171.075 ;
        RECT 58.625 170.395 65.935 171.075 ;
        RECT 58.625 170.165 59.975 170.395 ;
        RECT 61.510 170.175 62.420 170.395 ;
        RECT 65.945 170.265 69.615 171.075 ;
        RECT 69.635 170.165 72.365 171.075 ;
        RECT 72.385 170.265 74.215 171.075 ;
        RECT 74.235 170.205 74.665 170.990 ;
        RECT 74.685 170.265 78.355 171.075 ;
        RECT 78.835 170.165 81.565 171.075 ;
        RECT 82.735 170.395 86.635 171.075 ;
        RECT 86.645 170.395 93.955 171.075 ;
        RECT 85.705 170.165 86.635 170.395 ;
        RECT 90.160 170.175 91.070 170.395 ;
        RECT 92.605 170.165 93.955 170.395 ;
        RECT 94.005 170.265 95.835 171.075 ;
        RECT 96.305 170.295 97.675 171.075 ;
        RECT 97.845 170.255 99.775 171.075 ;
        RECT 98.825 170.165 99.775 170.255 ;
        RECT 99.995 170.205 100.425 170.990 ;
        RECT 100.445 170.395 104.345 171.075 ;
        RECT 105.045 170.395 108.945 171.075 ;
        RECT 100.445 170.165 101.375 170.395 ;
        RECT 105.045 170.165 105.975 170.395 ;
        RECT 109.185 170.265 111.935 171.075 ;
        RECT 111.945 170.395 115.845 171.075 ;
        RECT 111.945 170.165 112.875 170.395 ;
        RECT 117.005 170.295 118.375 171.075 ;
        RECT 118.385 170.395 125.695 171.075 ;
        RECT 121.900 170.175 122.810 170.395 ;
        RECT 124.345 170.165 125.695 170.395 ;
        RECT 125.755 170.205 126.185 170.990 ;
        RECT 126.205 170.165 129.415 171.075 ;
        RECT 129.425 170.165 132.635 171.075 ;
        RECT 132.645 170.265 138.155 171.075 ;
        RECT 138.175 170.165 139.525 171.075 ;
        RECT 139.545 170.265 141.375 171.075 ;
        RECT 141.385 170.395 143.675 171.075 ;
        RECT 142.755 170.165 143.675 170.395 ;
        RECT 143.685 170.265 149.195 171.075 ;
        RECT 149.205 170.265 151.035 171.075 ;
        RECT 151.515 170.205 151.945 170.990 ;
        RECT 152.060 170.395 155.525 171.075 ;
        RECT 152.060 170.165 152.980 170.395 ;
        RECT 155.645 170.265 157.015 171.075 ;
      LAYER nwell ;
        RECT 22.510 167.045 157.210 169.875 ;
      LAYER pwell ;
        RECT 22.705 165.845 24.075 166.655 ;
        RECT 24.085 165.845 29.595 166.655 ;
        RECT 29.605 165.845 31.435 166.655 ;
        RECT 31.905 166.525 33.040 166.755 ;
        RECT 31.905 165.845 35.115 166.525 ;
        RECT 35.595 165.930 36.025 166.715 ;
        RECT 37.850 166.555 38.795 166.755 ;
        RECT 36.045 165.875 38.795 166.555 ;
        RECT 22.845 165.635 23.015 165.845 ;
        RECT 24.225 165.635 24.395 165.845 ;
        RECT 29.745 165.655 29.915 165.845 ;
        RECT 29.745 165.635 29.910 165.655 ;
        RECT 30.205 165.635 30.375 165.825 ;
        RECT 31.580 165.685 31.700 165.795 ;
        RECT 33.885 165.635 34.055 165.825 ;
        RECT 34.805 165.655 34.975 165.845 ;
        RECT 35.265 165.795 35.435 165.825 ;
        RECT 35.260 165.685 35.435 165.795 ;
        RECT 35.265 165.635 35.435 165.685 ;
        RECT 36.190 165.655 36.360 165.875 ;
        RECT 37.850 165.845 38.795 165.875 ;
        RECT 38.805 165.845 42.475 166.655 ;
        RECT 42.495 165.845 45.225 166.755 ;
        RECT 45.245 166.555 46.200 166.755 ;
        RECT 45.245 165.875 47.525 166.555 ;
        RECT 51.060 166.525 51.970 166.745 ;
        RECT 53.505 166.525 54.855 166.755 ;
        RECT 45.245 165.845 46.200 165.875 ;
        RECT 36.645 165.635 36.815 165.825 ;
        RECT 38.945 165.655 39.115 165.845 ;
        RECT 42.165 165.635 42.335 165.825 ;
        RECT 44.000 165.685 44.120 165.795 ;
        RECT 44.460 165.635 44.630 165.825 ;
        RECT 44.925 165.655 45.095 165.845 ;
        RECT 47.230 165.655 47.400 165.875 ;
        RECT 47.545 165.845 54.855 166.525 ;
        RECT 54.905 166.525 55.825 166.755 ;
        RECT 57.300 166.525 58.220 166.755 ;
        RECT 54.905 165.845 57.195 166.525 ;
        RECT 57.300 165.845 60.765 166.525 ;
        RECT 61.355 165.930 61.785 166.715 ;
        RECT 65.780 166.525 66.690 166.745 ;
        RECT 68.225 166.525 69.575 166.755 ;
        RECT 62.265 165.845 69.575 166.525 ;
        RECT 70.640 166.525 71.560 166.755 ;
        RECT 74.225 166.525 75.155 166.755 ;
        RECT 70.640 165.845 74.105 166.525 ;
        RECT 74.225 165.845 78.125 166.525 ;
        RECT 78.365 165.845 79.735 166.655 ;
        RECT 81.115 166.555 82.470 166.755 ;
        RECT 85.945 166.665 86.895 166.755 ;
        RECT 79.790 166.525 82.470 166.555 ;
        RECT 79.790 165.875 82.955 166.525 ;
        RECT 81.115 165.845 82.955 165.875 ;
        RECT 82.965 165.845 84.795 166.655 ;
        RECT 84.965 165.845 86.895 166.665 ;
        RECT 87.115 165.930 87.545 166.715 ;
        RECT 87.565 165.845 89.775 166.755 ;
        RECT 90.770 166.525 92.140 166.755 ;
        RECT 89.865 165.845 92.140 166.525 ;
        RECT 92.165 165.845 95.835 166.655 ;
        RECT 99.360 166.525 100.270 166.745 ;
        RECT 101.805 166.525 103.155 166.755 ;
        RECT 95.845 165.845 103.155 166.525 ;
        RECT 103.220 166.525 104.590 166.755 ;
        RECT 106.410 166.525 107.780 166.755 ;
        RECT 103.220 165.845 105.495 166.525 ;
        RECT 105.505 165.845 107.780 166.525 ;
        RECT 107.805 165.845 110.015 166.755 ;
        RECT 110.105 165.845 112.855 166.655 ;
        RECT 112.875 165.930 113.305 166.715 ;
        RECT 113.325 165.845 116.995 166.655 ;
        RECT 117.925 166.525 118.855 166.755 ;
        RECT 117.925 165.845 121.825 166.525 ;
        RECT 122.065 165.845 127.575 166.655 ;
        RECT 127.585 165.845 131.255 166.655 ;
        RECT 131.725 165.845 133.075 166.755 ;
        RECT 133.115 165.845 135.845 166.755 ;
        RECT 135.865 165.845 137.235 166.625 ;
        RECT 137.245 165.845 138.615 166.655 ;
        RECT 138.635 165.930 139.065 166.715 ;
        RECT 139.085 165.845 140.455 166.625 ;
        RECT 140.465 165.845 145.975 166.655 ;
        RECT 145.985 165.845 147.355 166.655 ;
        RECT 150.880 166.525 151.790 166.745 ;
        RECT 153.325 166.525 154.675 166.755 ;
        RECT 147.365 165.845 154.675 166.525 ;
        RECT 155.645 165.845 157.015 166.655 ;
        RECT 47.685 165.655 47.855 165.845 ;
        RECT 48.140 165.635 48.310 165.825 ;
        RECT 51.360 165.635 51.530 165.825 ;
        RECT 55.045 165.635 55.215 165.825 ;
        RECT 55.505 165.635 55.675 165.825 ;
        RECT 56.885 165.655 57.055 165.845 ;
        RECT 60.565 165.655 60.735 165.845 ;
        RECT 61.020 165.685 61.140 165.795 ;
        RECT 61.940 165.685 62.060 165.795 ;
        RECT 62.405 165.655 62.575 165.845 ;
        RECT 64.245 165.635 64.415 165.825 ;
        RECT 64.700 165.685 64.820 165.795 ;
        RECT 65.165 165.635 65.335 165.825 ;
        RECT 67.935 165.680 68.095 165.790 ;
        RECT 69.775 165.690 69.935 165.800 ;
        RECT 70.685 165.635 70.855 165.825 ;
        RECT 71.145 165.655 71.315 165.825 ;
        RECT 73.455 165.680 73.615 165.790 ;
        RECT 73.905 165.655 74.075 165.845 ;
        RECT 74.640 165.655 74.810 165.845 ;
        RECT 78.505 165.825 78.675 165.845 ;
        RECT 71.165 165.635 71.315 165.655 ;
        RECT 74.825 165.635 74.995 165.825 ;
        RECT 76.205 165.635 76.375 165.825 ;
        RECT 78.040 165.685 78.160 165.795 ;
        RECT 78.505 165.655 78.680 165.825 ;
        RECT 82.645 165.655 82.815 165.845 ;
        RECT 83.105 165.655 83.275 165.845 ;
        RECT 84.965 165.825 85.115 165.845 ;
        RECT 84.945 165.655 85.115 165.825 ;
        RECT 85.860 165.685 85.980 165.795 ;
        RECT 87.710 165.655 87.880 165.845 ;
        RECT 78.510 165.635 78.680 165.655 ;
        RECT 22.705 164.825 24.075 165.635 ;
        RECT 24.085 164.825 27.755 165.635 ;
        RECT 28.075 164.955 29.910 165.635 ;
        RECT 28.075 164.725 29.005 164.955 ;
        RECT 30.065 164.825 33.735 165.635 ;
        RECT 33.745 164.825 35.115 165.635 ;
        RECT 35.135 164.725 36.485 165.635 ;
        RECT 36.505 164.825 42.015 165.635 ;
        RECT 42.025 164.825 43.855 165.635 ;
        RECT 44.345 164.725 45.695 165.635 ;
        RECT 45.845 164.725 48.455 165.635 ;
        RECT 48.475 164.765 48.905 165.550 ;
        RECT 49.065 164.725 51.675 165.635 ;
        RECT 51.780 164.955 55.245 165.635 ;
        RECT 51.780 164.725 52.700 164.955 ;
        RECT 55.365 164.825 57.195 165.635 ;
        RECT 57.245 164.955 64.555 165.635 ;
        RECT 57.245 164.725 58.595 164.955 ;
        RECT 60.130 164.735 61.040 164.955 ;
        RECT 65.035 164.725 67.765 165.635 ;
        RECT 68.705 164.955 70.995 165.635 ;
        RECT 68.705 164.725 69.625 164.955 ;
        RECT 71.165 164.815 73.095 165.635 ;
        RECT 72.145 164.725 73.095 164.815 ;
        RECT 74.235 164.765 74.665 165.550 ;
        RECT 74.685 164.855 76.055 165.635 ;
        RECT 76.065 164.825 77.895 165.635 ;
        RECT 78.365 164.725 85.475 165.635 ;
        RECT 86.190 165.605 87.595 165.635 ;
        RECT 89.085 165.605 89.255 165.825 ;
        RECT 89.545 165.635 89.715 165.825 ;
        RECT 90.010 165.655 90.180 165.845 ;
        RECT 92.305 165.655 92.475 165.845 ;
        RECT 94.610 165.635 94.780 165.825 ;
        RECT 95.985 165.655 96.155 165.845 ;
        RECT 97.825 165.655 97.995 165.825 ;
        RECT 97.830 165.635 97.995 165.655 ;
        RECT 100.585 165.635 100.755 165.825 ;
        RECT 102.425 165.635 102.595 165.825 ;
        RECT 105.180 165.655 105.350 165.845 ;
        RECT 105.650 165.825 105.820 165.845 ;
        RECT 105.645 165.655 105.820 165.825 ;
        RECT 107.495 165.680 107.655 165.790 ;
        RECT 107.950 165.655 108.120 165.845 ;
        RECT 105.645 165.635 105.815 165.655 ;
        RECT 109.325 165.635 109.495 165.825 ;
        RECT 109.785 165.635 109.955 165.825 ;
        RECT 110.245 165.655 110.415 165.845 ;
        RECT 113.465 165.795 113.635 165.845 ;
        RECT 113.460 165.685 113.635 165.795 ;
        RECT 113.465 165.655 113.635 165.685 ;
        RECT 113.925 165.635 114.095 165.825 ;
        RECT 117.155 165.690 117.315 165.800 ;
        RECT 118.340 165.655 118.510 165.845 ;
        RECT 121.285 165.635 121.455 165.825 ;
        RECT 122.205 165.655 122.375 165.845 ;
        RECT 124.975 165.680 125.135 165.790 ;
        RECT 126.345 165.635 126.515 165.825 ;
        RECT 127.725 165.655 127.895 165.845 ;
        RECT 129.110 165.635 129.280 165.825 ;
        RECT 130.945 165.635 131.115 165.825 ;
        RECT 131.400 165.685 131.520 165.795 ;
        RECT 132.790 165.655 132.960 165.845 ;
        RECT 134.165 165.635 134.335 165.825 ;
        RECT 135.545 165.655 135.715 165.845 ;
        RECT 136.005 165.655 136.175 165.845 ;
        RECT 137.385 165.655 137.555 165.845 ;
        RECT 139.225 165.655 139.395 165.845 ;
        RECT 140.605 165.655 140.775 165.845 ;
        RECT 143.365 165.635 143.535 165.825 ;
        RECT 143.825 165.635 143.995 165.825 ;
        RECT 146.125 165.655 146.295 165.845 ;
        RECT 147.505 165.655 147.675 165.845 ;
        RECT 149.345 165.635 149.515 165.825 ;
        RECT 151.180 165.685 151.300 165.795 ;
        RECT 152.105 165.635 152.275 165.825 ;
        RECT 154.875 165.690 155.035 165.800 ;
        RECT 156.705 165.635 156.875 165.845 ;
        RECT 86.190 164.925 89.395 165.605 ;
        RECT 89.405 164.955 94.220 165.635 ;
        RECT 94.610 165.405 97.665 165.635 ;
        RECT 86.190 164.725 87.595 164.925 ;
        RECT 94.465 164.725 97.665 165.405 ;
        RECT 97.830 164.955 99.665 165.635 ;
        RECT 98.735 164.725 99.665 164.955 ;
        RECT 99.995 164.765 100.425 165.550 ;
        RECT 100.445 164.955 102.275 165.635 ;
        RECT 100.930 164.725 102.275 164.955 ;
        RECT 102.285 164.825 105.035 165.635 ;
        RECT 105.505 164.955 107.335 165.635 ;
        RECT 105.990 164.725 107.335 164.955 ;
        RECT 108.275 164.725 109.625 165.635 ;
        RECT 109.645 164.825 113.315 165.635 ;
        RECT 113.785 164.955 121.095 165.635 ;
        RECT 121.255 164.955 124.720 165.635 ;
        RECT 117.300 164.735 118.210 164.955 ;
        RECT 119.745 164.725 121.095 164.955 ;
        RECT 123.800 164.725 124.720 164.955 ;
        RECT 125.755 164.765 126.185 165.550 ;
        RECT 126.205 164.825 128.955 165.635 ;
        RECT 128.965 164.725 130.795 165.635 ;
        RECT 130.805 164.955 134.015 165.635 ;
        RECT 134.025 164.955 136.315 165.635 ;
        RECT 132.880 164.725 134.015 164.955 ;
        RECT 135.395 164.725 136.315 164.955 ;
        RECT 136.365 164.955 143.675 165.635 ;
        RECT 136.365 164.725 137.715 164.955 ;
        RECT 139.250 164.735 140.160 164.955 ;
        RECT 143.685 164.825 149.195 165.635 ;
        RECT 149.205 164.825 151.035 165.635 ;
        RECT 151.515 164.765 151.945 165.550 ;
        RECT 151.965 164.825 155.635 165.635 ;
        RECT 155.645 164.825 157.015 165.635 ;
      LAYER nwell ;
        RECT 22.510 161.605 157.210 164.435 ;
      LAYER pwell ;
        RECT 22.705 160.405 24.075 161.215 ;
        RECT 27.600 161.085 28.510 161.305 ;
        RECT 30.045 161.085 31.395 161.315 ;
        RECT 24.085 160.405 31.395 161.085 ;
        RECT 31.445 161.115 32.375 161.315 ;
        RECT 33.705 161.115 34.655 161.315 ;
        RECT 31.445 160.635 34.655 161.115 ;
        RECT 31.590 160.435 34.655 160.635 ;
        RECT 35.595 160.490 36.025 161.275 ;
        RECT 39.560 161.085 40.470 161.305 ;
        RECT 42.005 161.085 43.355 161.315 ;
        RECT 22.845 160.195 23.015 160.405 ;
        RECT 24.225 160.355 24.395 160.405 ;
        RECT 24.220 160.245 24.395 160.355 ;
        RECT 24.225 160.215 24.395 160.245 ;
        RECT 25.605 160.195 25.775 160.385 ;
        RECT 27.905 160.195 28.075 160.385 ;
        RECT 31.590 160.215 31.760 160.435 ;
        RECT 33.720 160.405 34.655 160.435 ;
        RECT 36.045 160.405 43.355 161.085 ;
        RECT 43.405 161.085 44.325 161.315 ;
        RECT 43.405 160.405 45.695 161.085 ;
        RECT 46.635 160.405 49.365 161.315 ;
        RECT 49.385 160.405 52.595 161.315 ;
        RECT 55.260 161.085 56.180 161.315 ;
        RECT 58.940 161.085 59.860 161.315 ;
        RECT 52.715 160.405 56.180 161.085 ;
        RECT 56.395 160.405 59.860 161.085 ;
        RECT 59.965 160.405 61.335 161.215 ;
        RECT 61.355 160.490 61.785 161.275 ;
        RECT 61.805 161.085 62.725 161.315 ;
        RECT 61.805 160.405 64.095 161.085 ;
        RECT 64.105 160.405 69.615 161.215 ;
        RECT 70.585 161.085 71.935 161.315 ;
        RECT 73.470 161.085 74.380 161.305 ;
        RECT 70.585 160.405 77.895 161.085 ;
        RECT 77.905 160.405 79.735 161.215 ;
        RECT 79.985 160.405 87.095 161.315 ;
        RECT 87.115 160.490 87.545 161.275 ;
        RECT 87.565 161.085 88.495 161.315 ;
        RECT 87.565 160.405 91.465 161.085 ;
        RECT 92.265 160.405 94.455 161.315 ;
        RECT 94.465 160.405 99.975 161.215 ;
        RECT 100.930 161.085 102.275 161.315 ;
        RECT 109.020 161.085 109.930 161.305 ;
        RECT 111.465 161.085 112.815 161.315 ;
        RECT 100.445 160.405 102.275 161.085 ;
        RECT 102.285 160.405 105.025 161.085 ;
        RECT 105.505 160.405 112.815 161.085 ;
        RECT 112.875 160.490 113.305 161.275 ;
        RECT 113.420 161.085 114.340 161.315 ;
        RECT 117.560 161.085 118.480 161.315 ;
        RECT 113.420 160.405 116.885 161.085 ;
        RECT 117.560 160.405 121.025 161.085 ;
        RECT 121.145 160.405 124.355 161.315 ;
        RECT 125.285 160.405 128.940 161.315 ;
        RECT 128.965 160.405 130.795 161.215 ;
        RECT 130.815 160.405 132.165 161.315 ;
        RECT 132.185 160.405 133.555 161.215 ;
        RECT 133.565 161.115 134.495 161.315 ;
        RECT 135.825 161.115 136.775 161.315 ;
        RECT 133.565 160.635 136.775 161.115 ;
        RECT 133.710 160.435 136.775 160.635 ;
        RECT 32.965 160.195 33.135 160.385 ;
        RECT 33.425 160.195 33.595 160.385 ;
        RECT 34.815 160.355 34.975 160.360 ;
        RECT 34.800 160.250 34.975 160.355 ;
        RECT 34.800 160.245 34.920 160.250 ;
        RECT 36.185 160.195 36.355 160.405 ;
        RECT 36.645 160.195 36.815 160.385 ;
        RECT 22.705 159.385 24.075 160.195 ;
        RECT 24.545 159.415 25.915 160.195 ;
        RECT 25.925 159.515 28.215 160.195 ;
        RECT 28.460 159.515 33.275 160.195 ;
        RECT 25.925 159.285 26.845 159.515 ;
        RECT 33.285 159.415 34.655 160.195 ;
        RECT 35.135 159.285 36.485 160.195 ;
        RECT 36.505 159.385 38.335 160.195 ;
        RECT 38.490 160.165 38.660 160.385 ;
        RECT 44.005 160.215 44.175 160.385 ;
        RECT 45.385 160.215 45.555 160.405 ;
        RECT 45.855 160.250 46.015 160.360 ;
        RECT 46.765 160.215 46.935 160.405 ;
        RECT 44.005 160.195 44.075 160.215 ;
        RECT 47.225 160.195 47.395 160.385 ;
        RECT 47.695 160.240 47.855 160.350 ;
        RECT 49.075 160.240 49.235 160.350 ;
        RECT 52.285 160.215 52.455 160.405 ;
        RECT 52.745 160.215 52.915 160.405 ;
        RECT 54.585 160.195 54.755 160.385 ;
        RECT 56.425 160.215 56.595 160.405 ;
        RECT 60.105 160.215 60.275 160.405 ;
        RECT 61.945 160.195 62.115 160.385 ;
        RECT 62.405 160.195 62.575 160.385 ;
        RECT 63.785 160.215 63.955 160.405 ;
        RECT 64.245 160.215 64.415 160.405 ;
        RECT 64.705 160.195 64.875 160.385 ;
        RECT 68.380 160.195 68.550 160.385 ;
        RECT 68.845 160.195 69.015 160.385 ;
        RECT 69.775 160.250 69.935 160.360 ;
        RECT 70.685 160.215 70.855 160.385 ;
        RECT 70.705 160.195 70.855 160.215 ;
        RECT 73.905 160.195 74.075 160.385 ;
        RECT 74.820 160.245 74.940 160.355 ;
        RECT 75.560 160.195 75.730 160.385 ;
        RECT 77.585 160.215 77.755 160.405 ;
        RECT 78.045 160.215 78.215 160.405 ;
        RECT 86.780 160.385 86.950 160.405 ;
        RECT 79.425 160.195 79.595 160.385 ;
        RECT 81.725 160.195 81.895 160.385 ;
        RECT 83.105 160.195 83.275 160.385 ;
        RECT 84.485 160.215 84.655 160.385 ;
        RECT 86.780 160.215 86.955 160.385 ;
        RECT 87.980 160.215 88.150 160.405 ;
        RECT 91.840 160.245 91.960 160.355 ;
        RECT 94.140 160.350 94.310 160.405 ;
        RECT 94.140 160.240 94.315 160.350 ;
        RECT 94.140 160.215 94.310 160.240 ;
        RECT 94.605 160.215 94.775 160.405 ;
        RECT 84.505 160.195 84.655 160.215 ;
        RECT 86.785 160.195 86.955 160.215 ;
        RECT 95.065 160.195 95.235 160.385 ;
        RECT 97.825 160.195 97.995 160.385 ;
        RECT 100.585 160.355 100.755 160.405 ;
        RECT 99.660 160.245 99.780 160.355 ;
        RECT 100.120 160.245 100.240 160.355 ;
        RECT 100.580 160.245 100.755 160.355 ;
        RECT 100.585 160.215 100.755 160.245 ;
        RECT 101.040 160.195 101.210 160.385 ;
        RECT 102.425 160.195 102.595 160.405 ;
        RECT 104.260 160.245 104.380 160.355 ;
        RECT 104.730 160.195 104.900 160.385 ;
        RECT 105.180 160.245 105.300 160.355 ;
        RECT 105.645 160.215 105.815 160.405 ;
        RECT 109.785 160.195 109.955 160.385 ;
        RECT 110.245 160.195 110.415 160.385 ;
        RECT 112.085 160.195 112.255 160.385 ;
        RECT 115.305 160.195 115.475 160.385 ;
        RECT 116.685 160.215 116.855 160.405 ;
        RECT 117.140 160.245 117.260 160.355 ;
        RECT 120.825 160.215 120.995 160.405 ;
        RECT 40.150 160.165 41.095 160.195 ;
        RECT 38.345 159.485 41.095 160.165 ;
        RECT 41.805 159.965 44.075 160.195 ;
        RECT 40.150 159.285 41.095 159.485 ;
        RECT 41.320 159.285 44.075 159.965 ;
        RECT 44.325 159.285 47.535 160.195 ;
        RECT 48.475 159.325 48.905 160.110 ;
        RECT 50.080 159.515 54.895 160.195 ;
        RECT 54.945 159.515 62.255 160.195 ;
        RECT 62.265 159.515 64.555 160.195 ;
        RECT 54.945 159.285 56.295 159.515 ;
        RECT 57.830 159.295 58.740 159.515 ;
        RECT 63.635 159.285 64.555 159.515 ;
        RECT 64.565 159.385 66.395 160.195 ;
        RECT 66.420 159.515 68.695 160.195 ;
        RECT 66.420 159.285 67.790 159.515 ;
        RECT 68.705 159.385 70.535 160.195 ;
        RECT 70.705 159.375 72.635 160.195 ;
        RECT 72.845 159.415 74.215 160.195 ;
        RECT 71.685 159.285 72.635 159.375 ;
        RECT 74.235 159.325 74.665 160.110 ;
        RECT 75.145 159.515 79.045 160.195 ;
        RECT 79.285 159.515 81.575 160.195 ;
        RECT 75.145 159.285 76.075 159.515 ;
        RECT 80.655 159.285 81.575 159.515 ;
        RECT 81.595 159.285 82.945 160.195 ;
        RECT 82.965 159.385 84.335 160.195 ;
        RECT 84.505 159.375 86.435 160.195 ;
        RECT 86.645 159.515 93.955 160.195 ;
        RECT 85.485 159.285 86.435 159.375 ;
        RECT 90.160 159.295 91.070 159.515 ;
        RECT 92.605 159.285 93.955 159.515 ;
        RECT 94.935 159.285 97.665 160.195 ;
        RECT 97.685 159.385 99.515 160.195 ;
        RECT 99.995 159.325 100.425 160.110 ;
        RECT 100.925 159.285 102.275 160.195 ;
        RECT 102.285 159.385 104.115 160.195 ;
        RECT 104.585 159.285 106.795 160.195 ;
        RECT 106.885 159.285 110.095 160.195 ;
        RECT 110.105 159.385 111.935 160.195 ;
        RECT 111.945 159.285 115.155 160.195 ;
        RECT 115.165 159.515 122.475 160.195 ;
        RECT 122.670 160.165 122.840 160.385 ;
        RECT 124.045 160.215 124.215 160.405 ;
        RECT 124.515 160.250 124.675 160.360 ;
        RECT 125.430 160.355 125.600 160.405 ;
        RECT 125.420 160.245 125.600 160.355 ;
        RECT 125.430 160.215 125.600 160.245 ;
        RECT 128.645 160.195 128.815 160.385 ;
        RECT 129.105 160.215 129.275 160.405 ;
        RECT 130.945 160.215 131.115 160.405 ;
        RECT 131.405 160.195 131.575 160.385 ;
        RECT 132.325 160.215 132.495 160.405 ;
        RECT 132.785 160.195 132.955 160.385 ;
        RECT 133.245 160.195 133.415 160.385 ;
        RECT 133.710 160.215 133.880 160.435 ;
        RECT 135.840 160.405 136.775 160.435 ;
        RECT 136.785 160.405 138.615 161.215 ;
        RECT 138.635 160.490 139.065 161.275 ;
        RECT 139.125 161.085 140.475 161.315 ;
        RECT 142.010 161.085 142.920 161.305 ;
        RECT 149.960 161.085 150.870 161.305 ;
        RECT 152.405 161.085 153.755 161.315 ;
        RECT 139.125 160.405 146.435 161.085 ;
        RECT 146.445 160.405 153.755 161.085 ;
        RECT 153.805 160.405 155.635 161.215 ;
        RECT 155.645 160.405 157.015 161.215 ;
        RECT 136.000 160.245 136.120 160.355 ;
        RECT 136.465 160.195 136.635 160.385 ;
        RECT 136.925 160.215 137.095 160.405 ;
        RECT 138.765 160.195 138.935 160.385 ;
        RECT 142.455 160.240 142.615 160.350 ;
        RECT 143.365 160.195 143.535 160.385 ;
        RECT 146.125 160.215 146.295 160.405 ;
        RECT 146.585 160.355 146.755 160.405 ;
        RECT 146.580 160.245 146.755 160.355 ;
        RECT 146.585 160.215 146.755 160.245 ;
        RECT 147.040 160.195 147.210 160.385 ;
        RECT 148.425 160.195 148.595 160.385 ;
        RECT 151.180 160.245 151.300 160.355 ;
        RECT 153.945 160.215 154.115 160.405 ;
        RECT 155.325 160.195 155.495 160.385 ;
        RECT 156.705 160.195 156.875 160.405 ;
        RECT 124.330 160.165 125.275 160.195 ;
        RECT 118.680 159.295 119.590 159.515 ;
        RECT 121.125 159.285 122.475 159.515 ;
        RECT 122.525 159.485 125.275 160.165 ;
        RECT 124.330 159.285 125.275 159.485 ;
        RECT 125.755 159.325 126.185 160.110 ;
        RECT 126.205 159.515 128.955 160.195 ;
        RECT 128.965 159.515 131.715 160.195 ;
        RECT 126.205 159.285 127.135 159.515 ;
        RECT 128.965 159.285 129.895 159.515 ;
        RECT 131.735 159.285 133.085 160.195 ;
        RECT 133.105 159.385 135.855 160.195 ;
        RECT 136.325 159.515 138.615 160.195 ;
        RECT 137.695 159.285 138.615 159.515 ;
        RECT 138.625 159.385 142.295 160.195 ;
        RECT 143.325 159.285 146.435 160.195 ;
        RECT 146.925 159.285 148.275 160.195 ;
        RECT 148.285 159.385 151.035 160.195 ;
        RECT 151.515 159.325 151.945 160.110 ;
        RECT 152.060 159.515 155.525 160.195 ;
        RECT 152.060 159.285 152.980 159.515 ;
        RECT 155.645 159.385 157.015 160.195 ;
      LAYER nwell ;
        RECT 22.510 156.165 157.210 158.995 ;
      LAYER pwell ;
        RECT 22.705 154.965 24.075 155.775 ;
        RECT 24.085 154.965 27.755 155.775 ;
        RECT 28.225 155.645 29.145 155.875 ;
        RECT 28.225 154.965 30.515 155.645 ;
        RECT 30.525 154.965 31.875 155.875 ;
        RECT 31.925 154.965 33.275 155.875 ;
        RECT 33.285 154.965 34.635 155.875 ;
        RECT 35.595 155.050 36.025 155.835 ;
        RECT 36.045 154.965 37.875 155.775 ;
        RECT 39.690 155.675 40.635 155.875 ;
        RECT 37.885 154.995 40.635 155.675 ;
        RECT 22.845 154.755 23.015 154.965 ;
        RECT 24.225 154.755 24.395 154.965 ;
        RECT 27.900 154.805 28.020 154.915 ;
        RECT 30.205 154.775 30.375 154.965 ;
        RECT 31.590 154.775 31.760 154.965 ;
        RECT 32.040 154.775 32.210 154.965 ;
        RECT 33.425 154.775 33.595 154.945 ;
        RECT 33.425 154.755 33.590 154.775 ;
        RECT 33.885 154.755 34.055 154.945 ;
        RECT 34.350 154.775 34.520 154.965 ;
        RECT 34.815 154.810 34.975 154.920 ;
        RECT 35.265 154.755 35.435 154.945 ;
        RECT 36.185 154.775 36.355 154.965 ;
        RECT 38.030 154.945 38.200 154.995 ;
        RECT 39.690 154.965 40.635 154.995 ;
        RECT 41.585 154.965 42.935 155.875 ;
        RECT 43.405 154.965 46.155 155.875 ;
        RECT 46.165 154.965 47.995 155.775 ;
        RECT 51.520 155.645 52.430 155.865 ;
        RECT 53.965 155.645 55.315 155.875 ;
        RECT 48.005 154.965 55.315 155.645 ;
        RECT 55.365 154.965 57.195 155.775 ;
        RECT 57.215 154.965 59.945 155.875 ;
        RECT 59.965 154.965 61.335 155.775 ;
        RECT 61.355 155.050 61.785 155.835 ;
        RECT 61.845 155.645 63.195 155.875 ;
        RECT 64.730 155.645 65.640 155.865 ;
        RECT 73.140 155.645 74.050 155.865 ;
        RECT 75.585 155.645 76.935 155.875 ;
        RECT 61.845 154.965 69.155 155.645 ;
        RECT 69.625 154.965 76.935 155.645 ;
        RECT 76.985 154.965 82.495 155.775 ;
        RECT 82.505 154.965 86.175 155.775 ;
        RECT 87.115 155.050 87.545 155.835 ;
        RECT 87.565 154.965 88.935 155.745 ;
        RECT 89.865 154.965 91.235 155.745 ;
        RECT 94.760 155.645 95.670 155.865 ;
        RECT 97.205 155.645 98.555 155.875 ;
        RECT 91.245 154.965 98.555 155.645 ;
        RECT 99.565 155.645 100.915 155.875 ;
        RECT 102.450 155.645 103.360 155.865 ;
        RECT 99.565 154.965 106.875 155.645 ;
        RECT 107.805 154.965 110.015 155.875 ;
        RECT 110.105 154.965 112.855 155.775 ;
        RECT 112.875 155.050 113.305 155.835 ;
        RECT 113.420 155.645 114.340 155.875 ;
        RECT 113.420 154.965 116.885 155.645 ;
        RECT 117.005 154.965 120.215 155.875 ;
        RECT 123.800 155.645 124.720 155.875 ;
        RECT 121.255 154.965 124.720 155.645 ;
        RECT 124.825 154.965 128.035 155.875 ;
        RECT 128.045 154.965 131.255 155.875 ;
        RECT 131.275 154.965 134.005 155.875 ;
        RECT 135.995 155.645 136.925 155.875 ;
        RECT 135.090 154.965 136.925 155.645 ;
        RECT 137.265 154.965 138.615 155.875 ;
        RECT 138.635 155.050 139.065 155.835 ;
        RECT 139.545 154.965 140.915 155.745 ;
        RECT 140.965 155.645 142.315 155.875 ;
        RECT 143.850 155.645 144.760 155.865 ;
        RECT 140.965 154.965 148.275 155.645 ;
        RECT 148.285 154.965 149.655 155.775 ;
        RECT 149.665 154.965 154.480 155.645 ;
        RECT 155.645 154.965 157.015 155.775 ;
        RECT 36.645 154.755 36.815 154.945 ;
        RECT 38.025 154.775 38.200 154.945 ;
        RECT 40.795 154.810 40.955 154.920 ;
        RECT 38.025 154.755 38.195 154.775 ;
        RECT 41.245 154.755 41.415 154.945 ;
        RECT 41.700 154.775 41.870 154.965 ;
        RECT 43.085 154.915 43.255 154.945 ;
        RECT 43.080 154.805 43.255 154.915 ;
        RECT 43.085 154.755 43.255 154.805 ;
        RECT 43.545 154.775 43.715 154.965 ;
        RECT 45.845 154.755 46.015 154.945 ;
        RECT 46.305 154.775 46.475 154.965 ;
        RECT 48.145 154.775 48.315 154.965 ;
        RECT 49.060 154.805 49.180 154.915 ;
        RECT 49.525 154.755 49.695 154.945 ;
        RECT 55.505 154.775 55.675 154.965 ;
        RECT 56.885 154.755 57.055 154.945 ;
        RECT 58.725 154.755 58.895 154.945 ;
        RECT 59.645 154.775 59.815 154.965 ;
        RECT 60.105 154.775 60.275 154.965 ;
        RECT 62.400 154.805 62.520 154.915 ;
        RECT 65.165 154.755 65.335 154.945 ;
        RECT 65.635 154.800 65.795 154.910 ;
        RECT 68.380 154.755 68.550 154.945 ;
        RECT 68.845 154.755 69.015 154.965 ;
        RECT 69.300 154.805 69.420 154.915 ;
        RECT 69.765 154.775 69.935 154.965 ;
        RECT 77.125 154.775 77.295 154.965 ;
        RECT 78.230 154.755 78.400 154.945 ;
        RECT 78.970 154.755 79.140 154.945 ;
        RECT 81.265 154.755 81.435 154.945 ;
        RECT 82.645 154.775 82.815 154.965 ;
        RECT 84.485 154.755 84.655 154.945 ;
        RECT 86.335 154.810 86.495 154.920 ;
        RECT 87.705 154.775 87.875 154.965 ;
        RECT 88.165 154.755 88.335 154.945 ;
        RECT 89.095 154.810 89.255 154.920 ;
        RECT 89.545 154.755 89.715 154.945 ;
        RECT 90.005 154.775 90.175 154.965 ;
        RECT 91.385 154.775 91.555 154.965 ;
        RECT 93.225 154.755 93.395 154.945 ;
        RECT 93.680 154.805 93.800 154.915 ;
        RECT 22.705 153.945 24.075 154.755 ;
        RECT 24.085 154.075 31.395 154.755 ;
        RECT 27.600 153.855 28.510 154.075 ;
        RECT 30.045 153.845 31.395 154.075 ;
        RECT 31.755 154.075 33.590 154.755 ;
        RECT 31.755 153.845 32.685 154.075 ;
        RECT 33.745 153.975 35.115 154.755 ;
        RECT 35.125 153.945 36.495 154.755 ;
        RECT 36.515 153.845 37.865 154.755 ;
        RECT 37.885 153.845 41.095 154.755 ;
        RECT 41.105 153.945 42.935 154.755 ;
        RECT 42.945 153.845 45.665 154.755 ;
        RECT 45.705 153.945 48.455 154.755 ;
        RECT 48.475 153.885 48.905 154.670 ;
        RECT 49.385 154.075 56.695 154.755 ;
        RECT 52.900 153.855 53.810 154.075 ;
        RECT 55.345 153.845 56.695 154.075 ;
        RECT 56.745 153.945 58.575 154.755 ;
        RECT 58.695 154.075 62.160 154.755 ;
        RECT 61.240 153.845 62.160 154.075 ;
        RECT 62.735 153.845 65.465 154.755 ;
        RECT 66.485 153.845 68.695 154.755 ;
        RECT 68.705 153.945 74.215 154.755 ;
        RECT 74.235 153.885 74.665 154.670 ;
        RECT 74.915 154.075 78.815 154.755 ;
        RECT 77.885 153.845 78.815 154.075 ;
        RECT 78.825 153.845 81.035 154.755 ;
        RECT 81.125 153.945 82.495 154.755 ;
        RECT 82.505 154.075 84.795 154.755 ;
        RECT 84.900 154.075 88.365 154.755 ;
        RECT 82.505 153.845 83.425 154.075 ;
        RECT 84.900 153.845 85.820 154.075 ;
        RECT 88.495 153.845 89.845 154.755 ;
        RECT 89.960 154.075 93.425 154.755 ;
        RECT 94.005 154.725 94.940 154.755 ;
        RECT 96.900 154.725 97.070 154.945 ;
        RECT 97.360 154.805 97.480 154.915 ;
        RECT 97.825 154.755 97.995 154.945 ;
        RECT 98.755 154.810 98.915 154.920 ;
        RECT 100.580 154.805 100.700 154.915 ;
        RECT 101.045 154.755 101.215 154.945 ;
        RECT 104.725 154.755 104.895 154.945 ;
        RECT 106.565 154.755 106.735 154.965 ;
        RECT 107.035 154.810 107.195 154.920 ;
        RECT 107.950 154.775 108.120 154.965 ;
        RECT 110.245 154.775 110.415 154.965 ;
        RECT 113.925 154.755 114.095 154.945 ;
        RECT 115.765 154.755 115.935 154.945 ;
        RECT 116.685 154.775 116.855 154.965 ;
        RECT 119.905 154.775 120.075 154.965 ;
        RECT 120.375 154.810 120.535 154.920 ;
        RECT 121.285 154.775 121.455 154.965 ;
        RECT 123.125 154.755 123.295 154.945 ;
        RECT 126.345 154.755 126.515 154.945 ;
        RECT 127.725 154.775 127.895 154.965 ;
        RECT 129.565 154.755 129.735 154.945 ;
        RECT 130.945 154.775 131.115 154.965 ;
        RECT 132.330 154.755 132.500 154.945 ;
        RECT 133.705 154.775 133.875 154.965 ;
        RECT 135.090 154.945 135.255 154.965 ;
        RECT 134.175 154.810 134.335 154.920 ;
        RECT 134.625 154.755 134.795 154.945 ;
        RECT 135.085 154.775 135.260 154.945 ;
        RECT 137.380 154.775 137.550 154.965 ;
        RECT 139.225 154.915 139.395 154.945 ;
        RECT 139.220 154.805 139.395 154.915 ;
        RECT 94.005 154.525 97.070 154.725 ;
        RECT 89.960 153.845 90.880 154.075 ;
        RECT 94.005 154.045 97.215 154.525 ;
        RECT 97.685 154.075 99.975 154.755 ;
        RECT 94.005 153.845 94.955 154.045 ;
        RECT 96.285 153.845 97.215 154.045 ;
        RECT 99.055 153.845 99.975 154.075 ;
        RECT 99.995 153.885 100.425 154.670 ;
        RECT 101.015 154.075 104.480 154.755 ;
        RECT 103.560 153.845 104.480 154.075 ;
        RECT 104.585 153.945 106.415 154.755 ;
        RECT 106.425 154.075 113.735 154.755 ;
        RECT 109.940 153.855 110.850 154.075 ;
        RECT 112.385 153.845 113.735 154.075 ;
        RECT 113.785 153.945 115.615 154.755 ;
        RECT 115.625 154.075 122.935 154.755 ;
        RECT 119.140 153.855 120.050 154.075 ;
        RECT 121.585 153.845 122.935 154.075 ;
        RECT 122.985 153.945 125.735 154.755 ;
        RECT 125.755 153.885 126.185 154.670 ;
        RECT 126.205 153.845 129.415 154.755 ;
        RECT 129.425 153.945 131.255 154.755 ;
        RECT 131.265 153.845 132.615 154.755 ;
        RECT 132.645 154.075 134.935 154.755 ;
        RECT 135.090 154.725 135.260 154.775 ;
        RECT 139.225 154.755 139.395 154.805 ;
        RECT 139.685 154.755 139.855 154.965 ;
        RECT 147.965 154.755 148.135 154.965 ;
        RECT 148.425 154.755 148.595 154.965 ;
        RECT 149.805 154.775 149.975 154.965 ;
        RECT 151.180 154.805 151.300 154.915 ;
        RECT 152.105 154.755 152.275 154.945 ;
        RECT 154.875 154.810 155.035 154.920 ;
        RECT 156.705 154.755 156.875 154.965 ;
        RECT 137.220 154.725 138.155 154.755 ;
        RECT 135.090 154.525 138.155 154.725 ;
        RECT 132.645 153.845 133.565 154.075 ;
        RECT 134.945 154.045 138.155 154.525 ;
        RECT 134.945 153.845 135.875 154.045 ;
        RECT 137.205 153.845 138.155 154.045 ;
        RECT 138.175 153.845 139.525 154.755 ;
        RECT 139.545 153.975 140.915 154.755 ;
        RECT 140.965 154.075 148.275 154.755 ;
        RECT 140.965 153.845 142.315 154.075 ;
        RECT 143.850 153.855 144.760 154.075 ;
        RECT 148.285 153.945 151.035 154.755 ;
        RECT 151.515 153.885 151.945 154.670 ;
        RECT 151.965 153.945 155.635 154.755 ;
        RECT 155.645 153.945 157.015 154.755 ;
      LAYER nwell ;
        RECT 22.510 150.725 157.210 153.555 ;
      LAYER pwell ;
        RECT 22.705 149.525 24.075 150.335 ;
        RECT 25.005 149.525 26.375 150.305 ;
        RECT 26.385 149.525 28.215 150.335 ;
        RECT 28.705 149.525 30.055 150.435 ;
        RECT 30.065 150.235 30.995 150.435 ;
        RECT 32.325 150.235 33.275 150.435 ;
        RECT 30.065 149.755 33.275 150.235 ;
        RECT 30.210 149.555 33.275 149.755 ;
        RECT 22.845 149.315 23.015 149.525 ;
        RECT 24.225 149.315 24.395 149.505 ;
        RECT 26.065 149.335 26.235 149.525 ;
        RECT 26.525 149.335 26.695 149.525 ;
        RECT 28.360 149.365 28.480 149.475 ;
        RECT 28.820 149.335 28.990 149.525 ;
        RECT 29.745 149.315 29.915 149.505 ;
        RECT 30.210 149.335 30.380 149.555 ;
        RECT 32.340 149.525 33.275 149.555 ;
        RECT 33.285 150.205 34.205 150.435 ;
        RECT 33.285 149.525 35.575 150.205 ;
        RECT 35.595 149.610 36.025 150.395 ;
        RECT 36.055 149.525 37.405 150.435 ;
        RECT 37.425 149.525 39.255 150.335 ;
        RECT 41.530 150.235 42.475 150.435 ;
        RECT 39.725 149.555 42.475 150.235 ;
        RECT 35.265 149.335 35.435 149.525 ;
        RECT 37.105 149.335 37.275 149.525 ;
        RECT 37.565 149.335 37.735 149.525 ;
        RECT 39.870 149.505 40.040 149.555 ;
        RECT 41.530 149.525 42.475 149.555 ;
        RECT 43.405 150.205 46.230 150.435 ;
        RECT 43.405 149.525 46.935 150.205 ;
        RECT 47.115 149.525 49.835 150.435 ;
        RECT 49.845 149.525 53.515 150.335 ;
        RECT 53.535 149.525 56.265 150.435 ;
        RECT 57.655 150.205 58.575 150.435 ;
        RECT 56.285 149.525 58.575 150.205 ;
        RECT 58.585 150.205 59.505 150.435 ;
        RECT 58.585 149.525 60.875 150.205 ;
        RECT 61.355 149.610 61.785 150.395 ;
        RECT 64.095 150.205 65.015 150.435 ;
        RECT 62.725 149.525 65.015 150.205 ;
        RECT 65.025 149.525 66.395 150.335 ;
        RECT 66.490 149.525 75.595 150.205 ;
        RECT 75.605 149.525 77.435 150.335 ;
        RECT 80.960 150.205 81.870 150.425 ;
        RECT 83.405 150.205 84.755 150.435 ;
        RECT 86.175 150.205 87.095 150.435 ;
        RECT 77.445 149.525 84.755 150.205 ;
        RECT 84.805 149.525 87.095 150.205 ;
        RECT 87.115 149.610 87.545 150.395 ;
        RECT 91.080 150.205 91.990 150.425 ;
        RECT 93.525 150.205 94.875 150.435 ;
        RECT 87.565 149.525 94.875 150.205 ;
        RECT 94.925 149.525 98.135 150.435 ;
        RECT 98.345 150.345 99.295 150.435 ;
        RECT 98.345 149.525 100.275 150.345 ;
        RECT 100.445 149.525 103.555 150.435 ;
        RECT 104.585 149.525 107.795 150.435 ;
        RECT 107.805 149.525 112.620 150.205 ;
        RECT 112.875 149.610 113.305 150.395 ;
        RECT 113.325 149.525 115.155 150.335 ;
        RECT 119.140 150.205 120.050 150.425 ;
        RECT 121.585 150.205 122.935 150.435 ;
        RECT 115.625 149.525 122.935 150.205 ;
        RECT 123.080 150.205 124.000 150.435 ;
        RECT 129.320 150.205 130.240 150.435 ;
        RECT 123.080 149.525 126.545 150.205 ;
        RECT 126.775 149.525 130.240 150.205 ;
        RECT 130.345 149.525 133.555 150.435 ;
        RECT 133.575 149.525 136.305 150.435 ;
        RECT 136.325 149.525 138.155 150.205 ;
        RECT 138.635 149.610 139.065 150.395 ;
        RECT 139.085 149.525 144.595 150.335 ;
        RECT 144.605 149.525 147.355 150.335 ;
        RECT 147.865 150.205 149.215 150.435 ;
        RECT 150.750 150.205 151.660 150.425 ;
        RECT 147.865 149.525 155.175 150.205 ;
        RECT 155.645 149.525 157.015 150.335 ;
        RECT 46.735 149.505 46.935 149.525 ;
        RECT 39.405 149.475 39.575 149.505 ;
        RECT 39.400 149.365 39.575 149.475 ;
        RECT 39.405 149.315 39.575 149.365 ;
        RECT 39.865 149.335 40.040 149.505 ;
        RECT 42.635 149.370 42.795 149.480 ;
        RECT 39.865 149.315 40.035 149.335 ;
        RECT 45.385 149.315 45.555 149.505 ;
        RECT 46.765 149.335 46.935 149.505 ;
        RECT 48.140 149.365 48.260 149.475 ;
        RECT 49.525 149.335 49.695 149.525 ;
        RECT 49.985 149.505 50.155 149.525 ;
        RECT 49.985 149.335 50.160 149.505 ;
        RECT 49.990 149.315 50.160 149.335 ;
        RECT 51.370 149.315 51.540 149.505 ;
        RECT 51.820 149.365 51.940 149.475 ;
        RECT 53.665 149.335 53.835 149.525 ;
        RECT 56.425 149.335 56.595 149.525 ;
        RECT 59.185 149.315 59.355 149.505 ;
        RECT 60.565 149.335 60.735 149.525 ;
        RECT 61.020 149.365 61.140 149.475 ;
        RECT 61.955 149.370 62.115 149.480 ;
        RECT 62.865 149.335 63.035 149.525 ;
        RECT 65.165 149.335 65.335 149.525 ;
        RECT 66.545 149.315 66.715 149.505 ;
        RECT 73.905 149.315 74.075 149.505 ;
        RECT 74.820 149.365 74.940 149.475 ;
        RECT 75.285 149.335 75.455 149.525 ;
        RECT 75.745 149.335 75.915 149.525 ;
        RECT 77.585 149.335 77.755 149.525 ;
        RECT 75.305 149.315 75.455 149.335 ;
        RECT 78.505 149.315 78.675 149.505 ;
        RECT 78.965 149.315 79.135 149.505 ;
        RECT 80.800 149.365 80.920 149.475 ;
        RECT 81.265 149.315 81.435 149.505 ;
        RECT 84.025 149.315 84.195 149.505 ;
        RECT 84.945 149.335 85.115 149.525 ;
        RECT 87.705 149.315 87.875 149.525 ;
        RECT 88.165 149.315 88.335 149.505 ;
        RECT 95.065 149.335 95.235 149.525 ;
        RECT 100.125 149.505 100.275 149.525 ;
        RECT 98.285 149.315 98.455 149.505 ;
        RECT 98.745 149.315 98.915 149.505 ;
        RECT 100.125 149.335 100.295 149.505 ;
        RECT 103.345 149.335 103.515 149.525 ;
        RECT 103.815 149.370 103.975 149.480 ;
        RECT 107.485 149.315 107.655 149.525 ;
        RECT 107.945 149.315 108.115 149.525 ;
        RECT 113.465 149.335 113.635 149.525 ;
        RECT 115.300 149.470 115.420 149.475 ;
        RECT 115.300 149.365 115.475 149.470 ;
        RECT 115.315 149.360 115.475 149.365 ;
        RECT 115.765 149.335 115.935 149.525 ;
        RECT 116.225 149.315 116.395 149.505 ;
        RECT 125.420 149.365 125.540 149.475 ;
        RECT 126.345 149.335 126.515 149.525 ;
        RECT 126.805 149.335 126.975 149.525 ;
        RECT 129.105 149.315 129.275 149.505 ;
        RECT 132.325 149.315 132.495 149.505 ;
        RECT 132.785 149.335 132.955 149.505 ;
        RECT 133.245 149.335 133.415 149.525 ;
        RECT 132.805 149.315 132.955 149.335 ;
        RECT 136.005 149.315 136.175 149.525 ;
        RECT 136.465 149.315 136.635 149.525 ;
        RECT 138.300 149.365 138.420 149.475 ;
        RECT 139.225 149.335 139.395 149.525 ;
        RECT 141.985 149.315 142.155 149.505 ;
        RECT 144.745 149.335 144.915 149.525 ;
        RECT 147.500 149.365 147.620 149.475 ;
        RECT 147.965 149.315 148.135 149.505 ;
        RECT 149.345 149.315 149.515 149.505 ;
        RECT 151.180 149.365 151.300 149.475 ;
        RECT 152.105 149.315 152.275 149.505 ;
        RECT 154.865 149.335 155.035 149.525 ;
        RECT 155.320 149.365 155.440 149.475 ;
        RECT 156.705 149.315 156.875 149.525 ;
        RECT 22.705 148.505 24.075 149.315 ;
        RECT 24.085 148.505 29.595 149.315 ;
        RECT 29.605 148.505 32.355 149.315 ;
        RECT 32.405 148.635 39.715 149.315 ;
        RECT 32.405 148.405 33.755 148.635 ;
        RECT 35.290 148.415 36.200 148.635 ;
        RECT 39.725 148.505 45.235 149.315 ;
        RECT 45.245 148.505 47.995 149.315 ;
        RECT 48.475 148.445 48.905 149.230 ;
        RECT 48.925 148.405 50.275 149.315 ;
        RECT 50.305 148.405 51.655 149.315 ;
        RECT 52.185 148.635 59.495 149.315 ;
        RECT 59.545 148.635 66.855 149.315 ;
        RECT 66.905 148.635 74.215 149.315 ;
        RECT 52.185 148.405 53.535 148.635 ;
        RECT 55.070 148.415 55.980 148.635 ;
        RECT 59.545 148.405 60.895 148.635 ;
        RECT 62.430 148.415 63.340 148.635 ;
        RECT 66.905 148.405 68.255 148.635 ;
        RECT 69.790 148.415 70.700 148.635 ;
        RECT 74.235 148.445 74.665 149.230 ;
        RECT 75.305 148.495 77.235 149.315 ;
        RECT 77.445 148.535 78.815 149.315 ;
        RECT 78.825 148.505 80.655 149.315 ;
        RECT 76.285 148.405 77.235 148.495 ;
        RECT 81.135 148.405 83.865 149.315 ;
        RECT 83.885 148.505 85.255 149.315 ;
        RECT 85.275 148.405 88.005 149.315 ;
        RECT 88.035 148.405 89.385 149.315 ;
        RECT 89.490 148.635 98.595 149.315 ;
        RECT 98.605 148.505 99.975 149.315 ;
        RECT 99.995 148.445 100.425 149.230 ;
        RECT 100.485 148.635 107.795 149.315 ;
        RECT 107.805 148.635 115.115 149.315 ;
        RECT 116.085 148.635 125.190 149.315 ;
        RECT 100.485 148.405 101.835 148.635 ;
        RECT 103.370 148.415 104.280 148.635 ;
        RECT 111.320 148.415 112.230 148.635 ;
        RECT 113.765 148.405 115.115 148.635 ;
        RECT 125.755 148.445 126.185 149.230 ;
        RECT 126.205 148.405 129.415 149.315 ;
        RECT 129.425 148.405 132.635 149.315 ;
        RECT 132.805 148.495 134.735 149.315 ;
        RECT 133.785 148.405 134.735 148.495 ;
        RECT 134.955 148.405 136.305 149.315 ;
        RECT 136.325 148.505 141.835 149.315 ;
        RECT 141.845 148.505 147.355 149.315 ;
        RECT 147.825 148.535 149.195 149.315 ;
        RECT 149.205 148.505 151.035 149.315 ;
        RECT 151.515 148.445 151.945 149.230 ;
        RECT 151.965 148.505 155.635 149.315 ;
        RECT 155.645 148.505 157.015 149.315 ;
      LAYER nwell ;
        RECT 22.510 145.285 157.210 148.115 ;
      LAYER pwell ;
        RECT 29.345 144.905 30.295 144.995 ;
        RECT 22.705 144.085 24.075 144.895 ;
        RECT 24.085 144.085 25.455 144.895 ;
        RECT 25.465 144.085 26.835 144.865 ;
        RECT 26.845 144.085 28.675 144.895 ;
        RECT 29.345 144.085 31.275 144.905 ;
        RECT 31.755 144.765 32.685 144.995 ;
        RECT 31.755 144.085 33.590 144.765 ;
        RECT 33.745 144.085 35.575 144.895 ;
        RECT 35.595 144.170 36.025 144.955 ;
        RECT 36.045 144.085 41.555 144.895 ;
        RECT 42.485 144.085 46.615 144.995 ;
        RECT 47.085 144.085 50.740 144.995 ;
        RECT 50.775 144.085 52.125 144.995 ;
        RECT 52.155 144.085 53.505 144.995 ;
        RECT 53.525 144.085 56.275 144.895 ;
        RECT 56.295 144.085 59.025 144.995 ;
        RECT 59.045 144.085 60.875 144.895 ;
        RECT 61.355 144.170 61.785 144.955 ;
        RECT 62.735 144.085 65.465 144.995 ;
        RECT 74.520 144.765 75.430 144.985 ;
        RECT 76.965 144.765 78.315 144.995 ;
        RECT 65.945 144.085 70.760 144.765 ;
        RECT 71.005 144.085 78.315 144.765 ;
        RECT 78.365 144.765 79.295 144.995 ;
        RECT 78.365 144.085 82.265 144.765 ;
        RECT 82.505 144.085 85.255 144.895 ;
        RECT 85.735 144.085 87.085 144.995 ;
        RECT 87.115 144.170 87.545 144.955 ;
        RECT 88.025 144.765 88.945 144.995 ;
        RECT 88.025 144.085 90.315 144.765 ;
        RECT 90.800 144.085 94.455 144.995 ;
        RECT 95.515 144.765 96.445 144.995 ;
        RECT 94.610 144.085 96.445 144.765 ;
        RECT 96.765 144.795 97.695 144.995 ;
        RECT 99.025 144.795 99.975 144.995 ;
        RECT 96.765 144.315 99.975 144.795 ;
        RECT 101.035 144.765 101.965 144.995 ;
        RECT 96.910 144.115 99.975 144.315 ;
        RECT 22.845 143.875 23.015 144.085 ;
        RECT 24.225 143.875 24.395 144.085 ;
        RECT 26.525 143.895 26.695 144.085 ;
        RECT 26.985 143.895 27.155 144.085 ;
        RECT 31.125 144.065 31.275 144.085 ;
        RECT 33.425 144.065 33.590 144.085 ;
        RECT 28.820 143.925 28.940 144.035 ;
        RECT 31.125 143.895 31.295 144.065 ;
        RECT 33.425 143.895 33.595 144.065 ;
        RECT 33.885 143.895 34.055 144.085 ;
        RECT 34.340 143.875 34.510 144.065 ;
        RECT 34.805 143.875 34.975 144.065 ;
        RECT 36.185 143.895 36.355 144.085 ;
        RECT 39.865 143.875 40.035 144.065 ;
        RECT 40.325 143.875 40.495 144.065 ;
        RECT 41.705 143.875 41.875 144.065 ;
        RECT 43.085 143.875 43.255 144.065 ;
        RECT 44.465 143.875 44.635 144.065 ;
        RECT 46.305 143.895 46.475 144.085 ;
        RECT 46.760 143.925 46.880 144.035 ;
        RECT 47.230 143.895 47.400 144.085 ;
        RECT 47.695 143.920 47.855 144.030 ;
        RECT 22.705 143.065 24.075 143.875 ;
        RECT 24.085 143.195 31.395 143.875 ;
        RECT 27.600 142.975 28.510 143.195 ;
        RECT 30.045 142.965 31.395 143.195 ;
        RECT 31.735 142.965 34.655 143.875 ;
        RECT 34.665 143.065 36.495 143.875 ;
        RECT 36.600 143.195 40.065 143.875 ;
        RECT 36.600 142.965 37.520 143.195 ;
        RECT 40.185 143.095 41.555 143.875 ;
        RECT 41.575 142.965 42.925 143.875 ;
        RECT 42.955 142.965 44.305 143.875 ;
        RECT 44.325 142.965 47.535 143.875 ;
        RECT 48.925 143.845 49.870 143.875 ;
        RECT 51.360 143.845 51.530 144.065 ;
        RECT 51.825 144.035 51.995 144.085 ;
        RECT 51.820 143.925 51.995 144.035 ;
        RECT 51.825 143.895 51.995 143.925 ;
        RECT 52.285 143.895 52.455 144.085 ;
        RECT 53.665 143.895 53.835 144.085 ;
        RECT 54.125 143.875 54.295 144.065 ;
        RECT 54.585 143.875 54.755 144.065 ;
        RECT 56.425 143.895 56.595 144.085 ;
        RECT 59.185 143.895 59.355 144.085 ;
        RECT 60.105 143.875 60.275 144.065 ;
        RECT 61.020 143.925 61.140 144.035 ;
        RECT 61.955 143.930 62.115 144.040 ;
        RECT 62.865 143.895 63.035 144.085 ;
        RECT 63.785 143.875 63.955 144.065 ;
        RECT 64.245 143.875 64.415 144.065 ;
        RECT 65.620 143.925 65.740 144.035 ;
        RECT 66.085 143.895 66.255 144.085 ;
        RECT 67.005 143.875 67.175 144.065 ;
        RECT 67.460 143.925 67.580 144.035 ;
        RECT 68.200 143.875 68.370 144.065 ;
        RECT 71.145 143.895 71.315 144.085 ;
        RECT 72.065 143.875 72.235 144.065 ;
        RECT 73.900 143.925 74.020 144.035 ;
        RECT 75.745 143.875 75.915 144.065 ;
        RECT 76.200 143.925 76.320 144.035 ;
        RECT 76.665 143.895 76.835 144.065 ;
        RECT 78.780 143.895 78.950 144.085 ;
        RECT 76.685 143.875 76.835 143.895 ;
        RECT 78.965 143.875 79.135 144.065 ;
        RECT 80.805 143.875 80.975 144.065 ;
        RECT 82.645 143.895 82.815 144.085 ;
        RECT 85.400 143.925 85.520 144.035 ;
        RECT 86.785 143.895 86.955 144.085 ;
        RECT 87.700 143.925 87.820 144.035 ;
        RECT 88.175 143.920 88.335 144.030 ;
        RECT 89.085 143.875 89.255 144.065 ;
        RECT 90.005 143.895 90.175 144.085 ;
        RECT 90.460 143.925 90.580 144.035 ;
        RECT 92.765 143.875 92.935 144.065 ;
        RECT 94.140 143.895 94.310 144.085 ;
        RECT 94.610 144.065 94.775 144.085 ;
        RECT 94.605 143.895 94.775 144.065 ;
        RECT 95.985 143.895 96.155 144.065 ;
        RECT 96.910 143.895 97.080 144.115 ;
        RECT 99.040 144.085 99.975 144.115 ;
        RECT 100.130 144.085 101.965 144.765 ;
        RECT 102.285 144.085 103.655 144.865 ;
        RECT 104.135 144.085 106.875 144.765 ;
        RECT 106.885 144.085 110.095 144.995 ;
        RECT 110.105 144.085 112.845 144.765 ;
        RECT 112.875 144.170 113.305 144.955 ;
        RECT 113.325 144.085 114.695 144.895 ;
        RECT 118.220 144.765 119.130 144.985 ;
        RECT 120.665 144.765 122.015 144.995 ;
        RECT 114.705 144.085 122.015 144.765 ;
        RECT 122.065 144.085 123.435 144.895 ;
        RECT 123.445 144.085 126.655 144.995 ;
        RECT 126.680 144.085 128.495 144.995 ;
        RECT 128.505 144.085 129.875 144.895 ;
        RECT 129.895 144.085 132.625 144.995 ;
        RECT 132.645 144.795 133.595 144.995 ;
        RECT 134.925 144.795 135.855 144.995 ;
        RECT 137.005 144.905 137.955 144.995 ;
        RECT 132.645 144.315 135.855 144.795 ;
        RECT 132.645 144.115 135.710 144.315 ;
        RECT 132.645 144.085 133.580 144.115 ;
        RECT 100.130 144.065 100.295 144.085 ;
        RECT 96.135 143.875 96.155 143.895 ;
        RECT 98.740 143.875 98.910 144.065 ;
        RECT 100.125 143.895 100.295 144.065 ;
        RECT 100.595 143.920 100.755 144.030 ;
        RECT 102.425 143.895 102.595 144.085 ;
        RECT 103.800 143.925 103.920 144.035 ;
        RECT 104.725 143.875 104.895 144.065 ;
        RECT 105.185 143.875 105.355 144.065 ;
        RECT 106.565 143.875 106.735 144.085 ;
        RECT 108.400 143.925 108.520 144.035 ;
        RECT 108.870 143.875 109.040 144.065 ;
        RECT 109.785 143.895 109.955 144.085 ;
        RECT 110.245 143.875 110.415 144.085 ;
        RECT 112.080 143.925 112.200 144.035 ;
        RECT 113.465 143.895 113.635 144.085 ;
        RECT 114.845 143.895 115.015 144.085 ;
        RECT 115.765 143.875 115.935 144.065 ;
        RECT 116.235 143.920 116.395 144.030 ;
        RECT 119.905 143.875 120.075 144.065 ;
        RECT 120.365 143.875 120.535 144.065 ;
        RECT 122.205 143.895 122.375 144.085 ;
        RECT 123.585 143.895 123.755 144.085 ;
        RECT 126.805 143.895 126.975 144.085 ;
        RECT 128.645 143.895 128.815 144.085 ;
        RECT 129.560 143.875 129.730 144.065 ;
        RECT 130.030 143.875 130.200 144.065 ;
        RECT 132.325 143.875 132.495 144.085 ;
        RECT 135.540 143.895 135.710 144.115 ;
        RECT 136.025 144.085 137.955 144.905 ;
        RECT 138.635 144.170 139.065 144.955 ;
        RECT 139.085 144.085 140.455 144.865 ;
        RECT 140.475 144.085 141.825 144.995 ;
        RECT 141.865 144.085 143.215 144.995 ;
        RECT 144.275 144.765 145.205 144.995 ;
        RECT 146.895 144.765 147.815 144.995 ;
        RECT 143.370 144.085 145.205 144.765 ;
        RECT 145.525 144.085 147.815 144.765 ;
        RECT 148.325 144.765 149.675 144.995 ;
        RECT 151.210 144.765 152.120 144.985 ;
        RECT 148.325 144.085 155.635 144.765 ;
        RECT 155.645 144.085 157.015 144.895 ;
        RECT 136.025 144.065 136.175 144.085 ;
        RECT 136.005 143.895 136.175 144.065 ;
        RECT 138.300 143.925 138.420 144.035 ;
        RECT 139.225 143.895 139.395 144.085 ;
        RECT 141.065 143.875 141.235 144.065 ;
        RECT 141.525 143.895 141.695 144.085 ;
        RECT 141.980 143.895 142.150 144.085 ;
        RECT 143.370 144.065 143.535 144.085 ;
        RECT 145.665 144.065 145.835 144.085 ;
        RECT 143.365 143.895 143.535 144.065 ;
        RECT 144.285 143.875 144.455 144.065 ;
        RECT 144.755 143.920 144.915 144.030 ;
        RECT 145.665 143.895 145.840 144.065 ;
        RECT 147.960 143.925 148.080 144.035 ;
        RECT 48.475 143.005 48.905 143.790 ;
        RECT 48.925 143.165 51.675 143.845 ;
        RECT 52.145 143.195 54.435 143.875 ;
        RECT 54.445 143.195 56.735 143.875 ;
        RECT 48.925 142.965 49.870 143.165 ;
        RECT 52.145 142.965 53.065 143.195 ;
        RECT 55.815 142.965 56.735 143.195 ;
        RECT 56.840 143.195 60.305 143.875 ;
        RECT 60.520 143.195 63.985 143.875 ;
        RECT 56.840 142.965 57.760 143.195 ;
        RECT 60.520 142.965 61.440 143.195 ;
        RECT 64.105 143.065 65.935 143.875 ;
        RECT 65.945 143.095 67.315 143.875 ;
        RECT 67.785 143.195 71.685 143.875 ;
        RECT 67.785 142.965 68.715 143.195 ;
        RECT 71.925 143.065 73.755 143.875 ;
        RECT 74.235 143.005 74.665 143.790 ;
        RECT 74.685 143.095 76.055 143.875 ;
        RECT 76.685 143.055 78.615 143.875 ;
        RECT 78.825 143.065 80.655 143.875 ;
        RECT 80.665 143.195 87.975 143.875 ;
        RECT 89.055 143.195 92.520 143.875 ;
        RECT 77.665 142.965 78.615 143.055 ;
        RECT 84.180 142.975 85.090 143.195 ;
        RECT 86.625 142.965 87.975 143.195 ;
        RECT 91.600 142.965 92.520 143.195 ;
        RECT 92.625 142.965 95.835 143.875 ;
        RECT 96.135 143.195 98.585 143.875 ;
        RECT 96.625 142.965 98.585 143.195 ;
        RECT 98.625 142.965 99.975 143.875 ;
        RECT 99.995 143.005 100.425 143.790 ;
        RECT 101.460 143.195 104.925 143.875 ;
        RECT 101.460 142.965 102.380 143.195 ;
        RECT 105.045 143.095 106.415 143.875 ;
        RECT 106.425 143.065 108.255 143.875 ;
        RECT 108.725 142.965 110.075 143.875 ;
        RECT 110.105 143.065 111.935 143.875 ;
        RECT 112.500 143.195 115.965 143.875 ;
        RECT 112.500 142.965 113.420 143.195 ;
        RECT 117.005 142.965 120.215 143.875 ;
        RECT 120.225 143.065 125.735 143.875 ;
        RECT 125.755 143.005 126.185 143.790 ;
        RECT 126.220 142.965 129.875 143.875 ;
        RECT 130.030 143.645 131.720 143.875 ;
        RECT 129.885 142.965 131.720 143.645 ;
        RECT 132.185 143.065 134.015 143.875 ;
        RECT 134.065 143.195 141.375 143.875 ;
        RECT 141.385 143.195 144.595 143.875 ;
        RECT 145.670 143.845 145.840 143.895 ;
        RECT 148.890 143.875 149.060 144.065 ;
        RECT 151.190 143.875 151.360 144.065 ;
        RECT 152.105 143.875 152.275 144.065 ;
        RECT 153.485 143.875 153.655 144.065 ;
        RECT 155.325 144.035 155.495 144.085 ;
        RECT 155.320 143.925 155.495 144.035 ;
        RECT 155.325 143.895 155.495 143.925 ;
        RECT 156.705 143.875 156.875 144.085 ;
        RECT 147.800 143.845 148.735 143.875 ;
        RECT 145.670 143.645 148.735 143.845 ;
        RECT 134.065 142.965 135.415 143.195 ;
        RECT 136.950 142.975 137.860 143.195 ;
        RECT 141.385 142.965 142.520 143.195 ;
        RECT 145.525 143.165 148.735 143.645 ;
        RECT 145.525 142.965 146.455 143.165 ;
        RECT 147.785 142.965 148.735 143.165 ;
        RECT 148.745 142.965 150.095 143.875 ;
        RECT 150.125 142.965 151.475 143.875 ;
        RECT 151.515 143.005 151.945 143.790 ;
        RECT 151.965 143.095 153.335 143.875 ;
        RECT 153.345 143.065 155.175 143.875 ;
        RECT 155.645 143.065 157.015 143.875 ;
      LAYER nwell ;
        RECT 22.510 139.845 157.210 142.675 ;
      LAYER pwell ;
        RECT 22.705 138.645 24.075 139.455 ;
        RECT 24.085 138.645 25.915 139.455 ;
        RECT 26.385 139.355 27.335 139.555 ;
        RECT 28.665 139.355 29.595 139.555 ;
        RECT 26.385 138.875 29.595 139.355 ;
        RECT 31.435 139.325 32.355 139.555 ;
        RECT 26.385 138.675 29.450 138.875 ;
        RECT 26.385 138.645 27.320 138.675 ;
        RECT 22.845 138.435 23.015 138.645 ;
        RECT 24.225 138.435 24.395 138.645 ;
        RECT 26.060 138.485 26.180 138.595 ;
        RECT 29.280 138.455 29.450 138.675 ;
        RECT 30.065 138.645 32.355 139.325 ;
        RECT 32.365 139.355 33.295 139.555 ;
        RECT 34.625 139.355 35.575 139.555 ;
        RECT 32.365 138.875 35.575 139.355 ;
        RECT 32.510 138.675 35.575 138.875 ;
        RECT 35.595 138.730 36.025 139.515 ;
        RECT 36.085 139.325 37.435 139.555 ;
        RECT 38.970 139.325 39.880 139.545 ;
        RECT 29.740 138.590 29.860 138.595 ;
        RECT 29.740 138.485 29.915 138.590 ;
        RECT 29.755 138.480 29.915 138.485 ;
        RECT 30.205 138.455 30.375 138.645 ;
        RECT 30.665 138.435 30.835 138.625 ;
        RECT 32.510 138.455 32.680 138.675 ;
        RECT 34.640 138.645 35.575 138.675 ;
        RECT 36.085 138.645 43.395 139.325 ;
        RECT 44.335 138.645 45.685 139.555 ;
        RECT 45.705 138.645 49.835 139.555 ;
        RECT 49.845 138.645 51.215 139.455 ;
        RECT 51.235 138.645 53.965 139.555 ;
        RECT 54.025 139.325 55.375 139.555 ;
        RECT 56.910 139.325 57.820 139.545 ;
        RECT 54.025 138.645 61.335 139.325 ;
        RECT 61.355 138.730 61.785 139.515 ;
        RECT 61.805 138.645 63.635 139.455 ;
        RECT 67.160 139.325 68.070 139.545 ;
        RECT 69.605 139.325 70.955 139.555 ;
        RECT 63.645 138.645 70.955 139.325 ;
        RECT 71.015 138.645 72.365 139.555 ;
        RECT 73.305 138.645 76.415 139.555 ;
        RECT 76.525 138.645 82.035 139.455 ;
        RECT 82.975 138.645 85.705 139.555 ;
        RECT 85.725 138.645 87.095 139.455 ;
        RECT 87.115 138.730 87.545 139.515 ;
        RECT 92.000 139.325 92.910 139.545 ;
        RECT 94.445 139.325 95.795 139.555 ;
        RECT 88.485 138.645 95.795 139.325 ;
        RECT 95.940 139.325 96.860 139.555 ;
        RECT 95.940 138.645 99.405 139.325 ;
        RECT 99.525 138.645 101.355 139.455 ;
        RECT 101.405 139.325 102.755 139.555 ;
        RECT 104.290 139.325 105.200 139.545 ;
        RECT 101.405 138.645 108.715 139.325 ;
        RECT 109.645 138.645 112.855 139.555 ;
        RECT 112.875 138.730 113.305 139.515 ;
        RECT 117.760 139.325 118.670 139.545 ;
        RECT 120.205 139.325 121.555 139.555 ;
        RECT 114.245 138.645 121.555 139.325 ;
        RECT 121.700 139.325 122.620 139.555 ;
        RECT 121.700 138.645 125.165 139.325 ;
        RECT 125.285 138.645 127.115 139.455 ;
        RECT 127.125 138.645 128.940 139.555 ;
        RECT 128.965 138.645 132.635 139.455 ;
        RECT 134.345 139.325 136.305 139.555 ;
        RECT 133.855 138.645 136.305 139.325 ;
        RECT 136.325 138.645 138.155 139.455 ;
        RECT 138.635 138.730 139.065 139.515 ;
        RECT 139.095 138.645 140.445 139.555 ;
        RECT 143.580 139.325 144.500 139.555 ;
        RECT 146.115 139.325 147.045 139.555 ;
        RECT 151.800 139.325 152.710 139.545 ;
        RECT 154.245 139.325 155.595 139.555 ;
        RECT 141.035 138.645 144.500 139.325 ;
        RECT 145.210 138.645 147.045 139.325 ;
        RECT 148.285 138.645 155.595 139.325 ;
        RECT 155.645 138.645 157.015 139.455 ;
        RECT 33.425 138.435 33.595 138.625 ;
        RECT 40.785 138.435 40.955 138.625 ;
        RECT 22.705 137.625 24.075 138.435 ;
        RECT 24.085 137.625 29.595 138.435 ;
        RECT 30.525 137.525 33.275 138.435 ;
        RECT 33.285 137.755 40.595 138.435 ;
        RECT 36.800 137.535 37.710 137.755 ;
        RECT 39.245 137.525 40.595 137.755 ;
        RECT 40.645 137.625 42.015 138.435 ;
        RECT 42.170 138.405 42.340 138.625 ;
        RECT 43.085 138.455 43.255 138.645 ;
        RECT 43.555 138.490 43.715 138.600 ;
        RECT 44.465 138.455 44.635 138.645 ;
        RECT 43.830 138.405 44.775 138.435 ;
        RECT 44.930 138.405 45.100 138.625 ;
        RECT 45.845 138.455 46.015 138.645 ;
        RECT 47.695 138.480 47.855 138.590 ;
        RECT 49.065 138.435 49.235 138.625 ;
        RECT 49.985 138.455 50.155 138.645 ;
        RECT 50.445 138.435 50.615 138.625 ;
        RECT 51.365 138.455 51.535 138.645 ;
        RECT 57.800 138.485 57.920 138.595 ;
        RECT 58.265 138.435 58.435 138.625 ;
        RECT 61.025 138.435 61.195 138.645 ;
        RECT 61.945 138.455 62.115 138.645 ;
        RECT 63.785 138.455 63.955 138.645 ;
        RECT 66.820 138.435 66.990 138.625 ;
        RECT 70.690 138.435 70.860 138.625 ;
        RECT 71.145 138.455 71.315 138.645 ;
        RECT 72.065 138.435 72.235 138.625 ;
        RECT 72.535 138.490 72.695 138.600 ;
        RECT 73.900 138.485 74.020 138.595 ;
        RECT 74.820 138.485 74.940 138.595 ;
        RECT 75.560 138.435 75.730 138.625 ;
        RECT 76.205 138.455 76.375 138.645 ;
        RECT 76.665 138.455 76.835 138.645 ;
        RECT 79.425 138.435 79.595 138.625 ;
        RECT 82.195 138.490 82.355 138.600 ;
        RECT 83.105 138.455 83.275 138.645 ;
        RECT 85.865 138.435 86.035 138.645 ;
        RECT 87.715 138.490 87.875 138.600 ;
        RECT 88.625 138.455 88.795 138.645 ;
        RECT 89.545 138.435 89.715 138.625 ;
        RECT 91.845 138.455 92.015 138.625 ;
        RECT 91.845 138.435 92.010 138.455 ;
        RECT 92.305 138.435 92.475 138.625 ;
        RECT 93.685 138.455 93.855 138.625 ;
        RECT 93.695 138.435 93.855 138.455 ;
        RECT 97.830 138.435 98.000 138.625 ;
        RECT 99.205 138.455 99.375 138.645 ;
        RECT 99.665 138.595 99.835 138.645 ;
        RECT 99.660 138.485 99.835 138.595 ;
        RECT 99.665 138.455 99.835 138.485 ;
        RECT 100.585 138.455 100.755 138.625 ;
        RECT 100.590 138.435 100.755 138.455 ;
        RECT 102.885 138.435 103.055 138.625 ;
        RECT 106.100 138.435 106.270 138.625 ;
        RECT 106.565 138.435 106.735 138.625 ;
        RECT 108.405 138.455 108.575 138.645 ;
        RECT 108.875 138.490 109.035 138.600 ;
        RECT 109.785 138.455 109.955 138.645 ;
        RECT 113.475 138.490 113.635 138.600 ;
        RECT 114.385 138.455 114.555 138.645 ;
        RECT 117.145 138.435 117.315 138.625 ;
        RECT 117.600 138.485 117.720 138.595 ;
        RECT 121.285 138.435 121.455 138.625 ;
        RECT 124.965 138.435 125.135 138.645 ;
        RECT 125.425 138.595 125.595 138.645 ;
        RECT 125.420 138.485 125.595 138.595 ;
        RECT 125.425 138.455 125.595 138.485 ;
        RECT 128.645 138.455 128.815 138.645 ;
        RECT 129.105 138.455 129.275 138.645 ;
        RECT 133.855 138.625 133.875 138.645 ;
        RECT 129.560 138.435 129.730 138.625 ;
        RECT 132.785 138.435 132.955 138.625 ;
        RECT 133.240 138.485 133.360 138.595 ;
        RECT 133.705 138.435 133.875 138.625 ;
        RECT 136.465 138.455 136.635 138.645 ;
        RECT 138.300 138.485 138.420 138.595 ;
        RECT 140.145 138.455 140.315 138.645 ;
        RECT 140.600 138.485 140.720 138.595 ;
        RECT 141.065 138.455 141.235 138.645 ;
        RECT 145.210 138.625 145.375 138.645 ;
        RECT 141.985 138.435 142.155 138.625 ;
        RECT 142.455 138.480 142.615 138.590 ;
        RECT 144.285 138.435 144.455 138.625 ;
        RECT 144.750 138.595 144.920 138.625 ;
        RECT 144.740 138.485 144.920 138.595 ;
        RECT 46.590 138.405 47.535 138.435 ;
        RECT 42.025 137.725 44.775 138.405 ;
        RECT 44.785 137.725 47.535 138.405 ;
        RECT 43.830 137.525 44.775 137.725 ;
        RECT 46.590 137.525 47.535 137.725 ;
        RECT 48.475 137.565 48.905 138.350 ;
        RECT 48.925 137.625 50.295 138.435 ;
        RECT 50.305 137.755 57.615 138.435 ;
        RECT 53.820 137.535 54.730 137.755 ;
        RECT 56.265 137.525 57.615 137.755 ;
        RECT 58.135 137.525 60.865 138.435 ;
        RECT 60.885 137.625 66.395 138.435 ;
        RECT 66.405 137.755 70.305 138.435 ;
        RECT 66.405 137.525 67.335 137.755 ;
        RECT 70.545 137.525 71.895 138.435 ;
        RECT 71.925 137.625 73.755 138.435 ;
        RECT 74.235 137.565 74.665 138.350 ;
        RECT 75.145 137.755 79.045 138.435 ;
        RECT 75.145 137.525 76.075 137.755 ;
        RECT 79.285 137.625 82.955 138.435 ;
        RECT 83.885 137.755 86.175 138.435 ;
        RECT 86.280 137.755 89.745 138.435 ;
        RECT 90.175 137.755 92.010 138.435 ;
        RECT 83.885 137.525 84.805 137.755 ;
        RECT 86.280 137.525 87.200 137.755 ;
        RECT 90.175 137.525 91.105 137.755 ;
        RECT 92.175 137.525 93.525 138.435 ;
        RECT 93.695 137.525 97.350 138.435 ;
        RECT 97.685 137.525 99.515 138.435 ;
        RECT 99.995 137.565 100.425 138.350 ;
        RECT 100.590 137.755 102.425 138.435 ;
        RECT 102.745 137.755 105.035 138.435 ;
        RECT 101.495 137.525 102.425 137.755 ;
        RECT 104.115 137.525 105.035 137.755 ;
        RECT 105.065 137.525 106.415 138.435 ;
        RECT 106.425 137.755 113.735 138.435 ;
        RECT 109.940 137.535 110.850 137.755 ;
        RECT 112.385 137.525 113.735 137.755 ;
        RECT 113.880 137.755 117.345 138.435 ;
        RECT 118.020 137.755 121.485 138.435 ;
        RECT 121.700 137.755 125.165 138.435 ;
        RECT 113.880 137.525 114.800 137.755 ;
        RECT 118.020 137.525 118.940 137.755 ;
        RECT 121.700 137.525 122.620 137.755 ;
        RECT 125.755 137.565 126.185 138.350 ;
        RECT 126.290 137.755 129.875 138.435 ;
        RECT 128.955 137.525 129.875 137.755 ;
        RECT 129.885 137.525 133.095 138.435 ;
        RECT 133.565 137.755 140.875 138.435 ;
        RECT 137.080 137.535 137.990 137.755 ;
        RECT 139.525 137.525 140.875 137.755 ;
        RECT 140.935 137.525 142.285 138.435 ;
        RECT 143.235 137.525 144.585 138.435 ;
        RECT 144.750 138.405 144.920 138.485 ;
        RECT 145.205 138.455 145.375 138.625 ;
        RECT 147.515 138.490 147.675 138.600 ;
        RECT 147.965 138.435 148.135 138.625 ;
        RECT 148.425 138.455 148.595 138.645 ;
        RECT 149.345 138.435 149.515 138.625 ;
        RECT 150.735 138.480 150.895 138.590 ;
        RECT 152.105 138.435 152.275 138.625 ;
        RECT 156.705 138.435 156.875 138.645 ;
        RECT 146.880 138.405 147.815 138.435 ;
        RECT 144.750 138.205 147.815 138.405 ;
        RECT 144.605 137.725 147.815 138.205 ;
        RECT 144.605 137.525 145.535 137.725 ;
        RECT 146.865 137.525 147.815 137.725 ;
        RECT 147.825 137.625 149.195 138.435 ;
        RECT 149.205 137.655 150.575 138.435 ;
        RECT 151.515 137.565 151.945 138.350 ;
        RECT 151.965 137.625 155.635 138.435 ;
        RECT 155.645 137.625 157.015 138.435 ;
      LAYER nwell ;
        RECT 22.510 134.405 157.210 137.235 ;
      LAYER pwell ;
        RECT 22.705 133.205 24.075 134.015 ;
        RECT 24.085 133.205 26.835 134.015 ;
        RECT 27.155 133.885 28.085 134.115 ;
        RECT 29.145 133.885 30.065 134.115 ;
        RECT 27.155 133.205 28.990 133.885 ;
        RECT 29.145 133.205 31.435 133.885 ;
        RECT 31.465 133.205 32.815 134.115 ;
        RECT 32.825 133.205 35.575 134.015 ;
        RECT 35.595 133.290 36.025 134.075 ;
        RECT 36.140 133.885 37.060 134.115 ;
        RECT 41.115 134.025 42.705 134.115 ;
        RECT 36.140 133.205 39.605 133.885 ;
        RECT 39.725 133.205 41.095 134.015 ;
        RECT 41.115 133.205 43.685 134.025 ;
        RECT 43.960 133.885 44.880 134.115 ;
        RECT 43.960 133.205 47.425 133.885 ;
        RECT 47.545 133.205 51.215 134.015 ;
        RECT 51.225 133.205 52.595 134.015 ;
        RECT 52.700 133.885 53.620 134.115 ;
        RECT 52.700 133.205 56.165 133.885 ;
        RECT 56.285 133.205 59.955 134.015 ;
        RECT 59.965 133.205 61.335 134.015 ;
        RECT 61.355 133.290 61.785 134.075 ;
        RECT 61.805 133.205 67.315 134.015 ;
        RECT 67.325 133.205 70.075 134.015 ;
        RECT 70.545 133.205 71.915 133.985 ;
        RECT 75.440 133.885 76.350 134.105 ;
        RECT 77.885 133.885 79.235 134.115 ;
        RECT 82.800 133.885 83.710 134.105 ;
        RECT 85.245 133.885 86.595 134.115 ;
        RECT 71.925 133.205 79.235 133.885 ;
        RECT 79.285 133.205 86.595 133.885 ;
        RECT 87.115 133.290 87.545 134.075 ;
        RECT 87.565 133.885 88.485 134.115 ;
        RECT 87.565 133.205 89.855 133.885 ;
        RECT 90.335 133.205 91.685 134.115 ;
        RECT 91.705 133.205 95.375 134.015 ;
        RECT 95.855 133.205 97.205 134.115 ;
        RECT 97.225 133.205 98.575 134.115 ;
        RECT 98.605 133.205 104.115 134.015 ;
        RECT 104.125 133.205 106.875 134.015 ;
        RECT 107.345 133.205 110.555 134.115 ;
        RECT 110.565 133.205 112.395 134.015 ;
        RECT 112.875 133.290 113.305 134.075 ;
        RECT 113.325 133.205 116.075 134.015 ;
        RECT 119.600 133.885 120.510 134.105 ;
        RECT 122.045 133.885 123.395 134.115 ;
        RECT 116.085 133.205 123.395 133.885 ;
        RECT 123.455 133.205 124.805 134.115 ;
        RECT 125.305 133.205 126.655 134.115 ;
        RECT 126.815 133.205 130.470 134.115 ;
        RECT 130.805 133.885 131.735 134.115 ;
        RECT 130.805 133.205 133.555 133.885 ;
        RECT 133.565 133.205 134.935 134.015 ;
        RECT 135.040 133.885 135.960 134.115 ;
        RECT 135.040 133.205 138.505 133.885 ;
        RECT 138.635 133.290 139.065 134.075 ;
        RECT 140.225 134.025 141.175 134.115 ;
        RECT 139.245 133.205 141.175 134.025 ;
        RECT 141.580 133.205 145.055 134.115 ;
        RECT 148.580 133.885 149.490 134.105 ;
        RECT 151.025 133.885 152.375 134.115 ;
        RECT 145.065 133.205 152.375 133.885 ;
        RECT 152.425 133.205 155.175 134.015 ;
        RECT 155.645 133.205 157.015 134.015 ;
        RECT 22.845 132.995 23.015 133.205 ;
        RECT 24.225 132.995 24.395 133.205 ;
        RECT 28.825 133.185 28.990 133.205 ;
        RECT 26.985 132.995 27.155 133.185 ;
        RECT 27.455 133.040 27.615 133.150 ;
        RECT 28.370 132.995 28.540 133.185 ;
        RECT 28.825 133.015 28.995 133.185 ;
        RECT 29.745 132.995 29.915 133.185 ;
        RECT 31.125 133.015 31.295 133.205 ;
        RECT 31.580 133.015 31.750 133.205 ;
        RECT 32.965 133.015 33.135 133.205 ;
        RECT 37.115 133.040 37.275 133.150 ;
        RECT 38.025 132.995 38.195 133.185 ;
        RECT 39.405 133.015 39.575 133.205 ;
        RECT 39.865 133.015 40.035 133.205 ;
        RECT 43.545 133.185 43.685 133.205 ;
        RECT 43.545 133.015 43.715 133.185 ;
        RECT 46.305 132.995 46.475 133.185 ;
        RECT 46.765 132.995 46.935 133.185 ;
        RECT 47.225 133.015 47.395 133.205 ;
        RECT 47.685 133.015 47.855 133.205 ;
        RECT 49.065 132.995 49.235 133.185 ;
        RECT 50.905 133.015 51.075 133.185 ;
        RECT 51.365 133.015 51.535 133.205 ;
        RECT 51.055 132.995 51.075 133.015 ;
        RECT 22.705 132.185 24.075 132.995 ;
        RECT 24.085 132.185 25.915 132.995 ;
        RECT 25.925 132.215 27.295 132.995 ;
        RECT 28.225 132.085 29.575 132.995 ;
        RECT 29.605 132.315 36.915 132.995 ;
        RECT 37.885 132.315 45.195 132.995 ;
        RECT 33.120 132.095 34.030 132.315 ;
        RECT 35.565 132.085 36.915 132.315 ;
        RECT 41.400 132.095 42.310 132.315 ;
        RECT 43.845 132.085 45.195 132.315 ;
        RECT 45.245 132.215 46.615 132.995 ;
        RECT 46.625 132.185 48.455 132.995 ;
        RECT 48.475 132.125 48.905 132.910 ;
        RECT 48.925 132.185 50.755 132.995 ;
        RECT 51.055 132.315 53.505 132.995 ;
        RECT 53.665 132.765 53.835 133.185 ;
        RECT 55.965 133.015 56.135 133.205 ;
        RECT 56.425 133.015 56.595 133.205 ;
        RECT 57.805 132.995 57.975 133.185 ;
        RECT 60.105 133.015 60.275 133.205 ;
        RECT 61.485 132.995 61.655 133.185 ;
        RECT 61.945 133.015 62.115 133.205 ;
        RECT 64.705 133.015 64.875 133.185 ;
        RECT 64.705 132.995 64.870 133.015 ;
        RECT 65.440 132.995 65.610 133.185 ;
        RECT 67.465 133.015 67.635 133.205 ;
        RECT 69.305 132.995 69.475 133.185 ;
        RECT 70.220 133.045 70.340 133.155 ;
        RECT 70.685 133.015 70.855 133.205 ;
        RECT 72.065 133.015 72.235 133.205 ;
        RECT 72.985 132.995 73.155 133.185 ;
        RECT 74.825 132.995 74.995 133.185 ;
        RECT 76.205 133.015 76.375 133.185 ;
        RECT 76.225 132.995 76.375 133.015 ;
        RECT 78.505 132.995 78.675 133.185 ;
        RECT 79.425 133.015 79.595 133.205 ;
        RECT 82.185 132.995 82.355 133.185 ;
        RECT 86.780 133.045 86.900 133.155 ;
        RECT 87.245 132.995 87.415 133.185 ;
        RECT 87.705 132.995 87.875 133.185 ;
        RECT 89.545 133.015 89.715 133.205 ;
        RECT 90.000 133.045 90.120 133.155 ;
        RECT 90.465 133.015 90.635 133.205 ;
        RECT 91.845 133.015 92.015 133.205 ;
        RECT 95.065 132.995 95.235 133.185 ;
        RECT 95.520 133.045 95.640 133.155 ;
        RECT 95.985 133.015 96.155 133.205 ;
        RECT 96.905 133.015 97.075 133.185 ;
        RECT 97.370 133.015 97.540 133.205 ;
        RECT 98.745 133.015 98.915 133.205 ;
        RECT 104.265 133.185 104.435 133.205 ;
        RECT 99.215 133.040 99.375 133.150 ;
        RECT 96.925 132.995 97.075 133.015 ;
        RECT 100.585 132.995 100.755 133.185 ;
        RECT 104.265 133.015 104.440 133.185 ;
        RECT 106.565 133.015 106.735 133.185 ;
        RECT 107.020 133.045 107.140 133.155 ;
        RECT 104.270 132.995 104.440 133.015 ;
        RECT 106.570 132.995 106.735 133.015 ;
        RECT 108.865 132.995 109.035 133.185 ;
        RECT 110.245 133.015 110.415 133.205 ;
        RECT 110.705 133.015 110.875 133.205 ;
        RECT 112.540 133.045 112.660 133.155 ;
        RECT 113.005 132.995 113.175 133.185 ;
        RECT 113.465 133.015 113.635 133.205 ;
        RECT 116.225 132.995 116.395 133.205 ;
        RECT 123.585 132.995 123.755 133.205 ;
        RECT 124.960 133.045 125.080 133.155 ;
        RECT 125.420 133.015 125.590 133.205 ;
        RECT 126.815 133.185 126.975 133.205 ;
        RECT 126.350 132.995 126.520 133.185 ;
        RECT 126.805 133.015 126.975 133.185 ;
        RECT 130.025 132.995 130.195 133.185 ;
        RECT 131.405 132.995 131.575 133.185 ;
        RECT 132.785 132.995 132.955 133.185 ;
        RECT 133.245 133.015 133.415 133.205 ;
        RECT 133.705 133.015 133.875 133.205 ;
        RECT 136.920 133.045 137.040 133.155 ;
        RECT 137.385 132.995 137.555 133.185 ;
        RECT 138.305 133.015 138.475 133.205 ;
        RECT 139.245 133.185 139.395 133.205 ;
        RECT 139.225 133.015 139.395 133.185 ;
        RECT 141.990 132.995 142.160 133.185 ;
        RECT 142.440 133.045 142.560 133.155 ;
        RECT 142.900 132.995 143.070 133.185 ;
        RECT 144.285 132.995 144.455 133.185 ;
        RECT 144.740 133.015 144.910 133.205 ;
        RECT 145.205 133.015 145.375 133.205 ;
        RECT 145.665 133.015 145.835 133.185 ;
        RECT 145.670 132.995 145.835 133.015 ;
        RECT 151.185 132.995 151.355 133.185 ;
        RECT 152.565 133.015 152.735 133.205 ;
        RECT 155.325 133.155 155.495 133.185 ;
        RECT 155.320 133.045 155.495 133.155 ;
        RECT 155.325 132.995 155.495 133.045 ;
        RECT 156.705 132.995 156.875 133.205 ;
        RECT 54.945 132.765 57.655 132.995 ;
        RECT 51.545 132.085 53.505 132.315 ;
        RECT 53.560 132.315 57.655 132.765 ;
        RECT 53.560 132.085 54.935 132.315 ;
        RECT 56.705 132.085 57.655 132.315 ;
        RECT 57.665 132.185 61.335 132.995 ;
        RECT 61.345 132.215 62.715 132.995 ;
        RECT 63.035 132.315 64.870 132.995 ;
        RECT 65.025 132.315 68.925 132.995 ;
        RECT 63.035 132.085 63.965 132.315 ;
        RECT 65.025 132.085 65.955 132.315 ;
        RECT 69.165 132.185 72.835 132.995 ;
        RECT 72.845 132.185 74.215 132.995 ;
        RECT 74.235 132.125 74.665 132.910 ;
        RECT 74.685 132.185 76.055 132.995 ;
        RECT 76.225 132.175 78.155 132.995 ;
        RECT 78.365 132.185 82.035 132.995 ;
        RECT 77.205 132.085 78.155 132.175 ;
        RECT 82.055 132.085 84.785 132.995 ;
        RECT 84.815 132.085 87.545 132.995 ;
        RECT 87.565 132.315 94.875 132.995 ;
        RECT 91.080 132.095 91.990 132.315 ;
        RECT 93.525 132.085 94.875 132.315 ;
        RECT 94.925 132.185 96.755 132.995 ;
        RECT 96.925 132.175 98.855 132.995 ;
        RECT 97.905 132.085 98.855 132.175 ;
        RECT 99.995 132.125 100.425 132.910 ;
        RECT 100.445 132.185 104.115 132.995 ;
        RECT 104.125 132.085 106.335 132.995 ;
        RECT 106.570 132.315 108.405 132.995 ;
        RECT 107.475 132.085 108.405 132.315 ;
        RECT 108.725 132.185 112.395 132.995 ;
        RECT 112.865 132.085 116.075 132.995 ;
        RECT 116.085 132.315 123.395 132.995 ;
        RECT 119.600 132.095 120.510 132.315 ;
        RECT 122.045 132.085 123.395 132.315 ;
        RECT 123.445 132.185 125.275 132.995 ;
        RECT 125.755 132.125 126.185 132.910 ;
        RECT 126.205 132.315 129.790 132.995 ;
        RECT 126.205 132.085 127.125 132.315 ;
        RECT 129.895 132.085 131.245 132.995 ;
        RECT 131.265 132.185 132.635 132.995 ;
        RECT 132.645 132.085 136.775 132.995 ;
        RECT 137.355 132.315 140.820 132.995 ;
        RECT 139.900 132.085 140.820 132.315 ;
        RECT 140.925 132.085 142.275 132.995 ;
        RECT 142.785 132.085 144.135 132.995 ;
        RECT 144.145 132.185 145.515 132.995 ;
        RECT 145.670 132.315 147.505 132.995 ;
        RECT 146.575 132.085 147.505 132.315 ;
        RECT 147.920 132.315 151.385 132.995 ;
        RECT 147.920 132.085 148.840 132.315 ;
        RECT 151.515 132.125 151.945 132.910 ;
        RECT 152.060 132.315 155.525 132.995 ;
        RECT 152.060 132.085 152.980 132.315 ;
        RECT 155.645 132.185 157.015 132.995 ;
      LAYER nwell ;
        RECT 22.510 128.965 157.210 131.795 ;
      LAYER pwell ;
        RECT 22.705 127.765 24.075 128.575 ;
        RECT 27.600 128.445 28.510 128.665 ;
        RECT 30.045 128.445 31.395 128.675 ;
        RECT 24.085 127.765 31.395 128.445 ;
        RECT 31.445 127.765 35.115 128.575 ;
        RECT 35.595 127.850 36.025 128.635 ;
        RECT 36.045 127.765 39.715 128.575 ;
        RECT 40.185 128.445 41.105 128.675 ;
        RECT 47.380 128.445 48.290 128.665 ;
        RECT 49.825 128.445 51.175 128.675 ;
        RECT 54.740 128.445 55.650 128.665 ;
        RECT 57.185 128.445 58.535 128.675 ;
        RECT 40.185 127.765 43.770 128.445 ;
        RECT 43.865 127.765 51.175 128.445 ;
        RECT 51.225 127.765 58.535 128.445 ;
        RECT 58.605 127.765 59.955 128.675 ;
        RECT 59.965 127.765 61.335 128.575 ;
        RECT 61.355 127.850 61.785 128.635 ;
        RECT 65.320 128.445 66.230 128.665 ;
        RECT 67.765 128.445 69.115 128.675 ;
        RECT 72.680 128.445 73.590 128.665 ;
        RECT 75.125 128.445 76.475 128.675 ;
        RECT 79.180 128.445 80.100 128.675 ;
        RECT 61.805 127.765 69.115 128.445 ;
        RECT 69.165 127.765 76.475 128.445 ;
        RECT 76.635 127.765 80.100 128.445 ;
        RECT 80.515 128.445 81.445 128.675 ;
        RECT 80.515 127.765 82.350 128.445 ;
        RECT 82.505 127.765 83.855 128.675 ;
        RECT 84.345 127.765 85.695 128.675 ;
        RECT 85.725 127.765 87.095 128.575 ;
        RECT 87.115 127.850 87.545 128.635 ;
        RECT 87.565 127.765 93.075 128.575 ;
        RECT 93.085 127.765 94.915 128.575 ;
        RECT 101.660 128.445 102.570 128.665 ;
        RECT 104.105 128.445 105.455 128.675 ;
        RECT 108.160 128.445 109.080 128.675 ;
        RECT 110.325 128.585 111.275 128.675 ;
        RECT 95.385 127.765 97.215 128.445 ;
        RECT 98.145 127.765 105.455 128.445 ;
        RECT 105.615 127.765 109.080 128.445 ;
        RECT 109.345 127.765 111.275 128.585 ;
        RECT 111.485 127.765 112.855 128.545 ;
        RECT 112.875 127.850 113.305 128.635 ;
        RECT 113.325 127.765 118.835 128.575 ;
        RECT 118.845 127.765 124.355 128.575 ;
        RECT 124.365 127.765 129.875 128.575 ;
        RECT 129.885 127.765 131.255 128.575 ;
        RECT 134.780 128.445 135.690 128.665 ;
        RECT 137.225 128.445 138.575 128.675 ;
        RECT 131.265 127.765 138.575 128.445 ;
        RECT 138.635 127.850 139.065 128.635 ;
        RECT 139.085 127.765 140.915 128.575 ;
        RECT 141.020 128.445 141.940 128.675 ;
        RECT 145.655 128.445 146.585 128.675 ;
        RECT 141.020 127.765 144.485 128.445 ;
        RECT 144.750 127.765 146.585 128.445 ;
        RECT 146.905 127.765 148.275 128.575 ;
        RECT 151.800 128.445 152.710 128.665 ;
        RECT 154.245 128.445 155.595 128.675 ;
        RECT 148.285 127.765 155.595 128.445 ;
        RECT 155.645 127.765 157.015 128.575 ;
        RECT 22.845 127.555 23.015 127.765 ;
        RECT 24.225 127.555 24.395 127.765 ;
        RECT 27.900 127.605 28.020 127.715 ;
        RECT 28.365 127.555 28.535 127.745 ;
        RECT 30.205 127.555 30.375 127.745 ;
        RECT 31.585 127.575 31.755 127.765 ;
        RECT 32.960 127.605 33.080 127.715 ;
        RECT 33.425 127.555 33.595 127.745 ;
        RECT 35.260 127.605 35.380 127.715 ;
        RECT 22.705 126.745 24.075 127.555 ;
        RECT 24.085 126.745 27.755 127.555 ;
        RECT 28.240 126.645 30.055 127.555 ;
        RECT 30.065 126.745 32.815 127.555 ;
        RECT 33.285 126.875 35.575 127.555 ;
        RECT 35.725 127.525 35.895 127.745 ;
        RECT 36.185 127.575 36.355 127.765 ;
        RECT 38.485 127.555 38.655 127.745 ;
        RECT 39.860 127.605 39.980 127.715 ;
        RECT 40.330 127.575 40.500 127.765 ;
        RECT 43.545 127.575 43.715 127.745 ;
        RECT 44.005 127.575 44.175 127.765 ;
        RECT 43.565 127.555 43.715 127.575 ;
        RECT 45.845 127.555 46.015 127.745 ;
        RECT 36.925 127.525 38.305 127.555 ;
        RECT 34.655 126.645 35.575 126.875 ;
        RECT 35.600 126.845 38.305 127.525 ;
        RECT 38.345 126.875 43.160 127.555 ;
        RECT 36.925 126.645 38.305 126.845 ;
        RECT 43.565 126.735 45.495 127.555 ;
        RECT 45.705 126.745 48.455 127.555 ;
        RECT 49.070 127.525 49.240 127.745 ;
        RECT 51.365 127.575 51.535 127.765 ;
        RECT 58.720 127.745 58.890 127.765 ;
        RECT 51.200 127.525 52.135 127.555 ;
        RECT 52.290 127.525 52.460 127.745 ;
        RECT 55.965 127.555 56.135 127.745 ;
        RECT 58.720 127.575 58.895 127.745 ;
        RECT 60.105 127.575 60.275 127.765 ;
        RECT 61.945 127.575 62.115 127.765 ;
        RECT 62.415 127.600 62.575 127.710 ;
        RECT 58.725 127.555 58.895 127.575 ;
        RECT 63.325 127.555 63.495 127.745 ;
        RECT 67.925 127.555 68.095 127.745 ;
        RECT 68.385 127.555 68.555 127.745 ;
        RECT 69.305 127.575 69.475 127.765 ;
        RECT 73.900 127.605 74.020 127.715 ;
        RECT 74.825 127.555 74.995 127.745 ;
        RECT 76.665 127.575 76.835 127.765 ;
        RECT 82.185 127.745 82.350 127.765 ;
        RECT 78.500 127.555 78.670 127.745 ;
        RECT 78.965 127.555 79.135 127.745 ;
        RECT 82.185 127.575 82.355 127.745 ;
        RECT 82.650 127.575 82.820 127.765 ;
        RECT 84.020 127.605 84.140 127.715 ;
        RECT 84.490 127.575 84.660 127.765 ;
        RECT 85.865 127.575 86.035 127.765 ;
        RECT 87.705 127.575 87.875 127.765 ;
        RECT 89.545 127.555 89.715 127.745 ;
        RECT 90.005 127.555 90.175 127.745 ;
        RECT 91.385 127.555 91.555 127.745 ;
        RECT 93.225 127.575 93.395 127.765 ;
        RECT 95.060 127.605 95.180 127.715 ;
        RECT 96.905 127.575 97.075 127.765 ;
        RECT 97.375 127.610 97.535 127.720 ;
        RECT 98.285 127.575 98.455 127.765 ;
        RECT 98.745 127.555 98.915 127.745 ;
        RECT 103.805 127.555 103.975 127.745 ;
        RECT 104.270 127.555 104.440 127.745 ;
        RECT 105.645 127.575 105.815 127.765 ;
        RECT 109.345 127.745 109.495 127.765 ;
        RECT 109.325 127.575 109.495 127.745 ;
        RECT 111.625 127.575 111.795 127.765 ;
        RECT 113.465 127.575 113.635 127.765 ;
        RECT 114.845 127.555 115.015 127.745 ;
        RECT 115.305 127.555 115.475 127.745 ;
        RECT 118.985 127.575 119.155 127.765 ;
        RECT 122.660 127.605 122.780 127.715 ;
        RECT 54.865 127.525 55.815 127.555 ;
        RECT 44.545 126.645 45.495 126.735 ;
        RECT 48.475 126.685 48.905 127.470 ;
        RECT 49.070 127.325 52.135 127.525 ;
        RECT 48.925 126.845 52.135 127.325 ;
        RECT 52.145 126.845 55.815 127.525 ;
        RECT 48.925 126.645 49.855 126.845 ;
        RECT 51.185 126.645 52.135 126.845 ;
        RECT 54.865 126.645 55.815 126.845 ;
        RECT 55.825 126.745 58.575 127.555 ;
        RECT 58.695 126.875 62.160 127.555 ;
        RECT 61.240 126.645 62.160 126.875 ;
        RECT 63.285 126.645 66.395 127.555 ;
        RECT 66.405 126.875 68.235 127.555 ;
        RECT 66.405 126.645 67.750 126.875 ;
        RECT 68.245 126.745 73.755 127.555 ;
        RECT 74.235 126.685 74.665 127.470 ;
        RECT 74.685 126.745 76.515 127.555 ;
        RECT 76.605 126.645 78.815 127.555 ;
        RECT 78.825 126.875 86.135 127.555 ;
        RECT 82.340 126.655 83.250 126.875 ;
        RECT 84.785 126.645 86.135 126.875 ;
        RECT 86.280 126.875 89.745 127.555 ;
        RECT 86.280 126.645 87.200 126.875 ;
        RECT 89.865 126.745 91.235 127.555 ;
        RECT 91.245 126.875 98.555 127.555 ;
        RECT 94.760 126.655 95.670 126.875 ;
        RECT 97.205 126.645 98.555 126.875 ;
        RECT 98.605 126.745 99.975 127.555 ;
        RECT 99.995 126.685 100.425 127.470 ;
        RECT 100.540 126.875 104.005 127.555 ;
        RECT 104.125 126.875 107.710 127.555 ;
        RECT 107.845 126.875 115.155 127.555 ;
        RECT 115.165 126.875 122.475 127.555 ;
        RECT 123.130 127.525 123.300 127.745 ;
        RECT 124.505 127.575 124.675 127.765 ;
        RECT 126.345 127.555 126.515 127.745 ;
        RECT 130.025 127.575 130.195 127.765 ;
        RECT 131.405 127.555 131.575 127.765 ;
        RECT 133.245 127.555 133.415 127.745 ;
        RECT 137.840 127.555 138.010 127.745 ;
        RECT 138.305 127.555 138.475 127.745 ;
        RECT 139.225 127.575 139.395 127.765 ;
        RECT 144.285 127.575 144.455 127.765 ;
        RECT 144.750 127.745 144.915 127.765 ;
        RECT 144.745 127.575 144.915 127.745 ;
        RECT 145.675 127.600 145.835 127.710 ;
        RECT 146.585 127.555 146.755 127.745 ;
        RECT 147.045 127.575 147.215 127.765 ;
        RECT 148.425 127.575 148.595 127.765 ;
        RECT 152.110 127.555 152.280 127.745 ;
        RECT 156.705 127.555 156.875 127.765 ;
        RECT 124.790 127.525 125.735 127.555 ;
        RECT 100.540 126.645 101.460 126.875 ;
        RECT 104.125 126.645 105.045 126.875 ;
        RECT 107.845 126.645 109.195 126.875 ;
        RECT 110.730 126.655 111.640 126.875 ;
        RECT 118.680 126.655 119.590 126.875 ;
        RECT 121.125 126.645 122.475 126.875 ;
        RECT 122.985 126.845 125.735 127.525 ;
        RECT 124.790 126.645 125.735 126.845 ;
        RECT 125.755 126.685 126.185 127.470 ;
        RECT 126.205 126.875 131.020 127.555 ;
        RECT 131.265 126.875 133.095 127.555 ;
        RECT 131.750 126.645 133.095 126.875 ;
        RECT 133.105 126.745 134.475 127.555 ;
        RECT 134.680 126.645 138.155 127.555 ;
        RECT 138.165 126.875 145.475 127.555 ;
        RECT 146.445 126.875 151.260 127.555 ;
        RECT 141.680 126.655 142.590 126.875 ;
        RECT 144.125 126.645 145.475 126.875 ;
        RECT 151.515 126.685 151.945 127.470 ;
        RECT 151.965 126.645 155.440 127.555 ;
        RECT 155.645 126.745 157.015 127.555 ;
      LAYER nwell ;
        RECT 22.510 123.525 157.210 126.355 ;
      LAYER pwell ;
        RECT 22.705 122.325 24.075 123.135 ;
        RECT 27.600 123.005 28.510 123.225 ;
        RECT 30.045 123.005 31.395 123.235 ;
        RECT 24.085 122.325 31.395 123.005 ;
        RECT 31.540 123.005 32.460 123.235 ;
        RECT 31.540 122.325 35.005 123.005 ;
        RECT 35.595 122.410 36.025 123.195 ;
        RECT 36.085 123.005 37.435 123.235 ;
        RECT 38.970 123.005 39.880 123.225 ;
        RECT 44.525 123.145 45.475 123.235 ;
        RECT 36.085 122.325 43.395 123.005 ;
        RECT 44.525 122.325 46.455 123.145 ;
        RECT 46.625 122.325 52.135 123.135 ;
        RECT 52.605 122.325 53.955 123.235 ;
        RECT 53.985 122.325 59.495 123.135 ;
        RECT 59.505 123.005 60.850 123.235 ;
        RECT 59.505 122.325 61.335 123.005 ;
        RECT 61.355 122.410 61.785 123.195 ;
        RECT 62.290 123.005 63.635 123.235 ;
        RECT 64.130 123.005 65.475 123.235 ;
        RECT 61.805 122.325 63.635 123.005 ;
        RECT 63.645 122.325 65.475 123.005 ;
        RECT 65.485 122.325 68.235 123.135 ;
        RECT 68.285 123.005 69.635 123.235 ;
        RECT 71.170 123.005 72.080 123.225 ;
        RECT 75.915 123.005 76.845 123.235 ;
        RECT 68.285 122.325 75.595 123.005 ;
        RECT 75.915 122.325 77.750 123.005 ;
        RECT 77.905 122.325 80.655 123.135 ;
        RECT 80.675 122.325 83.405 123.235 ;
        RECT 83.425 123.005 84.345 123.235 ;
        RECT 83.425 122.325 85.715 123.005 ;
        RECT 85.745 122.325 87.095 123.235 ;
        RECT 87.115 122.410 87.545 123.195 ;
        RECT 88.485 122.325 93.300 123.005 ;
        RECT 93.555 122.325 96.285 123.235 ;
        RECT 96.305 123.005 97.225 123.235 ;
        RECT 96.305 122.325 98.595 123.005 ;
        RECT 98.605 122.325 100.435 123.135 ;
        RECT 101.000 123.005 101.920 123.235 ;
        RECT 101.000 122.325 104.465 123.005 ;
        RECT 104.595 122.325 107.325 123.235 ;
        RECT 107.345 122.325 110.095 123.135 ;
        RECT 110.115 122.325 112.845 123.235 ;
        RECT 112.875 122.410 113.305 123.195 ;
        RECT 115.980 123.005 116.900 123.235 ;
        RECT 113.435 122.325 116.900 123.005 ;
        RECT 117.005 123.005 117.925 123.235 ;
        RECT 119.765 123.035 120.695 123.235 ;
        RECT 122.030 123.035 122.975 123.235 ;
        RECT 117.005 122.325 119.295 123.005 ;
        RECT 119.765 122.555 122.975 123.035 ;
        RECT 119.905 122.355 122.975 122.555 ;
        RECT 22.845 122.115 23.015 122.325 ;
        RECT 24.225 122.115 24.395 122.325 ;
        RECT 26.060 122.165 26.180 122.275 ;
        RECT 29.745 122.115 29.915 122.305 ;
        RECT 30.205 122.115 30.375 122.305 ;
        RECT 22.705 121.305 24.075 122.115 ;
        RECT 24.085 121.305 25.915 122.115 ;
        RECT 26.480 121.435 29.945 122.115 ;
        RECT 26.480 121.205 27.400 121.435 ;
        RECT 30.065 121.305 31.435 122.115 ;
        RECT 31.590 122.085 31.760 122.305 ;
        RECT 34.805 122.115 34.975 122.325 ;
        RECT 35.260 122.165 35.380 122.275 ;
        RECT 37.565 122.115 37.735 122.305 ;
        RECT 38.940 122.165 39.060 122.275 ;
        RECT 40.320 122.115 40.490 122.305 ;
        RECT 40.785 122.115 40.955 122.305 ;
        RECT 43.085 122.135 43.255 122.325 ;
        RECT 46.305 122.305 46.455 122.325 ;
        RECT 43.555 122.170 43.715 122.280 ;
        RECT 46.305 122.135 46.475 122.305 ;
        RECT 46.765 122.135 46.935 122.325 ;
        RECT 48.140 122.165 48.260 122.275 ;
        RECT 49.065 122.115 49.235 122.305 ;
        RECT 51.820 122.115 51.990 122.305 ;
        RECT 52.285 122.275 52.455 122.305 ;
        RECT 52.280 122.165 52.455 122.275 ;
        RECT 52.285 122.115 52.455 122.165 ;
        RECT 52.750 122.135 52.920 122.325 ;
        RECT 54.125 122.135 54.295 122.325 ;
        RECT 59.645 122.115 59.815 122.305 ;
        RECT 61.025 122.135 61.195 122.325 ;
        RECT 61.945 122.135 62.115 122.325 ;
        RECT 63.785 122.135 63.955 122.325 ;
        RECT 65.625 122.135 65.795 122.325 ;
        RECT 67.005 122.115 67.175 122.305 ;
        RECT 69.765 122.115 69.935 122.305 ;
        RECT 73.455 122.160 73.615 122.270 ;
        RECT 75.285 122.135 75.455 122.325 ;
        RECT 77.585 122.305 77.750 122.325 ;
        RECT 75.740 122.115 75.910 122.305 ;
        RECT 76.205 122.115 76.375 122.305 ;
        RECT 77.585 122.135 77.755 122.305 ;
        RECT 78.045 122.135 78.215 122.325 ;
        RECT 80.805 122.135 80.975 122.325 ;
        RECT 81.725 122.115 81.895 122.305 ;
        RECT 85.405 122.135 85.575 122.325 ;
        RECT 86.780 122.305 86.950 122.325 ;
        RECT 86.780 122.135 86.955 122.305 ;
        RECT 86.785 122.115 86.955 122.135 ;
        RECT 87.245 122.115 87.415 122.305 ;
        RECT 87.715 122.170 87.875 122.280 ;
        RECT 88.625 122.135 88.795 122.325 ;
        RECT 88.630 122.115 88.795 122.135 ;
        RECT 92.765 122.115 92.935 122.305 ;
        RECT 93.220 122.165 93.340 122.275 ;
        RECT 93.685 122.135 93.855 122.325 ;
        RECT 96.905 122.115 97.075 122.305 ;
        RECT 97.365 122.115 97.535 122.305 ;
        RECT 98.285 122.135 98.455 122.325 ;
        RECT 98.745 122.135 98.915 122.325 ;
        RECT 100.585 122.275 100.755 122.305 ;
        RECT 100.580 122.165 100.755 122.275 ;
        RECT 100.585 122.115 100.755 122.165 ;
        RECT 101.965 122.115 102.135 122.305 ;
        RECT 104.265 122.135 104.435 122.325 ;
        RECT 104.725 122.135 104.895 122.325 ;
        RECT 107.485 122.135 107.655 122.325 ;
        RECT 109.320 122.165 109.440 122.275 ;
        RECT 109.785 122.115 109.955 122.305 ;
        RECT 110.245 122.135 110.415 122.325 ;
        RECT 113.465 122.135 113.635 122.325 ;
        RECT 115.305 122.115 115.475 122.305 ;
        RECT 115.775 122.160 115.935 122.270 ;
        RECT 118.985 122.135 119.155 122.325 ;
        RECT 119.440 122.165 119.560 122.275 ;
        RECT 119.905 122.135 120.075 122.355 ;
        RECT 122.030 122.325 122.975 122.355 ;
        RECT 122.985 123.005 124.330 123.235 ;
        RECT 122.985 122.325 124.815 123.005 ;
        RECT 124.825 122.325 126.195 123.135 ;
        RECT 128.025 123.005 128.955 123.235 ;
        RECT 132.480 123.005 133.390 123.225 ;
        RECT 134.925 123.005 136.275 123.235 ;
        RECT 126.205 122.325 128.955 123.005 ;
        RECT 128.965 122.325 136.275 123.005 ;
        RECT 136.635 123.005 137.565 123.235 ;
        RECT 136.635 122.325 138.470 123.005 ;
        RECT 138.635 122.410 139.065 123.195 ;
        RECT 139.180 123.005 140.100 123.235 ;
        RECT 142.765 123.035 143.710 123.235 ;
        RECT 139.180 122.325 142.645 123.005 ;
        RECT 142.765 122.355 145.515 123.035 ;
        RECT 142.765 122.325 143.710 122.355 ;
        RECT 123.585 122.115 123.755 122.305 ;
        RECT 124.505 122.135 124.675 122.325 ;
        RECT 124.965 122.115 125.135 122.325 ;
        RECT 125.420 122.165 125.540 122.275 ;
        RECT 126.345 122.135 126.515 122.325 ;
        RECT 127.270 122.115 127.440 122.305 ;
        RECT 127.725 122.135 127.895 122.305 ;
        RECT 129.105 122.135 129.275 122.325 ;
        RECT 138.305 122.305 138.470 122.325 ;
        RECT 127.730 122.115 127.895 122.135 ;
        RECT 133.245 122.115 133.415 122.305 ;
        RECT 133.710 122.115 133.880 122.305 ;
        RECT 138.305 122.135 138.475 122.305 ;
        RECT 140.600 122.115 140.770 122.305 ;
        RECT 142.445 122.135 142.615 122.325 ;
        RECT 144.285 122.115 144.455 122.305 ;
        RECT 145.200 122.135 145.370 122.355 ;
        RECT 145.525 122.325 147.355 123.135 ;
        RECT 150.880 123.005 151.790 123.225 ;
        RECT 153.325 123.005 154.675 123.235 ;
        RECT 147.365 122.325 154.675 123.005 ;
        RECT 155.645 122.325 157.015 123.135 ;
        RECT 145.665 122.135 145.835 122.325 ;
        RECT 147.505 122.135 147.675 122.325 ;
        RECT 147.965 122.115 148.135 122.305 ;
        RECT 33.720 122.085 34.655 122.115 ;
        RECT 31.590 121.885 34.655 122.085 ;
        RECT 31.445 121.405 34.655 121.885 ;
        RECT 31.445 121.205 32.375 121.405 ;
        RECT 33.705 121.205 34.655 121.405 ;
        RECT 34.675 121.205 37.405 122.115 ;
        RECT 37.425 121.335 38.795 122.115 ;
        RECT 39.285 121.205 40.635 122.115 ;
        RECT 40.645 121.435 47.955 122.115 ;
        RECT 44.160 121.215 45.070 121.435 ;
        RECT 46.605 121.205 47.955 121.435 ;
        RECT 48.475 121.245 48.905 122.030 ;
        RECT 48.925 121.305 50.295 122.115 ;
        RECT 50.305 121.205 52.135 122.115 ;
        RECT 52.145 121.435 59.455 122.115 ;
        RECT 59.505 121.435 66.815 122.115 ;
        RECT 55.660 121.215 56.570 121.435 ;
        RECT 58.105 121.205 59.455 121.435 ;
        RECT 63.020 121.215 63.930 121.435 ;
        RECT 65.465 121.205 66.815 121.435 ;
        RECT 66.875 121.205 69.605 122.115 ;
        RECT 69.735 121.435 73.200 122.115 ;
        RECT 72.280 121.205 73.200 121.435 ;
        RECT 74.235 121.245 74.665 122.030 ;
        RECT 74.705 121.205 76.055 122.115 ;
        RECT 76.065 121.305 81.575 122.115 ;
        RECT 81.585 121.305 83.415 122.115 ;
        RECT 83.520 121.435 86.985 122.115 ;
        RECT 83.520 121.205 84.440 121.435 ;
        RECT 87.105 121.305 88.475 122.115 ;
        RECT 88.630 121.435 90.465 122.115 ;
        RECT 89.535 121.205 90.465 121.435 ;
        RECT 90.785 121.435 93.075 122.115 ;
        RECT 93.640 121.435 97.105 122.115 ;
        RECT 90.785 121.205 91.705 121.435 ;
        RECT 93.640 121.205 94.560 121.435 ;
        RECT 97.235 121.205 99.965 122.115 ;
        RECT 99.995 121.245 100.425 122.030 ;
        RECT 100.445 121.305 101.815 122.115 ;
        RECT 101.825 121.435 109.135 122.115 ;
        RECT 109.755 121.435 113.220 122.115 ;
        RECT 105.340 121.215 106.250 121.435 ;
        RECT 107.785 121.205 109.135 121.435 ;
        RECT 112.300 121.205 113.220 121.435 ;
        RECT 113.325 121.435 115.615 122.115 ;
        RECT 116.585 121.435 123.895 122.115 ;
        RECT 113.325 121.205 114.245 121.435 ;
        RECT 116.585 121.205 117.935 121.435 ;
        RECT 119.470 121.215 120.380 121.435 ;
        RECT 123.905 121.335 125.275 122.115 ;
        RECT 125.755 121.245 126.185 122.030 ;
        RECT 126.205 121.205 127.555 122.115 ;
        RECT 127.730 121.435 129.565 122.115 ;
        RECT 128.635 121.205 129.565 121.435 ;
        RECT 129.980 121.435 133.445 122.115 ;
        RECT 129.980 121.205 130.900 121.435 ;
        RECT 133.565 121.205 137.040 122.115 ;
        RECT 137.440 121.205 140.915 122.115 ;
        RECT 141.020 121.435 144.485 122.115 ;
        RECT 144.700 121.435 148.165 122.115 ;
        RECT 148.285 122.085 149.230 122.115 ;
        RECT 150.720 122.085 150.890 122.305 ;
        RECT 151.180 122.165 151.300 122.275 ;
        RECT 154.875 122.170 155.035 122.280 ;
        RECT 155.325 122.115 155.495 122.305 ;
        RECT 156.705 122.115 156.875 122.325 ;
        RECT 141.020 121.205 141.940 121.435 ;
        RECT 144.700 121.205 145.620 121.435 ;
        RECT 148.285 121.405 151.035 122.085 ;
        RECT 148.285 121.205 149.230 121.405 ;
        RECT 151.515 121.245 151.945 122.030 ;
        RECT 152.060 121.435 155.525 122.115 ;
        RECT 152.060 121.205 152.980 121.435 ;
        RECT 155.645 121.305 157.015 122.115 ;
      LAYER nwell ;
        RECT 22.510 118.085 157.210 120.915 ;
      LAYER pwell ;
        RECT 22.705 116.885 24.075 117.695 ;
        RECT 24.085 116.885 26.835 117.695 ;
        RECT 26.845 116.885 29.595 117.795 ;
        RECT 29.620 116.885 31.435 117.795 ;
        RECT 31.445 116.885 32.815 117.695 ;
        RECT 32.825 116.885 34.195 117.665 ;
        RECT 34.205 116.885 35.575 117.695 ;
        RECT 35.595 116.970 36.025 117.755 ;
        RECT 36.055 116.885 38.785 117.795 ;
        RECT 38.805 116.885 40.635 117.695 ;
        RECT 40.645 116.885 43.565 117.795 ;
        RECT 45.670 117.595 47.070 117.795 ;
        RECT 43.865 116.915 47.070 117.595 ;
        RECT 50.200 117.565 51.120 117.795 ;
        RECT 52.825 117.705 53.775 117.795 ;
        RECT 22.845 116.675 23.015 116.885 ;
        RECT 24.225 116.675 24.395 116.885 ;
        RECT 26.985 116.695 27.155 116.885 ;
        RECT 29.745 116.695 29.915 116.885 ;
        RECT 31.585 116.675 31.755 116.885 ;
        RECT 33.885 116.695 34.055 116.885 ;
        RECT 34.345 116.695 34.515 116.885 ;
        RECT 36.185 116.695 36.355 116.885 ;
        RECT 38.945 116.675 39.115 116.885 ;
        RECT 40.325 116.675 40.495 116.865 ;
        RECT 40.790 116.695 40.960 116.885 ;
        RECT 44.010 116.835 44.180 116.915 ;
        RECT 45.670 116.885 47.070 116.915 ;
        RECT 47.655 116.885 51.120 117.565 ;
        RECT 51.845 116.885 53.775 117.705 ;
        RECT 53.985 116.885 55.815 117.795 ;
        RECT 55.825 116.885 61.335 117.695 ;
        RECT 61.355 116.970 61.785 117.755 ;
        RECT 61.805 116.885 63.635 117.695 ;
        RECT 65.015 117.565 65.935 117.795 ;
        RECT 63.645 116.885 65.935 117.565 ;
        RECT 66.040 117.565 66.960 117.795 ;
        RECT 66.040 116.885 69.505 117.565 ;
        RECT 69.635 116.885 72.365 117.795 ;
        RECT 72.385 117.565 73.305 117.795 ;
        RECT 79.120 117.565 80.030 117.785 ;
        RECT 81.565 117.565 82.915 117.795 ;
        RECT 72.385 116.885 74.675 117.565 ;
        RECT 75.605 116.885 82.915 117.565 ;
        RECT 82.965 117.565 83.885 117.795 ;
        RECT 82.965 116.885 85.255 117.565 ;
        RECT 85.265 116.885 86.615 117.795 ;
        RECT 87.115 116.970 87.545 117.755 ;
        RECT 91.080 117.565 91.990 117.785 ;
        RECT 93.525 117.565 94.875 117.795 ;
        RECT 99.360 117.565 100.270 117.785 ;
        RECT 101.805 117.565 103.155 117.795 ;
        RECT 87.565 116.885 94.875 117.565 ;
        RECT 95.845 116.885 103.155 117.565 ;
        RECT 103.205 116.885 106.875 117.695 ;
        RECT 106.885 117.565 107.805 117.795 ;
        RECT 106.885 116.885 110.470 117.565 ;
        RECT 111.495 116.885 112.845 117.795 ;
        RECT 112.875 116.970 113.305 117.755 ;
        RECT 116.840 117.565 117.750 117.785 ;
        RECT 119.285 117.565 120.635 117.795 ;
        RECT 113.325 116.885 120.635 117.565 ;
        RECT 120.705 116.885 122.055 117.795 ;
        RECT 122.065 116.885 123.435 117.695 ;
        RECT 126.960 117.565 127.870 117.785 ;
        RECT 129.405 117.565 130.755 117.795 ;
        RECT 123.445 116.885 130.755 117.565 ;
        RECT 130.805 116.885 134.935 117.795 ;
        RECT 135.040 117.565 135.960 117.795 ;
        RECT 135.040 116.885 138.505 117.565 ;
        RECT 138.635 116.970 139.065 117.755 ;
        RECT 139.125 117.565 140.475 117.795 ;
        RECT 142.010 117.565 142.920 117.785 ;
        RECT 139.125 116.885 146.435 117.565 ;
        RECT 146.445 116.885 148.275 117.695 ;
        RECT 151.800 117.565 152.710 117.785 ;
        RECT 154.245 117.565 155.595 117.795 ;
        RECT 148.285 116.885 155.595 117.565 ;
        RECT 155.645 116.885 157.015 117.695 ;
        RECT 44.000 116.725 44.180 116.835 ;
        RECT 47.220 116.725 47.340 116.835 ;
        RECT 44.010 116.695 44.180 116.725 ;
        RECT 47.685 116.675 47.855 116.885 ;
        RECT 51.845 116.865 51.995 116.885 ;
        RECT 48.140 116.725 48.260 116.835 ;
        RECT 49.065 116.675 49.235 116.865 ;
        RECT 51.360 116.725 51.480 116.835 ;
        RECT 51.825 116.695 51.995 116.865 ;
        RECT 54.130 116.695 54.300 116.885 ;
        RECT 55.965 116.695 56.135 116.885 ;
        RECT 59.645 116.675 59.815 116.865 ;
        RECT 61.945 116.695 62.115 116.885 ;
        RECT 63.785 116.695 63.955 116.885 ;
        RECT 67.465 116.675 67.635 116.865 ;
        RECT 67.925 116.675 68.095 116.865 ;
        RECT 69.305 116.695 69.475 116.885 ;
        RECT 72.065 116.695 72.235 116.885 ;
        RECT 73.445 116.675 73.615 116.865 ;
        RECT 73.900 116.725 74.020 116.835 ;
        RECT 74.365 116.695 74.535 116.885 ;
        RECT 74.825 116.675 74.995 116.865 ;
        RECT 75.745 116.695 75.915 116.885 ;
        RECT 77.585 116.675 77.755 116.865 ;
        RECT 80.345 116.675 80.515 116.865 ;
        RECT 84.945 116.695 85.115 116.885 ;
        RECT 85.410 116.695 85.580 116.885 ;
        RECT 86.780 116.725 86.900 116.835 ;
        RECT 87.705 116.695 87.875 116.885 ;
        RECT 88.175 116.720 88.335 116.830 ;
        RECT 89.085 116.675 89.255 116.865 ;
        RECT 91.845 116.675 92.015 116.865 ;
        RECT 94.605 116.675 94.775 116.865 ;
        RECT 95.065 116.675 95.235 116.865 ;
        RECT 95.985 116.695 96.155 116.885 ;
        RECT 97.820 116.725 97.940 116.835 ;
        RECT 99.660 116.675 99.830 116.865 ;
        RECT 100.585 116.675 100.755 116.865 ;
        RECT 103.345 116.695 103.515 116.885 ;
        RECT 106.105 116.675 106.275 116.865 ;
        RECT 107.030 116.695 107.200 116.885 ;
        RECT 109.780 116.725 109.900 116.835 ;
        RECT 110.245 116.675 110.415 116.865 ;
        RECT 110.715 116.730 110.875 116.840 ;
        RECT 112.545 116.695 112.715 116.885 ;
        RECT 113.465 116.695 113.635 116.885 ;
        RECT 121.740 116.865 121.910 116.885 ;
        RECT 116.225 116.675 116.395 116.865 ;
        RECT 116.685 116.675 116.855 116.865 ;
        RECT 121.740 116.695 121.915 116.865 ;
        RECT 121.745 116.675 121.915 116.695 ;
        RECT 122.205 116.675 122.375 116.885 ;
        RECT 123.585 116.695 123.755 116.885 ;
        RECT 126.355 116.720 126.515 116.830 ;
        RECT 22.705 115.865 24.075 116.675 ;
        RECT 24.085 115.995 31.395 116.675 ;
        RECT 31.445 115.995 38.755 116.675 ;
        RECT 27.600 115.775 28.510 115.995 ;
        RECT 30.045 115.765 31.395 115.995 ;
        RECT 34.960 115.775 35.870 115.995 ;
        RECT 37.405 115.765 38.755 115.995 ;
        RECT 38.805 115.865 40.175 116.675 ;
        RECT 40.265 115.765 43.715 116.675 ;
        RECT 44.420 115.995 47.885 116.675 ;
        RECT 44.420 115.765 45.340 115.995 ;
        RECT 48.475 115.805 48.905 116.590 ;
        RECT 48.925 115.995 56.235 116.675 ;
        RECT 52.440 115.775 53.350 115.995 ;
        RECT 54.885 115.765 56.235 115.995 ;
        RECT 56.380 115.995 59.845 116.675 ;
        RECT 60.045 115.995 67.775 116.675 ;
        RECT 67.785 115.995 70.075 116.675 ;
        RECT 56.380 115.765 57.300 115.995 ;
        RECT 60.045 115.765 61.815 115.995 ;
        RECT 63.350 115.775 64.260 115.995 ;
        RECT 69.155 115.765 70.075 115.995 ;
        RECT 70.180 115.995 73.645 116.675 ;
        RECT 70.180 115.765 71.100 115.995 ;
        RECT 74.235 115.805 74.665 116.590 ;
        RECT 74.695 115.765 77.425 116.675 ;
        RECT 77.455 115.765 80.185 116.675 ;
        RECT 80.205 115.995 87.935 116.675 ;
        RECT 83.720 115.775 84.630 115.995 ;
        RECT 86.165 115.765 87.935 115.995 ;
        RECT 88.955 115.765 91.685 116.675 ;
        RECT 91.705 115.865 93.075 116.675 ;
        RECT 93.085 115.995 94.915 116.675 ;
        RECT 94.925 115.865 97.675 116.675 ;
        RECT 98.145 115.765 99.975 116.675 ;
        RECT 99.995 115.805 100.425 116.590 ;
        RECT 100.445 115.865 105.955 116.675 ;
        RECT 105.965 115.865 109.635 116.675 ;
        RECT 110.215 115.995 113.680 116.675 ;
        RECT 112.760 115.765 113.680 115.995 ;
        RECT 113.795 115.765 116.525 116.675 ;
        RECT 116.545 115.865 118.375 116.675 ;
        RECT 118.480 115.995 121.945 116.675 ;
        RECT 118.480 115.765 119.400 115.995 ;
        RECT 122.065 115.865 125.735 116.675 ;
        RECT 127.125 116.645 128.080 116.675 ;
        RECT 129.110 116.645 129.280 116.865 ;
        RECT 129.565 116.645 129.735 116.865 ;
        RECT 130.945 116.695 131.115 116.885 ;
        RECT 134.625 116.695 134.795 116.865 ;
        RECT 135.085 116.695 135.255 116.865 ;
        RECT 134.625 116.675 134.790 116.695 ;
        RECT 131.690 116.645 132.635 116.675 ;
        RECT 125.755 115.805 126.185 116.590 ;
        RECT 127.125 115.965 129.405 116.645 ;
        RECT 129.565 116.445 132.635 116.645 ;
        RECT 129.425 115.965 132.635 116.445 ;
        RECT 127.125 115.765 128.080 115.965 ;
        RECT 129.425 115.765 130.355 115.965 ;
        RECT 131.690 115.765 132.635 115.965 ;
        RECT 132.955 115.995 134.790 116.675 ;
        RECT 135.090 116.675 135.255 116.695 ;
        RECT 137.385 116.675 137.555 116.865 ;
        RECT 138.305 116.695 138.475 116.885 ;
        RECT 141.065 116.695 141.235 116.865 ;
        RECT 141.065 116.675 141.230 116.695 ;
        RECT 141.525 116.675 141.695 116.865 ;
        RECT 142.905 116.675 143.075 116.865 ;
        RECT 146.125 116.695 146.295 116.885 ;
        RECT 146.585 116.865 146.755 116.885 ;
        RECT 146.585 116.695 146.760 116.865 ;
        RECT 148.425 116.695 148.595 116.885 ;
        RECT 146.590 116.675 146.760 116.695 ;
        RECT 150.265 116.675 150.435 116.865 ;
        RECT 152.110 116.675 152.280 116.865 ;
        RECT 156.705 116.675 156.875 116.885 ;
        RECT 135.090 115.995 136.925 116.675 ;
        RECT 137.245 115.995 139.075 116.675 ;
        RECT 139.395 115.995 141.230 116.675 ;
        RECT 132.955 115.765 133.885 115.995 ;
        RECT 135.995 115.765 136.925 115.995 ;
        RECT 139.395 115.765 140.325 115.995 ;
        RECT 141.385 115.865 142.755 116.675 ;
        RECT 142.875 115.995 146.340 116.675 ;
        RECT 145.420 115.765 146.340 115.995 ;
        RECT 146.445 115.765 149.920 116.675 ;
        RECT 150.125 115.865 151.495 116.675 ;
        RECT 151.515 115.805 151.945 116.590 ;
        RECT 151.965 115.765 155.440 116.675 ;
        RECT 155.645 115.865 157.015 116.675 ;
      LAYER nwell ;
        RECT 22.510 112.645 157.210 115.475 ;
      LAYER pwell ;
        RECT 22.705 111.445 24.075 112.255 ;
        RECT 24.085 111.445 25.915 112.255 ;
        RECT 26.480 112.125 27.400 112.355 ;
        RECT 30.160 112.125 31.080 112.355 ;
        RECT 26.480 111.445 29.945 112.125 ;
        RECT 30.160 111.445 33.625 112.125 ;
        RECT 33.745 111.445 35.575 112.255 ;
        RECT 35.595 111.530 36.025 112.315 ;
        RECT 36.045 112.125 36.965 112.355 ;
        RECT 41.860 112.125 42.770 112.345 ;
        RECT 44.305 112.125 45.655 112.355 ;
        RECT 36.045 111.445 38.335 112.125 ;
        RECT 38.345 111.445 45.655 112.125 ;
        RECT 45.705 111.445 47.075 112.255 ;
        RECT 47.105 111.445 48.455 112.355 ;
        RECT 48.465 111.445 51.215 112.255 ;
        RECT 51.320 112.125 52.240 112.355 ;
        RECT 54.905 112.125 55.825 112.355 ;
        RECT 51.320 111.445 54.785 112.125 ;
        RECT 54.905 111.445 57.195 112.125 ;
        RECT 57.205 111.445 59.035 112.355 ;
        RECT 59.045 111.445 60.875 112.255 ;
        RECT 61.355 111.530 61.785 112.315 ;
        RECT 61.805 111.445 67.645 112.355 ;
        RECT 67.825 112.125 69.175 112.355 ;
        RECT 70.710 112.125 71.620 112.345 ;
        RECT 67.825 111.445 75.135 112.125 ;
        RECT 75.145 111.445 80.655 112.255 ;
        RECT 80.675 111.445 83.405 112.355 ;
        RECT 83.425 112.125 84.345 112.355 ;
        RECT 83.425 111.445 85.715 112.125 ;
        RECT 85.725 111.445 87.095 112.255 ;
        RECT 87.115 111.530 87.545 112.315 ;
        RECT 87.565 111.445 91.235 112.255 ;
        RECT 92.615 112.125 93.535 112.355 ;
        RECT 97.060 112.125 97.970 112.345 ;
        RECT 99.505 112.125 101.275 112.355 ;
        RECT 105.800 112.125 106.710 112.345 ;
        RECT 108.245 112.125 109.595 112.355 ;
        RECT 91.245 111.445 93.535 112.125 ;
        RECT 93.545 111.445 101.275 112.125 ;
        RECT 102.285 111.445 109.595 112.125 ;
        RECT 109.645 112.125 110.565 112.355 ;
        RECT 109.645 111.445 111.935 112.125 ;
        RECT 112.875 111.530 113.305 112.315 ;
        RECT 113.325 111.445 114.695 112.255 ;
        RECT 114.705 112.125 115.625 112.355 ;
        RECT 114.705 111.445 116.995 112.125 ;
        RECT 117.475 111.445 118.825 112.355 ;
        RECT 122.420 112.125 123.340 112.355 ;
        RECT 119.875 111.445 123.340 112.125 ;
        RECT 123.445 111.445 125.275 112.355 ;
        RECT 125.285 111.445 127.115 112.255 ;
        RECT 127.585 111.445 129.415 112.355 ;
        RECT 130.475 112.125 131.405 112.355 ;
        RECT 129.570 111.445 131.405 112.125 ;
        RECT 131.920 111.445 135.395 112.355 ;
        RECT 136.915 112.125 137.845 112.355 ;
        RECT 136.010 111.445 137.845 112.125 ;
        RECT 138.635 111.530 139.065 112.315 ;
        RECT 139.180 112.125 140.100 112.355 ;
        RECT 142.765 112.125 144.110 112.355 ;
        RECT 139.180 111.445 142.645 112.125 ;
        RECT 142.765 111.445 144.595 112.125 ;
        RECT 144.800 111.445 148.275 112.355 ;
        RECT 151.800 112.125 152.710 112.345 ;
        RECT 154.245 112.125 155.595 112.355 ;
        RECT 148.285 111.445 155.595 112.125 ;
        RECT 155.645 111.445 157.015 112.255 ;
        RECT 22.845 111.235 23.015 111.445 ;
        RECT 24.225 111.235 24.395 111.445 ;
        RECT 26.060 111.285 26.180 111.395 ;
        RECT 26.985 111.235 27.155 111.425 ;
        RECT 29.745 111.235 29.915 111.445 ;
        RECT 31.580 111.285 31.700 111.395 ;
        RECT 33.425 111.255 33.595 111.445 ;
        RECT 33.885 111.255 34.055 111.445 ;
        RECT 22.705 110.425 24.075 111.235 ;
        RECT 24.085 110.425 26.835 111.235 ;
        RECT 26.845 110.325 29.595 111.235 ;
        RECT 29.605 110.425 31.435 111.235 ;
        RECT 31.905 111.205 32.840 111.235 ;
        RECT 34.800 111.205 34.970 111.425 ;
        RECT 35.265 111.235 35.435 111.425 ;
        RECT 38.025 111.255 38.195 111.445 ;
        RECT 38.485 111.255 38.655 111.445 ;
        RECT 40.785 111.235 40.955 111.425 ;
        RECT 45.845 111.255 46.015 111.445 ;
        RECT 46.305 111.235 46.475 111.425 ;
        RECT 48.140 111.255 48.310 111.445 ;
        RECT 48.605 111.255 48.775 111.445 ;
        RECT 49.065 111.235 49.235 111.425 ;
        RECT 52.745 111.255 52.915 111.425 ;
        RECT 53.200 111.285 53.320 111.395 ;
        RECT 54.585 111.255 54.755 111.445 ;
        RECT 52.745 111.235 52.910 111.255 ;
        RECT 55.040 111.235 55.210 111.425 ;
        RECT 55.505 111.235 55.675 111.425 ;
        RECT 56.885 111.255 57.055 111.445 ;
        RECT 58.720 111.425 58.890 111.445 ;
        RECT 58.720 111.255 58.895 111.425 ;
        RECT 59.185 111.255 59.355 111.445 ;
        RECT 61.020 111.285 61.140 111.395 ;
        RECT 61.945 111.255 62.115 111.445 ;
        RECT 64.255 111.280 64.415 111.390 ;
        RECT 58.725 111.235 58.895 111.255 ;
        RECT 65.165 111.235 65.335 111.425 ;
        RECT 68.380 111.235 68.550 111.425 ;
        RECT 68.855 111.280 69.015 111.390 ;
        RECT 72.065 111.235 72.235 111.425 ;
        RECT 72.525 111.235 72.695 111.425 ;
        RECT 74.825 111.395 74.995 111.445 ;
        RECT 74.820 111.285 74.995 111.395 ;
        RECT 74.825 111.255 74.995 111.285 ;
        RECT 75.285 111.235 75.455 111.445 ;
        RECT 80.805 111.255 80.975 111.445 ;
        RECT 82.645 111.235 82.815 111.425 ;
        RECT 85.405 111.395 85.575 111.445 ;
        RECT 85.400 111.285 85.575 111.395 ;
        RECT 85.405 111.255 85.575 111.285 ;
        RECT 85.865 111.235 86.035 111.445 ;
        RECT 87.705 111.255 87.875 111.445 ;
        RECT 91.385 111.255 91.555 111.445 ;
        RECT 93.685 111.255 93.855 111.445 ;
        RECT 96.445 111.235 96.615 111.425 ;
        RECT 96.905 111.235 97.075 111.425 ;
        RECT 99.660 111.285 99.780 111.395 ;
        RECT 100.590 111.235 100.760 111.425 ;
        RECT 101.515 111.290 101.675 111.400 ;
        RECT 101.965 111.235 102.135 111.425 ;
        RECT 102.425 111.255 102.595 111.445 ;
        RECT 104.725 111.235 104.895 111.425 ;
        RECT 108.405 111.235 108.575 111.425 ;
        RECT 108.865 111.235 109.035 111.425 ;
        RECT 111.625 111.255 111.795 111.445 ;
        RECT 112.095 111.290 112.255 111.400 ;
        RECT 113.465 111.255 113.635 111.445 ;
        RECT 114.365 111.235 114.535 111.425 ;
        RECT 116.685 111.255 116.855 111.445 ;
        RECT 117.140 111.285 117.260 111.395 ;
        RECT 118.525 111.255 118.695 111.445 ;
        RECT 118.995 111.290 119.155 111.400 ;
        RECT 119.905 111.255 120.075 111.445 ;
        RECT 124.960 111.255 125.130 111.445 ;
        RECT 125.425 111.235 125.595 111.445 ;
        RECT 126.345 111.235 126.515 111.425 ;
        RECT 127.260 111.285 127.380 111.395 ;
        RECT 127.730 111.255 127.900 111.445 ;
        RECT 129.570 111.425 129.735 111.445 ;
        RECT 129.105 111.235 129.275 111.425 ;
        RECT 129.565 111.255 129.735 111.425 ;
        RECT 132.785 111.235 132.955 111.425 ;
        RECT 135.080 111.255 135.250 111.445 ;
        RECT 136.010 111.425 136.175 111.445 ;
        RECT 135.540 111.285 135.660 111.395 ;
        RECT 136.005 111.255 136.175 111.425 ;
        RECT 138.300 111.285 138.420 111.395 ;
        RECT 142.445 111.255 142.615 111.445 ;
        RECT 144.285 111.255 144.455 111.445 ;
        RECT 147.045 111.235 147.215 111.425 ;
        RECT 147.960 111.255 148.130 111.445 ;
        RECT 148.425 111.255 148.595 111.445 ;
        RECT 150.725 111.235 150.895 111.425 ;
        RECT 151.180 111.285 151.300 111.395 ;
        RECT 155.325 111.235 155.495 111.425 ;
        RECT 156.705 111.235 156.875 111.445 ;
        RECT 31.905 111.005 34.970 111.205 ;
        RECT 31.905 110.525 35.115 111.005 ;
        RECT 31.905 110.325 32.855 110.525 ;
        RECT 34.185 110.325 35.115 110.525 ;
        RECT 35.125 110.425 40.635 111.235 ;
        RECT 40.645 110.425 46.155 111.235 ;
        RECT 46.165 110.425 47.995 111.235 ;
        RECT 48.475 110.365 48.905 111.150 ;
        RECT 48.925 110.425 50.755 111.235 ;
        RECT 51.075 110.555 52.910 111.235 ;
        RECT 51.075 110.325 52.005 110.555 ;
        RECT 53.525 110.325 55.355 111.235 ;
        RECT 55.465 110.325 58.575 111.235 ;
        RECT 58.585 110.425 64.095 111.235 ;
        RECT 65.025 110.555 67.315 111.235 ;
        RECT 66.395 110.325 67.315 110.555 ;
        RECT 67.345 110.325 68.695 111.235 ;
        RECT 69.635 110.325 72.365 111.235 ;
        RECT 72.385 110.425 74.215 111.235 ;
        RECT 74.235 110.365 74.665 111.150 ;
        RECT 75.145 110.555 82.455 111.235 ;
        RECT 78.660 110.335 79.570 110.555 ;
        RECT 81.105 110.325 82.455 110.555 ;
        RECT 82.505 110.425 85.255 111.235 ;
        RECT 85.725 110.555 93.035 111.235 ;
        RECT 89.240 110.335 90.150 110.555 ;
        RECT 91.685 110.325 93.035 110.555 ;
        RECT 93.180 110.555 96.645 111.235 ;
        RECT 93.180 110.325 94.100 110.555 ;
        RECT 96.775 110.325 99.505 111.235 ;
        RECT 99.995 110.365 100.425 111.150 ;
        RECT 100.445 110.325 101.795 111.235 ;
        RECT 101.825 110.425 104.575 111.235 ;
        RECT 104.595 110.325 107.325 111.235 ;
        RECT 107.355 110.325 108.705 111.235 ;
        RECT 108.725 110.425 114.235 111.235 ;
        RECT 114.255 110.555 118.280 111.235 ;
        RECT 118.425 110.555 125.735 111.235 ;
        RECT 114.255 110.325 115.600 110.555 ;
        RECT 118.425 110.325 119.775 110.555 ;
        RECT 121.310 110.335 122.220 110.555 ;
        RECT 125.755 110.365 126.185 111.150 ;
        RECT 126.205 110.425 128.955 111.235 ;
        RECT 129.075 110.555 132.540 111.235 ;
        RECT 132.645 110.555 139.955 111.235 ;
        RECT 131.620 110.325 132.540 110.555 ;
        RECT 136.160 110.335 137.070 110.555 ;
        RECT 138.605 110.325 139.955 110.555 ;
        RECT 140.045 110.555 147.355 111.235 ;
        RECT 147.460 110.555 150.925 111.235 ;
        RECT 140.045 110.325 141.395 110.555 ;
        RECT 142.930 110.335 143.840 110.555 ;
        RECT 147.460 110.325 148.380 110.555 ;
        RECT 151.515 110.365 151.945 111.150 ;
        RECT 152.060 110.555 155.525 111.235 ;
        RECT 152.060 110.325 152.980 110.555 ;
        RECT 155.645 110.425 157.015 111.235 ;
      LAYER nwell ;
        RECT 22.510 107.205 157.210 110.035 ;
      LAYER pwell ;
        RECT 22.705 106.005 24.075 106.815 ;
        RECT 24.085 106.005 29.595 106.815 ;
        RECT 29.605 106.005 32.355 106.815 ;
        RECT 32.375 106.005 35.105 106.915 ;
        RECT 35.595 106.090 36.025 106.875 ;
        RECT 36.045 106.005 37.860 106.915 ;
        RECT 37.885 106.005 39.715 106.815 ;
        RECT 39.725 106.005 41.075 106.915 ;
        RECT 41.200 106.685 42.120 106.915 ;
        RECT 45.705 106.685 46.625 106.915 ;
        RECT 41.200 106.005 44.665 106.685 ;
        RECT 45.705 106.005 47.995 106.685 ;
        RECT 48.005 106.005 50.755 106.915 ;
        RECT 51.545 106.685 53.505 106.915 ;
        RECT 51.055 106.005 53.505 106.685 ;
        RECT 54.545 106.005 57.655 106.915 ;
        RECT 57.665 106.005 61.335 106.815 ;
        RECT 61.355 106.090 61.785 106.875 ;
        RECT 61.805 106.005 63.175 106.815 ;
        RECT 63.185 106.005 66.855 106.915 ;
        RECT 66.865 106.005 68.215 106.915 ;
        RECT 68.245 106.005 70.075 106.815 ;
        RECT 70.555 106.005 73.285 106.915 ;
        RECT 76.880 106.685 77.800 106.915 ;
        RECT 74.335 106.005 77.800 106.685 ;
        RECT 77.905 106.005 81.575 106.915 ;
        RECT 81.680 106.685 82.600 106.915 ;
        RECT 81.680 106.005 85.145 106.685 ;
        RECT 85.265 106.005 86.615 106.915 ;
        RECT 87.115 106.090 87.545 106.875 ;
        RECT 88.035 106.005 90.765 106.915 ;
        RECT 90.785 106.685 91.705 106.915 ;
        RECT 90.785 106.005 93.075 106.685 ;
        RECT 93.085 106.005 95.835 106.815 ;
        RECT 96.305 106.005 99.975 106.915 ;
        RECT 101.355 106.685 102.275 106.915 ;
        RECT 99.985 106.005 102.275 106.685 ;
        RECT 102.380 106.685 103.300 106.915 ;
        RECT 105.965 106.685 106.885 106.915 ;
        RECT 102.380 106.005 105.845 106.685 ;
        RECT 105.965 106.005 109.550 106.685 ;
        RECT 109.655 106.005 112.385 106.915 ;
        RECT 112.875 106.090 113.305 106.875 ;
        RECT 116.840 106.685 117.750 106.905 ;
        RECT 119.285 106.685 120.635 106.915 ;
        RECT 113.325 106.005 120.635 106.685 ;
        RECT 120.700 106.005 122.515 106.915 ;
        RECT 123.025 106.685 124.375 106.915 ;
        RECT 125.910 106.685 126.820 106.905 ;
        RECT 133.000 106.685 133.920 106.915 ;
        RECT 123.025 106.005 130.335 106.685 ;
        RECT 130.455 106.005 133.920 106.685 ;
        RECT 134.025 106.005 137.500 106.915 ;
        RECT 138.635 106.090 139.065 106.875 ;
        RECT 139.085 106.005 140.915 106.815 ;
        RECT 143.580 106.685 144.500 106.915 ;
        RECT 141.035 106.005 144.500 106.685 ;
        RECT 144.605 106.715 145.550 106.915 ;
        RECT 144.605 106.035 147.355 106.715 ;
        RECT 150.880 106.685 151.790 106.905 ;
        RECT 153.325 106.685 154.675 106.915 ;
        RECT 144.605 106.005 145.550 106.035 ;
        RECT 22.845 105.795 23.015 106.005 ;
        RECT 24.225 105.795 24.395 106.005 ;
        RECT 29.745 105.815 29.915 106.005 ;
        RECT 33.420 105.795 33.590 105.985 ;
        RECT 33.885 105.795 34.055 105.985 ;
        RECT 34.805 105.815 34.975 106.005 ;
        RECT 35.260 105.845 35.380 105.955 ;
        RECT 37.565 105.815 37.735 106.005 ;
        RECT 38.025 105.815 38.195 106.005 ;
        RECT 40.790 105.815 40.960 106.005 ;
        RECT 41.245 105.795 41.415 105.985 ;
        RECT 44.465 105.815 44.635 106.005 ;
        RECT 44.935 105.850 45.095 105.960 ;
        RECT 47.685 105.815 47.855 106.005 ;
        RECT 48.145 105.815 48.315 106.005 ;
        RECT 51.055 105.985 51.075 106.005 ;
        RECT 54.585 105.985 54.755 106.005 ;
        RECT 49.065 105.795 49.235 105.985 ;
        RECT 50.905 105.795 51.075 105.985 ;
        RECT 53.675 105.850 53.835 105.960 ;
        RECT 54.580 105.815 54.755 105.985 ;
        RECT 54.580 105.795 54.750 105.815 ;
        RECT 56.885 105.795 57.055 105.985 ;
        RECT 57.805 105.815 57.975 106.005 ;
        RECT 61.945 105.985 62.115 106.005 ;
        RECT 60.565 105.795 60.735 105.985 ;
        RECT 61.035 105.840 61.195 105.950 ;
        RECT 61.935 105.815 62.115 105.985 ;
        RECT 63.330 105.815 63.500 106.005 ;
        RECT 67.010 105.985 67.180 106.005 ;
        RECT 65.160 105.845 65.280 105.955 ;
        RECT 61.935 105.795 62.105 105.815 ;
        RECT 66.540 105.795 66.710 105.985 ;
        RECT 67.005 105.815 67.180 105.985 ;
        RECT 68.385 105.815 68.555 106.005 ;
        RECT 70.220 105.845 70.340 105.955 ;
        RECT 70.685 105.815 70.855 106.005 ;
        RECT 73.455 105.850 73.615 105.960 ;
        RECT 74.365 105.815 74.535 106.005 ;
        RECT 67.005 105.795 67.175 105.815 ;
        RECT 76.665 105.795 76.835 105.985 ;
        RECT 77.120 105.845 77.240 105.955 ;
        RECT 77.585 105.795 77.755 105.985 ;
        RECT 78.050 105.815 78.220 106.005 ;
        RECT 84.945 105.985 85.115 106.005 ;
        RECT 82.185 105.795 82.355 105.985 ;
        RECT 82.645 105.795 82.815 105.985 ;
        RECT 84.480 105.845 84.600 105.955 ;
        RECT 84.945 105.815 85.120 105.985 ;
        RECT 85.410 105.815 85.580 106.005 ;
        RECT 84.950 105.795 85.120 105.815 ;
        RECT 86.325 105.795 86.495 105.985 ;
        RECT 86.780 105.845 86.900 105.955 ;
        RECT 87.700 105.845 87.820 105.955 ;
        RECT 88.165 105.815 88.335 106.005 ;
        RECT 91.840 105.845 91.960 105.955 ;
        RECT 92.295 105.795 92.465 105.985 ;
        RECT 92.765 105.815 92.935 106.005 ;
        RECT 93.225 105.815 93.395 106.005 ;
        RECT 95.980 105.845 96.100 105.955 ;
        RECT 96.450 105.815 96.620 106.005 ;
        RECT 98.745 105.795 98.915 105.985 ;
        RECT 99.215 105.840 99.375 105.950 ;
        RECT 100.125 105.815 100.295 106.005 ;
        RECT 100.590 105.795 100.760 105.985 ;
        RECT 105.645 105.815 105.815 106.005 ;
        RECT 106.110 105.815 106.280 106.005 ;
        RECT 108.865 105.795 109.035 105.985 ;
        RECT 109.335 105.840 109.495 105.950 ;
        RECT 109.785 105.815 109.955 106.005 ;
        RECT 112.545 105.955 112.715 105.985 ;
        RECT 112.540 105.845 112.715 105.955 ;
        RECT 112.545 105.795 112.715 105.845 ;
        RECT 113.465 105.815 113.635 106.005 ;
        RECT 114.845 105.795 115.015 105.985 ;
        RECT 115.305 105.795 115.475 105.985 ;
        RECT 120.365 105.795 120.535 105.985 ;
        RECT 120.825 105.795 120.995 106.005 ;
        RECT 122.660 105.845 122.780 105.955 ;
        RECT 124.505 105.795 124.675 105.985 ;
        RECT 126.345 105.795 126.515 105.985 ;
        RECT 128.185 105.815 128.355 105.985 ;
        RECT 130.025 105.815 130.195 106.005 ;
        RECT 130.485 105.985 130.655 106.005 ;
        RECT 130.485 105.815 130.660 105.985 ;
        RECT 134.170 105.815 134.340 106.005 ;
        RECT 128.190 105.795 128.355 105.815 ;
        RECT 130.490 105.795 130.660 105.815 ;
        RECT 137.380 105.795 137.550 105.985 ;
        RECT 137.845 105.795 138.015 105.985 ;
        RECT 139.225 105.815 139.395 106.005 ;
        RECT 141.065 105.815 141.235 106.005 ;
        RECT 144.740 105.795 144.910 105.985 ;
        RECT 147.040 105.815 147.210 106.035 ;
        RECT 147.365 106.005 154.675 106.685 ;
        RECT 155.645 106.005 157.015 106.815 ;
        RECT 147.505 105.815 147.675 106.005 ;
        RECT 148.425 105.795 148.595 105.985 ;
        RECT 150.725 105.815 150.895 105.985 ;
        RECT 151.180 105.845 151.300 105.955 ;
        RECT 154.875 105.850 155.035 105.960 ;
        RECT 150.725 105.795 150.890 105.815 ;
        RECT 155.325 105.795 155.495 105.985 ;
        RECT 156.705 105.795 156.875 106.005 ;
        RECT 22.705 104.985 24.075 105.795 ;
        RECT 24.085 104.985 29.595 105.795 ;
        RECT 30.815 104.885 33.735 105.795 ;
        RECT 33.745 105.115 41.055 105.795 ;
        RECT 41.105 105.115 48.415 105.795 ;
        RECT 37.260 104.895 38.170 105.115 ;
        RECT 39.705 104.885 41.055 105.115 ;
        RECT 44.620 104.895 45.530 105.115 ;
        RECT 47.065 104.885 48.415 105.115 ;
        RECT 48.475 104.925 48.905 105.710 ;
        RECT 48.925 104.985 50.755 105.795 ;
        RECT 50.875 105.115 54.340 105.795 ;
        RECT 53.420 104.885 54.340 105.115 ;
        RECT 54.465 104.885 55.815 105.795 ;
        RECT 55.835 104.885 57.185 105.795 ;
        RECT 57.300 105.115 60.765 105.795 ;
        RECT 57.300 104.885 58.220 105.115 ;
        RECT 61.805 104.885 65.015 105.795 ;
        RECT 65.505 104.885 66.855 105.795 ;
        RECT 66.865 105.115 74.175 105.795 ;
        RECT 70.380 104.895 71.290 105.115 ;
        RECT 72.825 104.885 74.175 105.115 ;
        RECT 74.235 104.925 74.665 105.710 ;
        RECT 74.685 105.115 76.975 105.795 ;
        RECT 74.685 104.885 75.605 105.115 ;
        RECT 77.455 104.885 80.185 105.795 ;
        RECT 80.205 105.115 82.495 105.795 ;
        RECT 80.205 104.885 81.125 105.115 ;
        RECT 82.505 104.985 84.335 105.795 ;
        RECT 84.805 104.885 86.155 105.795 ;
        RECT 86.185 104.985 91.695 105.795 ;
        RECT 92.165 104.885 95.375 105.795 ;
        RECT 95.480 105.115 98.945 105.795 ;
        RECT 95.480 104.885 96.400 105.115 ;
        RECT 99.995 104.925 100.425 105.710 ;
        RECT 100.445 104.885 101.795 105.795 ;
        RECT 101.865 105.115 109.175 105.795 ;
        RECT 101.865 104.885 103.215 105.115 ;
        RECT 104.750 104.895 105.660 105.115 ;
        RECT 110.115 104.885 112.845 105.795 ;
        RECT 112.865 105.115 115.155 105.795 ;
        RECT 112.865 104.885 113.785 105.115 ;
        RECT 115.165 104.985 116.995 105.795 ;
        RECT 117.100 105.115 120.565 105.795 ;
        RECT 117.100 104.885 118.020 105.115 ;
        RECT 120.685 104.985 124.355 105.795 ;
        RECT 124.365 104.985 125.735 105.795 ;
        RECT 125.755 104.925 126.185 105.710 ;
        RECT 126.205 104.985 128.035 105.795 ;
        RECT 128.190 105.115 130.025 105.795 ;
        RECT 129.095 104.885 130.025 105.115 ;
        RECT 130.345 104.885 133.820 105.795 ;
        RECT 134.220 104.885 137.695 105.795 ;
        RECT 137.815 105.115 141.280 105.795 ;
        RECT 140.360 104.885 141.280 105.115 ;
        RECT 141.580 104.885 145.055 105.795 ;
        RECT 145.160 105.115 148.625 105.795 ;
        RECT 149.055 105.115 150.890 105.795 ;
        RECT 145.160 104.885 146.080 105.115 ;
        RECT 149.055 104.885 149.985 105.115 ;
        RECT 151.515 104.925 151.945 105.710 ;
        RECT 152.060 105.115 155.525 105.795 ;
        RECT 152.060 104.885 152.980 105.115 ;
        RECT 155.645 104.985 157.015 105.795 ;
      LAYER nwell ;
        RECT 22.510 101.765 157.210 104.595 ;
      LAYER pwell ;
        RECT 22.705 100.565 24.075 101.375 ;
        RECT 24.085 100.565 29.595 101.375 ;
        RECT 30.655 101.245 31.585 101.475 ;
        RECT 34.645 101.245 35.575 101.475 ;
        RECT 29.750 100.565 31.585 101.245 ;
        RECT 32.825 100.565 35.575 101.245 ;
        RECT 35.595 100.650 36.025 101.435 ;
        RECT 36.045 100.565 37.415 101.345 ;
        RECT 37.425 100.565 39.255 101.375 ;
        RECT 39.725 100.565 41.075 101.475 ;
        RECT 41.415 101.245 42.345 101.475 ;
        RECT 41.415 100.565 43.250 101.245 ;
        RECT 44.325 100.565 45.695 101.345 ;
        RECT 45.705 100.565 49.375 101.375 ;
        RECT 49.425 101.245 50.775 101.475 ;
        RECT 52.310 101.245 53.220 101.465 ;
        RECT 49.425 100.565 56.735 101.245 ;
        RECT 56.745 100.565 58.115 101.375 ;
        RECT 58.125 100.565 61.335 101.475 ;
        RECT 61.355 100.650 61.785 101.435 ;
        RECT 61.805 100.565 63.635 101.375 ;
        RECT 63.695 100.565 68.165 101.475 ;
        RECT 68.265 100.565 69.615 101.475 ;
        RECT 69.625 100.565 75.135 101.375 ;
        RECT 75.145 100.565 76.515 101.375 ;
        RECT 76.535 100.565 79.265 101.475 ;
        RECT 79.745 100.565 82.955 101.475 ;
        RECT 82.965 100.565 86.635 101.475 ;
        RECT 87.115 100.650 87.545 101.435 ;
        RECT 91.080 101.245 91.990 101.465 ;
        RECT 93.525 101.245 94.875 101.475 ;
        RECT 87.565 100.565 94.875 101.245 ;
        RECT 94.925 101.245 95.845 101.475 ;
        RECT 94.925 100.565 97.215 101.245 ;
        RECT 97.225 100.565 100.895 101.475 ;
        RECT 100.925 100.565 102.275 101.475 ;
        RECT 102.285 100.565 103.635 101.475 ;
        RECT 103.665 100.565 109.175 101.375 ;
        RECT 109.185 100.565 112.855 101.375 ;
        RECT 112.875 100.650 113.305 101.435 ;
        RECT 113.325 100.565 114.675 101.475 ;
        RECT 115.665 101.245 117.015 101.475 ;
        RECT 118.550 101.245 119.460 101.465 ;
        RECT 115.665 100.565 122.975 101.245 ;
        RECT 122.985 100.565 124.815 101.375 ;
        RECT 128.340 101.245 129.250 101.465 ;
        RECT 130.785 101.245 132.135 101.475 ;
        RECT 124.825 100.565 132.135 101.245 ;
        RECT 132.280 101.245 133.200 101.475 ;
        RECT 135.865 101.275 136.810 101.475 ;
        RECT 132.280 100.565 135.745 101.245 ;
        RECT 135.865 100.595 138.615 101.275 ;
        RECT 138.635 100.650 139.065 101.435 ;
        RECT 135.865 100.565 136.810 100.595 ;
        RECT 22.845 100.355 23.015 100.565 ;
        RECT 24.225 100.355 24.395 100.565 ;
        RECT 29.750 100.545 29.915 100.565 ;
        RECT 29.745 100.375 29.915 100.545 ;
        RECT 31.595 100.400 31.755 100.510 ;
        RECT 32.055 100.410 32.215 100.520 ;
        RECT 32.965 100.375 33.135 100.565 ;
        RECT 34.345 100.355 34.515 100.545 ;
        RECT 34.805 100.375 34.975 100.545 ;
        RECT 37.105 100.375 37.275 100.565 ;
        RECT 37.565 100.375 37.735 100.565 ;
        RECT 34.825 100.355 34.975 100.375 ;
        RECT 38.030 100.355 38.200 100.545 ;
        RECT 38.485 100.355 38.655 100.545 ;
        RECT 39.400 100.405 39.520 100.515 ;
        RECT 40.790 100.375 40.960 100.565 ;
        RECT 43.085 100.545 43.250 100.565 ;
        RECT 43.085 100.375 43.255 100.545 ;
        RECT 43.555 100.410 43.715 100.520 ;
        RECT 44.005 100.355 44.175 100.545 ;
        RECT 45.385 100.375 45.555 100.565 ;
        RECT 45.845 100.375 46.015 100.565 ;
        RECT 47.695 100.400 47.855 100.510 ;
        RECT 49.065 100.355 49.235 100.545 ;
        RECT 54.595 100.400 54.755 100.510 ;
        RECT 55.505 100.355 55.675 100.545 ;
        RECT 56.425 100.375 56.595 100.565 ;
        RECT 56.885 100.375 57.055 100.565 ;
        RECT 58.255 100.375 58.425 100.565 ;
        RECT 58.725 100.355 58.895 100.545 ;
        RECT 61.945 100.375 62.115 100.565 ;
        RECT 62.410 100.355 62.580 100.545 ;
        RECT 63.765 100.375 63.935 100.565 ;
        RECT 66.085 100.355 66.255 100.545 ;
        RECT 69.300 100.375 69.470 100.565 ;
        RECT 69.765 100.355 69.935 100.565 ;
        RECT 72.070 100.355 72.240 100.545 ;
        RECT 72.525 100.355 72.695 100.545 ;
        RECT 74.825 100.355 74.995 100.545 ;
        RECT 75.285 100.375 75.455 100.565 ;
        RECT 76.665 100.375 76.835 100.565 ;
        RECT 79.420 100.405 79.540 100.515 ;
        RECT 79.875 100.375 80.045 100.565 ;
        RECT 82.190 100.355 82.360 100.545 ;
        RECT 83.110 100.375 83.280 100.565 ;
        RECT 85.865 100.355 86.035 100.545 ;
        RECT 86.780 100.405 86.900 100.515 ;
        RECT 87.705 100.375 87.875 100.565 ;
        RECT 89.545 100.355 89.715 100.545 ;
        RECT 92.305 100.355 92.475 100.545 ;
        RECT 95.980 100.405 96.100 100.515 ;
        RECT 96.450 100.355 96.620 100.545 ;
        RECT 96.905 100.375 97.075 100.565 ;
        RECT 97.370 100.375 97.540 100.565 ;
        RECT 100.585 100.355 100.755 100.545 ;
        RECT 101.960 100.375 102.130 100.565 ;
        RECT 102.430 100.375 102.600 100.565 ;
        RECT 103.805 100.375 103.975 100.565 ;
        RECT 104.275 100.400 104.435 100.510 ;
        RECT 105.185 100.355 105.355 100.545 ;
        RECT 109.325 100.375 109.495 100.565 ;
        RECT 112.540 100.405 112.660 100.515 ;
        RECT 114.390 100.375 114.560 100.565 ;
        RECT 114.855 100.410 115.015 100.520 ;
        RECT 116.225 100.355 116.395 100.545 ;
        RECT 116.685 100.355 116.855 100.545 ;
        RECT 119.905 100.355 120.075 100.545 ;
        RECT 122.665 100.375 122.835 100.565 ;
        RECT 123.125 100.375 123.295 100.565 ;
        RECT 124.965 100.375 125.135 100.565 ;
        RECT 125.420 100.405 125.540 100.515 ;
        RECT 124.965 100.355 125.115 100.375 ;
        RECT 126.345 100.355 126.515 100.545 ;
        RECT 128.180 100.405 128.300 100.515 ;
        RECT 128.645 100.355 128.815 100.545 ;
        RECT 130.485 100.355 130.655 100.545 ;
        RECT 135.545 100.375 135.715 100.565 ;
        RECT 138.300 100.375 138.470 100.595 ;
        RECT 139.085 100.565 143.900 101.245 ;
        RECT 144.340 100.565 147.815 101.475 ;
        RECT 151.800 101.245 152.710 101.465 ;
        RECT 154.245 101.245 155.595 101.475 ;
        RECT 148.285 100.565 155.595 101.245 ;
        RECT 155.645 100.565 157.015 101.375 ;
        RECT 139.225 100.375 139.395 100.565 ;
        RECT 140.145 100.355 140.315 100.545 ;
        RECT 143.820 100.355 143.990 100.545 ;
        RECT 144.285 100.355 144.455 100.545 ;
        RECT 147.500 100.375 147.670 100.565 ;
        RECT 147.970 100.515 148.140 100.545 ;
        RECT 147.960 100.405 148.140 100.515 ;
        RECT 147.970 100.355 148.140 100.405 ;
        RECT 148.425 100.375 148.595 100.565 ;
        RECT 155.325 100.355 155.495 100.545 ;
        RECT 156.705 100.355 156.875 100.565 ;
        RECT 22.705 99.545 24.075 100.355 ;
        RECT 24.085 99.675 31.395 100.355 ;
        RECT 27.600 99.455 28.510 99.675 ;
        RECT 30.045 99.445 31.395 99.675 ;
        RECT 32.365 99.675 34.655 100.355 ;
        RECT 32.365 99.445 33.285 99.675 ;
        RECT 34.825 99.535 36.755 100.355 ;
        RECT 35.805 99.445 36.755 99.535 ;
        RECT 36.965 99.445 38.315 100.355 ;
        RECT 38.345 99.545 43.855 100.355 ;
        RECT 43.865 99.545 47.535 100.355 ;
        RECT 48.475 99.485 48.905 100.270 ;
        RECT 48.925 99.545 54.435 100.355 ;
        RECT 55.465 99.445 58.575 100.355 ;
        RECT 58.585 99.545 62.255 100.355 ;
        RECT 62.265 99.445 65.935 100.355 ;
        RECT 65.945 99.545 69.615 100.355 ;
        RECT 69.625 99.545 70.995 100.355 ;
        RECT 71.005 99.445 72.355 100.355 ;
        RECT 72.385 99.545 74.215 100.355 ;
        RECT 74.235 99.485 74.665 100.270 ;
        RECT 74.685 99.675 81.995 100.355 ;
        RECT 78.200 99.455 79.110 99.675 ;
        RECT 80.645 99.445 81.995 99.675 ;
        RECT 82.045 99.445 85.715 100.355 ;
        RECT 85.725 99.545 89.395 100.355 ;
        RECT 89.415 99.445 92.145 100.355 ;
        RECT 92.165 99.545 95.835 100.355 ;
        RECT 96.305 99.445 99.975 100.355 ;
        RECT 99.995 99.485 100.425 100.270 ;
        RECT 100.445 99.545 104.115 100.355 ;
        RECT 105.045 99.675 112.355 100.355 ;
        RECT 108.560 99.455 109.470 99.675 ;
        RECT 111.005 99.445 112.355 99.675 ;
        RECT 112.960 99.675 116.425 100.355 ;
        RECT 112.960 99.445 113.880 99.675 ;
        RECT 116.545 99.445 119.755 100.355 ;
        RECT 119.845 99.445 122.845 100.355 ;
        RECT 123.185 99.535 125.115 100.355 ;
        RECT 123.185 99.445 124.135 99.535 ;
        RECT 125.755 99.485 126.185 100.270 ;
        RECT 126.205 99.545 128.035 100.355 ;
        RECT 128.505 99.675 130.335 100.355 ;
        RECT 128.990 99.445 130.335 99.675 ;
        RECT 130.345 99.545 133.095 100.355 ;
        RECT 133.145 99.675 140.455 100.355 ;
        RECT 133.145 99.445 134.495 99.675 ;
        RECT 136.030 99.455 136.940 99.675 ;
        RECT 140.660 99.445 144.135 100.355 ;
        RECT 144.255 99.675 147.720 100.355 ;
        RECT 146.800 99.445 147.720 99.675 ;
        RECT 147.825 99.445 151.300 100.355 ;
        RECT 151.515 99.485 151.945 100.270 ;
        RECT 152.060 99.675 155.525 100.355 ;
        RECT 152.060 99.445 152.980 99.675 ;
        RECT 155.645 99.545 157.015 100.355 ;
      LAYER nwell ;
        RECT 22.510 96.325 157.210 99.155 ;
      LAYER pwell ;
        RECT 22.705 95.125 24.075 95.935 ;
        RECT 24.085 95.125 25.455 95.935 ;
        RECT 25.465 95.125 26.835 95.905 ;
        RECT 26.845 95.125 29.595 95.935 ;
        RECT 29.605 95.355 32.355 96.035 ;
        RECT 32.365 95.835 33.310 96.035 ;
        RECT 34.645 95.835 35.575 96.035 ;
        RECT 32.365 95.355 35.575 95.835 ;
        RECT 29.605 95.125 32.215 95.355 ;
        RECT 32.365 95.155 35.435 95.355 ;
        RECT 35.595 95.210 36.025 95.995 ;
        RECT 40.480 95.805 41.390 96.025 ;
        RECT 42.925 95.805 44.275 96.035 ;
        RECT 47.840 95.805 48.750 96.025 ;
        RECT 50.285 95.805 51.635 96.035 ;
        RECT 32.365 95.125 33.310 95.155 ;
        RECT 22.845 94.915 23.015 95.125 ;
        RECT 24.225 94.915 24.395 95.125 ;
        RECT 26.525 94.935 26.695 95.125 ;
        RECT 26.985 94.935 27.155 95.125 ;
        RECT 29.745 94.915 29.915 95.105 ;
        RECT 32.045 94.935 32.215 95.125 ;
        RECT 32.510 94.915 32.680 95.105 ;
        RECT 33.885 94.915 34.055 95.105 ;
        RECT 35.265 94.935 35.435 95.155 ;
        RECT 36.965 95.125 44.275 95.805 ;
        RECT 44.325 95.125 51.635 95.805 ;
        RECT 51.685 95.125 55.355 95.935 ;
        RECT 55.365 95.125 56.735 95.905 ;
        RECT 56.745 95.125 60.415 95.935 ;
        RECT 61.355 95.210 61.785 95.995 ;
        RECT 61.805 95.125 65.475 95.935 ;
        RECT 65.485 95.125 68.695 96.035 ;
        RECT 71.360 95.805 72.280 96.035 ;
        RECT 78.365 95.805 79.285 96.035 ;
        RECT 80.760 95.805 81.680 96.035 ;
        RECT 68.815 95.125 72.280 95.805 ;
        RECT 72.385 95.125 77.200 95.805 ;
        RECT 78.365 95.125 80.655 95.805 ;
        RECT 80.760 95.125 84.225 95.805 ;
        RECT 84.345 95.125 85.695 96.035 ;
        RECT 85.725 95.125 87.095 95.935 ;
        RECT 87.115 95.210 87.545 95.995 ;
        RECT 87.565 95.125 89.395 95.935 ;
        RECT 91.235 95.805 92.155 96.035 ;
        RECT 89.865 95.125 92.155 95.805 ;
        RECT 92.165 95.125 93.995 95.935 ;
        RECT 95.515 95.805 96.445 96.035 ;
        RECT 94.610 95.125 96.445 95.805 ;
        RECT 96.765 95.125 98.115 96.035 ;
        RECT 98.145 95.125 100.895 95.935 ;
        RECT 101.365 95.125 102.735 95.905 ;
        RECT 102.745 95.125 106.415 95.935 ;
        RECT 107.345 95.125 108.715 95.905 ;
        RECT 109.185 95.805 110.115 96.035 ;
        RECT 109.185 95.125 111.935 95.805 ;
        RECT 112.875 95.210 113.305 95.995 ;
        RECT 113.325 95.125 114.675 96.035 ;
        RECT 116.675 95.805 117.605 96.035 ;
        RECT 115.770 95.125 117.605 95.805 ;
        RECT 117.925 95.125 119.275 96.035 ;
        RECT 121.275 95.805 122.205 96.035 ;
        RECT 120.370 95.125 122.205 95.805 ;
        RECT 122.540 95.125 124.355 96.035 ;
        RECT 124.365 95.125 126.195 95.935 ;
        RECT 126.215 95.125 127.565 96.035 ;
        RECT 127.605 95.125 128.955 96.035 ;
        RECT 128.965 95.125 134.475 95.935 ;
        RECT 134.485 95.125 135.855 95.935 ;
        RECT 136.175 95.805 137.105 96.035 ;
        RECT 136.175 95.125 138.010 95.805 ;
        RECT 138.635 95.210 139.065 95.995 ;
        RECT 139.125 95.805 140.475 96.035 ;
        RECT 142.010 95.805 142.920 96.025 ;
        RECT 139.125 95.125 146.435 95.805 ;
        RECT 146.445 95.125 147.815 95.935 ;
        RECT 151.340 95.805 152.250 96.025 ;
        RECT 153.785 95.805 155.135 96.035 ;
        RECT 147.825 95.125 155.135 95.805 ;
        RECT 155.645 95.125 157.015 95.935 ;
        RECT 35.720 94.965 35.840 95.075 ;
        RECT 36.195 94.970 36.355 95.080 ;
        RECT 37.105 94.935 37.275 95.125 ;
        RECT 40.785 94.915 40.955 95.105 ;
        RECT 42.165 94.915 42.335 95.105 ;
        RECT 42.625 94.915 42.795 95.105 ;
        RECT 44.465 94.935 44.635 95.125 ;
        RECT 48.140 94.965 48.260 95.075 ;
        RECT 49.985 94.915 50.155 95.105 ;
        RECT 50.455 94.960 50.615 95.070 ;
        RECT 22.705 94.105 24.075 94.915 ;
        RECT 24.085 94.105 29.595 94.915 ;
        RECT 29.605 94.105 32.355 94.915 ;
        RECT 32.365 94.005 33.715 94.915 ;
        RECT 33.745 94.105 35.575 94.915 ;
        RECT 36.280 94.235 41.095 94.915 ;
        RECT 41.105 94.135 42.475 94.915 ;
        RECT 42.485 94.105 47.995 94.915 ;
        RECT 48.475 94.045 48.905 94.830 ;
        RECT 48.925 94.135 50.295 94.915 ;
        RECT 51.370 94.885 51.540 95.105 ;
        RECT 51.825 94.935 51.995 95.125 ;
        RECT 54.585 94.915 54.755 95.105 ;
        RECT 55.505 94.935 55.675 95.125 ;
        RECT 56.885 94.935 57.055 95.125 ;
        RECT 60.575 94.970 60.735 95.080 ;
        RECT 61.945 94.915 62.115 95.125 ;
        RECT 65.625 94.915 65.795 95.105 ;
        RECT 66.085 94.915 66.255 95.105 ;
        RECT 68.385 94.935 68.555 95.125 ;
        RECT 68.845 94.935 69.015 95.125 ;
        RECT 72.525 94.935 72.695 95.125 ;
        RECT 73.455 94.960 73.615 95.070 ;
        RECT 74.825 94.935 74.995 95.105 ;
        RECT 74.830 94.915 74.995 94.935 ;
        RECT 77.125 94.915 77.295 95.105 ;
        RECT 77.595 94.970 77.755 95.080 ;
        RECT 80.345 94.935 80.515 95.125 ;
        RECT 81.725 94.935 81.895 95.105 ;
        RECT 81.725 94.915 81.875 94.935 ;
        RECT 82.185 94.915 82.355 95.105 ;
        RECT 84.025 94.935 84.195 95.125 ;
        RECT 84.490 94.935 84.660 95.125 ;
        RECT 85.865 94.935 86.035 95.125 ;
        RECT 87.705 95.105 87.875 95.125 ;
        RECT 87.700 94.935 87.875 95.105 ;
        RECT 87.700 94.915 87.870 94.935 ;
        RECT 88.165 94.915 88.335 95.105 ;
        RECT 89.540 94.965 89.660 95.075 ;
        RECT 90.005 94.935 90.175 95.125 ;
        RECT 92.305 94.935 92.475 95.125 ;
        RECT 94.610 95.105 94.775 95.125 ;
        RECT 94.140 94.965 94.260 95.075 ;
        RECT 94.605 94.935 94.775 95.105 ;
        RECT 95.525 94.915 95.695 95.105 ;
        RECT 97.830 94.935 98.000 95.125 ;
        RECT 98.285 94.935 98.455 95.125 ;
        RECT 100.585 94.915 100.755 95.105 ;
        RECT 101.040 94.965 101.160 95.075 ;
        RECT 102.425 94.935 102.595 95.125 ;
        RECT 102.885 94.935 103.055 95.125 ;
        RECT 106.575 94.970 106.735 95.080 ;
        RECT 108.405 94.935 108.575 95.125 ;
        RECT 108.860 94.965 108.980 95.075 ;
        RECT 111.625 94.935 111.795 95.125 ;
        RECT 112.095 94.970 112.255 95.080 ;
        RECT 112.545 94.915 112.715 95.105 ;
        RECT 113.010 94.915 113.180 95.105 ;
        RECT 114.390 94.935 114.560 95.125 ;
        RECT 115.770 95.105 115.935 95.125 ;
        RECT 114.855 94.970 115.015 95.080 ;
        RECT 115.765 94.935 115.935 95.105 ;
        RECT 116.220 94.965 116.340 95.075 ;
        RECT 116.675 94.915 116.845 95.105 ;
        RECT 118.070 94.935 118.240 95.125 ;
        RECT 120.370 95.105 120.535 95.125 ;
        RECT 119.455 94.970 119.615 95.080 ;
        RECT 119.915 94.960 120.075 95.070 ;
        RECT 120.365 94.935 120.535 95.105 ;
        RECT 120.825 94.915 120.995 95.105 ;
        RECT 122.665 94.935 122.835 95.125 ;
        RECT 124.505 95.105 124.675 95.125 ;
        RECT 124.505 94.935 124.680 95.105 ;
        RECT 124.510 94.915 124.680 94.935 ;
        RECT 126.345 94.915 126.515 95.105 ;
        RECT 127.265 94.935 127.435 95.125 ;
        RECT 128.640 94.935 128.810 95.125 ;
        RECT 129.105 94.935 129.275 95.125 ;
        RECT 133.705 94.935 133.875 95.105 ;
        RECT 134.625 94.935 134.795 95.125 ;
        RECT 137.845 95.105 138.010 95.125 ;
        RECT 136.000 94.965 136.120 95.075 ;
        RECT 137.845 94.935 138.015 95.105 ;
        RECT 138.305 95.075 138.475 95.105 ;
        RECT 138.300 94.965 138.475 95.075 ;
        RECT 138.305 94.935 138.475 94.965 ;
        RECT 133.710 94.915 133.875 94.935 ;
        RECT 138.305 94.915 138.470 94.935 ;
        RECT 139.690 94.915 139.860 95.105 ;
        RECT 141.070 94.915 141.240 95.105 ;
        RECT 141.520 94.965 141.640 95.075 ;
        RECT 141.985 94.935 142.155 95.105 ;
        RECT 146.125 94.935 146.295 95.125 ;
        RECT 146.585 94.935 146.755 95.125 ;
        RECT 147.965 95.105 148.135 95.125 ;
        RECT 141.990 94.915 142.155 94.935 ;
        RECT 147.505 94.915 147.675 95.105 ;
        RECT 147.965 94.935 148.140 95.105 ;
        RECT 155.325 95.075 155.495 95.105 ;
        RECT 155.320 94.965 155.495 95.075 ;
        RECT 147.970 94.915 148.140 94.935 ;
        RECT 155.325 94.915 155.495 94.965 ;
        RECT 156.705 94.915 156.875 95.125 ;
        RECT 53.500 94.885 54.435 94.915 ;
        RECT 51.370 94.685 54.435 94.885 ;
        RECT 51.225 94.205 54.435 94.685 ;
        RECT 54.445 94.235 61.755 94.915 ;
        RECT 51.225 94.005 52.155 94.205 ;
        RECT 53.485 94.005 54.435 94.205 ;
        RECT 57.960 94.015 58.870 94.235 ;
        RECT 60.405 94.005 61.755 94.235 ;
        RECT 61.805 94.135 63.175 94.915 ;
        RECT 63.185 94.235 65.935 94.915 ;
        RECT 65.945 94.235 73.255 94.915 ;
        RECT 63.185 94.005 64.115 94.235 ;
        RECT 69.460 94.015 70.370 94.235 ;
        RECT 71.905 94.005 73.255 94.235 ;
        RECT 74.235 94.045 74.665 94.830 ;
        RECT 74.830 94.235 76.665 94.915 ;
        RECT 75.735 94.005 76.665 94.235 ;
        RECT 76.985 94.105 79.735 94.915 ;
        RECT 79.945 94.095 81.875 94.915 ;
        RECT 79.945 94.005 80.895 94.095 ;
        RECT 82.055 94.005 84.785 94.915 ;
        RECT 85.095 94.005 88.015 94.915 ;
        RECT 88.025 94.235 95.335 94.915 ;
        RECT 91.540 94.015 92.450 94.235 ;
        RECT 93.985 94.005 95.335 94.235 ;
        RECT 95.385 94.005 99.935 94.915 ;
        RECT 99.995 94.045 100.425 94.830 ;
        RECT 100.445 94.235 107.755 94.915 ;
        RECT 108.040 94.235 112.855 94.915 ;
        RECT 103.960 94.015 104.870 94.235 ;
        RECT 106.405 94.005 107.755 94.235 ;
        RECT 112.865 94.005 115.785 94.915 ;
        RECT 116.545 94.005 119.755 94.915 ;
        RECT 120.765 94.005 124.215 94.915 ;
        RECT 124.365 94.005 125.715 94.915 ;
        RECT 125.755 94.045 126.185 94.830 ;
        RECT 126.205 94.235 133.515 94.915 ;
        RECT 133.710 94.235 135.545 94.915 ;
        RECT 129.720 94.015 130.630 94.235 ;
        RECT 132.165 94.005 133.515 94.235 ;
        RECT 134.615 94.005 135.545 94.235 ;
        RECT 136.635 94.235 138.470 94.915 ;
        RECT 136.635 94.005 137.565 94.235 ;
        RECT 138.625 94.005 139.975 94.915 ;
        RECT 140.005 94.005 141.355 94.915 ;
        RECT 141.990 94.235 143.825 94.915 ;
        RECT 142.895 94.005 143.825 94.235 ;
        RECT 144.240 94.235 147.705 94.915 ;
        RECT 144.240 94.005 145.160 94.235 ;
        RECT 147.825 94.005 151.300 94.915 ;
        RECT 151.515 94.045 151.945 94.830 ;
        RECT 152.060 94.235 155.525 94.915 ;
        RECT 152.060 94.005 152.980 94.235 ;
        RECT 155.645 94.105 157.015 94.915 ;
      LAYER nwell ;
        RECT 22.510 90.885 157.210 93.715 ;
      LAYER pwell ;
        RECT 22.705 89.685 24.075 90.495 ;
        RECT 27.600 90.365 28.510 90.585 ;
        RECT 30.045 90.365 31.395 90.595 ;
        RECT 34.170 90.395 35.115 90.595 ;
        RECT 24.085 89.685 31.395 90.365 ;
        RECT 32.365 89.715 35.115 90.395 ;
        RECT 35.595 89.770 36.025 90.555 ;
        RECT 22.845 89.475 23.015 89.685 ;
        RECT 24.225 89.475 24.395 89.685 ;
        RECT 29.740 89.525 29.860 89.635 ;
        RECT 31.120 89.475 31.290 89.665 ;
        RECT 31.580 89.640 31.750 89.665 ;
        RECT 31.580 89.530 31.755 89.640 ;
        RECT 31.580 89.475 31.750 89.530 ;
        RECT 32.510 89.495 32.680 89.715 ;
        RECT 34.170 89.685 35.115 89.715 ;
        RECT 36.045 89.685 38.965 90.595 ;
        RECT 41.555 90.365 42.475 90.595 ;
        RECT 40.185 89.685 42.475 90.365 ;
        RECT 42.485 89.685 45.695 90.595 ;
        RECT 46.175 89.685 47.525 90.595 ;
        RECT 47.545 90.395 48.475 90.595 ;
        RECT 49.805 90.395 50.755 90.595 ;
        RECT 47.545 89.915 50.755 90.395 ;
        RECT 47.690 89.715 50.755 89.915 ;
        RECT 32.970 89.475 33.140 89.665 ;
        RECT 35.260 89.525 35.380 89.635 ;
        RECT 36.190 89.495 36.360 89.685 ;
        RECT 36.645 89.475 36.815 89.665 ;
        RECT 38.485 89.475 38.655 89.665 ;
        RECT 39.415 89.530 39.575 89.640 ;
        RECT 40.325 89.495 40.495 89.685 ;
        RECT 42.165 89.495 42.335 89.665 ;
        RECT 42.615 89.495 42.785 89.685 ;
        RECT 42.165 89.475 42.315 89.495 ;
        RECT 44.925 89.475 45.095 89.665 ;
        RECT 45.385 89.495 45.555 89.665 ;
        RECT 45.840 89.525 45.960 89.635 ;
        RECT 47.225 89.495 47.395 89.685 ;
        RECT 47.690 89.495 47.860 89.715 ;
        RECT 49.820 89.685 50.755 89.715 ;
        RECT 50.765 89.685 54.240 90.595 ;
        RECT 54.915 89.685 56.265 90.595 ;
        RECT 56.285 90.365 59.110 90.595 ;
        RECT 56.285 89.685 59.815 90.365 ;
        RECT 59.965 89.685 61.315 90.595 ;
        RECT 61.355 89.770 61.785 90.555 ;
        RECT 62.855 90.365 63.785 90.595 ;
        RECT 61.950 89.685 63.785 90.365 ;
        RECT 64.105 89.685 65.935 90.495 ;
        RECT 66.405 89.685 69.325 90.595 ;
        RECT 69.635 89.685 72.365 90.595 ;
        RECT 72.385 89.685 73.735 90.595 ;
        RECT 73.765 89.685 77.435 90.495 ;
        RECT 77.985 89.685 81.435 90.595 ;
        RECT 81.585 89.685 84.505 90.595 ;
        RECT 84.805 89.685 86.635 90.495 ;
        RECT 87.115 89.770 87.545 90.555 ;
        RECT 87.565 90.365 88.495 90.595 ;
        RECT 87.565 89.685 90.315 90.365 ;
        RECT 90.325 89.685 91.695 90.465 ;
        RECT 91.705 89.685 93.535 90.495 ;
        RECT 94.005 89.685 97.215 90.595 ;
        RECT 97.695 89.685 99.045 90.595 ;
        RECT 99.065 90.395 99.995 90.595 ;
        RECT 101.325 90.395 102.275 90.595 ;
        RECT 99.065 89.915 102.275 90.395 ;
        RECT 99.210 89.715 102.275 89.915 ;
        RECT 49.075 89.520 49.235 89.630 ;
        RECT 45.390 89.475 45.555 89.495 ;
        RECT 49.975 89.475 50.145 89.665 ;
        RECT 50.910 89.495 51.080 89.685 ;
        RECT 53.205 89.495 53.375 89.665 ;
        RECT 54.580 89.525 54.700 89.635 ;
        RECT 53.210 89.475 53.375 89.495 ;
        RECT 55.505 89.475 55.675 89.665 ;
        RECT 55.965 89.495 56.135 89.685 ;
        RECT 59.615 89.665 59.815 89.685 ;
        RECT 59.645 89.495 59.815 89.665 ;
        RECT 22.705 88.665 24.075 89.475 ;
        RECT 24.085 88.665 29.595 89.475 ;
        RECT 30.085 88.565 31.435 89.475 ;
        RECT 31.465 88.565 32.815 89.475 ;
        RECT 32.825 88.565 36.300 89.475 ;
        RECT 36.520 88.565 38.335 89.475 ;
        RECT 38.345 88.665 40.175 89.475 ;
        RECT 40.385 88.655 42.315 89.475 ;
        RECT 40.385 88.565 41.335 88.655 ;
        RECT 42.515 88.565 45.235 89.475 ;
        RECT 45.390 88.795 47.225 89.475 ;
        RECT 46.295 88.565 47.225 88.795 ;
        RECT 48.475 88.605 48.905 89.390 ;
        RECT 49.845 88.565 53.055 89.475 ;
        RECT 53.210 88.795 55.045 89.475 ;
        RECT 54.115 88.565 55.045 88.795 ;
        RECT 55.365 88.665 57.195 89.475 ;
        RECT 57.205 89.445 58.140 89.475 ;
        RECT 60.100 89.445 60.270 89.665 ;
        RECT 60.565 89.475 60.735 89.665 ;
        RECT 61.030 89.495 61.200 89.685 ;
        RECT 61.950 89.665 62.115 89.685 ;
        RECT 61.945 89.495 62.115 89.665 ;
        RECT 64.245 89.495 64.415 89.685 ;
        RECT 66.085 89.635 66.255 89.665 ;
        RECT 66.080 89.525 66.255 89.635 ;
        RECT 66.085 89.475 66.255 89.525 ;
        RECT 66.550 89.495 66.720 89.685 ;
        RECT 69.765 89.495 69.935 89.685 ;
        RECT 71.605 89.475 71.775 89.665 ;
        RECT 73.450 89.495 73.620 89.685 ;
        RECT 73.905 89.495 74.075 89.685 ;
        RECT 74.825 89.475 74.995 89.665 ;
        RECT 77.580 89.525 77.700 89.635 ;
        RECT 78.045 89.495 78.215 89.685 ;
        RECT 81.730 89.495 81.900 89.685 ;
        RECT 82.185 89.495 82.355 89.665 ;
        RECT 84.495 89.520 84.655 89.630 ;
        RECT 84.945 89.495 85.115 89.685 ;
        RECT 82.190 89.475 82.355 89.495 ;
        RECT 85.405 89.475 85.575 89.665 ;
        RECT 86.780 89.630 86.900 89.635 ;
        RECT 86.780 89.525 86.955 89.630 ;
        RECT 86.795 89.520 86.955 89.525 ;
        RECT 87.700 89.475 87.870 89.665 ;
        RECT 89.085 89.475 89.255 89.665 ;
        RECT 90.005 89.495 90.175 89.685 ;
        RECT 91.385 89.495 91.555 89.685 ;
        RECT 91.845 89.495 92.015 89.685 ;
        RECT 93.680 89.525 93.800 89.635 ;
        RECT 94.135 89.495 94.305 89.685 ;
        RECT 94.605 89.475 94.775 89.665 ;
        RECT 97.360 89.525 97.480 89.635 ;
        RECT 98.745 89.495 98.915 89.685 ;
        RECT 99.210 89.495 99.380 89.715 ;
        RECT 101.340 89.685 102.275 89.715 ;
        RECT 103.205 89.685 106.680 90.595 ;
        RECT 106.885 89.685 108.255 90.495 ;
        RECT 108.275 89.685 111.005 90.595 ;
        RECT 111.025 89.685 112.375 90.595 ;
        RECT 112.875 89.770 113.305 90.555 ;
        RECT 113.325 90.365 114.245 90.595 ;
        RECT 113.325 89.685 115.615 90.365 ;
        RECT 115.625 89.685 116.995 90.495 ;
        RECT 117.005 89.685 121.555 90.595 ;
        RECT 121.605 89.685 125.275 90.495 ;
        RECT 125.285 89.685 126.655 90.495 ;
        RECT 126.665 89.685 128.480 90.595 ;
        RECT 128.505 89.685 131.425 90.595 ;
        RECT 131.725 89.685 134.475 90.495 ;
        RECT 134.945 89.685 138.155 90.595 ;
        RECT 138.635 89.770 139.065 90.555 ;
        RECT 139.085 89.685 141.835 90.495 ;
        RECT 141.845 89.685 143.215 90.465 ;
        RECT 146.740 90.365 147.650 90.585 ;
        RECT 149.185 90.365 150.535 90.595 ;
        RECT 143.225 89.685 150.535 90.365 ;
        RECT 151.600 90.365 152.520 90.595 ;
        RECT 151.600 89.685 155.065 90.365 ;
        RECT 155.645 89.685 157.015 90.495 ;
        RECT 100.585 89.475 100.755 89.665 ;
        RECT 102.415 89.640 102.585 89.665 ;
        RECT 102.415 89.530 102.595 89.640 ;
        RECT 102.415 89.475 102.585 89.530 ;
        RECT 103.350 89.495 103.520 89.685 ;
        RECT 106.565 89.475 106.735 89.665 ;
        RECT 107.025 89.495 107.195 89.685 ;
        RECT 108.405 89.495 108.575 89.685 ;
        RECT 108.865 89.495 109.035 89.665 ;
        RECT 108.865 89.475 109.030 89.495 ;
        RECT 109.325 89.475 109.495 89.665 ;
        RECT 110.705 89.475 110.875 89.665 ;
        RECT 112.090 89.495 112.260 89.685 ;
        RECT 112.540 89.525 112.660 89.635 ;
        RECT 115.305 89.495 115.475 89.685 ;
        RECT 115.765 89.495 115.935 89.685 ;
        RECT 117.145 89.495 117.315 89.685 ;
        RECT 119.905 89.495 120.075 89.665 ;
        RECT 119.905 89.475 120.070 89.495 ;
        RECT 120.360 89.475 120.530 89.665 ;
        RECT 121.745 89.475 121.915 89.685 ;
        RECT 125.425 89.635 125.595 89.685 ;
        RECT 125.420 89.525 125.595 89.635 ;
        RECT 126.340 89.525 126.460 89.635 ;
        RECT 125.425 89.495 125.595 89.525 ;
        RECT 126.805 89.475 126.975 89.665 ;
        RECT 128.185 89.495 128.355 89.685 ;
        RECT 128.650 89.495 128.820 89.685 ;
        RECT 129.105 89.475 129.275 89.665 ;
        RECT 131.865 89.495 132.035 89.685 ;
        RECT 135.075 89.665 135.245 89.685 ;
        RECT 134.620 89.525 134.740 89.635 ;
        RECT 135.075 89.495 135.255 89.665 ;
        RECT 138.300 89.525 138.420 89.635 ;
        RECT 139.225 89.495 139.395 89.685 ;
        RECT 141.985 89.665 142.155 89.685 ;
        RECT 139.680 89.525 139.800 89.635 ;
        RECT 135.085 89.475 135.255 89.495 ;
        RECT 141.065 89.475 141.235 89.665 ;
        RECT 141.520 89.525 141.640 89.635 ;
        RECT 141.985 89.495 142.160 89.665 ;
        RECT 143.365 89.495 143.535 89.685 ;
        RECT 141.990 89.475 142.160 89.495 ;
        RECT 148.435 89.475 148.605 89.665 ;
        RECT 148.885 89.495 149.055 89.665 ;
        RECT 150.735 89.530 150.895 89.640 ;
        RECT 151.180 89.525 151.300 89.635 ;
        RECT 152.105 89.495 152.275 89.665 ;
        RECT 148.890 89.475 149.055 89.495 ;
        RECT 152.110 89.475 152.275 89.495 ;
        RECT 154.405 89.475 154.575 89.665 ;
        RECT 154.865 89.495 155.035 89.685 ;
        RECT 155.320 89.525 155.440 89.635 ;
        RECT 156.705 89.475 156.875 89.685 ;
        RECT 57.205 89.245 60.270 89.445 ;
        RECT 57.205 88.765 60.415 89.245 ;
        RECT 57.205 88.565 58.155 88.765 ;
        RECT 59.485 88.565 60.415 88.765 ;
        RECT 60.425 88.665 65.935 89.475 ;
        RECT 65.945 88.665 71.455 89.475 ;
        RECT 71.465 88.665 74.215 89.475 ;
        RECT 74.235 88.605 74.665 89.390 ;
        RECT 74.685 88.795 81.995 89.475 ;
        RECT 82.190 88.795 84.025 89.475 ;
        RECT 78.200 88.575 79.110 88.795 ;
        RECT 80.645 88.565 81.995 88.795 ;
        RECT 83.095 88.565 84.025 88.795 ;
        RECT 85.265 88.695 86.635 89.475 ;
        RECT 87.585 88.565 88.935 89.475 ;
        RECT 88.945 88.665 94.455 89.475 ;
        RECT 94.465 88.665 99.975 89.475 ;
        RECT 99.995 88.605 100.425 89.390 ;
        RECT 100.445 88.665 102.275 89.475 ;
        RECT 102.285 88.565 105.495 89.475 ;
        RECT 105.515 88.565 106.865 89.475 ;
        RECT 107.195 88.795 109.030 89.475 ;
        RECT 107.195 88.565 108.125 88.795 ;
        RECT 109.185 88.695 110.555 89.475 ;
        RECT 110.565 88.795 117.875 89.475 ;
        RECT 114.080 88.575 114.990 88.795 ;
        RECT 116.525 88.565 117.875 88.795 ;
        RECT 118.235 88.795 120.070 89.475 ;
        RECT 118.235 88.565 119.165 88.795 ;
        RECT 120.245 88.565 121.595 89.475 ;
        RECT 121.605 88.665 125.275 89.475 ;
        RECT 125.755 88.605 126.185 89.390 ;
        RECT 126.665 88.795 128.955 89.475 ;
        RECT 128.035 88.565 128.955 88.795 ;
        RECT 128.965 88.665 134.475 89.475 ;
        RECT 134.945 88.565 139.495 89.475 ;
        RECT 140.015 88.565 141.365 89.475 ;
        RECT 141.845 88.565 145.320 89.475 ;
        RECT 145.525 88.565 148.735 89.475 ;
        RECT 148.890 88.795 150.725 89.475 ;
        RECT 149.795 88.565 150.725 88.795 ;
        RECT 151.515 88.605 151.945 89.390 ;
        RECT 152.110 88.795 153.945 89.475 ;
        RECT 153.015 88.565 153.945 88.795 ;
        RECT 154.265 88.665 155.635 89.475 ;
        RECT 155.645 88.665 157.015 89.475 ;
      LAYER nwell ;
        RECT 22.510 85.445 157.210 88.275 ;
      LAYER pwell ;
        RECT 22.705 84.245 24.075 85.055 ;
        RECT 24.085 84.245 29.595 85.055 ;
        RECT 29.605 84.245 33.275 85.055 ;
        RECT 34.205 84.245 35.555 85.155 ;
        RECT 35.595 84.330 36.025 85.115 ;
        RECT 37.095 84.925 38.025 85.155 ;
        RECT 36.190 84.245 38.025 84.925 ;
        RECT 38.345 84.925 39.265 85.155 ;
        RECT 38.345 84.245 40.635 84.925 ;
        RECT 42.945 84.245 44.295 85.155 ;
        RECT 45.705 84.245 49.375 85.055 ;
        RECT 49.385 84.245 50.735 85.155 ;
        RECT 53.065 84.245 54.895 85.055 ;
        RECT 56.415 84.925 57.345 85.155 ;
        RECT 59.035 84.925 59.955 85.155 ;
        RECT 55.510 84.245 57.345 84.925 ;
        RECT 57.665 84.245 59.955 84.925 ;
        RECT 59.965 84.245 61.335 85.055 ;
        RECT 61.355 84.330 61.785 85.115 ;
        RECT 61.805 84.245 64.555 85.055 ;
        RECT 65.935 84.925 66.855 85.155 ;
        RECT 64.565 84.245 66.855 84.925 ;
        RECT 66.865 84.245 70.075 85.155 ;
        RECT 70.085 84.245 74.635 85.155 ;
        RECT 77.645 85.065 78.595 85.155 ;
        RECT 74.685 84.245 77.435 85.055 ;
        RECT 77.645 84.245 79.575 85.065 ;
        RECT 79.760 84.245 81.575 85.155 ;
        RECT 81.605 84.245 82.955 85.155 ;
        RECT 82.965 84.245 85.715 85.055 ;
        RECT 85.725 84.245 87.075 85.155 ;
        RECT 87.115 84.330 87.545 85.115 ;
        RECT 87.605 84.925 88.955 85.155 ;
        RECT 90.490 84.925 91.400 85.145 ;
        RECT 95.695 84.925 96.625 85.155 ;
        RECT 87.605 84.245 94.915 84.925 ;
        RECT 95.695 84.245 97.530 84.925 ;
        RECT 97.685 84.245 99.035 85.155 ;
        RECT 99.985 84.955 100.935 85.155 ;
        RECT 102.265 84.955 103.195 85.155 ;
        RECT 99.985 84.475 103.195 84.955 ;
        RECT 99.985 84.275 103.050 84.475 ;
        RECT 99.985 84.245 100.920 84.275 ;
        RECT 22.845 84.035 23.015 84.245 ;
        RECT 24.225 84.035 24.395 84.245 ;
        RECT 26.985 84.055 27.155 84.225 ;
        RECT 27.445 84.035 27.615 84.225 ;
        RECT 29.745 84.055 29.915 84.245 ;
        RECT 35.270 84.225 35.440 84.245 ;
        RECT 36.190 84.225 36.355 84.245 ;
        RECT 31.135 84.080 31.295 84.190 ;
        RECT 32.965 84.035 33.135 84.225 ;
        RECT 33.425 84.035 33.595 84.225 ;
        RECT 35.260 84.055 35.440 84.225 ;
        RECT 36.185 84.055 36.355 84.225 ;
        RECT 36.655 84.080 36.815 84.190 ;
        RECT 40.325 84.055 40.495 84.245 ;
        RECT 40.785 84.055 40.955 84.225 ;
        RECT 42.175 84.090 42.335 84.200 ;
        RECT 35.260 84.035 35.430 84.055 ;
        RECT 42.620 84.035 42.790 84.225 ;
        RECT 43.090 84.035 43.260 84.225 ;
        RECT 44.010 84.055 44.180 84.245 ;
        RECT 45.385 84.055 45.555 84.225 ;
        RECT 45.845 84.055 46.015 84.245 ;
        RECT 49.075 84.080 49.235 84.190 ;
        RECT 49.990 84.035 50.160 84.225 ;
        RECT 50.450 84.055 50.620 84.245 ;
        RECT 50.915 84.090 51.075 84.200 ;
        RECT 52.745 84.055 52.915 84.225 ;
        RECT 53.205 84.055 53.375 84.245 ;
        RECT 55.510 84.225 55.675 84.245 ;
        RECT 55.040 84.085 55.160 84.195 ;
        RECT 55.505 84.055 55.675 84.225 ;
        RECT 57.805 84.055 57.975 84.245 ;
        RECT 60.105 84.055 60.275 84.245 ;
        RECT 61.945 84.055 62.115 84.245 ;
        RECT 62.405 84.035 62.575 84.225 ;
        RECT 62.865 84.035 63.035 84.225 ;
        RECT 64.705 84.055 64.875 84.245 ;
        RECT 66.995 84.055 67.165 84.245 ;
        RECT 70.225 84.055 70.395 84.245 ;
        RECT 72.065 84.055 72.235 84.225 ;
        RECT 72.065 84.035 72.230 84.055 ;
        RECT 73.450 84.035 73.620 84.225 ;
        RECT 73.900 84.085 74.020 84.195 ;
        RECT 74.825 84.035 74.995 84.245 ;
        RECT 79.425 84.225 79.575 84.245 ;
        RECT 79.425 84.055 79.595 84.225 ;
        RECT 79.885 84.055 80.055 84.245 ;
        RECT 80.345 84.035 80.515 84.225 ;
        RECT 82.640 84.055 82.810 84.245 ;
        RECT 83.105 84.055 83.275 84.245 ;
        RECT 83.565 84.035 83.735 84.225 ;
        RECT 86.790 84.055 86.960 84.245 ;
        RECT 89.085 84.055 89.255 84.225 ;
        RECT 91.380 84.085 91.500 84.195 ;
        RECT 94.605 84.055 94.775 84.245 ;
        RECT 97.365 84.225 97.530 84.245 ;
        RECT 98.750 84.225 98.920 84.245 ;
        RECT 95.060 84.085 95.180 84.195 ;
        RECT 97.365 84.055 97.535 84.225 ;
        RECT 98.745 84.055 98.920 84.225 ;
        RECT 99.215 84.080 99.375 84.200 ;
        RECT 100.580 84.085 100.700 84.195 ;
        RECT 89.090 84.035 89.255 84.055 ;
        RECT 98.745 84.035 98.915 84.055 ;
        RECT 101.045 84.035 101.215 84.225 ;
        RECT 102.880 84.055 103.050 84.275 ;
        RECT 103.205 84.245 105.955 85.055 ;
        RECT 105.965 84.245 107.315 85.155 ;
        RECT 107.345 84.245 112.855 85.055 ;
        RECT 112.875 84.330 113.305 85.115 ;
        RECT 113.325 84.245 118.835 85.055 ;
        RECT 118.845 84.245 124.355 85.055 ;
        RECT 124.365 84.245 127.115 85.055 ;
        RECT 127.125 84.245 128.495 85.025 ;
        RECT 132.020 84.925 132.930 85.145 ;
        RECT 134.465 84.925 135.815 85.155 ;
        RECT 136.915 84.925 137.845 85.155 ;
        RECT 128.505 84.245 135.815 84.925 ;
        RECT 136.010 84.245 137.845 84.925 ;
        RECT 138.635 84.330 139.065 85.115 ;
        RECT 140.005 84.955 140.935 85.155 ;
        RECT 142.265 84.955 143.215 85.155 ;
        RECT 140.005 84.475 143.215 84.955 ;
        RECT 140.150 84.275 143.215 84.475 ;
        RECT 103.345 84.055 103.515 84.245 ;
        RECT 105.645 84.055 105.815 84.225 ;
        RECT 107.030 84.055 107.200 84.245 ;
        RECT 107.485 84.055 107.655 84.245 ;
        RECT 105.615 84.035 105.815 84.055 ;
        RECT 22.705 83.225 24.075 84.035 ;
        RECT 24.085 83.225 25.915 84.035 ;
        RECT 27.305 83.225 30.975 84.035 ;
        RECT 31.905 83.255 33.275 84.035 ;
        RECT 33.285 83.225 35.115 84.035 ;
        RECT 35.145 83.125 36.495 84.035 ;
        RECT 37.425 83.355 42.935 84.035 ;
        RECT 42.945 83.355 48.455 84.035 ;
        RECT 37.425 83.125 38.815 83.355 ;
        RECT 47.065 83.125 48.455 83.355 ;
        RECT 48.475 83.165 48.905 83.950 ;
        RECT 49.845 83.355 55.355 84.035 ;
        RECT 53.965 83.125 55.355 83.355 ;
        RECT 55.405 83.355 62.715 84.035 ;
        RECT 62.725 83.355 70.035 84.035 ;
        RECT 55.405 83.125 56.755 83.355 ;
        RECT 58.290 83.135 59.200 83.355 ;
        RECT 66.240 83.135 67.150 83.355 ;
        RECT 68.685 83.125 70.035 83.355 ;
        RECT 70.395 83.355 72.230 84.035 ;
        RECT 70.395 83.125 71.325 83.355 ;
        RECT 72.385 83.125 73.735 84.035 ;
        RECT 74.235 83.165 74.665 83.950 ;
        RECT 74.685 83.225 80.195 84.035 ;
        RECT 80.205 83.225 82.035 84.035 ;
        RECT 83.425 83.225 88.935 84.035 ;
        RECT 89.090 83.355 90.925 84.035 ;
        RECT 89.995 83.125 90.925 83.355 ;
        RECT 91.745 83.355 99.055 84.035 ;
        RECT 91.745 83.125 93.095 83.355 ;
        RECT 94.630 83.135 95.540 83.355 ;
        RECT 99.995 83.165 100.425 83.950 ;
        RECT 100.905 83.255 102.275 84.035 ;
        RECT 102.285 83.355 105.815 84.035 ;
        RECT 105.965 84.005 106.900 84.035 ;
        RECT 108.860 84.005 109.030 84.225 ;
        RECT 109.325 84.055 109.495 84.225 ;
        RECT 112.545 84.055 112.715 84.225 ;
        RECT 105.965 83.805 109.030 84.005 ;
        RECT 109.330 84.035 109.495 84.055 ;
        RECT 113.005 84.035 113.175 84.225 ;
        RECT 113.465 84.055 113.635 84.245 ;
        RECT 115.765 84.055 115.935 84.225 ;
        RECT 116.220 84.085 116.340 84.195 ;
        RECT 117.605 84.055 117.775 84.225 ;
        RECT 118.060 84.085 118.180 84.195 ;
        RECT 118.530 84.035 118.700 84.225 ;
        RECT 118.985 84.055 119.155 84.245 ;
        RECT 124.040 84.085 124.160 84.195 ;
        RECT 124.505 84.055 124.675 84.245 ;
        RECT 125.425 84.035 125.595 84.225 ;
        RECT 127.265 84.055 127.435 84.245 ;
        RECT 128.185 84.035 128.355 84.225 ;
        RECT 128.645 84.055 128.815 84.245 ;
        RECT 136.010 84.225 136.175 84.245 ;
        RECT 128.650 84.035 128.815 84.055 ;
        RECT 130.945 84.035 131.115 84.225 ;
        RECT 133.705 84.055 133.875 84.225 ;
        RECT 134.160 84.085 134.280 84.195 ;
        RECT 135.550 84.035 135.720 84.225 ;
        RECT 136.005 84.035 136.175 84.225 ;
        RECT 138.300 84.085 138.420 84.195 ;
        RECT 139.235 84.090 139.395 84.200 ;
        RECT 140.150 84.055 140.320 84.275 ;
        RECT 142.280 84.245 143.215 84.275 ;
        RECT 143.225 84.245 145.975 85.055 ;
        RECT 145.985 84.245 147.335 85.155 ;
        RECT 147.365 84.245 148.735 85.055 ;
        RECT 149.055 84.925 149.985 85.155 ;
        RECT 149.055 84.245 150.890 84.925 ;
        RECT 151.045 84.245 154.715 85.055 ;
        RECT 155.645 84.245 157.015 85.055 ;
        RECT 102.285 83.125 105.110 83.355 ;
        RECT 105.965 83.325 109.175 83.805 ;
        RECT 109.330 83.355 111.165 84.035 ;
        RECT 105.965 83.125 106.915 83.325 ;
        RECT 108.245 83.125 109.175 83.325 ;
        RECT 110.235 83.125 111.165 83.355 ;
        RECT 112.865 83.225 114.695 84.035 ;
        RECT 118.385 83.355 123.895 84.035 ;
        RECT 122.505 83.125 123.895 83.355 ;
        RECT 124.365 83.255 125.735 84.035 ;
        RECT 125.755 83.165 126.185 83.950 ;
        RECT 126.205 83.355 128.495 84.035 ;
        RECT 128.650 83.355 130.485 84.035 ;
        RECT 126.205 83.125 127.125 83.355 ;
        RECT 129.555 83.125 130.485 83.355 ;
        RECT 130.805 83.225 132.635 84.035 ;
        RECT 134.485 83.125 135.835 84.035 ;
        RECT 135.865 83.225 141.375 84.035 ;
        RECT 141.530 84.005 141.700 84.225 ;
        RECT 143.365 84.055 143.535 84.245 ;
        RECT 145.665 84.035 145.835 84.225 ;
        RECT 146.125 84.035 146.295 84.225 ;
        RECT 147.050 84.055 147.220 84.245 ;
        RECT 147.505 84.055 147.675 84.245 ;
        RECT 150.725 84.225 150.890 84.245 ;
        RECT 148.430 84.035 148.600 84.225 ;
        RECT 148.885 84.035 149.055 84.225 ;
        RECT 150.725 84.055 150.895 84.225 ;
        RECT 151.185 84.055 151.355 84.245 ;
        RECT 152.105 84.035 152.275 84.225 ;
        RECT 154.875 84.090 155.035 84.200 ;
        RECT 156.705 84.035 156.875 84.245 ;
        RECT 143.660 84.005 144.595 84.035 ;
        RECT 141.530 83.805 144.595 84.005 ;
        RECT 141.385 83.325 144.595 83.805 ;
        RECT 141.385 83.125 142.315 83.325 ;
        RECT 143.645 83.125 144.595 83.325 ;
        RECT 144.615 83.125 145.965 84.035 ;
        RECT 145.985 83.255 147.355 84.035 ;
        RECT 147.365 83.125 148.715 84.035 ;
        RECT 148.745 83.225 151.495 84.035 ;
        RECT 151.515 83.165 151.945 83.950 ;
        RECT 151.965 83.225 155.635 84.035 ;
        RECT 155.645 83.225 157.015 84.035 ;
      LAYER nwell ;
        RECT 22.510 80.005 157.210 82.835 ;
      LAYER pwell ;
        RECT 22.705 78.805 24.075 79.615 ;
        RECT 24.085 78.805 26.835 79.615 ;
        RECT 26.845 78.805 28.215 79.585 ;
        RECT 31.740 79.485 32.650 79.705 ;
        RECT 34.185 79.485 35.535 79.715 ;
        RECT 28.225 78.805 35.535 79.485 ;
        RECT 35.595 78.890 36.025 79.675 ;
        RECT 37.095 79.485 38.025 79.715 ;
        RECT 44.765 79.485 46.155 79.715 ;
        RECT 36.190 78.805 38.025 79.485 ;
        RECT 40.645 78.805 46.155 79.485 ;
        RECT 46.185 78.805 47.535 79.715 ;
        RECT 47.545 78.805 49.375 79.615 ;
        RECT 49.845 78.805 51.195 79.715 ;
        RECT 51.225 78.805 54.145 79.715 ;
        RECT 54.445 78.805 55.795 79.715 ;
        RECT 55.825 78.805 57.195 79.615 ;
        RECT 57.225 78.805 58.575 79.715 ;
        RECT 59.045 78.805 60.415 79.585 ;
        RECT 61.355 78.890 61.785 79.675 ;
        RECT 61.805 78.805 64.555 79.615 ;
        RECT 65.025 78.805 66.395 79.585 ;
        RECT 66.405 78.805 70.075 79.615 ;
        RECT 70.085 78.805 71.455 79.615 ;
        RECT 76.965 79.485 78.355 79.715 ;
        RECT 80.335 79.485 81.265 79.715 ;
        RECT 85.705 79.485 87.095 79.715 ;
        RECT 72.845 78.805 78.355 79.485 ;
        RECT 79.430 78.805 81.265 79.485 ;
        RECT 81.585 78.805 87.095 79.485 ;
        RECT 87.115 78.890 87.545 79.675 ;
        RECT 91.685 79.485 93.075 79.715 ;
        RECT 87.565 78.805 93.075 79.485 ;
        RECT 93.085 78.805 94.915 79.615 ;
        RECT 96.755 79.485 97.675 79.715 ;
        RECT 95.385 78.805 97.675 79.485 ;
        RECT 97.685 78.805 99.055 79.585 ;
        RECT 99.065 78.805 100.895 79.615 ;
        RECT 104.420 79.485 105.330 79.705 ;
        RECT 106.865 79.485 108.215 79.715 ;
        RECT 100.905 78.805 108.215 79.485 ;
        RECT 108.265 78.805 109.635 79.615 ;
        RECT 109.645 78.805 110.995 79.715 ;
        RECT 111.025 78.805 112.855 79.615 ;
        RECT 112.875 78.890 113.305 79.675 ;
        RECT 118.365 79.485 119.755 79.715 ;
        RECT 124.660 79.485 125.570 79.705 ;
        RECT 127.105 79.485 128.455 79.715 ;
        RECT 114.245 78.805 119.755 79.485 ;
        RECT 121.145 78.805 128.455 79.485 ;
        RECT 128.525 78.805 129.875 79.715 ;
        RECT 136.765 79.485 138.155 79.715 ;
        RECT 132.645 78.805 138.155 79.485 ;
        RECT 138.635 78.890 139.065 79.675 ;
        RECT 139.085 78.805 140.915 79.615 ;
        RECT 141.770 79.485 144.595 79.715 ;
        RECT 148.580 79.485 149.490 79.705 ;
        RECT 151.025 79.485 152.375 79.715 ;
        RECT 141.065 78.805 144.595 79.485 ;
        RECT 145.065 78.805 152.375 79.485 ;
        RECT 152.425 78.805 155.175 79.615 ;
        RECT 155.645 78.805 157.015 79.615 ;
        RECT 22.845 78.595 23.015 78.805 ;
        RECT 24.225 78.595 24.395 78.805 ;
        RECT 25.610 78.595 25.780 78.785 ;
        RECT 27.905 78.615 28.075 78.805 ;
        RECT 28.365 78.615 28.535 78.805 ;
        RECT 36.190 78.785 36.355 78.805 ;
        RECT 31.125 78.595 31.295 78.785 ;
        RECT 32.505 78.615 32.675 78.785 ;
        RECT 33.895 78.640 34.055 78.750 ;
        RECT 35.730 78.595 35.900 78.785 ;
        RECT 36.185 78.595 36.355 78.785 ;
        RECT 38.495 78.650 38.655 78.760 ;
        RECT 39.405 78.615 39.575 78.785 ;
        RECT 40.790 78.615 40.960 78.805 ;
        RECT 41.705 78.595 41.875 78.785 ;
        RECT 43.545 78.595 43.715 78.785 ;
        RECT 45.845 78.595 46.015 78.785 ;
        RECT 46.305 78.595 46.475 78.785 ;
        RECT 47.220 78.615 47.390 78.805 ;
        RECT 47.685 78.615 47.855 78.805 ;
        RECT 48.140 78.645 48.260 78.755 ;
        RECT 49.520 78.645 49.640 78.755 ;
        RECT 50.910 78.615 51.080 78.805 ;
        RECT 51.370 78.615 51.540 78.805 ;
        RECT 22.705 77.785 24.075 78.595 ;
        RECT 24.085 77.785 25.455 78.595 ;
        RECT 25.465 77.915 30.975 78.595 ;
        RECT 29.585 77.685 30.975 77.915 ;
        RECT 30.985 77.785 32.355 78.595 ;
        RECT 34.665 77.685 36.015 78.595 ;
        RECT 36.045 77.785 41.555 78.595 ;
        RECT 41.565 77.785 43.395 78.595 ;
        RECT 43.405 77.815 44.775 78.595 ;
        RECT 44.785 77.815 46.155 78.595 ;
        RECT 46.165 77.785 47.995 78.595 ;
        RECT 48.925 78.565 49.860 78.595 ;
        RECT 51.820 78.565 51.990 78.785 ;
        RECT 52.285 78.615 52.455 78.785 ;
        RECT 54.590 78.615 54.760 78.805 ;
        RECT 48.475 77.725 48.905 78.510 ;
        RECT 48.925 78.365 51.990 78.565 ;
        RECT 52.290 78.595 52.455 78.615 ;
        RECT 55.965 78.595 56.135 78.805 ;
        RECT 56.420 78.645 56.540 78.755 ;
        RECT 56.890 78.595 57.060 78.785 ;
        RECT 57.340 78.615 57.510 78.805 ;
        RECT 58.720 78.645 58.840 78.755 ;
        RECT 59.185 78.615 59.355 78.805 ;
        RECT 60.575 78.650 60.735 78.760 ;
        RECT 61.945 78.615 62.115 78.805 ;
        RECT 63.325 78.615 63.495 78.785 ;
        RECT 63.785 78.595 63.955 78.785 ;
        RECT 64.700 78.645 64.820 78.755 ;
        RECT 66.085 78.615 66.255 78.805 ;
        RECT 66.545 78.755 66.715 78.805 ;
        RECT 66.540 78.645 66.715 78.755 ;
        RECT 66.545 78.615 66.715 78.645 ;
        RECT 67.925 78.615 68.095 78.785 ;
        RECT 69.305 78.615 69.475 78.785 ;
        RECT 69.765 78.595 69.935 78.785 ;
        RECT 70.225 78.615 70.395 78.805 ;
        RECT 72.990 78.785 73.160 78.805 ;
        RECT 79.430 78.785 79.595 78.805 ;
        RECT 71.605 78.615 71.775 78.785 ;
        RECT 72.520 78.645 72.640 78.755 ;
        RECT 72.985 78.615 73.160 78.785 ;
        RECT 74.820 78.645 74.940 78.755 ;
        RECT 72.985 78.595 73.155 78.615 ;
        RECT 75.280 78.595 75.450 78.785 ;
        RECT 76.670 78.595 76.840 78.785 ;
        RECT 78.515 78.650 78.675 78.760 ;
        RECT 79.425 78.615 79.595 78.785 ;
        RECT 80.800 78.595 80.970 78.785 ;
        RECT 81.265 78.595 81.435 78.785 ;
        RECT 81.730 78.615 81.900 78.805 ;
        RECT 83.105 78.595 83.275 78.785 ;
        RECT 84.955 78.640 85.115 78.750 ;
        RECT 85.865 78.595 86.035 78.785 ;
        RECT 87.710 78.615 87.880 78.805 ;
        RECT 88.165 78.615 88.335 78.785 ;
        RECT 88.635 78.640 88.795 78.750 ;
        RECT 89.545 78.615 89.715 78.785 ;
        RECT 90.930 78.595 91.100 78.785 ;
        RECT 93.225 78.615 93.395 78.805 ;
        RECT 95.060 78.645 95.180 78.755 ;
        RECT 95.525 78.615 95.695 78.805 ;
        RECT 96.445 78.595 96.615 78.785 ;
        RECT 98.745 78.615 98.915 78.805 ;
        RECT 99.205 78.615 99.375 78.805 ;
        RECT 100.585 78.595 100.755 78.785 ;
        RECT 101.045 78.615 101.215 78.805 ;
        RECT 102.885 78.615 103.055 78.785 ;
        RECT 103.345 78.595 103.515 78.785 ;
        RECT 108.405 78.615 108.575 78.805 ;
        RECT 108.870 78.595 109.040 78.785 ;
        RECT 109.790 78.615 109.960 78.805 ;
        RECT 111.165 78.615 111.335 78.805 ;
        RECT 113.475 78.650 113.635 78.760 ;
        RECT 114.390 78.755 114.560 78.805 ;
        RECT 114.380 78.645 114.560 78.755 ;
        RECT 114.390 78.615 114.560 78.645 ;
        RECT 114.845 78.595 115.015 78.785 ;
        RECT 116.230 78.595 116.400 78.785 ;
        RECT 120.825 78.615 120.995 78.785 ;
        RECT 121.285 78.615 121.455 78.805 ;
        RECT 121.745 78.595 121.915 78.785 ;
        RECT 125.420 78.645 125.540 78.755 ;
        RECT 126.345 78.595 126.515 78.785 ;
        RECT 128.640 78.615 128.810 78.805 ;
        RECT 129.105 78.595 129.275 78.785 ;
        RECT 130.035 78.650 130.195 78.760 ;
        RECT 130.490 78.595 130.660 78.785 ;
        RECT 131.865 78.615 132.035 78.785 ;
        RECT 132.320 78.645 132.440 78.755 ;
        RECT 132.790 78.615 132.960 78.805 ;
        RECT 136.925 78.595 137.095 78.785 ;
        RECT 137.385 78.595 137.555 78.785 ;
        RECT 138.300 78.645 138.420 78.755 ;
        RECT 139.225 78.615 139.395 78.805 ;
        RECT 141.065 78.785 141.265 78.805 ;
        RECT 48.925 77.885 52.135 78.365 ;
        RECT 52.290 77.915 54.125 78.595 ;
        RECT 54.445 77.915 56.275 78.595 ;
        RECT 56.745 77.915 62.255 78.595 ;
        RECT 48.925 77.685 49.875 77.885 ;
        RECT 51.205 77.685 52.135 77.885 ;
        RECT 53.195 77.685 54.125 77.915 ;
        RECT 60.865 77.685 62.255 77.915 ;
        RECT 63.645 77.785 66.395 78.595 ;
        RECT 69.625 77.785 72.375 78.595 ;
        RECT 72.845 77.815 74.215 78.595 ;
        RECT 74.235 77.725 74.665 78.510 ;
        RECT 75.165 77.685 76.515 78.595 ;
        RECT 76.525 77.685 77.875 78.595 ;
        RECT 78.195 77.685 81.115 78.595 ;
        RECT 81.125 77.915 82.955 78.595 ;
        RECT 82.965 77.915 84.795 78.595 ;
        RECT 85.725 77.815 87.095 78.595 ;
        RECT 90.785 77.915 96.295 78.595 ;
        RECT 94.905 77.685 96.295 77.915 ;
        RECT 96.305 77.785 99.975 78.595 ;
        RECT 99.995 77.725 100.425 78.510 ;
        RECT 100.445 77.785 101.815 78.595 ;
        RECT 103.205 77.785 108.715 78.595 ;
        RECT 108.725 77.915 114.235 78.595 ;
        RECT 112.845 77.685 114.235 77.915 ;
        RECT 114.705 77.815 116.075 78.595 ;
        RECT 116.085 77.915 121.595 78.595 ;
        RECT 120.205 77.685 121.595 77.915 ;
        RECT 121.605 77.785 125.275 78.595 ;
        RECT 125.755 77.725 126.185 78.510 ;
        RECT 126.205 77.785 128.955 78.595 ;
        RECT 128.965 77.815 130.335 78.595 ;
        RECT 130.345 77.915 135.855 78.595 ;
        RECT 134.465 77.685 135.855 77.915 ;
        RECT 135.865 77.815 137.235 78.595 ;
        RECT 137.245 77.785 139.995 78.595 ;
        RECT 140.150 78.565 140.320 78.785 ;
        RECT 141.065 78.615 141.235 78.785 ;
        RECT 143.365 78.595 143.535 78.785 ;
        RECT 145.205 78.755 145.375 78.805 ;
        RECT 144.740 78.645 144.860 78.755 ;
        RECT 145.200 78.645 145.375 78.755 ;
        RECT 145.205 78.615 145.375 78.645 ;
        RECT 147.505 78.615 147.675 78.785 ;
        RECT 147.505 78.595 147.670 78.615 ;
        RECT 147.965 78.595 148.135 78.785 ;
        RECT 152.105 78.595 152.275 78.785 ;
        RECT 152.565 78.615 152.735 78.805 ;
        RECT 155.320 78.645 155.440 78.755 ;
        RECT 156.705 78.595 156.875 78.805 ;
        RECT 142.280 78.565 143.215 78.595 ;
        RECT 140.150 78.365 143.215 78.565 ;
        RECT 140.005 77.885 143.215 78.365 ;
        RECT 140.005 77.685 140.935 77.885 ;
        RECT 142.265 77.685 143.215 77.885 ;
        RECT 143.225 77.785 145.055 78.595 ;
        RECT 145.835 77.915 147.670 78.595 ;
        RECT 145.835 77.685 146.765 77.915 ;
        RECT 147.825 77.785 151.495 78.595 ;
        RECT 151.515 77.725 151.945 78.510 ;
        RECT 151.965 77.785 155.635 78.595 ;
        RECT 155.645 77.785 157.015 78.595 ;
      LAYER nwell ;
        RECT 22.510 74.565 157.210 77.395 ;
      LAYER pwell ;
        RECT 22.705 73.365 24.075 74.175 ;
        RECT 24.085 73.365 25.915 74.175 ;
        RECT 31.885 74.045 33.275 74.275 ;
        RECT 27.765 73.365 33.275 74.045 ;
        RECT 34.205 73.365 35.575 74.145 ;
        RECT 35.595 73.450 36.025 74.235 ;
        RECT 40.165 74.045 41.555 74.275 ;
        RECT 36.045 73.365 41.555 74.045 ;
        RECT 41.585 73.365 42.935 74.275 ;
        RECT 42.945 73.365 48.455 74.175 ;
        RECT 48.465 73.365 50.295 74.175 ;
        RECT 50.325 73.365 51.675 74.275 ;
        RECT 51.685 73.365 55.355 74.175 ;
        RECT 55.380 74.045 56.750 74.275 ;
        RECT 55.380 73.365 57.655 74.045 ;
        RECT 57.665 73.365 60.875 74.275 ;
        RECT 61.355 73.450 61.785 74.235 ;
        RECT 62.115 74.045 63.045 74.275 ;
        RECT 62.115 73.365 63.950 74.045 ;
        RECT 64.105 73.365 65.455 74.275 ;
        RECT 65.485 73.365 66.855 74.175 ;
        RECT 70.985 74.045 72.375 74.275 ;
        RECT 66.865 73.365 72.375 74.045 ;
        RECT 72.385 73.365 73.735 74.275 ;
        RECT 73.765 73.365 75.135 74.175 ;
        RECT 75.145 74.075 76.095 74.275 ;
        RECT 77.425 74.075 78.355 74.275 ;
        RECT 75.145 73.595 78.355 74.075 ;
        RECT 75.145 73.395 78.210 73.595 ;
        RECT 75.145 73.365 76.080 73.395 ;
        RECT 22.845 73.155 23.015 73.365 ;
        RECT 24.225 73.155 24.395 73.365 ;
        RECT 26.060 73.205 26.180 73.315 ;
        RECT 26.525 73.175 26.695 73.345 ;
        RECT 27.910 73.175 28.080 73.365 ;
        RECT 29.745 73.155 29.915 73.345 ;
        RECT 33.435 73.210 33.595 73.320 ;
        RECT 34.345 73.175 34.515 73.365 ;
        RECT 35.265 73.155 35.435 73.345 ;
        RECT 36.190 73.175 36.360 73.365 ;
        RECT 38.025 73.155 38.195 73.345 ;
        RECT 41.705 73.155 41.875 73.345 ;
        RECT 42.175 73.200 42.335 73.310 ;
        RECT 42.620 73.175 42.790 73.365 ;
        RECT 43.085 73.345 43.255 73.365 ;
        RECT 43.080 73.175 43.255 73.345 ;
        RECT 22.705 72.345 24.075 73.155 ;
        RECT 24.085 72.345 29.595 73.155 ;
        RECT 29.605 72.345 35.115 73.155 ;
        RECT 35.125 72.345 37.875 73.155 ;
        RECT 37.895 72.245 39.245 73.155 ;
        RECT 39.275 72.245 42.005 73.155 ;
        RECT 43.080 73.125 43.250 73.175 ;
        RECT 45.385 73.155 45.555 73.345 ;
        RECT 48.140 73.205 48.260 73.315 ;
        RECT 48.605 73.175 48.775 73.365 ;
        RECT 49.065 73.155 49.235 73.345 ;
        RECT 50.440 73.175 50.610 73.365 ;
        RECT 51.360 73.155 51.530 73.345 ;
        RECT 51.825 73.315 51.995 73.365 ;
        RECT 51.820 73.205 51.995 73.315 ;
        RECT 51.825 73.175 51.995 73.205 ;
        RECT 44.280 73.125 45.235 73.155 ;
        RECT 42.955 72.445 45.235 73.125 ;
        RECT 44.280 72.245 45.235 72.445 ;
        RECT 45.245 72.345 47.995 73.155 ;
        RECT 48.475 72.285 48.905 73.070 ;
        RECT 48.925 72.345 50.295 73.155 ;
        RECT 50.325 72.245 51.675 73.155 ;
        RECT 52.145 73.125 53.100 73.155 ;
        RECT 54.130 73.125 54.300 73.345 ;
        RECT 54.585 73.155 54.755 73.345 ;
        RECT 55.965 73.155 56.135 73.345 ;
        RECT 57.340 73.175 57.510 73.365 ;
        RECT 57.795 73.175 57.965 73.365 ;
        RECT 63.785 73.345 63.950 73.365 ;
        RECT 58.260 73.155 58.430 73.345 ;
        RECT 58.725 73.155 58.895 73.345 ;
        RECT 60.560 73.205 60.680 73.315 ;
        RECT 61.020 73.155 61.190 73.345 ;
        RECT 62.405 73.155 62.575 73.345 ;
        RECT 63.785 73.175 63.955 73.345 ;
        RECT 64.250 73.175 64.420 73.365 ;
        RECT 65.625 73.345 65.795 73.365 ;
        RECT 65.160 73.205 65.280 73.315 ;
        RECT 65.625 73.175 65.800 73.345 ;
        RECT 67.010 73.175 67.180 73.365 ;
        RECT 65.630 73.155 65.800 73.175 ;
        RECT 71.145 73.155 71.315 73.345 ;
        RECT 72.530 73.175 72.700 73.365 ;
        RECT 73.905 73.315 74.075 73.365 ;
        RECT 73.900 73.205 74.075 73.315 ;
        RECT 73.905 73.175 74.075 73.205 ;
        RECT 74.820 73.155 74.990 73.345 ;
        RECT 76.205 73.155 76.375 73.345 ;
        RECT 78.040 73.175 78.210 73.395 ;
        RECT 78.365 73.365 82.035 74.175 ;
        RECT 82.985 73.365 84.335 74.275 ;
        RECT 84.345 73.365 85.715 74.175 ;
        RECT 85.735 73.365 87.085 74.275 ;
        RECT 87.115 73.450 87.545 74.235 ;
        RECT 88.025 74.075 88.980 74.275 ;
        RECT 88.025 73.395 90.305 74.075 ;
        RECT 88.025 73.365 88.980 73.395 ;
        RECT 78.505 73.175 78.675 73.365 ;
        RECT 78.960 73.205 79.080 73.315 ;
        RECT 79.425 73.155 79.595 73.345 ;
        RECT 82.185 73.175 82.355 73.345 ;
        RECT 84.020 73.175 84.190 73.365 ;
        RECT 82.205 73.155 82.355 73.175 ;
        RECT 84.485 73.155 84.655 73.365 ;
        RECT 85.865 73.175 86.035 73.365 ;
        RECT 90.010 73.345 90.180 73.395 ;
        RECT 90.325 73.365 91.695 74.145 ;
        RECT 91.705 73.365 94.455 74.175 ;
        RECT 94.945 73.365 96.295 74.275 ;
        RECT 97.445 74.185 98.395 74.275 ;
        RECT 96.465 73.365 98.395 74.185 ;
        RECT 100.400 74.075 101.355 74.275 ;
        RECT 99.075 73.395 101.355 74.075 ;
        RECT 105.485 74.045 106.875 74.275 ;
        RECT 107.935 74.045 108.865 74.275 ;
        RECT 52.145 72.445 54.425 73.125 ;
        RECT 52.145 72.245 53.100 72.445 ;
        RECT 54.455 72.245 55.805 73.155 ;
        RECT 55.825 72.345 57.195 73.155 ;
        RECT 57.225 72.245 58.575 73.155 ;
        RECT 58.585 72.345 60.415 73.155 ;
        RECT 60.905 72.245 62.255 73.155 ;
        RECT 62.265 72.345 65.015 73.155 ;
        RECT 65.485 72.475 70.995 73.155 ;
        RECT 69.605 72.245 70.995 72.475 ;
        RECT 71.005 72.345 73.755 73.155 ;
        RECT 74.235 72.285 74.665 73.070 ;
        RECT 74.705 72.245 76.055 73.155 ;
        RECT 76.065 72.345 78.815 73.155 ;
        RECT 79.285 72.475 82.035 73.155 ;
        RECT 81.105 72.245 82.035 72.475 ;
        RECT 82.205 72.335 84.135 73.155 ;
        RECT 84.345 72.345 87.095 73.155 ;
        RECT 87.250 73.125 87.420 73.345 ;
        RECT 87.700 73.205 87.820 73.315 ;
        RECT 90.005 73.175 90.180 73.345 ;
        RECT 90.465 73.175 90.635 73.365 ;
        RECT 91.845 73.175 92.015 73.365 ;
        RECT 94.600 73.205 94.720 73.315 ;
        RECT 95.535 73.200 95.695 73.310 ;
        RECT 95.980 73.175 96.150 73.365 ;
        RECT 96.465 73.345 96.615 73.365 ;
        RECT 90.005 73.155 90.175 73.175 ;
        RECT 96.445 73.155 96.615 73.345 ;
        RECT 98.745 73.315 98.915 73.345 ;
        RECT 98.740 73.205 98.915 73.315 ;
        RECT 98.745 73.155 98.915 73.205 ;
        RECT 99.200 73.175 99.370 73.395 ;
        RECT 100.400 73.365 101.355 73.395 ;
        RECT 101.365 73.365 106.875 74.045 ;
        RECT 107.030 73.365 108.865 74.045 ;
        RECT 109.645 74.075 110.575 74.275 ;
        RECT 111.905 74.075 112.855 74.275 ;
        RECT 109.645 73.595 112.855 74.075 ;
        RECT 109.790 73.395 112.855 73.595 ;
        RECT 112.875 73.450 113.305 74.235 ;
        RECT 101.510 73.345 101.680 73.365 ;
        RECT 107.030 73.345 107.195 73.365 ;
        RECT 100.595 73.200 100.755 73.310 ;
        RECT 101.505 73.175 101.680 73.345 ;
        RECT 103.805 73.175 103.975 73.345 ;
        RECT 101.505 73.155 101.675 73.175 ;
        RECT 104.265 73.155 104.435 73.345 ;
        RECT 107.025 73.175 107.195 73.345 ;
        RECT 107.955 73.200 108.115 73.310 ;
        RECT 108.865 73.155 109.035 73.345 ;
        RECT 109.320 73.205 109.440 73.315 ;
        RECT 109.790 73.175 109.960 73.395 ;
        RECT 111.920 73.365 112.855 73.395 ;
        RECT 113.325 73.365 114.675 74.275 ;
        RECT 114.705 73.365 117.625 74.275 ;
        RECT 117.925 73.365 119.275 74.275 ;
        RECT 119.305 73.365 122.975 74.175 ;
        RECT 123.005 73.365 124.355 74.275 ;
        RECT 124.365 73.365 127.115 74.175 ;
        RECT 127.595 73.365 128.945 74.275 ;
        RECT 128.965 73.365 130.795 74.175 ;
        RECT 132.140 74.075 133.095 74.275 ;
        RECT 130.815 73.395 133.095 74.075 ;
        RECT 110.705 73.155 110.875 73.345 ;
        RECT 112.545 73.155 112.715 73.345 ;
        RECT 113.920 73.155 114.090 73.345 ;
        RECT 114.390 73.175 114.560 73.365 ;
        RECT 114.850 73.175 115.020 73.365 ;
        RECT 115.305 73.155 115.475 73.345 ;
        RECT 117.140 73.205 117.260 73.315 ;
        RECT 117.605 73.155 117.775 73.345 ;
        RECT 118.070 73.175 118.240 73.365 ;
        RECT 119.445 73.175 119.615 73.365 ;
        RECT 120.370 73.155 120.540 73.345 ;
        RECT 123.590 73.155 123.760 73.345 ;
        RECT 124.040 73.175 124.210 73.365 ;
        RECT 124.505 73.175 124.675 73.365 ;
        RECT 124.975 73.200 125.135 73.310 ;
        RECT 126.340 73.205 126.460 73.315 ;
        RECT 88.910 73.125 89.855 73.155 ;
        RECT 87.105 72.445 89.855 73.125 ;
        RECT 83.185 72.245 84.135 72.335 ;
        RECT 88.910 72.245 89.855 72.445 ;
        RECT 89.865 72.345 95.375 73.155 ;
        RECT 96.305 72.475 98.595 73.155 ;
        RECT 97.675 72.245 98.595 72.475 ;
        RECT 98.605 72.375 99.975 73.155 ;
        RECT 99.995 72.285 100.425 73.070 ;
        RECT 101.365 72.375 102.735 73.155 ;
        RECT 104.125 72.345 107.795 73.155 ;
        RECT 108.725 72.475 110.555 73.155 ;
        RECT 110.565 72.475 112.395 73.155 ;
        RECT 112.405 72.345 113.775 73.155 ;
        RECT 113.805 72.245 115.155 73.155 ;
        RECT 115.165 72.345 116.995 73.155 ;
        RECT 117.465 72.475 120.215 73.155 ;
        RECT 120.370 72.925 123.425 73.155 ;
        RECT 119.285 72.245 120.215 72.475 ;
        RECT 120.225 72.245 123.425 72.925 ;
        RECT 123.445 72.245 124.795 73.155 ;
        RECT 126.810 73.125 126.980 73.345 ;
        RECT 127.260 73.205 127.380 73.315 ;
        RECT 127.725 73.175 127.895 73.365 ;
        RECT 129.105 73.175 129.275 73.365 ;
        RECT 129.565 73.155 129.735 73.345 ;
        RECT 130.940 73.175 131.110 73.395 ;
        RECT 132.140 73.365 133.095 73.395 ;
        RECT 133.105 73.365 134.935 74.175 ;
        RECT 134.965 73.365 136.315 74.275 ;
        RECT 137.245 73.365 138.615 74.145 ;
        RECT 138.635 73.450 139.065 74.235 ;
        RECT 145.505 74.045 146.895 74.275 ;
        RECT 141.385 73.365 146.895 74.045 ;
        RECT 146.905 73.365 152.415 74.175 ;
        RECT 152.425 73.365 155.175 74.175 ;
        RECT 155.645 73.365 157.015 74.175 ;
        RECT 133.245 73.175 133.415 73.365 ;
        RECT 135.085 73.155 135.255 73.345 ;
        RECT 136.000 73.175 136.170 73.365 ;
        RECT 136.465 73.175 136.635 73.345 ;
        RECT 137.385 73.175 137.555 73.365 ;
        RECT 136.485 73.155 136.635 73.175 ;
        RECT 138.765 73.155 138.935 73.345 ;
        RECT 139.235 73.210 139.395 73.320 ;
        RECT 140.145 73.175 140.315 73.345 ;
        RECT 141.065 73.175 141.235 73.345 ;
        RECT 141.530 73.175 141.700 73.365 ;
        RECT 142.450 73.155 142.620 73.345 ;
        RECT 147.045 73.175 147.215 73.365 ;
        RECT 147.965 73.155 148.135 73.345 ;
        RECT 152.105 73.155 152.275 73.345 ;
        RECT 152.565 73.175 152.735 73.365 ;
        RECT 155.320 73.205 155.440 73.315 ;
        RECT 156.705 73.155 156.875 73.365 ;
        RECT 128.470 73.125 129.415 73.155 ;
        RECT 125.755 72.285 126.185 73.070 ;
        RECT 126.665 72.445 129.415 73.125 ;
        RECT 128.470 72.245 129.415 72.445 ;
        RECT 129.425 72.345 134.935 73.155 ;
        RECT 134.945 72.345 136.315 73.155 ;
        RECT 136.485 72.335 138.415 73.155 ;
        RECT 138.625 72.475 140.915 73.155 ;
        RECT 142.305 72.475 147.815 73.155 ;
        RECT 137.465 72.245 138.415 72.335 ;
        RECT 139.995 72.245 140.915 72.475 ;
        RECT 146.425 72.245 147.815 72.475 ;
        RECT 147.825 72.345 151.495 73.155 ;
        RECT 151.515 72.285 151.945 73.070 ;
        RECT 151.965 72.345 155.635 73.155 ;
        RECT 155.645 72.345 157.015 73.155 ;
      LAYER nwell ;
        RECT 22.510 69.125 157.210 71.955 ;
      LAYER pwell ;
        RECT 22.705 67.925 24.075 68.735 ;
        RECT 24.085 67.925 29.595 68.735 ;
        RECT 29.605 67.925 35.115 68.735 ;
        RECT 35.595 68.010 36.025 68.795 ;
        RECT 36.525 67.925 37.875 68.835 ;
        RECT 37.885 67.925 39.715 68.735 ;
        RECT 41.520 68.635 42.475 68.835 ;
        RECT 40.195 67.955 42.475 68.635 ;
        RECT 22.845 67.715 23.015 67.925 ;
        RECT 24.225 67.715 24.395 67.925 ;
        RECT 29.745 67.875 29.915 67.925 ;
        RECT 29.740 67.765 29.915 67.875 ;
        RECT 29.745 67.735 29.915 67.765 ;
        RECT 30.205 67.735 30.375 67.905 ;
        RECT 31.590 67.715 31.760 67.905 ;
        RECT 35.260 67.765 35.380 67.875 ;
        RECT 36.180 67.765 36.300 67.875 ;
        RECT 37.560 67.735 37.730 67.925 ;
        RECT 38.025 67.735 38.195 67.925 ;
        RECT 38.480 67.715 38.650 67.905 ;
        RECT 38.945 67.715 39.115 67.905 ;
        RECT 39.860 67.765 39.980 67.875 ;
        RECT 40.320 67.735 40.490 67.955 ;
        RECT 41.520 67.925 42.475 67.955 ;
        RECT 42.485 67.925 45.695 68.835 ;
        RECT 45.705 67.925 47.055 68.835 ;
        RECT 47.095 68.155 50.295 68.835 ;
        RECT 51.680 68.155 53.515 68.835 ;
        RECT 47.095 67.925 50.150 68.155 ;
        RECT 51.680 67.925 53.370 68.155 ;
        RECT 53.525 67.925 54.875 68.835 ;
        RECT 54.905 67.925 58.575 68.735 ;
        RECT 59.045 67.925 60.395 68.835 ;
        RECT 61.355 68.010 61.785 68.795 ;
        RECT 63.185 67.925 66.855 68.735 ;
        RECT 68.095 68.605 69.025 68.835 ;
        RECT 70.085 68.635 71.030 68.835 ;
        RECT 68.095 67.925 69.930 68.605 ;
        RECT 70.085 67.955 72.835 68.635 ;
        RECT 72.845 68.155 74.680 68.835 ;
        RECT 70.085 67.925 71.030 67.955 ;
        RECT 42.615 67.905 42.785 67.925 ;
        RECT 42.615 67.735 42.800 67.905 ;
        RECT 42.630 67.715 42.800 67.735 ;
        RECT 44.925 67.715 45.095 67.905 ;
        RECT 45.385 67.715 45.555 67.905 ;
        RECT 45.850 67.735 46.020 67.925 ;
        RECT 48.140 67.715 48.310 67.905 ;
        RECT 49.980 67.735 50.150 67.925 ;
        RECT 50.455 67.770 50.615 67.880 ;
        RECT 53.200 67.735 53.370 67.925 ;
        RECT 53.670 67.735 53.840 67.925 ;
        RECT 54.580 67.715 54.750 67.905 ;
        RECT 55.045 67.735 55.215 67.925 ;
        RECT 60.110 67.905 60.280 67.925 ;
        RECT 55.965 67.735 56.135 67.905 ;
        RECT 57.340 67.715 57.510 67.905 ;
        RECT 58.720 67.715 58.890 67.905 ;
        RECT 60.100 67.735 60.280 67.905 ;
        RECT 60.100 67.715 60.270 67.735 ;
        RECT 60.570 67.715 60.740 67.905 ;
        RECT 62.865 67.735 63.035 67.905 ;
        RECT 63.325 67.735 63.495 67.925 ;
        RECT 69.765 67.905 69.930 67.925 ;
        RECT 72.520 67.905 72.690 67.955 ;
        RECT 72.990 67.925 74.680 68.155 ;
        RECT 75.145 67.925 76.975 68.735 ;
        RECT 77.455 68.155 80.655 68.835 ;
        RECT 77.455 67.925 80.510 68.155 ;
        RECT 80.665 67.925 82.035 68.735 ;
        RECT 82.045 67.925 83.875 68.835 ;
        RECT 83.885 67.925 85.235 68.835 ;
        RECT 85.745 67.925 87.095 68.835 ;
        RECT 87.115 68.010 87.545 68.795 ;
        RECT 87.585 67.925 88.935 68.835 ;
        RECT 89.400 68.155 91.235 68.835 ;
        RECT 89.400 67.925 91.090 68.155 ;
        RECT 91.245 67.925 92.595 68.835 ;
        RECT 93.545 68.635 94.475 68.835 ;
        RECT 95.805 68.635 96.755 68.835 ;
        RECT 93.545 68.155 96.755 68.635 ;
        RECT 96.765 68.635 97.695 68.835 ;
        RECT 99.025 68.635 99.975 68.835 ;
        RECT 96.765 68.155 99.975 68.635 ;
        RECT 93.690 67.955 96.755 68.155 ;
        RECT 66.545 67.715 66.715 67.905 ;
        RECT 67.015 67.770 67.175 67.880 ;
        RECT 68.390 67.715 68.560 67.905 ;
        RECT 69.765 67.735 69.935 67.905 ;
        RECT 70.680 67.715 70.850 67.905 ;
        RECT 71.150 67.715 71.320 67.905 ;
        RECT 72.520 67.735 72.695 67.905 ;
        RECT 72.990 67.735 73.160 67.925 ;
        RECT 75.285 67.735 75.455 67.925 ;
        RECT 72.525 67.715 72.695 67.735 ;
        RECT 75.740 67.715 75.910 67.905 ;
        RECT 76.200 67.765 76.320 67.875 ;
        RECT 77.120 67.765 77.240 67.875 ;
        RECT 77.580 67.715 77.750 67.905 ;
        RECT 78.960 67.715 79.130 67.905 ;
        RECT 79.425 67.715 79.595 67.905 ;
        RECT 80.340 67.735 80.510 67.925 ;
        RECT 80.805 67.735 80.975 67.925 ;
        RECT 81.260 67.765 81.380 67.875 ;
        RECT 82.190 67.735 82.360 67.925 ;
        RECT 82.645 67.735 82.815 67.905 ;
        RECT 83.105 67.715 83.275 67.905 ;
        RECT 84.030 67.735 84.200 67.925 ;
        RECT 85.400 67.765 85.520 67.875 ;
        RECT 86.780 67.735 86.950 67.925 ;
        RECT 88.620 67.870 88.790 67.925 ;
        RECT 90.920 67.905 91.090 67.925 ;
        RECT 88.620 67.760 88.795 67.870 ;
        RECT 88.620 67.735 88.790 67.760 ;
        RECT 90.460 67.715 90.630 67.905 ;
        RECT 90.920 67.735 91.095 67.905 ;
        RECT 91.390 67.735 91.560 67.925 ;
        RECT 92.775 67.770 92.935 67.880 ;
        RECT 93.690 67.735 93.860 67.955 ;
        RECT 95.820 67.925 96.755 67.955 ;
        RECT 96.910 67.955 99.975 68.155 ;
        RECT 96.910 67.735 97.080 67.955 ;
        RECT 99.040 67.925 99.975 67.955 ;
        RECT 100.445 67.925 101.815 68.705 ;
        RECT 105.945 68.605 107.335 68.835 ;
        RECT 109.150 68.635 110.095 68.835 ;
        RECT 101.825 67.925 107.335 68.605 ;
        RECT 107.345 67.955 110.095 68.635 ;
        RECT 97.365 67.735 97.535 67.905 ;
        RECT 90.925 67.715 91.095 67.735 ;
        RECT 22.705 66.905 24.075 67.715 ;
        RECT 24.085 66.905 29.595 67.715 ;
        RECT 31.445 67.035 37.415 67.715 ;
        RECT 35.630 66.805 37.415 67.035 ;
        RECT 37.445 66.805 38.795 67.715 ;
        RECT 38.805 66.905 42.475 67.715 ;
        RECT 42.485 66.805 43.835 67.715 ;
        RECT 43.875 66.805 45.225 67.715 ;
        RECT 45.245 66.905 47.075 67.715 ;
        RECT 47.105 66.805 48.455 67.715 ;
        RECT 48.475 66.845 48.905 67.630 ;
        RECT 48.925 67.035 54.895 67.715 ;
        RECT 48.925 66.805 50.710 67.035 ;
        RECT 56.305 66.805 57.655 67.715 ;
        RECT 57.685 66.805 59.035 67.715 ;
        RECT 59.065 66.805 60.415 67.715 ;
        RECT 60.425 67.035 66.395 67.715 ;
        RECT 64.610 66.805 66.395 67.035 ;
        RECT 66.405 66.905 68.235 67.715 ;
        RECT 68.245 66.805 69.595 67.715 ;
        RECT 69.645 66.805 70.995 67.715 ;
        RECT 71.005 66.805 72.355 67.715 ;
        RECT 72.385 66.905 74.215 67.715 ;
        RECT 74.235 66.845 74.665 67.630 ;
        RECT 74.705 66.805 76.055 67.715 ;
        RECT 76.545 66.805 77.895 67.715 ;
        RECT 77.925 66.805 79.275 67.715 ;
        RECT 79.285 66.905 81.115 67.715 ;
        RECT 82.965 66.905 88.475 67.715 ;
        RECT 89.425 66.805 90.775 67.715 ;
        RECT 90.785 66.905 96.295 67.715 ;
        RECT 97.820 67.685 97.990 67.905 ;
        RECT 100.120 67.765 100.240 67.875 ;
        RECT 100.585 67.715 100.755 67.925 ;
        RECT 101.970 67.905 102.140 67.925 ;
        RECT 101.965 67.735 102.140 67.905 ;
        RECT 101.965 67.715 102.135 67.735 ;
        RECT 103.345 67.715 103.515 67.905 ;
        RECT 107.025 67.715 107.195 67.905 ;
        RECT 107.490 67.735 107.660 67.955 ;
        RECT 109.150 67.925 110.095 67.955 ;
        RECT 110.415 68.605 111.345 68.835 ;
        RECT 110.415 67.925 112.250 68.605 ;
        RECT 112.875 68.010 113.305 68.795 ;
        RECT 113.325 68.155 115.160 68.835 ;
        RECT 119.065 68.745 120.015 68.835 ;
        RECT 112.085 67.905 112.250 67.925 ;
        RECT 113.470 67.925 115.160 68.155 ;
        RECT 115.625 67.925 117.455 68.735 ;
        RECT 118.085 67.925 120.015 68.745 ;
        RECT 120.225 67.925 122.055 68.735 ;
        RECT 122.525 67.925 124.355 68.835 ;
        RECT 124.365 67.925 128.035 68.735 ;
        RECT 128.045 68.155 129.880 68.835 ;
        RECT 128.190 67.925 129.880 68.155 ;
        RECT 130.365 67.925 131.715 68.835 ;
        RECT 131.725 67.925 133.075 68.835 ;
        RECT 133.105 68.635 134.035 68.835 ;
        RECT 135.365 68.635 136.315 68.835 ;
        RECT 133.105 68.155 136.315 68.635 ;
        RECT 133.250 67.955 136.315 68.155 ;
        RECT 108.410 67.715 108.580 67.905 ;
        RECT 110.700 67.715 110.870 67.905 ;
        RECT 111.165 67.715 111.335 67.905 ;
        RECT 112.085 67.735 112.255 67.905 ;
        RECT 112.540 67.765 112.660 67.875 ;
        RECT 113.470 67.735 113.640 67.925 ;
        RECT 113.920 67.715 114.090 67.905 ;
        RECT 115.300 67.715 115.470 67.905 ;
        RECT 115.765 67.715 115.935 67.925 ;
        RECT 118.085 67.905 118.235 67.925 ;
        RECT 117.600 67.765 117.720 67.875 ;
        RECT 118.065 67.735 118.235 67.905 ;
        RECT 118.520 67.765 118.640 67.875 ;
        RECT 119.900 67.715 120.070 67.905 ;
        RECT 120.365 67.735 120.535 67.925 ;
        RECT 121.280 67.715 121.450 67.905 ;
        RECT 121.745 67.715 121.915 67.905 ;
        RECT 122.200 67.765 122.320 67.875 ;
        RECT 122.670 67.735 122.840 67.925 ;
        RECT 124.040 67.715 124.210 67.905 ;
        RECT 124.505 67.715 124.675 67.925 ;
        RECT 126.345 67.715 126.515 67.905 ;
        RECT 128.190 67.735 128.360 67.925 ;
        RECT 129.100 67.765 129.220 67.875 ;
        RECT 130.480 67.715 130.650 67.905 ;
        RECT 131.400 67.735 131.570 67.925 ;
        RECT 131.870 67.905 132.040 67.925 ;
        RECT 131.860 67.735 132.040 67.905 ;
        RECT 132.335 67.760 132.495 67.870 ;
        RECT 131.860 67.715 132.030 67.735 ;
        RECT 99.020 67.685 99.975 67.715 ;
        RECT 97.695 67.005 99.975 67.685 ;
        RECT 99.020 66.805 99.975 67.005 ;
        RECT 99.995 66.845 100.425 67.630 ;
        RECT 100.445 66.935 101.815 67.715 ;
        RECT 101.825 66.935 103.195 67.715 ;
        RECT 103.205 66.905 106.875 67.715 ;
        RECT 106.885 66.905 108.255 67.715 ;
        RECT 108.265 66.805 109.615 67.715 ;
        RECT 109.665 66.805 111.015 67.715 ;
        RECT 111.025 66.905 112.855 67.715 ;
        RECT 112.885 66.805 114.235 67.715 ;
        RECT 114.265 66.805 115.615 67.715 ;
        RECT 115.625 66.905 118.375 67.715 ;
        RECT 118.865 66.805 120.215 67.715 ;
        RECT 120.245 66.805 121.595 67.715 ;
        RECT 121.605 66.905 122.975 67.715 ;
        RECT 123.005 66.805 124.355 67.715 ;
        RECT 124.365 66.905 125.735 67.715 ;
        RECT 125.755 66.845 126.185 67.630 ;
        RECT 126.205 66.905 128.955 67.715 ;
        RECT 129.445 66.805 130.795 67.715 ;
        RECT 130.825 66.805 132.175 67.715 ;
        RECT 133.250 67.685 133.420 67.955 ;
        RECT 135.380 67.925 136.315 67.955 ;
        RECT 137.245 67.925 138.615 68.705 ;
        RECT 138.635 68.010 139.065 68.795 ;
        RECT 140.420 68.635 141.375 68.835 ;
        RECT 142.720 68.635 143.675 68.835 ;
        RECT 139.095 67.955 141.375 68.635 ;
        RECT 141.395 67.955 143.675 68.635 ;
        RECT 136.465 67.715 136.635 67.905 ;
        RECT 137.385 67.735 137.555 67.925 ;
        RECT 139.220 67.905 139.390 67.955 ;
        RECT 140.420 67.925 141.375 67.955 ;
        RECT 137.845 67.715 138.015 67.905 ;
        RECT 139.220 67.735 139.395 67.905 ;
        RECT 141.520 67.735 141.690 67.955 ;
        RECT 142.720 67.925 143.675 67.955 ;
        RECT 143.685 67.925 145.055 68.705 ;
        RECT 145.065 67.925 146.435 68.705 ;
        RECT 146.445 67.925 151.955 68.735 ;
        RECT 151.965 67.925 155.635 68.735 ;
        RECT 155.645 67.925 157.015 68.735 ;
        RECT 139.225 67.715 139.395 67.735 ;
        RECT 144.745 67.715 144.915 67.925 ;
        RECT 145.205 67.735 145.375 67.925 ;
        RECT 146.585 67.735 146.755 67.925 ;
        RECT 150.265 67.715 150.435 67.905 ;
        RECT 152.105 67.715 152.275 67.925 ;
        RECT 156.705 67.715 156.875 67.925 ;
        RECT 135.380 67.685 136.315 67.715 ;
        RECT 133.250 67.485 136.315 67.685 ;
        RECT 133.105 67.005 136.315 67.485 ;
        RECT 133.105 66.805 134.035 67.005 ;
        RECT 135.365 66.805 136.315 67.005 ;
        RECT 136.325 66.905 137.695 67.715 ;
        RECT 137.705 66.935 139.075 67.715 ;
        RECT 139.085 66.905 144.595 67.715 ;
        RECT 144.605 66.905 150.115 67.715 ;
        RECT 150.125 66.905 151.495 67.715 ;
        RECT 151.515 66.845 151.945 67.630 ;
        RECT 151.965 66.905 155.635 67.715 ;
        RECT 155.645 66.905 157.015 67.715 ;
      LAYER nwell ;
        RECT 22.510 63.685 157.210 66.515 ;
      LAYER pwell ;
        RECT 22.705 62.485 24.075 63.295 ;
        RECT 28.730 63.165 30.515 63.395 ;
        RECT 24.545 62.485 30.515 63.165 ;
        RECT 31.905 62.485 33.735 63.295 ;
        RECT 33.745 62.485 35.095 63.395 ;
        RECT 35.595 62.570 36.025 63.355 ;
        RECT 36.065 62.485 37.415 63.395 ;
        RECT 37.445 62.485 38.795 63.395 ;
        RECT 38.805 62.485 40.175 63.295 ;
        RECT 41.565 62.485 42.915 63.395 ;
        RECT 42.965 62.485 44.315 63.395 ;
        RECT 49.430 63.165 51.215 63.395 ;
        RECT 55.410 63.165 57.195 63.395 ;
        RECT 45.245 62.485 51.215 63.165 ;
        RECT 51.225 62.485 57.195 63.165 ;
        RECT 58.585 62.485 61.335 63.295 ;
        RECT 61.355 62.570 61.785 63.355 ;
        RECT 61.805 62.485 64.555 63.295 ;
        RECT 69.210 63.165 70.995 63.395 ;
        RECT 65.025 62.485 70.995 63.165 ;
        RECT 71.005 62.485 72.835 63.295 ;
        RECT 82.090 63.165 83.875 63.395 ;
        RECT 77.905 62.485 83.875 63.165 ;
        RECT 83.885 62.485 85.235 63.395 ;
        RECT 85.265 62.485 86.615 63.395 ;
        RECT 87.115 62.570 87.545 63.355 ;
        RECT 88.945 62.485 90.315 63.295 ;
        RECT 94.005 62.485 95.835 63.295 ;
        RECT 100.030 63.165 101.815 63.395 ;
        RECT 95.845 62.485 101.815 63.165 ;
        RECT 104.585 62.485 106.415 63.295 ;
        RECT 109.645 62.485 112.395 63.295 ;
        RECT 112.875 62.570 113.305 63.355 ;
        RECT 121.650 63.165 123.435 63.395 ;
        RECT 117.465 62.485 123.435 63.165 ;
        RECT 124.385 62.485 125.735 63.395 ;
        RECT 129.930 63.165 131.715 63.395 ;
        RECT 125.745 62.485 131.715 63.165 ;
        RECT 135.865 62.485 137.235 63.295 ;
        RECT 138.635 62.570 139.065 63.355 ;
        RECT 143.730 63.165 145.515 63.395 ;
        RECT 139.545 62.485 145.515 63.165 ;
        RECT 148.285 62.485 153.795 63.295 ;
        RECT 153.805 62.485 155.635 63.295 ;
        RECT 155.645 62.485 157.015 63.295 ;
        RECT 22.845 62.275 23.015 62.485 ;
        RECT 24.220 62.325 24.340 62.435 ;
        RECT 24.690 62.275 24.860 62.485 ;
        RECT 31.585 62.295 31.755 62.465 ;
        RECT 32.045 62.295 32.215 62.485 ;
        RECT 33.890 62.295 34.060 62.485 ;
        RECT 35.260 62.325 35.380 62.435 ;
        RECT 36.180 62.275 36.350 62.465 ;
        RECT 36.650 62.275 36.820 62.465 ;
        RECT 37.100 62.295 37.270 62.485 ;
        RECT 38.480 62.295 38.650 62.485 ;
        RECT 38.945 62.295 39.115 62.485 ;
        RECT 40.325 62.295 40.495 62.465 ;
        RECT 41.710 62.295 41.880 62.485 ;
        RECT 42.630 62.275 42.800 62.465 ;
        RECT 44.000 62.295 44.170 62.485 ;
        RECT 44.475 62.330 44.635 62.440 ;
        RECT 45.390 62.295 45.560 62.485 ;
        RECT 51.370 62.465 51.540 62.485 ;
        RECT 49.065 62.295 49.235 62.465 ;
        RECT 51.365 62.295 51.540 62.465 ;
        RECT 51.820 62.325 51.940 62.435 ;
        RECT 52.285 62.295 52.455 62.465 ;
        RECT 53.670 62.275 53.840 62.465 ;
        RECT 58.265 62.295 58.435 62.465 ;
        RECT 58.725 62.295 58.895 62.485 ;
        RECT 59.650 62.275 59.820 62.465 ;
        RECT 61.945 62.295 62.115 62.485 ;
        RECT 64.700 62.325 64.820 62.435 ;
        RECT 65.170 62.295 65.340 62.485 ;
        RECT 65.625 62.295 65.795 62.465 ;
        RECT 67.005 62.295 67.175 62.465 ;
        RECT 68.390 62.275 68.560 62.465 ;
        RECT 71.145 62.295 71.315 62.485 ;
        RECT 72.980 62.325 73.100 62.435 ;
        RECT 73.445 62.295 73.615 62.465 ;
        RECT 74.830 62.435 75.000 62.465 ;
        RECT 74.820 62.325 75.000 62.435 ;
        RECT 74.830 62.275 75.000 62.325 ;
        RECT 76.205 62.295 76.375 62.465 ;
        RECT 76.665 62.295 76.835 62.465 ;
        RECT 78.050 62.295 78.220 62.485 ;
        RECT 84.030 62.295 84.200 62.485 ;
        RECT 85.410 62.295 85.580 62.485 ;
        RECT 86.320 62.275 86.490 62.465 ;
        RECT 86.790 62.435 86.960 62.465 ;
        RECT 86.780 62.325 86.960 62.435 ;
        RECT 86.790 62.275 86.960 62.325 ;
        RECT 88.625 62.295 88.795 62.465 ;
        RECT 89.085 62.295 89.255 62.485 ;
        RECT 91.385 62.295 91.555 62.465 ;
        RECT 91.855 62.330 92.015 62.440 ;
        RECT 92.770 62.275 92.940 62.465 ;
        RECT 93.685 62.295 93.855 62.465 ;
        RECT 94.145 62.295 94.315 62.485 ;
        RECT 95.990 62.295 96.160 62.485 ;
        RECT 98.745 62.295 98.915 62.465 ;
        RECT 100.590 62.275 100.760 62.465 ;
        RECT 102.885 62.295 103.055 62.465 ;
        RECT 103.345 62.295 103.515 62.465 ;
        RECT 104.725 62.295 104.895 62.485 ;
        RECT 106.570 62.435 106.740 62.465 ;
        RECT 106.560 62.325 106.740 62.435 ;
        RECT 106.570 62.275 106.740 62.325 ;
        RECT 107.945 62.295 108.115 62.465 ;
        RECT 108.405 62.295 108.575 62.465 ;
        RECT 109.785 62.295 109.955 62.485 ;
        RECT 112.550 62.435 112.720 62.465 ;
        RECT 112.540 62.325 112.720 62.435 ;
        RECT 112.550 62.275 112.720 62.325 ;
        RECT 114.385 62.295 114.555 62.465 ;
        RECT 114.845 62.295 115.015 62.465 ;
        RECT 116.225 62.295 116.395 62.465 ;
        RECT 117.610 62.295 117.780 62.485 ;
        RECT 125.420 62.465 125.590 62.485 ;
        RECT 118.530 62.275 118.700 62.465 ;
        RECT 123.595 62.330 123.755 62.440 ;
        RECT 125.420 62.295 125.595 62.465 ;
        RECT 125.890 62.295 126.060 62.485 ;
        RECT 126.350 62.275 126.520 62.465 ;
        RECT 132.330 62.275 132.500 62.465 ;
        RECT 132.785 62.295 132.955 62.465 ;
        RECT 134.165 62.295 134.335 62.465 ;
        RECT 134.625 62.295 134.795 62.465 ;
        RECT 136.005 62.295 136.175 62.485 ;
        RECT 137.385 62.295 137.555 62.465 ;
        RECT 138.310 62.275 138.480 62.465 ;
        RECT 139.220 62.325 139.340 62.435 ;
        RECT 139.690 62.295 139.860 62.485 ;
        RECT 144.290 62.275 144.460 62.465 ;
        RECT 146.585 62.295 146.755 62.465 ;
        RECT 147.965 62.295 148.135 62.465 ;
        RECT 148.425 62.295 148.595 62.485 ;
        RECT 150.265 62.275 150.435 62.465 ;
        RECT 152.105 62.275 152.275 62.465 ;
        RECT 153.945 62.295 154.115 62.485 ;
        RECT 156.705 62.275 156.875 62.485 ;
        RECT 22.705 61.465 24.075 62.275 ;
        RECT 24.545 61.595 30.515 62.275 ;
        RECT 28.730 61.365 30.515 61.595 ;
        RECT 30.525 61.595 36.495 62.275 ;
        RECT 36.505 61.595 42.475 62.275 ;
        RECT 42.485 61.595 48.455 62.275 ;
        RECT 30.525 61.365 32.310 61.595 ;
        RECT 40.690 61.365 42.475 61.595 ;
        RECT 46.670 61.365 48.455 61.595 ;
        RECT 48.475 61.405 48.905 62.190 ;
        RECT 53.525 61.595 59.495 62.275 ;
        RECT 59.505 61.595 65.475 62.275 ;
        RECT 68.245 61.595 74.215 62.275 ;
        RECT 57.710 61.365 59.495 61.595 ;
        RECT 63.690 61.365 65.475 61.595 ;
        RECT 72.430 61.365 74.215 61.595 ;
        RECT 74.235 61.405 74.665 62.190 ;
        RECT 74.685 61.595 80.655 62.275 ;
        RECT 78.870 61.365 80.655 61.595 ;
        RECT 80.665 61.595 86.635 62.275 ;
        RECT 86.645 61.595 92.615 62.275 ;
        RECT 92.625 61.595 98.595 62.275 ;
        RECT 80.665 61.365 82.450 61.595 ;
        RECT 90.830 61.365 92.615 61.595 ;
        RECT 96.810 61.365 98.595 61.595 ;
        RECT 99.995 61.405 100.425 62.190 ;
        RECT 100.445 61.595 106.415 62.275 ;
        RECT 106.425 61.595 112.395 62.275 ;
        RECT 112.405 61.595 118.375 62.275 ;
        RECT 118.385 61.595 124.355 62.275 ;
        RECT 104.630 61.365 106.415 61.595 ;
        RECT 110.610 61.365 112.395 61.595 ;
        RECT 116.590 61.365 118.375 61.595 ;
        RECT 122.570 61.365 124.355 61.595 ;
        RECT 125.755 61.405 126.185 62.190 ;
        RECT 126.205 61.595 132.175 62.275 ;
        RECT 132.185 61.595 138.155 62.275 ;
        RECT 138.165 61.595 144.135 62.275 ;
        RECT 144.145 61.595 150.115 62.275 ;
        RECT 130.390 61.365 132.175 61.595 ;
        RECT 136.370 61.365 138.155 61.595 ;
        RECT 142.350 61.365 144.135 61.595 ;
        RECT 148.330 61.365 150.115 61.595 ;
        RECT 150.125 61.465 151.495 62.275 ;
        RECT 151.515 61.405 151.945 62.190 ;
        RECT 151.965 61.465 155.635 62.275 ;
        RECT 155.645 61.465 157.015 62.275 ;
      LAYER nwell ;
        RECT 22.510 58.245 157.210 61.075 ;
      LAYER pwell ;
        RECT 22.705 57.045 24.075 57.855 ;
        RECT 28.225 57.045 29.595 57.855 ;
        RECT 33.790 57.725 35.575 57.955 ;
        RECT 29.605 57.045 35.575 57.725 ;
        RECT 35.595 57.130 36.025 57.915 ;
        RECT 39.725 57.045 41.095 57.855 ;
        RECT 45.290 57.725 47.075 57.955 ;
        RECT 41.105 57.045 47.075 57.725 ;
        RECT 48.475 57.130 48.905 57.915 ;
        RECT 48.925 57.045 52.595 57.855 ;
        RECT 57.710 57.725 59.495 57.955 ;
        RECT 53.525 57.045 59.495 57.725 ;
        RECT 61.355 57.130 61.785 57.915 ;
        RECT 61.805 57.045 64.555 57.855 ;
        RECT 71.050 57.725 72.835 57.955 ;
        RECT 66.865 57.045 72.835 57.725 ;
        RECT 72.845 57.045 74.215 57.855 ;
        RECT 74.235 57.130 74.665 57.915 ;
        RECT 78.870 57.725 80.655 57.955 ;
        RECT 85.310 57.725 87.095 57.955 ;
        RECT 74.685 57.045 80.655 57.725 ;
        RECT 81.125 57.045 87.095 57.725 ;
        RECT 87.115 57.130 87.545 57.915 ;
        RECT 94.050 57.725 95.835 57.955 ;
        RECT 89.865 57.045 95.835 57.725 ;
        RECT 95.845 57.045 99.515 57.855 ;
        RECT 99.995 57.130 100.425 57.915 ;
        RECT 105.090 57.725 106.875 57.955 ;
        RECT 111.070 57.725 112.855 57.955 ;
        RECT 100.905 57.045 106.875 57.725 ;
        RECT 106.885 57.045 112.855 57.725 ;
        RECT 112.875 57.130 113.305 57.915 ;
        RECT 117.510 57.725 119.295 57.955 ;
        RECT 123.950 57.725 125.735 57.955 ;
        RECT 113.325 57.045 119.295 57.725 ;
        RECT 119.765 57.045 125.735 57.725 ;
        RECT 125.755 57.130 126.185 57.915 ;
        RECT 128.965 57.045 130.795 57.855 ;
        RECT 134.990 57.725 136.775 57.955 ;
        RECT 130.805 57.045 136.775 57.725 ;
        RECT 138.635 57.130 139.065 57.915 ;
        RECT 143.270 57.725 145.055 57.955 ;
        RECT 149.250 57.725 151.035 57.955 ;
        RECT 139.085 57.045 145.055 57.725 ;
        RECT 145.065 57.045 151.035 57.725 ;
        RECT 151.515 57.130 151.945 57.915 ;
        RECT 151.965 57.045 155.635 57.855 ;
        RECT 155.645 57.045 157.015 57.855 ;
        RECT 22.845 56.855 23.015 57.045 ;
        RECT 24.235 56.890 24.395 57.000 ;
        RECT 26.065 56.855 26.235 57.025 ;
        RECT 26.520 56.885 26.640 56.995 ;
        RECT 27.905 56.855 28.075 57.025 ;
        RECT 28.365 56.855 28.535 57.045 ;
        RECT 29.750 56.855 29.920 57.045 ;
        RECT 36.195 56.890 36.355 57.000 ;
        RECT 38.025 56.855 38.195 57.025 ;
        RECT 39.405 56.855 39.575 57.025 ;
        RECT 39.865 56.855 40.035 57.045 ;
        RECT 41.250 56.855 41.420 57.045 ;
        RECT 48.145 56.855 48.315 57.025 ;
        RECT 49.065 56.855 49.235 57.045 ;
        RECT 52.755 56.890 52.915 57.000 ;
        RECT 53.670 56.855 53.840 57.045 ;
        RECT 60.565 56.855 60.735 57.025 ;
        RECT 61.020 56.885 61.140 56.995 ;
        RECT 61.945 56.855 62.115 57.045 ;
        RECT 64.700 56.885 64.820 56.995 ;
        RECT 66.085 56.855 66.255 57.025 ;
        RECT 66.540 56.885 66.660 56.995 ;
        RECT 67.010 56.855 67.180 57.045 ;
        RECT 72.985 56.855 73.155 57.045 ;
        RECT 74.830 56.855 75.000 57.045 ;
        RECT 80.800 56.885 80.920 56.995 ;
        RECT 81.270 56.855 81.440 57.045 ;
        RECT 87.700 56.885 87.820 56.995 ;
        RECT 89.085 56.855 89.255 57.025 ;
        RECT 89.540 56.885 89.660 56.995 ;
        RECT 90.010 56.855 90.180 57.045 ;
        RECT 95.985 56.855 96.155 57.045 ;
        RECT 99.660 56.885 99.780 56.995 ;
        RECT 100.580 56.885 100.700 56.995 ;
        RECT 101.050 56.855 101.220 57.045 ;
        RECT 107.030 56.855 107.200 57.045 ;
        RECT 113.470 56.855 113.640 57.045 ;
        RECT 119.440 56.885 119.560 56.995 ;
        RECT 119.910 56.855 120.080 57.045 ;
        RECT 127.265 56.855 127.435 57.025 ;
        RECT 128.645 56.855 128.815 57.025 ;
        RECT 129.105 56.855 129.275 57.045 ;
        RECT 130.950 56.855 131.120 57.045 ;
        RECT 136.920 56.885 137.040 56.995 ;
        RECT 137.385 56.855 137.555 57.025 ;
        RECT 139.230 56.855 139.400 57.045 ;
        RECT 145.210 56.855 145.380 57.045 ;
        RECT 151.180 56.885 151.300 56.995 ;
        RECT 152.105 56.855 152.275 57.045 ;
        RECT 156.705 56.855 156.875 57.045 ;
        RECT 32.820 33.660 35.780 47.760 ;
        RECT 39.820 37.910 42.780 38.760 ;
        RECT 43.520 37.910 46.480 38.310 ;
        RECT 39.820 36.460 46.480 37.910 ;
        RECT 39.820 33.660 42.780 36.460 ;
        RECT 43.520 34.090 46.480 36.460 ;
        RECT 32.980 29.260 33.280 29.860 ;
        RECT 34.820 22.680 37.780 33.260 ;
        RECT 46.530 32.150 50.130 35.110 ;
        RECT 50.230 28.700 53.330 35.110 ;
        RECT 74.040 34.500 77.000 48.600 ;
        RECT 81.040 38.750 84.000 39.600 ;
        RECT 84.740 38.750 87.700 39.150 ;
        RECT 81.040 37.300 87.700 38.750 ;
        RECT 81.040 34.500 84.000 37.300 ;
        RECT 84.740 34.930 87.700 37.300 ;
        RECT 74.200 30.100 74.500 30.700 ;
        RECT 49.800 25.310 53.880 28.410 ;
        RECT 50.350 24.860 53.420 25.310 ;
        RECT 36.320 14.160 39.280 22.260 ;
        RECT 49.970 21.760 54.930 24.860 ;
        RECT 76.040 23.520 79.000 34.100 ;
        RECT 87.750 32.990 91.350 35.950 ;
        RECT 91.450 29.540 94.550 35.950 ;
        RECT 113.920 35.900 116.880 50.000 ;
        RECT 120.920 40.150 123.880 41.000 ;
        RECT 124.620 40.150 127.580 40.550 ;
        RECT 120.920 38.700 127.580 40.150 ;
        RECT 120.920 35.900 123.880 38.700 ;
        RECT 124.620 36.330 127.580 38.700 ;
        RECT 114.080 31.500 114.380 32.100 ;
        RECT 91.020 26.150 95.100 29.250 ;
        RECT 91.570 25.700 94.640 26.150 ;
        RECT 50.350 21.280 53.420 21.760 ;
        RECT 49.940 18.180 56.140 21.280 ;
        RECT 50.350 17.700 53.420 18.180 ;
        RECT 49.810 14.600 57.770 17.700 ;
        RECT 77.540 15.000 80.500 23.100 ;
        RECT 91.190 22.600 96.150 25.700 ;
        RECT 115.920 24.920 118.880 35.500 ;
        RECT 127.630 34.390 131.230 37.350 ;
        RECT 131.330 30.940 134.430 37.350 ;
        RECT 130.900 27.550 134.980 30.650 ;
        RECT 131.450 27.100 134.520 27.550 ;
        RECT 91.570 22.120 94.640 22.600 ;
        RECT 91.160 19.020 97.360 22.120 ;
        RECT 91.570 18.540 94.640 19.020 ;
        RECT 91.030 15.440 98.990 18.540 ;
        RECT 117.420 16.400 120.380 24.500 ;
        RECT 131.070 24.000 136.030 27.100 ;
        RECT 131.450 23.520 134.520 24.000 ;
        RECT 131.040 20.420 137.240 23.520 ;
        RECT 131.450 19.940 134.520 20.420 ;
        RECT 130.910 16.840 138.870 19.940 ;
        RECT 131.450 16.360 134.520 16.840 ;
        RECT 91.570 14.960 94.640 15.440 ;
        RECT 50.350 14.120 53.420 14.600 ;
        RECT 38.320 7.420 41.280 13.760 ;
        RECT 49.830 11.020 60.270 14.120 ;
        RECT 50.350 10.540 53.420 11.020 ;
        RECT 49.840 7.440 63.800 10.540 ;
        RECT 79.540 8.260 82.500 14.600 ;
        RECT 91.050 11.860 101.490 14.960 ;
        RECT 91.570 11.380 94.640 11.860 ;
        RECT 91.060 8.280 105.020 11.380 ;
        RECT 119.420 9.660 122.380 16.000 ;
        RECT 130.930 13.260 141.370 16.360 ;
        RECT 131.450 12.780 134.520 13.260 ;
        RECT 130.940 9.680 144.900 12.780 ;
      LAYER li1 ;
        RECT 22.700 209.175 157.020 209.345 ;
        RECT 22.785 208.425 23.995 209.175 ;
        RECT 24.165 208.630 29.510 209.175 ;
        RECT 29.685 208.630 35.030 209.175 ;
        RECT 22.785 207.885 23.305 208.425 ;
        RECT 23.475 207.715 23.995 208.255 ;
        RECT 25.750 207.800 26.090 208.630 ;
        RECT 22.785 206.625 23.995 207.715 ;
        RECT 27.570 207.060 27.920 208.310 ;
        RECT 31.270 207.800 31.610 208.630 ;
        RECT 35.665 208.450 35.955 209.175 ;
        RECT 36.125 208.630 41.470 209.175 ;
        RECT 41.645 208.630 46.990 209.175 ;
        RECT 33.090 207.060 33.440 208.310 ;
        RECT 37.710 207.800 38.050 208.630 ;
        RECT 24.165 206.625 29.510 207.060 ;
        RECT 29.685 206.625 35.030 207.060 ;
        RECT 35.665 206.625 35.955 207.790 ;
        RECT 39.530 207.060 39.880 208.310 ;
        RECT 43.230 207.800 43.570 208.630 ;
        RECT 47.165 208.425 48.375 209.175 ;
        RECT 48.545 208.450 48.835 209.175 ;
        RECT 49.030 208.525 49.340 208.995 ;
        RECT 49.510 208.695 50.245 209.175 ;
        RECT 50.415 208.605 50.585 208.955 ;
        RECT 50.755 208.775 51.135 209.175 ;
        RECT 45.050 207.060 45.400 208.310 ;
        RECT 47.165 207.885 47.685 208.425 ;
        RECT 49.030 208.355 49.765 208.525 ;
        RECT 50.415 208.435 51.155 208.605 ;
        RECT 51.325 208.500 51.595 208.845 ;
        RECT 49.515 208.265 49.765 208.355 ;
        RECT 50.985 208.265 51.155 208.435 ;
        RECT 47.855 207.715 48.375 208.255 ;
        RECT 49.010 207.935 49.345 208.185 ;
        RECT 49.515 207.935 50.255 208.265 ;
        RECT 50.985 207.935 51.215 208.265 ;
        RECT 36.125 206.625 41.470 207.060 ;
        RECT 41.645 206.625 46.990 207.060 ;
        RECT 47.165 206.625 48.375 207.715 ;
        RECT 48.545 206.625 48.835 207.790 ;
        RECT 49.010 206.625 49.265 207.765 ;
        RECT 49.515 207.375 49.685 207.935 ;
        RECT 50.985 207.765 51.155 207.935 ;
        RECT 51.425 207.765 51.595 208.500 ;
        RECT 51.765 208.375 52.075 209.175 ;
        RECT 52.280 208.375 52.975 209.005 ;
        RECT 53.145 208.435 53.465 208.915 ;
        RECT 53.635 208.605 53.865 209.005 ;
        RECT 54.035 208.785 54.385 209.175 ;
        RECT 53.635 208.525 54.145 208.605 ;
        RECT 54.555 208.525 54.885 209.005 ;
        RECT 53.635 208.435 54.885 208.525 ;
        RECT 51.775 207.935 52.110 208.205 ;
        RECT 52.280 207.775 52.450 208.375 ;
        RECT 52.620 207.935 52.955 208.185 ;
        RECT 49.910 207.595 51.155 207.765 ;
        RECT 49.910 207.345 50.330 207.595 ;
        RECT 49.460 206.845 50.655 207.175 ;
        RECT 50.835 206.625 51.115 207.425 ;
        RECT 51.325 206.795 51.595 207.765 ;
        RECT 51.765 206.625 52.045 207.765 ;
        RECT 52.215 206.795 52.545 207.775 ;
        RECT 52.715 206.625 52.975 207.765 ;
        RECT 53.145 207.505 53.315 208.435 ;
        RECT 53.975 208.355 54.885 208.435 ;
        RECT 55.055 208.355 55.225 209.175 ;
        RECT 55.730 208.435 56.195 208.980 ;
        RECT 53.485 207.845 53.655 208.265 ;
        RECT 53.885 208.015 54.485 208.185 ;
        RECT 53.485 207.675 54.145 207.845 ;
        RECT 53.145 207.305 53.805 207.505 ;
        RECT 53.975 207.475 54.145 207.675 ;
        RECT 54.315 207.815 54.485 208.015 ;
        RECT 54.655 207.985 55.350 208.185 ;
        RECT 55.610 207.815 55.855 208.265 ;
        RECT 54.315 207.645 55.855 207.815 ;
        RECT 56.025 207.475 56.195 208.435 ;
        RECT 53.975 207.305 56.195 207.475 ;
        RECT 57.285 208.435 57.670 209.005 ;
        RECT 57.840 208.715 58.165 209.175 ;
        RECT 58.685 208.545 58.965 209.005 ;
        RECT 57.285 207.765 57.565 208.435 ;
        RECT 57.840 208.375 58.965 208.545 ;
        RECT 57.840 208.265 58.290 208.375 ;
        RECT 57.735 207.935 58.290 208.265 ;
        RECT 59.155 208.205 59.555 209.005 ;
        RECT 59.955 208.715 60.225 209.175 ;
        RECT 60.395 208.545 60.680 209.005 ;
        RECT 53.635 207.135 53.805 207.305 ;
        RECT 53.165 206.625 53.465 207.135 ;
        RECT 53.635 206.965 54.015 207.135 ;
        RECT 54.595 206.625 55.225 207.135 ;
        RECT 55.395 206.795 55.725 207.305 ;
        RECT 55.895 206.625 56.195 207.135 ;
        RECT 57.285 206.795 57.670 207.765 ;
        RECT 57.840 207.475 58.290 207.935 ;
        RECT 58.460 207.645 59.555 208.205 ;
        RECT 57.840 207.255 58.965 207.475 ;
        RECT 57.840 206.625 58.165 207.085 ;
        RECT 58.685 206.795 58.965 207.255 ;
        RECT 59.155 206.795 59.555 207.645 ;
        RECT 59.725 208.375 60.680 208.545 ;
        RECT 61.425 208.450 61.715 209.175 ;
        RECT 61.885 208.500 62.145 209.005 ;
        RECT 62.325 208.795 62.655 209.175 ;
        RECT 62.835 208.625 63.005 209.005 ;
        RECT 59.725 207.475 59.935 208.375 ;
        RECT 60.105 207.645 60.795 208.205 ;
        RECT 59.725 207.255 60.680 207.475 ;
        RECT 59.955 206.625 60.225 207.085 ;
        RECT 60.395 206.795 60.680 207.255 ;
        RECT 61.425 206.625 61.715 207.790 ;
        RECT 61.885 207.700 62.055 208.500 ;
        RECT 62.340 208.455 63.005 208.625 ;
        RECT 64.275 208.625 64.445 209.005 ;
        RECT 64.625 208.795 64.955 209.175 ;
        RECT 64.275 208.455 64.940 208.625 ;
        RECT 65.135 208.500 65.395 209.005 ;
        RECT 62.340 208.200 62.510 208.455 ;
        RECT 62.225 207.870 62.510 208.200 ;
        RECT 62.745 207.905 63.075 208.275 ;
        RECT 64.205 207.905 64.535 208.275 ;
        RECT 64.770 208.200 64.940 208.455 ;
        RECT 62.340 207.725 62.510 207.870 ;
        RECT 64.770 207.870 65.055 208.200 ;
        RECT 64.770 207.725 64.940 207.870 ;
        RECT 61.885 206.795 62.155 207.700 ;
        RECT 62.340 207.555 63.005 207.725 ;
        RECT 62.325 206.625 62.655 207.385 ;
        RECT 62.835 206.795 63.005 207.555 ;
        RECT 64.275 207.555 64.940 207.725 ;
        RECT 65.225 207.700 65.395 208.500 ;
        RECT 65.565 208.405 69.075 209.175 ;
        RECT 69.705 208.525 69.965 209.005 ;
        RECT 70.135 208.635 70.385 209.175 ;
        RECT 65.565 207.885 67.215 208.405 ;
        RECT 67.385 207.715 69.075 208.235 ;
        RECT 64.275 206.795 64.445 207.555 ;
        RECT 64.625 206.625 64.955 207.385 ;
        RECT 65.125 206.795 65.395 207.700 ;
        RECT 65.565 206.625 69.075 207.715 ;
        RECT 69.705 207.495 69.875 208.525 ;
        RECT 70.555 208.470 70.775 208.955 ;
        RECT 70.045 207.875 70.275 208.270 ;
        RECT 70.445 208.045 70.775 208.470 ;
        RECT 70.945 208.795 71.835 208.965 ;
        RECT 70.945 208.070 71.115 208.795 ;
        RECT 72.095 208.625 72.265 209.005 ;
        RECT 72.445 208.795 72.775 209.175 ;
        RECT 71.285 208.240 71.835 208.625 ;
        RECT 72.095 208.455 72.760 208.625 ;
        RECT 72.955 208.500 73.215 209.005 ;
        RECT 70.945 208.000 71.835 208.070 ;
        RECT 70.940 207.975 71.835 208.000 ;
        RECT 70.930 207.960 71.835 207.975 ;
        RECT 70.925 207.945 71.835 207.960 ;
        RECT 70.915 207.940 71.835 207.945 ;
        RECT 70.910 207.930 71.835 207.940 ;
        RECT 70.905 207.920 71.835 207.930 ;
        RECT 70.895 207.915 71.835 207.920 ;
        RECT 70.885 207.905 71.835 207.915 ;
        RECT 72.025 207.905 72.355 208.275 ;
        RECT 72.590 208.200 72.760 208.455 ;
        RECT 70.875 207.900 71.835 207.905 ;
        RECT 70.875 207.895 71.210 207.900 ;
        RECT 70.860 207.890 71.210 207.895 ;
        RECT 70.845 207.880 71.210 207.890 ;
        RECT 70.820 207.875 71.210 207.880 ;
        RECT 70.045 207.870 71.210 207.875 ;
        RECT 70.045 207.835 71.180 207.870 ;
        RECT 70.045 207.810 71.145 207.835 ;
        RECT 70.045 207.780 71.115 207.810 ;
        RECT 70.045 207.750 71.095 207.780 ;
        RECT 70.045 207.720 71.075 207.750 ;
        RECT 70.045 207.710 71.005 207.720 ;
        RECT 70.045 207.700 70.980 207.710 ;
        RECT 70.045 207.685 70.960 207.700 ;
        RECT 70.045 207.670 70.940 207.685 ;
        RECT 70.150 207.660 70.935 207.670 ;
        RECT 70.150 207.625 70.920 207.660 ;
        RECT 69.705 206.795 69.980 207.495 ;
        RECT 70.150 207.375 70.905 207.625 ;
        RECT 71.075 207.305 71.405 207.550 ;
        RECT 71.575 207.450 71.835 207.900 ;
        RECT 72.590 207.870 72.875 208.200 ;
        RECT 72.590 207.725 72.760 207.870 ;
        RECT 72.095 207.555 72.760 207.725 ;
        RECT 73.045 207.700 73.215 208.500 ;
        RECT 74.305 208.450 74.595 209.175 ;
        RECT 74.765 208.405 78.275 209.175 ;
        RECT 78.995 208.625 79.165 209.005 ;
        RECT 79.380 208.795 79.710 209.175 ;
        RECT 78.995 208.455 79.710 208.625 ;
        RECT 74.765 207.885 76.415 208.405 ;
        RECT 71.220 207.280 71.405 207.305 ;
        RECT 71.220 207.180 71.835 207.280 ;
        RECT 70.150 206.625 70.405 207.170 ;
        RECT 70.575 206.795 71.055 207.135 ;
        RECT 71.230 206.625 71.835 207.180 ;
        RECT 72.095 206.795 72.265 207.555 ;
        RECT 72.445 206.625 72.775 207.385 ;
        RECT 72.945 206.795 73.215 207.700 ;
        RECT 74.305 206.625 74.595 207.790 ;
        RECT 76.585 207.715 78.275 208.235 ;
        RECT 78.905 207.905 79.260 208.275 ;
        RECT 79.540 208.265 79.710 208.455 ;
        RECT 79.880 208.430 80.135 209.005 ;
        RECT 79.540 207.935 79.795 208.265 ;
        RECT 79.540 207.725 79.710 207.935 ;
        RECT 74.765 206.625 78.275 207.715 ;
        RECT 78.995 207.555 79.710 207.725 ;
        RECT 79.965 207.700 80.135 208.430 ;
        RECT 80.310 208.335 80.570 209.175 ;
        RECT 80.745 208.375 81.055 209.175 ;
        RECT 81.260 208.375 81.955 209.005 ;
        RECT 82.585 208.435 82.970 209.005 ;
        RECT 83.140 208.715 83.465 209.175 ;
        RECT 83.985 208.545 84.265 209.005 ;
        RECT 80.755 207.935 81.090 208.205 ;
        RECT 81.260 207.775 81.430 208.375 ;
        RECT 81.600 207.935 81.935 208.185 ;
        RECT 78.995 206.795 79.165 207.555 ;
        RECT 79.380 206.625 79.710 207.385 ;
        RECT 79.880 206.795 80.135 207.700 ;
        RECT 80.310 206.625 80.570 207.775 ;
        RECT 80.745 206.625 81.025 207.765 ;
        RECT 81.195 206.795 81.525 207.775 ;
        RECT 82.585 207.765 82.865 208.435 ;
        RECT 83.140 208.375 84.265 208.545 ;
        RECT 83.140 208.265 83.590 208.375 ;
        RECT 83.035 207.935 83.590 208.265 ;
        RECT 84.455 208.205 84.855 209.005 ;
        RECT 85.255 208.715 85.525 209.175 ;
        RECT 85.695 208.545 85.980 209.005 ;
        RECT 81.695 206.625 81.955 207.765 ;
        RECT 82.585 206.795 82.970 207.765 ;
        RECT 83.140 207.475 83.590 207.935 ;
        RECT 83.760 207.645 84.855 208.205 ;
        RECT 83.140 207.255 84.265 207.475 ;
        RECT 83.140 206.625 83.465 207.085 ;
        RECT 83.985 206.795 84.265 207.255 ;
        RECT 84.455 206.795 84.855 207.645 ;
        RECT 85.025 208.375 85.980 208.545 ;
        RECT 87.185 208.450 87.475 209.175 ;
        RECT 87.750 208.705 87.920 209.175 ;
        RECT 88.090 208.535 88.420 209.005 ;
        RECT 88.590 208.705 88.760 209.175 ;
        RECT 88.930 208.535 89.180 209.005 ;
        RECT 89.360 208.775 89.740 209.175 ;
        RECT 89.960 208.605 90.130 208.955 ;
        RECT 90.300 208.775 90.630 209.175 ;
        RECT 90.830 208.605 91.000 208.955 ;
        RECT 91.330 208.675 91.580 209.175 ;
        RECT 85.025 207.475 85.235 208.375 ;
        RECT 87.645 208.355 89.180 208.535 ;
        RECT 89.350 208.435 91.160 208.605 ;
        RECT 85.405 207.645 86.095 208.205 ;
        RECT 87.645 207.805 87.890 208.355 ;
        RECT 89.350 208.185 89.520 208.435 ;
        RECT 88.060 208.015 89.520 208.185 ;
        RECT 89.690 207.815 89.860 208.265 ;
        RECT 85.025 207.255 85.980 207.475 ;
        RECT 85.255 206.625 85.525 207.085 ;
        RECT 85.695 206.795 85.980 207.255 ;
        RECT 87.185 206.625 87.475 207.790 ;
        RECT 87.645 207.635 89.220 207.805 ;
        RECT 89.425 207.645 89.860 207.815 ;
        RECT 90.090 207.810 90.420 208.265 ;
        RECT 87.710 206.625 87.960 207.465 ;
        RECT 88.130 206.795 88.380 207.635 ;
        RECT 88.550 206.625 88.800 207.465 ;
        RECT 88.970 206.795 89.220 207.635 ;
        RECT 90.090 207.475 90.300 207.810 ;
        RECT 90.650 207.640 90.820 208.265 ;
        RECT 89.445 206.625 89.695 207.465 ;
        RECT 89.980 206.885 90.300 207.475 ;
        RECT 90.470 206.885 90.820 207.640 ;
        RECT 90.990 207.765 91.160 208.435 ;
        RECT 91.330 207.935 91.615 208.505 ;
        RECT 91.785 208.405 93.455 209.175 ;
        RECT 93.715 208.625 93.885 209.005 ;
        RECT 94.100 208.795 94.430 209.175 ;
        RECT 93.715 208.455 94.430 208.625 ;
        RECT 91.785 207.885 92.535 208.405 ;
        RECT 90.990 207.595 91.585 207.765 ;
        RECT 92.705 207.715 93.455 208.235 ;
        RECT 93.625 207.905 93.980 208.275 ;
        RECT 94.260 208.265 94.430 208.455 ;
        RECT 94.600 208.430 94.855 209.005 ;
        RECT 94.260 207.935 94.515 208.265 ;
        RECT 94.260 207.725 94.430 207.935 ;
        RECT 91.250 206.810 91.585 207.595 ;
        RECT 91.785 206.625 93.455 207.715 ;
        RECT 93.715 207.555 94.430 207.725 ;
        RECT 94.685 207.700 94.855 208.430 ;
        RECT 95.030 208.335 95.290 209.175 ;
        RECT 95.465 208.405 98.975 209.175 ;
        RECT 100.065 208.450 100.355 209.175 ;
        RECT 100.525 208.500 100.800 208.845 ;
        RECT 100.990 208.775 101.365 209.175 ;
        RECT 101.535 208.605 101.705 208.955 ;
        RECT 101.875 208.775 102.205 209.175 ;
        RECT 102.375 208.605 102.635 209.005 ;
        RECT 95.465 207.885 97.115 208.405 ;
        RECT 93.715 206.795 93.885 207.555 ;
        RECT 94.100 206.625 94.430 207.385 ;
        RECT 94.600 206.795 94.855 207.700 ;
        RECT 95.030 206.625 95.290 207.775 ;
        RECT 97.285 207.715 98.975 208.235 ;
        RECT 95.465 206.625 98.975 207.715 ;
        RECT 100.065 206.625 100.355 207.790 ;
        RECT 100.525 207.765 100.695 208.500 ;
        RECT 100.970 208.435 102.635 208.605 ;
        RECT 100.970 208.265 101.140 208.435 ;
        RECT 102.815 208.355 103.145 208.775 ;
        RECT 103.315 208.355 103.575 209.175 ;
        RECT 103.835 208.625 104.005 209.005 ;
        RECT 104.185 208.795 104.515 209.175 ;
        RECT 103.835 208.455 104.500 208.625 ;
        RECT 104.695 208.500 104.955 209.005 ;
        RECT 102.815 208.265 103.065 208.355 ;
        RECT 100.865 207.935 101.140 208.265 ;
        RECT 101.310 207.935 102.135 208.265 ;
        RECT 102.350 207.935 103.065 208.265 ;
        RECT 103.235 207.935 103.570 208.185 ;
        RECT 100.970 207.765 101.140 207.935 ;
        RECT 100.525 206.795 100.800 207.765 ;
        RECT 100.970 207.595 101.630 207.765 ;
        RECT 101.890 207.645 102.135 207.935 ;
        RECT 101.460 207.475 101.630 207.595 ;
        RECT 102.305 207.475 102.635 207.765 ;
        RECT 101.010 206.625 101.290 207.425 ;
        RECT 101.460 207.305 102.635 207.475 ;
        RECT 102.895 207.375 103.065 207.935 ;
        RECT 103.765 207.905 104.095 208.275 ;
        RECT 104.330 208.200 104.500 208.455 ;
        RECT 104.330 207.870 104.615 208.200 ;
        RECT 101.460 206.805 103.075 207.135 ;
        RECT 103.315 206.625 103.575 207.765 ;
        RECT 104.330 207.725 104.500 207.870 ;
        RECT 103.835 207.555 104.500 207.725 ;
        RECT 104.785 207.700 104.955 208.500 ;
        RECT 105.125 208.405 106.795 209.175 ;
        RECT 107.425 208.675 107.685 209.005 ;
        RECT 107.855 208.815 108.185 209.175 ;
        RECT 108.440 208.795 109.740 209.005 ;
        RECT 105.125 207.885 105.875 208.405 ;
        RECT 106.045 207.715 106.795 208.235 ;
        RECT 103.835 206.795 104.005 207.555 ;
        RECT 104.185 206.625 104.515 207.385 ;
        RECT 104.685 206.795 104.955 207.700 ;
        RECT 105.125 206.625 106.795 207.715 ;
        RECT 107.425 207.475 107.595 208.675 ;
        RECT 108.440 208.645 108.610 208.795 ;
        RECT 107.855 208.520 108.610 208.645 ;
        RECT 107.765 208.475 108.610 208.520 ;
        RECT 107.765 208.355 108.035 208.475 ;
        RECT 107.765 207.780 107.935 208.355 ;
        RECT 108.165 207.915 108.575 208.220 ;
        RECT 108.865 208.185 109.075 208.585 ;
        RECT 108.745 207.975 109.075 208.185 ;
        RECT 109.320 208.185 109.540 208.585 ;
        RECT 110.015 208.410 110.470 209.175 ;
        RECT 110.650 208.775 110.985 209.175 ;
        RECT 111.155 208.605 111.360 209.005 ;
        RECT 111.570 208.695 111.845 209.175 ;
        RECT 112.055 208.675 112.315 209.005 ;
        RECT 110.675 208.435 111.360 208.605 ;
        RECT 109.320 207.975 109.795 208.185 ;
        RECT 109.985 207.985 110.475 208.185 ;
        RECT 107.765 207.745 107.965 207.780 ;
        RECT 109.295 207.745 110.470 207.805 ;
        RECT 107.765 207.635 110.470 207.745 ;
        RECT 107.825 207.575 109.625 207.635 ;
        RECT 109.295 207.545 109.625 207.575 ;
        RECT 107.425 206.795 107.685 207.475 ;
        RECT 107.855 206.625 108.105 207.405 ;
        RECT 108.355 207.375 109.190 207.385 ;
        RECT 109.780 207.375 109.965 207.465 ;
        RECT 108.355 207.175 109.965 207.375 ;
        RECT 108.355 206.795 108.605 207.175 ;
        RECT 109.735 207.135 109.965 207.175 ;
        RECT 110.215 207.015 110.470 207.635 ;
        RECT 110.675 207.405 111.015 208.435 ;
        RECT 111.185 207.765 111.435 208.265 ;
        RECT 111.615 207.935 111.975 208.515 ;
        RECT 112.145 207.765 112.315 208.675 ;
        RECT 112.945 208.450 113.235 209.175 ;
        RECT 113.410 208.410 113.865 209.175 ;
        RECT 114.140 208.795 115.440 209.005 ;
        RECT 115.695 208.815 116.025 209.175 ;
        RECT 115.270 208.645 115.440 208.795 ;
        RECT 116.195 208.675 116.455 209.005 ;
        RECT 114.340 208.185 114.560 208.585 ;
        RECT 113.405 207.985 113.895 208.185 ;
        RECT 114.085 207.975 114.560 208.185 ;
        RECT 114.805 208.185 115.015 208.585 ;
        RECT 115.270 208.520 116.025 208.645 ;
        RECT 115.270 208.475 116.115 208.520 ;
        RECT 115.845 208.355 116.115 208.475 ;
        RECT 114.805 207.975 115.135 208.185 ;
        RECT 115.305 207.915 115.715 208.220 ;
        RECT 111.185 207.595 112.315 207.765 ;
        RECT 110.675 207.230 111.340 207.405 ;
        RECT 108.775 206.625 109.130 207.005 ;
        RECT 110.135 206.795 110.470 207.015 ;
        RECT 110.650 206.625 110.985 207.050 ;
        RECT 111.155 206.825 111.340 207.230 ;
        RECT 111.545 206.625 111.875 207.405 ;
        RECT 112.045 206.825 112.315 207.595 ;
        RECT 112.945 206.625 113.235 207.790 ;
        RECT 113.410 207.745 114.585 207.805 ;
        RECT 115.945 207.780 116.115 208.355 ;
        RECT 115.915 207.745 116.115 207.780 ;
        RECT 113.410 207.635 116.115 207.745 ;
        RECT 113.410 207.015 113.665 207.635 ;
        RECT 114.255 207.575 116.055 207.635 ;
        RECT 114.255 207.545 114.585 207.575 ;
        RECT 116.285 207.475 116.455 208.675 ;
        RECT 113.915 207.375 114.100 207.465 ;
        RECT 114.690 207.375 115.525 207.385 ;
        RECT 113.915 207.175 115.525 207.375 ;
        RECT 113.915 207.135 114.145 207.175 ;
        RECT 113.410 206.795 113.745 207.015 ;
        RECT 114.750 206.625 115.105 207.005 ;
        RECT 115.275 206.795 115.525 207.175 ;
        RECT 115.775 206.625 116.025 207.405 ;
        RECT 116.195 206.795 116.455 207.475 ;
        RECT 117.545 208.435 117.930 209.005 ;
        RECT 118.100 208.715 118.425 209.175 ;
        RECT 118.945 208.545 119.225 209.005 ;
        RECT 117.545 207.765 117.825 208.435 ;
        RECT 118.100 208.375 119.225 208.545 ;
        RECT 118.100 208.265 118.550 208.375 ;
        RECT 117.995 207.935 118.550 208.265 ;
        RECT 119.415 208.205 119.815 209.005 ;
        RECT 120.215 208.715 120.485 209.175 ;
        RECT 120.655 208.545 120.940 209.005 ;
        RECT 121.230 208.775 121.565 209.175 ;
        RECT 121.735 208.605 121.940 209.005 ;
        RECT 122.150 208.695 122.425 209.175 ;
        RECT 122.635 208.675 122.895 209.005 ;
        RECT 123.070 208.775 123.405 209.175 ;
        RECT 117.545 206.795 117.930 207.765 ;
        RECT 118.100 207.475 118.550 207.935 ;
        RECT 118.720 207.645 119.815 208.205 ;
        RECT 118.100 207.255 119.225 207.475 ;
        RECT 118.100 206.625 118.425 207.085 ;
        RECT 118.945 206.795 119.225 207.255 ;
        RECT 119.415 206.795 119.815 207.645 ;
        RECT 119.985 208.375 120.940 208.545 ;
        RECT 121.255 208.435 121.940 208.605 ;
        RECT 119.985 207.475 120.195 208.375 ;
        RECT 120.365 207.645 121.055 208.205 ;
        RECT 119.985 207.255 120.940 207.475 ;
        RECT 120.215 206.625 120.485 207.085 ;
        RECT 120.655 206.795 120.940 207.255 ;
        RECT 121.255 207.405 121.595 208.435 ;
        RECT 121.765 207.765 122.015 208.265 ;
        RECT 122.195 207.935 122.555 208.515 ;
        RECT 122.725 207.765 122.895 208.675 ;
        RECT 123.575 208.605 123.780 209.005 ;
        RECT 123.990 208.695 124.265 209.175 ;
        RECT 124.475 208.675 124.735 209.005 ;
        RECT 121.765 207.595 122.895 207.765 ;
        RECT 121.255 207.230 121.920 207.405 ;
        RECT 121.230 206.625 121.565 207.050 ;
        RECT 121.735 206.825 121.920 207.230 ;
        RECT 122.125 206.625 122.455 207.405 ;
        RECT 122.625 206.825 122.895 207.595 ;
        RECT 123.095 208.435 123.780 208.605 ;
        RECT 123.095 207.405 123.435 208.435 ;
        RECT 123.605 207.765 123.855 208.265 ;
        RECT 124.035 207.935 124.395 208.515 ;
        RECT 124.565 207.765 124.735 208.675 ;
        RECT 125.825 208.450 126.115 209.175 ;
        RECT 126.285 208.405 129.795 209.175 ;
        RECT 130.430 208.775 130.765 209.175 ;
        RECT 130.935 208.605 131.140 209.005 ;
        RECT 131.350 208.695 131.625 209.175 ;
        RECT 131.835 208.675 132.095 209.005 ;
        RECT 130.455 208.435 131.140 208.605 ;
        RECT 126.285 207.885 127.935 208.405 ;
        RECT 123.605 207.595 124.735 207.765 ;
        RECT 123.095 207.230 123.760 207.405 ;
        RECT 123.070 206.625 123.405 207.050 ;
        RECT 123.575 206.825 123.760 207.230 ;
        RECT 123.965 206.625 124.295 207.405 ;
        RECT 124.465 206.825 124.735 207.595 ;
        RECT 125.825 206.625 126.115 207.790 ;
        RECT 128.105 207.715 129.795 208.235 ;
        RECT 126.285 206.625 129.795 207.715 ;
        RECT 130.455 207.405 130.795 208.435 ;
        RECT 130.965 207.765 131.215 208.265 ;
        RECT 131.395 207.935 131.755 208.515 ;
        RECT 131.925 207.765 132.095 208.675 ;
        RECT 132.265 208.425 133.475 209.175 ;
        RECT 133.645 208.500 133.905 209.005 ;
        RECT 134.085 208.795 134.415 209.175 ;
        RECT 134.595 208.625 134.765 209.005 ;
        RECT 132.265 207.885 132.785 208.425 ;
        RECT 130.965 207.595 132.095 207.765 ;
        RECT 132.955 207.715 133.475 208.255 ;
        RECT 130.455 207.230 131.120 207.405 ;
        RECT 130.430 206.625 130.765 207.050 ;
        RECT 130.935 206.825 131.120 207.230 ;
        RECT 131.325 206.625 131.655 207.405 ;
        RECT 131.825 206.825 132.095 207.595 ;
        RECT 132.265 206.625 133.475 207.715 ;
        RECT 133.645 207.700 133.815 208.500 ;
        RECT 134.100 208.455 134.765 208.625 ;
        RECT 134.100 208.200 134.270 208.455 ;
        RECT 135.025 208.405 138.535 209.175 ;
        RECT 138.705 208.450 138.995 209.175 ;
        RECT 139.165 208.605 139.600 209.005 ;
        RECT 139.770 208.775 140.155 209.175 ;
        RECT 139.165 208.435 140.155 208.605 ;
        RECT 140.325 208.435 140.750 209.005 ;
        RECT 140.940 208.605 141.195 209.005 ;
        RECT 141.365 208.775 141.750 209.175 ;
        RECT 140.940 208.435 141.750 208.605 ;
        RECT 141.920 208.435 142.165 209.005 ;
        RECT 142.355 208.605 142.610 209.005 ;
        RECT 142.780 208.775 143.165 209.175 ;
        RECT 142.355 208.435 143.165 208.605 ;
        RECT 143.335 208.435 143.595 209.005 ;
        RECT 143.765 208.630 149.110 209.175 ;
        RECT 133.985 207.870 134.270 208.200 ;
        RECT 134.505 207.905 134.835 208.275 ;
        RECT 135.025 207.885 136.675 208.405 ;
        RECT 139.820 208.265 140.155 208.435 ;
        RECT 140.400 208.265 140.750 208.435 ;
        RECT 141.400 208.265 141.750 208.435 ;
        RECT 141.995 208.265 142.165 208.435 ;
        RECT 142.815 208.265 143.165 208.435 ;
        RECT 134.100 207.725 134.270 207.870 ;
        RECT 133.645 206.795 133.915 207.700 ;
        RECT 134.100 207.555 134.765 207.725 ;
        RECT 136.845 207.715 138.535 208.235 ;
        RECT 134.085 206.625 134.415 207.385 ;
        RECT 134.595 206.795 134.765 207.555 ;
        RECT 135.025 206.625 138.535 207.715 ;
        RECT 138.705 206.625 138.995 207.790 ;
        RECT 139.165 207.560 139.650 208.265 ;
        RECT 139.820 207.935 140.230 208.265 ;
        RECT 139.820 207.390 140.155 207.935 ;
        RECT 140.400 207.765 141.230 208.265 ;
        RECT 139.165 207.220 140.155 207.390 ;
        RECT 140.325 207.585 141.230 207.765 ;
        RECT 141.400 207.935 141.825 208.265 ;
        RECT 139.165 206.795 139.600 207.220 ;
        RECT 139.770 206.625 140.155 207.050 ;
        RECT 140.325 206.795 140.750 207.585 ;
        RECT 141.400 207.415 141.750 207.935 ;
        RECT 141.995 207.765 142.645 208.265 ;
        RECT 140.920 207.220 141.750 207.415 ;
        RECT 141.920 207.585 142.645 207.765 ;
        RECT 142.815 207.935 143.240 208.265 ;
        RECT 140.920 206.795 141.195 207.220 ;
        RECT 141.365 206.625 141.750 207.050 ;
        RECT 141.920 206.795 142.165 207.585 ;
        RECT 142.815 207.415 143.165 207.935 ;
        RECT 143.410 207.765 143.595 208.435 ;
        RECT 145.350 207.800 145.690 208.630 ;
        RECT 149.285 208.405 150.955 209.175 ;
        RECT 151.585 208.450 151.875 209.175 ;
        RECT 152.505 208.500 152.765 209.005 ;
        RECT 152.945 208.795 153.275 209.175 ;
        RECT 153.455 208.625 153.625 209.005 ;
        RECT 142.355 207.220 143.165 207.415 ;
        RECT 142.355 206.795 142.610 207.220 ;
        RECT 142.780 206.625 143.165 207.050 ;
        RECT 143.335 206.795 143.595 207.765 ;
        RECT 147.170 207.060 147.520 208.310 ;
        RECT 149.285 207.885 150.035 208.405 ;
        RECT 150.205 207.715 150.955 208.235 ;
        RECT 143.765 206.625 149.110 207.060 ;
        RECT 149.285 206.625 150.955 207.715 ;
        RECT 151.585 206.625 151.875 207.790 ;
        RECT 152.505 207.700 152.675 208.500 ;
        RECT 152.960 208.455 153.625 208.625 ;
        RECT 152.960 208.200 153.130 208.455 ;
        RECT 153.885 208.405 155.555 209.175 ;
        RECT 155.725 208.425 156.935 209.175 ;
        RECT 152.845 207.870 153.130 208.200 ;
        RECT 153.365 207.905 153.695 208.275 ;
        RECT 153.885 207.885 154.635 208.405 ;
        RECT 152.960 207.725 153.130 207.870 ;
        RECT 152.505 206.795 152.775 207.700 ;
        RECT 152.960 207.555 153.625 207.725 ;
        RECT 154.805 207.715 155.555 208.235 ;
        RECT 152.945 206.625 153.275 207.385 ;
        RECT 153.455 206.795 153.625 207.555 ;
        RECT 153.885 206.625 155.555 207.715 ;
        RECT 155.725 207.715 156.245 208.255 ;
        RECT 156.415 207.885 156.935 208.425 ;
        RECT 155.725 206.625 156.935 207.715 ;
        RECT 22.700 206.455 157.020 206.625 ;
        RECT 22.785 205.365 23.995 206.455 ;
        RECT 24.165 205.365 27.675 206.455 ;
        RECT 28.025 205.540 28.195 206.455 ;
        RECT 28.365 205.395 28.695 206.240 ;
        RECT 28.865 205.445 29.035 206.455 ;
        RECT 29.205 205.725 29.545 206.285 ;
        RECT 29.775 205.955 30.090 206.455 ;
        RECT 30.270 205.985 31.155 206.155 ;
        RECT 22.785 204.655 23.305 205.195 ;
        RECT 23.475 204.825 23.995 205.365 ;
        RECT 24.165 204.675 25.815 205.195 ;
        RECT 25.985 204.845 27.675 205.365 ;
        RECT 28.305 205.315 28.695 205.395 ;
        RECT 29.205 205.350 30.100 205.725 ;
        RECT 28.305 205.265 28.520 205.315 ;
        RECT 28.305 204.685 28.475 205.265 ;
        RECT 29.205 205.145 29.395 205.350 ;
        RECT 30.270 205.145 30.440 205.985 ;
        RECT 31.380 205.955 31.630 206.285 ;
        RECT 28.645 204.815 29.395 205.145 ;
        RECT 29.565 204.815 30.440 205.145 ;
        RECT 22.785 203.905 23.995 204.655 ;
        RECT 24.165 203.905 27.675 204.675 ;
        RECT 28.305 204.645 28.530 204.685 ;
        RECT 29.195 204.645 29.395 204.815 ;
        RECT 28.305 204.560 28.685 204.645 ;
        RECT 28.015 203.905 28.185 204.420 ;
        RECT 28.355 204.125 28.685 204.560 ;
        RECT 28.855 203.905 29.025 204.515 ;
        RECT 29.195 204.120 29.525 204.645 ;
        RECT 29.785 203.905 29.995 204.435 ;
        RECT 30.270 204.355 30.440 204.815 ;
        RECT 30.610 204.855 30.930 205.815 ;
        RECT 31.100 205.065 31.290 205.785 ;
        RECT 31.460 204.885 31.630 205.955 ;
        RECT 31.800 205.655 31.970 206.455 ;
        RECT 32.140 206.010 33.245 206.180 ;
        RECT 32.140 205.395 32.310 206.010 ;
        RECT 33.455 205.860 33.705 206.285 ;
        RECT 33.875 205.995 34.140 206.455 ;
        RECT 32.480 205.475 33.010 205.840 ;
        RECT 33.455 205.730 33.760 205.860 ;
        RECT 31.800 205.305 32.310 205.395 ;
        RECT 31.800 205.135 32.670 205.305 ;
        RECT 31.800 205.065 31.970 205.135 ;
        RECT 32.090 204.885 32.290 204.915 ;
        RECT 30.610 204.525 31.075 204.855 ;
        RECT 31.460 204.585 32.290 204.885 ;
        RECT 31.460 204.355 31.630 204.585 ;
        RECT 30.270 204.185 31.055 204.355 ;
        RECT 31.225 204.185 31.630 204.355 ;
        RECT 31.810 203.905 32.180 204.405 ;
        RECT 32.500 204.355 32.670 205.135 ;
        RECT 32.840 204.775 33.010 205.475 ;
        RECT 33.180 204.945 33.420 205.540 ;
        RECT 32.840 204.555 33.365 204.775 ;
        RECT 33.590 204.625 33.760 205.730 ;
        RECT 33.535 204.495 33.760 204.625 ;
        RECT 33.930 204.535 34.210 205.485 ;
        RECT 33.535 204.355 33.705 204.495 ;
        RECT 32.500 204.185 33.175 204.355 ;
        RECT 33.370 204.185 33.705 204.355 ;
        RECT 33.875 203.905 34.125 204.365 ;
        RECT 34.380 204.165 34.565 206.285 ;
        RECT 34.735 205.955 35.065 206.455 ;
        RECT 35.235 205.785 35.405 206.285 ;
        RECT 34.740 205.615 35.405 205.785 ;
        RECT 34.740 204.625 34.970 205.615 ;
        RECT 35.140 204.795 35.490 205.445 ;
        RECT 35.665 205.290 35.955 206.455 ;
        RECT 36.215 205.785 36.385 206.285 ;
        RECT 36.555 205.955 36.885 206.455 ;
        RECT 36.215 205.615 36.880 205.785 ;
        RECT 36.130 204.795 36.480 205.445 ;
        RECT 34.740 204.455 35.405 204.625 ;
        RECT 34.735 203.905 35.065 204.285 ;
        RECT 35.235 204.165 35.405 204.455 ;
        RECT 35.665 203.905 35.955 204.630 ;
        RECT 36.650 204.625 36.880 205.615 ;
        RECT 36.215 204.455 36.880 204.625 ;
        RECT 36.215 204.165 36.385 204.455 ;
        RECT 36.555 203.905 36.885 204.285 ;
        RECT 37.055 204.165 37.240 206.285 ;
        RECT 37.480 205.995 37.745 206.455 ;
        RECT 37.915 205.860 38.165 206.285 ;
        RECT 38.375 206.010 39.480 206.180 ;
        RECT 37.860 205.730 38.165 205.860 ;
        RECT 37.410 204.535 37.690 205.485 ;
        RECT 37.860 204.625 38.030 205.730 ;
        RECT 38.200 204.945 38.440 205.540 ;
        RECT 38.610 205.475 39.140 205.840 ;
        RECT 38.610 204.775 38.780 205.475 ;
        RECT 39.310 205.395 39.480 206.010 ;
        RECT 39.650 205.655 39.820 206.455 ;
        RECT 39.990 205.955 40.240 206.285 ;
        RECT 40.465 205.985 41.350 206.155 ;
        RECT 39.310 205.305 39.820 205.395 ;
        RECT 37.860 204.495 38.085 204.625 ;
        RECT 38.255 204.555 38.780 204.775 ;
        RECT 38.950 205.135 39.820 205.305 ;
        RECT 37.495 203.905 37.745 204.365 ;
        RECT 37.915 204.355 38.085 204.495 ;
        RECT 38.950 204.355 39.120 205.135 ;
        RECT 39.650 205.065 39.820 205.135 ;
        RECT 39.330 204.885 39.530 204.915 ;
        RECT 39.990 204.885 40.160 205.955 ;
        RECT 40.330 205.065 40.520 205.785 ;
        RECT 39.330 204.585 40.160 204.885 ;
        RECT 40.690 204.855 41.010 205.815 ;
        RECT 37.915 204.185 38.250 204.355 ;
        RECT 38.445 204.185 39.120 204.355 ;
        RECT 39.440 203.905 39.810 204.405 ;
        RECT 39.990 204.355 40.160 204.585 ;
        RECT 40.545 204.525 41.010 204.855 ;
        RECT 41.180 205.145 41.350 205.985 ;
        RECT 41.530 205.955 41.845 206.455 ;
        RECT 42.075 205.725 42.415 206.285 ;
        RECT 41.520 205.350 42.415 205.725 ;
        RECT 42.585 205.445 42.755 206.455 ;
        RECT 42.225 205.145 42.415 205.350 ;
        RECT 42.925 205.395 43.255 206.240 ;
        RECT 43.425 205.540 43.595 206.455 ;
        RECT 44.035 205.785 44.205 206.285 ;
        RECT 44.375 205.955 44.705 206.455 ;
        RECT 44.035 205.615 44.700 205.785 ;
        RECT 42.925 205.315 43.315 205.395 ;
        RECT 43.100 205.265 43.315 205.315 ;
        RECT 41.180 204.815 42.055 205.145 ;
        RECT 42.225 204.815 42.975 205.145 ;
        RECT 41.180 204.355 41.350 204.815 ;
        RECT 42.225 204.645 42.425 204.815 ;
        RECT 43.145 204.685 43.315 205.265 ;
        RECT 43.950 204.795 44.300 205.445 ;
        RECT 43.090 204.645 43.315 204.685 ;
        RECT 39.990 204.185 40.395 204.355 ;
        RECT 40.565 204.185 41.350 204.355 ;
        RECT 41.625 203.905 41.835 204.435 ;
        RECT 42.095 204.120 42.425 204.645 ;
        RECT 42.935 204.560 43.315 204.645 ;
        RECT 44.470 204.625 44.700 205.615 ;
        RECT 42.595 203.905 42.765 204.515 ;
        RECT 42.935 204.125 43.265 204.560 ;
        RECT 44.035 204.455 44.700 204.625 ;
        RECT 43.435 203.905 43.605 204.420 ;
        RECT 44.035 204.165 44.205 204.455 ;
        RECT 44.375 203.905 44.705 204.285 ;
        RECT 44.875 204.165 45.060 206.285 ;
        RECT 45.300 205.995 45.565 206.455 ;
        RECT 45.735 205.860 45.985 206.285 ;
        RECT 46.195 206.010 47.300 206.180 ;
        RECT 45.680 205.730 45.985 205.860 ;
        RECT 45.230 204.535 45.510 205.485 ;
        RECT 45.680 204.625 45.850 205.730 ;
        RECT 46.020 204.945 46.260 205.540 ;
        RECT 46.430 205.475 46.960 205.840 ;
        RECT 46.430 204.775 46.600 205.475 ;
        RECT 47.130 205.395 47.300 206.010 ;
        RECT 47.470 205.655 47.640 206.455 ;
        RECT 47.810 205.955 48.060 206.285 ;
        RECT 48.285 205.985 49.170 206.155 ;
        RECT 47.130 205.305 47.640 205.395 ;
        RECT 45.680 204.495 45.905 204.625 ;
        RECT 46.075 204.555 46.600 204.775 ;
        RECT 46.770 205.135 47.640 205.305 ;
        RECT 45.315 203.905 45.565 204.365 ;
        RECT 45.735 204.355 45.905 204.495 ;
        RECT 46.770 204.355 46.940 205.135 ;
        RECT 47.470 205.065 47.640 205.135 ;
        RECT 47.150 204.885 47.350 204.915 ;
        RECT 47.810 204.885 47.980 205.955 ;
        RECT 48.150 205.065 48.340 205.785 ;
        RECT 47.150 204.585 47.980 204.885 ;
        RECT 48.510 204.855 48.830 205.815 ;
        RECT 45.735 204.185 46.070 204.355 ;
        RECT 46.265 204.185 46.940 204.355 ;
        RECT 47.260 203.905 47.630 204.405 ;
        RECT 47.810 204.355 47.980 204.585 ;
        RECT 48.365 204.525 48.830 204.855 ;
        RECT 49.000 205.145 49.170 205.985 ;
        RECT 49.350 205.955 49.665 206.455 ;
        RECT 49.895 205.725 50.235 206.285 ;
        RECT 49.340 205.350 50.235 205.725 ;
        RECT 50.405 205.445 50.575 206.455 ;
        RECT 50.045 205.145 50.235 205.350 ;
        RECT 50.745 205.395 51.075 206.240 ;
        RECT 50.745 205.315 51.135 205.395 ;
        RECT 50.920 205.265 51.135 205.315 ;
        RECT 49.000 204.815 49.875 205.145 ;
        RECT 50.045 204.815 50.795 205.145 ;
        RECT 49.000 204.355 49.170 204.815 ;
        RECT 50.045 204.645 50.245 204.815 ;
        RECT 50.965 204.685 51.135 205.265 ;
        RECT 50.910 204.645 51.135 204.685 ;
        RECT 47.810 204.185 48.215 204.355 ;
        RECT 48.385 204.185 49.170 204.355 ;
        RECT 49.445 203.905 49.655 204.435 ;
        RECT 49.915 204.120 50.245 204.645 ;
        RECT 50.755 204.560 51.135 204.645 ;
        RECT 51.765 205.380 52.035 206.285 ;
        RECT 52.205 205.695 52.535 206.455 ;
        RECT 52.715 205.525 52.885 206.285 ;
        RECT 53.235 205.785 53.405 206.285 ;
        RECT 53.575 205.955 53.905 206.455 ;
        RECT 53.235 205.615 53.900 205.785 ;
        RECT 51.765 204.580 51.935 205.380 ;
        RECT 52.220 205.355 52.885 205.525 ;
        RECT 52.220 205.210 52.390 205.355 ;
        RECT 52.105 204.880 52.390 205.210 ;
        RECT 52.220 204.625 52.390 204.880 ;
        RECT 52.625 204.805 52.955 205.175 ;
        RECT 53.150 204.795 53.500 205.445 ;
        RECT 53.670 204.625 53.900 205.615 ;
        RECT 50.415 203.905 50.585 204.515 ;
        RECT 50.755 204.125 51.085 204.560 ;
        RECT 51.765 204.075 52.025 204.580 ;
        RECT 52.220 204.455 52.885 204.625 ;
        RECT 52.205 203.905 52.535 204.285 ;
        RECT 52.715 204.075 52.885 204.455 ;
        RECT 53.235 204.455 53.900 204.625 ;
        RECT 53.235 204.165 53.405 204.455 ;
        RECT 53.575 203.905 53.905 204.285 ;
        RECT 54.075 204.165 54.260 206.285 ;
        RECT 54.500 205.995 54.765 206.455 ;
        RECT 54.935 205.860 55.185 206.285 ;
        RECT 55.395 206.010 56.500 206.180 ;
        RECT 54.880 205.730 55.185 205.860 ;
        RECT 54.430 204.535 54.710 205.485 ;
        RECT 54.880 204.625 55.050 205.730 ;
        RECT 55.220 204.945 55.460 205.540 ;
        RECT 55.630 205.475 56.160 205.840 ;
        RECT 55.630 204.775 55.800 205.475 ;
        RECT 56.330 205.395 56.500 206.010 ;
        RECT 56.670 205.655 56.840 206.455 ;
        RECT 57.010 205.955 57.260 206.285 ;
        RECT 57.485 205.985 58.370 206.155 ;
        RECT 56.330 205.305 56.840 205.395 ;
        RECT 54.880 204.495 55.105 204.625 ;
        RECT 55.275 204.555 55.800 204.775 ;
        RECT 55.970 205.135 56.840 205.305 ;
        RECT 54.515 203.905 54.765 204.365 ;
        RECT 54.935 204.355 55.105 204.495 ;
        RECT 55.970 204.355 56.140 205.135 ;
        RECT 56.670 205.065 56.840 205.135 ;
        RECT 56.350 204.885 56.550 204.915 ;
        RECT 57.010 204.885 57.180 205.955 ;
        RECT 57.350 205.065 57.540 205.785 ;
        RECT 56.350 204.585 57.180 204.885 ;
        RECT 57.710 204.855 58.030 205.815 ;
        RECT 54.935 204.185 55.270 204.355 ;
        RECT 55.465 204.185 56.140 204.355 ;
        RECT 56.460 203.905 56.830 204.405 ;
        RECT 57.010 204.355 57.180 204.585 ;
        RECT 57.565 204.525 58.030 204.855 ;
        RECT 58.200 205.145 58.370 205.985 ;
        RECT 58.550 205.955 58.865 206.455 ;
        RECT 59.095 205.725 59.435 206.285 ;
        RECT 58.540 205.350 59.435 205.725 ;
        RECT 59.605 205.445 59.775 206.455 ;
        RECT 59.245 205.145 59.435 205.350 ;
        RECT 59.945 205.395 60.275 206.240 ;
        RECT 59.945 205.315 60.335 205.395 ;
        RECT 60.120 205.265 60.335 205.315 ;
        RECT 61.425 205.290 61.715 206.455 ;
        RECT 61.885 205.315 62.165 206.455 ;
        RECT 62.335 205.305 62.665 206.285 ;
        RECT 62.835 205.315 63.095 206.455 ;
        RECT 63.265 205.380 63.535 206.285 ;
        RECT 63.705 205.695 64.035 206.455 ;
        RECT 64.215 205.525 64.385 206.285 ;
        RECT 58.200 204.815 59.075 205.145 ;
        RECT 59.245 204.815 59.995 205.145 ;
        RECT 58.200 204.355 58.370 204.815 ;
        RECT 59.245 204.645 59.445 204.815 ;
        RECT 60.165 204.685 60.335 205.265 ;
        RECT 61.895 204.875 62.230 205.145 ;
        RECT 62.400 204.705 62.570 205.305 ;
        RECT 62.740 204.895 63.075 205.145 ;
        RECT 60.110 204.645 60.335 204.685 ;
        RECT 57.010 204.185 57.415 204.355 ;
        RECT 57.585 204.185 58.370 204.355 ;
        RECT 58.645 203.905 58.855 204.435 ;
        RECT 59.115 204.120 59.445 204.645 ;
        RECT 59.955 204.560 60.335 204.645 ;
        RECT 59.615 203.905 59.785 204.515 ;
        RECT 59.955 204.125 60.285 204.560 ;
        RECT 61.425 203.905 61.715 204.630 ;
        RECT 61.885 203.905 62.195 204.705 ;
        RECT 62.400 204.075 63.095 204.705 ;
        RECT 63.265 204.580 63.435 205.380 ;
        RECT 63.720 205.355 64.385 205.525 ;
        RECT 63.720 205.210 63.890 205.355 ;
        RECT 64.705 205.315 64.915 206.455 ;
        RECT 63.605 204.880 63.890 205.210 ;
        RECT 65.085 205.305 65.415 206.285 ;
        RECT 65.585 205.315 65.815 206.455 ;
        RECT 66.115 205.525 66.285 206.285 ;
        RECT 66.465 205.695 66.795 206.455 ;
        RECT 66.115 205.355 66.780 205.525 ;
        RECT 66.965 205.380 67.235 206.285 ;
        RECT 67.495 205.785 67.665 206.285 ;
        RECT 67.835 205.955 68.165 206.455 ;
        RECT 67.495 205.615 68.160 205.785 ;
        RECT 63.720 204.625 63.890 204.880 ;
        RECT 64.125 204.805 64.455 205.175 ;
        RECT 63.265 204.075 63.525 204.580 ;
        RECT 63.720 204.455 64.385 204.625 ;
        RECT 63.705 203.905 64.035 204.285 ;
        RECT 64.215 204.075 64.385 204.455 ;
        RECT 64.705 203.905 64.915 204.725 ;
        RECT 65.085 204.705 65.335 205.305 ;
        RECT 66.610 205.210 66.780 205.355 ;
        RECT 65.505 204.895 65.835 205.145 ;
        RECT 66.045 204.805 66.375 205.175 ;
        RECT 66.610 204.880 66.895 205.210 ;
        RECT 65.085 204.075 65.415 204.705 ;
        RECT 65.585 203.905 65.815 204.725 ;
        RECT 66.610 204.625 66.780 204.880 ;
        RECT 66.115 204.455 66.780 204.625 ;
        RECT 67.065 204.580 67.235 205.380 ;
        RECT 67.410 204.795 67.760 205.445 ;
        RECT 67.930 204.625 68.160 205.615 ;
        RECT 66.115 204.075 66.285 204.455 ;
        RECT 66.465 203.905 66.795 204.285 ;
        RECT 66.975 204.075 67.235 204.580 ;
        RECT 67.495 204.455 68.160 204.625 ;
        RECT 67.495 204.165 67.665 204.455 ;
        RECT 67.835 203.905 68.165 204.285 ;
        RECT 68.335 204.165 68.520 206.285 ;
        RECT 68.760 205.995 69.025 206.455 ;
        RECT 69.195 205.860 69.445 206.285 ;
        RECT 69.655 206.010 70.760 206.180 ;
        RECT 69.140 205.730 69.445 205.860 ;
        RECT 68.690 204.535 68.970 205.485 ;
        RECT 69.140 204.625 69.310 205.730 ;
        RECT 69.480 204.945 69.720 205.540 ;
        RECT 69.890 205.475 70.420 205.840 ;
        RECT 69.890 204.775 70.060 205.475 ;
        RECT 70.590 205.395 70.760 206.010 ;
        RECT 70.930 205.655 71.100 206.455 ;
        RECT 71.270 205.955 71.520 206.285 ;
        RECT 71.745 205.985 72.630 206.155 ;
        RECT 70.590 205.305 71.100 205.395 ;
        RECT 69.140 204.495 69.365 204.625 ;
        RECT 69.535 204.555 70.060 204.775 ;
        RECT 70.230 205.135 71.100 205.305 ;
        RECT 68.775 203.905 69.025 204.365 ;
        RECT 69.195 204.355 69.365 204.495 ;
        RECT 70.230 204.355 70.400 205.135 ;
        RECT 70.930 205.065 71.100 205.135 ;
        RECT 70.610 204.885 70.810 204.915 ;
        RECT 71.270 204.885 71.440 205.955 ;
        RECT 71.610 205.065 71.800 205.785 ;
        RECT 70.610 204.585 71.440 204.885 ;
        RECT 71.970 204.855 72.290 205.815 ;
        RECT 69.195 204.185 69.530 204.355 ;
        RECT 69.725 204.185 70.400 204.355 ;
        RECT 70.720 203.905 71.090 204.405 ;
        RECT 71.270 204.355 71.440 204.585 ;
        RECT 71.825 204.525 72.290 204.855 ;
        RECT 72.460 205.145 72.630 205.985 ;
        RECT 72.810 205.955 73.125 206.455 ;
        RECT 73.355 205.725 73.695 206.285 ;
        RECT 72.800 205.350 73.695 205.725 ;
        RECT 73.865 205.445 74.035 206.455 ;
        RECT 73.505 205.145 73.695 205.350 ;
        RECT 74.205 205.395 74.535 206.240 ;
        RECT 74.205 205.315 74.595 205.395 ;
        RECT 75.225 205.315 75.505 206.455 ;
        RECT 74.380 205.265 74.595 205.315 ;
        RECT 75.675 205.305 76.005 206.285 ;
        RECT 76.175 205.315 76.435 206.455 ;
        RECT 76.695 205.785 76.865 206.285 ;
        RECT 77.035 205.955 77.365 206.455 ;
        RECT 76.695 205.615 77.360 205.785 ;
        RECT 72.460 204.815 73.335 205.145 ;
        RECT 73.505 204.815 74.255 205.145 ;
        RECT 72.460 204.355 72.630 204.815 ;
        RECT 73.505 204.645 73.705 204.815 ;
        RECT 74.425 204.685 74.595 205.265 ;
        RECT 75.235 204.875 75.570 205.145 ;
        RECT 75.740 204.705 75.910 205.305 ;
        RECT 76.080 204.895 76.415 205.145 ;
        RECT 76.610 204.795 76.960 205.445 ;
        RECT 74.370 204.645 74.595 204.685 ;
        RECT 71.270 204.185 71.675 204.355 ;
        RECT 71.845 204.185 72.630 204.355 ;
        RECT 72.905 203.905 73.115 204.435 ;
        RECT 73.375 204.120 73.705 204.645 ;
        RECT 74.215 204.560 74.595 204.645 ;
        RECT 73.875 203.905 74.045 204.515 ;
        RECT 74.215 204.125 74.545 204.560 ;
        RECT 75.225 203.905 75.535 204.705 ;
        RECT 75.740 204.075 76.435 204.705 ;
        RECT 77.130 204.625 77.360 205.615 ;
        RECT 76.695 204.455 77.360 204.625 ;
        RECT 76.695 204.165 76.865 204.455 ;
        RECT 77.035 203.905 77.365 204.285 ;
        RECT 77.535 204.165 77.720 206.285 ;
        RECT 77.960 205.995 78.225 206.455 ;
        RECT 78.395 205.860 78.645 206.285 ;
        RECT 78.855 206.010 79.960 206.180 ;
        RECT 78.340 205.730 78.645 205.860 ;
        RECT 77.890 204.535 78.170 205.485 ;
        RECT 78.340 204.625 78.510 205.730 ;
        RECT 78.680 204.945 78.920 205.540 ;
        RECT 79.090 205.475 79.620 205.840 ;
        RECT 79.090 204.775 79.260 205.475 ;
        RECT 79.790 205.395 79.960 206.010 ;
        RECT 80.130 205.655 80.300 206.455 ;
        RECT 80.470 205.955 80.720 206.285 ;
        RECT 80.945 205.985 81.830 206.155 ;
        RECT 79.790 205.305 80.300 205.395 ;
        RECT 78.340 204.495 78.565 204.625 ;
        RECT 78.735 204.555 79.260 204.775 ;
        RECT 79.430 205.135 80.300 205.305 ;
        RECT 77.975 203.905 78.225 204.365 ;
        RECT 78.395 204.355 78.565 204.495 ;
        RECT 79.430 204.355 79.600 205.135 ;
        RECT 80.130 205.065 80.300 205.135 ;
        RECT 79.810 204.885 80.010 204.915 ;
        RECT 80.470 204.885 80.640 205.955 ;
        RECT 80.810 205.065 81.000 205.785 ;
        RECT 79.810 204.585 80.640 204.885 ;
        RECT 81.170 204.855 81.490 205.815 ;
        RECT 78.395 204.185 78.730 204.355 ;
        RECT 78.925 204.185 79.600 204.355 ;
        RECT 79.920 203.905 80.290 204.405 ;
        RECT 80.470 204.355 80.640 204.585 ;
        RECT 81.025 204.525 81.490 204.855 ;
        RECT 81.660 205.145 81.830 205.985 ;
        RECT 82.010 205.955 82.325 206.455 ;
        RECT 82.555 205.725 82.895 206.285 ;
        RECT 82.000 205.350 82.895 205.725 ;
        RECT 83.065 205.445 83.235 206.455 ;
        RECT 82.705 205.145 82.895 205.350 ;
        RECT 83.405 205.395 83.735 206.240 ;
        RECT 83.405 205.315 83.795 205.395 ;
        RECT 83.965 205.365 85.175 206.455 ;
        RECT 83.580 205.265 83.795 205.315 ;
        RECT 81.660 204.815 82.535 205.145 ;
        RECT 82.705 204.815 83.455 205.145 ;
        RECT 81.660 204.355 81.830 204.815 ;
        RECT 82.705 204.645 82.905 204.815 ;
        RECT 83.625 204.685 83.795 205.265 ;
        RECT 83.570 204.645 83.795 204.685 ;
        RECT 80.470 204.185 80.875 204.355 ;
        RECT 81.045 204.185 81.830 204.355 ;
        RECT 82.105 203.905 82.315 204.435 ;
        RECT 82.575 204.120 82.905 204.645 ;
        RECT 83.415 204.560 83.795 204.645 ;
        RECT 83.965 204.655 84.485 205.195 ;
        RECT 84.655 204.825 85.175 205.365 ;
        RECT 85.435 205.525 85.605 206.285 ;
        RECT 85.820 205.695 86.150 206.455 ;
        RECT 85.435 205.355 86.150 205.525 ;
        RECT 86.320 205.380 86.575 206.285 ;
        RECT 85.345 204.805 85.700 205.175 ;
        RECT 85.980 205.145 86.150 205.355 ;
        RECT 85.980 204.815 86.235 205.145 ;
        RECT 83.075 203.905 83.245 204.515 ;
        RECT 83.415 204.125 83.745 204.560 ;
        RECT 83.965 203.905 85.175 204.655 ;
        RECT 85.980 204.625 86.150 204.815 ;
        RECT 86.405 204.650 86.575 205.380 ;
        RECT 86.750 205.305 87.010 206.455 ;
        RECT 87.185 205.290 87.475 206.455 ;
        RECT 87.645 205.380 87.915 206.285 ;
        RECT 88.085 205.695 88.415 206.455 ;
        RECT 88.595 205.525 88.765 206.285 ;
        RECT 85.435 204.455 86.150 204.625 ;
        RECT 85.435 204.075 85.605 204.455 ;
        RECT 85.820 203.905 86.150 204.285 ;
        RECT 86.320 204.075 86.575 204.650 ;
        RECT 86.750 203.905 87.010 204.745 ;
        RECT 87.185 203.905 87.475 204.630 ;
        RECT 87.645 204.580 87.815 205.380 ;
        RECT 88.100 205.355 88.765 205.525 ;
        RECT 89.545 205.395 89.875 206.240 ;
        RECT 90.045 205.445 90.215 206.455 ;
        RECT 90.385 205.725 90.725 206.285 ;
        RECT 90.955 205.955 91.270 206.455 ;
        RECT 91.450 205.985 92.335 206.155 ;
        RECT 88.100 205.210 88.270 205.355 ;
        RECT 87.985 204.880 88.270 205.210 ;
        RECT 89.485 205.315 89.875 205.395 ;
        RECT 90.385 205.350 91.280 205.725 ;
        RECT 89.485 205.265 89.700 205.315 ;
        RECT 88.100 204.625 88.270 204.880 ;
        RECT 88.505 204.805 88.835 205.175 ;
        RECT 89.485 204.685 89.655 205.265 ;
        RECT 90.385 205.145 90.575 205.350 ;
        RECT 91.450 205.145 91.620 205.985 ;
        RECT 92.560 205.955 92.810 206.285 ;
        RECT 89.825 204.815 90.575 205.145 ;
        RECT 90.745 204.815 91.620 205.145 ;
        RECT 89.485 204.645 89.710 204.685 ;
        RECT 90.375 204.645 90.575 204.815 ;
        RECT 87.645 204.075 87.905 204.580 ;
        RECT 88.100 204.455 88.765 204.625 ;
        RECT 89.485 204.560 89.865 204.645 ;
        RECT 88.085 203.905 88.415 204.285 ;
        RECT 88.595 204.075 88.765 204.455 ;
        RECT 89.535 204.125 89.865 204.560 ;
        RECT 90.035 203.905 90.205 204.515 ;
        RECT 90.375 204.120 90.705 204.645 ;
        RECT 90.965 203.905 91.175 204.435 ;
        RECT 91.450 204.355 91.620 204.815 ;
        RECT 91.790 204.855 92.110 205.815 ;
        RECT 92.280 205.065 92.470 205.785 ;
        RECT 92.640 204.885 92.810 205.955 ;
        RECT 92.980 205.655 93.150 206.455 ;
        RECT 93.320 206.010 94.425 206.180 ;
        RECT 93.320 205.395 93.490 206.010 ;
        RECT 94.635 205.860 94.885 206.285 ;
        RECT 95.055 205.995 95.320 206.455 ;
        RECT 93.660 205.475 94.190 205.840 ;
        RECT 94.635 205.730 94.940 205.860 ;
        RECT 92.980 205.305 93.490 205.395 ;
        RECT 92.980 205.135 93.850 205.305 ;
        RECT 92.980 205.065 93.150 205.135 ;
        RECT 93.270 204.885 93.470 204.915 ;
        RECT 91.790 204.525 92.255 204.855 ;
        RECT 92.640 204.585 93.470 204.885 ;
        RECT 92.640 204.355 92.810 204.585 ;
        RECT 91.450 204.185 92.235 204.355 ;
        RECT 92.405 204.185 92.810 204.355 ;
        RECT 92.990 203.905 93.360 204.405 ;
        RECT 93.680 204.355 93.850 205.135 ;
        RECT 94.020 204.775 94.190 205.475 ;
        RECT 94.360 204.945 94.600 205.540 ;
        RECT 94.020 204.555 94.545 204.775 ;
        RECT 94.770 204.625 94.940 205.730 ;
        RECT 94.715 204.495 94.940 204.625 ;
        RECT 95.110 204.535 95.390 205.485 ;
        RECT 94.715 204.355 94.885 204.495 ;
        RECT 93.680 204.185 94.355 204.355 ;
        RECT 94.550 204.185 94.885 204.355 ;
        RECT 95.055 203.905 95.305 204.365 ;
        RECT 95.560 204.165 95.745 206.285 ;
        RECT 95.915 205.955 96.245 206.455 ;
        RECT 96.415 205.785 96.585 206.285 ;
        RECT 95.920 205.615 96.585 205.785 ;
        RECT 95.920 204.625 96.150 205.615 ;
        RECT 96.320 204.795 96.670 205.445 ;
        RECT 96.845 205.380 97.115 206.285 ;
        RECT 97.285 205.695 97.615 206.455 ;
        RECT 97.795 205.525 97.965 206.285 ;
        RECT 95.920 204.455 96.585 204.625 ;
        RECT 95.915 203.905 96.245 204.285 ;
        RECT 96.415 204.165 96.585 204.455 ;
        RECT 96.845 204.580 97.015 205.380 ;
        RECT 97.300 205.355 97.965 205.525 ;
        RECT 98.775 205.525 98.945 206.285 ;
        RECT 99.125 205.695 99.455 206.455 ;
        RECT 98.775 205.355 99.440 205.525 ;
        RECT 99.625 205.380 99.895 206.285 ;
        RECT 100.125 205.395 100.455 206.240 ;
        RECT 100.625 205.445 100.795 206.455 ;
        RECT 100.965 205.725 101.305 206.285 ;
        RECT 101.535 205.955 101.850 206.455 ;
        RECT 102.030 205.985 102.915 206.155 ;
        RECT 97.300 205.210 97.470 205.355 ;
        RECT 97.185 204.880 97.470 205.210 ;
        RECT 99.270 205.210 99.440 205.355 ;
        RECT 97.300 204.625 97.470 204.880 ;
        RECT 97.705 204.805 98.035 205.175 ;
        RECT 98.705 204.805 99.035 205.175 ;
        RECT 99.270 204.880 99.555 205.210 ;
        RECT 99.270 204.625 99.440 204.880 ;
        RECT 96.845 204.075 97.105 204.580 ;
        RECT 97.300 204.455 97.965 204.625 ;
        RECT 97.285 203.905 97.615 204.285 ;
        RECT 97.795 204.075 97.965 204.455 ;
        RECT 98.775 204.455 99.440 204.625 ;
        RECT 99.725 204.580 99.895 205.380 ;
        RECT 98.775 204.075 98.945 204.455 ;
        RECT 99.125 203.905 99.455 204.285 ;
        RECT 99.635 204.075 99.895 204.580 ;
        RECT 100.065 205.315 100.455 205.395 ;
        RECT 100.965 205.350 101.860 205.725 ;
        RECT 100.065 205.265 100.280 205.315 ;
        RECT 100.065 204.685 100.235 205.265 ;
        RECT 100.965 205.145 101.155 205.350 ;
        RECT 102.030 205.145 102.200 205.985 ;
        RECT 103.140 205.955 103.390 206.285 ;
        RECT 100.405 204.815 101.155 205.145 ;
        RECT 101.325 204.815 102.200 205.145 ;
        RECT 100.065 204.645 100.290 204.685 ;
        RECT 100.955 204.645 101.155 204.815 ;
        RECT 100.065 204.560 100.445 204.645 ;
        RECT 100.115 204.125 100.445 204.560 ;
        RECT 100.615 203.905 100.785 204.515 ;
        RECT 100.955 204.120 101.285 204.645 ;
        RECT 101.545 203.905 101.755 204.435 ;
        RECT 102.030 204.355 102.200 204.815 ;
        RECT 102.370 204.855 102.690 205.815 ;
        RECT 102.860 205.065 103.050 205.785 ;
        RECT 103.220 204.885 103.390 205.955 ;
        RECT 103.560 205.655 103.730 206.455 ;
        RECT 103.900 206.010 105.005 206.180 ;
        RECT 103.900 205.395 104.070 206.010 ;
        RECT 105.215 205.860 105.465 206.285 ;
        RECT 105.635 205.995 105.900 206.455 ;
        RECT 104.240 205.475 104.770 205.840 ;
        RECT 105.215 205.730 105.520 205.860 ;
        RECT 103.560 205.305 104.070 205.395 ;
        RECT 103.560 205.135 104.430 205.305 ;
        RECT 103.560 205.065 103.730 205.135 ;
        RECT 103.850 204.885 104.050 204.915 ;
        RECT 102.370 204.525 102.835 204.855 ;
        RECT 103.220 204.585 104.050 204.885 ;
        RECT 103.220 204.355 103.390 204.585 ;
        RECT 102.030 204.185 102.815 204.355 ;
        RECT 102.985 204.185 103.390 204.355 ;
        RECT 103.570 203.905 103.940 204.405 ;
        RECT 104.260 204.355 104.430 205.135 ;
        RECT 104.600 204.775 104.770 205.475 ;
        RECT 104.940 204.945 105.180 205.540 ;
        RECT 104.600 204.555 105.125 204.775 ;
        RECT 105.350 204.625 105.520 205.730 ;
        RECT 105.295 204.495 105.520 204.625 ;
        RECT 105.690 204.535 105.970 205.485 ;
        RECT 105.295 204.355 105.465 204.495 ;
        RECT 104.260 204.185 104.935 204.355 ;
        RECT 105.130 204.185 105.465 204.355 ;
        RECT 105.635 203.905 105.885 204.365 ;
        RECT 106.140 204.165 106.325 206.285 ;
        RECT 106.495 205.955 106.825 206.455 ;
        RECT 106.995 205.785 107.165 206.285 ;
        RECT 106.500 205.615 107.165 205.785 ;
        RECT 106.500 204.625 106.730 205.615 ;
        RECT 106.900 204.795 107.250 205.445 ;
        RECT 107.425 205.365 109.095 206.455 ;
        RECT 107.425 204.675 108.175 205.195 ;
        RECT 108.345 204.845 109.095 205.365 ;
        RECT 109.265 205.315 109.650 206.285 ;
        RECT 109.820 205.995 110.145 206.455 ;
        RECT 110.665 205.825 110.945 206.285 ;
        RECT 109.820 205.605 110.945 205.825 ;
        RECT 106.500 204.455 107.165 204.625 ;
        RECT 106.495 203.905 106.825 204.285 ;
        RECT 106.995 204.165 107.165 204.455 ;
        RECT 107.425 203.905 109.095 204.675 ;
        RECT 109.265 204.645 109.545 205.315 ;
        RECT 109.820 205.145 110.270 205.605 ;
        RECT 111.135 205.435 111.535 206.285 ;
        RECT 111.935 205.995 112.205 206.455 ;
        RECT 112.375 205.825 112.660 206.285 ;
        RECT 109.715 204.815 110.270 205.145 ;
        RECT 110.440 204.875 111.535 205.435 ;
        RECT 109.820 204.705 110.270 204.815 ;
        RECT 109.265 204.075 109.650 204.645 ;
        RECT 109.820 204.535 110.945 204.705 ;
        RECT 109.820 203.905 110.145 204.365 ;
        RECT 110.665 204.075 110.945 204.535 ;
        RECT 111.135 204.075 111.535 204.875 ;
        RECT 111.705 205.605 112.660 205.825 ;
        RECT 111.705 204.705 111.915 205.605 ;
        RECT 112.085 204.875 112.775 205.435 ;
        RECT 112.945 205.290 113.235 206.455 ;
        RECT 114.415 205.785 114.585 206.285 ;
        RECT 114.755 205.955 115.085 206.455 ;
        RECT 114.415 205.615 115.080 205.785 ;
        RECT 114.330 204.795 114.680 205.445 ;
        RECT 111.705 204.535 112.660 204.705 ;
        RECT 111.935 203.905 112.205 204.365 ;
        RECT 112.375 204.075 112.660 204.535 ;
        RECT 112.945 203.905 113.235 204.630 ;
        RECT 114.850 204.625 115.080 205.615 ;
        RECT 114.415 204.455 115.080 204.625 ;
        RECT 114.415 204.165 114.585 204.455 ;
        RECT 114.755 203.905 115.085 204.285 ;
        RECT 115.255 204.165 115.440 206.285 ;
        RECT 115.680 205.995 115.945 206.455 ;
        RECT 116.115 205.860 116.365 206.285 ;
        RECT 116.575 206.010 117.680 206.180 ;
        RECT 116.060 205.730 116.365 205.860 ;
        RECT 115.610 204.535 115.890 205.485 ;
        RECT 116.060 204.625 116.230 205.730 ;
        RECT 116.400 204.945 116.640 205.540 ;
        RECT 116.810 205.475 117.340 205.840 ;
        RECT 116.810 204.775 116.980 205.475 ;
        RECT 117.510 205.395 117.680 206.010 ;
        RECT 117.850 205.655 118.020 206.455 ;
        RECT 118.190 205.955 118.440 206.285 ;
        RECT 118.665 205.985 119.550 206.155 ;
        RECT 117.510 205.305 118.020 205.395 ;
        RECT 116.060 204.495 116.285 204.625 ;
        RECT 116.455 204.555 116.980 204.775 ;
        RECT 117.150 205.135 118.020 205.305 ;
        RECT 115.695 203.905 115.945 204.365 ;
        RECT 116.115 204.355 116.285 204.495 ;
        RECT 117.150 204.355 117.320 205.135 ;
        RECT 117.850 205.065 118.020 205.135 ;
        RECT 117.530 204.885 117.730 204.915 ;
        RECT 118.190 204.885 118.360 205.955 ;
        RECT 118.530 205.065 118.720 205.785 ;
        RECT 117.530 204.585 118.360 204.885 ;
        RECT 118.890 204.855 119.210 205.815 ;
        RECT 116.115 204.185 116.450 204.355 ;
        RECT 116.645 204.185 117.320 204.355 ;
        RECT 117.640 203.905 118.010 204.405 ;
        RECT 118.190 204.355 118.360 204.585 ;
        RECT 118.745 204.525 119.210 204.855 ;
        RECT 119.380 205.145 119.550 205.985 ;
        RECT 119.730 205.955 120.045 206.455 ;
        RECT 120.275 205.725 120.615 206.285 ;
        RECT 119.720 205.350 120.615 205.725 ;
        RECT 120.785 205.445 120.955 206.455 ;
        RECT 120.425 205.145 120.615 205.350 ;
        RECT 121.125 205.395 121.455 206.240 ;
        RECT 121.685 205.605 122.065 206.285 ;
        RECT 122.655 205.605 122.825 206.455 ;
        RECT 122.995 205.775 123.325 206.285 ;
        RECT 123.495 205.945 123.665 206.455 ;
        RECT 123.835 205.775 124.235 206.285 ;
        RECT 122.995 205.605 124.235 205.775 ;
        RECT 121.125 205.315 121.515 205.395 ;
        RECT 121.300 205.265 121.515 205.315 ;
        RECT 119.380 204.815 120.255 205.145 ;
        RECT 120.425 204.815 121.175 205.145 ;
        RECT 119.380 204.355 119.550 204.815 ;
        RECT 120.425 204.645 120.625 204.815 ;
        RECT 121.345 204.685 121.515 205.265 ;
        RECT 121.290 204.645 121.515 204.685 ;
        RECT 118.190 204.185 118.595 204.355 ;
        RECT 118.765 204.185 119.550 204.355 ;
        RECT 119.825 203.905 120.035 204.435 ;
        RECT 120.295 204.120 120.625 204.645 ;
        RECT 121.135 204.560 121.515 204.645 ;
        RECT 121.685 204.645 121.855 205.605 ;
        RECT 122.025 205.265 123.330 205.435 ;
        RECT 124.415 205.355 124.735 206.285 ;
        RECT 122.025 204.815 122.270 205.265 ;
        RECT 122.440 204.895 122.990 205.095 ;
        RECT 123.160 205.065 123.330 205.265 ;
        RECT 124.105 205.185 124.735 205.355 ;
        RECT 124.925 205.400 125.230 206.185 ;
        RECT 125.410 205.985 126.095 206.455 ;
        RECT 125.405 205.465 126.100 205.775 ;
        RECT 123.160 204.895 123.535 205.065 ;
        RECT 123.705 204.645 123.935 205.145 ;
        RECT 120.795 203.905 120.965 204.515 ;
        RECT 121.135 204.125 121.465 204.560 ;
        RECT 121.685 204.475 123.935 204.645 ;
        RECT 121.735 203.905 122.065 204.295 ;
        RECT 122.235 204.155 122.405 204.475 ;
        RECT 124.105 204.305 124.275 205.185 ;
        RECT 122.575 203.905 122.905 204.295 ;
        RECT 123.320 204.135 124.275 204.305 ;
        RECT 124.445 203.905 124.735 204.740 ;
        RECT 124.925 204.595 125.100 205.400 ;
        RECT 126.275 205.295 126.560 206.240 ;
        RECT 126.735 206.005 127.065 206.455 ;
        RECT 127.235 205.835 127.405 206.265 ;
        RECT 125.700 205.145 126.560 205.295 ;
        RECT 125.275 205.125 126.560 205.145 ;
        RECT 126.730 205.605 127.405 205.835 ;
        RECT 127.755 205.835 127.925 206.265 ;
        RECT 128.095 206.005 128.425 206.455 ;
        RECT 127.755 205.605 128.430 205.835 ;
        RECT 125.275 204.765 126.260 205.125 ;
        RECT 126.730 204.955 126.965 205.605 ;
        RECT 124.925 204.075 125.165 204.595 ;
        RECT 126.090 204.430 126.260 204.765 ;
        RECT 126.430 204.625 126.965 204.955 ;
        RECT 126.745 204.475 126.965 204.625 ;
        RECT 127.135 204.585 127.435 205.435 ;
        RECT 127.725 204.585 128.025 205.435 ;
        RECT 128.195 204.955 128.430 205.605 ;
        RECT 128.600 205.295 128.885 206.240 ;
        RECT 129.065 205.985 129.750 206.455 ;
        RECT 129.060 205.465 129.755 205.775 ;
        RECT 129.930 205.400 130.235 206.185 ;
        RECT 131.435 205.785 131.605 206.285 ;
        RECT 131.775 205.955 132.105 206.455 ;
        RECT 131.435 205.615 132.100 205.785 ;
        RECT 128.600 205.145 129.460 205.295 ;
        RECT 128.600 205.125 129.885 205.145 ;
        RECT 128.195 204.625 128.730 204.955 ;
        RECT 128.900 204.765 129.885 205.125 ;
        RECT 128.195 204.475 128.415 204.625 ;
        RECT 125.335 203.905 125.730 204.400 ;
        RECT 126.090 204.235 126.465 204.430 ;
        RECT 126.295 204.090 126.465 204.235 ;
        RECT 126.745 204.100 126.985 204.475 ;
        RECT 127.155 203.905 127.490 204.410 ;
        RECT 127.670 203.905 128.005 204.410 ;
        RECT 128.175 204.100 128.415 204.475 ;
        RECT 128.900 204.430 129.070 204.765 ;
        RECT 130.060 204.595 130.235 205.400 ;
        RECT 131.350 204.795 131.700 205.445 ;
        RECT 131.870 204.625 132.100 205.615 ;
        RECT 128.695 204.235 129.070 204.430 ;
        RECT 128.695 204.090 128.865 204.235 ;
        RECT 129.430 203.905 129.825 204.400 ;
        RECT 129.995 204.075 130.235 204.595 ;
        RECT 131.435 204.455 132.100 204.625 ;
        RECT 131.435 204.165 131.605 204.455 ;
        RECT 131.775 203.905 132.105 204.285 ;
        RECT 132.275 204.165 132.460 206.285 ;
        RECT 132.700 205.995 132.965 206.455 ;
        RECT 133.135 205.860 133.385 206.285 ;
        RECT 133.595 206.010 134.700 206.180 ;
        RECT 133.080 205.730 133.385 205.860 ;
        RECT 132.630 204.535 132.910 205.485 ;
        RECT 133.080 204.625 133.250 205.730 ;
        RECT 133.420 204.945 133.660 205.540 ;
        RECT 133.830 205.475 134.360 205.840 ;
        RECT 133.830 204.775 134.000 205.475 ;
        RECT 134.530 205.395 134.700 206.010 ;
        RECT 134.870 205.655 135.040 206.455 ;
        RECT 135.210 205.955 135.460 206.285 ;
        RECT 135.685 205.985 136.570 206.155 ;
        RECT 134.530 205.305 135.040 205.395 ;
        RECT 133.080 204.495 133.305 204.625 ;
        RECT 133.475 204.555 134.000 204.775 ;
        RECT 134.170 205.135 135.040 205.305 ;
        RECT 132.715 203.905 132.965 204.365 ;
        RECT 133.135 204.355 133.305 204.495 ;
        RECT 134.170 204.355 134.340 205.135 ;
        RECT 134.870 205.065 135.040 205.135 ;
        RECT 134.550 204.885 134.750 204.915 ;
        RECT 135.210 204.885 135.380 205.955 ;
        RECT 135.550 205.065 135.740 205.785 ;
        RECT 134.550 204.585 135.380 204.885 ;
        RECT 135.910 204.855 136.230 205.815 ;
        RECT 133.135 204.185 133.470 204.355 ;
        RECT 133.665 204.185 134.340 204.355 ;
        RECT 134.660 203.905 135.030 204.405 ;
        RECT 135.210 204.355 135.380 204.585 ;
        RECT 135.765 204.525 136.230 204.855 ;
        RECT 136.400 205.145 136.570 205.985 ;
        RECT 136.750 205.955 137.065 206.455 ;
        RECT 137.295 205.725 137.635 206.285 ;
        RECT 136.740 205.350 137.635 205.725 ;
        RECT 137.805 205.445 137.975 206.455 ;
        RECT 137.445 205.145 137.635 205.350 ;
        RECT 138.145 205.395 138.475 206.240 ;
        RECT 138.145 205.315 138.535 205.395 ;
        RECT 138.320 205.265 138.535 205.315 ;
        RECT 138.705 205.290 138.995 206.455 ;
        RECT 139.255 205.525 139.425 206.285 ;
        RECT 139.605 205.695 139.935 206.455 ;
        RECT 139.255 205.355 139.920 205.525 ;
        RECT 140.105 205.380 140.375 206.285 ;
        RECT 140.605 205.395 140.935 206.240 ;
        RECT 141.105 205.445 141.275 206.455 ;
        RECT 141.445 205.725 141.785 206.285 ;
        RECT 142.015 205.955 142.330 206.455 ;
        RECT 142.510 205.985 143.395 206.155 ;
        RECT 136.400 204.815 137.275 205.145 ;
        RECT 137.445 204.815 138.195 205.145 ;
        RECT 136.400 204.355 136.570 204.815 ;
        RECT 137.445 204.645 137.645 204.815 ;
        RECT 138.365 204.685 138.535 205.265 ;
        RECT 139.750 205.210 139.920 205.355 ;
        RECT 139.185 204.805 139.515 205.175 ;
        RECT 139.750 204.880 140.035 205.210 ;
        RECT 138.310 204.645 138.535 204.685 ;
        RECT 135.210 204.185 135.615 204.355 ;
        RECT 135.785 204.185 136.570 204.355 ;
        RECT 136.845 203.905 137.055 204.435 ;
        RECT 137.315 204.120 137.645 204.645 ;
        RECT 138.155 204.560 138.535 204.645 ;
        RECT 137.815 203.905 137.985 204.515 ;
        RECT 138.155 204.125 138.485 204.560 ;
        RECT 138.705 203.905 138.995 204.630 ;
        RECT 139.750 204.625 139.920 204.880 ;
        RECT 139.255 204.455 139.920 204.625 ;
        RECT 140.205 204.580 140.375 205.380 ;
        RECT 139.255 204.075 139.425 204.455 ;
        RECT 139.605 203.905 139.935 204.285 ;
        RECT 140.115 204.075 140.375 204.580 ;
        RECT 140.545 205.315 140.935 205.395 ;
        RECT 141.445 205.350 142.340 205.725 ;
        RECT 140.545 205.265 140.760 205.315 ;
        RECT 140.545 204.685 140.715 205.265 ;
        RECT 141.445 205.145 141.635 205.350 ;
        RECT 142.510 205.145 142.680 205.985 ;
        RECT 143.620 205.955 143.870 206.285 ;
        RECT 140.885 204.815 141.635 205.145 ;
        RECT 141.805 204.815 142.680 205.145 ;
        RECT 140.545 204.645 140.770 204.685 ;
        RECT 141.435 204.645 141.635 204.815 ;
        RECT 140.545 204.560 140.925 204.645 ;
        RECT 140.595 204.125 140.925 204.560 ;
        RECT 141.095 203.905 141.265 204.515 ;
        RECT 141.435 204.120 141.765 204.645 ;
        RECT 142.025 203.905 142.235 204.435 ;
        RECT 142.510 204.355 142.680 204.815 ;
        RECT 142.850 204.855 143.170 205.815 ;
        RECT 143.340 205.065 143.530 205.785 ;
        RECT 143.700 204.885 143.870 205.955 ;
        RECT 144.040 205.655 144.210 206.455 ;
        RECT 144.380 206.010 145.485 206.180 ;
        RECT 144.380 205.395 144.550 206.010 ;
        RECT 145.695 205.860 145.945 206.285 ;
        RECT 146.115 205.995 146.380 206.455 ;
        RECT 144.720 205.475 145.250 205.840 ;
        RECT 145.695 205.730 146.000 205.860 ;
        RECT 144.040 205.305 144.550 205.395 ;
        RECT 144.040 205.135 144.910 205.305 ;
        RECT 144.040 205.065 144.210 205.135 ;
        RECT 144.330 204.885 144.530 204.915 ;
        RECT 142.850 204.525 143.315 204.855 ;
        RECT 143.700 204.585 144.530 204.885 ;
        RECT 143.700 204.355 143.870 204.585 ;
        RECT 142.510 204.185 143.295 204.355 ;
        RECT 143.465 204.185 143.870 204.355 ;
        RECT 144.050 203.905 144.420 204.405 ;
        RECT 144.740 204.355 144.910 205.135 ;
        RECT 145.080 204.775 145.250 205.475 ;
        RECT 145.420 204.945 145.660 205.540 ;
        RECT 145.080 204.555 145.605 204.775 ;
        RECT 145.830 204.625 146.000 205.730 ;
        RECT 145.775 204.495 146.000 204.625 ;
        RECT 146.170 204.535 146.450 205.485 ;
        RECT 145.775 204.355 145.945 204.495 ;
        RECT 144.740 204.185 145.415 204.355 ;
        RECT 145.610 204.185 145.945 204.355 ;
        RECT 146.115 203.905 146.365 204.365 ;
        RECT 146.620 204.165 146.805 206.285 ;
        RECT 146.975 205.955 147.305 206.455 ;
        RECT 147.475 205.785 147.645 206.285 ;
        RECT 147.905 206.020 153.250 206.455 ;
        RECT 146.980 205.615 147.645 205.785 ;
        RECT 146.980 204.625 147.210 205.615 ;
        RECT 147.380 204.795 147.730 205.445 ;
        RECT 146.980 204.455 147.645 204.625 ;
        RECT 146.975 203.905 147.305 204.285 ;
        RECT 147.475 204.165 147.645 204.455 ;
        RECT 149.490 204.450 149.830 205.280 ;
        RECT 151.310 204.770 151.660 206.020 ;
        RECT 153.425 205.365 155.095 206.455 ;
        RECT 153.425 204.675 154.175 205.195 ;
        RECT 154.345 204.845 155.095 205.365 ;
        RECT 155.725 205.365 156.935 206.455 ;
        RECT 155.725 204.825 156.245 205.365 ;
        RECT 147.905 203.905 153.250 204.450 ;
        RECT 153.425 203.905 155.095 204.675 ;
        RECT 156.415 204.655 156.935 205.195 ;
        RECT 155.725 203.905 156.935 204.655 ;
        RECT 22.700 203.735 157.020 203.905 ;
        RECT 22.785 202.985 23.995 203.735 ;
        RECT 24.335 203.220 24.505 203.735 ;
        RECT 24.675 203.080 25.005 203.515 ;
        RECT 25.175 203.125 25.345 203.735 ;
        RECT 24.625 202.995 25.005 203.080 ;
        RECT 25.515 202.995 25.845 203.520 ;
        RECT 26.105 203.205 26.315 203.735 ;
        RECT 26.590 203.285 27.375 203.455 ;
        RECT 27.545 203.285 27.950 203.455 ;
        RECT 22.785 202.445 23.305 202.985 ;
        RECT 24.625 202.955 24.850 202.995 ;
        RECT 23.475 202.275 23.995 202.815 ;
        RECT 22.785 201.185 23.995 202.275 ;
        RECT 24.625 202.375 24.795 202.955 ;
        RECT 25.515 202.825 25.715 202.995 ;
        RECT 26.590 202.825 26.760 203.285 ;
        RECT 24.965 202.495 25.715 202.825 ;
        RECT 25.885 202.495 26.760 202.825 ;
        RECT 24.625 202.325 24.840 202.375 ;
        RECT 24.625 202.245 25.015 202.325 ;
        RECT 24.345 201.185 24.515 202.100 ;
        RECT 24.685 201.400 25.015 202.245 ;
        RECT 25.525 202.290 25.715 202.495 ;
        RECT 25.185 201.185 25.355 202.195 ;
        RECT 25.525 201.915 26.420 202.290 ;
        RECT 25.525 201.355 25.865 201.915 ;
        RECT 26.095 201.185 26.410 201.685 ;
        RECT 26.590 201.655 26.760 202.495 ;
        RECT 26.930 202.785 27.395 203.115 ;
        RECT 27.780 203.055 27.950 203.285 ;
        RECT 28.130 203.235 28.500 203.735 ;
        RECT 28.820 203.285 29.495 203.455 ;
        RECT 29.690 203.285 30.025 203.455 ;
        RECT 26.930 201.825 27.250 202.785 ;
        RECT 27.780 202.755 28.610 203.055 ;
        RECT 27.420 201.855 27.610 202.575 ;
        RECT 27.780 201.685 27.950 202.755 ;
        RECT 28.410 202.725 28.610 202.755 ;
        RECT 28.120 202.505 28.290 202.575 ;
        RECT 28.820 202.505 28.990 203.285 ;
        RECT 29.855 203.145 30.025 203.285 ;
        RECT 30.195 203.275 30.445 203.735 ;
        RECT 28.120 202.335 28.990 202.505 ;
        RECT 29.160 202.865 29.685 203.085 ;
        RECT 29.855 203.015 30.080 203.145 ;
        RECT 28.120 202.245 28.630 202.335 ;
        RECT 26.590 201.485 27.475 201.655 ;
        RECT 27.700 201.355 27.950 201.685 ;
        RECT 28.120 201.185 28.290 201.985 ;
        RECT 28.460 201.630 28.630 202.245 ;
        RECT 29.160 202.165 29.330 202.865 ;
        RECT 28.800 201.800 29.330 202.165 ;
        RECT 29.500 202.100 29.740 202.695 ;
        RECT 29.910 201.910 30.080 203.015 ;
        RECT 30.250 202.155 30.530 203.105 ;
        RECT 29.775 201.780 30.080 201.910 ;
        RECT 28.460 201.460 29.565 201.630 ;
        RECT 29.775 201.355 30.025 201.780 ;
        RECT 30.195 201.185 30.460 201.645 ;
        RECT 30.700 201.355 30.885 203.475 ;
        RECT 31.055 203.355 31.385 203.735 ;
        RECT 31.555 203.185 31.725 203.475 ;
        RECT 31.060 203.015 31.725 203.185 ;
        RECT 31.060 202.025 31.290 203.015 ;
        RECT 31.460 202.195 31.810 202.845 ;
        RECT 31.060 201.855 31.725 202.025 ;
        RECT 31.055 201.185 31.385 201.685 ;
        RECT 31.555 201.355 31.725 201.855 ;
        RECT 32.905 201.355 33.655 203.565 ;
        RECT 33.825 202.965 37.335 203.735 ;
        RECT 37.505 202.985 38.715 203.735 ;
        RECT 33.825 202.445 35.475 202.965 ;
        RECT 35.645 202.275 37.335 202.795 ;
        RECT 37.505 202.445 38.025 202.985 ;
        RECT 38.885 202.935 39.580 203.565 ;
        RECT 39.785 202.935 40.095 203.735 ;
        RECT 40.815 203.185 40.985 203.565 ;
        RECT 41.165 203.355 41.495 203.735 ;
        RECT 40.815 203.015 41.480 203.185 ;
        RECT 41.675 203.060 41.935 203.565 ;
        RECT 42.350 203.255 42.650 203.735 ;
        RECT 42.820 203.085 43.080 203.540 ;
        RECT 43.250 203.255 43.510 203.735 ;
        RECT 43.680 203.085 43.940 203.540 ;
        RECT 44.110 203.255 44.370 203.735 ;
        RECT 44.540 203.085 44.800 203.540 ;
        RECT 44.970 203.255 45.230 203.735 ;
        RECT 45.400 203.085 45.660 203.540 ;
        RECT 45.830 203.210 46.090 203.735 ;
        RECT 38.195 202.275 38.715 202.815 ;
        RECT 38.905 202.495 39.240 202.745 ;
        RECT 39.410 202.335 39.580 202.935 ;
        RECT 39.750 202.495 40.085 202.765 ;
        RECT 40.745 202.465 41.075 202.835 ;
        RECT 41.310 202.760 41.480 203.015 ;
        RECT 41.310 202.430 41.595 202.760 ;
        RECT 33.825 201.185 37.335 202.275 ;
        RECT 37.505 201.185 38.715 202.275 ;
        RECT 38.885 201.185 39.145 202.325 ;
        RECT 39.315 201.355 39.645 202.335 ;
        RECT 39.815 201.185 40.095 202.325 ;
        RECT 41.310 202.285 41.480 202.430 ;
        RECT 40.815 202.115 41.480 202.285 ;
        RECT 41.765 202.260 41.935 203.060 ;
        RECT 40.815 201.355 40.985 202.115 ;
        RECT 41.165 201.185 41.495 201.945 ;
        RECT 41.665 201.355 41.935 202.260 ;
        RECT 42.350 202.915 45.660 203.085 ;
        RECT 42.350 202.325 43.320 202.915 ;
        RECT 46.260 202.745 46.510 203.555 ;
        RECT 46.690 203.275 46.935 203.735 ;
        RECT 43.490 202.495 46.510 202.745 ;
        RECT 46.680 202.495 46.995 203.105 ;
        RECT 47.165 202.985 48.375 203.735 ;
        RECT 48.545 203.010 48.835 203.735 ;
        RECT 49.075 203.095 49.405 203.565 ;
        RECT 49.575 203.265 49.745 203.735 ;
        RECT 49.915 203.095 50.245 203.565 ;
        RECT 50.415 203.265 50.585 203.735 ;
        RECT 50.755 203.345 52.765 203.565 ;
        RECT 52.955 203.345 54.965 203.565 ;
        RECT 50.755 203.095 51.005 203.345 ;
        RECT 42.350 202.085 45.660 202.325 ;
        RECT 42.355 201.185 42.650 201.915 ;
        RECT 42.820 201.360 43.080 202.085 ;
        RECT 43.250 201.185 43.510 201.915 ;
        RECT 43.680 201.360 43.940 202.085 ;
        RECT 44.110 201.185 44.370 201.915 ;
        RECT 44.540 201.360 44.800 202.085 ;
        RECT 44.970 201.185 45.230 201.915 ;
        RECT 45.400 201.360 45.660 202.085 ;
        RECT 45.830 201.185 46.090 202.295 ;
        RECT 46.260 201.360 46.510 202.495 ;
        RECT 47.165 202.445 47.685 202.985 ;
        RECT 49.075 202.915 51.005 203.095 ;
        RECT 51.175 202.935 54.545 203.175 ;
        RECT 46.690 201.185 46.985 202.295 ;
        RECT 47.855 202.275 48.375 202.815 ;
        RECT 49.005 202.535 50.830 202.745 ;
        RECT 51.055 202.535 52.465 202.745 ;
        RECT 52.700 202.545 54.125 202.745 ;
        RECT 54.295 202.375 54.545 202.935 ;
        RECT 54.715 203.095 54.965 203.345 ;
        RECT 55.135 203.265 55.305 203.735 ;
        RECT 55.475 203.095 55.805 203.565 ;
        RECT 55.975 203.265 56.145 203.735 ;
        RECT 56.315 203.095 56.645 203.565 ;
        RECT 54.715 202.915 56.645 203.095 ;
        RECT 56.825 202.965 59.415 203.735 ;
        RECT 60.135 203.185 60.305 203.475 ;
        RECT 60.475 203.355 60.805 203.735 ;
        RECT 60.135 203.015 60.800 203.185 ;
        RECT 54.845 202.545 56.650 202.745 ;
        RECT 56.825 202.445 58.035 202.965 ;
        RECT 47.165 201.185 48.375 202.275 ;
        RECT 48.545 201.185 48.835 202.350 ;
        RECT 49.115 202.195 53.245 202.365 ;
        RECT 49.115 201.355 49.365 202.195 ;
        RECT 49.535 201.185 49.785 202.025 ;
        RECT 49.955 201.355 50.205 202.195 ;
        RECT 50.375 201.185 50.625 202.025 ;
        RECT 50.795 201.355 51.045 202.195 ;
        RECT 51.215 201.185 51.465 202.025 ;
        RECT 51.635 201.355 51.885 202.195 ;
        RECT 52.055 201.185 52.305 202.025 ;
        RECT 52.475 201.525 53.245 202.195 ;
        RECT 53.415 202.195 56.145 202.375 ;
        RECT 53.415 201.695 53.665 202.195 ;
        RECT 53.835 201.525 54.085 202.025 ;
        RECT 54.255 201.695 54.505 202.195 ;
        RECT 54.675 201.525 54.925 202.025 ;
        RECT 55.095 201.695 55.345 202.195 ;
        RECT 55.515 201.525 55.765 202.025 ;
        RECT 55.935 201.695 56.145 202.195 ;
        RECT 56.315 201.525 56.650 202.365 ;
        RECT 58.205 202.275 59.415 202.795 ;
        RECT 52.475 201.355 56.650 201.525 ;
        RECT 56.825 201.185 59.415 202.275 ;
        RECT 60.050 202.195 60.400 202.845 ;
        RECT 60.570 202.025 60.800 203.015 ;
        RECT 60.135 201.855 60.800 202.025 ;
        RECT 60.135 201.355 60.305 201.855 ;
        RECT 60.475 201.185 60.805 201.685 ;
        RECT 60.975 201.355 61.160 203.475 ;
        RECT 61.415 203.275 61.665 203.735 ;
        RECT 61.835 203.285 62.170 203.455 ;
        RECT 62.365 203.285 63.040 203.455 ;
        RECT 61.835 203.145 62.005 203.285 ;
        RECT 61.330 202.155 61.610 203.105 ;
        RECT 61.780 203.015 62.005 203.145 ;
        RECT 61.780 201.910 61.950 203.015 ;
        RECT 62.175 202.865 62.700 203.085 ;
        RECT 62.120 202.100 62.360 202.695 ;
        RECT 62.530 202.165 62.700 202.865 ;
        RECT 62.870 202.505 63.040 203.285 ;
        RECT 63.360 203.235 63.730 203.735 ;
        RECT 63.910 203.285 64.315 203.455 ;
        RECT 64.485 203.285 65.270 203.455 ;
        RECT 63.910 203.055 64.080 203.285 ;
        RECT 63.250 202.755 64.080 203.055 ;
        RECT 64.465 202.785 64.930 203.115 ;
        RECT 63.250 202.725 63.450 202.755 ;
        RECT 63.570 202.505 63.740 202.575 ;
        RECT 62.870 202.335 63.740 202.505 ;
        RECT 63.230 202.245 63.740 202.335 ;
        RECT 61.780 201.780 62.085 201.910 ;
        RECT 62.530 201.800 63.060 202.165 ;
        RECT 61.400 201.185 61.665 201.645 ;
        RECT 61.835 201.355 62.085 201.780 ;
        RECT 63.230 201.630 63.400 202.245 ;
        RECT 62.295 201.460 63.400 201.630 ;
        RECT 63.570 201.185 63.740 201.985 ;
        RECT 63.910 201.685 64.080 202.755 ;
        RECT 64.250 201.855 64.440 202.575 ;
        RECT 64.610 201.825 64.930 202.785 ;
        RECT 65.100 202.825 65.270 203.285 ;
        RECT 65.545 203.205 65.755 203.735 ;
        RECT 66.015 202.995 66.345 203.520 ;
        RECT 66.515 203.125 66.685 203.735 ;
        RECT 66.855 203.080 67.185 203.515 ;
        RECT 66.855 202.995 67.235 203.080 ;
        RECT 66.145 202.825 66.345 202.995 ;
        RECT 67.010 202.955 67.235 202.995 ;
        RECT 65.100 202.495 65.975 202.825 ;
        RECT 66.145 202.495 66.895 202.825 ;
        RECT 63.910 201.355 64.160 201.685 ;
        RECT 65.100 201.655 65.270 202.495 ;
        RECT 66.145 202.290 66.335 202.495 ;
        RECT 67.065 202.375 67.235 202.955 ;
        RECT 67.405 202.965 69.995 203.735 ;
        RECT 70.660 202.995 71.275 203.565 ;
        RECT 71.445 203.225 71.660 203.735 ;
        RECT 71.890 203.225 72.170 203.555 ;
        RECT 72.350 203.225 72.590 203.735 ;
        RECT 67.405 202.445 68.615 202.965 ;
        RECT 67.020 202.325 67.235 202.375 ;
        RECT 65.440 201.915 66.335 202.290 ;
        RECT 66.845 202.245 67.235 202.325 ;
        RECT 68.785 202.275 69.995 202.795 ;
        RECT 64.385 201.485 65.270 201.655 ;
        RECT 65.450 201.185 65.765 201.685 ;
        RECT 65.995 201.355 66.335 201.915 ;
        RECT 66.505 201.185 66.675 202.195 ;
        RECT 66.845 201.400 67.175 202.245 ;
        RECT 67.405 201.185 69.995 202.275 ;
        RECT 70.660 201.975 70.975 202.995 ;
        RECT 71.145 202.325 71.315 202.825 ;
        RECT 71.565 202.495 71.830 203.055 ;
        RECT 72.000 202.325 72.170 203.225 ;
        RECT 72.340 202.495 72.695 203.055 ;
        RECT 72.925 202.935 73.620 203.565 ;
        RECT 73.825 202.935 74.135 203.735 ;
        RECT 74.305 203.010 74.595 203.735 ;
        RECT 74.765 202.985 75.975 203.735 ;
        RECT 72.945 202.495 73.280 202.745 ;
        RECT 73.450 202.335 73.620 202.935 ;
        RECT 73.790 202.495 74.125 202.765 ;
        RECT 74.765 202.445 75.285 202.985 ;
        RECT 71.145 202.155 72.570 202.325 ;
        RECT 70.660 201.355 71.195 201.975 ;
        RECT 71.365 201.185 71.695 201.985 ;
        RECT 72.180 201.980 72.570 202.155 ;
        RECT 72.925 201.185 73.185 202.325 ;
        RECT 73.355 201.355 73.685 202.335 ;
        RECT 73.855 201.185 74.135 202.325 ;
        RECT 74.305 201.185 74.595 202.350 ;
        RECT 75.455 202.275 75.975 202.815 ;
        RECT 74.765 201.185 75.975 202.275 ;
        RECT 76.145 201.355 76.895 203.565 ;
        RECT 77.995 203.355 78.325 203.735 ;
        RECT 78.495 203.235 78.705 203.565 ;
        RECT 78.995 203.235 79.215 203.565 ;
        RECT 78.035 202.190 78.235 203.080 ;
        RECT 78.535 202.825 78.705 203.235 ;
        RECT 78.535 202.495 78.875 202.825 ;
        RECT 78.535 201.990 78.705 202.495 ;
        RECT 79.045 202.160 79.215 203.235 ;
        RECT 78.075 201.820 78.705 201.990 ;
        RECT 78.915 201.905 79.215 202.160 ;
        RECT 79.425 202.075 79.645 203.400 ;
        RECT 79.860 202.125 80.175 203.400 ;
        RECT 80.660 203.355 80.990 203.735 ;
        RECT 81.160 203.180 81.445 203.565 ;
        RECT 81.615 203.355 81.950 203.735 ;
        RECT 80.345 202.205 80.675 203.175 ;
        RECT 81.160 202.995 81.955 203.180 ;
        RECT 80.895 202.495 81.155 202.825 ;
        RECT 80.895 202.025 81.065 202.495 ;
        RECT 81.325 202.285 81.955 202.995 ;
        RECT 82.125 202.985 83.335 203.735 ;
        RECT 83.595 203.185 83.765 203.475 ;
        RECT 83.935 203.355 84.265 203.735 ;
        RECT 83.595 203.015 84.260 203.185 ;
        RECT 82.125 202.445 82.645 202.985 ;
        RECT 80.340 201.905 81.065 202.025 ;
        RECT 78.915 201.855 81.065 201.905 ;
        RECT 81.240 202.075 81.955 202.285 ;
        RECT 82.815 202.275 83.335 202.815 ;
        RECT 78.075 201.355 78.245 201.820 ;
        RECT 78.915 201.735 80.510 201.855 ;
        RECT 78.415 201.185 78.745 201.625 ;
        RECT 78.915 201.355 79.085 201.735 ;
        RECT 79.455 201.185 80.125 201.565 ;
        RECT 80.340 201.355 80.510 201.735 ;
        RECT 80.740 201.185 81.070 201.625 ;
        RECT 81.240 201.355 81.445 202.075 ;
        RECT 81.615 201.185 81.950 201.905 ;
        RECT 82.125 201.185 83.335 202.275 ;
        RECT 83.510 202.195 83.860 202.845 ;
        RECT 84.030 202.025 84.260 203.015 ;
        RECT 83.595 201.855 84.260 202.025 ;
        RECT 83.595 201.355 83.765 201.855 ;
        RECT 83.935 201.185 84.265 201.685 ;
        RECT 84.435 201.355 84.620 203.475 ;
        RECT 84.875 203.275 85.125 203.735 ;
        RECT 85.295 203.285 85.630 203.455 ;
        RECT 85.825 203.285 86.500 203.455 ;
        RECT 85.295 203.145 85.465 203.285 ;
        RECT 84.790 202.155 85.070 203.105 ;
        RECT 85.240 203.015 85.465 203.145 ;
        RECT 85.240 201.910 85.410 203.015 ;
        RECT 85.635 202.865 86.160 203.085 ;
        RECT 85.580 202.100 85.820 202.695 ;
        RECT 85.990 202.165 86.160 202.865 ;
        RECT 86.330 202.505 86.500 203.285 ;
        RECT 86.820 203.235 87.190 203.735 ;
        RECT 87.370 203.285 87.775 203.455 ;
        RECT 87.945 203.285 88.730 203.455 ;
        RECT 87.370 203.055 87.540 203.285 ;
        RECT 86.710 202.755 87.540 203.055 ;
        RECT 87.925 202.785 88.390 203.115 ;
        RECT 86.710 202.725 86.910 202.755 ;
        RECT 87.030 202.505 87.200 202.575 ;
        RECT 86.330 202.335 87.200 202.505 ;
        RECT 86.690 202.245 87.200 202.335 ;
        RECT 85.240 201.780 85.545 201.910 ;
        RECT 85.990 201.800 86.520 202.165 ;
        RECT 84.860 201.185 85.125 201.645 ;
        RECT 85.295 201.355 85.545 201.780 ;
        RECT 86.690 201.630 86.860 202.245 ;
        RECT 85.755 201.460 86.860 201.630 ;
        RECT 87.030 201.185 87.200 201.985 ;
        RECT 87.370 201.685 87.540 202.755 ;
        RECT 87.710 201.855 87.900 202.575 ;
        RECT 88.070 201.825 88.390 202.785 ;
        RECT 88.560 202.825 88.730 203.285 ;
        RECT 89.005 203.205 89.215 203.735 ;
        RECT 89.475 202.995 89.805 203.520 ;
        RECT 89.975 203.125 90.145 203.735 ;
        RECT 90.315 203.080 90.645 203.515 ;
        RECT 91.950 203.225 92.190 203.735 ;
        RECT 92.370 203.225 92.650 203.555 ;
        RECT 92.880 203.225 93.095 203.735 ;
        RECT 90.315 202.995 90.695 203.080 ;
        RECT 89.605 202.825 89.805 202.995 ;
        RECT 90.470 202.955 90.695 202.995 ;
        RECT 88.560 202.495 89.435 202.825 ;
        RECT 89.605 202.495 90.355 202.825 ;
        RECT 87.370 201.355 87.620 201.685 ;
        RECT 88.560 201.655 88.730 202.495 ;
        RECT 89.605 202.290 89.795 202.495 ;
        RECT 90.525 202.375 90.695 202.955 ;
        RECT 91.845 202.495 92.200 203.055 ;
        RECT 90.480 202.325 90.695 202.375 ;
        RECT 92.370 202.325 92.540 203.225 ;
        RECT 92.710 202.495 92.975 203.055 ;
        RECT 93.265 202.995 93.880 203.565 ;
        RECT 93.225 202.325 93.395 202.825 ;
        RECT 88.900 201.915 89.795 202.290 ;
        RECT 90.305 202.245 90.695 202.325 ;
        RECT 87.845 201.485 88.730 201.655 ;
        RECT 88.910 201.185 89.225 201.685 ;
        RECT 89.455 201.355 89.795 201.915 ;
        RECT 89.965 201.185 90.135 202.195 ;
        RECT 90.305 201.400 90.635 202.245 ;
        RECT 91.970 202.155 93.395 202.325 ;
        RECT 91.970 201.980 92.360 202.155 ;
        RECT 92.845 201.185 93.175 201.985 ;
        RECT 93.565 201.975 93.880 202.995 ;
        RECT 94.085 202.915 94.345 203.735 ;
        RECT 94.515 202.915 94.845 203.335 ;
        RECT 95.025 203.250 95.815 203.515 ;
        RECT 94.595 202.825 94.845 202.915 ;
        RECT 93.345 201.355 93.880 201.975 ;
        RECT 94.085 201.865 94.425 202.745 ;
        RECT 94.595 202.575 95.390 202.825 ;
        RECT 94.085 201.185 94.345 201.695 ;
        RECT 94.595 201.355 94.765 202.575 ;
        RECT 95.560 202.395 95.815 203.250 ;
        RECT 95.985 203.095 96.185 203.515 ;
        RECT 96.375 203.275 96.705 203.735 ;
        RECT 95.985 202.575 96.395 203.095 ;
        RECT 96.875 203.085 97.135 203.565 ;
        RECT 96.565 202.395 96.795 202.825 ;
        RECT 95.005 202.225 96.795 202.395 ;
        RECT 95.005 201.860 95.255 202.225 ;
        RECT 95.425 201.865 95.755 202.055 ;
        RECT 95.975 201.930 96.690 202.225 ;
        RECT 96.965 202.055 97.135 203.085 ;
        RECT 95.425 201.690 95.620 201.865 ;
        RECT 95.005 201.185 95.620 201.690 ;
        RECT 95.790 201.355 96.265 201.695 ;
        RECT 96.435 201.185 96.650 201.730 ;
        RECT 96.860 201.355 97.135 202.055 ;
        RECT 97.305 203.275 97.865 203.565 ;
        RECT 98.035 203.275 98.285 203.735 ;
        RECT 97.305 201.905 97.555 203.275 ;
        RECT 98.905 203.105 99.235 203.465 ;
        RECT 97.845 202.915 99.235 203.105 ;
        RECT 100.065 203.010 100.355 203.735 ;
        RECT 100.525 203.085 100.785 203.565 ;
        RECT 100.955 203.275 101.285 203.735 ;
        RECT 101.475 203.095 101.675 203.515 ;
        RECT 97.845 202.825 98.015 202.915 ;
        RECT 97.725 202.495 98.015 202.825 ;
        RECT 98.185 202.495 98.525 202.745 ;
        RECT 98.745 202.495 99.420 202.745 ;
        RECT 97.845 202.245 98.015 202.495 ;
        RECT 97.845 202.075 98.785 202.245 ;
        RECT 99.155 202.135 99.420 202.495 ;
        RECT 97.305 201.355 97.765 201.905 ;
        RECT 97.955 201.185 98.285 201.905 ;
        RECT 98.485 201.525 98.785 202.075 ;
        RECT 98.955 201.185 99.235 201.855 ;
        RECT 100.065 201.185 100.355 202.350 ;
        RECT 100.525 202.055 100.695 203.085 ;
        RECT 100.865 202.395 101.095 202.825 ;
        RECT 101.265 202.575 101.675 203.095 ;
        RECT 101.845 203.250 102.635 203.515 ;
        RECT 101.845 202.395 102.100 203.250 ;
        RECT 102.815 202.915 103.145 203.335 ;
        RECT 103.315 202.915 103.575 203.735 ;
        RECT 103.745 203.235 104.045 203.565 ;
        RECT 104.215 203.255 104.490 203.735 ;
        RECT 102.815 202.825 103.065 202.915 ;
        RECT 102.270 202.575 103.065 202.825 ;
        RECT 100.865 202.225 102.655 202.395 ;
        RECT 100.525 201.355 100.800 202.055 ;
        RECT 100.970 201.930 101.685 202.225 ;
        RECT 101.905 201.865 102.235 202.055 ;
        RECT 101.010 201.185 101.225 201.730 ;
        RECT 101.395 201.355 101.870 201.695 ;
        RECT 102.040 201.690 102.235 201.865 ;
        RECT 102.405 201.860 102.655 202.225 ;
        RECT 102.040 201.185 102.655 201.690 ;
        RECT 102.895 201.355 103.065 202.575 ;
        RECT 103.235 201.865 103.575 202.745 ;
        RECT 103.745 202.325 103.915 203.235 ;
        RECT 104.670 203.085 104.965 203.475 ;
        RECT 105.135 203.255 105.390 203.735 ;
        RECT 105.565 203.085 105.825 203.475 ;
        RECT 105.995 203.255 106.275 203.735 ;
        RECT 106.595 203.185 106.765 203.475 ;
        RECT 106.935 203.355 107.265 203.735 ;
        RECT 104.085 202.495 104.435 203.065 ;
        RECT 104.670 202.915 106.320 203.085 ;
        RECT 106.595 203.015 107.260 203.185 ;
        RECT 104.605 202.575 105.745 202.745 ;
        RECT 104.605 202.325 104.775 202.575 ;
        RECT 105.915 202.405 106.320 202.915 ;
        RECT 103.745 202.155 104.775 202.325 ;
        RECT 105.565 202.235 106.320 202.405 ;
        RECT 103.315 201.185 103.575 201.695 ;
        RECT 103.745 201.355 104.055 202.155 ;
        RECT 105.565 201.985 105.825 202.235 ;
        RECT 106.510 202.195 106.860 202.845 ;
        RECT 104.225 201.185 104.535 201.985 ;
        RECT 104.705 201.815 105.825 201.985 ;
        RECT 104.705 201.355 104.965 201.815 ;
        RECT 105.135 201.185 105.390 201.645 ;
        RECT 105.565 201.355 105.825 201.815 ;
        RECT 105.995 201.185 106.280 202.055 ;
        RECT 107.030 202.025 107.260 203.015 ;
        RECT 106.595 201.855 107.260 202.025 ;
        RECT 106.595 201.355 106.765 201.855 ;
        RECT 106.935 201.185 107.265 201.685 ;
        RECT 107.435 201.355 107.620 203.475 ;
        RECT 107.875 203.275 108.125 203.735 ;
        RECT 108.295 203.285 108.630 203.455 ;
        RECT 108.825 203.285 109.500 203.455 ;
        RECT 108.295 203.145 108.465 203.285 ;
        RECT 107.790 202.155 108.070 203.105 ;
        RECT 108.240 203.015 108.465 203.145 ;
        RECT 108.240 201.910 108.410 203.015 ;
        RECT 108.635 202.865 109.160 203.085 ;
        RECT 108.580 202.100 108.820 202.695 ;
        RECT 108.990 202.165 109.160 202.865 ;
        RECT 109.330 202.505 109.500 203.285 ;
        RECT 109.820 203.235 110.190 203.735 ;
        RECT 110.370 203.285 110.775 203.455 ;
        RECT 110.945 203.285 111.730 203.455 ;
        RECT 110.370 203.055 110.540 203.285 ;
        RECT 109.710 202.755 110.540 203.055 ;
        RECT 110.925 202.785 111.390 203.115 ;
        RECT 109.710 202.725 109.910 202.755 ;
        RECT 110.030 202.505 110.200 202.575 ;
        RECT 109.330 202.335 110.200 202.505 ;
        RECT 109.690 202.245 110.200 202.335 ;
        RECT 108.240 201.780 108.545 201.910 ;
        RECT 108.990 201.800 109.520 202.165 ;
        RECT 107.860 201.185 108.125 201.645 ;
        RECT 108.295 201.355 108.545 201.780 ;
        RECT 109.690 201.630 109.860 202.245 ;
        RECT 108.755 201.460 109.860 201.630 ;
        RECT 110.030 201.185 110.200 201.985 ;
        RECT 110.370 201.685 110.540 202.755 ;
        RECT 110.710 201.855 110.900 202.575 ;
        RECT 111.070 201.825 111.390 202.785 ;
        RECT 111.560 202.825 111.730 203.285 ;
        RECT 112.005 203.205 112.215 203.735 ;
        RECT 112.475 202.995 112.805 203.520 ;
        RECT 112.975 203.125 113.145 203.735 ;
        RECT 113.315 203.080 113.645 203.515 ;
        RECT 113.955 203.185 114.125 203.475 ;
        RECT 114.295 203.355 114.625 203.735 ;
        RECT 113.315 202.995 113.695 203.080 ;
        RECT 113.955 203.015 114.620 203.185 ;
        RECT 112.605 202.825 112.805 202.995 ;
        RECT 113.470 202.955 113.695 202.995 ;
        RECT 111.560 202.495 112.435 202.825 ;
        RECT 112.605 202.495 113.355 202.825 ;
        RECT 110.370 201.355 110.620 201.685 ;
        RECT 111.560 201.655 111.730 202.495 ;
        RECT 112.605 202.290 112.795 202.495 ;
        RECT 113.525 202.375 113.695 202.955 ;
        RECT 113.480 202.325 113.695 202.375 ;
        RECT 111.900 201.915 112.795 202.290 ;
        RECT 113.305 202.245 113.695 202.325 ;
        RECT 110.845 201.485 111.730 201.655 ;
        RECT 111.910 201.185 112.225 201.685 ;
        RECT 112.455 201.355 112.795 201.915 ;
        RECT 112.965 201.185 113.135 202.195 ;
        RECT 113.305 201.400 113.635 202.245 ;
        RECT 113.870 202.195 114.220 202.845 ;
        RECT 114.390 202.025 114.620 203.015 ;
        RECT 113.955 201.855 114.620 202.025 ;
        RECT 113.955 201.355 114.125 201.855 ;
        RECT 114.295 201.185 114.625 201.685 ;
        RECT 114.795 201.355 114.980 203.475 ;
        RECT 115.235 203.275 115.485 203.735 ;
        RECT 115.655 203.285 115.990 203.455 ;
        RECT 116.185 203.285 116.860 203.455 ;
        RECT 115.655 203.145 115.825 203.285 ;
        RECT 115.150 202.155 115.430 203.105 ;
        RECT 115.600 203.015 115.825 203.145 ;
        RECT 115.600 201.910 115.770 203.015 ;
        RECT 115.995 202.865 116.520 203.085 ;
        RECT 115.940 202.100 116.180 202.695 ;
        RECT 116.350 202.165 116.520 202.865 ;
        RECT 116.690 202.505 116.860 203.285 ;
        RECT 117.180 203.235 117.550 203.735 ;
        RECT 117.730 203.285 118.135 203.455 ;
        RECT 118.305 203.285 119.090 203.455 ;
        RECT 117.730 203.055 117.900 203.285 ;
        RECT 117.070 202.755 117.900 203.055 ;
        RECT 118.285 202.785 118.750 203.115 ;
        RECT 117.070 202.725 117.270 202.755 ;
        RECT 117.390 202.505 117.560 202.575 ;
        RECT 116.690 202.335 117.560 202.505 ;
        RECT 117.050 202.245 117.560 202.335 ;
        RECT 115.600 201.780 115.905 201.910 ;
        RECT 116.350 201.800 116.880 202.165 ;
        RECT 115.220 201.185 115.485 201.645 ;
        RECT 115.655 201.355 115.905 201.780 ;
        RECT 117.050 201.630 117.220 202.245 ;
        RECT 116.115 201.460 117.220 201.630 ;
        RECT 117.390 201.185 117.560 201.985 ;
        RECT 117.730 201.685 117.900 202.755 ;
        RECT 118.070 201.855 118.260 202.575 ;
        RECT 118.430 201.825 118.750 202.785 ;
        RECT 118.920 202.825 119.090 203.285 ;
        RECT 119.365 203.205 119.575 203.735 ;
        RECT 119.835 202.995 120.165 203.520 ;
        RECT 120.335 203.125 120.505 203.735 ;
        RECT 120.675 203.080 121.005 203.515 ;
        RECT 120.675 202.995 121.055 203.080 ;
        RECT 119.965 202.825 120.165 202.995 ;
        RECT 120.830 202.955 121.055 202.995 ;
        RECT 118.920 202.495 119.795 202.825 ;
        RECT 119.965 202.495 120.715 202.825 ;
        RECT 117.730 201.355 117.980 201.685 ;
        RECT 118.920 201.655 119.090 202.495 ;
        RECT 119.965 202.290 120.155 202.495 ;
        RECT 120.885 202.375 121.055 202.955 ;
        RECT 120.840 202.325 121.055 202.375 ;
        RECT 119.260 201.915 120.155 202.290 ;
        RECT 120.665 202.245 121.055 202.325 ;
        RECT 121.225 202.995 121.610 203.565 ;
        RECT 121.780 203.275 122.105 203.735 ;
        RECT 122.625 203.105 122.905 203.565 ;
        RECT 121.225 202.325 121.505 202.995 ;
        RECT 121.780 202.935 122.905 203.105 ;
        RECT 121.780 202.825 122.230 202.935 ;
        RECT 121.675 202.495 122.230 202.825 ;
        RECT 123.095 202.765 123.495 203.565 ;
        RECT 123.895 203.275 124.165 203.735 ;
        RECT 124.335 203.105 124.620 203.565 ;
        RECT 118.205 201.485 119.090 201.655 ;
        RECT 119.270 201.185 119.585 201.685 ;
        RECT 119.815 201.355 120.155 201.915 ;
        RECT 120.325 201.185 120.495 202.195 ;
        RECT 120.665 201.400 120.995 202.245 ;
        RECT 121.225 201.355 121.610 202.325 ;
        RECT 121.780 202.035 122.230 202.495 ;
        RECT 122.400 202.205 123.495 202.765 ;
        RECT 121.780 201.815 122.905 202.035 ;
        RECT 121.780 201.185 122.105 201.645 ;
        RECT 122.625 201.355 122.905 201.815 ;
        RECT 123.095 201.355 123.495 202.205 ;
        RECT 123.665 202.935 124.620 203.105 ;
        RECT 125.825 203.010 126.115 203.735 ;
        RECT 126.610 203.165 126.780 203.415 ;
        RECT 126.285 202.995 126.780 203.165 ;
        RECT 127.015 202.995 127.345 203.735 ;
        RECT 127.515 203.165 127.685 203.510 ;
        RECT 127.855 203.335 128.185 203.735 ;
        RECT 128.355 203.165 128.875 203.565 ;
        RECT 127.515 202.995 128.875 203.165 ;
        RECT 129.060 203.165 129.315 203.515 ;
        RECT 129.485 203.335 129.815 203.735 ;
        RECT 129.985 203.165 130.155 203.515 ;
        RECT 130.325 203.335 130.705 203.735 ;
        RECT 129.060 202.995 130.725 203.165 ;
        RECT 130.895 203.060 131.170 203.405 ;
        RECT 131.430 203.235 131.925 203.565 ;
        RECT 123.665 202.035 123.875 202.935 ;
        RECT 124.045 202.205 124.735 202.765 ;
        RECT 123.665 201.815 124.620 202.035 ;
        RECT 123.895 201.185 124.165 201.645 ;
        RECT 124.335 201.355 124.620 201.815 ;
        RECT 125.825 201.185 126.115 202.350 ;
        RECT 126.285 202.035 126.455 202.995 ;
        RECT 126.625 202.205 126.975 202.825 ;
        RECT 127.145 202.205 127.485 202.825 ;
        RECT 127.655 202.205 127.895 202.825 ;
        RECT 128.075 202.575 128.535 202.745 ;
        RECT 128.075 202.035 128.245 202.575 ;
        RECT 128.705 202.375 128.875 202.995 ;
        RECT 130.555 202.825 130.725 202.995 ;
        RECT 129.045 202.495 129.390 202.825 ;
        RECT 129.560 202.495 130.385 202.825 ;
        RECT 130.555 202.495 130.830 202.825 ;
        RECT 126.285 201.865 128.245 202.035 ;
        RECT 127.015 201.185 127.345 201.695 ;
        RECT 128.415 201.365 128.875 202.375 ;
        RECT 129.065 202.035 129.390 202.325 ;
        RECT 129.560 202.205 129.755 202.495 ;
        RECT 130.555 202.325 130.725 202.495 ;
        RECT 131.000 202.325 131.170 203.060 ;
        RECT 130.065 202.155 130.725 202.325 ;
        RECT 130.065 202.035 130.235 202.155 ;
        RECT 129.065 201.865 130.235 202.035 ;
        RECT 129.045 201.405 130.235 201.695 ;
        RECT 130.405 201.185 130.685 201.985 ;
        RECT 130.895 201.355 131.170 202.325 ;
        RECT 131.345 201.745 131.585 203.055 ;
        RECT 131.755 202.325 131.925 203.235 ;
        RECT 132.145 202.495 132.495 203.460 ;
        RECT 132.675 202.495 132.975 203.465 ;
        RECT 133.155 202.495 133.435 203.465 ;
        RECT 133.615 202.935 133.885 203.735 ;
        RECT 134.055 203.015 134.395 203.525 ;
        RECT 133.630 202.495 133.960 202.745 ;
        RECT 133.630 202.325 133.945 202.495 ;
        RECT 131.755 202.155 133.945 202.325 ;
        RECT 131.350 201.185 131.685 201.565 ;
        RECT 131.855 201.355 132.105 202.155 ;
        RECT 132.325 201.185 132.655 201.905 ;
        RECT 132.840 201.355 133.090 202.155 ;
        RECT 133.555 201.185 133.885 201.985 ;
        RECT 134.135 201.615 134.395 203.015 ;
        RECT 134.055 201.355 134.395 201.615 ;
        RECT 134.565 203.085 134.825 203.565 ;
        RECT 134.995 203.275 135.325 203.735 ;
        RECT 135.515 203.095 135.715 203.515 ;
        RECT 134.565 202.055 134.735 203.085 ;
        RECT 134.905 202.395 135.135 202.825 ;
        RECT 135.305 202.575 135.715 203.095 ;
        RECT 135.885 203.250 136.675 203.515 ;
        RECT 135.885 202.395 136.140 203.250 ;
        RECT 136.855 202.915 137.185 203.335 ;
        RECT 137.355 202.915 137.615 203.735 ;
        RECT 137.785 202.915 138.045 203.735 ;
        RECT 138.215 202.915 138.545 203.335 ;
        RECT 138.725 203.250 139.515 203.515 ;
        RECT 136.855 202.825 137.105 202.915 ;
        RECT 136.310 202.575 137.105 202.825 ;
        RECT 138.295 202.825 138.545 202.915 ;
        RECT 134.905 202.225 136.695 202.395 ;
        RECT 134.565 201.355 134.840 202.055 ;
        RECT 135.010 201.930 135.725 202.225 ;
        RECT 135.945 201.865 136.275 202.055 ;
        RECT 135.050 201.185 135.265 201.730 ;
        RECT 135.435 201.355 135.910 201.695 ;
        RECT 136.080 201.690 136.275 201.865 ;
        RECT 136.445 201.860 136.695 202.225 ;
        RECT 136.080 201.185 136.695 201.690 ;
        RECT 136.935 201.355 137.105 202.575 ;
        RECT 137.275 201.865 137.615 202.745 ;
        RECT 137.785 201.865 138.125 202.745 ;
        RECT 138.295 202.575 139.090 202.825 ;
        RECT 137.355 201.185 137.615 201.695 ;
        RECT 137.785 201.185 138.045 201.695 ;
        RECT 138.295 201.355 138.465 202.575 ;
        RECT 139.260 202.395 139.515 203.250 ;
        RECT 139.685 203.095 139.885 203.515 ;
        RECT 140.075 203.275 140.405 203.735 ;
        RECT 139.685 202.575 140.095 203.095 ;
        RECT 140.575 203.085 140.835 203.565 ;
        RECT 140.265 202.395 140.495 202.825 ;
        RECT 138.705 202.225 140.495 202.395 ;
        RECT 138.705 201.860 138.955 202.225 ;
        RECT 139.125 201.865 139.455 202.055 ;
        RECT 139.675 201.930 140.390 202.225 ;
        RECT 140.665 202.055 140.835 203.085 ;
        RECT 141.005 202.965 142.675 203.735 ;
        RECT 142.845 202.995 143.310 203.540 ;
        RECT 141.005 202.445 141.755 202.965 ;
        RECT 141.925 202.275 142.675 202.795 ;
        RECT 139.125 201.690 139.320 201.865 ;
        RECT 138.705 201.185 139.320 201.690 ;
        RECT 139.490 201.355 139.965 201.695 ;
        RECT 140.135 201.185 140.350 201.730 ;
        RECT 140.560 201.355 140.835 202.055 ;
        RECT 141.005 201.185 142.675 202.275 ;
        RECT 142.845 202.035 143.015 202.995 ;
        RECT 143.815 202.915 143.985 203.735 ;
        RECT 144.155 203.085 144.485 203.565 ;
        RECT 144.655 203.345 145.005 203.735 ;
        RECT 145.175 203.165 145.405 203.565 ;
        RECT 144.895 203.085 145.405 203.165 ;
        RECT 144.155 202.995 145.405 203.085 ;
        RECT 145.575 202.995 145.895 203.475 ;
        RECT 146.065 203.190 151.410 203.735 ;
        RECT 144.155 202.915 145.065 202.995 ;
        RECT 143.185 202.375 143.430 202.825 ;
        RECT 143.690 202.545 144.385 202.745 ;
        RECT 144.555 202.575 145.155 202.745 ;
        RECT 144.555 202.375 144.725 202.575 ;
        RECT 145.385 202.405 145.555 202.825 ;
        RECT 143.185 202.205 144.725 202.375 ;
        RECT 144.895 202.235 145.555 202.405 ;
        RECT 144.895 202.035 145.065 202.235 ;
        RECT 145.725 202.065 145.895 202.995 ;
        RECT 147.650 202.360 147.990 203.190 ;
        RECT 151.585 203.010 151.875 203.735 ;
        RECT 152.045 202.995 152.430 203.565 ;
        RECT 152.600 203.275 152.925 203.735 ;
        RECT 153.445 203.105 153.725 203.565 ;
        RECT 142.845 201.865 145.065 202.035 ;
        RECT 145.235 201.865 145.895 202.065 ;
        RECT 142.845 201.185 143.145 201.695 ;
        RECT 143.315 201.355 143.645 201.865 ;
        RECT 145.235 201.695 145.405 201.865 ;
        RECT 143.815 201.185 144.445 201.695 ;
        RECT 145.025 201.525 145.405 201.695 ;
        RECT 145.575 201.185 145.875 201.695 ;
        RECT 149.470 201.620 149.820 202.870 ;
        RECT 146.065 201.185 151.410 201.620 ;
        RECT 151.585 201.185 151.875 202.350 ;
        RECT 152.045 202.325 152.325 202.995 ;
        RECT 152.600 202.935 153.725 203.105 ;
        RECT 152.600 202.825 153.050 202.935 ;
        RECT 152.495 202.495 153.050 202.825 ;
        RECT 153.915 202.765 154.315 203.565 ;
        RECT 154.715 203.275 154.985 203.735 ;
        RECT 155.155 203.105 155.440 203.565 ;
        RECT 152.045 201.355 152.430 202.325 ;
        RECT 152.600 202.035 153.050 202.495 ;
        RECT 153.220 202.205 154.315 202.765 ;
        RECT 152.600 201.815 153.725 202.035 ;
        RECT 152.600 201.185 152.925 201.645 ;
        RECT 153.445 201.355 153.725 201.815 ;
        RECT 153.915 201.355 154.315 202.205 ;
        RECT 154.485 202.935 155.440 203.105 ;
        RECT 155.725 202.985 156.935 203.735 ;
        RECT 154.485 202.035 154.695 202.935 ;
        RECT 154.865 202.205 155.555 202.765 ;
        RECT 155.725 202.275 156.245 202.815 ;
        RECT 156.415 202.445 156.935 202.985 ;
        RECT 154.485 201.815 155.440 202.035 ;
        RECT 154.715 201.185 154.985 201.645 ;
        RECT 155.155 201.355 155.440 201.815 ;
        RECT 155.725 201.185 156.935 202.275 ;
        RECT 22.700 201.015 157.020 201.185 ;
        RECT 22.785 199.925 23.995 201.015 ;
        RECT 24.165 200.580 29.510 201.015 ;
        RECT 29.685 200.580 35.030 201.015 ;
        RECT 22.785 199.215 23.305 199.755 ;
        RECT 23.475 199.385 23.995 199.925 ;
        RECT 22.785 198.465 23.995 199.215 ;
        RECT 25.750 199.010 26.090 199.840 ;
        RECT 27.570 199.330 27.920 200.580 ;
        RECT 31.270 199.010 31.610 199.840 ;
        RECT 33.090 199.330 33.440 200.580 ;
        RECT 35.665 199.850 35.955 201.015 ;
        RECT 36.125 199.925 37.335 201.015 ;
        RECT 37.595 200.345 37.765 200.845 ;
        RECT 37.935 200.515 38.265 201.015 ;
        RECT 37.595 200.175 38.260 200.345 ;
        RECT 36.125 199.215 36.645 199.755 ;
        RECT 36.815 199.385 37.335 199.925 ;
        RECT 37.510 199.355 37.860 200.005 ;
        RECT 24.165 198.465 29.510 199.010 ;
        RECT 29.685 198.465 35.030 199.010 ;
        RECT 35.665 198.465 35.955 199.190 ;
        RECT 36.125 198.465 37.335 199.215 ;
        RECT 38.030 199.185 38.260 200.175 ;
        RECT 37.595 199.015 38.260 199.185 ;
        RECT 37.595 198.725 37.765 199.015 ;
        RECT 37.935 198.465 38.265 198.845 ;
        RECT 38.435 198.725 38.620 200.845 ;
        RECT 38.860 200.555 39.125 201.015 ;
        RECT 39.295 200.420 39.545 200.845 ;
        RECT 39.755 200.570 40.860 200.740 ;
        RECT 39.240 200.290 39.545 200.420 ;
        RECT 38.790 199.095 39.070 200.045 ;
        RECT 39.240 199.185 39.410 200.290 ;
        RECT 39.580 199.505 39.820 200.100 ;
        RECT 39.990 200.035 40.520 200.400 ;
        RECT 39.990 199.335 40.160 200.035 ;
        RECT 40.690 199.955 40.860 200.570 ;
        RECT 41.030 200.215 41.200 201.015 ;
        RECT 41.370 200.515 41.620 200.845 ;
        RECT 41.845 200.545 42.730 200.715 ;
        RECT 40.690 199.865 41.200 199.955 ;
        RECT 39.240 199.055 39.465 199.185 ;
        RECT 39.635 199.115 40.160 199.335 ;
        RECT 40.330 199.695 41.200 199.865 ;
        RECT 38.875 198.465 39.125 198.925 ;
        RECT 39.295 198.915 39.465 199.055 ;
        RECT 40.330 198.915 40.500 199.695 ;
        RECT 41.030 199.625 41.200 199.695 ;
        RECT 40.710 199.445 40.910 199.475 ;
        RECT 41.370 199.445 41.540 200.515 ;
        RECT 41.710 199.625 41.900 200.345 ;
        RECT 40.710 199.145 41.540 199.445 ;
        RECT 42.070 199.415 42.390 200.375 ;
        RECT 39.295 198.745 39.630 198.915 ;
        RECT 39.825 198.745 40.500 198.915 ;
        RECT 40.820 198.465 41.190 198.965 ;
        RECT 41.370 198.915 41.540 199.145 ;
        RECT 41.925 199.085 42.390 199.415 ;
        RECT 42.560 199.705 42.730 200.545 ;
        RECT 42.910 200.515 43.225 201.015 ;
        RECT 43.455 200.285 43.795 200.845 ;
        RECT 42.900 199.910 43.795 200.285 ;
        RECT 43.965 200.005 44.135 201.015 ;
        RECT 43.605 199.705 43.795 199.910 ;
        RECT 44.305 199.955 44.635 200.800 ;
        RECT 44.305 199.875 44.695 199.955 ;
        RECT 44.480 199.825 44.695 199.875 ;
        RECT 42.560 199.375 43.435 199.705 ;
        RECT 43.605 199.375 44.355 199.705 ;
        RECT 42.560 198.915 42.730 199.375 ;
        RECT 43.605 199.205 43.805 199.375 ;
        RECT 44.525 199.245 44.695 199.825 ;
        RECT 44.470 199.205 44.695 199.245 ;
        RECT 41.370 198.745 41.775 198.915 ;
        RECT 41.945 198.745 42.730 198.915 ;
        RECT 43.005 198.465 43.215 198.995 ;
        RECT 43.475 198.680 43.805 199.205 ;
        RECT 44.315 199.120 44.695 199.205 ;
        RECT 43.975 198.465 44.145 199.075 ;
        RECT 44.315 198.685 44.645 199.120 ;
        RECT 44.875 198.645 45.135 200.835 ;
        RECT 45.305 200.285 45.645 201.015 ;
        RECT 45.825 200.105 46.095 200.835 ;
        RECT 45.325 199.885 46.095 200.105 ;
        RECT 46.275 200.125 46.505 200.835 ;
        RECT 46.675 200.305 47.005 201.015 ;
        RECT 47.175 200.125 47.435 200.835 ;
        RECT 47.715 200.395 47.885 200.825 ;
        RECT 48.055 200.565 48.385 201.015 ;
        RECT 47.715 200.165 48.390 200.395 ;
        RECT 46.275 199.885 47.435 200.125 ;
        RECT 45.325 199.215 45.615 199.885 ;
        RECT 45.795 199.395 46.260 199.705 ;
        RECT 46.440 199.395 46.965 199.705 ;
        RECT 45.325 199.015 46.555 199.215 ;
        RECT 45.395 198.465 46.065 198.835 ;
        RECT 46.245 198.645 46.555 199.015 ;
        RECT 46.735 198.755 46.965 199.395 ;
        RECT 47.145 199.375 47.445 199.705 ;
        RECT 47.145 198.465 47.435 199.195 ;
        RECT 47.685 199.145 47.985 199.995 ;
        RECT 48.155 199.515 48.390 200.165 ;
        RECT 48.560 199.855 48.845 200.800 ;
        RECT 49.025 200.545 49.710 201.015 ;
        RECT 49.020 200.025 49.715 200.335 ;
        RECT 49.890 199.960 50.195 200.745 ;
        RECT 48.560 199.705 49.420 199.855 ;
        RECT 48.560 199.685 49.845 199.705 ;
        RECT 48.155 199.185 48.690 199.515 ;
        RECT 48.860 199.325 49.845 199.685 ;
        RECT 48.155 199.035 48.375 199.185 ;
        RECT 47.630 198.465 47.965 198.970 ;
        RECT 48.135 198.660 48.375 199.035 ;
        RECT 48.860 198.990 49.030 199.325 ;
        RECT 50.020 199.155 50.195 199.960 ;
        RECT 50.395 200.045 50.725 200.845 ;
        RECT 50.895 200.215 51.125 201.015 ;
        RECT 51.295 200.045 51.625 200.845 ;
        RECT 50.395 199.875 51.625 200.045 ;
        RECT 51.795 199.875 52.050 201.015 ;
        RECT 52.225 200.580 57.570 201.015 ;
        RECT 50.385 199.375 50.695 199.705 ;
        RECT 48.655 198.795 49.030 198.990 ;
        RECT 48.655 198.650 48.825 198.795 ;
        RECT 49.390 198.465 49.785 198.960 ;
        RECT 49.955 198.635 50.195 199.155 ;
        RECT 50.395 198.975 50.725 199.205 ;
        RECT 50.900 199.145 51.275 199.705 ;
        RECT 51.445 198.975 51.625 199.875 ;
        RECT 51.810 199.125 52.030 199.705 ;
        RECT 53.810 199.010 54.150 199.840 ;
        RECT 55.630 199.330 55.980 200.580 ;
        RECT 57.745 199.925 61.255 201.015 ;
        RECT 57.745 199.235 59.395 199.755 ;
        RECT 59.565 199.405 61.255 199.925 ;
        RECT 61.425 199.850 61.715 201.015 ;
        RECT 61.885 200.145 62.160 200.845 ;
        RECT 62.370 200.470 62.585 201.015 ;
        RECT 62.755 200.505 63.230 200.845 ;
        RECT 63.400 200.510 64.015 201.015 ;
        RECT 63.400 200.335 63.595 200.510 ;
        RECT 50.395 198.635 51.625 198.975 ;
        RECT 51.795 198.465 52.050 198.955 ;
        RECT 52.225 198.465 57.570 199.010 ;
        RECT 57.745 198.465 61.255 199.235 ;
        RECT 61.425 198.465 61.715 199.190 ;
        RECT 61.885 199.115 62.055 200.145 ;
        RECT 62.330 199.975 63.045 200.270 ;
        RECT 63.265 200.145 63.595 200.335 ;
        RECT 63.765 199.975 64.015 200.340 ;
        RECT 62.225 199.805 64.015 199.975 ;
        RECT 62.225 199.375 62.455 199.805 ;
        RECT 61.885 198.635 62.145 199.115 ;
        RECT 62.625 199.105 63.035 199.625 ;
        RECT 62.315 198.465 62.645 198.925 ;
        RECT 62.835 198.685 63.035 199.105 ;
        RECT 63.205 198.950 63.460 199.805 ;
        RECT 64.255 199.625 64.425 200.845 ;
        RECT 64.675 200.505 64.935 201.015 ;
        RECT 63.630 199.375 64.425 199.625 ;
        RECT 64.595 199.455 64.935 200.335 ;
        RECT 65.115 200.045 65.445 200.830 ;
        RECT 65.115 199.875 65.795 200.045 ;
        RECT 65.975 199.875 66.305 201.015 ;
        RECT 66.945 199.940 67.215 200.845 ;
        RECT 67.385 200.255 67.715 201.015 ;
        RECT 67.895 200.085 68.065 200.845 ;
        RECT 65.105 199.455 65.455 199.705 ;
        RECT 64.175 199.285 64.425 199.375 ;
        RECT 63.205 198.685 63.995 198.950 ;
        RECT 64.175 198.865 64.505 199.285 ;
        RECT 64.675 198.465 64.935 199.285 ;
        RECT 65.625 199.275 65.795 199.875 ;
        RECT 65.965 199.455 66.315 199.705 ;
        RECT 65.125 198.465 65.365 199.275 ;
        RECT 65.535 198.635 65.865 199.275 ;
        RECT 66.035 198.465 66.305 199.275 ;
        RECT 66.945 199.140 67.115 199.940 ;
        RECT 67.400 199.915 68.065 200.085 ;
        RECT 68.325 199.925 69.995 201.015 ;
        RECT 67.400 199.770 67.570 199.915 ;
        RECT 67.285 199.440 67.570 199.770 ;
        RECT 67.400 199.185 67.570 199.440 ;
        RECT 67.805 199.365 68.135 199.735 ;
        RECT 68.325 199.235 69.075 199.755 ;
        RECT 69.245 199.405 69.995 199.925 ;
        RECT 70.165 199.875 70.445 201.015 ;
        RECT 70.615 199.865 70.945 200.845 ;
        RECT 71.115 199.875 71.375 201.015 ;
        RECT 71.545 199.925 74.135 201.015 ;
        RECT 70.175 199.435 70.510 199.705 ;
        RECT 70.680 199.265 70.850 199.865 ;
        RECT 71.020 199.455 71.355 199.705 ;
        RECT 66.945 198.635 67.205 199.140 ;
        RECT 67.400 199.015 68.065 199.185 ;
        RECT 67.385 198.465 67.715 198.845 ;
        RECT 67.895 198.635 68.065 199.015 ;
        RECT 68.325 198.465 69.995 199.235 ;
        RECT 70.165 198.465 70.475 199.265 ;
        RECT 70.680 198.635 71.375 199.265 ;
        RECT 71.545 199.235 72.755 199.755 ;
        RECT 72.925 199.405 74.135 199.925 ;
        RECT 74.950 200.045 75.340 200.220 ;
        RECT 75.825 200.215 76.155 201.015 ;
        RECT 76.325 200.225 76.860 200.845 ;
        RECT 74.950 199.875 76.375 200.045 ;
        RECT 71.545 198.465 74.135 199.235 ;
        RECT 74.825 199.145 75.180 199.705 ;
        RECT 75.350 198.975 75.520 199.875 ;
        RECT 75.690 199.145 75.955 199.705 ;
        RECT 76.205 199.375 76.375 199.875 ;
        RECT 76.545 199.205 76.860 200.225 ;
        RECT 77.075 200.065 77.350 200.835 ;
        RECT 77.520 200.405 77.850 200.835 ;
        RECT 78.020 200.575 78.215 201.015 ;
        RECT 78.395 200.405 78.725 200.835 ;
        RECT 78.905 200.580 84.250 201.015 ;
        RECT 77.520 200.235 78.725 200.405 ;
        RECT 77.075 199.875 77.660 200.065 ;
        RECT 77.830 199.905 78.725 200.235 ;
        RECT 74.930 198.465 75.170 198.975 ;
        RECT 75.350 198.645 75.630 198.975 ;
        RECT 75.860 198.465 76.075 198.975 ;
        RECT 76.245 198.635 76.860 199.205 ;
        RECT 77.075 199.055 77.315 199.705 ;
        RECT 77.485 199.205 77.660 199.875 ;
        RECT 77.830 199.375 78.245 199.705 ;
        RECT 78.425 199.375 78.720 199.705 ;
        RECT 77.485 199.025 77.815 199.205 ;
        RECT 77.090 198.465 77.420 198.855 ;
        RECT 77.590 198.645 77.815 199.025 ;
        RECT 78.015 198.755 78.245 199.375 ;
        RECT 78.425 198.465 78.725 199.195 ;
        RECT 80.490 199.010 80.830 199.840 ;
        RECT 82.310 199.330 82.660 200.580 ;
        RECT 85.070 200.045 85.460 200.220 ;
        RECT 85.945 200.215 86.275 201.015 ;
        RECT 86.445 200.225 86.980 200.845 ;
        RECT 85.070 199.875 86.495 200.045 ;
        RECT 84.945 199.145 85.300 199.705 ;
        RECT 78.905 198.465 84.250 199.010 ;
        RECT 85.470 198.975 85.640 199.875 ;
        RECT 85.810 199.145 86.075 199.705 ;
        RECT 86.325 199.375 86.495 199.875 ;
        RECT 86.665 199.205 86.980 200.225 ;
        RECT 87.185 199.850 87.475 201.015 ;
        RECT 87.645 200.580 92.990 201.015 ;
        RECT 85.050 198.465 85.290 198.975 ;
        RECT 85.470 198.645 85.750 198.975 ;
        RECT 85.980 198.465 86.195 198.975 ;
        RECT 86.365 198.635 86.980 199.205 ;
        RECT 87.185 198.465 87.475 199.190 ;
        RECT 89.230 199.010 89.570 199.840 ;
        RECT 91.050 199.330 91.400 200.580 ;
        RECT 93.165 199.925 95.755 201.015 ;
        RECT 93.165 199.235 94.375 199.755 ;
        RECT 94.545 199.405 95.755 199.925 ;
        RECT 96.570 200.045 96.960 200.220 ;
        RECT 97.445 200.215 97.775 201.015 ;
        RECT 97.945 200.225 98.480 200.845 ;
        RECT 96.570 199.875 97.995 200.045 ;
        RECT 87.645 198.465 92.990 199.010 ;
        RECT 93.165 198.465 95.755 199.235 ;
        RECT 96.445 199.145 96.800 199.705 ;
        RECT 96.970 198.975 97.140 199.875 ;
        RECT 97.310 199.145 97.575 199.705 ;
        RECT 97.825 199.375 97.995 199.875 ;
        RECT 98.165 199.205 98.480 200.225 ;
        RECT 98.685 199.925 100.355 201.015 ;
        RECT 100.525 200.460 101.130 201.015 ;
        RECT 101.305 200.505 101.785 200.845 ;
        RECT 101.955 200.470 102.210 201.015 ;
        RECT 100.525 200.360 101.140 200.460 ;
        RECT 100.955 200.335 101.140 200.360 ;
        RECT 96.550 198.465 96.790 198.975 ;
        RECT 96.970 198.645 97.250 198.975 ;
        RECT 97.480 198.465 97.695 198.975 ;
        RECT 97.865 198.635 98.480 199.205 ;
        RECT 98.685 199.235 99.435 199.755 ;
        RECT 99.605 199.405 100.355 199.925 ;
        RECT 100.525 199.740 100.785 200.190 ;
        RECT 100.955 200.090 101.285 200.335 ;
        RECT 101.455 200.015 102.210 200.265 ;
        RECT 102.380 200.145 102.655 200.845 ;
        RECT 101.440 199.980 102.210 200.015 ;
        RECT 101.425 199.970 102.210 199.980 ;
        RECT 101.420 199.955 102.315 199.970 ;
        RECT 101.400 199.940 102.315 199.955 ;
        RECT 101.380 199.930 102.315 199.940 ;
        RECT 101.355 199.920 102.315 199.930 ;
        RECT 101.285 199.890 102.315 199.920 ;
        RECT 101.265 199.860 102.315 199.890 ;
        RECT 101.245 199.830 102.315 199.860 ;
        RECT 101.215 199.805 102.315 199.830 ;
        RECT 101.180 199.770 102.315 199.805 ;
        RECT 101.150 199.765 102.315 199.770 ;
        RECT 101.150 199.760 101.540 199.765 ;
        RECT 101.150 199.750 101.515 199.760 ;
        RECT 101.150 199.745 101.500 199.750 ;
        RECT 101.150 199.740 101.485 199.745 ;
        RECT 100.525 199.735 101.485 199.740 ;
        RECT 100.525 199.725 101.475 199.735 ;
        RECT 100.525 199.720 101.465 199.725 ;
        RECT 100.525 199.710 101.455 199.720 ;
        RECT 100.525 199.700 101.450 199.710 ;
        RECT 100.525 199.695 101.445 199.700 ;
        RECT 100.525 199.680 101.435 199.695 ;
        RECT 100.525 199.665 101.430 199.680 ;
        RECT 100.525 199.640 101.420 199.665 ;
        RECT 100.525 199.570 101.415 199.640 ;
        RECT 98.685 198.465 100.355 199.235 ;
        RECT 100.525 199.015 101.075 199.400 ;
        RECT 101.245 198.845 101.415 199.570 ;
        RECT 100.525 198.675 101.415 198.845 ;
        RECT 101.585 199.170 101.915 199.595 ;
        RECT 102.085 199.370 102.315 199.765 ;
        RECT 101.585 198.685 101.805 199.170 ;
        RECT 102.485 199.115 102.655 200.145 ;
        RECT 102.825 199.875 103.105 201.015 ;
        RECT 103.275 199.865 103.605 200.845 ;
        RECT 103.775 199.875 104.035 201.015 ;
        RECT 104.295 200.085 104.465 200.845 ;
        RECT 104.645 200.255 104.975 201.015 ;
        RECT 104.295 199.915 104.960 200.085 ;
        RECT 105.145 199.940 105.415 200.845 ;
        RECT 105.585 200.580 110.930 201.015 ;
        RECT 102.835 199.435 103.170 199.705 ;
        RECT 103.340 199.315 103.510 199.865 ;
        RECT 104.790 199.770 104.960 199.915 ;
        RECT 103.680 199.455 104.015 199.705 ;
        RECT 104.225 199.365 104.555 199.735 ;
        RECT 104.790 199.440 105.075 199.770 ;
        RECT 103.340 199.265 103.515 199.315 ;
        RECT 101.975 198.465 102.225 199.005 ;
        RECT 102.395 198.635 102.655 199.115 ;
        RECT 102.825 198.465 103.135 199.265 ;
        RECT 103.340 198.635 104.035 199.265 ;
        RECT 104.790 199.185 104.960 199.440 ;
        RECT 104.295 199.015 104.960 199.185 ;
        RECT 105.245 199.140 105.415 199.940 ;
        RECT 104.295 198.635 104.465 199.015 ;
        RECT 104.645 198.465 104.975 198.845 ;
        RECT 105.155 198.635 105.415 199.140 ;
        RECT 107.170 199.010 107.510 199.840 ;
        RECT 108.990 199.330 109.340 200.580 ;
        RECT 111.105 199.925 112.775 201.015 ;
        RECT 111.105 199.235 111.855 199.755 ;
        RECT 112.025 199.405 112.775 199.925 ;
        RECT 112.945 199.850 113.235 201.015 ;
        RECT 113.405 200.165 113.665 200.845 ;
        RECT 113.835 200.235 114.085 201.015 ;
        RECT 114.335 200.465 114.585 200.845 ;
        RECT 114.755 200.635 115.110 201.015 ;
        RECT 116.115 200.625 116.450 200.845 ;
        RECT 115.715 200.465 115.945 200.505 ;
        RECT 114.335 200.265 115.945 200.465 ;
        RECT 114.335 200.255 115.170 200.265 ;
        RECT 115.760 200.175 115.945 200.265 ;
        RECT 105.585 198.465 110.930 199.010 ;
        RECT 111.105 198.465 112.775 199.235 ;
        RECT 112.945 198.465 113.235 199.190 ;
        RECT 113.405 198.965 113.575 200.165 ;
        RECT 115.275 200.065 115.605 200.095 ;
        RECT 113.805 200.005 115.605 200.065 ;
        RECT 116.195 200.005 116.450 200.625 ;
        RECT 113.745 199.895 116.450 200.005 ;
        RECT 116.625 199.925 120.135 201.015 ;
        RECT 113.745 199.860 113.945 199.895 ;
        RECT 113.745 199.285 113.915 199.860 ;
        RECT 115.275 199.835 116.450 199.895 ;
        RECT 114.145 199.420 114.555 199.725 ;
        RECT 114.725 199.455 115.055 199.665 ;
        RECT 113.745 199.165 114.015 199.285 ;
        RECT 113.745 199.120 114.590 199.165 ;
        RECT 113.835 198.995 114.590 199.120 ;
        RECT 114.845 199.055 115.055 199.455 ;
        RECT 115.300 199.455 115.775 199.665 ;
        RECT 115.965 199.455 116.455 199.655 ;
        RECT 115.300 199.055 115.520 199.455 ;
        RECT 116.625 199.235 118.275 199.755 ;
        RECT 118.445 199.405 120.135 199.925 ;
        RECT 120.310 199.875 120.565 201.015 ;
        RECT 120.760 200.465 121.955 200.795 ;
        RECT 120.815 199.705 120.985 200.265 ;
        RECT 121.210 200.045 121.630 200.295 ;
        RECT 122.135 200.215 122.415 201.015 ;
        RECT 121.210 199.875 122.455 200.045 ;
        RECT 122.625 199.875 122.895 200.845 ;
        RECT 123.065 199.925 125.655 201.015 ;
        RECT 126.285 200.505 127.475 200.795 ;
        RECT 122.285 199.705 122.455 199.875 ;
        RECT 122.665 199.825 122.895 199.875 ;
        RECT 120.310 199.455 120.645 199.705 ;
        RECT 120.815 199.375 121.555 199.705 ;
        RECT 122.285 199.375 122.515 199.705 ;
        RECT 120.815 199.285 121.065 199.375 ;
        RECT 113.405 198.635 113.665 198.965 ;
        RECT 114.420 198.845 114.590 198.995 ;
        RECT 113.835 198.465 114.165 198.825 ;
        RECT 114.420 198.635 115.720 198.845 ;
        RECT 115.995 198.465 116.450 199.230 ;
        RECT 116.625 198.465 120.135 199.235 ;
        RECT 120.330 199.115 121.065 199.285 ;
        RECT 122.285 199.205 122.455 199.375 ;
        RECT 120.330 198.645 120.640 199.115 ;
        RECT 121.715 199.035 122.455 199.205 ;
        RECT 122.725 199.140 122.895 199.825 ;
        RECT 120.810 198.465 121.545 198.945 ;
        RECT 121.715 198.685 121.885 199.035 ;
        RECT 122.055 198.465 122.435 198.865 ;
        RECT 122.625 198.795 122.895 199.140 ;
        RECT 123.065 199.235 124.275 199.755 ;
        RECT 124.445 199.405 125.655 199.925 ;
        RECT 126.305 200.165 127.475 200.335 ;
        RECT 127.645 200.215 127.925 201.015 ;
        RECT 126.305 199.875 126.630 200.165 ;
        RECT 127.305 200.045 127.475 200.165 ;
        RECT 126.800 199.705 126.995 199.995 ;
        RECT 127.305 199.875 127.965 200.045 ;
        RECT 128.135 199.875 128.410 200.845 ;
        RECT 128.585 199.925 131.175 201.015 ;
        RECT 131.805 200.460 132.410 201.015 ;
        RECT 132.585 200.505 133.065 200.845 ;
        RECT 133.235 200.470 133.490 201.015 ;
        RECT 131.805 200.360 132.420 200.460 ;
        RECT 132.235 200.335 132.420 200.360 ;
        RECT 127.795 199.705 127.965 199.875 ;
        RECT 126.285 199.375 126.630 199.705 ;
        RECT 126.800 199.375 127.625 199.705 ;
        RECT 127.795 199.375 128.070 199.705 ;
        RECT 123.065 198.465 125.655 199.235 ;
        RECT 127.795 199.205 127.965 199.375 ;
        RECT 126.300 199.035 127.965 199.205 ;
        RECT 128.240 199.140 128.410 199.875 ;
        RECT 126.300 198.685 126.555 199.035 ;
        RECT 126.725 198.465 127.055 198.865 ;
        RECT 127.225 198.685 127.395 199.035 ;
        RECT 127.565 198.465 127.945 198.865 ;
        RECT 128.135 198.795 128.410 199.140 ;
        RECT 128.585 199.235 129.795 199.755 ;
        RECT 129.965 199.405 131.175 199.925 ;
        RECT 131.805 199.740 132.065 200.190 ;
        RECT 132.235 200.090 132.565 200.335 ;
        RECT 132.735 200.015 133.490 200.265 ;
        RECT 133.660 200.145 133.935 200.845 ;
        RECT 132.720 199.980 133.490 200.015 ;
        RECT 132.705 199.970 133.490 199.980 ;
        RECT 132.700 199.955 133.595 199.970 ;
        RECT 132.680 199.940 133.595 199.955 ;
        RECT 132.660 199.930 133.595 199.940 ;
        RECT 132.635 199.920 133.595 199.930 ;
        RECT 132.565 199.890 133.595 199.920 ;
        RECT 132.545 199.860 133.595 199.890 ;
        RECT 132.525 199.830 133.595 199.860 ;
        RECT 132.495 199.805 133.595 199.830 ;
        RECT 132.460 199.770 133.595 199.805 ;
        RECT 132.430 199.765 133.595 199.770 ;
        RECT 132.430 199.760 132.820 199.765 ;
        RECT 132.430 199.750 132.795 199.760 ;
        RECT 132.430 199.745 132.780 199.750 ;
        RECT 132.430 199.740 132.765 199.745 ;
        RECT 131.805 199.735 132.765 199.740 ;
        RECT 131.805 199.725 132.755 199.735 ;
        RECT 131.805 199.720 132.745 199.725 ;
        RECT 131.805 199.710 132.735 199.720 ;
        RECT 131.805 199.700 132.730 199.710 ;
        RECT 131.805 199.695 132.725 199.700 ;
        RECT 131.805 199.680 132.715 199.695 ;
        RECT 131.805 199.665 132.710 199.680 ;
        RECT 131.805 199.640 132.700 199.665 ;
        RECT 131.805 199.570 132.695 199.640 ;
        RECT 128.585 198.465 131.175 199.235 ;
        RECT 131.805 199.015 132.355 199.400 ;
        RECT 132.525 198.845 132.695 199.570 ;
        RECT 131.805 198.675 132.695 198.845 ;
        RECT 132.865 199.170 133.195 199.595 ;
        RECT 133.365 199.370 133.595 199.765 ;
        RECT 132.865 198.685 133.085 199.170 ;
        RECT 133.765 199.115 133.935 200.145 ;
        RECT 134.165 199.875 134.375 201.015 ;
        RECT 134.545 199.865 134.875 200.845 ;
        RECT 135.045 199.875 135.275 201.015 ;
        RECT 133.255 198.465 133.505 199.005 ;
        RECT 133.675 198.635 133.935 199.115 ;
        RECT 134.165 198.465 134.375 199.285 ;
        RECT 134.545 199.265 134.795 199.865 ;
        RECT 134.965 199.455 135.295 199.705 ;
        RECT 134.545 198.635 134.875 199.265 ;
        RECT 135.045 198.465 135.275 199.285 ;
        RECT 135.495 198.645 135.755 200.835 ;
        RECT 135.925 200.285 136.265 201.015 ;
        RECT 136.445 200.105 136.715 200.835 ;
        RECT 135.945 199.885 136.715 200.105 ;
        RECT 136.895 200.125 137.125 200.835 ;
        RECT 137.295 200.305 137.625 201.015 ;
        RECT 137.795 200.125 138.055 200.835 ;
        RECT 136.895 199.885 138.055 200.125 ;
        RECT 135.945 199.215 136.235 199.885 ;
        RECT 138.705 199.850 138.995 201.015 ;
        RECT 140.175 200.345 140.345 200.845 ;
        RECT 140.515 200.515 140.845 201.015 ;
        RECT 140.175 200.175 140.840 200.345 ;
        RECT 136.415 199.395 136.880 199.705 ;
        RECT 137.060 199.395 137.585 199.705 ;
        RECT 135.945 199.015 137.175 199.215 ;
        RECT 136.015 198.465 136.685 198.835 ;
        RECT 136.865 198.645 137.175 199.015 ;
        RECT 137.355 198.755 137.585 199.395 ;
        RECT 137.765 199.375 138.065 199.705 ;
        RECT 140.090 199.355 140.440 200.005 ;
        RECT 137.765 198.465 138.055 199.195 ;
        RECT 138.705 198.465 138.995 199.190 ;
        RECT 140.610 199.185 140.840 200.175 ;
        RECT 140.175 199.015 140.840 199.185 ;
        RECT 140.175 198.725 140.345 199.015 ;
        RECT 140.515 198.465 140.845 198.845 ;
        RECT 141.015 198.725 141.200 200.845 ;
        RECT 141.440 200.555 141.705 201.015 ;
        RECT 141.875 200.420 142.125 200.845 ;
        RECT 142.335 200.570 143.440 200.740 ;
        RECT 141.820 200.290 142.125 200.420 ;
        RECT 141.370 199.095 141.650 200.045 ;
        RECT 141.820 199.185 141.990 200.290 ;
        RECT 142.160 199.505 142.400 200.100 ;
        RECT 142.570 200.035 143.100 200.400 ;
        RECT 142.570 199.335 142.740 200.035 ;
        RECT 143.270 199.955 143.440 200.570 ;
        RECT 143.610 200.215 143.780 201.015 ;
        RECT 143.950 200.515 144.200 200.845 ;
        RECT 144.425 200.545 145.310 200.715 ;
        RECT 143.270 199.865 143.780 199.955 ;
        RECT 141.820 199.055 142.045 199.185 ;
        RECT 142.215 199.115 142.740 199.335 ;
        RECT 142.910 199.695 143.780 199.865 ;
        RECT 141.455 198.465 141.705 198.925 ;
        RECT 141.875 198.915 142.045 199.055 ;
        RECT 142.910 198.915 143.080 199.695 ;
        RECT 143.610 199.625 143.780 199.695 ;
        RECT 143.290 199.445 143.490 199.475 ;
        RECT 143.950 199.445 144.120 200.515 ;
        RECT 144.290 199.625 144.480 200.345 ;
        RECT 143.290 199.145 144.120 199.445 ;
        RECT 144.650 199.415 144.970 200.375 ;
        RECT 141.875 198.745 142.210 198.915 ;
        RECT 142.405 198.745 143.080 198.915 ;
        RECT 143.400 198.465 143.770 198.965 ;
        RECT 143.950 198.915 144.120 199.145 ;
        RECT 144.505 199.085 144.970 199.415 ;
        RECT 145.140 199.705 145.310 200.545 ;
        RECT 145.490 200.515 145.805 201.015 ;
        RECT 146.035 200.285 146.375 200.845 ;
        RECT 145.480 199.910 146.375 200.285 ;
        RECT 146.545 200.005 146.715 201.015 ;
        RECT 146.185 199.705 146.375 199.910 ;
        RECT 146.885 199.955 147.215 200.800 ;
        RECT 147.535 200.345 147.705 200.845 ;
        RECT 147.875 200.515 148.205 201.015 ;
        RECT 147.535 200.175 148.200 200.345 ;
        RECT 146.885 199.875 147.275 199.955 ;
        RECT 147.060 199.825 147.275 199.875 ;
        RECT 145.140 199.375 146.015 199.705 ;
        RECT 146.185 199.375 146.935 199.705 ;
        RECT 145.140 198.915 145.310 199.375 ;
        RECT 146.185 199.205 146.385 199.375 ;
        RECT 147.105 199.245 147.275 199.825 ;
        RECT 147.450 199.355 147.800 200.005 ;
        RECT 147.050 199.205 147.275 199.245 ;
        RECT 143.950 198.745 144.355 198.915 ;
        RECT 144.525 198.745 145.310 198.915 ;
        RECT 145.585 198.465 145.795 198.995 ;
        RECT 146.055 198.680 146.385 199.205 ;
        RECT 146.895 199.120 147.275 199.205 ;
        RECT 147.970 199.185 148.200 200.175 ;
        RECT 146.555 198.465 146.725 199.075 ;
        RECT 146.895 198.685 147.225 199.120 ;
        RECT 147.535 199.015 148.200 199.185 ;
        RECT 147.535 198.725 147.705 199.015 ;
        RECT 147.875 198.465 148.205 198.845 ;
        RECT 148.375 198.725 148.560 200.845 ;
        RECT 148.800 200.555 149.065 201.015 ;
        RECT 149.235 200.420 149.485 200.845 ;
        RECT 149.695 200.570 150.800 200.740 ;
        RECT 149.180 200.290 149.485 200.420 ;
        RECT 148.730 199.095 149.010 200.045 ;
        RECT 149.180 199.185 149.350 200.290 ;
        RECT 149.520 199.505 149.760 200.100 ;
        RECT 149.930 200.035 150.460 200.400 ;
        RECT 149.930 199.335 150.100 200.035 ;
        RECT 150.630 199.955 150.800 200.570 ;
        RECT 150.970 200.215 151.140 201.015 ;
        RECT 151.310 200.515 151.560 200.845 ;
        RECT 151.785 200.545 152.670 200.715 ;
        RECT 150.630 199.865 151.140 199.955 ;
        RECT 149.180 199.055 149.405 199.185 ;
        RECT 149.575 199.115 150.100 199.335 ;
        RECT 150.270 199.695 151.140 199.865 ;
        RECT 148.815 198.465 149.065 198.925 ;
        RECT 149.235 198.915 149.405 199.055 ;
        RECT 150.270 198.915 150.440 199.695 ;
        RECT 150.970 199.625 151.140 199.695 ;
        RECT 150.650 199.445 150.850 199.475 ;
        RECT 151.310 199.445 151.480 200.515 ;
        RECT 151.650 199.625 151.840 200.345 ;
        RECT 150.650 199.145 151.480 199.445 ;
        RECT 152.010 199.415 152.330 200.375 ;
        RECT 149.235 198.745 149.570 198.915 ;
        RECT 149.765 198.745 150.440 198.915 ;
        RECT 150.760 198.465 151.130 198.965 ;
        RECT 151.310 198.915 151.480 199.145 ;
        RECT 151.865 199.085 152.330 199.415 ;
        RECT 152.500 199.705 152.670 200.545 ;
        RECT 152.850 200.515 153.165 201.015 ;
        RECT 153.395 200.285 153.735 200.845 ;
        RECT 152.840 199.910 153.735 200.285 ;
        RECT 153.905 200.005 154.075 201.015 ;
        RECT 153.545 199.705 153.735 199.910 ;
        RECT 154.245 199.955 154.575 200.800 ;
        RECT 154.245 199.875 154.635 199.955 ;
        RECT 154.420 199.825 154.635 199.875 ;
        RECT 152.500 199.375 153.375 199.705 ;
        RECT 153.545 199.375 154.295 199.705 ;
        RECT 152.500 198.915 152.670 199.375 ;
        RECT 153.545 199.205 153.745 199.375 ;
        RECT 154.465 199.245 154.635 199.825 ;
        RECT 155.725 199.925 156.935 201.015 ;
        RECT 155.725 199.385 156.245 199.925 ;
        RECT 154.410 199.205 154.635 199.245 ;
        RECT 156.415 199.215 156.935 199.755 ;
        RECT 151.310 198.745 151.715 198.915 ;
        RECT 151.885 198.745 152.670 198.915 ;
        RECT 152.945 198.465 153.155 198.995 ;
        RECT 153.415 198.680 153.745 199.205 ;
        RECT 154.255 199.120 154.635 199.205 ;
        RECT 153.915 198.465 154.085 199.075 ;
        RECT 154.255 198.685 154.585 199.120 ;
        RECT 155.725 198.465 156.935 199.215 ;
        RECT 22.700 198.295 157.020 198.465 ;
        RECT 22.785 197.545 23.995 198.295 ;
        RECT 24.165 197.750 29.510 198.295 ;
        RECT 22.785 197.005 23.305 197.545 ;
        RECT 23.475 196.835 23.995 197.375 ;
        RECT 25.750 196.920 26.090 197.750 ;
        RECT 29.685 197.525 32.275 198.295 ;
        RECT 32.495 197.640 32.825 198.075 ;
        RECT 32.995 197.685 33.165 198.295 ;
        RECT 32.445 197.555 32.825 197.640 ;
        RECT 33.335 197.555 33.665 198.080 ;
        RECT 33.925 197.765 34.135 198.295 ;
        RECT 34.410 197.845 35.195 198.015 ;
        RECT 35.365 197.845 35.770 198.015 ;
        RECT 22.785 195.745 23.995 196.835 ;
        RECT 27.570 196.180 27.920 197.430 ;
        RECT 29.685 197.005 30.895 197.525 ;
        RECT 32.445 197.515 32.670 197.555 ;
        RECT 31.065 196.835 32.275 197.355 ;
        RECT 24.165 195.745 29.510 196.180 ;
        RECT 29.685 195.745 32.275 196.835 ;
        RECT 32.445 196.935 32.615 197.515 ;
        RECT 33.335 197.385 33.535 197.555 ;
        RECT 34.410 197.385 34.580 197.845 ;
        RECT 32.785 197.055 33.535 197.385 ;
        RECT 33.705 197.055 34.580 197.385 ;
        RECT 32.445 196.885 32.660 196.935 ;
        RECT 32.445 196.805 32.835 196.885 ;
        RECT 32.505 195.960 32.835 196.805 ;
        RECT 33.345 196.850 33.535 197.055 ;
        RECT 33.005 195.745 33.175 196.755 ;
        RECT 33.345 196.475 34.240 196.850 ;
        RECT 33.345 195.915 33.685 196.475 ;
        RECT 33.915 195.745 34.230 196.245 ;
        RECT 34.410 196.215 34.580 197.055 ;
        RECT 34.750 197.345 35.215 197.675 ;
        RECT 35.600 197.615 35.770 197.845 ;
        RECT 35.950 197.795 36.320 198.295 ;
        RECT 36.640 197.845 37.315 198.015 ;
        RECT 37.510 197.845 37.845 198.015 ;
        RECT 34.750 196.385 35.070 197.345 ;
        RECT 35.600 197.315 36.430 197.615 ;
        RECT 35.240 196.415 35.430 197.135 ;
        RECT 35.600 196.245 35.770 197.315 ;
        RECT 36.230 197.285 36.430 197.315 ;
        RECT 35.940 197.065 36.110 197.135 ;
        RECT 36.640 197.065 36.810 197.845 ;
        RECT 37.675 197.705 37.845 197.845 ;
        RECT 38.015 197.835 38.265 198.295 ;
        RECT 35.940 196.895 36.810 197.065 ;
        RECT 36.980 197.425 37.505 197.645 ;
        RECT 37.675 197.575 37.900 197.705 ;
        RECT 35.940 196.805 36.450 196.895 ;
        RECT 34.410 196.045 35.295 196.215 ;
        RECT 35.520 195.915 35.770 196.245 ;
        RECT 35.940 195.745 36.110 196.545 ;
        RECT 36.280 196.190 36.450 196.805 ;
        RECT 36.980 196.725 37.150 197.425 ;
        RECT 36.620 196.360 37.150 196.725 ;
        RECT 37.320 196.660 37.560 197.255 ;
        RECT 37.730 196.470 37.900 197.575 ;
        RECT 38.070 196.715 38.350 197.665 ;
        RECT 37.595 196.340 37.900 196.470 ;
        RECT 36.280 196.020 37.385 196.190 ;
        RECT 37.595 195.915 37.845 196.340 ;
        RECT 38.015 195.745 38.280 196.205 ;
        RECT 38.520 195.915 38.705 198.035 ;
        RECT 38.875 197.915 39.205 198.295 ;
        RECT 39.375 197.745 39.545 198.035 ;
        RECT 38.880 197.575 39.545 197.745 ;
        RECT 38.880 196.585 39.110 197.575 ;
        RECT 39.805 197.525 41.475 198.295 ;
        RECT 42.105 197.645 42.365 198.125 ;
        RECT 42.535 197.755 42.785 198.295 ;
        RECT 39.280 196.755 39.630 197.405 ;
        RECT 39.805 197.005 40.555 197.525 ;
        RECT 40.725 196.835 41.475 197.355 ;
        RECT 38.880 196.415 39.545 196.585 ;
        RECT 38.875 195.745 39.205 196.245 ;
        RECT 39.375 195.915 39.545 196.415 ;
        RECT 39.805 195.745 41.475 196.835 ;
        RECT 42.105 196.615 42.275 197.645 ;
        RECT 42.955 197.590 43.175 198.075 ;
        RECT 42.445 196.995 42.675 197.390 ;
        RECT 42.845 197.165 43.175 197.590 ;
        RECT 43.345 197.915 44.235 198.085 ;
        RECT 43.345 197.190 43.515 197.915 ;
        RECT 43.685 197.360 44.235 197.745 ;
        RECT 44.405 197.525 47.915 198.295 ;
        RECT 48.545 197.570 48.835 198.295 ;
        RECT 49.005 197.555 49.325 198.035 ;
        RECT 49.495 197.725 49.725 198.125 ;
        RECT 49.895 197.905 50.245 198.295 ;
        RECT 49.495 197.645 50.005 197.725 ;
        RECT 50.415 197.645 50.745 198.125 ;
        RECT 49.495 197.555 50.745 197.645 ;
        RECT 43.345 197.120 44.235 197.190 ;
        RECT 43.340 197.095 44.235 197.120 ;
        RECT 43.330 197.080 44.235 197.095 ;
        RECT 43.325 197.065 44.235 197.080 ;
        RECT 43.315 197.060 44.235 197.065 ;
        RECT 43.310 197.050 44.235 197.060 ;
        RECT 43.305 197.040 44.235 197.050 ;
        RECT 43.295 197.035 44.235 197.040 ;
        RECT 43.285 197.025 44.235 197.035 ;
        RECT 43.275 197.020 44.235 197.025 ;
        RECT 43.275 197.015 43.610 197.020 ;
        RECT 43.260 197.010 43.610 197.015 ;
        RECT 43.245 197.000 43.610 197.010 ;
        RECT 43.220 196.995 43.610 197.000 ;
        RECT 42.445 196.990 43.610 196.995 ;
        RECT 42.445 196.955 43.580 196.990 ;
        RECT 42.445 196.930 43.545 196.955 ;
        RECT 42.445 196.900 43.515 196.930 ;
        RECT 42.445 196.870 43.495 196.900 ;
        RECT 42.445 196.840 43.475 196.870 ;
        RECT 42.445 196.830 43.405 196.840 ;
        RECT 42.445 196.820 43.380 196.830 ;
        RECT 42.445 196.805 43.360 196.820 ;
        RECT 42.445 196.790 43.340 196.805 ;
        RECT 42.550 196.780 43.335 196.790 ;
        RECT 42.550 196.745 43.320 196.780 ;
        RECT 42.105 195.915 42.380 196.615 ;
        RECT 42.550 196.495 43.305 196.745 ;
        RECT 43.475 196.425 43.805 196.670 ;
        RECT 43.975 196.570 44.235 197.020 ;
        RECT 44.405 197.005 46.055 197.525 ;
        RECT 46.225 196.835 47.915 197.355 ;
        RECT 43.620 196.400 43.805 196.425 ;
        RECT 43.620 196.300 44.235 196.400 ;
        RECT 42.550 195.745 42.805 196.290 ;
        RECT 42.975 195.915 43.455 196.255 ;
        RECT 43.630 195.745 44.235 196.300 ;
        RECT 44.405 195.745 47.915 196.835 ;
        RECT 48.545 195.745 48.835 196.910 ;
        RECT 49.005 196.625 49.175 197.555 ;
        RECT 49.835 197.475 50.745 197.555 ;
        RECT 50.915 197.475 51.085 198.295 ;
        RECT 51.590 197.555 52.055 198.100 ;
        RECT 52.315 197.745 52.485 198.035 ;
        RECT 52.655 197.915 52.985 198.295 ;
        RECT 52.315 197.575 52.980 197.745 ;
        RECT 49.345 196.965 49.515 197.385 ;
        RECT 49.745 197.135 50.345 197.305 ;
        RECT 49.345 196.795 50.005 196.965 ;
        RECT 49.005 196.425 49.665 196.625 ;
        RECT 49.835 196.595 50.005 196.795 ;
        RECT 50.175 196.935 50.345 197.135 ;
        RECT 50.515 197.105 51.210 197.305 ;
        RECT 51.470 196.935 51.715 197.385 ;
        RECT 50.175 196.765 51.715 196.935 ;
        RECT 51.885 196.595 52.055 197.555 ;
        RECT 52.230 196.755 52.580 197.405 ;
        RECT 49.835 196.425 52.055 196.595 ;
        RECT 52.750 196.585 52.980 197.575 ;
        RECT 49.495 196.255 49.665 196.425 ;
        RECT 49.025 195.745 49.325 196.255 ;
        RECT 49.495 196.085 49.875 196.255 ;
        RECT 50.455 195.745 51.085 196.255 ;
        RECT 51.255 195.915 51.585 196.425 ;
        RECT 52.315 196.415 52.980 196.585 ;
        RECT 51.755 195.745 52.055 196.255 ;
        RECT 52.315 195.915 52.485 196.415 ;
        RECT 52.655 195.745 52.985 196.245 ;
        RECT 53.155 195.915 53.340 198.035 ;
        RECT 53.595 197.835 53.845 198.295 ;
        RECT 54.015 197.845 54.350 198.015 ;
        RECT 54.545 197.845 55.220 198.015 ;
        RECT 54.015 197.705 54.185 197.845 ;
        RECT 53.510 196.715 53.790 197.665 ;
        RECT 53.960 197.575 54.185 197.705 ;
        RECT 53.960 196.470 54.130 197.575 ;
        RECT 54.355 197.425 54.880 197.645 ;
        RECT 54.300 196.660 54.540 197.255 ;
        RECT 54.710 196.725 54.880 197.425 ;
        RECT 55.050 197.065 55.220 197.845 ;
        RECT 55.540 197.795 55.910 198.295 ;
        RECT 56.090 197.845 56.495 198.015 ;
        RECT 56.665 197.845 57.450 198.015 ;
        RECT 56.090 197.615 56.260 197.845 ;
        RECT 55.430 197.315 56.260 197.615 ;
        RECT 56.645 197.345 57.110 197.675 ;
        RECT 55.430 197.285 55.630 197.315 ;
        RECT 55.750 197.065 55.920 197.135 ;
        RECT 55.050 196.895 55.920 197.065 ;
        RECT 55.410 196.805 55.920 196.895 ;
        RECT 53.960 196.340 54.265 196.470 ;
        RECT 54.710 196.360 55.240 196.725 ;
        RECT 53.580 195.745 53.845 196.205 ;
        RECT 54.015 195.915 54.265 196.340 ;
        RECT 55.410 196.190 55.580 196.805 ;
        RECT 54.475 196.020 55.580 196.190 ;
        RECT 55.750 195.745 55.920 196.545 ;
        RECT 56.090 196.245 56.260 197.315 ;
        RECT 56.430 196.415 56.620 197.135 ;
        RECT 56.790 196.385 57.110 197.345 ;
        RECT 57.280 197.385 57.450 197.845 ;
        RECT 57.725 197.765 57.935 198.295 ;
        RECT 58.195 197.555 58.525 198.080 ;
        RECT 58.695 197.685 58.865 198.295 ;
        RECT 59.035 197.640 59.365 198.075 ;
        RECT 59.585 197.645 59.845 198.125 ;
        RECT 60.015 197.755 60.265 198.295 ;
        RECT 59.035 197.555 59.415 197.640 ;
        RECT 58.325 197.385 58.525 197.555 ;
        RECT 59.190 197.515 59.415 197.555 ;
        RECT 57.280 197.055 58.155 197.385 ;
        RECT 58.325 197.055 59.075 197.385 ;
        RECT 56.090 195.915 56.340 196.245 ;
        RECT 57.280 196.215 57.450 197.055 ;
        RECT 58.325 196.850 58.515 197.055 ;
        RECT 59.245 196.935 59.415 197.515 ;
        RECT 59.200 196.885 59.415 196.935 ;
        RECT 57.620 196.475 58.515 196.850 ;
        RECT 59.025 196.805 59.415 196.885 ;
        RECT 56.565 196.045 57.450 196.215 ;
        RECT 57.630 195.745 57.945 196.245 ;
        RECT 58.175 195.915 58.515 196.475 ;
        RECT 58.685 195.745 58.855 196.755 ;
        RECT 59.025 195.960 59.355 196.805 ;
        RECT 59.585 196.615 59.755 197.645 ;
        RECT 60.435 197.590 60.655 198.075 ;
        RECT 59.925 196.995 60.155 197.390 ;
        RECT 60.325 197.165 60.655 197.590 ;
        RECT 60.825 197.915 61.715 198.085 ;
        RECT 60.825 197.190 60.995 197.915 ;
        RECT 61.895 197.785 63.125 198.125 ;
        RECT 63.295 197.805 63.550 198.295 ;
        RECT 61.165 197.360 61.715 197.745 ;
        RECT 61.895 197.555 62.225 197.785 ;
        RECT 60.825 197.120 61.715 197.190 ;
        RECT 60.820 197.095 61.715 197.120 ;
        RECT 60.810 197.080 61.715 197.095 ;
        RECT 60.805 197.065 61.715 197.080 ;
        RECT 60.795 197.060 61.715 197.065 ;
        RECT 60.790 197.050 61.715 197.060 ;
        RECT 61.885 197.055 62.195 197.385 ;
        RECT 62.400 197.055 62.775 197.615 ;
        RECT 60.785 197.040 61.715 197.050 ;
        RECT 60.775 197.035 61.715 197.040 ;
        RECT 60.765 197.025 61.715 197.035 ;
        RECT 60.755 197.020 61.715 197.025 ;
        RECT 60.755 197.015 61.090 197.020 ;
        RECT 60.740 197.010 61.090 197.015 ;
        RECT 60.725 197.000 61.090 197.010 ;
        RECT 60.700 196.995 61.090 197.000 ;
        RECT 59.925 196.990 61.090 196.995 ;
        RECT 59.925 196.955 61.060 196.990 ;
        RECT 59.925 196.930 61.025 196.955 ;
        RECT 59.925 196.900 60.995 196.930 ;
        RECT 59.925 196.870 60.975 196.900 ;
        RECT 59.925 196.840 60.955 196.870 ;
        RECT 59.925 196.830 60.885 196.840 ;
        RECT 59.925 196.820 60.860 196.830 ;
        RECT 59.925 196.805 60.840 196.820 ;
        RECT 59.925 196.790 60.820 196.805 ;
        RECT 60.030 196.780 60.815 196.790 ;
        RECT 60.030 196.745 60.800 196.780 ;
        RECT 59.585 195.915 59.860 196.615 ;
        RECT 60.030 196.495 60.785 196.745 ;
        RECT 60.955 196.425 61.285 196.670 ;
        RECT 61.455 196.570 61.715 197.020 ;
        RECT 62.945 196.885 63.125 197.785 ;
        RECT 64.735 197.745 64.905 198.035 ;
        RECT 65.075 197.915 65.405 198.295 ;
        RECT 63.310 197.055 63.530 197.635 ;
        RECT 64.735 197.575 65.400 197.745 ;
        RECT 61.895 196.715 63.125 196.885 ;
        RECT 61.100 196.400 61.285 196.425 ;
        RECT 61.100 196.300 61.715 196.400 ;
        RECT 60.030 195.745 60.285 196.290 ;
        RECT 60.455 195.915 60.935 196.255 ;
        RECT 61.110 195.745 61.715 196.300 ;
        RECT 61.895 195.915 62.225 196.715 ;
        RECT 62.395 195.745 62.625 196.545 ;
        RECT 62.795 195.915 63.125 196.715 ;
        RECT 63.295 195.745 63.550 196.885 ;
        RECT 64.650 196.755 65.000 197.405 ;
        RECT 65.170 196.585 65.400 197.575 ;
        RECT 64.735 196.415 65.400 196.585 ;
        RECT 64.735 195.915 64.905 196.415 ;
        RECT 65.075 195.745 65.405 196.245 ;
        RECT 65.575 195.915 65.760 198.035 ;
        RECT 66.015 197.835 66.265 198.295 ;
        RECT 66.435 197.845 66.770 198.015 ;
        RECT 66.965 197.845 67.640 198.015 ;
        RECT 66.435 197.705 66.605 197.845 ;
        RECT 65.930 196.715 66.210 197.665 ;
        RECT 66.380 197.575 66.605 197.705 ;
        RECT 66.380 196.470 66.550 197.575 ;
        RECT 66.775 197.425 67.300 197.645 ;
        RECT 66.720 196.660 66.960 197.255 ;
        RECT 67.130 196.725 67.300 197.425 ;
        RECT 67.470 197.065 67.640 197.845 ;
        RECT 67.960 197.795 68.330 198.295 ;
        RECT 68.510 197.845 68.915 198.015 ;
        RECT 69.085 197.845 69.870 198.015 ;
        RECT 68.510 197.615 68.680 197.845 ;
        RECT 67.850 197.315 68.680 197.615 ;
        RECT 69.065 197.345 69.530 197.675 ;
        RECT 67.850 197.285 68.050 197.315 ;
        RECT 68.170 197.065 68.340 197.135 ;
        RECT 67.470 196.895 68.340 197.065 ;
        RECT 67.830 196.805 68.340 196.895 ;
        RECT 66.380 196.340 66.685 196.470 ;
        RECT 67.130 196.360 67.660 196.725 ;
        RECT 66.000 195.745 66.265 196.205 ;
        RECT 66.435 195.915 66.685 196.340 ;
        RECT 67.830 196.190 68.000 196.805 ;
        RECT 66.895 196.020 68.000 196.190 ;
        RECT 68.170 195.745 68.340 196.545 ;
        RECT 68.510 196.245 68.680 197.315 ;
        RECT 68.850 196.415 69.040 197.135 ;
        RECT 69.210 196.385 69.530 197.345 ;
        RECT 69.700 197.385 69.870 197.845 ;
        RECT 70.145 197.765 70.355 198.295 ;
        RECT 70.615 197.555 70.945 198.080 ;
        RECT 71.115 197.685 71.285 198.295 ;
        RECT 71.455 197.640 71.785 198.075 ;
        RECT 71.455 197.555 71.835 197.640 ;
        RECT 70.745 197.385 70.945 197.555 ;
        RECT 71.610 197.515 71.835 197.555 ;
        RECT 69.700 197.055 70.575 197.385 ;
        RECT 70.745 197.055 71.495 197.385 ;
        RECT 68.510 195.915 68.760 196.245 ;
        RECT 69.700 196.215 69.870 197.055 ;
        RECT 70.745 196.850 70.935 197.055 ;
        RECT 71.665 196.935 71.835 197.515 ;
        RECT 72.015 197.485 72.285 198.295 ;
        RECT 72.455 197.485 72.785 198.125 ;
        RECT 72.955 197.485 73.195 198.295 ;
        RECT 74.305 197.570 74.595 198.295 ;
        RECT 72.005 197.055 72.355 197.305 ;
        RECT 71.620 196.885 71.835 196.935 ;
        RECT 72.525 196.885 72.695 197.485 ;
        RECT 74.805 197.475 75.035 198.295 ;
        RECT 75.205 197.495 75.535 198.125 ;
        RECT 72.865 197.055 73.215 197.305 ;
        RECT 74.785 197.055 75.115 197.305 ;
        RECT 70.040 196.475 70.935 196.850 ;
        RECT 71.445 196.805 71.835 196.885 ;
        RECT 68.985 196.045 69.870 196.215 ;
        RECT 70.050 195.745 70.365 196.245 ;
        RECT 70.595 195.915 70.935 196.475 ;
        RECT 71.105 195.745 71.275 196.755 ;
        RECT 71.445 195.960 71.775 196.805 ;
        RECT 72.015 195.745 72.345 196.885 ;
        RECT 72.525 196.715 73.205 196.885 ;
        RECT 72.875 195.930 73.205 196.715 ;
        RECT 74.305 195.745 74.595 196.910 ;
        RECT 75.285 196.895 75.535 197.495 ;
        RECT 75.705 197.475 75.915 198.295 ;
        RECT 76.145 197.475 76.405 198.295 ;
        RECT 76.575 197.475 76.905 197.895 ;
        RECT 77.085 197.810 77.875 198.075 ;
        RECT 76.655 197.385 76.905 197.475 ;
        RECT 74.805 195.745 75.035 196.885 ;
        RECT 75.205 195.915 75.535 196.895 ;
        RECT 75.705 195.745 75.915 196.885 ;
        RECT 76.145 196.425 76.485 197.305 ;
        RECT 76.655 197.135 77.450 197.385 ;
        RECT 76.145 195.745 76.405 196.255 ;
        RECT 76.655 195.915 76.825 197.135 ;
        RECT 77.620 196.955 77.875 197.810 ;
        RECT 78.045 197.655 78.245 198.075 ;
        RECT 78.435 197.835 78.765 198.295 ;
        RECT 78.045 197.135 78.455 197.655 ;
        RECT 78.935 197.645 79.195 198.125 ;
        RECT 78.625 196.955 78.855 197.385 ;
        RECT 77.065 196.785 78.855 196.955 ;
        RECT 77.065 196.420 77.315 196.785 ;
        RECT 77.485 196.425 77.815 196.615 ;
        RECT 78.035 196.490 78.750 196.785 ;
        RECT 79.025 196.615 79.195 197.645 ;
        RECT 79.365 197.525 82.875 198.295 ;
        RECT 83.045 197.545 84.255 198.295 ;
        RECT 79.365 197.005 81.015 197.525 ;
        RECT 81.185 196.835 82.875 197.355 ;
        RECT 83.045 197.005 83.565 197.545 ;
        RECT 84.425 197.475 84.685 198.295 ;
        RECT 84.855 197.475 85.185 197.895 ;
        RECT 85.365 197.810 86.155 198.075 ;
        RECT 84.935 197.385 85.185 197.475 ;
        RECT 83.735 196.835 84.255 197.375 ;
        RECT 77.485 196.250 77.680 196.425 ;
        RECT 77.065 195.745 77.680 196.250 ;
        RECT 77.850 195.915 78.325 196.255 ;
        RECT 78.495 195.745 78.710 196.290 ;
        RECT 78.920 195.915 79.195 196.615 ;
        RECT 79.365 195.745 82.875 196.835 ;
        RECT 83.045 195.745 84.255 196.835 ;
        RECT 84.425 196.425 84.765 197.305 ;
        RECT 84.935 197.135 85.730 197.385 ;
        RECT 84.425 195.745 84.685 196.255 ;
        RECT 84.935 195.915 85.105 197.135 ;
        RECT 85.900 196.955 86.155 197.810 ;
        RECT 86.325 197.655 86.525 198.075 ;
        RECT 86.715 197.835 87.045 198.295 ;
        RECT 86.325 197.135 86.735 197.655 ;
        RECT 87.215 197.645 87.475 198.125 ;
        RECT 86.905 196.955 87.135 197.385 ;
        RECT 85.345 196.785 87.135 196.955 ;
        RECT 85.345 196.420 85.595 196.785 ;
        RECT 85.765 196.425 86.095 196.615 ;
        RECT 86.315 196.490 87.030 196.785 ;
        RECT 87.305 196.615 87.475 197.645 ;
        RECT 87.645 197.545 88.855 198.295 ;
        RECT 87.645 197.005 88.165 197.545 ;
        RECT 89.025 197.475 89.285 198.295 ;
        RECT 89.455 197.475 89.785 197.895 ;
        RECT 89.965 197.810 90.755 198.075 ;
        RECT 89.535 197.385 89.785 197.475 ;
        RECT 88.335 196.835 88.855 197.375 ;
        RECT 85.765 196.250 85.960 196.425 ;
        RECT 85.345 195.745 85.960 196.250 ;
        RECT 86.130 195.915 86.605 196.255 ;
        RECT 86.775 195.745 86.990 196.290 ;
        RECT 87.200 195.915 87.475 196.615 ;
        RECT 87.645 195.745 88.855 196.835 ;
        RECT 89.025 196.425 89.365 197.305 ;
        RECT 89.535 197.135 90.330 197.385 ;
        RECT 89.025 195.745 89.285 196.255 ;
        RECT 89.535 195.915 89.705 197.135 ;
        RECT 90.500 196.955 90.755 197.810 ;
        RECT 90.925 197.655 91.125 198.075 ;
        RECT 91.315 197.835 91.645 198.295 ;
        RECT 90.925 197.135 91.335 197.655 ;
        RECT 91.815 197.645 92.075 198.125 ;
        RECT 92.410 197.785 92.650 198.295 ;
        RECT 92.830 197.785 93.110 198.115 ;
        RECT 93.340 197.785 93.555 198.295 ;
        RECT 91.505 196.955 91.735 197.385 ;
        RECT 89.945 196.785 91.735 196.955 ;
        RECT 89.945 196.420 90.195 196.785 ;
        RECT 90.365 196.425 90.695 196.615 ;
        RECT 90.915 196.490 91.630 196.785 ;
        RECT 91.905 196.615 92.075 197.645 ;
        RECT 92.305 197.055 92.660 197.615 ;
        RECT 92.830 196.885 93.000 197.785 ;
        RECT 93.170 197.055 93.435 197.615 ;
        RECT 93.725 197.555 94.340 198.125 ;
        RECT 95.005 197.915 95.895 198.085 ;
        RECT 93.685 196.885 93.855 197.385 ;
        RECT 90.365 196.250 90.560 196.425 ;
        RECT 89.945 195.745 90.560 196.250 ;
        RECT 90.730 195.915 91.205 196.255 ;
        RECT 91.375 195.745 91.590 196.290 ;
        RECT 91.800 195.915 92.075 196.615 ;
        RECT 92.430 196.715 93.855 196.885 ;
        RECT 92.430 196.540 92.820 196.715 ;
        RECT 93.305 195.745 93.635 196.545 ;
        RECT 94.025 196.535 94.340 197.555 ;
        RECT 95.005 197.360 95.555 197.745 ;
        RECT 95.725 197.190 95.895 197.915 ;
        RECT 95.005 197.120 95.895 197.190 ;
        RECT 96.065 197.590 96.285 198.075 ;
        RECT 96.455 197.755 96.705 198.295 ;
        RECT 96.875 197.645 97.135 198.125 ;
        RECT 96.065 197.165 96.395 197.590 ;
        RECT 95.005 197.095 95.900 197.120 ;
        RECT 95.005 197.080 95.910 197.095 ;
        RECT 95.005 197.065 95.915 197.080 ;
        RECT 95.005 197.060 95.925 197.065 ;
        RECT 95.005 197.050 95.930 197.060 ;
        RECT 95.005 197.040 95.935 197.050 ;
        RECT 95.005 197.035 95.945 197.040 ;
        RECT 95.005 197.025 95.955 197.035 ;
        RECT 95.005 197.020 95.965 197.025 ;
        RECT 95.005 196.570 95.265 197.020 ;
        RECT 95.630 197.015 95.965 197.020 ;
        RECT 95.630 197.010 95.980 197.015 ;
        RECT 95.630 197.000 95.995 197.010 ;
        RECT 95.630 196.995 96.020 197.000 ;
        RECT 96.565 196.995 96.795 197.390 ;
        RECT 95.630 196.990 96.795 196.995 ;
        RECT 95.660 196.955 96.795 196.990 ;
        RECT 95.695 196.930 96.795 196.955 ;
        RECT 95.725 196.900 96.795 196.930 ;
        RECT 95.745 196.870 96.795 196.900 ;
        RECT 95.765 196.840 96.795 196.870 ;
        RECT 95.835 196.830 96.795 196.840 ;
        RECT 95.860 196.820 96.795 196.830 ;
        RECT 95.880 196.805 96.795 196.820 ;
        RECT 95.900 196.790 96.795 196.805 ;
        RECT 95.905 196.780 96.690 196.790 ;
        RECT 95.920 196.745 96.690 196.780 ;
        RECT 93.805 195.915 94.340 196.535 ;
        RECT 95.435 196.425 95.765 196.670 ;
        RECT 95.935 196.495 96.690 196.745 ;
        RECT 96.965 196.615 97.135 197.645 ;
        RECT 95.435 196.400 95.620 196.425 ;
        RECT 95.005 196.300 95.620 196.400 ;
        RECT 95.005 195.745 95.610 196.300 ;
        RECT 95.785 195.915 96.265 196.255 ;
        RECT 96.435 195.745 96.690 196.290 ;
        RECT 96.860 195.915 97.135 196.615 ;
        RECT 97.305 197.795 97.565 198.125 ;
        RECT 97.775 197.815 98.050 198.295 ;
        RECT 97.305 196.885 97.475 197.795 ;
        RECT 98.260 197.725 98.465 198.125 ;
        RECT 98.635 197.895 98.970 198.295 ;
        RECT 97.645 197.055 98.005 197.635 ;
        RECT 98.260 197.555 98.945 197.725 ;
        RECT 100.065 197.570 100.355 198.295 ;
        RECT 100.690 197.785 100.930 198.295 ;
        RECT 101.110 197.785 101.390 198.115 ;
        RECT 101.620 197.785 101.835 198.295 ;
        RECT 98.185 196.885 98.435 197.385 ;
        RECT 97.305 196.715 98.435 196.885 ;
        RECT 97.305 195.945 97.575 196.715 ;
        RECT 98.605 196.525 98.945 197.555 ;
        RECT 100.585 197.055 100.940 197.615 ;
        RECT 97.745 195.745 98.075 196.525 ;
        RECT 98.280 196.350 98.945 196.525 ;
        RECT 98.280 195.945 98.465 196.350 ;
        RECT 98.635 195.745 98.970 196.170 ;
        RECT 100.065 195.745 100.355 196.910 ;
        RECT 101.110 196.885 101.280 197.785 ;
        RECT 101.450 197.055 101.715 197.615 ;
        RECT 102.005 197.555 102.620 198.125 ;
        RECT 103.835 197.745 104.005 198.035 ;
        RECT 104.175 197.915 104.505 198.295 ;
        RECT 103.835 197.575 104.500 197.745 ;
        RECT 101.965 196.885 102.135 197.385 ;
        RECT 100.710 196.715 102.135 196.885 ;
        RECT 100.710 196.540 101.100 196.715 ;
        RECT 101.585 195.745 101.915 196.545 ;
        RECT 102.305 196.535 102.620 197.555 ;
        RECT 103.750 196.755 104.100 197.405 ;
        RECT 104.270 196.585 104.500 197.575 ;
        RECT 102.085 195.915 102.620 196.535 ;
        RECT 103.835 196.415 104.500 196.585 ;
        RECT 103.835 195.915 104.005 196.415 ;
        RECT 104.175 195.745 104.505 196.245 ;
        RECT 104.675 195.915 104.860 198.035 ;
        RECT 105.115 197.835 105.365 198.295 ;
        RECT 105.535 197.845 105.870 198.015 ;
        RECT 106.065 197.845 106.740 198.015 ;
        RECT 105.535 197.705 105.705 197.845 ;
        RECT 105.030 196.715 105.310 197.665 ;
        RECT 105.480 197.575 105.705 197.705 ;
        RECT 105.480 196.470 105.650 197.575 ;
        RECT 105.875 197.425 106.400 197.645 ;
        RECT 105.820 196.660 106.060 197.255 ;
        RECT 106.230 196.725 106.400 197.425 ;
        RECT 106.570 197.065 106.740 197.845 ;
        RECT 107.060 197.795 107.430 198.295 ;
        RECT 107.610 197.845 108.015 198.015 ;
        RECT 108.185 197.845 108.970 198.015 ;
        RECT 107.610 197.615 107.780 197.845 ;
        RECT 106.950 197.315 107.780 197.615 ;
        RECT 108.165 197.345 108.630 197.675 ;
        RECT 106.950 197.285 107.150 197.315 ;
        RECT 107.270 197.065 107.440 197.135 ;
        RECT 106.570 196.895 107.440 197.065 ;
        RECT 106.930 196.805 107.440 196.895 ;
        RECT 105.480 196.340 105.785 196.470 ;
        RECT 106.230 196.360 106.760 196.725 ;
        RECT 105.100 195.745 105.365 196.205 ;
        RECT 105.535 195.915 105.785 196.340 ;
        RECT 106.930 196.190 107.100 196.805 ;
        RECT 105.995 196.020 107.100 196.190 ;
        RECT 107.270 195.745 107.440 196.545 ;
        RECT 107.610 196.245 107.780 197.315 ;
        RECT 107.950 196.415 108.140 197.135 ;
        RECT 108.310 196.385 108.630 197.345 ;
        RECT 108.800 197.385 108.970 197.845 ;
        RECT 109.245 197.765 109.455 198.295 ;
        RECT 109.715 197.555 110.045 198.080 ;
        RECT 110.215 197.685 110.385 198.295 ;
        RECT 110.555 197.640 110.885 198.075 ;
        RECT 110.555 197.555 110.935 197.640 ;
        RECT 109.845 197.385 110.045 197.555 ;
        RECT 110.710 197.515 110.935 197.555 ;
        RECT 108.800 197.055 109.675 197.385 ;
        RECT 109.845 197.055 110.595 197.385 ;
        RECT 107.610 195.915 107.860 196.245 ;
        RECT 108.800 196.215 108.970 197.055 ;
        RECT 109.845 196.850 110.035 197.055 ;
        RECT 110.765 196.935 110.935 197.515 ;
        RECT 111.165 197.475 111.375 198.295 ;
        RECT 111.545 197.495 111.875 198.125 ;
        RECT 110.720 196.885 110.935 196.935 ;
        RECT 111.545 196.895 111.795 197.495 ;
        RECT 112.045 197.475 112.275 198.295 ;
        RECT 113.495 197.745 113.665 198.035 ;
        RECT 113.835 197.915 114.165 198.295 ;
        RECT 113.495 197.575 114.160 197.745 ;
        RECT 111.965 197.055 112.295 197.305 ;
        RECT 109.140 196.475 110.035 196.850 ;
        RECT 110.545 196.805 110.935 196.885 ;
        RECT 108.085 196.045 108.970 196.215 ;
        RECT 109.150 195.745 109.465 196.245 ;
        RECT 109.695 195.915 110.035 196.475 ;
        RECT 110.205 195.745 110.375 196.755 ;
        RECT 110.545 195.960 110.875 196.805 ;
        RECT 111.165 195.745 111.375 196.885 ;
        RECT 111.545 195.915 111.875 196.895 ;
        RECT 112.045 195.745 112.275 196.885 ;
        RECT 113.410 196.755 113.760 197.405 ;
        RECT 113.930 196.585 114.160 197.575 ;
        RECT 113.495 196.415 114.160 196.585 ;
        RECT 113.495 195.915 113.665 196.415 ;
        RECT 113.835 195.745 114.165 196.245 ;
        RECT 114.335 195.915 114.520 198.035 ;
        RECT 114.775 197.835 115.025 198.295 ;
        RECT 115.195 197.845 115.530 198.015 ;
        RECT 115.725 197.845 116.400 198.015 ;
        RECT 115.195 197.705 115.365 197.845 ;
        RECT 114.690 196.715 114.970 197.665 ;
        RECT 115.140 197.575 115.365 197.705 ;
        RECT 115.140 196.470 115.310 197.575 ;
        RECT 115.535 197.425 116.060 197.645 ;
        RECT 115.480 196.660 115.720 197.255 ;
        RECT 115.890 196.725 116.060 197.425 ;
        RECT 116.230 197.065 116.400 197.845 ;
        RECT 116.720 197.795 117.090 198.295 ;
        RECT 117.270 197.845 117.675 198.015 ;
        RECT 117.845 197.845 118.630 198.015 ;
        RECT 117.270 197.615 117.440 197.845 ;
        RECT 116.610 197.315 117.440 197.615 ;
        RECT 117.825 197.345 118.290 197.675 ;
        RECT 116.610 197.285 116.810 197.315 ;
        RECT 116.930 197.065 117.100 197.135 ;
        RECT 116.230 196.895 117.100 197.065 ;
        RECT 116.590 196.805 117.100 196.895 ;
        RECT 115.140 196.340 115.445 196.470 ;
        RECT 115.890 196.360 116.420 196.725 ;
        RECT 114.760 195.745 115.025 196.205 ;
        RECT 115.195 195.915 115.445 196.340 ;
        RECT 116.590 196.190 116.760 196.805 ;
        RECT 115.655 196.020 116.760 196.190 ;
        RECT 116.930 195.745 117.100 196.545 ;
        RECT 117.270 196.245 117.440 197.315 ;
        RECT 117.610 196.415 117.800 197.135 ;
        RECT 117.970 196.385 118.290 197.345 ;
        RECT 118.460 197.385 118.630 197.845 ;
        RECT 118.905 197.765 119.115 198.295 ;
        RECT 119.375 197.555 119.705 198.080 ;
        RECT 119.875 197.685 120.045 198.295 ;
        RECT 120.215 197.640 120.545 198.075 ;
        RECT 120.215 197.555 120.595 197.640 ;
        RECT 119.505 197.385 119.705 197.555 ;
        RECT 120.370 197.515 120.595 197.555 ;
        RECT 118.460 197.055 119.335 197.385 ;
        RECT 119.505 197.055 120.255 197.385 ;
        RECT 117.270 195.915 117.520 196.245 ;
        RECT 118.460 196.215 118.630 197.055 ;
        RECT 119.505 196.850 119.695 197.055 ;
        RECT 120.425 196.935 120.595 197.515 ;
        RECT 120.380 196.885 120.595 196.935 ;
        RECT 118.800 196.475 119.695 196.850 ;
        RECT 120.205 196.805 120.595 196.885 ;
        RECT 120.765 197.555 121.150 198.125 ;
        RECT 121.320 197.835 121.645 198.295 ;
        RECT 122.165 197.665 122.445 198.125 ;
        RECT 120.765 196.885 121.045 197.555 ;
        RECT 121.320 197.495 122.445 197.665 ;
        RECT 121.320 197.385 121.770 197.495 ;
        RECT 121.215 197.055 121.770 197.385 ;
        RECT 122.635 197.325 123.035 198.125 ;
        RECT 123.435 197.835 123.705 198.295 ;
        RECT 123.875 197.665 124.160 198.125 ;
        RECT 117.745 196.045 118.630 196.215 ;
        RECT 118.810 195.745 119.125 196.245 ;
        RECT 119.355 195.915 119.695 196.475 ;
        RECT 119.865 195.745 120.035 196.755 ;
        RECT 120.205 195.960 120.535 196.805 ;
        RECT 120.765 195.915 121.150 196.885 ;
        RECT 121.320 196.595 121.770 197.055 ;
        RECT 121.940 196.765 123.035 197.325 ;
        RECT 121.320 196.375 122.445 196.595 ;
        RECT 121.320 195.745 121.645 196.205 ;
        RECT 122.165 195.915 122.445 196.375 ;
        RECT 122.635 195.915 123.035 196.765 ;
        RECT 123.205 197.495 124.160 197.665 ;
        RECT 124.445 197.545 125.655 198.295 ;
        RECT 125.825 197.570 126.115 198.295 ;
        RECT 126.530 197.815 126.830 198.295 ;
        RECT 127.000 197.645 127.260 198.100 ;
        RECT 127.430 197.815 127.690 198.295 ;
        RECT 127.860 197.645 128.120 198.100 ;
        RECT 128.290 197.815 128.550 198.295 ;
        RECT 128.720 197.645 128.980 198.100 ;
        RECT 129.150 197.815 129.410 198.295 ;
        RECT 129.580 197.645 129.840 198.100 ;
        RECT 130.010 197.770 130.270 198.295 ;
        RECT 123.205 196.595 123.415 197.495 ;
        RECT 123.585 196.765 124.275 197.325 ;
        RECT 124.445 197.005 124.965 197.545 ;
        RECT 126.530 197.475 129.840 197.645 ;
        RECT 125.135 196.835 125.655 197.375 ;
        RECT 123.205 196.375 124.160 196.595 ;
        RECT 123.435 195.745 123.705 196.205 ;
        RECT 123.875 195.915 124.160 196.375 ;
        RECT 124.445 195.745 125.655 196.835 ;
        RECT 125.825 195.745 126.115 196.910 ;
        RECT 126.530 196.885 127.500 197.475 ;
        RECT 130.440 197.305 130.690 198.115 ;
        RECT 130.870 197.835 131.115 198.295 ;
        RECT 131.345 197.835 131.905 198.125 ;
        RECT 132.075 197.835 132.325 198.295 ;
        RECT 127.670 197.055 130.690 197.305 ;
        RECT 130.860 197.055 131.175 197.665 ;
        RECT 126.530 196.645 129.840 196.885 ;
        RECT 126.535 195.745 126.830 196.475 ;
        RECT 127.000 195.920 127.260 196.645 ;
        RECT 127.430 195.745 127.690 196.475 ;
        RECT 127.860 195.920 128.120 196.645 ;
        RECT 128.290 195.745 128.550 196.475 ;
        RECT 128.720 195.920 128.980 196.645 ;
        RECT 129.150 195.745 129.410 196.475 ;
        RECT 129.580 195.920 129.840 196.645 ;
        RECT 130.010 195.745 130.270 196.855 ;
        RECT 130.440 195.920 130.690 197.055 ;
        RECT 130.870 195.745 131.165 196.855 ;
        RECT 131.345 196.465 131.595 197.835 ;
        RECT 132.945 197.665 133.275 198.025 ;
        RECT 131.885 197.475 133.275 197.665 ;
        RECT 133.645 197.525 136.235 198.295 ;
        RECT 137.030 197.785 137.270 198.295 ;
        RECT 137.450 197.785 137.730 198.115 ;
        RECT 137.960 197.785 138.175 198.295 ;
        RECT 131.885 197.385 132.055 197.475 ;
        RECT 131.765 197.055 132.055 197.385 ;
        RECT 132.225 197.055 132.565 197.305 ;
        RECT 132.785 197.055 133.460 197.305 ;
        RECT 131.885 196.805 132.055 197.055 ;
        RECT 131.885 196.635 132.825 196.805 ;
        RECT 133.195 196.695 133.460 197.055 ;
        RECT 133.645 197.005 134.855 197.525 ;
        RECT 135.025 196.835 136.235 197.355 ;
        RECT 136.925 197.055 137.280 197.615 ;
        RECT 137.450 196.885 137.620 197.785 ;
        RECT 137.790 197.055 138.055 197.615 ;
        RECT 138.345 197.555 138.960 198.125 ;
        RECT 140.175 197.745 140.345 198.125 ;
        RECT 140.525 197.915 140.855 198.295 ;
        RECT 140.175 197.575 140.840 197.745 ;
        RECT 141.035 197.620 141.295 198.125 ;
        RECT 141.465 197.750 146.810 198.295 ;
        RECT 138.305 196.885 138.475 197.385 ;
        RECT 131.345 195.915 131.805 196.465 ;
        RECT 131.995 195.745 132.325 196.465 ;
        RECT 132.525 196.085 132.825 196.635 ;
        RECT 132.995 195.745 133.275 196.415 ;
        RECT 133.645 195.745 136.235 196.835 ;
        RECT 137.050 196.715 138.475 196.885 ;
        RECT 137.050 196.540 137.440 196.715 ;
        RECT 137.925 195.745 138.255 196.545 ;
        RECT 138.645 196.535 138.960 197.555 ;
        RECT 140.105 197.025 140.435 197.395 ;
        RECT 140.670 197.320 140.840 197.575 ;
        RECT 140.670 196.990 140.955 197.320 ;
        RECT 140.670 196.845 140.840 196.990 ;
        RECT 138.425 195.915 138.960 196.535 ;
        RECT 140.175 196.675 140.840 196.845 ;
        RECT 141.125 196.820 141.295 197.620 ;
        RECT 143.050 196.920 143.390 197.750 ;
        RECT 146.985 197.495 147.295 198.295 ;
        RECT 147.500 197.495 148.195 198.125 ;
        RECT 148.365 197.525 150.955 198.295 ;
        RECT 151.585 197.570 151.875 198.295 ;
        RECT 152.045 197.525 155.555 198.295 ;
        RECT 155.725 197.545 156.935 198.295 ;
        RECT 140.175 195.915 140.345 196.675 ;
        RECT 140.525 195.745 140.855 196.505 ;
        RECT 141.025 195.915 141.295 196.820 ;
        RECT 144.870 196.180 145.220 197.430 ;
        RECT 146.995 197.055 147.330 197.325 ;
        RECT 147.500 196.895 147.670 197.495 ;
        RECT 147.840 197.055 148.175 197.305 ;
        RECT 148.365 197.005 149.575 197.525 ;
        RECT 141.465 195.745 146.810 196.180 ;
        RECT 146.985 195.745 147.265 196.885 ;
        RECT 147.435 195.915 147.765 196.895 ;
        RECT 147.935 195.745 148.195 196.885 ;
        RECT 149.745 196.835 150.955 197.355 ;
        RECT 152.045 197.005 153.695 197.525 ;
        RECT 148.365 195.745 150.955 196.835 ;
        RECT 151.585 195.745 151.875 196.910 ;
        RECT 153.865 196.835 155.555 197.355 ;
        RECT 152.045 195.745 155.555 196.835 ;
        RECT 155.725 196.835 156.245 197.375 ;
        RECT 156.415 197.005 156.935 197.545 ;
        RECT 155.725 195.745 156.935 196.835 ;
        RECT 22.700 195.575 157.020 195.745 ;
        RECT 22.785 194.485 23.995 195.575 ;
        RECT 24.165 195.140 29.510 195.575 ;
        RECT 22.785 193.775 23.305 194.315 ;
        RECT 23.475 193.945 23.995 194.485 ;
        RECT 22.785 193.025 23.995 193.775 ;
        RECT 25.750 193.570 26.090 194.400 ;
        RECT 27.570 193.890 27.920 195.140 ;
        RECT 29.685 194.485 32.275 195.575 ;
        RECT 29.685 193.795 30.895 194.315 ;
        RECT 31.065 193.965 32.275 194.485 ;
        RECT 32.940 194.785 33.475 195.405 ;
        RECT 24.165 193.025 29.510 193.570 ;
        RECT 29.685 193.025 32.275 193.795 ;
        RECT 32.940 193.765 33.255 194.785 ;
        RECT 33.645 194.775 33.975 195.575 ;
        RECT 34.460 194.605 34.850 194.780 ;
        RECT 33.425 194.435 34.850 194.605 ;
        RECT 33.425 193.935 33.595 194.435 ;
        RECT 32.940 193.195 33.555 193.765 ;
        RECT 33.845 193.705 34.110 194.265 ;
        RECT 34.280 193.535 34.450 194.435 ;
        RECT 35.665 194.410 35.955 195.575 ;
        RECT 36.215 194.645 36.385 195.405 ;
        RECT 36.565 194.815 36.895 195.575 ;
        RECT 36.215 194.475 36.880 194.645 ;
        RECT 37.065 194.500 37.335 195.405 ;
        RECT 36.710 194.330 36.880 194.475 ;
        RECT 34.620 193.705 34.975 194.265 ;
        RECT 36.145 193.925 36.475 194.295 ;
        RECT 36.710 194.000 36.995 194.330 ;
        RECT 33.725 193.025 33.940 193.535 ;
        RECT 34.170 193.205 34.450 193.535 ;
        RECT 34.630 193.025 34.870 193.535 ;
        RECT 35.665 193.025 35.955 193.750 ;
        RECT 36.710 193.745 36.880 194.000 ;
        RECT 36.215 193.575 36.880 193.745 ;
        RECT 37.165 193.700 37.335 194.500 ;
        RECT 37.505 194.485 39.175 195.575 ;
        RECT 36.215 193.195 36.385 193.575 ;
        RECT 36.565 193.025 36.895 193.405 ;
        RECT 37.075 193.195 37.335 193.700 ;
        RECT 37.505 193.795 38.255 194.315 ;
        RECT 38.425 193.965 39.175 194.485 ;
        RECT 39.345 194.500 39.615 195.405 ;
        RECT 39.785 194.815 40.115 195.575 ;
        RECT 40.295 194.645 40.465 195.405 ;
        RECT 40.725 195.140 46.070 195.575 ;
        RECT 37.505 193.025 39.175 193.795 ;
        RECT 39.345 193.700 39.515 194.500 ;
        RECT 39.800 194.475 40.465 194.645 ;
        RECT 39.800 194.330 39.970 194.475 ;
        RECT 39.685 194.000 39.970 194.330 ;
        RECT 39.800 193.745 39.970 194.000 ;
        RECT 40.205 193.925 40.535 194.295 ;
        RECT 39.345 193.195 39.605 193.700 ;
        RECT 39.800 193.575 40.465 193.745 ;
        RECT 39.785 193.025 40.115 193.405 ;
        RECT 40.295 193.195 40.465 193.575 ;
        RECT 42.310 193.570 42.650 194.400 ;
        RECT 44.130 193.890 44.480 195.140 ;
        RECT 46.245 194.485 47.455 195.575 ;
        RECT 46.245 193.775 46.765 194.315 ;
        RECT 46.935 193.945 47.455 194.485 ;
        RECT 47.665 194.435 47.895 195.575 ;
        RECT 48.065 194.425 48.395 195.405 ;
        RECT 48.565 194.435 48.775 195.575 ;
        RECT 49.010 194.435 49.265 195.575 ;
        RECT 49.460 195.025 50.655 195.355 ;
        RECT 47.645 194.015 47.975 194.265 ;
        RECT 40.725 193.025 46.070 193.570 ;
        RECT 46.245 193.025 47.455 193.775 ;
        RECT 47.665 193.025 47.895 193.845 ;
        RECT 48.145 193.825 48.395 194.425 ;
        RECT 49.515 194.265 49.685 194.825 ;
        RECT 49.910 194.605 50.330 194.855 ;
        RECT 50.835 194.775 51.115 195.575 ;
        RECT 49.910 194.435 51.155 194.605 ;
        RECT 51.325 194.435 51.595 195.405 ;
        RECT 50.985 194.265 51.155 194.435 ;
        RECT 49.010 194.015 49.345 194.265 ;
        RECT 49.515 193.935 50.255 194.265 ;
        RECT 50.985 193.935 51.215 194.265 ;
        RECT 49.515 193.845 49.765 193.935 ;
        RECT 48.065 193.195 48.395 193.825 ;
        RECT 48.565 193.025 48.775 193.845 ;
        RECT 49.030 193.675 49.765 193.845 ;
        RECT 50.985 193.765 51.155 193.935 ;
        RECT 49.030 193.205 49.340 193.675 ;
        RECT 50.415 193.595 51.155 193.765 ;
        RECT 51.425 193.700 51.595 194.435 ;
        RECT 49.510 193.025 50.245 193.505 ;
        RECT 50.415 193.245 50.585 193.595 ;
        RECT 50.755 193.025 51.135 193.425 ;
        RECT 51.325 193.355 51.595 193.700 ;
        RECT 51.765 194.605 52.075 195.405 ;
        RECT 52.245 194.775 52.555 195.575 ;
        RECT 52.725 194.945 52.985 195.405 ;
        RECT 53.155 195.115 53.410 195.575 ;
        RECT 53.585 194.945 53.845 195.405 ;
        RECT 52.725 194.775 53.845 194.945 ;
        RECT 51.765 194.435 52.795 194.605 ;
        RECT 51.765 193.525 51.935 194.435 ;
        RECT 52.105 193.695 52.455 194.265 ;
        RECT 52.625 194.185 52.795 194.435 ;
        RECT 53.585 194.525 53.845 194.775 ;
        RECT 54.015 194.705 54.300 195.575 ;
        RECT 53.585 194.355 54.340 194.525 ;
        RECT 52.625 194.015 53.765 194.185 ;
        RECT 53.935 193.845 54.340 194.355 ;
        RECT 52.690 193.675 54.340 193.845 ;
        RECT 54.525 194.500 54.795 195.405 ;
        RECT 54.965 194.815 55.295 195.575 ;
        RECT 55.475 194.645 55.645 195.405 ;
        RECT 54.525 193.700 54.695 194.500 ;
        RECT 54.980 194.475 55.645 194.645 ;
        RECT 55.905 194.485 57.575 195.575 ;
        RECT 54.980 194.330 55.150 194.475 ;
        RECT 54.865 194.000 55.150 194.330 ;
        RECT 54.980 193.745 55.150 194.000 ;
        RECT 55.385 193.925 55.715 194.295 ;
        RECT 55.905 193.795 56.655 194.315 ;
        RECT 56.825 193.965 57.575 194.485 ;
        RECT 58.225 194.685 58.485 195.395 ;
        RECT 58.655 194.865 58.985 195.575 ;
        RECT 59.155 194.685 59.385 195.395 ;
        RECT 58.225 194.445 59.385 194.685 ;
        RECT 59.565 194.665 59.835 195.395 ;
        RECT 60.015 194.845 60.355 195.575 ;
        RECT 59.565 194.445 60.335 194.665 ;
        RECT 58.215 193.935 58.515 194.265 ;
        RECT 58.695 193.955 59.220 194.265 ;
        RECT 59.400 193.955 59.865 194.265 ;
        RECT 51.765 193.195 52.065 193.525 ;
        RECT 52.235 193.025 52.510 193.505 ;
        RECT 52.690 193.285 52.985 193.675 ;
        RECT 53.155 193.025 53.410 193.505 ;
        RECT 53.585 193.285 53.845 193.675 ;
        RECT 54.015 193.025 54.295 193.505 ;
        RECT 54.525 193.195 54.785 193.700 ;
        RECT 54.980 193.575 55.645 193.745 ;
        RECT 54.965 193.025 55.295 193.405 ;
        RECT 55.475 193.195 55.645 193.575 ;
        RECT 55.905 193.025 57.575 193.795 ;
        RECT 58.225 193.025 58.515 193.755 ;
        RECT 58.695 193.315 58.925 193.955 ;
        RECT 60.045 193.775 60.335 194.445 ;
        RECT 59.105 193.575 60.335 193.775 ;
        RECT 59.105 193.205 59.415 193.575 ;
        RECT 59.595 193.025 60.265 193.395 ;
        RECT 60.525 193.205 60.785 195.395 ;
        RECT 61.425 194.410 61.715 195.575 ;
        RECT 61.885 194.485 64.475 195.575 ;
        RECT 61.885 193.795 63.095 194.315 ;
        RECT 63.265 193.965 64.475 194.485 ;
        RECT 64.655 194.465 64.950 195.575 ;
        RECT 65.130 194.265 65.380 195.400 ;
        RECT 65.550 194.465 65.810 195.575 ;
        RECT 65.980 194.675 66.240 195.400 ;
        RECT 66.410 194.845 66.670 195.575 ;
        RECT 66.840 194.675 67.100 195.400 ;
        RECT 67.270 194.845 67.530 195.575 ;
        RECT 67.700 194.675 67.960 195.400 ;
        RECT 68.130 194.845 68.390 195.575 ;
        RECT 68.560 194.675 68.820 195.400 ;
        RECT 68.990 194.845 69.285 195.575 ;
        RECT 69.705 194.705 69.980 195.405 ;
        RECT 70.190 195.030 70.405 195.575 ;
        RECT 70.575 195.065 71.050 195.405 ;
        RECT 71.220 195.070 71.835 195.575 ;
        RECT 71.220 194.895 71.415 195.070 ;
        RECT 65.980 194.435 69.290 194.675 ;
        RECT 61.425 193.025 61.715 193.750 ;
        RECT 61.885 193.025 64.475 193.795 ;
        RECT 64.645 193.655 64.960 194.265 ;
        RECT 65.130 194.015 68.150 194.265 ;
        RECT 64.705 193.025 64.950 193.485 ;
        RECT 65.130 193.205 65.380 194.015 ;
        RECT 68.320 193.845 69.290 194.435 ;
        RECT 65.980 193.675 69.290 193.845 ;
        RECT 69.705 193.675 69.875 194.705 ;
        RECT 70.150 194.535 70.865 194.830 ;
        RECT 71.085 194.705 71.415 194.895 ;
        RECT 71.585 194.535 71.835 194.900 ;
        RECT 70.045 194.365 71.835 194.535 ;
        RECT 70.045 193.935 70.275 194.365 ;
        RECT 65.550 193.025 65.810 193.550 ;
        RECT 65.980 193.220 66.240 193.675 ;
        RECT 66.410 193.025 66.670 193.505 ;
        RECT 66.840 193.220 67.100 193.675 ;
        RECT 67.270 193.025 67.530 193.505 ;
        RECT 67.700 193.220 67.960 193.675 ;
        RECT 68.130 193.025 68.390 193.505 ;
        RECT 68.560 193.220 68.820 193.675 ;
        RECT 68.990 193.025 69.290 193.505 ;
        RECT 69.705 193.195 69.965 193.675 ;
        RECT 70.445 193.665 70.855 194.185 ;
        RECT 70.135 193.025 70.465 193.485 ;
        RECT 70.655 193.245 70.855 193.665 ;
        RECT 71.025 193.510 71.280 194.365 ;
        RECT 72.075 194.185 72.245 195.405 ;
        RECT 72.495 195.065 72.755 195.575 ;
        RECT 72.925 195.145 73.265 195.405 ;
        RECT 71.450 193.935 72.245 194.185 ;
        RECT 72.415 194.015 72.755 194.895 ;
        RECT 71.995 193.845 72.245 193.935 ;
        RECT 71.025 193.245 71.815 193.510 ;
        RECT 71.995 193.425 72.325 193.845 ;
        RECT 72.495 193.025 72.755 193.845 ;
        RECT 72.925 193.745 73.185 195.145 ;
        RECT 73.435 194.775 73.765 195.575 ;
        RECT 74.230 194.605 74.480 195.405 ;
        RECT 74.665 194.855 74.995 195.575 ;
        RECT 75.215 194.605 75.465 195.405 ;
        RECT 75.635 195.195 75.970 195.575 ;
        RECT 73.375 194.435 75.565 194.605 ;
        RECT 73.375 194.265 73.690 194.435 ;
        RECT 73.360 194.015 73.690 194.265 ;
        RECT 72.925 193.235 73.265 193.745 ;
        RECT 73.435 193.025 73.705 193.825 ;
        RECT 73.885 193.295 74.165 194.265 ;
        RECT 74.345 193.295 74.645 194.265 ;
        RECT 74.825 193.300 75.175 194.265 ;
        RECT 75.395 193.525 75.565 194.435 ;
        RECT 75.735 193.705 75.975 195.015 ;
        RECT 76.695 194.905 76.865 195.405 ;
        RECT 77.035 195.075 77.365 195.575 ;
        RECT 76.695 194.735 77.360 194.905 ;
        RECT 76.610 193.915 76.960 194.565 ;
        RECT 77.130 193.745 77.360 194.735 ;
        RECT 76.695 193.575 77.360 193.745 ;
        RECT 75.395 193.195 75.890 193.525 ;
        RECT 76.695 193.285 76.865 193.575 ;
        RECT 77.035 193.025 77.365 193.405 ;
        RECT 77.535 193.285 77.720 195.405 ;
        RECT 77.960 195.115 78.225 195.575 ;
        RECT 78.395 194.980 78.645 195.405 ;
        RECT 78.855 195.130 79.960 195.300 ;
        RECT 78.340 194.850 78.645 194.980 ;
        RECT 77.890 193.655 78.170 194.605 ;
        RECT 78.340 193.745 78.510 194.850 ;
        RECT 78.680 194.065 78.920 194.660 ;
        RECT 79.090 194.595 79.620 194.960 ;
        RECT 79.090 193.895 79.260 194.595 ;
        RECT 79.790 194.515 79.960 195.130 ;
        RECT 80.130 194.775 80.300 195.575 ;
        RECT 80.470 195.075 80.720 195.405 ;
        RECT 80.945 195.105 81.830 195.275 ;
        RECT 79.790 194.425 80.300 194.515 ;
        RECT 78.340 193.615 78.565 193.745 ;
        RECT 78.735 193.675 79.260 193.895 ;
        RECT 79.430 194.255 80.300 194.425 ;
        RECT 77.975 193.025 78.225 193.485 ;
        RECT 78.395 193.475 78.565 193.615 ;
        RECT 79.430 193.475 79.600 194.255 ;
        RECT 80.130 194.185 80.300 194.255 ;
        RECT 79.810 194.005 80.010 194.035 ;
        RECT 80.470 194.005 80.640 195.075 ;
        RECT 80.810 194.185 81.000 194.905 ;
        RECT 79.810 193.705 80.640 194.005 ;
        RECT 81.170 193.975 81.490 194.935 ;
        RECT 78.395 193.305 78.730 193.475 ;
        RECT 78.925 193.305 79.600 193.475 ;
        RECT 79.920 193.025 80.290 193.525 ;
        RECT 80.470 193.475 80.640 193.705 ;
        RECT 81.025 193.645 81.490 193.975 ;
        RECT 81.660 194.265 81.830 195.105 ;
        RECT 82.010 195.075 82.325 195.575 ;
        RECT 82.555 194.845 82.895 195.405 ;
        RECT 82.000 194.470 82.895 194.845 ;
        RECT 83.065 194.565 83.235 195.575 ;
        RECT 82.705 194.265 82.895 194.470 ;
        RECT 83.405 194.515 83.735 195.360 ;
        RECT 84.885 194.855 85.345 195.405 ;
        RECT 85.535 194.855 85.865 195.575 ;
        RECT 83.405 194.435 83.795 194.515 ;
        RECT 83.580 194.385 83.795 194.435 ;
        RECT 81.660 193.935 82.535 194.265 ;
        RECT 82.705 193.935 83.455 194.265 ;
        RECT 81.660 193.475 81.830 193.935 ;
        RECT 82.705 193.765 82.905 193.935 ;
        RECT 83.625 193.805 83.795 194.385 ;
        RECT 83.570 193.765 83.795 193.805 ;
        RECT 80.470 193.305 80.875 193.475 ;
        RECT 81.045 193.305 81.830 193.475 ;
        RECT 82.105 193.025 82.315 193.555 ;
        RECT 82.575 193.240 82.905 193.765 ;
        RECT 83.415 193.680 83.795 193.765 ;
        RECT 83.075 193.025 83.245 193.635 ;
        RECT 83.415 193.245 83.745 193.680 ;
        RECT 84.885 193.485 85.135 194.855 ;
        RECT 86.065 194.685 86.365 195.235 ;
        RECT 86.535 194.905 86.815 195.575 ;
        RECT 85.425 194.515 86.365 194.685 ;
        RECT 85.425 194.265 85.595 194.515 ;
        RECT 86.735 194.265 87.000 194.625 ;
        RECT 87.185 194.410 87.475 195.575 ;
        RECT 87.645 195.020 88.250 195.575 ;
        RECT 88.425 195.065 88.905 195.405 ;
        RECT 89.075 195.030 89.330 195.575 ;
        RECT 87.645 194.920 88.260 195.020 ;
        RECT 88.075 194.895 88.260 194.920 ;
        RECT 85.305 193.935 85.595 194.265 ;
        RECT 85.765 194.015 86.105 194.265 ;
        RECT 86.325 194.015 87.000 194.265 ;
        RECT 87.645 194.300 87.905 194.750 ;
        RECT 88.075 194.650 88.405 194.895 ;
        RECT 88.575 194.575 89.330 194.825 ;
        RECT 89.500 194.705 89.775 195.405 ;
        RECT 88.560 194.540 89.330 194.575 ;
        RECT 88.545 194.530 89.330 194.540 ;
        RECT 88.540 194.515 89.435 194.530 ;
        RECT 88.520 194.500 89.435 194.515 ;
        RECT 88.500 194.490 89.435 194.500 ;
        RECT 88.475 194.480 89.435 194.490 ;
        RECT 88.405 194.450 89.435 194.480 ;
        RECT 88.385 194.420 89.435 194.450 ;
        RECT 88.365 194.390 89.435 194.420 ;
        RECT 88.335 194.365 89.435 194.390 ;
        RECT 88.300 194.330 89.435 194.365 ;
        RECT 88.270 194.325 89.435 194.330 ;
        RECT 88.270 194.320 88.660 194.325 ;
        RECT 88.270 194.310 88.635 194.320 ;
        RECT 88.270 194.305 88.620 194.310 ;
        RECT 88.270 194.300 88.605 194.305 ;
        RECT 87.645 194.295 88.605 194.300 ;
        RECT 87.645 194.285 88.595 194.295 ;
        RECT 87.645 194.280 88.585 194.285 ;
        RECT 87.645 194.270 88.575 194.280 ;
        RECT 87.645 194.260 88.570 194.270 ;
        RECT 87.645 194.255 88.565 194.260 ;
        RECT 87.645 194.240 88.555 194.255 ;
        RECT 87.645 194.225 88.550 194.240 ;
        RECT 87.645 194.200 88.540 194.225 ;
        RECT 87.645 194.130 88.535 194.200 ;
        RECT 85.425 193.845 85.595 193.935 ;
        RECT 85.425 193.655 86.815 193.845 ;
        RECT 84.885 193.195 85.445 193.485 ;
        RECT 85.615 193.025 85.865 193.485 ;
        RECT 86.485 193.295 86.815 193.655 ;
        RECT 87.185 193.025 87.475 193.750 ;
        RECT 87.645 193.575 88.195 193.960 ;
        RECT 88.365 193.405 88.535 194.130 ;
        RECT 87.645 193.235 88.535 193.405 ;
        RECT 88.705 193.730 89.035 194.155 ;
        RECT 89.205 193.930 89.435 194.325 ;
        RECT 88.705 193.245 88.925 193.730 ;
        RECT 89.605 193.675 89.775 194.705 ;
        RECT 90.005 194.515 90.335 195.360 ;
        RECT 90.505 194.565 90.675 195.575 ;
        RECT 90.845 194.845 91.185 195.405 ;
        RECT 91.415 195.075 91.730 195.575 ;
        RECT 91.910 195.105 92.795 195.275 ;
        RECT 89.945 194.435 90.335 194.515 ;
        RECT 90.845 194.470 91.740 194.845 ;
        RECT 89.945 194.385 90.160 194.435 ;
        RECT 89.945 193.805 90.115 194.385 ;
        RECT 90.845 194.265 91.035 194.470 ;
        RECT 91.910 194.265 92.080 195.105 ;
        RECT 93.020 195.075 93.270 195.405 ;
        RECT 90.285 193.935 91.035 194.265 ;
        RECT 91.205 193.935 92.080 194.265 ;
        RECT 89.945 193.765 90.170 193.805 ;
        RECT 90.835 193.765 91.035 193.935 ;
        RECT 89.945 193.680 90.325 193.765 ;
        RECT 89.095 193.025 89.345 193.565 ;
        RECT 89.515 193.195 89.775 193.675 ;
        RECT 89.995 193.245 90.325 193.680 ;
        RECT 90.495 193.025 90.665 193.635 ;
        RECT 90.835 193.240 91.165 193.765 ;
        RECT 91.425 193.025 91.635 193.555 ;
        RECT 91.910 193.475 92.080 193.935 ;
        RECT 92.250 193.975 92.570 194.935 ;
        RECT 92.740 194.185 92.930 194.905 ;
        RECT 93.100 194.005 93.270 195.075 ;
        RECT 93.440 194.775 93.610 195.575 ;
        RECT 93.780 195.130 94.885 195.300 ;
        RECT 93.780 194.515 93.950 195.130 ;
        RECT 95.095 194.980 95.345 195.405 ;
        RECT 95.515 195.115 95.780 195.575 ;
        RECT 94.120 194.595 94.650 194.960 ;
        RECT 95.095 194.850 95.400 194.980 ;
        RECT 93.440 194.425 93.950 194.515 ;
        RECT 93.440 194.255 94.310 194.425 ;
        RECT 93.440 194.185 93.610 194.255 ;
        RECT 93.730 194.005 93.930 194.035 ;
        RECT 92.250 193.645 92.715 193.975 ;
        RECT 93.100 193.705 93.930 194.005 ;
        RECT 93.100 193.475 93.270 193.705 ;
        RECT 91.910 193.305 92.695 193.475 ;
        RECT 92.865 193.305 93.270 193.475 ;
        RECT 93.450 193.025 93.820 193.525 ;
        RECT 94.140 193.475 94.310 194.255 ;
        RECT 94.480 193.895 94.650 194.595 ;
        RECT 94.820 194.065 95.060 194.660 ;
        RECT 94.480 193.675 95.005 193.895 ;
        RECT 95.230 193.745 95.400 194.850 ;
        RECT 95.175 193.615 95.400 193.745 ;
        RECT 95.570 193.655 95.850 194.605 ;
        RECT 95.175 193.475 95.345 193.615 ;
        RECT 94.140 193.305 94.815 193.475 ;
        RECT 95.010 193.305 95.345 193.475 ;
        RECT 95.515 193.025 95.765 193.485 ;
        RECT 96.020 193.285 96.205 195.405 ;
        RECT 96.375 195.075 96.705 195.575 ;
        RECT 96.875 194.905 97.045 195.405 ;
        RECT 96.380 194.735 97.045 194.905 ;
        RECT 97.880 194.945 98.165 195.405 ;
        RECT 98.335 195.115 98.605 195.575 ;
        RECT 96.380 193.745 96.610 194.735 ;
        RECT 97.880 194.725 98.835 194.945 ;
        RECT 96.780 193.915 97.130 194.565 ;
        RECT 97.765 193.995 98.455 194.555 ;
        RECT 98.625 193.825 98.835 194.725 ;
        RECT 96.380 193.575 97.045 193.745 ;
        RECT 96.375 193.025 96.705 193.405 ;
        RECT 96.875 193.285 97.045 193.575 ;
        RECT 97.880 193.655 98.835 193.825 ;
        RECT 99.005 194.555 99.405 195.405 ;
        RECT 99.595 194.945 99.875 195.405 ;
        RECT 100.395 195.115 100.720 195.575 ;
        RECT 99.595 194.725 100.720 194.945 ;
        RECT 99.005 193.995 100.100 194.555 ;
        RECT 100.270 194.265 100.720 194.725 ;
        RECT 100.890 194.435 101.275 195.405 ;
        RECT 101.535 194.905 101.705 195.405 ;
        RECT 101.875 195.075 102.205 195.575 ;
        RECT 101.535 194.735 102.200 194.905 ;
        RECT 97.880 193.195 98.165 193.655 ;
        RECT 98.335 193.025 98.605 193.485 ;
        RECT 99.005 193.195 99.405 193.995 ;
        RECT 100.270 193.935 100.825 194.265 ;
        RECT 100.270 193.825 100.720 193.935 ;
        RECT 99.595 193.655 100.720 193.825 ;
        RECT 100.995 193.765 101.275 194.435 ;
        RECT 101.450 193.915 101.800 194.565 ;
        RECT 99.595 193.195 99.875 193.655 ;
        RECT 100.395 193.025 100.720 193.485 ;
        RECT 100.890 193.195 101.275 193.765 ;
        RECT 101.970 193.745 102.200 194.735 ;
        RECT 101.535 193.575 102.200 193.745 ;
        RECT 101.535 193.285 101.705 193.575 ;
        RECT 101.875 193.025 102.205 193.405 ;
        RECT 102.375 193.285 102.560 195.405 ;
        RECT 102.800 195.115 103.065 195.575 ;
        RECT 103.235 194.980 103.485 195.405 ;
        RECT 103.695 195.130 104.800 195.300 ;
        RECT 103.180 194.850 103.485 194.980 ;
        RECT 102.730 193.655 103.010 194.605 ;
        RECT 103.180 193.745 103.350 194.850 ;
        RECT 103.520 194.065 103.760 194.660 ;
        RECT 103.930 194.595 104.460 194.960 ;
        RECT 103.930 193.895 104.100 194.595 ;
        RECT 104.630 194.515 104.800 195.130 ;
        RECT 104.970 194.775 105.140 195.575 ;
        RECT 105.310 195.075 105.560 195.405 ;
        RECT 105.785 195.105 106.670 195.275 ;
        RECT 104.630 194.425 105.140 194.515 ;
        RECT 103.180 193.615 103.405 193.745 ;
        RECT 103.575 193.675 104.100 193.895 ;
        RECT 104.270 194.255 105.140 194.425 ;
        RECT 102.815 193.025 103.065 193.485 ;
        RECT 103.235 193.475 103.405 193.615 ;
        RECT 104.270 193.475 104.440 194.255 ;
        RECT 104.970 194.185 105.140 194.255 ;
        RECT 104.650 194.005 104.850 194.035 ;
        RECT 105.310 194.005 105.480 195.075 ;
        RECT 105.650 194.185 105.840 194.905 ;
        RECT 104.650 193.705 105.480 194.005 ;
        RECT 106.010 193.975 106.330 194.935 ;
        RECT 103.235 193.305 103.570 193.475 ;
        RECT 103.765 193.305 104.440 193.475 ;
        RECT 104.760 193.025 105.130 193.525 ;
        RECT 105.310 193.475 105.480 193.705 ;
        RECT 105.865 193.645 106.330 193.975 ;
        RECT 106.500 194.265 106.670 195.105 ;
        RECT 106.850 195.075 107.165 195.575 ;
        RECT 107.395 194.845 107.735 195.405 ;
        RECT 106.840 194.470 107.735 194.845 ;
        RECT 107.905 194.565 108.075 195.575 ;
        RECT 107.545 194.265 107.735 194.470 ;
        RECT 108.245 194.515 108.575 195.360 ;
        RECT 108.920 194.945 109.205 195.405 ;
        RECT 109.375 195.115 109.645 195.575 ;
        RECT 108.920 194.725 109.875 194.945 ;
        RECT 108.245 194.435 108.635 194.515 ;
        RECT 108.420 194.385 108.635 194.435 ;
        RECT 106.500 193.935 107.375 194.265 ;
        RECT 107.545 193.935 108.295 194.265 ;
        RECT 106.500 193.475 106.670 193.935 ;
        RECT 107.545 193.765 107.745 193.935 ;
        RECT 108.465 193.805 108.635 194.385 ;
        RECT 108.805 193.995 109.495 194.555 ;
        RECT 109.665 193.825 109.875 194.725 ;
        RECT 108.410 193.765 108.635 193.805 ;
        RECT 105.310 193.305 105.715 193.475 ;
        RECT 105.885 193.305 106.670 193.475 ;
        RECT 106.945 193.025 107.155 193.555 ;
        RECT 107.415 193.240 107.745 193.765 ;
        RECT 108.255 193.680 108.635 193.765 ;
        RECT 107.915 193.025 108.085 193.635 ;
        RECT 108.255 193.245 108.585 193.680 ;
        RECT 108.920 193.655 109.875 193.825 ;
        RECT 110.045 194.555 110.445 195.405 ;
        RECT 110.635 194.945 110.915 195.405 ;
        RECT 111.435 195.115 111.760 195.575 ;
        RECT 110.635 194.725 111.760 194.945 ;
        RECT 110.045 193.995 111.140 194.555 ;
        RECT 111.310 194.265 111.760 194.725 ;
        RECT 111.930 194.435 112.315 195.405 ;
        RECT 108.920 193.195 109.205 193.655 ;
        RECT 109.375 193.025 109.645 193.485 ;
        RECT 110.045 193.195 110.445 193.995 ;
        RECT 111.310 193.935 111.865 194.265 ;
        RECT 111.310 193.825 111.760 193.935 ;
        RECT 110.635 193.655 111.760 193.825 ;
        RECT 112.035 193.765 112.315 194.435 ;
        RECT 112.945 194.410 113.235 195.575 ;
        RECT 113.405 194.725 113.665 195.405 ;
        RECT 113.835 194.795 114.085 195.575 ;
        RECT 114.335 195.025 114.585 195.405 ;
        RECT 114.755 195.195 115.110 195.575 ;
        RECT 116.115 195.185 116.450 195.405 ;
        RECT 115.715 195.025 115.945 195.065 ;
        RECT 114.335 194.825 115.945 195.025 ;
        RECT 114.335 194.815 115.170 194.825 ;
        RECT 115.760 194.735 115.945 194.825 ;
        RECT 110.635 193.195 110.915 193.655 ;
        RECT 111.435 193.025 111.760 193.485 ;
        RECT 111.930 193.195 112.315 193.765 ;
        RECT 112.945 193.025 113.235 193.750 ;
        RECT 113.405 193.525 113.575 194.725 ;
        RECT 115.275 194.625 115.605 194.655 ;
        RECT 113.805 194.565 115.605 194.625 ;
        RECT 116.195 194.565 116.450 195.185 ;
        RECT 113.745 194.455 116.450 194.565 ;
        RECT 116.625 194.485 120.135 195.575 ;
        RECT 113.745 194.420 113.945 194.455 ;
        RECT 113.745 193.845 113.915 194.420 ;
        RECT 115.275 194.395 116.450 194.455 ;
        RECT 114.145 193.980 114.555 194.285 ;
        RECT 114.725 194.015 115.055 194.225 ;
        RECT 113.745 193.725 114.015 193.845 ;
        RECT 113.745 193.680 114.590 193.725 ;
        RECT 113.835 193.555 114.590 193.680 ;
        RECT 114.845 193.615 115.055 194.015 ;
        RECT 115.300 194.015 115.775 194.225 ;
        RECT 115.965 194.015 116.455 194.215 ;
        RECT 115.300 193.615 115.520 194.015 ;
        RECT 116.625 193.795 118.275 194.315 ;
        RECT 118.445 193.965 120.135 194.485 ;
        RECT 120.770 194.435 121.025 195.575 ;
        RECT 121.220 195.025 122.415 195.355 ;
        RECT 121.275 194.265 121.445 194.825 ;
        RECT 121.670 194.605 122.090 194.855 ;
        RECT 122.595 194.775 122.875 195.575 ;
        RECT 121.670 194.435 122.915 194.605 ;
        RECT 123.085 194.435 123.355 195.405 ;
        RECT 123.995 194.965 124.325 195.395 ;
        RECT 124.505 195.135 124.700 195.575 ;
        RECT 124.870 194.965 125.200 195.395 ;
        RECT 123.995 194.795 125.200 194.965 ;
        RECT 123.995 194.465 124.890 194.795 ;
        RECT 125.370 194.625 125.645 195.395 ;
        RECT 122.745 194.265 122.915 194.435 ;
        RECT 123.125 194.385 123.355 194.435 ;
        RECT 120.770 194.015 121.105 194.265 ;
        RECT 121.275 193.935 122.015 194.265 ;
        RECT 122.745 193.935 122.975 194.265 ;
        RECT 121.275 193.845 121.525 193.935 ;
        RECT 113.405 193.195 113.665 193.525 ;
        RECT 114.420 193.405 114.590 193.555 ;
        RECT 113.835 193.025 114.165 193.385 ;
        RECT 114.420 193.195 115.720 193.405 ;
        RECT 115.995 193.025 116.450 193.790 ;
        RECT 116.625 193.025 120.135 193.795 ;
        RECT 120.790 193.675 121.525 193.845 ;
        RECT 122.745 193.765 122.915 193.935 ;
        RECT 120.790 193.205 121.100 193.675 ;
        RECT 122.175 193.595 122.915 193.765 ;
        RECT 123.185 193.700 123.355 194.385 ;
        RECT 125.060 194.435 125.645 194.625 ;
        RECT 126.285 194.985 126.985 195.405 ;
        RECT 127.185 195.215 127.515 195.575 ;
        RECT 127.685 194.985 128.015 195.385 ;
        RECT 126.285 194.755 128.015 194.985 ;
        RECT 124.000 193.935 124.295 194.265 ;
        RECT 124.475 193.935 124.890 194.265 ;
        RECT 121.270 193.025 122.005 193.505 ;
        RECT 122.175 193.245 122.345 193.595 ;
        RECT 122.515 193.025 122.895 193.425 ;
        RECT 123.085 193.355 123.355 193.700 ;
        RECT 123.995 193.025 124.295 193.755 ;
        RECT 124.475 193.315 124.705 193.935 ;
        RECT 125.060 193.765 125.235 194.435 ;
        RECT 124.905 193.585 125.235 193.765 ;
        RECT 125.405 193.615 125.645 194.265 ;
        RECT 126.285 193.875 126.490 194.755 ;
        RECT 126.660 194.015 126.990 194.555 ;
        RECT 127.165 194.265 127.490 194.555 ;
        RECT 127.685 194.535 128.015 194.755 ;
        RECT 128.185 194.265 128.355 195.235 ;
        RECT 128.535 194.515 128.865 195.575 ;
        RECT 129.045 194.485 130.715 195.575 ;
        RECT 127.165 193.935 127.660 194.265 ;
        RECT 127.980 193.935 128.355 194.265 ;
        RECT 128.565 193.935 128.875 194.265 ;
        RECT 126.285 193.785 126.515 193.875 ;
        RECT 129.045 193.795 129.795 194.315 ;
        RECT 129.965 193.965 130.715 194.485 ;
        RECT 130.895 194.605 131.225 195.390 ;
        RECT 130.895 194.435 131.575 194.605 ;
        RECT 131.755 194.435 132.085 195.575 ;
        RECT 132.265 194.485 134.855 195.575 ;
        RECT 130.885 194.015 131.235 194.265 ;
        RECT 131.405 193.835 131.575 194.435 ;
        RECT 131.745 194.015 132.095 194.265 ;
        RECT 124.905 193.205 125.130 193.585 ;
        RECT 125.300 193.025 125.630 193.415 ;
        RECT 126.285 193.195 126.995 193.785 ;
        RECT 127.505 193.555 128.865 193.765 ;
        RECT 127.505 193.195 127.835 193.555 ;
        RECT 128.035 193.025 128.365 193.385 ;
        RECT 128.535 193.195 128.865 193.555 ;
        RECT 129.045 193.025 130.715 193.795 ;
        RECT 130.905 193.025 131.145 193.835 ;
        RECT 131.315 193.195 131.645 193.835 ;
        RECT 131.815 193.025 132.085 193.835 ;
        RECT 132.265 193.795 133.475 194.315 ;
        RECT 133.645 193.965 134.855 194.485 ;
        RECT 135.025 194.435 135.285 195.575 ;
        RECT 135.455 194.425 135.785 195.405 ;
        RECT 135.955 194.435 136.235 195.575 ;
        RECT 136.590 194.605 136.980 194.780 ;
        RECT 137.465 194.775 137.795 195.575 ;
        RECT 137.965 194.785 138.500 195.405 ;
        RECT 136.590 194.435 138.015 194.605 ;
        RECT 135.545 194.385 135.720 194.425 ;
        RECT 135.045 194.015 135.380 194.265 ;
        RECT 135.550 193.825 135.720 194.385 ;
        RECT 135.890 193.995 136.225 194.265 ;
        RECT 132.265 193.025 134.855 193.795 ;
        RECT 135.025 193.195 135.720 193.825 ;
        RECT 135.925 193.025 136.235 193.825 ;
        RECT 136.465 193.705 136.820 194.265 ;
        RECT 136.990 193.535 137.160 194.435 ;
        RECT 137.330 193.705 137.595 194.265 ;
        RECT 137.845 193.935 138.015 194.435 ;
        RECT 138.185 193.765 138.500 194.785 ;
        RECT 138.705 194.410 138.995 195.575 ;
        RECT 139.165 194.705 139.440 195.405 ;
        RECT 139.610 195.030 139.865 195.575 ;
        RECT 140.035 195.065 140.515 195.405 ;
        RECT 140.690 195.020 141.295 195.575 ;
        RECT 140.680 194.920 141.295 195.020 ;
        RECT 140.680 194.895 140.865 194.920 ;
        RECT 136.570 193.025 136.810 193.535 ;
        RECT 136.990 193.205 137.270 193.535 ;
        RECT 137.500 193.025 137.715 193.535 ;
        RECT 137.885 193.195 138.500 193.765 ;
        RECT 138.705 193.025 138.995 193.750 ;
        RECT 139.165 193.675 139.335 194.705 ;
        RECT 139.610 194.575 140.365 194.825 ;
        RECT 140.535 194.650 140.865 194.895 ;
        RECT 139.610 194.540 140.380 194.575 ;
        RECT 139.610 194.530 140.395 194.540 ;
        RECT 139.505 194.515 140.400 194.530 ;
        RECT 139.505 194.500 140.420 194.515 ;
        RECT 139.505 194.490 140.440 194.500 ;
        RECT 139.505 194.480 140.465 194.490 ;
        RECT 139.505 194.450 140.535 194.480 ;
        RECT 139.505 194.420 140.555 194.450 ;
        RECT 139.505 194.390 140.575 194.420 ;
        RECT 139.505 194.365 140.605 194.390 ;
        RECT 139.505 194.330 140.640 194.365 ;
        RECT 139.505 194.325 140.670 194.330 ;
        RECT 139.505 193.930 139.735 194.325 ;
        RECT 140.280 194.320 140.670 194.325 ;
        RECT 140.305 194.310 140.670 194.320 ;
        RECT 140.320 194.305 140.670 194.310 ;
        RECT 140.335 194.300 140.670 194.305 ;
        RECT 141.035 194.300 141.295 194.750 ;
        RECT 140.335 194.295 141.295 194.300 ;
        RECT 140.345 194.285 141.295 194.295 ;
        RECT 140.355 194.280 141.295 194.285 ;
        RECT 140.365 194.270 141.295 194.280 ;
        RECT 140.370 194.260 141.295 194.270 ;
        RECT 140.375 194.255 141.295 194.260 ;
        RECT 140.385 194.240 141.295 194.255 ;
        RECT 140.390 194.225 141.295 194.240 ;
        RECT 140.400 194.200 141.295 194.225 ;
        RECT 139.905 193.730 140.235 194.155 ;
        RECT 139.985 193.705 140.235 193.730 ;
        RECT 139.165 193.195 139.425 193.675 ;
        RECT 139.595 193.025 139.845 193.565 ;
        RECT 140.015 193.245 140.235 193.705 ;
        RECT 140.405 194.130 141.295 194.200 ;
        RECT 141.465 194.705 141.740 195.405 ;
        RECT 141.910 195.030 142.165 195.575 ;
        RECT 142.335 195.065 142.815 195.405 ;
        RECT 142.990 195.020 143.595 195.575 ;
        RECT 142.980 194.920 143.595 195.020 ;
        RECT 142.980 194.895 143.165 194.920 ;
        RECT 140.405 193.405 140.575 194.130 ;
        RECT 140.745 193.575 141.295 193.960 ;
        RECT 141.465 193.675 141.635 194.705 ;
        RECT 141.910 194.575 142.665 194.825 ;
        RECT 142.835 194.650 143.165 194.895 ;
        RECT 141.910 194.540 142.680 194.575 ;
        RECT 141.910 194.530 142.695 194.540 ;
        RECT 141.805 194.515 142.700 194.530 ;
        RECT 141.805 194.500 142.720 194.515 ;
        RECT 141.805 194.490 142.740 194.500 ;
        RECT 141.805 194.480 142.765 194.490 ;
        RECT 141.805 194.450 142.835 194.480 ;
        RECT 141.805 194.420 142.855 194.450 ;
        RECT 141.805 194.390 142.875 194.420 ;
        RECT 141.805 194.365 142.905 194.390 ;
        RECT 141.805 194.330 142.940 194.365 ;
        RECT 141.805 194.325 142.970 194.330 ;
        RECT 141.805 193.930 142.035 194.325 ;
        RECT 142.580 194.320 142.970 194.325 ;
        RECT 142.605 194.310 142.970 194.320 ;
        RECT 142.620 194.305 142.970 194.310 ;
        RECT 142.635 194.300 142.970 194.305 ;
        RECT 143.335 194.300 143.595 194.750 ;
        RECT 143.765 194.485 145.435 195.575 ;
        RECT 142.635 194.295 143.595 194.300 ;
        RECT 142.645 194.285 143.595 194.295 ;
        RECT 142.655 194.280 143.595 194.285 ;
        RECT 142.665 194.270 143.595 194.280 ;
        RECT 142.670 194.260 143.595 194.270 ;
        RECT 142.675 194.255 143.595 194.260 ;
        RECT 142.685 194.240 143.595 194.255 ;
        RECT 142.690 194.225 143.595 194.240 ;
        RECT 142.700 194.200 143.595 194.225 ;
        RECT 142.205 193.730 142.535 194.155 ;
        RECT 142.285 193.705 142.535 193.730 ;
        RECT 140.405 193.235 141.295 193.405 ;
        RECT 141.465 193.195 141.725 193.675 ;
        RECT 141.895 193.025 142.145 193.565 ;
        RECT 142.315 193.245 142.535 193.705 ;
        RECT 142.705 194.130 143.595 194.200 ;
        RECT 142.705 193.405 142.875 194.130 ;
        RECT 143.045 193.575 143.595 193.960 ;
        RECT 143.765 193.795 144.515 194.315 ;
        RECT 144.685 193.965 145.435 194.485 ;
        RECT 145.695 194.645 145.865 195.405 ;
        RECT 146.045 194.815 146.375 195.575 ;
        RECT 145.695 194.475 146.360 194.645 ;
        RECT 146.545 194.500 146.815 195.405 ;
        RECT 146.985 195.140 152.330 195.575 ;
        RECT 146.190 194.330 146.360 194.475 ;
        RECT 145.625 193.925 145.955 194.295 ;
        RECT 146.190 194.000 146.475 194.330 ;
        RECT 142.705 193.235 143.595 193.405 ;
        RECT 143.765 193.025 145.435 193.795 ;
        RECT 146.190 193.745 146.360 194.000 ;
        RECT 145.695 193.575 146.360 193.745 ;
        RECT 146.645 193.700 146.815 194.500 ;
        RECT 145.695 193.195 145.865 193.575 ;
        RECT 146.045 193.025 146.375 193.405 ;
        RECT 146.555 193.195 146.815 193.700 ;
        RECT 148.570 193.570 148.910 194.400 ;
        RECT 150.390 193.890 150.740 195.140 ;
        RECT 152.505 194.485 155.095 195.575 ;
        RECT 152.505 193.795 153.715 194.315 ;
        RECT 153.885 193.965 155.095 194.485 ;
        RECT 155.725 194.485 156.935 195.575 ;
        RECT 155.725 193.945 156.245 194.485 ;
        RECT 146.985 193.025 152.330 193.570 ;
        RECT 152.505 193.025 155.095 193.795 ;
        RECT 156.415 193.775 156.935 194.315 ;
        RECT 155.725 193.025 156.935 193.775 ;
        RECT 22.700 192.855 157.020 193.025 ;
        RECT 22.785 192.105 23.995 192.855 ;
        RECT 22.785 191.565 23.305 192.105 ;
        RECT 24.165 192.085 27.675 192.855 ;
        RECT 28.765 192.355 29.025 192.685 ;
        RECT 29.235 192.375 29.510 192.855 ;
        RECT 23.475 191.395 23.995 191.935 ;
        RECT 24.165 191.565 25.815 192.085 ;
        RECT 25.985 191.395 27.675 191.915 ;
        RECT 22.785 190.305 23.995 191.395 ;
        RECT 24.165 190.305 27.675 191.395 ;
        RECT 28.765 191.445 28.935 192.355 ;
        RECT 29.720 192.285 29.925 192.685 ;
        RECT 30.095 192.455 30.430 192.855 ;
        RECT 29.105 191.615 29.465 192.195 ;
        RECT 29.720 192.115 30.405 192.285 ;
        RECT 29.645 191.445 29.895 191.945 ;
        RECT 28.765 191.275 29.895 191.445 ;
        RECT 28.765 190.505 29.035 191.275 ;
        RECT 30.065 191.085 30.405 192.115 ;
        RECT 31.525 192.035 31.785 192.855 ;
        RECT 31.955 192.035 32.285 192.455 ;
        RECT 32.465 192.370 33.255 192.635 ;
        RECT 32.035 191.945 32.285 192.035 ;
        RECT 29.205 190.305 29.535 191.085 ;
        RECT 29.740 190.910 30.405 191.085 ;
        RECT 31.525 190.985 31.865 191.865 ;
        RECT 32.035 191.695 32.830 191.945 ;
        RECT 29.740 190.505 29.925 190.910 ;
        RECT 30.095 190.305 30.430 190.730 ;
        RECT 31.525 190.305 31.785 190.815 ;
        RECT 32.035 190.475 32.205 191.695 ;
        RECT 33.000 191.515 33.255 192.370 ;
        RECT 33.425 192.215 33.625 192.635 ;
        RECT 33.815 192.395 34.145 192.855 ;
        RECT 33.425 191.695 33.835 192.215 ;
        RECT 34.315 192.205 34.575 192.685 ;
        RECT 34.005 191.515 34.235 191.945 ;
        RECT 32.445 191.345 34.235 191.515 ;
        RECT 32.445 190.980 32.695 191.345 ;
        RECT 32.865 190.985 33.195 191.175 ;
        RECT 33.415 191.050 34.130 191.345 ;
        RECT 34.405 191.175 34.575 192.205 ;
        RECT 32.865 190.810 33.060 190.985 ;
        RECT 32.445 190.305 33.060 190.810 ;
        RECT 33.230 190.475 33.705 190.815 ;
        RECT 33.875 190.305 34.090 190.850 ;
        RECT 34.300 190.475 34.575 191.175 ;
        RECT 34.745 192.395 35.305 192.685 ;
        RECT 35.475 192.395 35.725 192.855 ;
        RECT 34.745 191.025 34.995 192.395 ;
        RECT 36.345 192.225 36.675 192.585 ;
        RECT 35.285 192.035 36.675 192.225 ;
        RECT 37.595 192.305 37.765 192.595 ;
        RECT 37.935 192.475 38.265 192.855 ;
        RECT 37.595 192.135 38.260 192.305 ;
        RECT 35.285 191.945 35.455 192.035 ;
        RECT 35.165 191.615 35.455 191.945 ;
        RECT 35.625 191.615 35.965 191.865 ;
        RECT 36.185 191.615 36.860 191.865 ;
        RECT 35.285 191.365 35.455 191.615 ;
        RECT 35.285 191.195 36.225 191.365 ;
        RECT 36.595 191.255 36.860 191.615 ;
        RECT 37.510 191.315 37.860 191.965 ;
        RECT 34.745 190.475 35.205 191.025 ;
        RECT 35.395 190.305 35.725 191.025 ;
        RECT 35.925 190.645 36.225 191.195 ;
        RECT 38.030 191.145 38.260 192.135 ;
        RECT 37.595 190.975 38.260 191.145 ;
        RECT 36.395 190.305 36.675 190.975 ;
        RECT 37.595 190.475 37.765 190.975 ;
        RECT 37.935 190.305 38.265 190.805 ;
        RECT 38.435 190.475 38.620 192.595 ;
        RECT 38.875 192.395 39.125 192.855 ;
        RECT 39.295 192.405 39.630 192.575 ;
        RECT 39.825 192.405 40.500 192.575 ;
        RECT 39.295 192.265 39.465 192.405 ;
        RECT 38.790 191.275 39.070 192.225 ;
        RECT 39.240 192.135 39.465 192.265 ;
        RECT 39.240 191.030 39.410 192.135 ;
        RECT 39.635 191.985 40.160 192.205 ;
        RECT 39.580 191.220 39.820 191.815 ;
        RECT 39.990 191.285 40.160 191.985 ;
        RECT 40.330 191.625 40.500 192.405 ;
        RECT 40.820 192.355 41.190 192.855 ;
        RECT 41.370 192.405 41.775 192.575 ;
        RECT 41.945 192.405 42.730 192.575 ;
        RECT 41.370 192.175 41.540 192.405 ;
        RECT 40.710 191.875 41.540 192.175 ;
        RECT 41.925 191.905 42.390 192.235 ;
        RECT 40.710 191.845 40.910 191.875 ;
        RECT 41.030 191.625 41.200 191.695 ;
        RECT 40.330 191.455 41.200 191.625 ;
        RECT 40.690 191.365 41.200 191.455 ;
        RECT 39.240 190.900 39.545 191.030 ;
        RECT 39.990 190.920 40.520 191.285 ;
        RECT 38.860 190.305 39.125 190.765 ;
        RECT 39.295 190.475 39.545 190.900 ;
        RECT 40.690 190.750 40.860 191.365 ;
        RECT 39.755 190.580 40.860 190.750 ;
        RECT 41.030 190.305 41.200 191.105 ;
        RECT 41.370 190.805 41.540 191.875 ;
        RECT 41.710 190.975 41.900 191.695 ;
        RECT 42.070 190.945 42.390 191.905 ;
        RECT 42.560 191.945 42.730 192.405 ;
        RECT 43.005 192.325 43.215 192.855 ;
        RECT 43.475 192.115 43.805 192.640 ;
        RECT 43.975 192.245 44.145 192.855 ;
        RECT 44.315 192.200 44.645 192.635 ;
        RECT 45.410 192.355 45.905 192.685 ;
        RECT 44.315 192.115 44.695 192.200 ;
        RECT 43.605 191.945 43.805 192.115 ;
        RECT 44.470 192.075 44.695 192.115 ;
        RECT 42.560 191.615 43.435 191.945 ;
        RECT 43.605 191.615 44.355 191.945 ;
        RECT 41.370 190.475 41.620 190.805 ;
        RECT 42.560 190.775 42.730 191.615 ;
        RECT 43.605 191.410 43.795 191.615 ;
        RECT 44.525 191.495 44.695 192.075 ;
        RECT 44.480 191.445 44.695 191.495 ;
        RECT 42.900 191.035 43.795 191.410 ;
        RECT 44.305 191.365 44.695 191.445 ;
        RECT 41.845 190.605 42.730 190.775 ;
        RECT 42.910 190.305 43.225 190.805 ;
        RECT 43.455 190.475 43.795 191.035 ;
        RECT 43.965 190.305 44.135 191.315 ;
        RECT 44.305 190.520 44.635 191.365 ;
        RECT 45.325 190.865 45.565 192.175 ;
        RECT 45.735 191.445 45.905 192.355 ;
        RECT 46.125 191.615 46.475 192.580 ;
        RECT 46.655 191.615 46.955 192.585 ;
        RECT 47.135 191.615 47.415 192.585 ;
        RECT 47.595 192.055 47.865 192.855 ;
        RECT 48.035 192.135 48.375 192.645 ;
        RECT 47.610 191.615 47.940 191.865 ;
        RECT 47.610 191.445 47.925 191.615 ;
        RECT 45.735 191.275 47.925 191.445 ;
        RECT 45.330 190.305 45.665 190.685 ;
        RECT 45.835 190.475 46.085 191.275 ;
        RECT 46.305 190.305 46.635 191.025 ;
        RECT 46.820 190.475 47.070 191.275 ;
        RECT 47.535 190.305 47.865 191.105 ;
        RECT 48.115 190.735 48.375 192.135 ;
        RECT 48.545 192.130 48.835 192.855 ;
        RECT 49.005 192.095 49.715 192.685 ;
        RECT 50.225 192.325 50.555 192.685 ;
        RECT 50.755 192.495 51.085 192.855 ;
        RECT 51.255 192.325 51.585 192.685 ;
        RECT 50.225 192.115 51.585 192.325 ;
        RECT 51.815 192.200 52.145 192.635 ;
        RECT 52.315 192.245 52.485 192.855 ;
        RECT 51.765 192.115 52.145 192.200 ;
        RECT 52.655 192.115 52.985 192.640 ;
        RECT 53.245 192.325 53.455 192.855 ;
        RECT 53.730 192.405 54.515 192.575 ;
        RECT 54.685 192.405 55.090 192.575 ;
        RECT 48.035 190.475 48.375 190.735 ;
        RECT 48.545 190.305 48.835 191.470 ;
        RECT 49.005 191.125 49.210 192.095 ;
        RECT 51.765 192.075 51.990 192.115 ;
        RECT 49.380 191.325 49.710 191.865 ;
        RECT 49.885 191.615 50.380 191.945 ;
        RECT 50.700 191.615 51.075 191.945 ;
        RECT 51.285 191.615 51.595 191.945 ;
        RECT 49.885 191.325 50.210 191.615 ;
        RECT 50.405 191.125 50.735 191.345 ;
        RECT 49.005 190.895 50.735 191.125 ;
        RECT 49.005 190.475 49.705 190.895 ;
        RECT 49.905 190.305 50.235 190.665 ;
        RECT 50.405 190.495 50.735 190.895 ;
        RECT 50.905 190.645 51.075 191.615 ;
        RECT 51.765 191.495 51.935 192.075 ;
        RECT 52.655 191.945 52.855 192.115 ;
        RECT 53.730 191.945 53.900 192.405 ;
        RECT 52.105 191.615 52.855 191.945 ;
        RECT 53.025 191.615 53.900 191.945 ;
        RECT 51.765 191.445 51.980 191.495 ;
        RECT 51.765 191.365 52.155 191.445 ;
        RECT 51.255 190.305 51.585 191.365 ;
        RECT 51.825 190.520 52.155 191.365 ;
        RECT 52.665 191.410 52.855 191.615 ;
        RECT 52.325 190.305 52.495 191.315 ;
        RECT 52.665 191.035 53.560 191.410 ;
        RECT 52.665 190.475 53.005 191.035 ;
        RECT 53.235 190.305 53.550 190.805 ;
        RECT 53.730 190.775 53.900 191.615 ;
        RECT 54.070 191.905 54.535 192.235 ;
        RECT 54.920 192.175 55.090 192.405 ;
        RECT 55.270 192.355 55.640 192.855 ;
        RECT 55.960 192.405 56.635 192.575 ;
        RECT 56.830 192.405 57.165 192.575 ;
        RECT 54.070 190.945 54.390 191.905 ;
        RECT 54.920 191.875 55.750 192.175 ;
        RECT 54.560 190.975 54.750 191.695 ;
        RECT 54.920 190.805 55.090 191.875 ;
        RECT 55.550 191.845 55.750 191.875 ;
        RECT 55.260 191.625 55.430 191.695 ;
        RECT 55.960 191.625 56.130 192.405 ;
        RECT 56.995 192.265 57.165 192.405 ;
        RECT 57.335 192.395 57.585 192.855 ;
        RECT 55.260 191.455 56.130 191.625 ;
        RECT 56.300 191.985 56.825 192.205 ;
        RECT 56.995 192.135 57.220 192.265 ;
        RECT 55.260 191.365 55.770 191.455 ;
        RECT 53.730 190.605 54.615 190.775 ;
        RECT 54.840 190.475 55.090 190.805 ;
        RECT 55.260 190.305 55.430 191.105 ;
        RECT 55.600 190.750 55.770 191.365 ;
        RECT 56.300 191.285 56.470 191.985 ;
        RECT 55.940 190.920 56.470 191.285 ;
        RECT 56.640 191.220 56.880 191.815 ;
        RECT 57.050 191.030 57.220 192.135 ;
        RECT 57.390 191.275 57.670 192.225 ;
        RECT 56.915 190.900 57.220 191.030 ;
        RECT 55.600 190.580 56.705 190.750 ;
        RECT 56.915 190.475 57.165 190.900 ;
        RECT 57.335 190.305 57.600 190.765 ;
        RECT 57.840 190.475 58.025 192.595 ;
        RECT 58.195 192.475 58.525 192.855 ;
        RECT 58.695 192.305 58.865 192.595 ;
        RECT 58.200 192.135 58.865 192.305 ;
        RECT 58.200 191.145 58.430 192.135 ;
        RECT 59.125 192.085 62.635 192.855 ;
        RECT 62.810 192.350 63.145 192.855 ;
        RECT 63.315 192.285 63.555 192.660 ;
        RECT 63.835 192.525 64.005 192.670 ;
        RECT 63.835 192.330 64.210 192.525 ;
        RECT 64.570 192.360 64.965 192.855 ;
        RECT 58.600 191.315 58.950 191.965 ;
        RECT 59.125 191.565 60.775 192.085 ;
        RECT 60.945 191.395 62.635 191.915 ;
        RECT 58.200 190.975 58.865 191.145 ;
        RECT 58.195 190.305 58.525 190.805 ;
        RECT 58.695 190.475 58.865 190.975 ;
        RECT 59.125 190.305 62.635 191.395 ;
        RECT 62.865 191.325 63.165 192.175 ;
        RECT 63.335 192.135 63.555 192.285 ;
        RECT 63.335 191.805 63.870 192.135 ;
        RECT 64.040 191.995 64.210 192.330 ;
        RECT 65.135 192.165 65.375 192.685 ;
        RECT 63.335 191.155 63.570 191.805 ;
        RECT 64.040 191.635 65.025 191.995 ;
        RECT 62.895 190.925 63.570 191.155 ;
        RECT 63.740 191.615 65.025 191.635 ;
        RECT 63.740 191.465 64.600 191.615 ;
        RECT 62.895 190.495 63.065 190.925 ;
        RECT 63.235 190.305 63.565 190.755 ;
        RECT 63.740 190.520 64.025 191.465 ;
        RECT 65.200 191.360 65.375 192.165 ;
        RECT 64.200 190.985 64.895 191.295 ;
        RECT 64.205 190.305 64.890 190.775 ;
        RECT 65.070 190.575 65.375 191.360 ;
        RECT 65.585 192.165 65.825 192.685 ;
        RECT 65.995 192.360 66.390 192.855 ;
        RECT 66.955 192.525 67.125 192.670 ;
        RECT 66.750 192.330 67.125 192.525 ;
        RECT 65.585 191.360 65.760 192.165 ;
        RECT 66.750 191.995 66.920 192.330 ;
        RECT 67.405 192.285 67.645 192.660 ;
        RECT 67.815 192.350 68.150 192.855 ;
        RECT 67.405 192.135 67.625 192.285 ;
        RECT 65.935 191.635 66.920 191.995 ;
        RECT 67.090 191.805 67.625 192.135 ;
        RECT 65.935 191.615 67.220 191.635 ;
        RECT 66.360 191.465 67.220 191.615 ;
        RECT 65.585 190.575 65.890 191.360 ;
        RECT 66.065 190.985 66.760 191.295 ;
        RECT 66.070 190.305 66.755 190.775 ;
        RECT 66.935 190.520 67.220 191.465 ;
        RECT 67.390 191.155 67.625 191.805 ;
        RECT 67.795 191.325 68.095 192.175 ;
        RECT 68.325 192.085 71.835 192.855 ;
        RECT 68.325 191.565 69.975 192.085 ;
        RECT 72.525 192.035 72.735 192.855 ;
        RECT 72.905 192.055 73.235 192.685 ;
        RECT 70.145 191.395 71.835 191.915 ;
        RECT 72.905 191.455 73.155 192.055 ;
        RECT 73.405 192.035 73.635 192.855 ;
        RECT 74.305 192.130 74.595 192.855 ;
        RECT 74.765 192.085 77.355 192.855 ;
        RECT 77.985 192.180 78.245 192.685 ;
        RECT 78.425 192.475 78.755 192.855 ;
        RECT 78.935 192.305 79.105 192.685 ;
        RECT 73.325 191.615 73.655 191.865 ;
        RECT 74.765 191.565 75.975 192.085 ;
        RECT 67.390 190.925 68.065 191.155 ;
        RECT 67.395 190.305 67.725 190.755 ;
        RECT 67.895 190.495 68.065 190.925 ;
        RECT 68.325 190.305 71.835 191.395 ;
        RECT 72.525 190.305 72.735 191.445 ;
        RECT 72.905 190.475 73.235 191.455 ;
        RECT 73.405 190.305 73.635 191.445 ;
        RECT 74.305 190.305 74.595 191.470 ;
        RECT 76.145 191.395 77.355 191.915 ;
        RECT 74.765 190.305 77.355 191.395 ;
        RECT 77.985 191.380 78.155 192.180 ;
        RECT 78.440 192.135 79.105 192.305 ;
        RECT 78.440 191.880 78.610 192.135 ;
        RECT 79.425 192.035 79.635 192.855 ;
        RECT 79.805 192.055 80.135 192.685 ;
        RECT 78.325 191.550 78.610 191.880 ;
        RECT 78.845 191.585 79.175 191.955 ;
        RECT 78.440 191.405 78.610 191.550 ;
        RECT 79.805 191.455 80.055 192.055 ;
        RECT 80.305 192.035 80.535 192.855 ;
        RECT 80.745 192.085 84.255 192.855 ;
        RECT 80.225 191.615 80.555 191.865 ;
        RECT 80.745 191.565 82.395 192.085 ;
        RECT 84.945 192.035 85.155 192.855 ;
        RECT 85.325 192.055 85.655 192.685 ;
        RECT 77.985 190.475 78.255 191.380 ;
        RECT 78.440 191.235 79.105 191.405 ;
        RECT 78.425 190.305 78.755 191.065 ;
        RECT 78.935 190.475 79.105 191.235 ;
        RECT 79.425 190.305 79.635 191.445 ;
        RECT 79.805 190.475 80.135 191.455 ;
        RECT 80.305 190.305 80.535 191.445 ;
        RECT 82.565 191.395 84.255 191.915 ;
        RECT 85.325 191.455 85.575 192.055 ;
        RECT 85.825 192.035 86.055 192.855 ;
        RECT 86.265 192.105 87.475 192.855 ;
        RECT 85.745 191.615 86.075 191.865 ;
        RECT 86.265 191.565 86.785 192.105 ;
        RECT 87.705 192.035 87.915 192.855 ;
        RECT 88.085 192.055 88.415 192.685 ;
        RECT 80.745 190.305 84.255 191.395 ;
        RECT 84.945 190.305 85.155 191.445 ;
        RECT 85.325 190.475 85.655 191.455 ;
        RECT 85.825 190.305 86.055 191.445 ;
        RECT 86.955 191.395 87.475 191.935 ;
        RECT 88.085 191.455 88.335 192.055 ;
        RECT 88.585 192.035 88.815 192.855 ;
        RECT 89.025 192.085 90.695 192.855 ;
        RECT 91.415 192.305 91.585 192.685 ;
        RECT 91.765 192.475 92.095 192.855 ;
        RECT 91.415 192.135 92.080 192.305 ;
        RECT 92.275 192.180 92.535 192.685 ;
        RECT 88.505 191.615 88.835 191.865 ;
        RECT 89.025 191.565 89.775 192.085 ;
        RECT 86.265 190.305 87.475 191.395 ;
        RECT 87.705 190.305 87.915 191.445 ;
        RECT 88.085 190.475 88.415 191.455 ;
        RECT 88.585 190.305 88.815 191.445 ;
        RECT 89.945 191.395 90.695 191.915 ;
        RECT 91.345 191.585 91.675 191.955 ;
        RECT 91.910 191.880 92.080 192.135 ;
        RECT 91.910 191.550 92.195 191.880 ;
        RECT 91.910 191.405 92.080 191.550 ;
        RECT 89.025 190.305 90.695 191.395 ;
        RECT 91.415 191.235 92.080 191.405 ;
        RECT 92.365 191.380 92.535 192.180 ;
        RECT 93.685 192.035 93.895 192.855 ;
        RECT 94.065 192.055 94.395 192.685 ;
        RECT 94.065 191.455 94.315 192.055 ;
        RECT 94.565 192.035 94.795 192.855 ;
        RECT 95.005 192.085 96.675 192.855 ;
        RECT 94.485 191.615 94.815 191.865 ;
        RECT 95.005 191.565 95.755 192.085 ;
        RECT 97.365 192.035 97.575 192.855 ;
        RECT 97.745 192.055 98.075 192.685 ;
        RECT 91.415 190.475 91.585 191.235 ;
        RECT 91.765 190.305 92.095 191.065 ;
        RECT 92.265 190.475 92.535 191.380 ;
        RECT 93.685 190.305 93.895 191.445 ;
        RECT 94.065 190.475 94.395 191.455 ;
        RECT 94.565 190.305 94.795 191.445 ;
        RECT 95.925 191.395 96.675 191.915 ;
        RECT 97.745 191.455 97.995 192.055 ;
        RECT 98.245 192.035 98.475 192.855 ;
        RECT 98.685 192.105 99.895 192.855 ;
        RECT 100.065 192.130 100.355 192.855 ;
        RECT 100.805 192.225 101.185 192.675 ;
        RECT 98.165 191.615 98.495 191.865 ;
        RECT 98.685 191.565 99.205 192.105 ;
        RECT 95.005 190.305 96.675 191.395 ;
        RECT 97.365 190.305 97.575 191.445 ;
        RECT 97.745 190.475 98.075 191.455 ;
        RECT 98.245 190.305 98.475 191.445 ;
        RECT 99.375 191.395 99.895 191.935 ;
        RECT 98.685 190.305 99.895 191.395 ;
        RECT 100.065 190.305 100.355 191.470 ;
        RECT 100.545 191.275 100.775 191.965 ;
        RECT 100.955 191.775 101.185 192.225 ;
        RECT 101.365 192.075 101.595 192.855 ;
        RECT 101.775 192.145 102.205 192.675 ;
        RECT 101.775 191.895 102.020 192.145 ;
        RECT 102.385 191.945 102.595 192.565 ;
        RECT 102.765 192.125 103.095 192.855 ;
        RECT 104.450 192.375 104.750 192.855 ;
        RECT 104.920 192.205 105.180 192.660 ;
        RECT 105.350 192.375 105.610 192.855 ;
        RECT 105.780 192.205 106.040 192.660 ;
        RECT 106.210 192.375 106.470 192.855 ;
        RECT 106.640 192.205 106.900 192.660 ;
        RECT 107.070 192.375 107.330 192.855 ;
        RECT 107.500 192.205 107.760 192.660 ;
        RECT 107.930 192.330 108.190 192.855 ;
        RECT 104.450 192.035 107.760 192.205 ;
        RECT 100.955 191.095 101.295 191.775 ;
        RECT 100.535 190.895 101.295 191.095 ;
        RECT 101.485 191.595 102.020 191.895 ;
        RECT 102.200 191.595 102.595 191.945 ;
        RECT 102.790 191.595 103.080 191.945 ;
        RECT 100.535 190.505 100.795 190.895 ;
        RECT 100.965 190.305 101.295 190.715 ;
        RECT 101.485 190.485 101.815 191.595 ;
        RECT 104.450 191.445 105.420 192.035 ;
        RECT 108.360 191.865 108.610 192.675 ;
        RECT 108.790 192.395 109.035 192.855 ;
        RECT 109.355 192.305 109.525 192.595 ;
        RECT 109.695 192.475 110.025 192.855 ;
        RECT 105.590 191.615 108.610 191.865 ;
        RECT 108.780 191.615 109.095 192.225 ;
        RECT 109.355 192.135 110.020 192.305 ;
        RECT 101.985 191.215 103.025 191.415 ;
        RECT 101.985 190.485 102.175 191.215 ;
        RECT 102.345 190.305 102.675 191.035 ;
        RECT 102.855 190.485 103.025 191.215 ;
        RECT 104.450 191.205 107.760 191.445 ;
        RECT 104.455 190.305 104.750 191.035 ;
        RECT 104.920 190.480 105.180 191.205 ;
        RECT 105.350 190.305 105.610 191.035 ;
        RECT 105.780 190.480 106.040 191.205 ;
        RECT 106.210 190.305 106.470 191.035 ;
        RECT 106.640 190.480 106.900 191.205 ;
        RECT 107.070 190.305 107.330 191.035 ;
        RECT 107.500 190.480 107.760 191.205 ;
        RECT 107.930 190.305 108.190 191.415 ;
        RECT 108.360 190.480 108.610 191.615 ;
        RECT 108.790 190.305 109.085 191.415 ;
        RECT 109.270 191.315 109.620 191.965 ;
        RECT 109.790 191.145 110.020 192.135 ;
        RECT 109.355 190.975 110.020 191.145 ;
        RECT 109.355 190.475 109.525 190.975 ;
        RECT 109.695 190.305 110.025 190.805 ;
        RECT 110.195 190.475 110.380 192.595 ;
        RECT 110.635 192.395 110.885 192.855 ;
        RECT 111.055 192.405 111.390 192.575 ;
        RECT 111.585 192.405 112.260 192.575 ;
        RECT 111.055 192.265 111.225 192.405 ;
        RECT 110.550 191.275 110.830 192.225 ;
        RECT 111.000 192.135 111.225 192.265 ;
        RECT 111.000 191.030 111.170 192.135 ;
        RECT 111.395 191.985 111.920 192.205 ;
        RECT 111.340 191.220 111.580 191.815 ;
        RECT 111.750 191.285 111.920 191.985 ;
        RECT 112.090 191.625 112.260 192.405 ;
        RECT 112.580 192.355 112.950 192.855 ;
        RECT 113.130 192.405 113.535 192.575 ;
        RECT 113.705 192.405 114.490 192.575 ;
        RECT 113.130 192.175 113.300 192.405 ;
        RECT 112.470 191.875 113.300 192.175 ;
        RECT 113.685 191.905 114.150 192.235 ;
        RECT 112.470 191.845 112.670 191.875 ;
        RECT 112.790 191.625 112.960 191.695 ;
        RECT 112.090 191.455 112.960 191.625 ;
        RECT 112.450 191.365 112.960 191.455 ;
        RECT 111.000 190.900 111.305 191.030 ;
        RECT 111.750 190.920 112.280 191.285 ;
        RECT 110.620 190.305 110.885 190.765 ;
        RECT 111.055 190.475 111.305 190.900 ;
        RECT 112.450 190.750 112.620 191.365 ;
        RECT 111.515 190.580 112.620 190.750 ;
        RECT 112.790 190.305 112.960 191.105 ;
        RECT 113.130 190.805 113.300 191.875 ;
        RECT 113.470 190.975 113.660 191.695 ;
        RECT 113.830 190.945 114.150 191.905 ;
        RECT 114.320 191.945 114.490 192.405 ;
        RECT 114.765 192.325 114.975 192.855 ;
        RECT 115.235 192.115 115.565 192.640 ;
        RECT 115.735 192.245 115.905 192.855 ;
        RECT 116.075 192.200 116.405 192.635 ;
        RECT 116.715 192.305 116.885 192.595 ;
        RECT 117.055 192.475 117.385 192.855 ;
        RECT 116.075 192.115 116.455 192.200 ;
        RECT 116.715 192.135 117.380 192.305 ;
        RECT 115.365 191.945 115.565 192.115 ;
        RECT 116.230 192.075 116.455 192.115 ;
        RECT 114.320 191.615 115.195 191.945 ;
        RECT 115.365 191.615 116.115 191.945 ;
        RECT 113.130 190.475 113.380 190.805 ;
        RECT 114.320 190.775 114.490 191.615 ;
        RECT 115.365 191.410 115.555 191.615 ;
        RECT 116.285 191.495 116.455 192.075 ;
        RECT 116.240 191.445 116.455 191.495 ;
        RECT 114.660 191.035 115.555 191.410 ;
        RECT 116.065 191.365 116.455 191.445 ;
        RECT 113.605 190.605 114.490 190.775 ;
        RECT 114.670 190.305 114.985 190.805 ;
        RECT 115.215 190.475 115.555 191.035 ;
        RECT 115.725 190.305 115.895 191.315 ;
        RECT 116.065 190.520 116.395 191.365 ;
        RECT 116.630 191.315 116.980 191.965 ;
        RECT 117.150 191.145 117.380 192.135 ;
        RECT 116.715 190.975 117.380 191.145 ;
        RECT 116.715 190.475 116.885 190.975 ;
        RECT 117.055 190.305 117.385 190.805 ;
        RECT 117.555 190.475 117.740 192.595 ;
        RECT 117.995 192.395 118.245 192.855 ;
        RECT 118.415 192.405 118.750 192.575 ;
        RECT 118.945 192.405 119.620 192.575 ;
        RECT 118.415 192.265 118.585 192.405 ;
        RECT 117.910 191.275 118.190 192.225 ;
        RECT 118.360 192.135 118.585 192.265 ;
        RECT 118.360 191.030 118.530 192.135 ;
        RECT 118.755 191.985 119.280 192.205 ;
        RECT 118.700 191.220 118.940 191.815 ;
        RECT 119.110 191.285 119.280 191.985 ;
        RECT 119.450 191.625 119.620 192.405 ;
        RECT 119.940 192.355 120.310 192.855 ;
        RECT 120.490 192.405 120.895 192.575 ;
        RECT 121.065 192.405 121.850 192.575 ;
        RECT 120.490 192.175 120.660 192.405 ;
        RECT 119.830 191.875 120.660 192.175 ;
        RECT 121.045 191.905 121.510 192.235 ;
        RECT 119.830 191.845 120.030 191.875 ;
        RECT 120.150 191.625 120.320 191.695 ;
        RECT 119.450 191.455 120.320 191.625 ;
        RECT 119.810 191.365 120.320 191.455 ;
        RECT 118.360 190.900 118.665 191.030 ;
        RECT 119.110 190.920 119.640 191.285 ;
        RECT 117.980 190.305 118.245 190.765 ;
        RECT 118.415 190.475 118.665 190.900 ;
        RECT 119.810 190.750 119.980 191.365 ;
        RECT 118.875 190.580 119.980 190.750 ;
        RECT 120.150 190.305 120.320 191.105 ;
        RECT 120.490 190.805 120.660 191.875 ;
        RECT 120.830 190.975 121.020 191.695 ;
        RECT 121.190 190.945 121.510 191.905 ;
        RECT 121.680 191.945 121.850 192.405 ;
        RECT 122.125 192.325 122.335 192.855 ;
        RECT 122.595 192.115 122.925 192.640 ;
        RECT 123.095 192.245 123.265 192.855 ;
        RECT 123.435 192.200 123.765 192.635 ;
        RECT 123.435 192.115 123.815 192.200 ;
        RECT 122.725 191.945 122.925 192.115 ;
        RECT 123.590 192.075 123.815 192.115 ;
        RECT 121.680 191.615 122.555 191.945 ;
        RECT 122.725 191.615 123.475 191.945 ;
        RECT 120.490 190.475 120.740 190.805 ;
        RECT 121.680 190.775 121.850 191.615 ;
        RECT 122.725 191.410 122.915 191.615 ;
        RECT 123.645 191.495 123.815 192.075 ;
        RECT 123.985 192.085 125.655 192.855 ;
        RECT 125.825 192.130 126.115 192.855 ;
        RECT 126.755 192.125 127.055 192.855 ;
        RECT 123.985 191.565 124.735 192.085 ;
        RECT 127.235 191.945 127.465 192.565 ;
        RECT 127.665 192.295 127.890 192.675 ;
        RECT 128.060 192.465 128.390 192.855 ;
        RECT 127.665 192.115 127.995 192.295 ;
        RECT 123.600 191.445 123.815 191.495 ;
        RECT 122.020 191.035 122.915 191.410 ;
        RECT 123.425 191.365 123.815 191.445 ;
        RECT 124.905 191.395 125.655 191.915 ;
        RECT 126.760 191.615 127.055 191.945 ;
        RECT 127.235 191.615 127.650 191.945 ;
        RECT 120.965 190.605 121.850 190.775 ;
        RECT 122.030 190.305 122.345 190.805 ;
        RECT 122.575 190.475 122.915 191.035 ;
        RECT 123.085 190.305 123.255 191.315 ;
        RECT 123.425 190.520 123.755 191.365 ;
        RECT 123.985 190.305 125.655 191.395 ;
        RECT 125.825 190.305 126.115 191.470 ;
        RECT 127.820 191.445 127.995 192.115 ;
        RECT 128.165 191.615 128.405 192.265 ;
        RECT 128.585 192.180 128.860 192.525 ;
        RECT 129.050 192.455 129.430 192.855 ;
        RECT 129.600 192.285 129.770 192.635 ;
        RECT 129.940 192.455 130.270 192.855 ;
        RECT 130.445 192.285 130.615 192.635 ;
        RECT 130.815 192.355 131.145 192.855 ;
        RECT 128.585 191.445 128.755 192.180 ;
        RECT 129.030 192.115 130.615 192.285 ;
        RECT 129.030 191.945 129.200 192.115 ;
        RECT 131.340 191.945 131.585 192.635 ;
        RECT 131.755 192.355 132.095 192.855 ;
        RECT 132.265 192.355 132.525 192.685 ;
        RECT 132.695 192.495 133.025 192.855 ;
        RECT 133.280 192.475 134.580 192.685 ;
        RECT 128.925 191.615 129.200 191.945 ;
        RECT 129.370 191.615 129.750 191.945 ;
        RECT 129.030 191.445 129.200 191.615 ;
        RECT 126.755 191.085 127.650 191.415 ;
        RECT 127.820 191.255 128.405 191.445 ;
        RECT 126.755 190.915 127.960 191.085 ;
        RECT 126.755 190.485 127.085 190.915 ;
        RECT 127.265 190.305 127.460 190.745 ;
        RECT 127.630 190.485 127.960 190.915 ;
        RECT 128.130 190.485 128.405 191.255 ;
        RECT 128.585 190.475 128.860 191.445 ;
        RECT 129.030 191.275 129.690 191.445 ;
        RECT 129.920 191.325 130.660 191.945 ;
        RECT 130.930 191.615 131.585 191.945 ;
        RECT 131.755 191.615 132.095 192.185 ;
        RECT 129.520 191.155 129.690 191.275 ;
        RECT 130.830 191.155 131.150 191.445 ;
        RECT 129.070 190.305 129.350 191.105 ;
        RECT 129.520 190.985 131.150 191.155 ;
        RECT 131.345 191.020 131.585 191.615 ;
        RECT 129.520 190.645 131.575 190.815 ;
        RECT 129.520 190.525 131.570 190.645 ;
        RECT 131.755 190.305 132.095 191.380 ;
        RECT 132.265 191.155 132.435 192.355 ;
        RECT 133.280 192.325 133.450 192.475 ;
        RECT 132.695 192.200 133.450 192.325 ;
        RECT 132.605 192.155 133.450 192.200 ;
        RECT 132.605 192.035 132.875 192.155 ;
        RECT 132.605 191.460 132.775 192.035 ;
        RECT 133.005 191.595 133.415 191.900 ;
        RECT 133.705 191.865 133.915 192.265 ;
        RECT 133.585 191.655 133.915 191.865 ;
        RECT 134.160 191.865 134.380 192.265 ;
        RECT 134.855 192.090 135.310 192.855 ;
        RECT 135.485 192.105 136.695 192.855 ;
        RECT 134.160 191.655 134.635 191.865 ;
        RECT 134.825 191.665 135.315 191.865 ;
        RECT 135.485 191.565 136.005 192.105 ;
        RECT 136.865 192.055 137.560 192.685 ;
        RECT 137.765 192.055 138.075 192.855 ;
        RECT 132.605 191.425 132.805 191.460 ;
        RECT 134.135 191.425 135.310 191.485 ;
        RECT 132.605 191.315 135.310 191.425 ;
        RECT 136.175 191.395 136.695 191.935 ;
        RECT 136.885 191.615 137.220 191.865 ;
        RECT 137.390 191.455 137.560 192.055 ;
        RECT 138.305 192.035 138.515 192.855 ;
        RECT 138.685 192.055 139.015 192.685 ;
        RECT 137.730 191.615 138.065 191.885 ;
        RECT 138.685 191.455 138.935 192.055 ;
        RECT 139.185 192.035 139.415 192.855 ;
        RECT 139.625 192.105 140.835 192.855 ;
        RECT 139.105 191.615 139.435 191.865 ;
        RECT 139.625 191.565 140.145 192.105 ;
        RECT 141.005 192.035 141.265 192.855 ;
        RECT 141.435 192.035 141.765 192.455 ;
        RECT 141.945 192.370 142.735 192.635 ;
        RECT 141.515 191.945 141.765 192.035 ;
        RECT 132.665 191.255 134.465 191.315 ;
        RECT 134.135 191.225 134.465 191.255 ;
        RECT 132.265 190.475 132.525 191.155 ;
        RECT 132.695 190.305 132.945 191.085 ;
        RECT 133.195 191.055 134.030 191.065 ;
        RECT 134.620 191.055 134.805 191.145 ;
        RECT 133.195 190.855 134.805 191.055 ;
        RECT 133.195 190.475 133.445 190.855 ;
        RECT 134.575 190.815 134.805 190.855 ;
        RECT 135.055 190.695 135.310 191.315 ;
        RECT 133.615 190.305 133.970 190.685 ;
        RECT 134.975 190.475 135.310 190.695 ;
        RECT 135.485 190.305 136.695 191.395 ;
        RECT 136.865 190.305 137.125 191.445 ;
        RECT 137.295 190.475 137.625 191.455 ;
        RECT 137.795 190.305 138.075 191.445 ;
        RECT 138.305 190.305 138.515 191.445 ;
        RECT 138.685 190.475 139.015 191.455 ;
        RECT 139.185 190.305 139.415 191.445 ;
        RECT 140.315 191.395 140.835 191.935 ;
        RECT 139.625 190.305 140.835 191.395 ;
        RECT 141.005 190.985 141.345 191.865 ;
        RECT 141.515 191.695 142.310 191.945 ;
        RECT 141.005 190.305 141.265 190.815 ;
        RECT 141.515 190.475 141.685 191.695 ;
        RECT 142.480 191.515 142.735 192.370 ;
        RECT 142.905 192.215 143.105 192.635 ;
        RECT 143.295 192.395 143.625 192.855 ;
        RECT 142.905 191.695 143.315 192.215 ;
        RECT 143.795 192.205 144.055 192.685 ;
        RECT 143.485 191.515 143.715 191.945 ;
        RECT 141.925 191.345 143.715 191.515 ;
        RECT 141.925 190.980 142.175 191.345 ;
        RECT 142.345 190.985 142.675 191.175 ;
        RECT 142.895 191.050 143.610 191.345 ;
        RECT 143.885 191.175 144.055 192.205 ;
        RECT 144.275 192.200 144.605 192.635 ;
        RECT 144.775 192.245 144.945 192.855 ;
        RECT 144.225 192.115 144.605 192.200 ;
        RECT 145.115 192.115 145.445 192.640 ;
        RECT 145.705 192.325 145.915 192.855 ;
        RECT 146.190 192.405 146.975 192.575 ;
        RECT 147.145 192.405 147.550 192.575 ;
        RECT 144.225 192.075 144.450 192.115 ;
        RECT 144.225 191.495 144.395 192.075 ;
        RECT 145.115 191.945 145.315 192.115 ;
        RECT 146.190 191.945 146.360 192.405 ;
        RECT 144.565 191.615 145.315 191.945 ;
        RECT 145.485 191.615 146.360 191.945 ;
        RECT 144.225 191.445 144.440 191.495 ;
        RECT 144.225 191.365 144.615 191.445 ;
        RECT 142.345 190.810 142.540 190.985 ;
        RECT 141.925 190.305 142.540 190.810 ;
        RECT 142.710 190.475 143.185 190.815 ;
        RECT 143.355 190.305 143.570 190.850 ;
        RECT 143.780 190.475 144.055 191.175 ;
        RECT 144.285 190.520 144.615 191.365 ;
        RECT 145.125 191.410 145.315 191.615 ;
        RECT 144.785 190.305 144.955 191.315 ;
        RECT 145.125 191.035 146.020 191.410 ;
        RECT 145.125 190.475 145.465 191.035 ;
        RECT 145.695 190.305 146.010 190.805 ;
        RECT 146.190 190.775 146.360 191.615 ;
        RECT 146.530 191.905 146.995 192.235 ;
        RECT 147.380 192.175 147.550 192.405 ;
        RECT 147.730 192.355 148.100 192.855 ;
        RECT 148.420 192.405 149.095 192.575 ;
        RECT 149.290 192.405 149.625 192.575 ;
        RECT 146.530 190.945 146.850 191.905 ;
        RECT 147.380 191.875 148.210 192.175 ;
        RECT 147.020 190.975 147.210 191.695 ;
        RECT 147.380 190.805 147.550 191.875 ;
        RECT 148.010 191.845 148.210 191.875 ;
        RECT 147.720 191.625 147.890 191.695 ;
        RECT 148.420 191.625 148.590 192.405 ;
        RECT 149.455 192.265 149.625 192.405 ;
        RECT 149.795 192.395 150.045 192.855 ;
        RECT 147.720 191.455 148.590 191.625 ;
        RECT 148.760 191.985 149.285 192.205 ;
        RECT 149.455 192.135 149.680 192.265 ;
        RECT 147.720 191.365 148.230 191.455 ;
        RECT 146.190 190.605 147.075 190.775 ;
        RECT 147.300 190.475 147.550 190.805 ;
        RECT 147.720 190.305 147.890 191.105 ;
        RECT 148.060 190.750 148.230 191.365 ;
        RECT 148.760 191.285 148.930 191.985 ;
        RECT 148.400 190.920 148.930 191.285 ;
        RECT 149.100 191.220 149.340 191.815 ;
        RECT 149.510 191.030 149.680 192.135 ;
        RECT 149.850 191.275 150.130 192.225 ;
        RECT 149.375 190.900 149.680 191.030 ;
        RECT 148.060 190.580 149.165 190.750 ;
        RECT 149.375 190.475 149.625 190.900 ;
        RECT 149.795 190.305 150.060 190.765 ;
        RECT 150.300 190.475 150.485 192.595 ;
        RECT 150.655 192.475 150.985 192.855 ;
        RECT 151.155 192.305 151.325 192.595 ;
        RECT 150.660 192.135 151.325 192.305 ;
        RECT 150.660 191.145 150.890 192.135 ;
        RECT 151.585 192.130 151.875 192.855 ;
        RECT 152.045 192.085 155.555 192.855 ;
        RECT 155.725 192.105 156.935 192.855 ;
        RECT 151.060 191.315 151.410 191.965 ;
        RECT 152.045 191.565 153.695 192.085 ;
        RECT 150.660 190.975 151.325 191.145 ;
        RECT 150.655 190.305 150.985 190.805 ;
        RECT 151.155 190.475 151.325 190.975 ;
        RECT 151.585 190.305 151.875 191.470 ;
        RECT 153.865 191.395 155.555 191.915 ;
        RECT 152.045 190.305 155.555 191.395 ;
        RECT 155.725 191.395 156.245 191.935 ;
        RECT 156.415 191.565 156.935 192.105 ;
        RECT 155.725 190.305 156.935 191.395 ;
        RECT 22.700 190.135 157.020 190.305 ;
        RECT 22.785 189.045 23.995 190.135 ;
        RECT 24.255 189.465 24.425 189.965 ;
        RECT 24.595 189.635 24.925 190.135 ;
        RECT 24.255 189.295 24.920 189.465 ;
        RECT 22.785 188.335 23.305 188.875 ;
        RECT 23.475 188.505 23.995 189.045 ;
        RECT 24.170 188.475 24.520 189.125 ;
        RECT 22.785 187.585 23.995 188.335 ;
        RECT 24.690 188.305 24.920 189.295 ;
        RECT 24.255 188.135 24.920 188.305 ;
        RECT 24.255 187.845 24.425 188.135 ;
        RECT 24.595 187.585 24.925 187.965 ;
        RECT 25.095 187.845 25.280 189.965 ;
        RECT 25.520 189.675 25.785 190.135 ;
        RECT 25.955 189.540 26.205 189.965 ;
        RECT 26.415 189.690 27.520 189.860 ;
        RECT 25.900 189.410 26.205 189.540 ;
        RECT 25.450 188.215 25.730 189.165 ;
        RECT 25.900 188.305 26.070 189.410 ;
        RECT 26.240 188.625 26.480 189.220 ;
        RECT 26.650 189.155 27.180 189.520 ;
        RECT 26.650 188.455 26.820 189.155 ;
        RECT 27.350 189.075 27.520 189.690 ;
        RECT 27.690 189.335 27.860 190.135 ;
        RECT 28.030 189.635 28.280 189.965 ;
        RECT 28.505 189.665 29.390 189.835 ;
        RECT 27.350 188.985 27.860 189.075 ;
        RECT 25.900 188.175 26.125 188.305 ;
        RECT 26.295 188.235 26.820 188.455 ;
        RECT 26.990 188.815 27.860 188.985 ;
        RECT 25.535 187.585 25.785 188.045 ;
        RECT 25.955 188.035 26.125 188.175 ;
        RECT 26.990 188.035 27.160 188.815 ;
        RECT 27.690 188.745 27.860 188.815 ;
        RECT 27.370 188.565 27.570 188.595 ;
        RECT 28.030 188.565 28.200 189.635 ;
        RECT 28.370 188.745 28.560 189.465 ;
        RECT 27.370 188.265 28.200 188.565 ;
        RECT 28.730 188.535 29.050 189.495 ;
        RECT 25.955 187.865 26.290 188.035 ;
        RECT 26.485 187.865 27.160 188.035 ;
        RECT 27.480 187.585 27.850 188.085 ;
        RECT 28.030 188.035 28.200 188.265 ;
        RECT 28.585 188.205 29.050 188.535 ;
        RECT 29.220 188.825 29.390 189.665 ;
        RECT 29.570 189.635 29.885 190.135 ;
        RECT 30.115 189.405 30.455 189.965 ;
        RECT 29.560 189.030 30.455 189.405 ;
        RECT 30.625 189.125 30.795 190.135 ;
        RECT 30.265 188.825 30.455 189.030 ;
        RECT 30.965 189.075 31.295 189.920 ;
        RECT 31.525 189.265 31.800 189.965 ;
        RECT 32.010 189.590 32.225 190.135 ;
        RECT 32.395 189.625 32.870 189.965 ;
        RECT 33.040 189.630 33.655 190.135 ;
        RECT 33.040 189.455 33.235 189.630 ;
        RECT 30.965 188.995 31.355 189.075 ;
        RECT 31.140 188.945 31.355 188.995 ;
        RECT 29.220 188.495 30.095 188.825 ;
        RECT 30.265 188.495 31.015 188.825 ;
        RECT 29.220 188.035 29.390 188.495 ;
        RECT 30.265 188.325 30.465 188.495 ;
        RECT 31.185 188.365 31.355 188.945 ;
        RECT 31.130 188.325 31.355 188.365 ;
        RECT 28.030 187.865 28.435 188.035 ;
        RECT 28.605 187.865 29.390 188.035 ;
        RECT 29.665 187.585 29.875 188.115 ;
        RECT 30.135 187.800 30.465 188.325 ;
        RECT 30.975 188.240 31.355 188.325 ;
        RECT 30.635 187.585 30.805 188.195 ;
        RECT 30.975 187.805 31.305 188.240 ;
        RECT 31.525 188.235 31.695 189.265 ;
        RECT 31.970 189.095 32.685 189.390 ;
        RECT 32.905 189.265 33.235 189.455 ;
        RECT 33.405 189.095 33.655 189.460 ;
        RECT 31.865 188.925 33.655 189.095 ;
        RECT 31.865 188.495 32.095 188.925 ;
        RECT 31.525 187.755 31.785 188.235 ;
        RECT 32.265 188.225 32.675 188.745 ;
        RECT 31.955 187.585 32.285 188.045 ;
        RECT 32.475 187.805 32.675 188.225 ;
        RECT 32.845 188.070 33.100 188.925 ;
        RECT 33.895 188.745 34.065 189.965 ;
        RECT 34.315 189.625 34.575 190.135 ;
        RECT 33.270 188.495 34.065 188.745 ;
        RECT 34.235 188.575 34.575 189.455 ;
        RECT 35.665 188.970 35.955 190.135 ;
        RECT 36.125 189.045 37.795 190.135 ;
        RECT 37.965 189.625 38.225 190.135 ;
        RECT 33.815 188.405 34.065 188.495 ;
        RECT 32.845 187.805 33.635 188.070 ;
        RECT 33.815 187.985 34.145 188.405 ;
        RECT 34.315 187.585 34.575 188.405 ;
        RECT 36.125 188.355 36.875 188.875 ;
        RECT 37.045 188.525 37.795 189.045 ;
        RECT 37.965 188.575 38.305 189.455 ;
        RECT 38.475 188.745 38.645 189.965 ;
        RECT 38.885 189.630 39.500 190.135 ;
        RECT 38.885 189.095 39.135 189.460 ;
        RECT 39.305 189.455 39.500 189.630 ;
        RECT 39.670 189.625 40.145 189.965 ;
        RECT 40.315 189.590 40.530 190.135 ;
        RECT 39.305 189.265 39.635 189.455 ;
        RECT 39.855 189.095 40.570 189.390 ;
        RECT 40.740 189.265 41.015 189.965 ;
        RECT 38.885 188.925 40.675 189.095 ;
        RECT 38.475 188.495 39.270 188.745 ;
        RECT 38.475 188.405 38.725 188.495 ;
        RECT 35.665 187.585 35.955 188.310 ;
        RECT 36.125 187.585 37.795 188.355 ;
        RECT 37.965 187.585 38.225 188.405 ;
        RECT 38.395 187.985 38.725 188.405 ;
        RECT 39.440 188.070 39.695 188.925 ;
        RECT 38.905 187.805 39.695 188.070 ;
        RECT 39.865 188.225 40.275 188.745 ;
        RECT 40.445 188.495 40.675 188.925 ;
        RECT 40.845 188.235 41.015 189.265 ;
        RECT 41.185 189.045 42.395 190.135 ;
        RECT 39.865 187.805 40.065 188.225 ;
        RECT 40.255 187.585 40.585 188.045 ;
        RECT 40.755 187.755 41.015 188.235 ;
        RECT 41.185 188.335 41.705 188.875 ;
        RECT 41.875 188.505 42.395 189.045 ;
        RECT 42.575 189.075 42.905 189.925 ;
        RECT 41.185 187.585 42.395 188.335 ;
        RECT 42.575 188.310 42.765 189.075 ;
        RECT 43.075 188.995 43.325 190.135 ;
        RECT 43.515 189.495 43.765 189.915 ;
        RECT 43.995 189.665 44.325 190.135 ;
        RECT 44.555 189.495 44.805 189.915 ;
        RECT 43.515 189.325 44.805 189.495 ;
        RECT 44.985 189.495 45.315 189.925 ;
        RECT 44.985 189.325 45.440 189.495 ;
        RECT 43.505 188.825 43.720 189.155 ;
        RECT 42.935 188.495 43.245 188.825 ;
        RECT 43.415 188.495 43.720 188.825 ;
        RECT 43.895 188.495 44.180 189.155 ;
        RECT 44.375 188.495 44.640 189.155 ;
        RECT 44.855 188.495 45.100 189.155 ;
        RECT 43.075 188.325 43.245 188.495 ;
        RECT 45.270 188.325 45.440 189.325 ;
        RECT 45.785 189.045 47.455 190.135 ;
        RECT 42.575 187.800 42.905 188.310 ;
        RECT 43.075 188.155 45.440 188.325 ;
        RECT 45.785 188.355 46.535 188.875 ;
        RECT 46.705 188.525 47.455 189.045 ;
        RECT 48.085 188.995 48.355 189.965 ;
        RECT 48.565 189.335 48.845 190.135 ;
        RECT 49.025 189.585 50.220 189.915 ;
        RECT 49.350 189.165 49.770 189.415 ;
        RECT 48.525 188.995 49.770 189.165 ;
        RECT 43.075 187.585 43.405 187.985 ;
        RECT 44.455 187.815 44.785 188.155 ;
        RECT 44.955 187.585 45.285 187.985 ;
        RECT 45.785 187.585 47.455 188.355 ;
        RECT 48.085 188.260 48.255 188.995 ;
        RECT 48.525 188.825 48.695 188.995 ;
        RECT 49.995 188.825 50.165 189.385 ;
        RECT 50.415 188.995 50.670 190.135 ;
        RECT 50.850 189.745 51.185 189.965 ;
        RECT 52.190 189.755 52.545 190.135 ;
        RECT 50.850 189.125 51.105 189.745 ;
        RECT 51.355 189.585 51.585 189.625 ;
        RECT 52.715 189.585 52.965 189.965 ;
        RECT 51.355 189.385 52.965 189.585 ;
        RECT 51.355 189.295 51.540 189.385 ;
        RECT 52.130 189.375 52.965 189.385 ;
        RECT 53.215 189.355 53.465 190.135 ;
        RECT 53.635 189.285 53.895 189.965 ;
        RECT 54.180 189.505 54.465 189.965 ;
        RECT 54.635 189.675 54.905 190.135 ;
        RECT 54.180 189.285 55.135 189.505 ;
        RECT 51.695 189.185 52.025 189.215 ;
        RECT 51.695 189.125 53.495 189.185 ;
        RECT 50.850 189.015 53.555 189.125 ;
        RECT 50.850 188.955 52.025 189.015 ;
        RECT 53.355 188.980 53.555 189.015 ;
        RECT 48.465 188.495 48.695 188.825 ;
        RECT 49.425 188.495 50.165 188.825 ;
        RECT 50.335 188.575 50.670 188.825 ;
        RECT 50.845 188.575 51.335 188.775 ;
        RECT 51.525 188.575 52.000 188.785 ;
        RECT 48.525 188.325 48.695 188.495 ;
        RECT 49.915 188.405 50.165 188.495 ;
        RECT 48.085 187.915 48.355 188.260 ;
        RECT 48.525 188.155 49.265 188.325 ;
        RECT 49.915 188.235 50.650 188.405 ;
        RECT 48.545 187.585 48.925 187.985 ;
        RECT 49.095 187.805 49.265 188.155 ;
        RECT 49.435 187.585 50.170 188.065 ;
        RECT 50.340 187.765 50.650 188.235 ;
        RECT 50.850 187.585 51.305 188.350 ;
        RECT 51.780 188.175 52.000 188.575 ;
        RECT 52.245 188.575 52.575 188.785 ;
        RECT 52.245 188.175 52.455 188.575 ;
        RECT 52.745 188.540 53.155 188.845 ;
        RECT 53.385 188.405 53.555 188.980 ;
        RECT 53.285 188.285 53.555 188.405 ;
        RECT 52.710 188.240 53.555 188.285 ;
        RECT 52.710 188.115 53.465 188.240 ;
        RECT 52.710 187.965 52.880 188.115 ;
        RECT 53.725 188.095 53.895 189.285 ;
        RECT 54.065 188.555 54.755 189.115 ;
        RECT 54.925 188.385 55.135 189.285 ;
        RECT 53.665 188.085 53.895 188.095 ;
        RECT 51.580 187.755 52.880 187.965 ;
        RECT 53.135 187.585 53.465 187.945 ;
        RECT 53.635 187.755 53.895 188.085 ;
        RECT 54.180 188.215 55.135 188.385 ;
        RECT 55.305 189.115 55.705 189.965 ;
        RECT 55.895 189.505 56.175 189.965 ;
        RECT 56.695 189.675 57.020 190.135 ;
        RECT 55.895 189.285 57.020 189.505 ;
        RECT 55.305 188.555 56.400 189.115 ;
        RECT 56.570 188.825 57.020 189.285 ;
        RECT 57.190 188.995 57.575 189.965 ;
        RECT 54.180 187.755 54.465 188.215 ;
        RECT 54.635 187.585 54.905 188.045 ;
        RECT 55.305 187.755 55.705 188.555 ;
        RECT 56.570 188.495 57.125 188.825 ;
        RECT 56.570 188.385 57.020 188.495 ;
        RECT 55.895 188.215 57.020 188.385 ;
        RECT 57.295 188.325 57.575 188.995 ;
        RECT 55.895 187.755 56.175 188.215 ;
        RECT 56.695 187.585 57.020 188.045 ;
        RECT 57.190 187.755 57.575 188.325 ;
        RECT 57.745 188.995 58.130 189.965 ;
        RECT 58.300 189.675 58.625 190.135 ;
        RECT 59.145 189.505 59.425 189.965 ;
        RECT 58.300 189.285 59.425 189.505 ;
        RECT 57.745 188.325 58.025 188.995 ;
        RECT 58.300 188.825 58.750 189.285 ;
        RECT 59.615 189.115 60.015 189.965 ;
        RECT 60.415 189.675 60.685 190.135 ;
        RECT 60.855 189.505 61.140 189.965 ;
        RECT 58.195 188.495 58.750 188.825 ;
        RECT 58.920 188.555 60.015 189.115 ;
        RECT 58.300 188.385 58.750 188.495 ;
        RECT 57.745 187.755 58.130 188.325 ;
        RECT 58.300 188.215 59.425 188.385 ;
        RECT 58.300 187.585 58.625 188.045 ;
        RECT 59.145 187.755 59.425 188.215 ;
        RECT 59.615 187.755 60.015 188.555 ;
        RECT 60.185 189.285 61.140 189.505 ;
        RECT 60.185 188.385 60.395 189.285 ;
        RECT 60.565 188.555 61.255 189.115 ;
        RECT 61.425 188.970 61.715 190.135 ;
        RECT 62.350 188.995 62.605 190.135 ;
        RECT 62.800 189.585 63.995 189.915 ;
        RECT 62.855 188.825 63.025 189.385 ;
        RECT 63.250 189.165 63.670 189.415 ;
        RECT 64.175 189.335 64.455 190.135 ;
        RECT 63.250 188.995 64.495 189.165 ;
        RECT 64.665 188.995 64.935 189.965 ;
        RECT 64.325 188.825 64.495 188.995 ;
        RECT 62.350 188.575 62.685 188.825 ;
        RECT 62.855 188.495 63.595 188.825 ;
        RECT 64.325 188.495 64.555 188.825 ;
        RECT 62.855 188.405 63.105 188.495 ;
        RECT 60.185 188.215 61.140 188.385 ;
        RECT 60.415 187.585 60.685 188.045 ;
        RECT 60.855 187.755 61.140 188.215 ;
        RECT 61.425 187.585 61.715 188.310 ;
        RECT 62.370 188.235 63.105 188.405 ;
        RECT 64.325 188.325 64.495 188.495 ;
        RECT 62.370 187.765 62.680 188.235 ;
        RECT 63.755 188.155 64.495 188.325 ;
        RECT 64.765 188.260 64.935 188.995 ;
        RECT 65.195 189.125 65.365 189.965 ;
        RECT 65.535 189.795 66.705 189.965 ;
        RECT 65.535 189.295 65.865 189.795 ;
        RECT 66.375 189.755 66.705 189.795 ;
        RECT 66.895 189.715 67.250 190.135 ;
        RECT 66.035 189.535 66.265 189.625 ;
        RECT 67.420 189.535 67.670 189.965 ;
        RECT 66.035 189.295 67.670 189.535 ;
        RECT 67.840 189.375 68.170 190.135 ;
        RECT 68.340 189.295 68.595 189.965 ;
        RECT 65.195 188.955 68.255 189.125 ;
        RECT 65.110 188.575 65.460 188.785 ;
        RECT 65.630 188.575 66.075 188.775 ;
        RECT 66.245 188.575 66.720 188.775 ;
        RECT 62.850 187.585 63.585 188.065 ;
        RECT 63.755 187.805 63.925 188.155 ;
        RECT 64.095 187.585 64.475 187.985 ;
        RECT 64.665 187.915 64.935 188.260 ;
        RECT 65.195 188.235 66.260 188.405 ;
        RECT 65.195 187.755 65.365 188.235 ;
        RECT 65.535 187.585 65.865 188.065 ;
        RECT 66.090 188.005 66.260 188.235 ;
        RECT 66.440 188.175 66.720 188.575 ;
        RECT 66.990 188.575 67.320 188.775 ;
        RECT 67.490 188.605 67.865 188.775 ;
        RECT 67.490 188.575 67.855 188.605 ;
        RECT 66.990 188.175 67.275 188.575 ;
        RECT 68.085 188.405 68.255 188.955 ;
        RECT 67.455 188.235 68.255 188.405 ;
        RECT 67.455 188.005 67.625 188.235 ;
        RECT 68.425 188.165 68.595 189.295 ;
        RECT 68.805 189.245 69.065 189.955 ;
        RECT 69.235 189.425 69.565 190.135 ;
        RECT 69.735 189.245 69.965 189.955 ;
        RECT 68.805 189.005 69.965 189.245 ;
        RECT 70.145 189.225 70.415 189.955 ;
        RECT 70.595 189.405 70.935 190.135 ;
        RECT 70.145 189.005 70.915 189.225 ;
        RECT 68.795 188.495 69.095 188.825 ;
        RECT 69.275 188.515 69.800 188.825 ;
        RECT 69.980 188.515 70.445 188.825 ;
        RECT 68.410 188.095 68.595 188.165 ;
        RECT 68.385 188.085 68.595 188.095 ;
        RECT 66.090 187.755 67.625 188.005 ;
        RECT 67.795 187.585 68.125 188.065 ;
        RECT 68.340 187.755 68.595 188.085 ;
        RECT 68.805 187.585 69.095 188.315 ;
        RECT 69.275 187.875 69.505 188.515 ;
        RECT 70.625 188.335 70.915 189.005 ;
        RECT 69.685 188.135 70.915 188.335 ;
        RECT 69.685 187.765 69.995 188.135 ;
        RECT 70.175 187.585 70.845 187.955 ;
        RECT 71.105 187.765 71.365 189.955 ;
        RECT 71.545 189.285 71.805 189.965 ;
        RECT 71.975 189.355 72.225 190.135 ;
        RECT 72.475 189.585 72.725 189.965 ;
        RECT 72.895 189.755 73.250 190.135 ;
        RECT 74.255 189.745 74.590 189.965 ;
        RECT 73.855 189.585 74.085 189.625 ;
        RECT 72.475 189.385 74.085 189.585 ;
        RECT 72.475 189.375 73.310 189.385 ;
        RECT 73.900 189.295 74.085 189.385 ;
        RECT 71.545 188.085 71.715 189.285 ;
        RECT 73.415 189.185 73.745 189.215 ;
        RECT 71.945 189.125 73.745 189.185 ;
        RECT 74.335 189.125 74.590 189.745 ;
        RECT 71.885 189.015 74.590 189.125 ;
        RECT 74.765 189.045 75.975 190.135 ;
        RECT 71.885 188.980 72.085 189.015 ;
        RECT 71.885 188.405 72.055 188.980 ;
        RECT 73.415 188.955 74.590 189.015 ;
        RECT 72.285 188.540 72.695 188.845 ;
        RECT 72.865 188.575 73.195 188.785 ;
        RECT 71.885 188.285 72.155 188.405 ;
        RECT 71.885 188.240 72.730 188.285 ;
        RECT 71.975 188.115 72.730 188.240 ;
        RECT 72.985 188.175 73.195 188.575 ;
        RECT 73.440 188.575 73.915 188.785 ;
        RECT 74.105 188.575 74.595 188.775 ;
        RECT 73.440 188.175 73.660 188.575 ;
        RECT 71.545 187.755 71.805 188.085 ;
        RECT 72.560 187.965 72.730 188.115 ;
        RECT 71.975 187.585 72.305 187.945 ;
        RECT 72.560 187.755 73.860 187.965 ;
        RECT 74.135 187.585 74.590 188.350 ;
        RECT 74.765 188.335 75.285 188.875 ;
        RECT 75.455 188.505 75.975 189.045 ;
        RECT 74.765 187.585 75.975 188.335 ;
        RECT 76.145 187.865 76.425 189.965 ;
        RECT 76.615 189.375 77.400 190.135 ;
        RECT 77.795 189.305 78.180 189.965 ;
        RECT 77.795 189.205 78.205 189.305 ;
        RECT 76.595 188.995 78.205 189.205 ;
        RECT 78.505 189.115 78.705 189.905 ;
        RECT 76.595 188.395 76.870 188.995 ;
        RECT 78.375 188.945 78.705 189.115 ;
        RECT 78.875 188.955 79.195 190.135 ;
        RECT 79.830 189.745 80.165 189.965 ;
        RECT 81.170 189.755 81.525 190.135 ;
        RECT 79.830 189.125 80.085 189.745 ;
        RECT 80.335 189.585 80.565 189.625 ;
        RECT 81.695 189.585 81.945 189.965 ;
        RECT 80.335 189.385 81.945 189.585 ;
        RECT 80.335 189.295 80.520 189.385 ;
        RECT 81.110 189.375 81.945 189.385 ;
        RECT 82.195 189.355 82.445 190.135 ;
        RECT 82.615 189.285 82.875 189.965 ;
        RECT 80.675 189.185 81.005 189.215 ;
        RECT 80.675 189.125 82.475 189.185 ;
        RECT 79.830 189.015 82.535 189.125 ;
        RECT 79.830 188.955 81.005 189.015 ;
        RECT 82.335 188.980 82.535 189.015 ;
        RECT 78.375 188.825 78.555 188.945 ;
        RECT 77.040 188.575 77.395 188.825 ;
        RECT 77.590 188.775 78.055 188.825 ;
        RECT 77.585 188.605 78.055 188.775 ;
        RECT 77.590 188.575 78.055 188.605 ;
        RECT 78.225 188.575 78.555 188.825 ;
        RECT 78.730 188.575 79.195 188.775 ;
        RECT 79.825 188.575 80.315 188.775 ;
        RECT 80.505 188.575 80.980 188.785 ;
        RECT 76.595 188.215 77.845 188.395 ;
        RECT 77.480 188.145 77.845 188.215 ;
        RECT 78.015 188.195 79.195 188.365 ;
        RECT 76.655 187.585 76.825 188.045 ;
        RECT 78.015 187.975 78.345 188.195 ;
        RECT 77.095 187.795 78.345 187.975 ;
        RECT 78.515 187.585 78.685 188.025 ;
        RECT 78.855 187.780 79.195 188.195 ;
        RECT 79.830 187.585 80.285 188.350 ;
        RECT 80.760 188.175 80.980 188.575 ;
        RECT 81.225 188.575 81.555 188.785 ;
        RECT 81.225 188.175 81.435 188.575 ;
        RECT 81.725 188.540 82.135 188.845 ;
        RECT 82.365 188.405 82.535 188.980 ;
        RECT 82.265 188.285 82.535 188.405 ;
        RECT 81.690 188.240 82.535 188.285 ;
        RECT 81.690 188.115 82.445 188.240 ;
        RECT 81.690 187.965 81.860 188.115 ;
        RECT 82.705 188.095 82.875 189.285 ;
        RECT 82.645 188.085 82.875 188.095 ;
        RECT 80.560 187.755 81.860 187.965 ;
        RECT 82.115 187.585 82.445 187.945 ;
        RECT 82.615 187.755 82.875 188.085 ;
        RECT 83.505 187.865 83.785 189.965 ;
        RECT 83.975 189.375 84.760 190.135 ;
        RECT 85.155 189.305 85.540 189.965 ;
        RECT 85.155 189.205 85.565 189.305 ;
        RECT 83.955 188.995 85.565 189.205 ;
        RECT 85.865 189.115 86.065 189.905 ;
        RECT 83.955 188.395 84.230 188.995 ;
        RECT 85.735 188.945 86.065 189.115 ;
        RECT 86.235 188.955 86.555 190.135 ;
        RECT 87.185 188.970 87.475 190.135 ;
        RECT 87.645 189.285 87.905 189.965 ;
        RECT 88.075 189.355 88.325 190.135 ;
        RECT 88.575 189.585 88.825 189.965 ;
        RECT 88.995 189.755 89.350 190.135 ;
        RECT 90.355 189.745 90.690 189.965 ;
        RECT 89.955 189.585 90.185 189.625 ;
        RECT 88.575 189.385 90.185 189.585 ;
        RECT 88.575 189.375 89.410 189.385 ;
        RECT 90.000 189.295 90.185 189.385 ;
        RECT 85.735 188.825 85.915 188.945 ;
        RECT 84.400 188.575 84.755 188.825 ;
        RECT 84.950 188.775 85.415 188.825 ;
        RECT 84.945 188.605 85.415 188.775 ;
        RECT 84.950 188.575 85.415 188.605 ;
        RECT 85.585 188.575 85.915 188.825 ;
        RECT 86.090 188.575 86.555 188.775 ;
        RECT 83.955 188.215 85.205 188.395 ;
        RECT 84.840 188.145 85.205 188.215 ;
        RECT 85.375 188.195 86.555 188.365 ;
        RECT 84.015 187.585 84.185 188.045 ;
        RECT 85.375 187.975 85.705 188.195 ;
        RECT 84.455 187.795 85.705 187.975 ;
        RECT 85.875 187.585 86.045 188.025 ;
        RECT 86.215 187.780 86.555 188.195 ;
        RECT 87.185 187.585 87.475 188.310 ;
        RECT 87.645 188.095 87.815 189.285 ;
        RECT 89.515 189.185 89.845 189.215 ;
        RECT 88.045 189.125 89.845 189.185 ;
        RECT 90.435 189.125 90.690 189.745 ;
        RECT 87.985 189.015 90.690 189.125 ;
        RECT 91.335 189.525 91.665 189.955 ;
        RECT 91.845 189.695 92.040 190.135 ;
        RECT 92.210 189.525 92.540 189.955 ;
        RECT 91.335 189.355 92.540 189.525 ;
        RECT 91.335 189.025 92.230 189.355 ;
        RECT 92.710 189.185 92.985 189.955 ;
        RECT 87.985 188.980 88.185 189.015 ;
        RECT 87.985 188.405 88.155 188.980 ;
        RECT 89.515 188.955 90.690 189.015 ;
        RECT 92.400 188.995 92.985 189.185 ;
        RECT 88.385 188.540 88.795 188.845 ;
        RECT 88.965 188.575 89.295 188.785 ;
        RECT 87.985 188.285 88.255 188.405 ;
        RECT 87.985 188.240 88.830 188.285 ;
        RECT 88.075 188.115 88.830 188.240 ;
        RECT 89.085 188.175 89.295 188.575 ;
        RECT 89.540 188.575 90.015 188.785 ;
        RECT 90.205 188.575 90.695 188.775 ;
        RECT 89.540 188.175 89.760 188.575 ;
        RECT 91.340 188.495 91.635 188.825 ;
        RECT 91.815 188.495 92.230 188.825 ;
        RECT 87.645 188.085 87.875 188.095 ;
        RECT 87.645 187.755 87.905 188.085 ;
        RECT 88.660 187.965 88.830 188.115 ;
        RECT 88.075 187.585 88.405 187.945 ;
        RECT 88.660 187.755 89.960 187.965 ;
        RECT 90.235 187.585 90.690 188.350 ;
        RECT 91.335 187.585 91.635 188.315 ;
        RECT 91.815 187.875 92.045 188.495 ;
        RECT 92.400 188.325 92.575 188.995 ;
        RECT 92.245 188.145 92.575 188.325 ;
        RECT 92.745 188.175 92.985 188.825 ;
        RECT 92.245 187.765 92.470 188.145 ;
        RECT 92.640 187.585 92.970 187.975 ;
        RECT 93.165 187.865 93.445 189.965 ;
        RECT 93.635 189.375 94.420 190.135 ;
        RECT 94.815 189.305 95.200 189.965 ;
        RECT 94.815 189.205 95.225 189.305 ;
        RECT 93.615 188.995 95.225 189.205 ;
        RECT 95.525 189.115 95.725 189.905 ;
        RECT 93.615 188.395 93.890 188.995 ;
        RECT 95.395 188.945 95.725 189.115 ;
        RECT 95.895 188.955 96.215 190.135 ;
        RECT 96.850 189.185 97.115 189.955 ;
        RECT 97.285 189.415 97.615 190.135 ;
        RECT 97.805 189.595 98.065 189.955 ;
        RECT 98.235 189.765 98.565 190.135 ;
        RECT 98.735 189.595 98.995 189.955 ;
        RECT 97.805 189.365 98.995 189.595 ;
        RECT 99.565 189.185 99.855 189.955 ;
        RECT 100.065 189.700 105.410 190.135 ;
        RECT 106.050 189.745 106.385 189.965 ;
        RECT 107.390 189.755 107.745 190.135 ;
        RECT 95.395 188.825 95.575 188.945 ;
        RECT 94.060 188.575 94.415 188.825 ;
        RECT 94.610 188.775 95.075 188.825 ;
        RECT 94.605 188.605 95.075 188.775 ;
        RECT 94.610 188.575 95.075 188.605 ;
        RECT 95.245 188.575 95.575 188.825 ;
        RECT 95.750 188.575 96.215 188.775 ;
        RECT 93.615 188.215 94.865 188.395 ;
        RECT 94.500 188.145 94.865 188.215 ;
        RECT 95.035 188.195 96.215 188.365 ;
        RECT 93.675 187.585 93.845 188.045 ;
        RECT 95.035 187.975 95.365 188.195 ;
        RECT 94.115 187.795 95.365 187.975 ;
        RECT 95.535 187.585 95.705 188.025 ;
        RECT 95.875 187.780 96.215 188.195 ;
        RECT 96.850 187.765 97.185 189.185 ;
        RECT 97.360 189.005 99.855 189.185 ;
        RECT 97.360 188.315 97.585 189.005 ;
        RECT 97.785 188.495 98.065 188.825 ;
        RECT 98.245 188.495 98.820 188.825 ;
        RECT 99.000 188.495 99.435 188.825 ;
        RECT 99.615 188.495 99.885 188.825 ;
        RECT 97.360 188.125 99.845 188.315 ;
        RECT 101.650 188.130 101.990 188.960 ;
        RECT 103.470 188.450 103.820 189.700 ;
        RECT 106.050 189.125 106.305 189.745 ;
        RECT 106.555 189.585 106.785 189.625 ;
        RECT 107.915 189.585 108.165 189.965 ;
        RECT 106.555 189.385 108.165 189.585 ;
        RECT 106.555 189.295 106.740 189.385 ;
        RECT 107.330 189.375 108.165 189.385 ;
        RECT 108.415 189.355 108.665 190.135 ;
        RECT 108.835 189.285 109.095 189.965 ;
        RECT 106.895 189.185 107.225 189.215 ;
        RECT 106.895 189.125 108.695 189.185 ;
        RECT 106.050 189.015 108.755 189.125 ;
        RECT 106.050 188.955 107.225 189.015 ;
        RECT 108.555 188.980 108.755 189.015 ;
        RECT 106.045 188.575 106.535 188.775 ;
        RECT 106.725 188.575 107.200 188.785 ;
        RECT 97.365 187.585 98.110 187.955 ;
        RECT 98.675 187.765 98.930 188.125 ;
        RECT 99.110 187.585 99.440 187.955 ;
        RECT 99.620 187.765 99.845 188.125 ;
        RECT 100.065 187.585 105.410 188.130 ;
        RECT 106.050 187.585 106.505 188.350 ;
        RECT 106.980 188.175 107.200 188.575 ;
        RECT 107.445 188.575 107.775 188.785 ;
        RECT 107.445 188.175 107.655 188.575 ;
        RECT 107.945 188.540 108.355 188.845 ;
        RECT 108.585 188.405 108.755 188.980 ;
        RECT 108.485 188.285 108.755 188.405 ;
        RECT 107.910 188.240 108.755 188.285 ;
        RECT 107.910 188.115 108.665 188.240 ;
        RECT 107.910 187.965 108.080 188.115 ;
        RECT 108.925 188.085 109.095 189.285 ;
        RECT 109.730 189.745 110.065 189.965 ;
        RECT 111.070 189.755 111.425 190.135 ;
        RECT 109.730 189.125 109.985 189.745 ;
        RECT 110.235 189.585 110.465 189.625 ;
        RECT 111.595 189.585 111.845 189.965 ;
        RECT 110.235 189.385 111.845 189.585 ;
        RECT 110.235 189.295 110.420 189.385 ;
        RECT 111.010 189.375 111.845 189.385 ;
        RECT 112.095 189.355 112.345 190.135 ;
        RECT 112.515 189.285 112.775 189.965 ;
        RECT 110.575 189.185 110.905 189.215 ;
        RECT 110.575 189.125 112.375 189.185 ;
        RECT 109.730 189.015 112.435 189.125 ;
        RECT 109.730 188.955 110.905 189.015 ;
        RECT 112.235 188.980 112.435 189.015 ;
        RECT 109.725 188.575 110.215 188.775 ;
        RECT 110.405 188.575 110.880 188.785 ;
        RECT 106.780 187.755 108.080 187.965 ;
        RECT 108.335 187.585 108.665 187.945 ;
        RECT 108.835 187.755 109.095 188.085 ;
        RECT 109.730 187.585 110.185 188.350 ;
        RECT 110.660 188.175 110.880 188.575 ;
        RECT 111.125 188.575 111.455 188.785 ;
        RECT 111.125 188.175 111.335 188.575 ;
        RECT 111.625 188.540 112.035 188.845 ;
        RECT 112.265 188.405 112.435 188.980 ;
        RECT 112.165 188.285 112.435 188.405 ;
        RECT 111.590 188.240 112.435 188.285 ;
        RECT 111.590 188.115 112.345 188.240 ;
        RECT 111.590 187.965 111.760 188.115 ;
        RECT 112.605 188.085 112.775 189.285 ;
        RECT 112.945 188.970 113.235 190.135 ;
        RECT 113.405 188.995 113.790 189.965 ;
        RECT 113.960 189.675 114.285 190.135 ;
        RECT 114.805 189.505 115.085 189.965 ;
        RECT 113.960 189.285 115.085 189.505 ;
        RECT 113.405 188.325 113.685 188.995 ;
        RECT 113.960 188.825 114.410 189.285 ;
        RECT 115.275 189.115 115.675 189.965 ;
        RECT 116.075 189.675 116.345 190.135 ;
        RECT 116.515 189.505 116.800 189.965 ;
        RECT 113.855 188.495 114.410 188.825 ;
        RECT 114.580 188.555 115.675 189.115 ;
        RECT 113.960 188.385 114.410 188.495 ;
        RECT 110.460 187.755 111.760 187.965 ;
        RECT 112.015 187.585 112.345 187.945 ;
        RECT 112.515 187.755 112.775 188.085 ;
        RECT 112.945 187.585 113.235 188.310 ;
        RECT 113.405 187.755 113.790 188.325 ;
        RECT 113.960 188.215 115.085 188.385 ;
        RECT 113.960 187.585 114.285 188.045 ;
        RECT 114.805 187.755 115.085 188.215 ;
        RECT 115.275 187.755 115.675 188.555 ;
        RECT 115.845 189.285 116.800 189.505 ;
        RECT 115.845 188.385 116.055 189.285 ;
        RECT 116.225 188.555 116.915 189.115 ;
        RECT 117.085 189.045 118.755 190.135 ;
        RECT 115.845 188.215 116.800 188.385 ;
        RECT 116.075 187.585 116.345 188.045 ;
        RECT 116.515 187.755 116.800 188.215 ;
        RECT 117.085 188.355 117.835 188.875 ;
        RECT 118.005 188.525 118.755 189.045 ;
        RECT 118.925 188.995 119.310 189.965 ;
        RECT 119.480 189.675 119.805 190.135 ;
        RECT 120.325 189.505 120.605 189.965 ;
        RECT 119.480 189.285 120.605 189.505 ;
        RECT 117.085 187.585 118.755 188.355 ;
        RECT 118.925 188.325 119.205 188.995 ;
        RECT 119.480 188.825 119.930 189.285 ;
        RECT 120.795 189.115 121.195 189.965 ;
        RECT 121.595 189.675 121.865 190.135 ;
        RECT 122.035 189.505 122.320 189.965 ;
        RECT 119.375 188.495 119.930 188.825 ;
        RECT 120.100 188.555 121.195 189.115 ;
        RECT 119.480 188.385 119.930 188.495 ;
        RECT 118.925 187.755 119.310 188.325 ;
        RECT 119.480 188.215 120.605 188.385 ;
        RECT 119.480 187.585 119.805 188.045 ;
        RECT 120.325 187.755 120.605 188.215 ;
        RECT 120.795 187.755 121.195 188.555 ;
        RECT 121.365 189.285 122.320 189.505 ;
        RECT 121.365 188.385 121.575 189.285 ;
        RECT 121.745 188.555 122.435 189.115 ;
        RECT 122.605 189.045 124.275 190.135 ;
        RECT 121.365 188.215 122.320 188.385 ;
        RECT 121.595 187.585 121.865 188.045 ;
        RECT 122.035 187.755 122.320 188.215 ;
        RECT 122.605 188.355 123.355 188.875 ;
        RECT 123.525 188.525 124.275 189.045 ;
        RECT 124.445 188.995 124.725 190.135 ;
        RECT 124.895 188.985 125.225 189.965 ;
        RECT 125.395 188.995 125.655 190.135 ;
        RECT 125.830 189.625 127.485 189.915 ;
        RECT 125.830 189.285 127.420 189.455 ;
        RECT 127.655 189.335 127.935 190.135 ;
        RECT 125.830 188.995 126.150 189.285 ;
        RECT 127.250 189.165 127.420 189.285 ;
        RECT 124.455 188.555 124.790 188.825 ;
        RECT 124.960 188.435 125.130 188.985 ;
        RECT 126.345 188.945 127.060 189.115 ;
        RECT 127.250 188.995 127.975 189.165 ;
        RECT 128.145 188.995 128.415 189.965 ;
        RECT 125.300 188.575 125.635 188.825 ;
        RECT 124.960 188.385 125.135 188.435 ;
        RECT 122.605 187.585 124.275 188.355 ;
        RECT 124.445 187.585 124.755 188.385 ;
        RECT 124.960 187.755 125.655 188.385 ;
        RECT 125.830 188.255 126.180 188.825 ;
        RECT 126.350 188.495 127.060 188.945 ;
        RECT 127.805 188.825 127.975 188.995 ;
        RECT 127.230 188.495 127.635 188.825 ;
        RECT 127.805 188.495 128.075 188.825 ;
        RECT 127.805 188.325 127.975 188.495 ;
        RECT 126.365 188.155 127.975 188.325 ;
        RECT 128.245 188.260 128.415 188.995 ;
        RECT 125.835 187.585 126.165 188.085 ;
        RECT 126.365 187.805 126.535 188.155 ;
        RECT 126.735 187.585 127.065 187.985 ;
        RECT 127.235 187.805 127.405 188.155 ;
        RECT 127.575 187.585 127.955 187.985 ;
        RECT 128.145 187.915 128.415 188.260 ;
        RECT 129.080 189.345 129.615 189.965 ;
        RECT 129.080 188.325 129.395 189.345 ;
        RECT 129.785 189.335 130.115 190.135 ;
        RECT 130.600 189.165 130.990 189.340 ;
        RECT 129.565 188.995 130.990 189.165 ;
        RECT 131.345 189.045 134.855 190.135 ;
        RECT 129.565 188.495 129.735 188.995 ;
        RECT 129.080 187.755 129.695 188.325 ;
        RECT 129.985 188.265 130.250 188.825 ;
        RECT 130.420 188.095 130.590 188.995 ;
        RECT 130.760 188.265 131.115 188.825 ;
        RECT 131.345 188.355 132.995 188.875 ;
        RECT 133.165 188.525 134.855 189.045 ;
        RECT 135.545 188.995 135.755 190.135 ;
        RECT 135.925 188.985 136.255 189.965 ;
        RECT 136.425 188.995 136.655 190.135 ;
        RECT 136.865 189.045 138.535 190.135 ;
        RECT 129.865 187.585 130.080 188.095 ;
        RECT 130.310 187.765 130.590 188.095 ;
        RECT 130.770 187.585 131.010 188.095 ;
        RECT 131.345 187.585 134.855 188.355 ;
        RECT 135.545 187.585 135.755 188.405 ;
        RECT 135.925 188.385 136.175 188.985 ;
        RECT 136.345 188.575 136.675 188.825 ;
        RECT 135.925 187.755 136.255 188.385 ;
        RECT 136.425 187.585 136.655 188.405 ;
        RECT 136.865 188.355 137.615 188.875 ;
        RECT 137.785 188.525 138.535 189.045 ;
        RECT 138.705 188.970 138.995 190.135 ;
        RECT 139.350 189.165 139.740 189.340 ;
        RECT 140.225 189.335 140.555 190.135 ;
        RECT 140.725 189.345 141.260 189.965 ;
        RECT 141.665 189.465 141.945 190.135 ;
        RECT 139.350 188.995 140.775 189.165 ;
        RECT 136.865 187.585 138.535 188.355 ;
        RECT 138.705 187.585 138.995 188.310 ;
        RECT 139.225 188.265 139.580 188.825 ;
        RECT 139.750 188.095 139.920 188.995 ;
        RECT 140.090 188.265 140.355 188.825 ;
        RECT 140.605 188.495 140.775 188.995 ;
        RECT 140.945 188.325 141.260 189.345 ;
        RECT 142.115 189.245 142.415 189.795 ;
        RECT 142.615 189.415 142.945 190.135 ;
        RECT 143.135 189.415 143.595 189.965 ;
        RECT 143.765 189.625 144.025 190.135 ;
        RECT 141.480 188.825 141.745 189.185 ;
        RECT 142.115 189.075 143.055 189.245 ;
        RECT 142.885 188.825 143.055 189.075 ;
        RECT 141.480 188.575 142.155 188.825 ;
        RECT 142.375 188.575 142.715 188.825 ;
        RECT 142.885 188.495 143.175 188.825 ;
        RECT 142.885 188.405 143.055 188.495 ;
        RECT 139.330 187.585 139.570 188.095 ;
        RECT 139.750 187.765 140.030 188.095 ;
        RECT 140.260 187.585 140.475 188.095 ;
        RECT 140.645 187.755 141.260 188.325 ;
        RECT 141.665 188.215 143.055 188.405 ;
        RECT 141.665 187.855 141.995 188.215 ;
        RECT 143.345 188.045 143.595 189.415 ;
        RECT 143.765 188.575 144.105 189.455 ;
        RECT 144.275 188.745 144.445 189.965 ;
        RECT 144.685 189.630 145.300 190.135 ;
        RECT 144.685 189.095 144.935 189.460 ;
        RECT 145.105 189.455 145.300 189.630 ;
        RECT 145.470 189.625 145.945 189.965 ;
        RECT 146.115 189.590 146.330 190.135 ;
        RECT 145.105 189.265 145.435 189.455 ;
        RECT 145.655 189.095 146.370 189.390 ;
        RECT 146.540 189.265 146.815 189.965 ;
        RECT 147.995 189.465 148.165 189.965 ;
        RECT 148.335 189.635 148.665 190.135 ;
        RECT 147.995 189.295 148.660 189.465 ;
        RECT 144.685 188.925 146.475 189.095 ;
        RECT 144.275 188.495 145.070 188.745 ;
        RECT 144.275 188.405 144.525 188.495 ;
        RECT 142.615 187.585 142.865 188.045 ;
        RECT 143.035 187.755 143.595 188.045 ;
        RECT 143.765 187.585 144.025 188.405 ;
        RECT 144.195 187.985 144.525 188.405 ;
        RECT 145.240 188.070 145.495 188.925 ;
        RECT 144.705 187.805 145.495 188.070 ;
        RECT 145.665 188.225 146.075 188.745 ;
        RECT 146.245 188.495 146.475 188.925 ;
        RECT 146.645 188.235 146.815 189.265 ;
        RECT 147.910 188.475 148.260 189.125 ;
        RECT 148.430 188.305 148.660 189.295 ;
        RECT 145.665 187.805 145.865 188.225 ;
        RECT 146.055 187.585 146.385 188.045 ;
        RECT 146.555 187.755 146.815 188.235 ;
        RECT 147.995 188.135 148.660 188.305 ;
        RECT 147.995 187.845 148.165 188.135 ;
        RECT 148.335 187.585 148.665 187.965 ;
        RECT 148.835 187.845 149.020 189.965 ;
        RECT 149.260 189.675 149.525 190.135 ;
        RECT 149.695 189.540 149.945 189.965 ;
        RECT 150.155 189.690 151.260 189.860 ;
        RECT 149.640 189.410 149.945 189.540 ;
        RECT 149.190 188.215 149.470 189.165 ;
        RECT 149.640 188.305 149.810 189.410 ;
        RECT 149.980 188.625 150.220 189.220 ;
        RECT 150.390 189.155 150.920 189.520 ;
        RECT 150.390 188.455 150.560 189.155 ;
        RECT 151.090 189.075 151.260 189.690 ;
        RECT 151.430 189.335 151.600 190.135 ;
        RECT 151.770 189.635 152.020 189.965 ;
        RECT 152.245 189.665 153.130 189.835 ;
        RECT 151.090 188.985 151.600 189.075 ;
        RECT 149.640 188.175 149.865 188.305 ;
        RECT 150.035 188.235 150.560 188.455 ;
        RECT 150.730 188.815 151.600 188.985 ;
        RECT 149.275 187.585 149.525 188.045 ;
        RECT 149.695 188.035 149.865 188.175 ;
        RECT 150.730 188.035 150.900 188.815 ;
        RECT 151.430 188.745 151.600 188.815 ;
        RECT 151.110 188.565 151.310 188.595 ;
        RECT 151.770 188.565 151.940 189.635 ;
        RECT 152.110 188.745 152.300 189.465 ;
        RECT 151.110 188.265 151.940 188.565 ;
        RECT 152.470 188.535 152.790 189.495 ;
        RECT 149.695 187.865 150.030 188.035 ;
        RECT 150.225 187.865 150.900 188.035 ;
        RECT 151.220 187.585 151.590 188.085 ;
        RECT 151.770 188.035 151.940 188.265 ;
        RECT 152.325 188.205 152.790 188.535 ;
        RECT 152.960 188.825 153.130 189.665 ;
        RECT 153.310 189.635 153.625 190.135 ;
        RECT 153.855 189.405 154.195 189.965 ;
        RECT 153.300 189.030 154.195 189.405 ;
        RECT 154.365 189.125 154.535 190.135 ;
        RECT 154.005 188.825 154.195 189.030 ;
        RECT 154.705 189.075 155.035 189.920 ;
        RECT 154.705 188.995 155.095 189.075 ;
        RECT 154.880 188.945 155.095 188.995 ;
        RECT 152.960 188.495 153.835 188.825 ;
        RECT 154.005 188.495 154.755 188.825 ;
        RECT 152.960 188.035 153.130 188.495 ;
        RECT 154.005 188.325 154.205 188.495 ;
        RECT 154.925 188.365 155.095 188.945 ;
        RECT 155.725 189.045 156.935 190.135 ;
        RECT 155.725 188.505 156.245 189.045 ;
        RECT 154.870 188.325 155.095 188.365 ;
        RECT 156.415 188.335 156.935 188.875 ;
        RECT 151.770 187.865 152.175 188.035 ;
        RECT 152.345 187.865 153.130 188.035 ;
        RECT 153.405 187.585 153.615 188.115 ;
        RECT 153.875 187.800 154.205 188.325 ;
        RECT 154.715 188.240 155.095 188.325 ;
        RECT 154.375 187.585 154.545 188.195 ;
        RECT 154.715 187.805 155.045 188.240 ;
        RECT 155.725 187.585 156.935 188.335 ;
        RECT 22.700 187.415 157.020 187.585 ;
        RECT 22.785 186.665 23.995 187.415 ;
        RECT 24.165 186.665 25.375 187.415 ;
        RECT 25.545 186.740 25.805 187.245 ;
        RECT 25.985 187.035 26.315 187.415 ;
        RECT 26.495 186.865 26.665 187.245 ;
        RECT 22.785 186.125 23.305 186.665 ;
        RECT 23.475 185.955 23.995 186.495 ;
        RECT 24.165 186.125 24.685 186.665 ;
        RECT 24.855 185.955 25.375 186.495 ;
        RECT 22.785 184.865 23.995 185.955 ;
        RECT 24.165 184.865 25.375 185.955 ;
        RECT 25.545 185.940 25.715 186.740 ;
        RECT 26.000 186.695 26.665 186.865 ;
        RECT 26.000 186.440 26.170 186.695 ;
        RECT 26.925 186.645 30.435 187.415 ;
        RECT 31.525 186.765 31.785 187.245 ;
        RECT 31.955 186.875 32.205 187.415 ;
        RECT 25.885 186.110 26.170 186.440 ;
        RECT 26.405 186.145 26.735 186.515 ;
        RECT 26.925 186.125 28.575 186.645 ;
        RECT 26.000 185.965 26.170 186.110 ;
        RECT 25.545 185.035 25.815 185.940 ;
        RECT 26.000 185.795 26.665 185.965 ;
        RECT 28.745 185.955 30.435 186.475 ;
        RECT 25.985 184.865 26.315 185.625 ;
        RECT 26.495 185.035 26.665 185.795 ;
        RECT 26.925 184.865 30.435 185.955 ;
        RECT 31.525 185.735 31.695 186.765 ;
        RECT 32.375 186.710 32.595 187.195 ;
        RECT 31.865 186.115 32.095 186.510 ;
        RECT 32.265 186.285 32.595 186.710 ;
        RECT 32.765 187.035 33.655 187.205 ;
        RECT 32.765 186.310 32.935 187.035 ;
        RECT 33.105 186.480 33.655 186.865 ;
        RECT 33.860 186.675 34.475 187.245 ;
        RECT 34.645 186.905 34.860 187.415 ;
        RECT 35.090 186.905 35.370 187.235 ;
        RECT 35.550 186.905 35.790 187.415 ;
        RECT 32.765 186.240 33.655 186.310 ;
        RECT 32.760 186.215 33.655 186.240 ;
        RECT 32.750 186.200 33.655 186.215 ;
        RECT 32.745 186.185 33.655 186.200 ;
        RECT 32.735 186.180 33.655 186.185 ;
        RECT 32.730 186.170 33.655 186.180 ;
        RECT 32.725 186.160 33.655 186.170 ;
        RECT 32.715 186.155 33.655 186.160 ;
        RECT 32.705 186.145 33.655 186.155 ;
        RECT 32.695 186.140 33.655 186.145 ;
        RECT 32.695 186.135 33.030 186.140 ;
        RECT 32.680 186.130 33.030 186.135 ;
        RECT 32.665 186.120 33.030 186.130 ;
        RECT 32.640 186.115 33.030 186.120 ;
        RECT 31.865 186.110 33.030 186.115 ;
        RECT 31.865 186.075 33.000 186.110 ;
        RECT 31.865 186.050 32.965 186.075 ;
        RECT 31.865 186.020 32.935 186.050 ;
        RECT 31.865 185.990 32.915 186.020 ;
        RECT 31.865 185.960 32.895 185.990 ;
        RECT 31.865 185.950 32.825 185.960 ;
        RECT 31.865 185.940 32.800 185.950 ;
        RECT 31.865 185.925 32.780 185.940 ;
        RECT 31.865 185.910 32.760 185.925 ;
        RECT 31.970 185.900 32.755 185.910 ;
        RECT 31.970 185.865 32.740 185.900 ;
        RECT 31.525 185.035 31.800 185.735 ;
        RECT 31.970 185.615 32.725 185.865 ;
        RECT 32.895 185.545 33.225 185.790 ;
        RECT 33.395 185.690 33.655 186.140 ;
        RECT 33.040 185.520 33.225 185.545 ;
        RECT 33.860 185.655 34.175 186.675 ;
        RECT 34.345 186.005 34.515 186.505 ;
        RECT 34.765 186.175 35.030 186.735 ;
        RECT 35.200 186.005 35.370 186.905 ;
        RECT 35.540 186.175 35.895 186.735 ;
        RECT 36.165 186.595 36.395 187.415 ;
        RECT 36.565 186.615 36.895 187.245 ;
        RECT 36.145 186.175 36.475 186.425 ;
        RECT 36.645 186.015 36.895 186.615 ;
        RECT 37.065 186.595 37.275 187.415 ;
        RECT 37.505 186.645 39.175 187.415 ;
        RECT 39.810 186.910 40.145 187.415 ;
        RECT 40.315 186.845 40.555 187.220 ;
        RECT 40.835 187.085 41.005 187.230 ;
        RECT 40.835 186.890 41.210 187.085 ;
        RECT 41.570 186.920 41.965 187.415 ;
        RECT 37.505 186.125 38.255 186.645 ;
        RECT 34.345 185.835 35.770 186.005 ;
        RECT 33.040 185.420 33.655 185.520 ;
        RECT 31.970 184.865 32.225 185.410 ;
        RECT 32.395 185.035 32.875 185.375 ;
        RECT 33.050 184.865 33.655 185.420 ;
        RECT 33.860 185.035 34.395 185.655 ;
        RECT 34.565 184.865 34.895 185.665 ;
        RECT 35.380 185.660 35.770 185.835 ;
        RECT 36.165 184.865 36.395 186.005 ;
        RECT 36.565 185.035 36.895 186.015 ;
        RECT 37.065 184.865 37.275 186.005 ;
        RECT 38.425 185.955 39.175 186.475 ;
        RECT 37.505 184.865 39.175 185.955 ;
        RECT 39.865 185.885 40.165 186.735 ;
        RECT 40.335 186.695 40.555 186.845 ;
        RECT 40.335 186.365 40.870 186.695 ;
        RECT 41.040 186.555 41.210 186.890 ;
        RECT 42.135 186.725 42.375 187.245 ;
        RECT 40.335 185.715 40.570 186.365 ;
        RECT 41.040 186.195 42.025 186.555 ;
        RECT 39.895 185.485 40.570 185.715 ;
        RECT 40.740 186.175 42.025 186.195 ;
        RECT 40.740 186.025 41.600 186.175 ;
        RECT 39.895 185.055 40.065 185.485 ;
        RECT 40.235 184.865 40.565 185.315 ;
        RECT 40.740 185.080 41.025 186.025 ;
        RECT 42.200 185.920 42.375 186.725 ;
        RECT 42.565 186.645 45.155 187.415 ;
        RECT 42.565 186.125 43.775 186.645 ;
        RECT 43.945 185.955 45.155 186.475 ;
        RECT 41.200 185.545 41.895 185.855 ;
        RECT 41.205 184.865 41.890 185.335 ;
        RECT 42.070 185.135 42.375 185.920 ;
        RECT 42.565 184.865 45.155 185.955 ;
        RECT 45.795 185.045 46.055 187.235 ;
        RECT 46.315 187.045 46.985 187.415 ;
        RECT 47.165 186.865 47.475 187.235 ;
        RECT 46.245 186.665 47.475 186.865 ;
        RECT 46.245 185.995 46.535 186.665 ;
        RECT 47.655 186.485 47.885 187.125 ;
        RECT 48.065 186.685 48.355 187.415 ;
        RECT 48.545 186.690 48.835 187.415 ;
        RECT 49.055 186.875 49.280 187.235 ;
        RECT 49.460 187.045 49.790 187.415 ;
        RECT 49.970 186.875 50.225 187.235 ;
        RECT 50.790 187.045 51.535 187.415 ;
        RECT 49.055 186.685 51.540 186.875 ;
        RECT 46.715 186.175 47.180 186.485 ;
        RECT 47.360 186.175 47.885 186.485 ;
        RECT 48.065 186.175 48.365 186.505 ;
        RECT 49.015 186.175 49.285 186.505 ;
        RECT 49.465 186.175 49.900 186.505 ;
        RECT 50.080 186.175 50.655 186.505 ;
        RECT 50.835 186.175 51.115 186.505 ;
        RECT 46.245 185.775 47.015 185.995 ;
        RECT 46.225 184.865 46.565 185.595 ;
        RECT 46.745 185.045 47.015 185.775 ;
        RECT 47.195 185.755 48.355 185.995 ;
        RECT 47.195 185.045 47.425 185.755 ;
        RECT 47.595 184.865 47.925 185.575 ;
        RECT 48.095 185.045 48.355 185.755 ;
        RECT 48.545 184.865 48.835 186.030 ;
        RECT 51.315 185.995 51.540 186.685 ;
        RECT 49.045 185.815 51.540 185.995 ;
        RECT 51.715 185.815 52.050 187.235 ;
        RECT 53.235 186.865 53.405 187.155 ;
        RECT 53.575 187.035 53.905 187.415 ;
        RECT 53.235 186.695 53.900 186.865 ;
        RECT 53.150 185.875 53.500 186.525 ;
        RECT 49.045 185.045 49.335 185.815 ;
        RECT 49.905 185.405 51.095 185.635 ;
        RECT 49.905 185.045 50.165 185.405 ;
        RECT 50.335 184.865 50.665 185.235 ;
        RECT 50.835 185.045 51.095 185.405 ;
        RECT 51.285 184.865 51.615 185.585 ;
        RECT 51.785 185.045 52.050 185.815 ;
        RECT 53.670 185.705 53.900 186.695 ;
        RECT 53.235 185.535 53.900 185.705 ;
        RECT 53.235 185.035 53.405 185.535 ;
        RECT 53.575 184.865 53.905 185.365 ;
        RECT 54.075 185.035 54.260 187.155 ;
        RECT 54.515 186.955 54.765 187.415 ;
        RECT 54.935 186.965 55.270 187.135 ;
        RECT 55.465 186.965 56.140 187.135 ;
        RECT 54.935 186.825 55.105 186.965 ;
        RECT 54.430 185.835 54.710 186.785 ;
        RECT 54.880 186.695 55.105 186.825 ;
        RECT 54.880 185.590 55.050 186.695 ;
        RECT 55.275 186.545 55.800 186.765 ;
        RECT 55.220 185.780 55.460 186.375 ;
        RECT 55.630 185.845 55.800 186.545 ;
        RECT 55.970 186.185 56.140 186.965 ;
        RECT 56.460 186.915 56.830 187.415 ;
        RECT 57.010 186.965 57.415 187.135 ;
        RECT 57.585 186.965 58.370 187.135 ;
        RECT 57.010 186.735 57.180 186.965 ;
        RECT 56.350 186.435 57.180 186.735 ;
        RECT 57.565 186.465 58.030 186.795 ;
        RECT 56.350 186.405 56.550 186.435 ;
        RECT 56.670 186.185 56.840 186.255 ;
        RECT 55.970 186.015 56.840 186.185 ;
        RECT 56.330 185.925 56.840 186.015 ;
        RECT 54.880 185.460 55.185 185.590 ;
        RECT 55.630 185.480 56.160 185.845 ;
        RECT 54.500 184.865 54.765 185.325 ;
        RECT 54.935 185.035 55.185 185.460 ;
        RECT 56.330 185.310 56.500 185.925 ;
        RECT 55.395 185.140 56.500 185.310 ;
        RECT 56.670 184.865 56.840 185.665 ;
        RECT 57.010 185.365 57.180 186.435 ;
        RECT 57.350 185.535 57.540 186.255 ;
        RECT 57.710 185.505 58.030 186.465 ;
        RECT 58.200 186.505 58.370 186.965 ;
        RECT 58.645 186.885 58.855 187.415 ;
        RECT 59.115 186.675 59.445 187.200 ;
        RECT 59.615 186.805 59.785 187.415 ;
        RECT 59.955 186.760 60.285 187.195 ;
        RECT 59.955 186.675 60.335 186.760 ;
        RECT 59.245 186.505 59.445 186.675 ;
        RECT 60.110 186.635 60.335 186.675 ;
        RECT 58.200 186.175 59.075 186.505 ;
        RECT 59.245 186.175 59.995 186.505 ;
        RECT 57.010 185.035 57.260 185.365 ;
        RECT 58.200 185.335 58.370 186.175 ;
        RECT 59.245 185.970 59.435 186.175 ;
        RECT 60.165 186.055 60.335 186.635 ;
        RECT 60.505 186.665 61.715 187.415 ;
        RECT 61.885 187.035 62.775 187.205 ;
        RECT 60.505 186.125 61.025 186.665 ;
        RECT 60.120 186.005 60.335 186.055 ;
        RECT 58.540 185.595 59.435 185.970 ;
        RECT 59.945 185.925 60.335 186.005 ;
        RECT 61.195 185.955 61.715 186.495 ;
        RECT 61.885 186.480 62.435 186.865 ;
        RECT 62.605 186.310 62.775 187.035 ;
        RECT 57.485 185.165 58.370 185.335 ;
        RECT 58.550 184.865 58.865 185.365 ;
        RECT 59.095 185.035 59.435 185.595 ;
        RECT 59.605 184.865 59.775 185.875 ;
        RECT 59.945 185.080 60.275 185.925 ;
        RECT 60.505 184.865 61.715 185.955 ;
        RECT 61.885 186.240 62.775 186.310 ;
        RECT 62.945 186.735 63.165 187.195 ;
        RECT 63.335 186.875 63.585 187.415 ;
        RECT 63.755 186.765 64.015 187.245 ;
        RECT 62.945 186.710 63.195 186.735 ;
        RECT 62.945 186.285 63.275 186.710 ;
        RECT 61.885 186.215 62.780 186.240 ;
        RECT 61.885 186.200 62.790 186.215 ;
        RECT 61.885 186.185 62.795 186.200 ;
        RECT 61.885 186.180 62.805 186.185 ;
        RECT 61.885 186.170 62.810 186.180 ;
        RECT 61.885 186.160 62.815 186.170 ;
        RECT 61.885 186.155 62.825 186.160 ;
        RECT 61.885 186.145 62.835 186.155 ;
        RECT 61.885 186.140 62.845 186.145 ;
        RECT 61.885 185.690 62.145 186.140 ;
        RECT 62.510 186.135 62.845 186.140 ;
        RECT 62.510 186.130 62.860 186.135 ;
        RECT 62.510 186.120 62.875 186.130 ;
        RECT 62.510 186.115 62.900 186.120 ;
        RECT 63.445 186.115 63.675 186.510 ;
        RECT 62.510 186.110 63.675 186.115 ;
        RECT 62.540 186.075 63.675 186.110 ;
        RECT 62.575 186.050 63.675 186.075 ;
        RECT 62.605 186.020 63.675 186.050 ;
        RECT 62.625 185.990 63.675 186.020 ;
        RECT 62.645 185.960 63.675 185.990 ;
        RECT 62.715 185.950 63.675 185.960 ;
        RECT 62.740 185.940 63.675 185.950 ;
        RECT 62.760 185.925 63.675 185.940 ;
        RECT 62.780 185.910 63.675 185.925 ;
        RECT 62.785 185.900 63.570 185.910 ;
        RECT 62.800 185.865 63.570 185.900 ;
        RECT 62.315 185.545 62.645 185.790 ;
        RECT 62.815 185.615 63.570 185.865 ;
        RECT 63.845 185.735 64.015 186.765 ;
        RECT 62.315 185.520 62.500 185.545 ;
        RECT 61.885 185.420 62.500 185.520 ;
        RECT 61.885 184.865 62.490 185.420 ;
        RECT 62.665 185.035 63.145 185.375 ;
        RECT 63.315 184.865 63.570 185.410 ;
        RECT 63.740 185.035 64.015 185.735 ;
        RECT 64.195 185.045 64.455 187.235 ;
        RECT 64.715 187.045 65.385 187.415 ;
        RECT 65.565 186.865 65.875 187.235 ;
        RECT 64.645 186.665 65.875 186.865 ;
        RECT 64.645 185.995 64.935 186.665 ;
        RECT 66.055 186.485 66.285 187.125 ;
        RECT 66.465 186.685 66.755 187.415 ;
        RECT 67.865 186.675 68.250 187.245 ;
        RECT 68.420 186.955 68.745 187.415 ;
        RECT 69.265 186.785 69.545 187.245 ;
        RECT 65.115 186.175 65.580 186.485 ;
        RECT 65.760 186.175 66.285 186.485 ;
        RECT 66.465 186.175 66.765 186.505 ;
        RECT 67.865 186.005 68.145 186.675 ;
        RECT 68.420 186.615 69.545 186.785 ;
        RECT 68.420 186.505 68.870 186.615 ;
        RECT 68.315 186.175 68.870 186.505 ;
        RECT 69.735 186.445 70.135 187.245 ;
        RECT 70.535 186.955 70.805 187.415 ;
        RECT 70.975 186.785 71.260 187.245 ;
        RECT 64.645 185.775 65.415 185.995 ;
        RECT 64.625 184.865 64.965 185.595 ;
        RECT 65.145 185.045 65.415 185.775 ;
        RECT 65.595 185.755 66.755 185.995 ;
        RECT 65.595 185.045 65.825 185.755 ;
        RECT 65.995 184.865 66.325 185.575 ;
        RECT 66.495 185.045 66.755 185.755 ;
        RECT 67.865 185.035 68.250 186.005 ;
        RECT 68.420 185.715 68.870 186.175 ;
        RECT 69.040 185.885 70.135 186.445 ;
        RECT 68.420 185.495 69.545 185.715 ;
        RECT 68.420 184.865 68.745 185.325 ;
        RECT 69.265 185.035 69.545 185.495 ;
        RECT 69.735 185.035 70.135 185.885 ;
        RECT 70.305 186.615 71.260 186.785 ;
        RECT 72.005 186.765 72.265 187.245 ;
        RECT 72.435 186.875 72.685 187.415 ;
        RECT 70.305 185.715 70.515 186.615 ;
        RECT 70.685 185.885 71.375 186.445 ;
        RECT 72.005 185.735 72.175 186.765 ;
        RECT 72.855 186.735 73.075 187.195 ;
        RECT 72.825 186.710 73.075 186.735 ;
        RECT 72.345 186.115 72.575 186.510 ;
        RECT 72.745 186.285 73.075 186.710 ;
        RECT 73.245 187.035 74.135 187.205 ;
        RECT 73.245 186.310 73.415 187.035 ;
        RECT 73.585 186.480 74.135 186.865 ;
        RECT 74.305 186.690 74.595 187.415 ;
        RECT 74.765 186.645 76.435 187.415 ;
        RECT 76.625 186.685 76.915 187.415 ;
        RECT 73.245 186.240 74.135 186.310 ;
        RECT 73.240 186.215 74.135 186.240 ;
        RECT 73.230 186.200 74.135 186.215 ;
        RECT 73.225 186.185 74.135 186.200 ;
        RECT 73.215 186.180 74.135 186.185 ;
        RECT 73.210 186.170 74.135 186.180 ;
        RECT 73.205 186.160 74.135 186.170 ;
        RECT 73.195 186.155 74.135 186.160 ;
        RECT 73.185 186.145 74.135 186.155 ;
        RECT 73.175 186.140 74.135 186.145 ;
        RECT 73.175 186.135 73.510 186.140 ;
        RECT 73.160 186.130 73.510 186.135 ;
        RECT 73.145 186.120 73.510 186.130 ;
        RECT 73.120 186.115 73.510 186.120 ;
        RECT 72.345 186.110 73.510 186.115 ;
        RECT 72.345 186.075 73.480 186.110 ;
        RECT 72.345 186.050 73.445 186.075 ;
        RECT 72.345 186.020 73.415 186.050 ;
        RECT 72.345 185.990 73.395 186.020 ;
        RECT 72.345 185.960 73.375 185.990 ;
        RECT 72.345 185.950 73.305 185.960 ;
        RECT 72.345 185.940 73.280 185.950 ;
        RECT 72.345 185.925 73.260 185.940 ;
        RECT 72.345 185.910 73.240 185.925 ;
        RECT 72.450 185.900 73.235 185.910 ;
        RECT 72.450 185.865 73.220 185.900 ;
        RECT 70.305 185.495 71.260 185.715 ;
        RECT 70.535 184.865 70.805 185.325 ;
        RECT 70.975 185.035 71.260 185.495 ;
        RECT 72.005 185.035 72.280 185.735 ;
        RECT 72.450 185.615 73.205 185.865 ;
        RECT 73.375 185.545 73.705 185.790 ;
        RECT 73.875 185.690 74.135 186.140 ;
        RECT 74.765 186.125 75.515 186.645 ;
        RECT 73.520 185.520 73.705 185.545 ;
        RECT 73.520 185.420 74.135 185.520 ;
        RECT 72.450 184.865 72.705 185.410 ;
        RECT 72.875 185.035 73.355 185.375 ;
        RECT 73.530 184.865 74.135 185.420 ;
        RECT 74.305 184.865 74.595 186.030 ;
        RECT 75.685 185.955 76.435 186.475 ;
        RECT 76.615 186.175 76.915 186.505 ;
        RECT 77.095 186.485 77.325 187.125 ;
        RECT 77.505 186.865 77.815 187.235 ;
        RECT 77.995 187.045 78.665 187.415 ;
        RECT 77.505 186.665 78.735 186.865 ;
        RECT 77.095 186.175 77.620 186.485 ;
        RECT 77.800 186.175 78.265 186.485 ;
        RECT 78.445 185.995 78.735 186.665 ;
        RECT 74.765 184.865 76.435 185.955 ;
        RECT 76.625 185.755 77.785 185.995 ;
        RECT 76.625 185.045 76.885 185.755 ;
        RECT 77.055 184.865 77.385 185.575 ;
        RECT 77.555 185.045 77.785 185.755 ;
        RECT 77.965 185.775 78.735 185.995 ;
        RECT 77.965 185.045 78.235 185.775 ;
        RECT 78.415 184.865 78.755 185.595 ;
        RECT 78.925 185.045 79.185 187.235 ;
        RECT 79.375 185.045 79.635 187.235 ;
        RECT 79.895 187.045 80.565 187.415 ;
        RECT 80.745 186.865 81.055 187.235 ;
        RECT 79.825 186.665 81.055 186.865 ;
        RECT 79.825 185.995 80.115 186.665 ;
        RECT 81.235 186.485 81.465 187.125 ;
        RECT 81.645 186.685 81.935 187.415 ;
        RECT 82.125 186.665 83.335 187.415 ;
        RECT 83.525 186.685 83.815 187.415 ;
        RECT 80.295 186.175 80.760 186.485 ;
        RECT 80.940 186.175 81.465 186.485 ;
        RECT 81.645 186.175 81.945 186.505 ;
        RECT 82.125 186.125 82.645 186.665 ;
        RECT 79.825 185.775 80.595 185.995 ;
        RECT 79.805 184.865 80.145 185.595 ;
        RECT 80.325 185.045 80.595 185.775 ;
        RECT 80.775 185.755 81.935 185.995 ;
        RECT 82.815 185.955 83.335 186.495 ;
        RECT 83.515 186.175 83.815 186.505 ;
        RECT 83.995 186.485 84.225 187.125 ;
        RECT 84.405 186.865 84.715 187.235 ;
        RECT 84.895 187.045 85.565 187.415 ;
        RECT 84.405 186.665 85.635 186.865 ;
        RECT 83.995 186.175 84.520 186.485 ;
        RECT 84.700 186.175 85.165 186.485 ;
        RECT 85.345 185.995 85.635 186.665 ;
        RECT 80.775 185.045 81.005 185.755 ;
        RECT 81.175 184.865 81.505 185.575 ;
        RECT 81.675 185.045 81.935 185.755 ;
        RECT 82.125 184.865 83.335 185.955 ;
        RECT 83.525 185.755 84.685 185.995 ;
        RECT 83.525 185.045 83.785 185.755 ;
        RECT 83.955 184.865 84.285 185.575 ;
        RECT 84.455 185.045 84.685 185.755 ;
        RECT 84.865 185.775 85.635 185.995 ;
        RECT 84.865 185.045 85.135 185.775 ;
        RECT 85.315 184.865 85.655 185.595 ;
        RECT 85.825 185.045 86.085 187.235 ;
        RECT 86.265 186.870 91.610 187.415 ;
        RECT 91.785 186.870 97.130 187.415 ;
        RECT 98.230 186.885 98.520 187.235 ;
        RECT 98.715 187.055 99.045 187.415 ;
        RECT 99.215 186.885 99.445 187.190 ;
        RECT 87.850 186.040 88.190 186.870 ;
        RECT 89.670 185.300 90.020 186.550 ;
        RECT 93.370 186.040 93.710 186.870 ;
        RECT 98.230 186.715 99.445 186.885 ;
        RECT 99.635 186.735 99.805 187.110 ;
        RECT 99.635 186.565 99.835 186.735 ;
        RECT 100.065 186.690 100.355 187.415 ;
        RECT 100.545 186.785 100.875 187.245 ;
        RECT 101.055 186.955 101.225 187.415 ;
        RECT 101.405 186.785 101.735 187.245 ;
        RECT 101.965 186.955 102.135 187.415 ;
        RECT 102.375 187.075 103.565 187.245 ;
        RECT 102.375 186.785 102.705 187.075 ;
        RECT 103.255 186.905 103.565 187.075 ;
        RECT 100.545 186.615 102.705 186.785 ;
        RECT 95.190 185.300 95.540 186.550 ;
        RECT 99.635 186.545 99.805 186.565 ;
        RECT 98.290 186.395 98.550 186.505 ;
        RECT 98.285 186.225 98.550 186.395 ;
        RECT 98.290 186.175 98.550 186.225 ;
        RECT 98.730 186.175 99.115 186.505 ;
        RECT 99.285 186.375 99.805 186.545 ;
        RECT 86.265 184.865 91.610 185.300 ;
        RECT 91.785 184.865 97.130 185.300 ;
        RECT 98.230 184.865 98.550 186.005 ;
        RECT 98.730 185.125 98.925 186.175 ;
        RECT 99.285 185.995 99.455 186.375 ;
        RECT 99.105 185.715 99.455 185.995 ;
        RECT 99.645 185.845 99.890 186.205 ;
        RECT 100.560 186.055 100.890 186.445 ;
        RECT 101.060 186.225 101.860 186.425 ;
        RECT 102.040 186.055 102.535 186.425 ;
        RECT 99.105 185.035 99.435 185.715 ;
        RECT 99.635 184.865 99.890 185.665 ;
        RECT 100.065 184.865 100.355 186.030 ;
        RECT 100.560 185.885 102.535 186.055 ;
        RECT 102.875 185.715 103.085 186.905 ;
        RECT 103.745 186.740 104.020 187.085 ;
        RECT 104.210 187.015 104.585 187.415 ;
        RECT 104.755 186.845 104.925 187.195 ;
        RECT 105.095 187.015 105.425 187.415 ;
        RECT 105.595 186.845 105.855 187.245 ;
        RECT 103.255 186.100 103.570 186.735 ;
        RECT 103.745 186.005 103.915 186.740 ;
        RECT 104.190 186.675 105.855 186.845 ;
        RECT 104.190 186.505 104.360 186.675 ;
        RECT 106.035 186.595 106.365 187.015 ;
        RECT 106.535 186.595 106.795 187.415 ;
        RECT 106.035 186.505 106.285 186.595 ;
        RECT 106.965 186.580 107.255 187.415 ;
        RECT 107.425 187.015 108.380 187.185 ;
        RECT 108.795 187.025 109.125 187.415 ;
        RECT 104.085 186.175 104.360 186.505 ;
        RECT 104.530 186.175 105.355 186.505 ;
        RECT 105.570 186.175 106.285 186.505 ;
        RECT 106.455 186.175 106.790 186.425 ;
        RECT 104.190 186.005 104.360 186.175 ;
        RECT 100.545 184.865 100.875 185.715 ;
        RECT 101.045 185.205 101.265 185.715 ;
        RECT 101.435 185.535 103.085 185.715 ;
        RECT 101.435 185.375 101.735 185.535 ;
        RECT 101.965 185.205 102.155 185.365 ;
        RECT 101.045 185.035 102.155 185.205 ;
        RECT 102.350 184.865 102.680 185.325 ;
        RECT 102.850 185.035 103.085 185.535 ;
        RECT 103.255 184.865 103.565 185.930 ;
        RECT 103.745 185.035 104.020 186.005 ;
        RECT 104.190 185.835 104.850 186.005 ;
        RECT 105.110 185.885 105.355 186.175 ;
        RECT 104.680 185.715 104.850 185.835 ;
        RECT 105.525 185.715 105.855 186.005 ;
        RECT 104.230 184.865 104.510 185.665 ;
        RECT 104.680 185.545 105.855 185.715 ;
        RECT 106.115 185.615 106.285 186.175 ;
        RECT 107.425 186.135 107.595 187.015 ;
        RECT 109.295 186.845 109.465 187.165 ;
        RECT 109.635 187.025 109.965 187.415 ;
        RECT 107.765 186.675 110.015 186.845 ;
        RECT 107.765 186.175 107.995 186.675 ;
        RECT 108.165 186.255 108.540 186.425 ;
        RECT 104.680 185.045 106.295 185.375 ;
        RECT 106.535 184.865 106.795 186.005 ;
        RECT 106.965 185.965 107.595 186.135 ;
        RECT 108.370 186.055 108.540 186.255 ;
        RECT 108.710 186.225 109.260 186.425 ;
        RECT 109.430 186.055 109.675 186.505 ;
        RECT 106.965 185.035 107.285 185.965 ;
        RECT 108.370 185.885 109.675 186.055 ;
        RECT 109.845 185.715 110.015 186.675 ;
        RECT 110.190 186.650 110.645 187.415 ;
        RECT 110.920 187.035 112.220 187.245 ;
        RECT 112.475 187.055 112.805 187.415 ;
        RECT 112.050 186.885 112.220 187.035 ;
        RECT 112.975 186.915 113.235 187.245 ;
        RECT 111.120 186.425 111.340 186.825 ;
        RECT 110.185 186.225 110.675 186.425 ;
        RECT 110.865 186.215 111.340 186.425 ;
        RECT 111.585 186.425 111.795 186.825 ;
        RECT 112.050 186.760 112.805 186.885 ;
        RECT 112.050 186.715 112.895 186.760 ;
        RECT 112.625 186.595 112.895 186.715 ;
        RECT 111.585 186.215 111.915 186.425 ;
        RECT 112.085 186.155 112.495 186.460 ;
        RECT 107.465 185.545 108.705 185.715 ;
        RECT 107.465 185.035 107.865 185.545 ;
        RECT 108.035 184.865 108.205 185.375 ;
        RECT 108.375 185.035 108.705 185.545 ;
        RECT 108.875 184.865 109.045 185.715 ;
        RECT 109.635 185.035 110.015 185.715 ;
        RECT 110.190 185.985 111.365 186.045 ;
        RECT 112.725 186.020 112.895 186.595 ;
        RECT 112.695 185.985 112.895 186.020 ;
        RECT 110.190 185.875 112.895 185.985 ;
        RECT 110.190 185.255 110.445 185.875 ;
        RECT 111.035 185.815 112.835 185.875 ;
        RECT 111.035 185.785 111.365 185.815 ;
        RECT 113.065 185.715 113.235 186.915 ;
        RECT 110.695 185.615 110.880 185.705 ;
        RECT 111.470 185.615 112.305 185.625 ;
        RECT 110.695 185.415 112.305 185.615 ;
        RECT 110.695 185.375 110.925 185.415 ;
        RECT 110.190 185.035 110.525 185.255 ;
        RECT 111.530 184.865 111.885 185.245 ;
        RECT 112.055 185.035 112.305 185.415 ;
        RECT 112.555 184.865 112.805 185.645 ;
        RECT 112.975 185.035 113.235 185.715 ;
        RECT 113.405 186.675 113.790 187.245 ;
        RECT 113.960 186.955 114.285 187.415 ;
        RECT 114.805 186.785 115.085 187.245 ;
        RECT 113.405 186.005 113.685 186.675 ;
        RECT 113.960 186.615 115.085 186.785 ;
        RECT 113.960 186.505 114.410 186.615 ;
        RECT 113.855 186.175 114.410 186.505 ;
        RECT 115.275 186.445 115.675 187.245 ;
        RECT 116.075 186.955 116.345 187.415 ;
        RECT 116.515 186.785 116.800 187.245 ;
        RECT 113.405 185.035 113.790 186.005 ;
        RECT 113.960 185.715 114.410 186.175 ;
        RECT 114.580 185.885 115.675 186.445 ;
        RECT 113.960 185.495 115.085 185.715 ;
        RECT 113.960 184.865 114.285 185.325 ;
        RECT 114.805 185.035 115.085 185.495 ;
        RECT 115.275 185.035 115.675 185.885 ;
        RECT 115.845 186.615 116.800 186.785 ;
        RECT 118.005 186.675 118.390 187.245 ;
        RECT 118.560 186.955 118.885 187.415 ;
        RECT 119.405 186.785 119.685 187.245 ;
        RECT 115.845 185.715 116.055 186.615 ;
        RECT 116.225 185.885 116.915 186.445 ;
        RECT 118.005 186.005 118.285 186.675 ;
        RECT 118.560 186.615 119.685 186.785 ;
        RECT 118.560 186.505 119.010 186.615 ;
        RECT 118.455 186.175 119.010 186.505 ;
        RECT 119.875 186.445 120.275 187.245 ;
        RECT 120.675 186.955 120.945 187.415 ;
        RECT 121.115 186.785 121.400 187.245 ;
        RECT 115.845 185.495 116.800 185.715 ;
        RECT 116.075 184.865 116.345 185.325 ;
        RECT 116.515 185.035 116.800 185.495 ;
        RECT 118.005 185.035 118.390 186.005 ;
        RECT 118.560 185.715 119.010 186.175 ;
        RECT 119.180 185.885 120.275 186.445 ;
        RECT 118.560 185.495 119.685 185.715 ;
        RECT 118.560 184.865 118.885 185.325 ;
        RECT 119.405 185.035 119.685 185.495 ;
        RECT 119.875 185.035 120.275 185.885 ;
        RECT 120.445 186.615 121.400 186.785 ;
        RECT 120.445 185.715 120.655 186.615 ;
        RECT 120.825 185.885 121.515 186.445 ;
        RECT 120.445 185.495 121.400 185.715 ;
        RECT 120.675 184.865 120.945 185.325 ;
        RECT 121.115 185.035 121.400 185.495 ;
        RECT 122.145 185.035 122.425 187.135 ;
        RECT 122.655 186.955 122.825 187.415 ;
        RECT 123.095 187.025 124.345 187.205 ;
        RECT 123.480 186.785 123.845 186.855 ;
        RECT 122.595 186.605 123.845 186.785 ;
        RECT 124.015 186.805 124.345 187.025 ;
        RECT 124.515 186.975 124.685 187.415 ;
        RECT 124.855 186.805 125.195 187.220 ;
        RECT 124.015 186.635 125.195 186.805 ;
        RECT 125.825 186.690 126.115 187.415 ;
        RECT 126.290 187.015 127.545 187.245 ;
        RECT 127.715 187.015 128.385 187.415 ;
        RECT 127.215 186.845 127.545 187.015 ;
        RECT 128.555 186.845 128.725 187.125 ;
        RECT 122.595 186.005 122.870 186.605 ;
        RECT 126.290 186.505 126.545 186.815 ;
        RECT 126.715 186.675 127.045 186.845 ;
        RECT 127.215 186.675 128.725 186.845 ;
        RECT 128.895 186.675 129.335 187.415 ;
        RECT 129.505 186.870 134.850 187.415 ;
        RECT 123.040 186.175 123.395 186.425 ;
        RECT 123.590 186.395 124.055 186.425 ;
        RECT 123.585 186.225 124.055 186.395 ;
        RECT 123.590 186.175 124.055 186.225 ;
        RECT 124.225 186.175 124.555 186.425 ;
        RECT 124.730 186.225 125.195 186.425 ;
        RECT 126.290 186.175 126.560 186.505 ;
        RECT 124.375 186.055 124.555 186.175 ;
        RECT 122.595 185.795 124.205 186.005 ;
        RECT 124.375 185.885 124.705 186.055 ;
        RECT 123.795 185.695 124.205 185.795 ;
        RECT 122.615 184.865 123.400 185.625 ;
        RECT 123.795 185.035 124.180 185.695 ;
        RECT 124.505 185.095 124.705 185.885 ;
        RECT 124.875 184.865 125.195 186.045 ;
        RECT 125.825 184.865 126.115 186.030 ;
        RECT 126.290 184.865 126.560 186.005 ;
        RECT 126.730 185.715 126.900 186.675 ;
        RECT 127.070 185.885 127.440 186.505 ;
        RECT 127.610 185.885 127.900 186.505 ;
        RECT 126.730 185.035 127.745 185.715 ;
        RECT 128.130 185.035 128.425 186.505 ;
        RECT 128.775 186.175 129.335 186.505 ;
        RECT 131.090 186.040 131.430 186.870 ;
        RECT 135.575 186.865 135.745 187.245 ;
        RECT 135.925 187.035 136.255 187.415 ;
        RECT 135.575 186.695 136.240 186.865 ;
        RECT 136.435 186.740 136.695 187.245 ;
        RECT 128.895 184.865 129.335 186.005 ;
        RECT 132.910 185.300 133.260 186.550 ;
        RECT 135.505 186.145 135.835 186.515 ;
        RECT 136.070 186.440 136.240 186.695 ;
        RECT 136.070 186.110 136.355 186.440 ;
        RECT 136.070 185.965 136.240 186.110 ;
        RECT 135.575 185.795 136.240 185.965 ;
        RECT 136.525 185.940 136.695 186.740 ;
        RECT 136.865 186.645 138.535 187.415 ;
        RECT 139.165 186.765 139.425 187.245 ;
        RECT 139.595 186.875 139.845 187.415 ;
        RECT 136.865 186.125 137.615 186.645 ;
        RECT 137.785 185.955 138.535 186.475 ;
        RECT 129.505 184.865 134.850 185.300 ;
        RECT 135.575 185.035 135.745 185.795 ;
        RECT 135.925 184.865 136.255 185.625 ;
        RECT 136.425 185.035 136.695 185.940 ;
        RECT 136.865 184.865 138.535 185.955 ;
        RECT 139.165 185.735 139.335 186.765 ;
        RECT 140.015 186.710 140.235 187.195 ;
        RECT 139.505 186.115 139.735 186.510 ;
        RECT 139.905 186.285 140.235 186.710 ;
        RECT 140.405 187.035 141.295 187.205 ;
        RECT 140.405 186.310 140.575 187.035 ;
        RECT 140.745 186.480 141.295 186.865 ;
        RECT 141.465 186.645 143.135 187.415 ;
        RECT 143.340 186.675 143.955 187.245 ;
        RECT 144.125 186.905 144.340 187.415 ;
        RECT 144.570 186.905 144.850 187.235 ;
        RECT 145.030 186.905 145.270 187.415 ;
        RECT 140.405 186.240 141.295 186.310 ;
        RECT 140.400 186.215 141.295 186.240 ;
        RECT 140.390 186.200 141.295 186.215 ;
        RECT 140.385 186.185 141.295 186.200 ;
        RECT 140.375 186.180 141.295 186.185 ;
        RECT 140.370 186.170 141.295 186.180 ;
        RECT 140.365 186.160 141.295 186.170 ;
        RECT 140.355 186.155 141.295 186.160 ;
        RECT 140.345 186.145 141.295 186.155 ;
        RECT 140.335 186.140 141.295 186.145 ;
        RECT 140.335 186.135 140.670 186.140 ;
        RECT 140.320 186.130 140.670 186.135 ;
        RECT 140.305 186.120 140.670 186.130 ;
        RECT 140.280 186.115 140.670 186.120 ;
        RECT 139.505 186.110 140.670 186.115 ;
        RECT 139.505 186.075 140.640 186.110 ;
        RECT 139.505 186.050 140.605 186.075 ;
        RECT 139.505 186.020 140.575 186.050 ;
        RECT 139.505 185.990 140.555 186.020 ;
        RECT 139.505 185.960 140.535 185.990 ;
        RECT 139.505 185.950 140.465 185.960 ;
        RECT 139.505 185.940 140.440 185.950 ;
        RECT 139.505 185.925 140.420 185.940 ;
        RECT 139.505 185.910 140.400 185.925 ;
        RECT 139.610 185.900 140.395 185.910 ;
        RECT 139.610 185.865 140.380 185.900 ;
        RECT 139.165 185.035 139.440 185.735 ;
        RECT 139.610 185.615 140.365 185.865 ;
        RECT 140.535 185.545 140.865 185.790 ;
        RECT 141.035 185.690 141.295 186.140 ;
        RECT 141.465 186.125 142.215 186.645 ;
        RECT 142.385 185.955 143.135 186.475 ;
        RECT 140.680 185.520 140.865 185.545 ;
        RECT 140.680 185.420 141.295 185.520 ;
        RECT 139.610 184.865 139.865 185.410 ;
        RECT 140.035 185.035 140.515 185.375 ;
        RECT 140.690 184.865 141.295 185.420 ;
        RECT 141.465 184.865 143.135 185.955 ;
        RECT 143.340 185.655 143.655 186.675 ;
        RECT 143.825 186.005 143.995 186.505 ;
        RECT 144.245 186.175 144.510 186.735 ;
        RECT 144.680 186.005 144.850 186.905 ;
        RECT 145.020 186.175 145.375 186.735 ;
        RECT 145.605 186.645 147.275 187.415 ;
        RECT 147.995 186.865 148.165 187.245 ;
        RECT 148.345 187.035 148.675 187.415 ;
        RECT 147.995 186.695 148.660 186.865 ;
        RECT 148.855 186.740 149.115 187.245 ;
        RECT 145.605 186.125 146.355 186.645 ;
        RECT 143.825 185.835 145.250 186.005 ;
        RECT 146.525 185.955 147.275 186.475 ;
        RECT 147.925 186.145 148.255 186.515 ;
        RECT 148.490 186.440 148.660 186.695 ;
        RECT 148.490 186.110 148.775 186.440 ;
        RECT 148.490 185.965 148.660 186.110 ;
        RECT 143.340 185.035 143.875 185.655 ;
        RECT 144.045 184.865 144.375 185.665 ;
        RECT 144.860 185.660 145.250 185.835 ;
        RECT 145.605 184.865 147.275 185.955 ;
        RECT 147.995 185.795 148.660 185.965 ;
        RECT 148.945 185.940 149.115 186.740 ;
        RECT 149.285 186.645 150.955 187.415 ;
        RECT 151.585 186.690 151.875 187.415 ;
        RECT 152.045 186.645 155.555 187.415 ;
        RECT 155.725 186.665 156.935 187.415 ;
        RECT 149.285 186.125 150.035 186.645 ;
        RECT 150.205 185.955 150.955 186.475 ;
        RECT 152.045 186.125 153.695 186.645 ;
        RECT 147.995 185.035 148.165 185.795 ;
        RECT 148.345 184.865 148.675 185.625 ;
        RECT 148.845 185.035 149.115 185.940 ;
        RECT 149.285 184.865 150.955 185.955 ;
        RECT 151.585 184.865 151.875 186.030 ;
        RECT 153.865 185.955 155.555 186.475 ;
        RECT 152.045 184.865 155.555 185.955 ;
        RECT 155.725 185.955 156.245 186.495 ;
        RECT 156.415 186.125 156.935 186.665 ;
        RECT 155.725 184.865 156.935 185.955 ;
        RECT 22.700 184.695 157.020 184.865 ;
        RECT 22.785 183.605 23.995 184.695 ;
        RECT 24.165 184.260 29.510 184.695 ;
        RECT 22.785 182.895 23.305 183.435 ;
        RECT 23.475 183.065 23.995 183.605 ;
        RECT 22.785 182.145 23.995 182.895 ;
        RECT 25.750 182.690 26.090 183.520 ;
        RECT 27.570 183.010 27.920 184.260 ;
        RECT 29.685 183.605 31.355 184.695 ;
        RECT 29.685 182.915 30.435 183.435 ;
        RECT 30.605 183.085 31.355 183.605 ;
        RECT 31.525 183.555 31.785 184.695 ;
        RECT 31.955 183.545 32.285 184.525 ;
        RECT 32.455 183.555 32.735 184.695 ;
        RECT 32.905 183.555 33.185 184.695 ;
        RECT 33.355 183.545 33.685 184.525 ;
        RECT 33.855 183.555 34.115 184.695 ;
        RECT 34.375 183.765 34.545 184.525 ;
        RECT 34.725 183.935 35.055 184.695 ;
        RECT 34.375 183.595 35.040 183.765 ;
        RECT 35.225 183.620 35.495 184.525 ;
        RECT 31.545 183.135 31.880 183.385 ;
        RECT 32.050 182.945 32.220 183.545 ;
        RECT 32.390 183.115 32.725 183.385 ;
        RECT 32.915 183.115 33.250 183.385 ;
        RECT 33.420 182.995 33.590 183.545 ;
        RECT 34.870 183.450 35.040 183.595 ;
        RECT 33.760 183.135 34.095 183.385 ;
        RECT 34.305 183.045 34.635 183.415 ;
        RECT 34.870 183.120 35.155 183.450 ;
        RECT 33.420 182.945 33.595 182.995 ;
        RECT 24.165 182.145 29.510 182.690 ;
        RECT 29.685 182.145 31.355 182.915 ;
        RECT 31.525 182.315 32.220 182.945 ;
        RECT 32.425 182.145 32.735 182.945 ;
        RECT 32.905 182.145 33.215 182.945 ;
        RECT 33.420 182.315 34.115 182.945 ;
        RECT 34.870 182.865 35.040 183.120 ;
        RECT 34.375 182.695 35.040 182.865 ;
        RECT 35.325 182.820 35.495 183.620 ;
        RECT 35.665 183.530 35.955 184.695 ;
        RECT 36.135 183.585 36.430 184.695 ;
        RECT 36.610 183.385 36.860 184.520 ;
        RECT 37.030 183.585 37.290 184.695 ;
        RECT 37.460 183.795 37.720 184.520 ;
        RECT 37.890 183.965 38.150 184.695 ;
        RECT 38.320 183.795 38.580 184.520 ;
        RECT 38.750 183.965 39.010 184.695 ;
        RECT 39.180 183.795 39.440 184.520 ;
        RECT 39.610 183.965 39.870 184.695 ;
        RECT 40.040 183.795 40.300 184.520 ;
        RECT 40.470 183.965 40.765 184.695 ;
        RECT 37.460 183.555 40.770 183.795 ;
        RECT 41.185 183.605 42.855 184.695 ;
        RECT 34.375 182.315 34.545 182.695 ;
        RECT 34.725 182.145 35.055 182.525 ;
        RECT 35.235 182.315 35.495 182.820 ;
        RECT 35.665 182.145 35.955 182.870 ;
        RECT 36.125 182.775 36.440 183.385 ;
        RECT 36.610 183.135 39.630 183.385 ;
        RECT 36.185 182.145 36.430 182.605 ;
        RECT 36.610 182.325 36.860 183.135 ;
        RECT 39.800 182.965 40.770 183.555 ;
        RECT 37.460 182.795 40.770 182.965 ;
        RECT 41.185 182.915 41.935 183.435 ;
        RECT 42.105 183.085 42.855 183.605 ;
        RECT 43.495 183.635 43.825 184.485 ;
        RECT 37.030 182.145 37.290 182.670 ;
        RECT 37.460 182.340 37.720 182.795 ;
        RECT 37.890 182.145 38.150 182.625 ;
        RECT 38.320 182.340 38.580 182.795 ;
        RECT 38.750 182.145 39.010 182.625 ;
        RECT 39.180 182.340 39.440 182.795 ;
        RECT 39.610 182.145 39.870 182.625 ;
        RECT 40.040 182.340 40.300 182.795 ;
        RECT 40.470 182.145 40.770 182.625 ;
        RECT 41.185 182.145 42.855 182.915 ;
        RECT 43.495 182.870 43.685 183.635 ;
        RECT 43.995 183.555 44.245 184.695 ;
        RECT 44.435 184.055 44.685 184.475 ;
        RECT 44.915 184.225 45.245 184.695 ;
        RECT 45.475 184.055 45.725 184.475 ;
        RECT 44.435 183.885 45.725 184.055 ;
        RECT 45.905 184.055 46.235 184.485 ;
        RECT 46.705 184.260 52.050 184.695 ;
        RECT 45.905 183.885 46.360 184.055 ;
        RECT 44.425 183.385 44.640 183.715 ;
        RECT 43.855 183.055 44.165 183.385 ;
        RECT 44.335 183.055 44.640 183.385 ;
        RECT 44.815 183.055 45.100 183.715 ;
        RECT 45.295 183.055 45.560 183.715 ;
        RECT 45.775 183.055 46.020 183.715 ;
        RECT 43.995 182.885 44.165 183.055 ;
        RECT 46.190 182.885 46.360 183.885 ;
        RECT 43.495 182.360 43.825 182.870 ;
        RECT 43.995 182.715 46.360 182.885 ;
        RECT 43.995 182.145 44.325 182.545 ;
        RECT 45.375 182.375 45.705 182.715 ;
        RECT 48.290 182.690 48.630 183.520 ;
        RECT 50.110 183.010 50.460 184.260 ;
        RECT 52.225 183.605 54.815 184.695 ;
        RECT 52.225 182.915 53.435 183.435 ;
        RECT 53.605 183.085 54.815 183.605 ;
        RECT 54.985 183.845 55.245 184.525 ;
        RECT 55.415 183.915 55.665 184.695 ;
        RECT 55.915 184.145 56.165 184.525 ;
        RECT 56.335 184.315 56.690 184.695 ;
        RECT 57.695 184.305 58.030 184.525 ;
        RECT 57.295 184.145 57.525 184.185 ;
        RECT 55.915 183.945 57.525 184.145 ;
        RECT 55.915 183.935 56.750 183.945 ;
        RECT 57.340 183.855 57.525 183.945 ;
        RECT 45.875 182.145 46.205 182.545 ;
        RECT 46.705 182.145 52.050 182.690 ;
        RECT 52.225 182.145 54.815 182.915 ;
        RECT 54.985 182.645 55.155 183.845 ;
        RECT 56.855 183.745 57.185 183.775 ;
        RECT 55.385 183.685 57.185 183.745 ;
        RECT 57.775 183.685 58.030 184.305 ;
        RECT 59.125 184.140 59.730 184.695 ;
        RECT 59.905 184.185 60.385 184.525 ;
        RECT 60.555 184.150 60.810 184.695 ;
        RECT 59.125 184.040 59.740 184.140 ;
        RECT 59.555 184.015 59.740 184.040 ;
        RECT 55.325 183.575 58.030 183.685 ;
        RECT 55.325 183.540 55.525 183.575 ;
        RECT 55.325 182.965 55.495 183.540 ;
        RECT 56.855 183.515 58.030 183.575 ;
        RECT 59.125 183.420 59.385 183.870 ;
        RECT 59.555 183.770 59.885 184.015 ;
        RECT 60.055 183.695 60.810 183.945 ;
        RECT 60.980 183.825 61.255 184.525 ;
        RECT 60.040 183.660 60.810 183.695 ;
        RECT 60.025 183.650 60.810 183.660 ;
        RECT 60.020 183.635 60.915 183.650 ;
        RECT 60.000 183.620 60.915 183.635 ;
        RECT 59.980 183.610 60.915 183.620 ;
        RECT 59.955 183.600 60.915 183.610 ;
        RECT 59.885 183.570 60.915 183.600 ;
        RECT 59.865 183.540 60.915 183.570 ;
        RECT 59.845 183.510 60.915 183.540 ;
        RECT 59.815 183.485 60.915 183.510 ;
        RECT 59.780 183.450 60.915 183.485 ;
        RECT 59.750 183.445 60.915 183.450 ;
        RECT 59.750 183.440 60.140 183.445 ;
        RECT 59.750 183.430 60.115 183.440 ;
        RECT 59.750 183.425 60.100 183.430 ;
        RECT 59.750 183.420 60.085 183.425 ;
        RECT 59.125 183.415 60.085 183.420 ;
        RECT 59.125 183.405 60.075 183.415 ;
        RECT 55.725 183.100 56.135 183.405 ;
        RECT 59.125 183.400 60.065 183.405 ;
        RECT 59.125 183.390 60.055 183.400 ;
        RECT 59.125 183.380 60.050 183.390 ;
        RECT 59.125 183.375 60.045 183.380 ;
        RECT 59.125 183.360 60.035 183.375 ;
        RECT 59.125 183.345 60.030 183.360 ;
        RECT 56.305 183.135 56.635 183.345 ;
        RECT 55.325 182.845 55.595 182.965 ;
        RECT 55.325 182.800 56.170 182.845 ;
        RECT 55.415 182.675 56.170 182.800 ;
        RECT 56.425 182.735 56.635 183.135 ;
        RECT 56.880 183.135 57.355 183.345 ;
        RECT 57.545 183.135 58.035 183.335 ;
        RECT 59.125 183.320 60.020 183.345 ;
        RECT 59.125 183.250 60.015 183.320 ;
        RECT 56.880 182.735 57.100 183.135 ;
        RECT 54.985 182.315 55.245 182.645 ;
        RECT 56.000 182.525 56.170 182.675 ;
        RECT 55.415 182.145 55.745 182.505 ;
        RECT 56.000 182.315 57.300 182.525 ;
        RECT 57.575 182.145 58.030 182.910 ;
        RECT 59.125 182.695 59.675 183.080 ;
        RECT 59.845 182.525 60.015 183.250 ;
        RECT 59.125 182.355 60.015 182.525 ;
        RECT 60.185 182.850 60.515 183.275 ;
        RECT 60.685 183.050 60.915 183.445 ;
        RECT 60.185 182.365 60.405 182.850 ;
        RECT 61.085 182.795 61.255 183.825 ;
        RECT 61.425 183.530 61.715 184.695 ;
        RECT 61.975 184.025 62.145 184.525 ;
        RECT 62.315 184.195 62.645 184.695 ;
        RECT 61.975 183.855 62.640 184.025 ;
        RECT 61.890 183.035 62.240 183.685 ;
        RECT 60.575 182.145 60.825 182.685 ;
        RECT 60.995 182.315 61.255 182.795 ;
        RECT 61.425 182.145 61.715 182.870 ;
        RECT 62.410 182.865 62.640 183.855 ;
        RECT 61.975 182.695 62.640 182.865 ;
        RECT 61.975 182.405 62.145 182.695 ;
        RECT 62.315 182.145 62.645 182.525 ;
        RECT 62.815 182.405 63.000 184.525 ;
        RECT 63.240 184.235 63.505 184.695 ;
        RECT 63.675 184.100 63.925 184.525 ;
        RECT 64.135 184.250 65.240 184.420 ;
        RECT 63.620 183.970 63.925 184.100 ;
        RECT 63.170 182.775 63.450 183.725 ;
        RECT 63.620 182.865 63.790 183.970 ;
        RECT 63.960 183.185 64.200 183.780 ;
        RECT 64.370 183.715 64.900 184.080 ;
        RECT 64.370 183.015 64.540 183.715 ;
        RECT 65.070 183.635 65.240 184.250 ;
        RECT 65.410 183.895 65.580 184.695 ;
        RECT 65.750 184.195 66.000 184.525 ;
        RECT 66.225 184.225 67.110 184.395 ;
        RECT 65.070 183.545 65.580 183.635 ;
        RECT 63.620 182.735 63.845 182.865 ;
        RECT 64.015 182.795 64.540 183.015 ;
        RECT 64.710 183.375 65.580 183.545 ;
        RECT 63.255 182.145 63.505 182.605 ;
        RECT 63.675 182.595 63.845 182.735 ;
        RECT 64.710 182.595 64.880 183.375 ;
        RECT 65.410 183.305 65.580 183.375 ;
        RECT 65.090 183.125 65.290 183.155 ;
        RECT 65.750 183.125 65.920 184.195 ;
        RECT 66.090 183.305 66.280 184.025 ;
        RECT 65.090 182.825 65.920 183.125 ;
        RECT 66.450 183.095 66.770 184.055 ;
        RECT 63.675 182.425 64.010 182.595 ;
        RECT 64.205 182.425 64.880 182.595 ;
        RECT 65.200 182.145 65.570 182.645 ;
        RECT 65.750 182.595 65.920 182.825 ;
        RECT 66.305 182.765 66.770 183.095 ;
        RECT 66.940 183.385 67.110 184.225 ;
        RECT 67.290 184.195 67.605 184.695 ;
        RECT 67.835 183.965 68.175 184.525 ;
        RECT 67.280 183.590 68.175 183.965 ;
        RECT 68.345 183.685 68.515 184.695 ;
        RECT 67.985 183.385 68.175 183.590 ;
        RECT 68.685 183.635 69.015 184.480 ;
        RECT 68.685 183.555 69.075 183.635 ;
        RECT 68.860 183.505 69.075 183.555 ;
        RECT 66.940 183.055 67.815 183.385 ;
        RECT 67.985 183.055 68.735 183.385 ;
        RECT 66.940 182.595 67.110 183.055 ;
        RECT 67.985 182.885 68.185 183.055 ;
        RECT 68.905 182.925 69.075 183.505 ;
        RECT 68.850 182.885 69.075 182.925 ;
        RECT 65.750 182.425 66.155 182.595 ;
        RECT 66.325 182.425 67.110 182.595 ;
        RECT 67.385 182.145 67.595 182.675 ;
        RECT 67.855 182.360 68.185 182.885 ;
        RECT 68.695 182.800 69.075 182.885 ;
        RECT 68.355 182.145 68.525 182.755 ;
        RECT 68.695 182.365 69.025 182.800 ;
        RECT 69.705 182.425 69.985 184.525 ;
        RECT 70.175 183.935 70.960 184.695 ;
        RECT 71.355 183.865 71.740 184.525 ;
        RECT 71.355 183.765 71.765 183.865 ;
        RECT 70.155 183.555 71.765 183.765 ;
        RECT 72.065 183.675 72.265 184.465 ;
        RECT 70.155 182.955 70.430 183.555 ;
        RECT 71.935 183.505 72.265 183.675 ;
        RECT 72.435 183.515 72.755 184.695 ;
        RECT 72.925 183.605 74.135 184.695 ;
        RECT 71.935 183.385 72.115 183.505 ;
        RECT 70.600 183.135 70.955 183.385 ;
        RECT 71.150 183.335 71.615 183.385 ;
        RECT 71.145 183.165 71.615 183.335 ;
        RECT 71.150 183.135 71.615 183.165 ;
        RECT 71.785 183.135 72.115 183.385 ;
        RECT 72.290 183.135 72.755 183.335 ;
        RECT 70.155 182.775 71.405 182.955 ;
        RECT 71.040 182.705 71.405 182.775 ;
        RECT 71.575 182.755 72.755 182.925 ;
        RECT 70.215 182.145 70.385 182.605 ;
        RECT 71.575 182.535 71.905 182.755 ;
        RECT 70.655 182.355 71.905 182.535 ;
        RECT 72.075 182.145 72.245 182.585 ;
        RECT 72.415 182.340 72.755 182.755 ;
        RECT 72.925 182.895 73.445 183.435 ;
        RECT 73.615 183.065 74.135 183.605 ;
        RECT 74.315 183.585 74.610 184.695 ;
        RECT 74.790 183.385 75.040 184.520 ;
        RECT 75.210 183.585 75.470 184.695 ;
        RECT 75.640 183.795 75.900 184.520 ;
        RECT 76.070 183.965 76.330 184.695 ;
        RECT 76.500 183.795 76.760 184.520 ;
        RECT 76.930 183.965 77.190 184.695 ;
        RECT 77.360 183.795 77.620 184.520 ;
        RECT 77.790 183.965 78.050 184.695 ;
        RECT 78.220 183.795 78.480 184.520 ;
        RECT 78.650 183.965 78.945 184.695 ;
        RECT 75.640 183.555 78.950 183.795 ;
        RECT 72.925 182.145 74.135 182.895 ;
        RECT 74.305 182.775 74.620 183.385 ;
        RECT 74.790 183.135 77.810 183.385 ;
        RECT 74.365 182.145 74.610 182.605 ;
        RECT 74.790 182.325 75.040 183.135 ;
        RECT 77.980 182.965 78.950 183.555 ;
        RECT 75.640 182.795 78.950 182.965 ;
        RECT 79.365 183.555 79.750 184.525 ;
        RECT 79.920 184.235 80.245 184.695 ;
        RECT 80.765 184.065 81.045 184.525 ;
        RECT 79.920 183.845 81.045 184.065 ;
        RECT 79.365 182.885 79.645 183.555 ;
        RECT 79.920 183.385 80.370 183.845 ;
        RECT 81.235 183.675 81.635 184.525 ;
        RECT 82.035 184.235 82.305 184.695 ;
        RECT 82.475 184.065 82.760 184.525 ;
        RECT 79.815 183.055 80.370 183.385 ;
        RECT 80.540 183.115 81.635 183.675 ;
        RECT 79.920 182.945 80.370 183.055 ;
        RECT 75.210 182.145 75.470 182.670 ;
        RECT 75.640 182.340 75.900 182.795 ;
        RECT 76.070 182.145 76.330 182.625 ;
        RECT 76.500 182.340 76.760 182.795 ;
        RECT 76.930 182.145 77.190 182.625 ;
        RECT 77.360 182.340 77.620 182.795 ;
        RECT 77.790 182.145 78.050 182.625 ;
        RECT 78.220 182.340 78.480 182.795 ;
        RECT 78.650 182.145 78.950 182.625 ;
        RECT 79.365 182.315 79.750 182.885 ;
        RECT 79.920 182.775 81.045 182.945 ;
        RECT 79.920 182.145 80.245 182.605 ;
        RECT 80.765 182.315 81.045 182.775 ;
        RECT 81.235 182.315 81.635 183.115 ;
        RECT 81.805 183.845 82.760 184.065 ;
        RECT 83.620 184.065 83.905 184.525 ;
        RECT 84.075 184.235 84.345 184.695 ;
        RECT 83.620 183.845 84.575 184.065 ;
        RECT 81.805 182.945 82.015 183.845 ;
        RECT 82.185 183.115 82.875 183.675 ;
        RECT 83.505 183.115 84.195 183.675 ;
        RECT 84.365 182.945 84.575 183.845 ;
        RECT 81.805 182.775 82.760 182.945 ;
        RECT 82.035 182.145 82.305 182.605 ;
        RECT 82.475 182.315 82.760 182.775 ;
        RECT 83.620 182.775 84.575 182.945 ;
        RECT 84.745 183.675 85.145 184.525 ;
        RECT 85.335 184.065 85.615 184.525 ;
        RECT 86.135 184.235 86.460 184.695 ;
        RECT 85.335 183.845 86.460 184.065 ;
        RECT 84.745 183.115 85.840 183.675 ;
        RECT 86.010 183.385 86.460 183.845 ;
        RECT 86.630 183.555 87.015 184.525 ;
        RECT 83.620 182.315 83.905 182.775 ;
        RECT 84.075 182.145 84.345 182.605 ;
        RECT 84.745 182.315 85.145 183.115 ;
        RECT 86.010 183.055 86.565 183.385 ;
        RECT 86.010 182.945 86.460 183.055 ;
        RECT 85.335 182.775 86.460 182.945 ;
        RECT 86.735 182.885 87.015 183.555 ;
        RECT 87.185 183.530 87.475 184.695 ;
        RECT 87.735 184.025 87.905 184.525 ;
        RECT 88.075 184.195 88.405 184.695 ;
        RECT 87.735 183.855 88.400 184.025 ;
        RECT 87.650 183.035 88.000 183.685 ;
        RECT 85.335 182.315 85.615 182.775 ;
        RECT 86.135 182.145 86.460 182.605 ;
        RECT 86.630 182.315 87.015 182.885 ;
        RECT 87.185 182.145 87.475 182.870 ;
        RECT 88.170 182.865 88.400 183.855 ;
        RECT 87.735 182.695 88.400 182.865 ;
        RECT 87.735 182.405 87.905 182.695 ;
        RECT 88.075 182.145 88.405 182.525 ;
        RECT 88.575 182.405 88.760 184.525 ;
        RECT 89.000 184.235 89.265 184.695 ;
        RECT 89.435 184.100 89.685 184.525 ;
        RECT 89.895 184.250 91.000 184.420 ;
        RECT 89.380 183.970 89.685 184.100 ;
        RECT 88.930 182.775 89.210 183.725 ;
        RECT 89.380 182.865 89.550 183.970 ;
        RECT 89.720 183.185 89.960 183.780 ;
        RECT 90.130 183.715 90.660 184.080 ;
        RECT 90.130 183.015 90.300 183.715 ;
        RECT 90.830 183.635 91.000 184.250 ;
        RECT 91.170 183.895 91.340 184.695 ;
        RECT 91.510 184.195 91.760 184.525 ;
        RECT 91.985 184.225 92.870 184.395 ;
        RECT 90.830 183.545 91.340 183.635 ;
        RECT 89.380 182.735 89.605 182.865 ;
        RECT 89.775 182.795 90.300 183.015 ;
        RECT 90.470 183.375 91.340 183.545 ;
        RECT 89.015 182.145 89.265 182.605 ;
        RECT 89.435 182.595 89.605 182.735 ;
        RECT 90.470 182.595 90.640 183.375 ;
        RECT 91.170 183.305 91.340 183.375 ;
        RECT 90.850 183.125 91.050 183.155 ;
        RECT 91.510 183.125 91.680 184.195 ;
        RECT 91.850 183.305 92.040 184.025 ;
        RECT 90.850 182.825 91.680 183.125 ;
        RECT 92.210 183.095 92.530 184.055 ;
        RECT 89.435 182.425 89.770 182.595 ;
        RECT 89.965 182.425 90.640 182.595 ;
        RECT 90.960 182.145 91.330 182.645 ;
        RECT 91.510 182.595 91.680 182.825 ;
        RECT 92.065 182.765 92.530 183.095 ;
        RECT 92.700 183.385 92.870 184.225 ;
        RECT 93.050 184.195 93.365 184.695 ;
        RECT 93.595 183.965 93.935 184.525 ;
        RECT 93.040 183.590 93.935 183.965 ;
        RECT 94.105 183.685 94.275 184.695 ;
        RECT 93.745 183.385 93.935 183.590 ;
        RECT 94.445 183.635 94.775 184.480 ;
        RECT 95.005 183.975 95.465 184.525 ;
        RECT 95.655 183.975 95.985 184.695 ;
        RECT 94.445 183.555 94.835 183.635 ;
        RECT 94.620 183.505 94.835 183.555 ;
        RECT 92.700 183.055 93.575 183.385 ;
        RECT 93.745 183.055 94.495 183.385 ;
        RECT 92.700 182.595 92.870 183.055 ;
        RECT 93.745 182.885 93.945 183.055 ;
        RECT 94.665 182.925 94.835 183.505 ;
        RECT 94.610 182.885 94.835 182.925 ;
        RECT 91.510 182.425 91.915 182.595 ;
        RECT 92.085 182.425 92.870 182.595 ;
        RECT 93.145 182.145 93.355 182.675 ;
        RECT 93.615 182.360 93.945 182.885 ;
        RECT 94.455 182.800 94.835 182.885 ;
        RECT 94.115 182.145 94.285 182.755 ;
        RECT 94.455 182.365 94.785 182.800 ;
        RECT 95.005 182.605 95.255 183.975 ;
        RECT 96.185 183.805 96.485 184.355 ;
        RECT 96.655 184.025 96.935 184.695 ;
        RECT 97.505 184.025 97.785 184.695 ;
        RECT 95.545 183.635 96.485 183.805 ;
        RECT 97.955 183.805 98.255 184.355 ;
        RECT 98.455 183.975 98.785 184.695 ;
        RECT 98.975 183.975 99.435 184.525 ;
        RECT 95.545 183.385 95.715 183.635 ;
        RECT 96.855 183.385 97.120 183.745 ;
        RECT 95.425 183.055 95.715 183.385 ;
        RECT 95.885 183.135 96.225 183.385 ;
        RECT 96.445 183.135 97.120 183.385 ;
        RECT 97.320 183.385 97.585 183.745 ;
        RECT 97.955 183.635 98.895 183.805 ;
        RECT 98.725 183.385 98.895 183.635 ;
        RECT 97.320 183.135 97.995 183.385 ;
        RECT 98.215 183.135 98.555 183.385 ;
        RECT 95.545 182.965 95.715 183.055 ;
        RECT 98.725 183.055 99.015 183.385 ;
        RECT 98.725 182.965 98.895 183.055 ;
        RECT 95.545 182.775 96.935 182.965 ;
        RECT 95.005 182.315 95.565 182.605 ;
        RECT 95.735 182.145 95.985 182.605 ;
        RECT 96.605 182.415 96.935 182.775 ;
        RECT 97.505 182.775 98.895 182.965 ;
        RECT 97.505 182.415 97.835 182.775 ;
        RECT 99.185 182.605 99.435 183.975 ;
        RECT 99.605 183.605 101.275 184.695 ;
        RECT 98.455 182.145 98.705 182.605 ;
        RECT 98.875 182.315 99.435 182.605 ;
        RECT 99.605 182.915 100.355 183.435 ;
        RECT 100.525 183.085 101.275 183.605 ;
        RECT 101.905 183.975 102.365 184.525 ;
        RECT 102.555 183.975 102.885 184.695 ;
        RECT 99.605 182.145 101.275 182.915 ;
        RECT 101.905 182.605 102.155 183.975 ;
        RECT 103.085 183.805 103.385 184.355 ;
        RECT 103.555 184.025 103.835 184.695 ;
        RECT 102.445 183.635 103.385 183.805 ;
        RECT 102.445 183.385 102.615 183.635 ;
        RECT 103.755 183.385 104.020 183.745 ;
        RECT 104.205 183.605 107.715 184.695 ;
        RECT 102.325 183.055 102.615 183.385 ;
        RECT 102.785 183.135 103.125 183.385 ;
        RECT 103.345 183.135 104.020 183.385 ;
        RECT 102.445 182.965 102.615 183.055 ;
        RECT 102.445 182.775 103.835 182.965 ;
        RECT 101.905 182.315 102.465 182.605 ;
        RECT 102.635 182.145 102.885 182.605 ;
        RECT 103.505 182.415 103.835 182.775 ;
        RECT 104.205 182.915 105.855 183.435 ;
        RECT 106.025 183.085 107.715 183.605 ;
        RECT 108.345 183.845 108.605 184.525 ;
        RECT 108.775 183.915 109.025 184.695 ;
        RECT 109.275 184.145 109.525 184.525 ;
        RECT 109.695 184.315 110.050 184.695 ;
        RECT 111.055 184.305 111.390 184.525 ;
        RECT 110.655 184.145 110.885 184.185 ;
        RECT 109.275 183.945 110.885 184.145 ;
        RECT 109.275 183.935 110.110 183.945 ;
        RECT 110.700 183.855 110.885 183.945 ;
        RECT 104.205 182.145 107.715 182.915 ;
        RECT 108.345 182.655 108.515 183.845 ;
        RECT 110.215 183.745 110.545 183.775 ;
        RECT 108.745 183.685 110.545 183.745 ;
        RECT 111.135 183.685 111.390 184.305 ;
        RECT 108.685 183.575 111.390 183.685 ;
        RECT 111.565 183.605 112.775 184.695 ;
        RECT 108.685 183.540 108.885 183.575 ;
        RECT 108.685 182.965 108.855 183.540 ;
        RECT 110.215 183.515 111.390 183.575 ;
        RECT 109.085 183.100 109.495 183.405 ;
        RECT 109.665 183.135 109.995 183.345 ;
        RECT 108.685 182.845 108.955 182.965 ;
        RECT 108.685 182.800 109.530 182.845 ;
        RECT 108.775 182.675 109.530 182.800 ;
        RECT 109.785 182.735 109.995 183.135 ;
        RECT 110.240 183.135 110.715 183.345 ;
        RECT 110.905 183.135 111.395 183.335 ;
        RECT 110.240 182.735 110.460 183.135 ;
        RECT 108.345 182.645 108.575 182.655 ;
        RECT 108.345 182.315 108.605 182.645 ;
        RECT 109.360 182.525 109.530 182.675 ;
        RECT 108.775 182.145 109.105 182.505 ;
        RECT 109.360 182.315 110.660 182.525 ;
        RECT 110.935 182.145 111.390 182.910 ;
        RECT 111.565 182.895 112.085 183.435 ;
        RECT 112.255 183.065 112.775 183.605 ;
        RECT 112.945 183.530 113.235 184.695 ;
        RECT 113.495 184.025 113.665 184.525 ;
        RECT 113.835 184.195 114.165 184.695 ;
        RECT 113.495 183.855 114.160 184.025 ;
        RECT 113.410 183.035 113.760 183.685 ;
        RECT 111.565 182.145 112.775 182.895 ;
        RECT 112.945 182.145 113.235 182.870 ;
        RECT 113.930 182.865 114.160 183.855 ;
        RECT 113.495 182.695 114.160 182.865 ;
        RECT 113.495 182.405 113.665 182.695 ;
        RECT 113.835 182.145 114.165 182.525 ;
        RECT 114.335 182.405 114.520 184.525 ;
        RECT 114.760 184.235 115.025 184.695 ;
        RECT 115.195 184.100 115.445 184.525 ;
        RECT 115.655 184.250 116.760 184.420 ;
        RECT 115.140 183.970 115.445 184.100 ;
        RECT 114.690 182.775 114.970 183.725 ;
        RECT 115.140 182.865 115.310 183.970 ;
        RECT 115.480 183.185 115.720 183.780 ;
        RECT 115.890 183.715 116.420 184.080 ;
        RECT 115.890 183.015 116.060 183.715 ;
        RECT 116.590 183.635 116.760 184.250 ;
        RECT 116.930 183.895 117.100 184.695 ;
        RECT 117.270 184.195 117.520 184.525 ;
        RECT 117.745 184.225 118.630 184.395 ;
        RECT 116.590 183.545 117.100 183.635 ;
        RECT 115.140 182.735 115.365 182.865 ;
        RECT 115.535 182.795 116.060 183.015 ;
        RECT 116.230 183.375 117.100 183.545 ;
        RECT 114.775 182.145 115.025 182.605 ;
        RECT 115.195 182.595 115.365 182.735 ;
        RECT 116.230 182.595 116.400 183.375 ;
        RECT 116.930 183.305 117.100 183.375 ;
        RECT 116.610 183.125 116.810 183.155 ;
        RECT 117.270 183.125 117.440 184.195 ;
        RECT 117.610 183.305 117.800 184.025 ;
        RECT 116.610 182.825 117.440 183.125 ;
        RECT 117.970 183.095 118.290 184.055 ;
        RECT 115.195 182.425 115.530 182.595 ;
        RECT 115.725 182.425 116.400 182.595 ;
        RECT 116.720 182.145 117.090 182.645 ;
        RECT 117.270 182.595 117.440 182.825 ;
        RECT 117.825 182.765 118.290 183.095 ;
        RECT 118.460 183.385 118.630 184.225 ;
        RECT 118.810 184.195 119.125 184.695 ;
        RECT 119.355 183.965 119.695 184.525 ;
        RECT 118.800 183.590 119.695 183.965 ;
        RECT 119.865 183.685 120.035 184.695 ;
        RECT 119.505 183.385 119.695 183.590 ;
        RECT 120.205 183.635 120.535 184.480 ;
        RECT 120.775 184.085 121.105 184.515 ;
        RECT 121.285 184.255 121.480 184.695 ;
        RECT 121.650 184.085 121.980 184.515 ;
        RECT 120.775 183.915 121.980 184.085 ;
        RECT 120.205 183.555 120.595 183.635 ;
        RECT 120.775 183.585 121.670 183.915 ;
        RECT 122.150 183.745 122.425 184.515 ;
        RECT 120.380 183.505 120.595 183.555 ;
        RECT 118.460 183.055 119.335 183.385 ;
        RECT 119.505 183.055 120.255 183.385 ;
        RECT 118.460 182.595 118.630 183.055 ;
        RECT 119.505 182.885 119.705 183.055 ;
        RECT 120.425 182.925 120.595 183.505 ;
        RECT 121.840 183.555 122.425 183.745 ;
        RECT 123.525 183.975 123.985 184.525 ;
        RECT 124.175 183.975 124.505 184.695 ;
        RECT 120.780 183.055 121.075 183.385 ;
        RECT 121.255 183.055 121.670 183.385 ;
        RECT 120.370 182.885 120.595 182.925 ;
        RECT 117.270 182.425 117.675 182.595 ;
        RECT 117.845 182.425 118.630 182.595 ;
        RECT 118.905 182.145 119.115 182.675 ;
        RECT 119.375 182.360 119.705 182.885 ;
        RECT 120.215 182.800 120.595 182.885 ;
        RECT 119.875 182.145 120.045 182.755 ;
        RECT 120.215 182.365 120.545 182.800 ;
        RECT 120.775 182.145 121.075 182.875 ;
        RECT 121.255 182.435 121.485 183.055 ;
        RECT 121.840 182.885 122.015 183.555 ;
        RECT 121.685 182.705 122.015 182.885 ;
        RECT 122.185 182.735 122.425 183.385 ;
        RECT 121.685 182.325 121.910 182.705 ;
        RECT 123.525 182.605 123.775 183.975 ;
        RECT 124.705 183.805 125.005 184.355 ;
        RECT 125.175 184.025 125.455 184.695 ;
        RECT 124.065 183.635 125.005 183.805 ;
        RECT 124.065 183.385 124.235 183.635 ;
        RECT 125.375 183.385 125.640 183.745 ;
        RECT 125.865 183.555 126.095 184.695 ;
        RECT 126.265 183.545 126.595 184.525 ;
        RECT 126.765 183.555 126.975 184.695 ;
        RECT 127.205 183.605 130.715 184.695 ;
        RECT 131.405 183.635 131.735 184.480 ;
        RECT 131.905 183.685 132.075 184.695 ;
        RECT 132.245 183.965 132.585 184.525 ;
        RECT 132.815 184.195 133.130 184.695 ;
        RECT 133.310 184.225 134.195 184.395 ;
        RECT 123.945 183.055 124.235 183.385 ;
        RECT 124.405 183.135 124.745 183.385 ;
        RECT 124.965 183.135 125.640 183.385 ;
        RECT 125.845 183.135 126.175 183.385 ;
        RECT 124.065 182.965 124.235 183.055 ;
        RECT 124.065 182.775 125.455 182.965 ;
        RECT 122.080 182.145 122.410 182.535 ;
        RECT 123.525 182.315 124.085 182.605 ;
        RECT 124.255 182.145 124.505 182.605 ;
        RECT 125.125 182.415 125.455 182.775 ;
        RECT 125.865 182.145 126.095 182.965 ;
        RECT 126.345 182.945 126.595 183.545 ;
        RECT 126.265 182.315 126.595 182.945 ;
        RECT 126.765 182.145 126.975 182.965 ;
        RECT 127.205 182.915 128.855 183.435 ;
        RECT 129.025 183.085 130.715 183.605 ;
        RECT 131.345 183.555 131.735 183.635 ;
        RECT 132.245 183.590 133.140 183.965 ;
        RECT 131.345 183.505 131.560 183.555 ;
        RECT 131.345 182.925 131.515 183.505 ;
        RECT 132.245 183.385 132.435 183.590 ;
        RECT 133.310 183.385 133.480 184.225 ;
        RECT 134.420 184.195 134.670 184.525 ;
        RECT 131.685 183.055 132.435 183.385 ;
        RECT 132.605 183.055 133.480 183.385 ;
        RECT 127.205 182.145 130.715 182.915 ;
        RECT 131.345 182.885 131.570 182.925 ;
        RECT 132.235 182.885 132.435 183.055 ;
        RECT 131.345 182.800 131.725 182.885 ;
        RECT 131.395 182.365 131.725 182.800 ;
        RECT 131.895 182.145 132.065 182.755 ;
        RECT 132.235 182.360 132.565 182.885 ;
        RECT 132.825 182.145 133.035 182.675 ;
        RECT 133.310 182.595 133.480 183.055 ;
        RECT 133.650 183.095 133.970 184.055 ;
        RECT 134.140 183.305 134.330 184.025 ;
        RECT 134.500 183.125 134.670 184.195 ;
        RECT 134.840 183.895 135.010 184.695 ;
        RECT 135.180 184.250 136.285 184.420 ;
        RECT 135.180 183.635 135.350 184.250 ;
        RECT 136.495 184.100 136.745 184.525 ;
        RECT 136.915 184.235 137.180 184.695 ;
        RECT 135.520 183.715 136.050 184.080 ;
        RECT 136.495 183.970 136.800 184.100 ;
        RECT 134.840 183.545 135.350 183.635 ;
        RECT 134.840 183.375 135.710 183.545 ;
        RECT 134.840 183.305 135.010 183.375 ;
        RECT 135.130 183.125 135.330 183.155 ;
        RECT 133.650 182.765 134.115 183.095 ;
        RECT 134.500 182.825 135.330 183.125 ;
        RECT 134.500 182.595 134.670 182.825 ;
        RECT 133.310 182.425 134.095 182.595 ;
        RECT 134.265 182.425 134.670 182.595 ;
        RECT 134.850 182.145 135.220 182.645 ;
        RECT 135.540 182.595 135.710 183.375 ;
        RECT 135.880 183.015 136.050 183.715 ;
        RECT 136.220 183.185 136.460 183.780 ;
        RECT 135.880 182.795 136.405 183.015 ;
        RECT 136.630 182.865 136.800 183.970 ;
        RECT 136.575 182.735 136.800 182.865 ;
        RECT 136.970 182.775 137.250 183.725 ;
        RECT 136.575 182.595 136.745 182.735 ;
        RECT 135.540 182.425 136.215 182.595 ;
        RECT 136.410 182.425 136.745 182.595 ;
        RECT 136.915 182.145 137.165 182.605 ;
        RECT 137.420 182.405 137.605 184.525 ;
        RECT 137.775 184.195 138.105 184.695 ;
        RECT 138.275 184.025 138.445 184.525 ;
        RECT 137.780 183.855 138.445 184.025 ;
        RECT 137.780 182.865 138.010 183.855 ;
        RECT 138.180 183.035 138.530 183.685 ;
        RECT 138.705 183.530 138.995 184.695 ;
        RECT 139.165 183.825 139.440 184.525 ;
        RECT 139.610 184.150 139.865 184.695 ;
        RECT 140.035 184.185 140.515 184.525 ;
        RECT 140.690 184.140 141.295 184.695 ;
        RECT 141.465 184.185 141.725 184.695 ;
        RECT 140.680 184.040 141.295 184.140 ;
        RECT 140.680 184.015 140.865 184.040 ;
        RECT 137.780 182.695 138.445 182.865 ;
        RECT 137.775 182.145 138.105 182.525 ;
        RECT 138.275 182.405 138.445 182.695 ;
        RECT 138.705 182.145 138.995 182.870 ;
        RECT 139.165 182.795 139.335 183.825 ;
        RECT 139.610 183.695 140.365 183.945 ;
        RECT 140.535 183.770 140.865 184.015 ;
        RECT 139.610 183.660 140.380 183.695 ;
        RECT 139.610 183.650 140.395 183.660 ;
        RECT 139.505 183.635 140.400 183.650 ;
        RECT 139.505 183.620 140.420 183.635 ;
        RECT 139.505 183.610 140.440 183.620 ;
        RECT 139.505 183.600 140.465 183.610 ;
        RECT 139.505 183.570 140.535 183.600 ;
        RECT 139.505 183.540 140.555 183.570 ;
        RECT 139.505 183.510 140.575 183.540 ;
        RECT 139.505 183.485 140.605 183.510 ;
        RECT 139.505 183.450 140.640 183.485 ;
        RECT 139.505 183.445 140.670 183.450 ;
        RECT 139.505 183.050 139.735 183.445 ;
        RECT 140.280 183.440 140.670 183.445 ;
        RECT 140.305 183.430 140.670 183.440 ;
        RECT 140.320 183.425 140.670 183.430 ;
        RECT 140.335 183.420 140.670 183.425 ;
        RECT 141.035 183.420 141.295 183.870 ;
        RECT 140.335 183.415 141.295 183.420 ;
        RECT 140.345 183.405 141.295 183.415 ;
        RECT 140.355 183.400 141.295 183.405 ;
        RECT 140.365 183.390 141.295 183.400 ;
        RECT 140.370 183.380 141.295 183.390 ;
        RECT 140.375 183.375 141.295 183.380 ;
        RECT 140.385 183.360 141.295 183.375 ;
        RECT 140.390 183.345 141.295 183.360 ;
        RECT 140.400 183.320 141.295 183.345 ;
        RECT 139.905 182.850 140.235 183.275 ;
        RECT 139.165 182.315 139.425 182.795 ;
        RECT 139.595 182.145 139.845 182.685 ;
        RECT 140.015 182.365 140.235 182.850 ;
        RECT 140.405 183.250 141.295 183.320 ;
        RECT 140.405 182.525 140.575 183.250 ;
        RECT 141.465 183.135 141.805 184.015 ;
        RECT 141.975 183.305 142.145 184.525 ;
        RECT 142.385 184.190 143.000 184.695 ;
        RECT 142.385 183.655 142.635 184.020 ;
        RECT 142.805 184.015 143.000 184.190 ;
        RECT 143.170 184.185 143.645 184.525 ;
        RECT 143.815 184.150 144.030 184.695 ;
        RECT 142.805 183.825 143.135 184.015 ;
        RECT 143.355 183.655 144.070 183.950 ;
        RECT 144.240 183.825 144.515 184.525 ;
        RECT 142.385 183.485 144.175 183.655 ;
        RECT 140.745 182.695 141.295 183.080 ;
        RECT 141.975 183.055 142.770 183.305 ;
        RECT 141.975 182.965 142.225 183.055 ;
        RECT 140.405 182.355 141.295 182.525 ;
        RECT 141.465 182.145 141.725 182.965 ;
        RECT 141.895 182.545 142.225 182.965 ;
        RECT 142.940 182.630 143.195 183.485 ;
        RECT 142.405 182.365 143.195 182.630 ;
        RECT 143.365 182.785 143.775 183.305 ;
        RECT 143.945 183.055 144.175 183.485 ;
        RECT 144.345 182.795 144.515 183.825 ;
        RECT 144.745 183.635 145.075 184.480 ;
        RECT 145.245 183.685 145.415 184.695 ;
        RECT 145.585 183.965 145.925 184.525 ;
        RECT 146.155 184.195 146.470 184.695 ;
        RECT 146.650 184.225 147.535 184.395 ;
        RECT 144.685 183.555 145.075 183.635 ;
        RECT 145.585 183.590 146.480 183.965 ;
        RECT 144.685 183.505 144.900 183.555 ;
        RECT 144.685 182.925 144.855 183.505 ;
        RECT 145.585 183.385 145.775 183.590 ;
        RECT 146.650 183.385 146.820 184.225 ;
        RECT 147.760 184.195 148.010 184.525 ;
        RECT 145.025 183.055 145.775 183.385 ;
        RECT 145.945 183.055 146.820 183.385 ;
        RECT 144.685 182.885 144.910 182.925 ;
        RECT 145.575 182.885 145.775 183.055 ;
        RECT 144.685 182.800 145.065 182.885 ;
        RECT 143.365 182.365 143.565 182.785 ;
        RECT 143.755 182.145 144.085 182.605 ;
        RECT 144.255 182.315 144.515 182.795 ;
        RECT 144.735 182.365 145.065 182.800 ;
        RECT 145.235 182.145 145.405 182.755 ;
        RECT 145.575 182.360 145.905 182.885 ;
        RECT 146.165 182.145 146.375 182.675 ;
        RECT 146.650 182.595 146.820 183.055 ;
        RECT 146.990 183.095 147.310 184.055 ;
        RECT 147.480 183.305 147.670 184.025 ;
        RECT 147.840 183.125 148.010 184.195 ;
        RECT 148.180 183.895 148.350 184.695 ;
        RECT 148.520 184.250 149.625 184.420 ;
        RECT 148.520 183.635 148.690 184.250 ;
        RECT 149.835 184.100 150.085 184.525 ;
        RECT 150.255 184.235 150.520 184.695 ;
        RECT 148.860 183.715 149.390 184.080 ;
        RECT 149.835 183.970 150.140 184.100 ;
        RECT 148.180 183.545 148.690 183.635 ;
        RECT 148.180 183.375 149.050 183.545 ;
        RECT 148.180 183.305 148.350 183.375 ;
        RECT 148.470 183.125 148.670 183.155 ;
        RECT 146.990 182.765 147.455 183.095 ;
        RECT 147.840 182.825 148.670 183.125 ;
        RECT 147.840 182.595 148.010 182.825 ;
        RECT 146.650 182.425 147.435 182.595 ;
        RECT 147.605 182.425 148.010 182.595 ;
        RECT 148.190 182.145 148.560 182.645 ;
        RECT 148.880 182.595 149.050 183.375 ;
        RECT 149.220 183.015 149.390 183.715 ;
        RECT 149.560 183.185 149.800 183.780 ;
        RECT 149.220 182.795 149.745 183.015 ;
        RECT 149.970 182.865 150.140 183.970 ;
        RECT 149.915 182.735 150.140 182.865 ;
        RECT 150.310 182.775 150.590 183.725 ;
        RECT 149.915 182.595 150.085 182.735 ;
        RECT 148.880 182.425 149.555 182.595 ;
        RECT 149.750 182.425 150.085 182.595 ;
        RECT 150.255 182.145 150.505 182.605 ;
        RECT 150.760 182.405 150.945 184.525 ;
        RECT 151.115 184.195 151.445 184.695 ;
        RECT 151.615 184.025 151.785 184.525 ;
        RECT 151.120 183.855 151.785 184.025 ;
        RECT 151.120 182.865 151.350 183.855 ;
        RECT 151.520 183.035 151.870 183.685 ;
        RECT 152.045 183.605 155.555 184.695 ;
        RECT 152.045 182.915 153.695 183.435 ;
        RECT 153.865 183.085 155.555 183.605 ;
        RECT 155.725 183.605 156.935 184.695 ;
        RECT 155.725 183.065 156.245 183.605 ;
        RECT 151.120 182.695 151.785 182.865 ;
        RECT 151.115 182.145 151.445 182.525 ;
        RECT 151.615 182.405 151.785 182.695 ;
        RECT 152.045 182.145 155.555 182.915 ;
        RECT 156.415 182.895 156.935 183.435 ;
        RECT 155.725 182.145 156.935 182.895 ;
        RECT 22.700 181.975 157.020 182.145 ;
        RECT 22.785 181.225 23.995 181.975 ;
        RECT 24.255 181.425 24.425 181.715 ;
        RECT 24.595 181.595 24.925 181.975 ;
        RECT 24.255 181.255 24.920 181.425 ;
        RECT 22.785 180.685 23.305 181.225 ;
        RECT 23.475 180.515 23.995 181.055 ;
        RECT 22.785 179.425 23.995 180.515 ;
        RECT 24.170 180.435 24.520 181.085 ;
        RECT 24.690 180.265 24.920 181.255 ;
        RECT 24.255 180.095 24.920 180.265 ;
        RECT 24.255 179.595 24.425 180.095 ;
        RECT 24.595 179.425 24.925 179.925 ;
        RECT 25.095 179.595 25.280 181.715 ;
        RECT 25.535 181.515 25.785 181.975 ;
        RECT 25.955 181.525 26.290 181.695 ;
        RECT 26.485 181.525 27.160 181.695 ;
        RECT 25.955 181.385 26.125 181.525 ;
        RECT 25.450 180.395 25.730 181.345 ;
        RECT 25.900 181.255 26.125 181.385 ;
        RECT 25.900 180.150 26.070 181.255 ;
        RECT 26.295 181.105 26.820 181.325 ;
        RECT 26.240 180.340 26.480 180.935 ;
        RECT 26.650 180.405 26.820 181.105 ;
        RECT 26.990 180.745 27.160 181.525 ;
        RECT 27.480 181.475 27.850 181.975 ;
        RECT 28.030 181.525 28.435 181.695 ;
        RECT 28.605 181.525 29.390 181.695 ;
        RECT 28.030 181.295 28.200 181.525 ;
        RECT 27.370 180.995 28.200 181.295 ;
        RECT 28.585 181.025 29.050 181.355 ;
        RECT 27.370 180.965 27.570 180.995 ;
        RECT 27.690 180.745 27.860 180.815 ;
        RECT 26.990 180.575 27.860 180.745 ;
        RECT 27.350 180.485 27.860 180.575 ;
        RECT 25.900 180.020 26.205 180.150 ;
        RECT 26.650 180.040 27.180 180.405 ;
        RECT 25.520 179.425 25.785 179.885 ;
        RECT 25.955 179.595 26.205 180.020 ;
        RECT 27.350 179.870 27.520 180.485 ;
        RECT 26.415 179.700 27.520 179.870 ;
        RECT 27.690 179.425 27.860 180.225 ;
        RECT 28.030 179.925 28.200 180.995 ;
        RECT 28.370 180.095 28.560 180.815 ;
        RECT 28.730 180.065 29.050 181.025 ;
        RECT 29.220 181.065 29.390 181.525 ;
        RECT 29.665 181.445 29.875 181.975 ;
        RECT 30.135 181.235 30.465 181.760 ;
        RECT 30.635 181.365 30.805 181.975 ;
        RECT 30.975 181.320 31.305 181.755 ;
        RECT 31.690 181.465 31.930 181.975 ;
        RECT 32.110 181.465 32.390 181.795 ;
        RECT 32.620 181.465 32.835 181.975 ;
        RECT 30.975 181.235 31.355 181.320 ;
        RECT 30.265 181.065 30.465 181.235 ;
        RECT 31.130 181.195 31.355 181.235 ;
        RECT 29.220 180.735 30.095 181.065 ;
        RECT 30.265 180.735 31.015 181.065 ;
        RECT 28.030 179.595 28.280 179.925 ;
        RECT 29.220 179.895 29.390 180.735 ;
        RECT 30.265 180.530 30.455 180.735 ;
        RECT 31.185 180.615 31.355 181.195 ;
        RECT 31.585 180.735 31.940 181.295 ;
        RECT 31.140 180.565 31.355 180.615 ;
        RECT 32.110 180.565 32.280 181.465 ;
        RECT 32.450 180.735 32.715 181.295 ;
        RECT 33.005 181.235 33.620 181.805 ;
        RECT 33.915 181.425 34.085 181.715 ;
        RECT 34.255 181.595 34.585 181.975 ;
        RECT 33.915 181.255 34.580 181.425 ;
        RECT 32.965 180.565 33.135 181.065 ;
        RECT 29.560 180.155 30.455 180.530 ;
        RECT 30.965 180.485 31.355 180.565 ;
        RECT 28.505 179.725 29.390 179.895 ;
        RECT 29.570 179.425 29.885 179.925 ;
        RECT 30.115 179.595 30.455 180.155 ;
        RECT 30.625 179.425 30.795 180.435 ;
        RECT 30.965 179.640 31.295 180.485 ;
        RECT 31.710 180.395 33.135 180.565 ;
        RECT 31.710 180.220 32.100 180.395 ;
        RECT 32.585 179.425 32.915 180.225 ;
        RECT 33.305 180.215 33.620 181.235 ;
        RECT 33.830 180.435 34.180 181.085 ;
        RECT 34.350 180.265 34.580 181.255 ;
        RECT 33.085 179.595 33.620 180.215 ;
        RECT 33.915 180.095 34.580 180.265 ;
        RECT 33.915 179.595 34.085 180.095 ;
        RECT 34.255 179.425 34.585 179.925 ;
        RECT 34.755 179.595 34.940 181.715 ;
        RECT 35.195 181.515 35.445 181.975 ;
        RECT 35.615 181.525 35.950 181.695 ;
        RECT 36.145 181.525 36.820 181.695 ;
        RECT 35.615 181.385 35.785 181.525 ;
        RECT 35.110 180.395 35.390 181.345 ;
        RECT 35.560 181.255 35.785 181.385 ;
        RECT 35.560 180.150 35.730 181.255 ;
        RECT 35.955 181.105 36.480 181.325 ;
        RECT 35.900 180.340 36.140 180.935 ;
        RECT 36.310 180.405 36.480 181.105 ;
        RECT 36.650 180.745 36.820 181.525 ;
        RECT 37.140 181.475 37.510 181.975 ;
        RECT 37.690 181.525 38.095 181.695 ;
        RECT 38.265 181.525 39.050 181.695 ;
        RECT 37.690 181.295 37.860 181.525 ;
        RECT 37.030 180.995 37.860 181.295 ;
        RECT 38.245 181.025 38.710 181.355 ;
        RECT 37.030 180.965 37.230 180.995 ;
        RECT 37.350 180.745 37.520 180.815 ;
        RECT 36.650 180.575 37.520 180.745 ;
        RECT 37.010 180.485 37.520 180.575 ;
        RECT 35.560 180.020 35.865 180.150 ;
        RECT 36.310 180.040 36.840 180.405 ;
        RECT 35.180 179.425 35.445 179.885 ;
        RECT 35.615 179.595 35.865 180.020 ;
        RECT 37.010 179.870 37.180 180.485 ;
        RECT 36.075 179.700 37.180 179.870 ;
        RECT 37.350 179.425 37.520 180.225 ;
        RECT 37.690 179.925 37.860 180.995 ;
        RECT 38.030 180.095 38.220 180.815 ;
        RECT 38.390 180.065 38.710 181.025 ;
        RECT 38.880 181.065 39.050 181.525 ;
        RECT 39.325 181.445 39.535 181.975 ;
        RECT 39.795 181.235 40.125 181.760 ;
        RECT 40.295 181.365 40.465 181.975 ;
        RECT 40.635 181.320 40.965 181.755 ;
        RECT 40.635 181.235 41.015 181.320 ;
        RECT 39.925 181.065 40.125 181.235 ;
        RECT 40.790 181.195 41.015 181.235 ;
        RECT 38.880 180.735 39.755 181.065 ;
        RECT 39.925 180.735 40.675 181.065 ;
        RECT 37.690 179.595 37.940 179.925 ;
        RECT 38.880 179.895 39.050 180.735 ;
        RECT 39.925 180.530 40.115 180.735 ;
        RECT 40.845 180.615 41.015 181.195 ;
        RECT 40.800 180.565 41.015 180.615 ;
        RECT 39.220 180.155 40.115 180.530 ;
        RECT 40.625 180.485 41.015 180.565 ;
        RECT 42.105 181.300 42.380 181.645 ;
        RECT 42.570 181.575 42.945 181.975 ;
        RECT 43.115 181.405 43.285 181.755 ;
        RECT 43.455 181.575 43.785 181.975 ;
        RECT 43.955 181.405 44.215 181.805 ;
        RECT 42.105 180.565 42.275 181.300 ;
        RECT 42.550 181.235 44.215 181.405 ;
        RECT 42.550 181.065 42.720 181.235 ;
        RECT 44.395 181.155 44.725 181.575 ;
        RECT 44.895 181.155 45.155 181.975 ;
        RECT 45.325 181.155 45.585 181.975 ;
        RECT 45.755 181.155 46.085 181.575 ;
        RECT 46.265 181.405 46.525 181.805 ;
        RECT 46.695 181.575 47.025 181.975 ;
        RECT 47.195 181.405 47.365 181.755 ;
        RECT 47.535 181.575 47.910 181.975 ;
        RECT 46.265 181.235 47.930 181.405 ;
        RECT 48.100 181.300 48.375 181.645 ;
        RECT 44.395 181.065 44.645 181.155 ;
        RECT 42.445 180.735 42.720 181.065 ;
        RECT 42.890 180.735 43.715 181.065 ;
        RECT 43.930 180.735 44.645 181.065 ;
        RECT 45.835 181.065 46.085 181.155 ;
        RECT 47.760 181.065 47.930 181.235 ;
        RECT 44.815 180.735 45.150 180.985 ;
        RECT 45.330 180.735 45.665 180.985 ;
        RECT 45.835 180.735 46.550 181.065 ;
        RECT 46.765 180.735 47.590 181.065 ;
        RECT 47.760 180.735 48.035 181.065 ;
        RECT 42.550 180.565 42.720 180.735 ;
        RECT 38.165 179.725 39.050 179.895 ;
        RECT 39.230 179.425 39.545 179.925 ;
        RECT 39.775 179.595 40.115 180.155 ;
        RECT 40.285 179.425 40.455 180.435 ;
        RECT 40.625 179.640 40.955 180.485 ;
        RECT 42.105 179.595 42.380 180.565 ;
        RECT 42.550 180.395 43.210 180.565 ;
        RECT 43.470 180.445 43.715 180.735 ;
        RECT 43.040 180.275 43.210 180.395 ;
        RECT 43.885 180.275 44.215 180.565 ;
        RECT 42.590 179.425 42.870 180.225 ;
        RECT 43.040 180.105 44.215 180.275 ;
        RECT 44.475 180.175 44.645 180.735 ;
        RECT 43.040 179.605 44.655 179.935 ;
        RECT 44.895 179.425 45.155 180.565 ;
        RECT 45.325 179.425 45.585 180.565 ;
        RECT 45.835 180.175 46.005 180.735 ;
        RECT 46.265 180.275 46.595 180.565 ;
        RECT 46.765 180.445 47.010 180.735 ;
        RECT 47.760 180.565 47.930 180.735 ;
        RECT 48.205 180.565 48.375 181.300 ;
        RECT 48.545 181.250 48.835 181.975 ;
        RECT 49.005 181.430 54.350 181.975 ;
        RECT 54.575 181.505 54.865 181.975 ;
        RECT 50.590 180.600 50.930 181.430 ;
        RECT 55.035 181.335 55.365 181.805 ;
        RECT 55.535 181.505 55.705 181.975 ;
        RECT 55.875 181.335 56.205 181.805 ;
        RECT 55.035 181.325 56.205 181.335 ;
        RECT 54.605 181.155 56.205 181.325 ;
        RECT 56.375 181.155 56.650 181.975 ;
        RECT 57.745 181.475 58.005 181.805 ;
        RECT 58.175 181.615 58.505 181.975 ;
        RECT 58.760 181.595 60.060 181.805 ;
        RECT 47.270 180.395 47.930 180.565 ;
        RECT 47.270 180.275 47.440 180.395 ;
        RECT 46.265 180.105 47.440 180.275 ;
        RECT 45.825 179.605 47.440 179.935 ;
        RECT 47.610 179.425 47.890 180.225 ;
        RECT 48.100 179.595 48.375 180.565 ;
        RECT 48.545 179.425 48.835 180.590 ;
        RECT 52.410 179.860 52.760 181.110 ;
        RECT 54.605 180.615 54.820 181.155 ;
        RECT 54.990 180.785 55.760 180.985 ;
        RECT 55.930 180.785 56.650 180.985 ;
        RECT 54.585 180.445 55.365 180.615 ;
        RECT 54.605 180.395 55.365 180.445 ;
        RECT 49.005 179.425 54.350 179.860 ;
        RECT 54.565 179.765 54.865 180.225 ;
        RECT 55.035 179.935 55.365 180.395 ;
        RECT 55.535 180.395 56.650 180.605 ;
        RECT 55.535 179.765 55.705 180.395 ;
        RECT 54.565 179.595 55.705 179.765 ;
        RECT 55.875 179.425 56.205 180.225 ;
        RECT 56.375 179.595 56.650 180.395 ;
        RECT 57.745 180.275 57.915 181.475 ;
        RECT 58.760 181.445 58.930 181.595 ;
        RECT 58.175 181.320 58.930 181.445 ;
        RECT 58.085 181.275 58.930 181.320 ;
        RECT 58.085 181.155 58.355 181.275 ;
        RECT 58.085 180.580 58.255 181.155 ;
        RECT 58.485 180.715 58.895 181.020 ;
        RECT 59.185 180.985 59.395 181.385 ;
        RECT 59.065 180.775 59.395 180.985 ;
        RECT 59.640 180.985 59.860 181.385 ;
        RECT 60.335 181.210 60.790 181.975 ;
        RECT 60.965 181.225 62.175 181.975 ;
        RECT 62.345 181.235 62.730 181.805 ;
        RECT 62.900 181.515 63.225 181.975 ;
        RECT 63.745 181.345 64.025 181.805 ;
        RECT 59.640 180.775 60.115 180.985 ;
        RECT 60.305 180.785 60.795 180.985 ;
        RECT 60.965 180.685 61.485 181.225 ;
        RECT 58.085 180.545 58.285 180.580 ;
        RECT 59.615 180.545 60.790 180.605 ;
        RECT 58.085 180.435 60.790 180.545 ;
        RECT 61.655 180.515 62.175 181.055 ;
        RECT 58.145 180.375 59.945 180.435 ;
        RECT 59.615 180.345 59.945 180.375 ;
        RECT 57.745 179.595 58.005 180.275 ;
        RECT 58.175 179.425 58.425 180.205 ;
        RECT 58.675 180.175 59.510 180.185 ;
        RECT 60.100 180.175 60.285 180.265 ;
        RECT 58.675 179.975 60.285 180.175 ;
        RECT 58.675 179.595 58.925 179.975 ;
        RECT 60.055 179.935 60.285 179.975 ;
        RECT 60.535 179.815 60.790 180.435 ;
        RECT 59.095 179.425 59.450 179.805 ;
        RECT 60.455 179.595 60.790 179.815 ;
        RECT 60.965 179.425 62.175 180.515 ;
        RECT 62.345 180.565 62.625 181.235 ;
        RECT 62.900 181.175 64.025 181.345 ;
        RECT 62.900 181.065 63.350 181.175 ;
        RECT 62.795 180.735 63.350 181.065 ;
        RECT 64.215 181.005 64.615 181.805 ;
        RECT 65.015 181.515 65.285 181.975 ;
        RECT 65.455 181.345 65.740 181.805 ;
        RECT 62.345 179.595 62.730 180.565 ;
        RECT 62.900 180.275 63.350 180.735 ;
        RECT 63.520 180.445 64.615 181.005 ;
        RECT 62.900 180.055 64.025 180.275 ;
        RECT 62.900 179.425 63.225 179.885 ;
        RECT 63.745 179.595 64.025 180.055 ;
        RECT 64.215 179.595 64.615 180.445 ;
        RECT 64.785 181.175 65.740 181.345 ;
        RECT 66.965 181.245 67.255 181.975 ;
        RECT 64.785 180.275 64.995 181.175 ;
        RECT 65.165 180.445 65.855 181.005 ;
        RECT 66.955 180.735 67.255 181.065 ;
        RECT 67.435 181.045 67.665 181.685 ;
        RECT 67.845 181.425 68.155 181.795 ;
        RECT 68.335 181.605 69.005 181.975 ;
        RECT 67.845 181.225 69.075 181.425 ;
        RECT 67.435 180.735 67.960 181.045 ;
        RECT 68.140 180.735 68.605 181.045 ;
        RECT 68.785 180.555 69.075 181.225 ;
        RECT 66.965 180.315 68.125 180.555 ;
        RECT 64.785 180.055 65.740 180.275 ;
        RECT 65.015 179.425 65.285 179.885 ;
        RECT 65.455 179.595 65.740 180.055 ;
        RECT 66.965 179.605 67.225 180.315 ;
        RECT 67.395 179.425 67.725 180.135 ;
        RECT 67.895 179.605 68.125 180.315 ;
        RECT 68.305 180.335 69.075 180.555 ;
        RECT 68.305 179.605 68.575 180.335 ;
        RECT 68.755 179.425 69.095 180.155 ;
        RECT 69.265 179.605 69.525 181.795 ;
        RECT 69.705 181.235 70.090 181.805 ;
        RECT 70.260 181.515 70.585 181.975 ;
        RECT 71.105 181.345 71.385 181.805 ;
        RECT 69.705 180.565 69.985 181.235 ;
        RECT 70.260 181.175 71.385 181.345 ;
        RECT 70.260 181.065 70.710 181.175 ;
        RECT 70.155 180.735 70.710 181.065 ;
        RECT 71.575 181.005 71.975 181.805 ;
        RECT 72.375 181.515 72.645 181.975 ;
        RECT 72.815 181.345 73.100 181.805 ;
        RECT 69.705 179.595 70.090 180.565 ;
        RECT 70.260 180.275 70.710 180.735 ;
        RECT 70.880 180.445 71.975 181.005 ;
        RECT 70.260 180.055 71.385 180.275 ;
        RECT 70.260 179.425 70.585 179.885 ;
        RECT 71.105 179.595 71.385 180.055 ;
        RECT 71.575 179.595 71.975 180.445 ;
        RECT 72.145 181.175 73.100 181.345 ;
        RECT 74.305 181.250 74.595 181.975 ;
        RECT 75.775 181.425 75.945 181.715 ;
        RECT 76.115 181.595 76.445 181.975 ;
        RECT 75.775 181.255 76.440 181.425 ;
        RECT 72.145 180.275 72.355 181.175 ;
        RECT 72.525 180.445 73.215 181.005 ;
        RECT 72.145 180.055 73.100 180.275 ;
        RECT 72.375 179.425 72.645 179.885 ;
        RECT 72.815 179.595 73.100 180.055 ;
        RECT 74.305 179.425 74.595 180.590 ;
        RECT 75.690 180.435 76.040 181.085 ;
        RECT 76.210 180.265 76.440 181.255 ;
        RECT 75.775 180.095 76.440 180.265 ;
        RECT 75.775 179.595 75.945 180.095 ;
        RECT 76.115 179.425 76.445 179.925 ;
        RECT 76.615 179.595 76.800 181.715 ;
        RECT 77.055 181.515 77.305 181.975 ;
        RECT 77.475 181.525 77.810 181.695 ;
        RECT 78.005 181.525 78.680 181.695 ;
        RECT 77.475 181.385 77.645 181.525 ;
        RECT 76.970 180.395 77.250 181.345 ;
        RECT 77.420 181.255 77.645 181.385 ;
        RECT 77.420 180.150 77.590 181.255 ;
        RECT 77.815 181.105 78.340 181.325 ;
        RECT 77.760 180.340 78.000 180.935 ;
        RECT 78.170 180.405 78.340 181.105 ;
        RECT 78.510 180.745 78.680 181.525 ;
        RECT 79.000 181.475 79.370 181.975 ;
        RECT 79.550 181.525 79.955 181.695 ;
        RECT 80.125 181.525 80.910 181.695 ;
        RECT 79.550 181.295 79.720 181.525 ;
        RECT 78.890 180.995 79.720 181.295 ;
        RECT 80.105 181.025 80.570 181.355 ;
        RECT 78.890 180.965 79.090 180.995 ;
        RECT 79.210 180.745 79.380 180.815 ;
        RECT 78.510 180.575 79.380 180.745 ;
        RECT 78.870 180.485 79.380 180.575 ;
        RECT 77.420 180.020 77.725 180.150 ;
        RECT 78.170 180.040 78.700 180.405 ;
        RECT 77.040 179.425 77.305 179.885 ;
        RECT 77.475 179.595 77.725 180.020 ;
        RECT 78.870 179.870 79.040 180.485 ;
        RECT 77.935 179.700 79.040 179.870 ;
        RECT 79.210 179.425 79.380 180.225 ;
        RECT 79.550 179.925 79.720 180.995 ;
        RECT 79.890 180.095 80.080 180.815 ;
        RECT 80.250 180.065 80.570 181.025 ;
        RECT 80.740 181.065 80.910 181.525 ;
        RECT 81.185 181.445 81.395 181.975 ;
        RECT 81.655 181.235 81.985 181.760 ;
        RECT 82.155 181.365 82.325 181.975 ;
        RECT 82.495 181.320 82.825 181.755 ;
        RECT 83.045 181.325 83.305 181.805 ;
        RECT 83.475 181.435 83.725 181.975 ;
        RECT 82.495 181.235 82.875 181.320 ;
        RECT 81.785 181.065 81.985 181.235 ;
        RECT 82.650 181.195 82.875 181.235 ;
        RECT 80.740 180.735 81.615 181.065 ;
        RECT 81.785 180.735 82.535 181.065 ;
        RECT 79.550 179.595 79.800 179.925 ;
        RECT 80.740 179.895 80.910 180.735 ;
        RECT 81.785 180.530 81.975 180.735 ;
        RECT 82.705 180.615 82.875 181.195 ;
        RECT 82.660 180.565 82.875 180.615 ;
        RECT 81.080 180.155 81.975 180.530 ;
        RECT 82.485 180.485 82.875 180.565 ;
        RECT 80.025 179.725 80.910 179.895 ;
        RECT 81.090 179.425 81.405 179.925 ;
        RECT 81.635 179.595 81.975 180.155 ;
        RECT 82.145 179.425 82.315 180.435 ;
        RECT 82.485 179.640 82.815 180.485 ;
        RECT 83.045 180.295 83.215 181.325 ;
        RECT 83.895 181.295 84.115 181.755 ;
        RECT 83.865 181.270 84.115 181.295 ;
        RECT 83.385 180.675 83.615 181.070 ;
        RECT 83.785 180.845 84.115 181.270 ;
        RECT 84.285 181.595 85.175 181.765 ;
        RECT 84.285 180.870 84.455 181.595 ;
        RECT 84.625 181.040 85.175 181.425 ;
        RECT 85.345 181.205 88.855 181.975 ;
        RECT 89.485 181.300 89.745 181.805 ;
        RECT 89.925 181.595 90.255 181.975 ;
        RECT 90.435 181.425 90.605 181.805 ;
        RECT 84.285 180.800 85.175 180.870 ;
        RECT 84.280 180.775 85.175 180.800 ;
        RECT 84.270 180.760 85.175 180.775 ;
        RECT 84.265 180.745 85.175 180.760 ;
        RECT 84.255 180.740 85.175 180.745 ;
        RECT 84.250 180.730 85.175 180.740 ;
        RECT 84.245 180.720 85.175 180.730 ;
        RECT 84.235 180.715 85.175 180.720 ;
        RECT 84.225 180.705 85.175 180.715 ;
        RECT 84.215 180.700 85.175 180.705 ;
        RECT 84.215 180.695 84.550 180.700 ;
        RECT 84.200 180.690 84.550 180.695 ;
        RECT 84.185 180.680 84.550 180.690 ;
        RECT 84.160 180.675 84.550 180.680 ;
        RECT 83.385 180.670 84.550 180.675 ;
        RECT 83.385 180.635 84.520 180.670 ;
        RECT 83.385 180.610 84.485 180.635 ;
        RECT 83.385 180.580 84.455 180.610 ;
        RECT 83.385 180.550 84.435 180.580 ;
        RECT 83.385 180.520 84.415 180.550 ;
        RECT 83.385 180.510 84.345 180.520 ;
        RECT 83.385 180.500 84.320 180.510 ;
        RECT 83.385 180.485 84.300 180.500 ;
        RECT 83.385 180.470 84.280 180.485 ;
        RECT 83.490 180.460 84.275 180.470 ;
        RECT 83.490 180.425 84.260 180.460 ;
        RECT 83.045 179.595 83.320 180.295 ;
        RECT 83.490 180.175 84.245 180.425 ;
        RECT 84.415 180.105 84.745 180.350 ;
        RECT 84.915 180.250 85.175 180.700 ;
        RECT 85.345 180.685 86.995 181.205 ;
        RECT 87.165 180.515 88.855 181.035 ;
        RECT 84.560 180.080 84.745 180.105 ;
        RECT 84.560 179.980 85.175 180.080 ;
        RECT 83.490 179.425 83.745 179.970 ;
        RECT 83.915 179.595 84.395 179.935 ;
        RECT 84.570 179.425 85.175 179.980 ;
        RECT 85.345 179.425 88.855 180.515 ;
        RECT 89.485 180.500 89.655 181.300 ;
        RECT 89.940 181.255 90.605 181.425 ;
        RECT 89.940 181.000 90.110 181.255 ;
        RECT 91.790 181.235 92.045 181.805 ;
        RECT 92.215 181.575 92.545 181.975 ;
        RECT 92.970 181.440 93.500 181.805 ;
        RECT 92.970 181.405 93.145 181.440 ;
        RECT 92.215 181.235 93.145 181.405 ;
        RECT 89.825 180.670 90.110 181.000 ;
        RECT 90.345 180.705 90.675 181.075 ;
        RECT 89.940 180.525 90.110 180.670 ;
        RECT 91.790 180.565 91.960 181.235 ;
        RECT 92.215 181.065 92.385 181.235 ;
        RECT 92.130 180.735 92.385 181.065 ;
        RECT 92.610 180.735 92.805 181.065 ;
        RECT 89.485 179.595 89.755 180.500 ;
        RECT 89.940 180.355 90.605 180.525 ;
        RECT 89.925 179.425 90.255 180.185 ;
        RECT 90.435 179.595 90.605 180.355 ;
        RECT 91.790 179.595 92.125 180.565 ;
        RECT 92.295 179.425 92.465 180.565 ;
        RECT 92.635 179.765 92.805 180.735 ;
        RECT 92.975 180.105 93.145 181.235 ;
        RECT 93.315 180.445 93.485 181.245 ;
        RECT 93.690 180.955 93.965 181.805 ;
        RECT 93.685 180.785 93.965 180.955 ;
        RECT 93.690 180.645 93.965 180.785 ;
        RECT 94.135 180.445 94.325 181.805 ;
        RECT 94.505 181.440 95.015 181.975 ;
        RECT 95.235 181.165 95.480 181.770 ;
        RECT 95.925 181.205 99.435 181.975 ;
        RECT 100.065 181.250 100.355 181.975 ;
        RECT 100.525 181.430 105.870 181.975 ;
        RECT 94.525 180.995 95.755 181.165 ;
        RECT 93.315 180.275 94.325 180.445 ;
        RECT 94.495 180.430 95.245 180.620 ;
        RECT 92.975 179.935 94.100 180.105 ;
        RECT 94.495 179.765 94.665 180.430 ;
        RECT 95.415 180.185 95.755 180.995 ;
        RECT 95.925 180.685 97.575 181.205 ;
        RECT 97.745 180.515 99.435 181.035 ;
        RECT 102.110 180.600 102.450 181.430 ;
        RECT 106.045 181.205 108.635 181.975 ;
        RECT 108.895 181.425 109.065 181.715 ;
        RECT 109.235 181.595 109.565 181.975 ;
        RECT 108.895 181.255 109.560 181.425 ;
        RECT 92.635 179.595 94.665 179.765 ;
        RECT 94.835 179.425 95.005 180.185 ;
        RECT 95.240 179.775 95.755 180.185 ;
        RECT 95.925 179.425 99.435 180.515 ;
        RECT 100.065 179.425 100.355 180.590 ;
        RECT 103.930 179.860 104.280 181.110 ;
        RECT 106.045 180.685 107.255 181.205 ;
        RECT 107.425 180.515 108.635 181.035 ;
        RECT 100.525 179.425 105.870 179.860 ;
        RECT 106.045 179.425 108.635 180.515 ;
        RECT 108.810 180.435 109.160 181.085 ;
        RECT 109.330 180.265 109.560 181.255 ;
        RECT 108.895 180.095 109.560 180.265 ;
        RECT 108.895 179.595 109.065 180.095 ;
        RECT 109.235 179.425 109.565 179.925 ;
        RECT 109.735 179.595 109.920 181.715 ;
        RECT 110.175 181.515 110.425 181.975 ;
        RECT 110.595 181.525 110.930 181.695 ;
        RECT 111.125 181.525 111.800 181.695 ;
        RECT 110.595 181.385 110.765 181.525 ;
        RECT 110.090 180.395 110.370 181.345 ;
        RECT 110.540 181.255 110.765 181.385 ;
        RECT 110.540 180.150 110.710 181.255 ;
        RECT 110.935 181.105 111.460 181.325 ;
        RECT 110.880 180.340 111.120 180.935 ;
        RECT 111.290 180.405 111.460 181.105 ;
        RECT 111.630 180.745 111.800 181.525 ;
        RECT 112.120 181.475 112.490 181.975 ;
        RECT 112.670 181.525 113.075 181.695 ;
        RECT 113.245 181.525 114.030 181.695 ;
        RECT 112.670 181.295 112.840 181.525 ;
        RECT 112.010 180.995 112.840 181.295 ;
        RECT 113.225 181.025 113.690 181.355 ;
        RECT 112.010 180.965 112.210 180.995 ;
        RECT 112.330 180.745 112.500 180.815 ;
        RECT 111.630 180.575 112.500 180.745 ;
        RECT 111.990 180.485 112.500 180.575 ;
        RECT 110.540 180.020 110.845 180.150 ;
        RECT 111.290 180.040 111.820 180.405 ;
        RECT 110.160 179.425 110.425 179.885 ;
        RECT 110.595 179.595 110.845 180.020 ;
        RECT 111.990 179.870 112.160 180.485 ;
        RECT 111.055 179.700 112.160 179.870 ;
        RECT 112.330 179.425 112.500 180.225 ;
        RECT 112.670 179.925 112.840 180.995 ;
        RECT 113.010 180.095 113.200 180.815 ;
        RECT 113.370 180.065 113.690 181.025 ;
        RECT 113.860 181.065 114.030 181.525 ;
        RECT 114.305 181.445 114.515 181.975 ;
        RECT 114.775 181.235 115.105 181.760 ;
        RECT 115.275 181.365 115.445 181.975 ;
        RECT 115.615 181.320 115.945 181.755 ;
        RECT 115.615 181.235 115.995 181.320 ;
        RECT 114.905 181.065 115.105 181.235 ;
        RECT 115.770 181.195 115.995 181.235 ;
        RECT 113.860 180.735 114.735 181.065 ;
        RECT 114.905 180.735 115.655 181.065 ;
        RECT 112.670 179.595 112.920 179.925 ;
        RECT 113.860 179.895 114.030 180.735 ;
        RECT 114.905 180.530 115.095 180.735 ;
        RECT 115.825 180.615 115.995 181.195 ;
        RECT 116.165 181.205 119.675 181.975 ;
        RECT 116.165 180.685 117.815 181.205 ;
        RECT 120.805 181.155 121.035 181.975 ;
        RECT 121.205 181.175 121.535 181.805 ;
        RECT 115.780 180.565 115.995 180.615 ;
        RECT 114.200 180.155 115.095 180.530 ;
        RECT 115.605 180.485 115.995 180.565 ;
        RECT 117.985 180.515 119.675 181.035 ;
        RECT 120.785 180.735 121.115 180.985 ;
        RECT 121.285 180.575 121.535 181.175 ;
        RECT 121.705 181.155 121.915 181.975 ;
        RECT 122.145 181.205 125.655 181.975 ;
        RECT 125.825 181.250 126.115 181.975 ;
        RECT 122.145 180.685 123.795 181.205 ;
        RECT 113.145 179.725 114.030 179.895 ;
        RECT 114.210 179.425 114.525 179.925 ;
        RECT 114.755 179.595 115.095 180.155 ;
        RECT 115.265 179.425 115.435 180.435 ;
        RECT 115.605 179.640 115.935 180.485 ;
        RECT 116.165 179.425 119.675 180.515 ;
        RECT 120.805 179.425 121.035 180.565 ;
        RECT 121.205 179.595 121.535 180.575 ;
        RECT 121.705 179.425 121.915 180.565 ;
        RECT 123.965 180.515 125.655 181.035 ;
        RECT 122.145 179.425 125.655 180.515 ;
        RECT 125.825 179.425 126.115 180.590 ;
        RECT 126.765 180.395 126.995 181.735 ;
        RECT 127.175 180.895 127.405 181.795 ;
        RECT 127.605 181.195 127.850 181.975 ;
        RECT 128.020 181.435 128.450 181.795 ;
        RECT 129.030 181.605 129.760 181.975 ;
        RECT 128.020 181.245 129.760 181.435 ;
        RECT 128.020 181.015 128.240 181.245 ;
        RECT 127.175 180.215 127.515 180.895 ;
        RECT 126.765 180.015 127.515 180.215 ;
        RECT 127.695 180.715 128.240 181.015 ;
        RECT 126.765 179.625 127.005 180.015 ;
        RECT 127.175 179.425 127.525 179.835 ;
        RECT 127.695 179.605 128.025 180.715 ;
        RECT 128.410 180.445 128.835 181.065 ;
        RECT 129.030 180.445 129.290 181.065 ;
        RECT 129.500 180.735 129.760 181.245 ;
        RECT 128.195 180.075 129.220 180.275 ;
        RECT 128.195 179.605 128.375 180.075 ;
        RECT 128.545 179.425 128.875 179.905 ;
        RECT 129.050 179.605 129.220 180.075 ;
        RECT 129.485 179.425 129.770 180.565 ;
        RECT 129.960 179.605 130.240 181.795 ;
        RECT 130.755 181.575 131.085 181.975 ;
        RECT 131.255 181.405 131.585 181.745 ;
        RECT 132.635 181.575 132.965 181.975 ;
        RECT 130.600 181.235 132.965 181.405 ;
        RECT 133.135 181.250 133.465 181.760 ;
        RECT 130.600 180.235 130.770 181.235 ;
        RECT 132.795 181.065 132.965 181.235 ;
        RECT 130.940 180.405 131.185 181.065 ;
        RECT 131.400 180.405 131.665 181.065 ;
        RECT 131.860 180.405 132.145 181.065 ;
        RECT 132.320 180.735 132.625 181.065 ;
        RECT 132.795 180.735 133.105 181.065 ;
        RECT 132.320 180.405 132.535 180.735 ;
        RECT 133.275 180.615 133.465 181.250 ;
        RECT 133.845 181.345 134.175 181.705 ;
        RECT 134.795 181.515 135.045 181.975 ;
        RECT 135.215 181.515 135.775 181.805 ;
        RECT 133.845 181.155 135.235 181.345 ;
        RECT 135.065 181.065 135.235 181.155 ;
        RECT 130.600 180.065 131.055 180.235 ;
        RECT 130.725 179.635 131.055 180.065 ;
        RECT 131.235 180.065 132.525 180.235 ;
        RECT 131.235 179.645 131.485 180.065 ;
        RECT 131.715 179.425 132.045 179.895 ;
        RECT 132.275 179.645 132.525 180.065 ;
        RECT 132.715 179.425 132.965 180.565 ;
        RECT 133.245 180.485 133.465 180.615 ;
        RECT 133.135 179.635 133.465 180.485 ;
        RECT 133.660 180.735 134.335 180.985 ;
        RECT 134.555 180.735 134.895 180.985 ;
        RECT 135.065 180.735 135.355 181.065 ;
        RECT 133.660 180.375 133.925 180.735 ;
        RECT 135.065 180.485 135.235 180.735 ;
        RECT 134.295 180.315 135.235 180.485 ;
        RECT 133.845 179.425 134.125 180.095 ;
        RECT 134.295 179.765 134.595 180.315 ;
        RECT 135.525 180.145 135.775 181.515 ;
        RECT 134.795 179.425 135.125 180.145 ;
        RECT 135.315 179.595 135.775 180.145 ;
        RECT 136.900 181.235 137.515 181.805 ;
        RECT 137.685 181.465 137.900 181.975 ;
        RECT 138.130 181.465 138.410 181.795 ;
        RECT 138.590 181.465 138.830 181.975 ;
        RECT 136.900 180.215 137.215 181.235 ;
        RECT 137.385 180.565 137.555 181.065 ;
        RECT 137.805 180.735 138.070 181.295 ;
        RECT 138.240 180.565 138.410 181.465 ;
        RECT 138.580 180.735 138.935 181.295 ;
        RECT 139.165 181.175 139.860 181.805 ;
        RECT 140.065 181.175 140.375 181.975 ;
        RECT 140.545 181.205 142.215 181.975 ;
        RECT 142.845 181.475 143.105 181.805 ;
        RECT 143.315 181.495 143.590 181.975 ;
        RECT 139.185 180.735 139.520 180.985 ;
        RECT 139.690 180.575 139.860 181.175 ;
        RECT 140.030 180.735 140.365 181.005 ;
        RECT 140.545 180.685 141.295 181.205 ;
        RECT 137.385 180.395 138.810 180.565 ;
        RECT 136.900 179.595 137.435 180.215 ;
        RECT 137.605 179.425 137.935 180.225 ;
        RECT 138.420 180.220 138.810 180.395 ;
        RECT 139.165 179.425 139.425 180.565 ;
        RECT 139.595 179.595 139.925 180.575 ;
        RECT 140.095 179.425 140.375 180.565 ;
        RECT 141.465 180.515 142.215 181.035 ;
        RECT 140.545 179.425 142.215 180.515 ;
        RECT 142.845 180.565 143.015 181.475 ;
        RECT 143.800 181.405 144.005 181.805 ;
        RECT 144.175 181.575 144.510 181.975 ;
        RECT 145.235 181.425 145.405 181.805 ;
        RECT 145.585 181.595 145.915 181.975 ;
        RECT 143.185 180.735 143.545 181.315 ;
        RECT 143.800 181.235 144.485 181.405 ;
        RECT 145.235 181.255 145.900 181.425 ;
        RECT 146.095 181.300 146.355 181.805 ;
        RECT 146.585 181.515 146.830 181.975 ;
        RECT 143.725 180.565 143.975 181.065 ;
        RECT 142.845 180.395 143.975 180.565 ;
        RECT 142.845 179.625 143.115 180.395 ;
        RECT 144.145 180.205 144.485 181.235 ;
        RECT 145.165 180.705 145.495 181.075 ;
        RECT 145.730 181.000 145.900 181.255 ;
        RECT 145.730 180.670 146.015 181.000 ;
        RECT 145.730 180.525 145.900 180.670 ;
        RECT 143.285 179.425 143.615 180.205 ;
        RECT 143.820 180.030 144.485 180.205 ;
        RECT 145.235 180.355 145.900 180.525 ;
        RECT 146.185 180.500 146.355 181.300 ;
        RECT 146.525 180.735 146.840 181.345 ;
        RECT 147.010 180.985 147.260 181.795 ;
        RECT 147.430 181.450 147.690 181.975 ;
        RECT 147.860 181.325 148.120 181.780 ;
        RECT 148.290 181.495 148.550 181.975 ;
        RECT 148.720 181.325 148.980 181.780 ;
        RECT 149.150 181.495 149.410 181.975 ;
        RECT 149.580 181.325 149.840 181.780 ;
        RECT 150.010 181.495 150.270 181.975 ;
        RECT 150.440 181.325 150.700 181.780 ;
        RECT 150.870 181.495 151.170 181.975 ;
        RECT 147.860 181.155 151.170 181.325 ;
        RECT 151.585 181.250 151.875 181.975 ;
        RECT 147.010 180.735 150.030 180.985 ;
        RECT 143.820 179.625 144.005 180.030 ;
        RECT 144.175 179.425 144.510 179.850 ;
        RECT 145.235 179.595 145.405 180.355 ;
        RECT 145.585 179.425 145.915 180.185 ;
        RECT 146.085 179.595 146.355 180.500 ;
        RECT 146.535 179.425 146.830 180.535 ;
        RECT 147.010 179.600 147.260 180.735 ;
        RECT 150.200 180.565 151.170 181.155 ;
        RECT 152.045 181.205 155.555 181.975 ;
        RECT 155.725 181.225 156.935 181.975 ;
        RECT 152.045 180.685 153.695 181.205 ;
        RECT 147.430 179.425 147.690 180.535 ;
        RECT 147.860 180.325 151.170 180.565 ;
        RECT 147.860 179.600 148.120 180.325 ;
        RECT 148.290 179.425 148.550 180.155 ;
        RECT 148.720 179.600 148.980 180.325 ;
        RECT 149.150 179.425 149.410 180.155 ;
        RECT 149.580 179.600 149.840 180.325 ;
        RECT 150.010 179.425 150.270 180.155 ;
        RECT 150.440 179.600 150.700 180.325 ;
        RECT 150.870 179.425 151.165 180.155 ;
        RECT 151.585 179.425 151.875 180.590 ;
        RECT 153.865 180.515 155.555 181.035 ;
        RECT 152.045 179.425 155.555 180.515 ;
        RECT 155.725 180.515 156.245 181.055 ;
        RECT 156.415 180.685 156.935 181.225 ;
        RECT 155.725 179.425 156.935 180.515 ;
        RECT 22.700 179.255 157.020 179.425 ;
        RECT 22.785 178.165 23.995 179.255 ;
        RECT 22.785 177.455 23.305 177.995 ;
        RECT 23.475 177.625 23.995 178.165 ;
        RECT 25.085 178.180 25.355 179.085 ;
        RECT 25.525 178.495 25.855 179.255 ;
        RECT 26.035 178.325 26.205 179.085 ;
        RECT 22.785 176.705 23.995 177.455 ;
        RECT 25.085 177.380 25.255 178.180 ;
        RECT 25.540 178.155 26.205 178.325 ;
        RECT 26.465 178.165 28.135 179.255 ;
        RECT 25.540 178.010 25.710 178.155 ;
        RECT 25.425 177.680 25.710 178.010 ;
        RECT 25.540 177.425 25.710 177.680 ;
        RECT 25.945 177.605 26.275 177.975 ;
        RECT 26.465 177.475 27.215 177.995 ;
        RECT 27.385 177.645 28.135 178.165 ;
        RECT 28.305 178.385 28.580 179.085 ;
        RECT 28.750 178.710 29.005 179.255 ;
        RECT 29.175 178.745 29.655 179.085 ;
        RECT 29.830 178.700 30.435 179.255 ;
        RECT 29.820 178.600 30.435 178.700 ;
        RECT 29.820 178.575 30.005 178.600 ;
        RECT 25.085 176.875 25.345 177.380 ;
        RECT 25.540 177.255 26.205 177.425 ;
        RECT 25.525 176.705 25.855 177.085 ;
        RECT 26.035 176.875 26.205 177.255 ;
        RECT 26.465 176.705 28.135 177.475 ;
        RECT 28.305 177.355 28.475 178.385 ;
        RECT 28.750 178.255 29.505 178.505 ;
        RECT 29.675 178.330 30.005 178.575 ;
        RECT 28.750 178.220 29.520 178.255 ;
        RECT 28.750 178.210 29.535 178.220 ;
        RECT 28.645 178.195 29.540 178.210 ;
        RECT 28.645 178.180 29.560 178.195 ;
        RECT 28.645 178.170 29.580 178.180 ;
        RECT 28.645 178.160 29.605 178.170 ;
        RECT 28.645 178.130 29.675 178.160 ;
        RECT 28.645 178.100 29.695 178.130 ;
        RECT 28.645 178.070 29.715 178.100 ;
        RECT 28.645 178.045 29.745 178.070 ;
        RECT 28.645 178.010 29.780 178.045 ;
        RECT 28.645 178.005 29.810 178.010 ;
        RECT 28.645 177.610 28.875 178.005 ;
        RECT 29.420 178.000 29.810 178.005 ;
        RECT 29.445 177.990 29.810 178.000 ;
        RECT 29.460 177.985 29.810 177.990 ;
        RECT 29.475 177.980 29.810 177.985 ;
        RECT 30.175 177.980 30.435 178.430 ;
        RECT 30.605 178.165 31.815 179.255 ;
        RECT 31.985 178.700 32.590 179.255 ;
        RECT 32.765 178.745 33.245 179.085 ;
        RECT 33.415 178.710 33.670 179.255 ;
        RECT 31.985 178.600 32.600 178.700 ;
        RECT 32.415 178.575 32.600 178.600 ;
        RECT 29.475 177.975 30.435 177.980 ;
        RECT 29.485 177.965 30.435 177.975 ;
        RECT 29.495 177.960 30.435 177.965 ;
        RECT 29.505 177.950 30.435 177.960 ;
        RECT 29.510 177.940 30.435 177.950 ;
        RECT 29.515 177.935 30.435 177.940 ;
        RECT 29.525 177.920 30.435 177.935 ;
        RECT 29.530 177.905 30.435 177.920 ;
        RECT 29.540 177.880 30.435 177.905 ;
        RECT 29.045 177.410 29.375 177.835 ;
        RECT 28.305 176.875 28.565 177.355 ;
        RECT 28.735 176.705 28.985 177.245 ;
        RECT 29.155 176.925 29.375 177.410 ;
        RECT 29.545 177.810 30.435 177.880 ;
        RECT 29.545 177.085 29.715 177.810 ;
        RECT 29.885 177.255 30.435 177.640 ;
        RECT 30.605 177.455 31.125 177.995 ;
        RECT 31.295 177.625 31.815 178.165 ;
        RECT 31.985 177.980 32.245 178.430 ;
        RECT 32.415 178.330 32.745 178.575 ;
        RECT 32.915 178.255 33.670 178.505 ;
        RECT 33.840 178.385 34.115 179.085 ;
        RECT 32.900 178.220 33.670 178.255 ;
        RECT 32.885 178.210 33.670 178.220 ;
        RECT 32.880 178.195 33.775 178.210 ;
        RECT 32.860 178.180 33.775 178.195 ;
        RECT 32.840 178.170 33.775 178.180 ;
        RECT 32.815 178.160 33.775 178.170 ;
        RECT 32.745 178.130 33.775 178.160 ;
        RECT 32.725 178.100 33.775 178.130 ;
        RECT 32.705 178.070 33.775 178.100 ;
        RECT 32.675 178.045 33.775 178.070 ;
        RECT 32.640 178.010 33.775 178.045 ;
        RECT 32.610 178.005 33.775 178.010 ;
        RECT 32.610 178.000 33.000 178.005 ;
        RECT 32.610 177.990 32.975 178.000 ;
        RECT 32.610 177.985 32.960 177.990 ;
        RECT 32.610 177.980 32.945 177.985 ;
        RECT 31.985 177.975 32.945 177.980 ;
        RECT 31.985 177.965 32.935 177.975 ;
        RECT 31.985 177.960 32.925 177.965 ;
        RECT 31.985 177.950 32.915 177.960 ;
        RECT 31.985 177.940 32.910 177.950 ;
        RECT 31.985 177.935 32.905 177.940 ;
        RECT 31.985 177.920 32.895 177.935 ;
        RECT 31.985 177.905 32.890 177.920 ;
        RECT 31.985 177.880 32.880 177.905 ;
        RECT 31.985 177.810 32.875 177.880 ;
        RECT 29.545 176.915 30.435 177.085 ;
        RECT 30.605 176.705 31.815 177.455 ;
        RECT 31.985 177.255 32.535 177.640 ;
        RECT 32.705 177.085 32.875 177.810 ;
        RECT 31.985 176.915 32.875 177.085 ;
        RECT 33.045 177.410 33.375 177.835 ;
        RECT 33.545 177.610 33.775 178.005 ;
        RECT 33.045 177.385 33.295 177.410 ;
        RECT 33.045 176.925 33.265 177.385 ;
        RECT 33.945 177.355 34.115 178.385 ;
        RECT 34.325 178.115 34.555 179.255 ;
        RECT 34.725 178.105 35.055 179.085 ;
        RECT 35.225 178.115 35.435 179.255 ;
        RECT 34.305 177.695 34.635 177.945 ;
        RECT 33.435 176.705 33.685 177.245 ;
        RECT 33.855 176.875 34.115 177.355 ;
        RECT 34.325 176.705 34.555 177.525 ;
        RECT 34.805 177.505 35.055 178.105 ;
        RECT 35.665 178.090 35.955 179.255 ;
        RECT 36.125 178.165 39.635 179.255 ;
        RECT 34.725 176.875 35.055 177.505 ;
        RECT 35.225 176.705 35.435 177.525 ;
        RECT 36.125 177.475 37.775 177.995 ;
        RECT 37.945 177.645 39.635 178.165 ;
        RECT 40.270 178.115 40.525 179.255 ;
        RECT 40.720 178.705 41.915 179.035 ;
        RECT 40.775 177.945 40.945 178.505 ;
        RECT 41.170 178.285 41.590 178.535 ;
        RECT 42.095 178.455 42.375 179.255 ;
        RECT 41.170 178.115 42.415 178.285 ;
        RECT 42.585 178.115 42.855 179.085 ;
        RECT 42.245 177.945 42.415 178.115 ;
        RECT 40.270 177.695 40.605 177.945 ;
        RECT 40.775 177.615 41.515 177.945 ;
        RECT 42.245 177.615 42.475 177.945 ;
        RECT 40.775 177.525 41.025 177.615 ;
        RECT 35.665 176.705 35.955 177.430 ;
        RECT 36.125 176.705 39.635 177.475 ;
        RECT 40.290 177.355 41.025 177.525 ;
        RECT 42.245 177.445 42.415 177.615 ;
        RECT 40.290 176.885 40.600 177.355 ;
        RECT 41.675 177.275 42.415 177.445 ;
        RECT 42.685 177.380 42.855 178.115 ;
        RECT 40.770 176.705 41.505 177.185 ;
        RECT 41.675 176.925 41.845 177.275 ;
        RECT 42.015 176.705 42.395 177.105 ;
        RECT 42.585 177.035 42.855 177.380 ;
        RECT 43.485 178.405 43.865 179.085 ;
        RECT 44.455 178.405 44.625 179.255 ;
        RECT 44.795 178.575 45.125 179.085 ;
        RECT 45.295 178.745 45.465 179.255 ;
        RECT 45.635 178.575 46.035 179.085 ;
        RECT 44.795 178.405 46.035 178.575 ;
        RECT 43.485 177.445 43.655 178.405 ;
        RECT 43.825 178.065 45.130 178.235 ;
        RECT 46.215 178.155 46.535 179.085 ;
        RECT 46.705 178.165 48.375 179.255 ;
        RECT 48.605 178.195 48.935 179.040 ;
        RECT 49.105 178.245 49.275 179.255 ;
        RECT 49.445 178.525 49.785 179.085 ;
        RECT 50.015 178.755 50.330 179.255 ;
        RECT 50.510 178.785 51.395 178.955 ;
        RECT 43.825 177.615 44.070 178.065 ;
        RECT 44.240 177.695 44.790 177.895 ;
        RECT 44.960 177.865 45.130 178.065 ;
        RECT 45.905 177.985 46.535 178.155 ;
        RECT 44.960 177.695 45.335 177.865 ;
        RECT 45.505 177.445 45.735 177.945 ;
        RECT 43.485 177.275 45.735 177.445 ;
        RECT 43.535 176.705 43.865 177.095 ;
        RECT 44.035 176.955 44.205 177.275 ;
        RECT 45.905 177.105 46.075 177.985 ;
        RECT 44.375 176.705 44.705 177.095 ;
        RECT 45.120 176.935 46.075 177.105 ;
        RECT 46.245 176.705 46.535 177.540 ;
        RECT 46.705 177.475 47.455 177.995 ;
        RECT 47.625 177.645 48.375 178.165 ;
        RECT 48.545 178.115 48.935 178.195 ;
        RECT 49.445 178.150 50.340 178.525 ;
        RECT 48.545 178.065 48.760 178.115 ;
        RECT 48.545 177.485 48.715 178.065 ;
        RECT 49.445 177.945 49.635 178.150 ;
        RECT 50.510 177.945 50.680 178.785 ;
        RECT 51.620 178.755 51.870 179.085 ;
        RECT 48.885 177.615 49.635 177.945 ;
        RECT 49.805 177.615 50.680 177.945 ;
        RECT 46.705 176.705 48.375 177.475 ;
        RECT 48.545 177.445 48.770 177.485 ;
        RECT 49.435 177.445 49.635 177.615 ;
        RECT 48.545 177.360 48.925 177.445 ;
        RECT 48.595 176.925 48.925 177.360 ;
        RECT 49.095 176.705 49.265 177.315 ;
        RECT 49.435 176.920 49.765 177.445 ;
        RECT 50.025 176.705 50.235 177.235 ;
        RECT 50.510 177.155 50.680 177.615 ;
        RECT 50.850 177.655 51.170 178.615 ;
        RECT 51.340 177.865 51.530 178.585 ;
        RECT 51.700 177.685 51.870 178.755 ;
        RECT 52.040 178.455 52.210 179.255 ;
        RECT 52.380 178.810 53.485 178.980 ;
        RECT 52.380 178.195 52.550 178.810 ;
        RECT 53.695 178.660 53.945 179.085 ;
        RECT 54.115 178.795 54.380 179.255 ;
        RECT 52.720 178.275 53.250 178.640 ;
        RECT 53.695 178.530 54.000 178.660 ;
        RECT 52.040 178.105 52.550 178.195 ;
        RECT 52.040 177.935 52.910 178.105 ;
        RECT 52.040 177.865 52.210 177.935 ;
        RECT 52.330 177.685 52.530 177.715 ;
        RECT 50.850 177.325 51.315 177.655 ;
        RECT 51.700 177.385 52.530 177.685 ;
        RECT 51.700 177.155 51.870 177.385 ;
        RECT 50.510 176.985 51.295 177.155 ;
        RECT 51.465 176.985 51.870 177.155 ;
        RECT 52.050 176.705 52.420 177.205 ;
        RECT 52.740 177.155 52.910 177.935 ;
        RECT 53.080 177.575 53.250 178.275 ;
        RECT 53.420 177.745 53.660 178.340 ;
        RECT 53.080 177.355 53.605 177.575 ;
        RECT 53.830 177.425 54.000 178.530 ;
        RECT 53.775 177.295 54.000 177.425 ;
        RECT 54.170 177.335 54.450 178.285 ;
        RECT 53.775 177.155 53.945 177.295 ;
        RECT 52.740 176.985 53.415 177.155 ;
        RECT 53.610 176.985 53.945 177.155 ;
        RECT 54.115 176.705 54.365 177.165 ;
        RECT 54.620 176.965 54.805 179.085 ;
        RECT 54.975 178.755 55.305 179.255 ;
        RECT 55.475 178.585 55.645 179.085 ;
        RECT 54.980 178.415 55.645 178.585 ;
        RECT 54.980 177.425 55.210 178.415 ;
        RECT 55.380 177.595 55.730 178.245 ;
        RECT 55.905 178.115 56.290 179.085 ;
        RECT 56.460 178.795 56.785 179.255 ;
        RECT 57.305 178.625 57.585 179.085 ;
        RECT 56.460 178.405 57.585 178.625 ;
        RECT 55.905 177.445 56.185 178.115 ;
        RECT 56.460 177.945 56.910 178.405 ;
        RECT 57.775 178.235 58.175 179.085 ;
        RECT 58.575 178.795 58.845 179.255 ;
        RECT 59.015 178.625 59.300 179.085 ;
        RECT 56.355 177.615 56.910 177.945 ;
        RECT 57.080 177.675 58.175 178.235 ;
        RECT 56.460 177.505 56.910 177.615 ;
        RECT 54.980 177.255 55.645 177.425 ;
        RECT 54.975 176.705 55.305 177.085 ;
        RECT 55.475 176.965 55.645 177.255 ;
        RECT 55.905 176.875 56.290 177.445 ;
        RECT 56.460 177.335 57.585 177.505 ;
        RECT 56.460 176.705 56.785 177.165 ;
        RECT 57.305 176.875 57.585 177.335 ;
        RECT 57.775 176.875 58.175 177.675 ;
        RECT 58.345 178.405 59.300 178.625 ;
        RECT 58.345 177.505 58.555 178.405 ;
        RECT 58.725 177.675 59.415 178.235 ;
        RECT 59.585 178.165 61.255 179.255 ;
        RECT 58.345 177.335 59.300 177.505 ;
        RECT 58.575 176.705 58.845 177.165 ;
        RECT 59.015 176.875 59.300 177.335 ;
        RECT 59.585 177.475 60.335 177.995 ;
        RECT 60.505 177.645 61.255 178.165 ;
        RECT 61.425 178.090 61.715 179.255 ;
        RECT 61.885 178.165 63.095 179.255 ;
        RECT 63.355 178.585 63.525 179.085 ;
        RECT 63.695 178.755 64.025 179.255 ;
        RECT 63.355 178.415 64.020 178.585 ;
        RECT 59.585 176.705 61.255 177.475 ;
        RECT 61.885 177.455 62.405 177.995 ;
        RECT 62.575 177.625 63.095 178.165 ;
        RECT 63.270 177.595 63.620 178.245 ;
        RECT 61.425 176.705 61.715 177.430 ;
        RECT 61.885 176.705 63.095 177.455 ;
        RECT 63.790 177.425 64.020 178.415 ;
        RECT 63.355 177.255 64.020 177.425 ;
        RECT 63.355 176.965 63.525 177.255 ;
        RECT 63.695 176.705 64.025 177.085 ;
        RECT 64.195 176.965 64.380 179.085 ;
        RECT 64.620 178.795 64.885 179.255 ;
        RECT 65.055 178.660 65.305 179.085 ;
        RECT 65.515 178.810 66.620 178.980 ;
        RECT 65.000 178.530 65.305 178.660 ;
        RECT 64.550 177.335 64.830 178.285 ;
        RECT 65.000 177.425 65.170 178.530 ;
        RECT 65.340 177.745 65.580 178.340 ;
        RECT 65.750 178.275 66.280 178.640 ;
        RECT 65.750 177.575 65.920 178.275 ;
        RECT 66.450 178.195 66.620 178.810 ;
        RECT 66.790 178.455 66.960 179.255 ;
        RECT 67.130 178.755 67.380 179.085 ;
        RECT 67.605 178.785 68.490 178.955 ;
        RECT 66.450 178.105 66.960 178.195 ;
        RECT 65.000 177.295 65.225 177.425 ;
        RECT 65.395 177.355 65.920 177.575 ;
        RECT 66.090 177.935 66.960 178.105 ;
        RECT 64.635 176.705 64.885 177.165 ;
        RECT 65.055 177.155 65.225 177.295 ;
        RECT 66.090 177.155 66.260 177.935 ;
        RECT 66.790 177.865 66.960 177.935 ;
        RECT 66.470 177.685 66.670 177.715 ;
        RECT 67.130 177.685 67.300 178.755 ;
        RECT 67.470 177.865 67.660 178.585 ;
        RECT 66.470 177.385 67.300 177.685 ;
        RECT 67.830 177.655 68.150 178.615 ;
        RECT 65.055 176.985 65.390 177.155 ;
        RECT 65.585 176.985 66.260 177.155 ;
        RECT 66.580 176.705 66.950 177.205 ;
        RECT 67.130 177.155 67.300 177.385 ;
        RECT 67.685 177.325 68.150 177.655 ;
        RECT 68.320 177.945 68.490 178.785 ;
        RECT 68.670 178.755 68.985 179.255 ;
        RECT 69.215 178.525 69.555 179.085 ;
        RECT 68.660 178.150 69.555 178.525 ;
        RECT 69.725 178.245 69.895 179.255 ;
        RECT 69.365 177.945 69.555 178.150 ;
        RECT 70.065 178.195 70.395 179.040 ;
        RECT 70.715 178.585 70.885 179.085 ;
        RECT 71.055 178.755 71.385 179.255 ;
        RECT 70.715 178.415 71.380 178.585 ;
        RECT 70.065 178.115 70.455 178.195 ;
        RECT 70.240 178.065 70.455 178.115 ;
        RECT 68.320 177.615 69.195 177.945 ;
        RECT 69.365 177.615 70.115 177.945 ;
        RECT 68.320 177.155 68.490 177.615 ;
        RECT 69.365 177.445 69.565 177.615 ;
        RECT 70.285 177.485 70.455 178.065 ;
        RECT 70.630 177.595 70.980 178.245 ;
        RECT 70.230 177.445 70.455 177.485 ;
        RECT 67.130 176.985 67.535 177.155 ;
        RECT 67.705 176.985 68.490 177.155 ;
        RECT 68.765 176.705 68.975 177.235 ;
        RECT 69.235 176.920 69.565 177.445 ;
        RECT 70.075 177.360 70.455 177.445 ;
        RECT 71.150 177.425 71.380 178.415 ;
        RECT 69.735 176.705 69.905 177.315 ;
        RECT 70.075 176.925 70.405 177.360 ;
        RECT 70.715 177.255 71.380 177.425 ;
        RECT 70.715 176.965 70.885 177.255 ;
        RECT 71.055 176.705 71.385 177.085 ;
        RECT 71.555 176.965 71.740 179.085 ;
        RECT 71.980 178.795 72.245 179.255 ;
        RECT 72.415 178.660 72.665 179.085 ;
        RECT 72.875 178.810 73.980 178.980 ;
        RECT 72.360 178.530 72.665 178.660 ;
        RECT 71.910 177.335 72.190 178.285 ;
        RECT 72.360 177.425 72.530 178.530 ;
        RECT 72.700 177.745 72.940 178.340 ;
        RECT 73.110 178.275 73.640 178.640 ;
        RECT 73.110 177.575 73.280 178.275 ;
        RECT 73.810 178.195 73.980 178.810 ;
        RECT 74.150 178.455 74.320 179.255 ;
        RECT 74.490 178.755 74.740 179.085 ;
        RECT 74.965 178.785 75.850 178.955 ;
        RECT 73.810 178.105 74.320 178.195 ;
        RECT 72.360 177.295 72.585 177.425 ;
        RECT 72.755 177.355 73.280 177.575 ;
        RECT 73.450 177.935 74.320 178.105 ;
        RECT 71.995 176.705 72.245 177.165 ;
        RECT 72.415 177.155 72.585 177.295 ;
        RECT 73.450 177.155 73.620 177.935 ;
        RECT 74.150 177.865 74.320 177.935 ;
        RECT 73.830 177.685 74.030 177.715 ;
        RECT 74.490 177.685 74.660 178.755 ;
        RECT 74.830 177.865 75.020 178.585 ;
        RECT 73.830 177.385 74.660 177.685 ;
        RECT 75.190 177.655 75.510 178.615 ;
        RECT 72.415 176.985 72.750 177.155 ;
        RECT 72.945 176.985 73.620 177.155 ;
        RECT 73.940 176.705 74.310 177.205 ;
        RECT 74.490 177.155 74.660 177.385 ;
        RECT 75.045 177.325 75.510 177.655 ;
        RECT 75.680 177.945 75.850 178.785 ;
        RECT 76.030 178.755 76.345 179.255 ;
        RECT 76.575 178.525 76.915 179.085 ;
        RECT 76.020 178.150 76.915 178.525 ;
        RECT 77.085 178.245 77.255 179.255 ;
        RECT 76.725 177.945 76.915 178.150 ;
        RECT 77.425 178.195 77.755 179.040 ;
        RECT 77.425 178.115 77.815 178.195 ;
        RECT 77.985 178.165 79.655 179.255 ;
        RECT 79.915 178.585 80.085 179.085 ;
        RECT 80.255 178.755 80.585 179.255 ;
        RECT 79.915 178.415 80.580 178.585 ;
        RECT 77.600 178.065 77.815 178.115 ;
        RECT 75.680 177.615 76.555 177.945 ;
        RECT 76.725 177.615 77.475 177.945 ;
        RECT 75.680 177.155 75.850 177.615 ;
        RECT 76.725 177.445 76.925 177.615 ;
        RECT 77.645 177.485 77.815 178.065 ;
        RECT 77.590 177.445 77.815 177.485 ;
        RECT 74.490 176.985 74.895 177.155 ;
        RECT 75.065 176.985 75.850 177.155 ;
        RECT 76.125 176.705 76.335 177.235 ;
        RECT 76.595 176.920 76.925 177.445 ;
        RECT 77.435 177.360 77.815 177.445 ;
        RECT 77.985 177.475 78.735 177.995 ;
        RECT 78.905 177.645 79.655 178.165 ;
        RECT 79.830 177.595 80.180 178.245 ;
        RECT 77.095 176.705 77.265 177.315 ;
        RECT 77.435 176.925 77.765 177.360 ;
        RECT 77.985 176.705 79.655 177.475 ;
        RECT 80.350 177.425 80.580 178.415 ;
        RECT 79.915 177.255 80.580 177.425 ;
        RECT 79.915 176.965 80.085 177.255 ;
        RECT 80.255 176.705 80.585 177.085 ;
        RECT 80.755 176.965 80.940 179.085 ;
        RECT 81.180 178.795 81.445 179.255 ;
        RECT 81.615 178.660 81.865 179.085 ;
        RECT 82.075 178.810 83.180 178.980 ;
        RECT 81.560 178.530 81.865 178.660 ;
        RECT 81.110 177.335 81.390 178.285 ;
        RECT 81.560 177.425 81.730 178.530 ;
        RECT 81.900 177.745 82.140 178.340 ;
        RECT 82.310 178.275 82.840 178.640 ;
        RECT 82.310 177.575 82.480 178.275 ;
        RECT 83.010 178.195 83.180 178.810 ;
        RECT 83.350 178.455 83.520 179.255 ;
        RECT 83.690 178.755 83.940 179.085 ;
        RECT 84.165 178.785 85.050 178.955 ;
        RECT 83.010 178.105 83.520 178.195 ;
        RECT 81.560 177.295 81.785 177.425 ;
        RECT 81.955 177.355 82.480 177.575 ;
        RECT 82.650 177.935 83.520 178.105 ;
        RECT 81.195 176.705 81.445 177.165 ;
        RECT 81.615 177.155 81.785 177.295 ;
        RECT 82.650 177.155 82.820 177.935 ;
        RECT 83.350 177.865 83.520 177.935 ;
        RECT 83.030 177.685 83.230 177.715 ;
        RECT 83.690 177.685 83.860 178.755 ;
        RECT 84.030 177.865 84.220 178.585 ;
        RECT 83.030 177.385 83.860 177.685 ;
        RECT 84.390 177.655 84.710 178.615 ;
        RECT 81.615 176.985 81.950 177.155 ;
        RECT 82.145 176.985 82.820 177.155 ;
        RECT 83.140 176.705 83.510 177.205 ;
        RECT 83.690 177.155 83.860 177.385 ;
        RECT 84.245 177.325 84.710 177.655 ;
        RECT 84.880 177.945 85.050 178.785 ;
        RECT 85.230 178.755 85.545 179.255 ;
        RECT 85.775 178.525 86.115 179.085 ;
        RECT 85.220 178.150 86.115 178.525 ;
        RECT 86.285 178.245 86.455 179.255 ;
        RECT 85.925 177.945 86.115 178.150 ;
        RECT 86.625 178.195 86.955 179.040 ;
        RECT 86.625 178.115 87.015 178.195 ;
        RECT 86.800 178.065 87.015 178.115 ;
        RECT 87.185 178.090 87.475 179.255 ;
        RECT 88.220 178.625 88.505 179.085 ;
        RECT 88.675 178.795 88.945 179.255 ;
        RECT 88.220 178.405 89.175 178.625 ;
        RECT 84.880 177.615 85.755 177.945 ;
        RECT 85.925 177.615 86.675 177.945 ;
        RECT 84.880 177.155 85.050 177.615 ;
        RECT 85.925 177.445 86.125 177.615 ;
        RECT 86.845 177.485 87.015 178.065 ;
        RECT 88.105 177.675 88.795 178.235 ;
        RECT 88.965 177.505 89.175 178.405 ;
        RECT 86.790 177.445 87.015 177.485 ;
        RECT 83.690 176.985 84.095 177.155 ;
        RECT 84.265 176.985 85.050 177.155 ;
        RECT 85.325 176.705 85.535 177.235 ;
        RECT 85.795 176.920 86.125 177.445 ;
        RECT 86.635 177.360 87.015 177.445 ;
        RECT 86.295 176.705 86.465 177.315 ;
        RECT 86.635 176.925 86.965 177.360 ;
        RECT 87.185 176.705 87.475 177.430 ;
        RECT 88.220 177.335 89.175 177.505 ;
        RECT 89.345 178.235 89.745 179.085 ;
        RECT 89.935 178.625 90.215 179.085 ;
        RECT 90.735 178.795 91.060 179.255 ;
        RECT 89.935 178.405 91.060 178.625 ;
        RECT 89.345 177.675 90.440 178.235 ;
        RECT 90.610 177.945 91.060 178.405 ;
        RECT 91.230 178.115 91.615 179.085 ;
        RECT 88.220 176.875 88.505 177.335 ;
        RECT 88.675 176.705 88.945 177.165 ;
        RECT 89.345 176.875 89.745 177.675 ;
        RECT 90.610 177.615 91.165 177.945 ;
        RECT 90.610 177.505 91.060 177.615 ;
        RECT 89.935 177.335 91.060 177.505 ;
        RECT 91.335 177.445 91.615 178.115 ;
        RECT 89.935 176.875 90.215 177.335 ;
        RECT 90.735 176.705 91.060 177.165 ;
        RECT 91.230 176.875 91.615 177.445 ;
        RECT 91.785 178.385 92.060 179.085 ;
        RECT 92.230 178.710 92.485 179.255 ;
        RECT 92.655 178.745 93.135 179.085 ;
        RECT 93.310 178.700 93.915 179.255 ;
        RECT 93.300 178.600 93.915 178.700 ;
        RECT 93.300 178.575 93.485 178.600 ;
        RECT 91.785 177.355 91.955 178.385 ;
        RECT 92.230 178.255 92.985 178.505 ;
        RECT 93.155 178.330 93.485 178.575 ;
        RECT 92.230 178.220 93.000 178.255 ;
        RECT 92.230 178.210 93.015 178.220 ;
        RECT 92.125 178.195 93.020 178.210 ;
        RECT 92.125 178.180 93.040 178.195 ;
        RECT 92.125 178.170 93.060 178.180 ;
        RECT 92.125 178.160 93.085 178.170 ;
        RECT 92.125 178.130 93.155 178.160 ;
        RECT 92.125 178.100 93.175 178.130 ;
        RECT 92.125 178.070 93.195 178.100 ;
        RECT 92.125 178.045 93.225 178.070 ;
        RECT 92.125 178.010 93.260 178.045 ;
        RECT 92.125 178.005 93.290 178.010 ;
        RECT 92.125 177.610 92.355 178.005 ;
        RECT 92.900 178.000 93.290 178.005 ;
        RECT 92.925 177.990 93.290 178.000 ;
        RECT 92.940 177.985 93.290 177.990 ;
        RECT 92.955 177.980 93.290 177.985 ;
        RECT 93.655 177.980 93.915 178.430 ;
        RECT 92.955 177.975 93.915 177.980 ;
        RECT 92.965 177.965 93.915 177.975 ;
        RECT 92.975 177.960 93.915 177.965 ;
        RECT 92.985 177.950 93.915 177.960 ;
        RECT 92.990 177.940 93.915 177.950 ;
        RECT 92.995 177.935 93.915 177.940 ;
        RECT 93.005 177.920 93.915 177.935 ;
        RECT 93.010 177.905 93.915 177.920 ;
        RECT 93.020 177.880 93.915 177.905 ;
        RECT 92.525 177.410 92.855 177.835 ;
        RECT 91.785 176.875 92.045 177.355 ;
        RECT 92.215 176.705 92.465 177.245 ;
        RECT 92.635 176.925 92.855 177.410 ;
        RECT 93.025 177.810 93.915 177.880 ;
        RECT 94.085 178.180 94.355 179.085 ;
        RECT 94.525 178.495 94.855 179.255 ;
        RECT 95.035 178.325 95.205 179.085 ;
        RECT 93.025 177.085 93.195 177.810 ;
        RECT 93.365 177.255 93.915 177.640 ;
        RECT 94.085 177.380 94.255 178.180 ;
        RECT 94.540 178.155 95.205 178.325 ;
        RECT 95.465 178.535 95.925 179.085 ;
        RECT 96.115 178.535 96.445 179.255 ;
        RECT 94.540 178.010 94.710 178.155 ;
        RECT 94.425 177.680 94.710 178.010 ;
        RECT 94.540 177.425 94.710 177.680 ;
        RECT 94.945 177.605 95.275 177.975 ;
        RECT 93.025 176.915 93.915 177.085 ;
        RECT 94.085 176.875 94.345 177.380 ;
        RECT 94.540 177.255 95.205 177.425 ;
        RECT 94.525 176.705 94.855 177.085 ;
        RECT 95.035 176.875 95.205 177.255 ;
        RECT 95.465 177.165 95.715 178.535 ;
        RECT 96.645 178.365 96.945 178.915 ;
        RECT 97.115 178.585 97.395 179.255 ;
        RECT 96.005 178.195 96.945 178.365 ;
        RECT 98.315 178.325 98.485 179.085 ;
        RECT 98.665 178.495 98.995 179.255 ;
        RECT 96.005 177.945 96.175 178.195 ;
        RECT 97.315 177.945 97.580 178.305 ;
        RECT 98.315 178.155 98.980 178.325 ;
        RECT 99.165 178.180 99.435 179.085 ;
        RECT 99.695 178.585 99.865 179.085 ;
        RECT 100.035 178.755 100.365 179.255 ;
        RECT 99.695 178.415 100.360 178.585 ;
        RECT 98.810 178.010 98.980 178.155 ;
        RECT 95.885 177.615 96.175 177.945 ;
        RECT 96.345 177.695 96.685 177.945 ;
        RECT 96.905 177.695 97.580 177.945 ;
        RECT 96.005 177.525 96.175 177.615 ;
        RECT 98.245 177.605 98.575 177.975 ;
        RECT 98.810 177.680 99.095 178.010 ;
        RECT 96.005 177.335 97.395 177.525 ;
        RECT 98.810 177.425 98.980 177.680 ;
        RECT 95.465 176.875 96.025 177.165 ;
        RECT 96.195 176.705 96.445 177.165 ;
        RECT 97.065 176.975 97.395 177.335 ;
        RECT 98.315 177.255 98.980 177.425 ;
        RECT 99.265 177.380 99.435 178.180 ;
        RECT 99.610 177.595 99.960 178.245 ;
        RECT 100.130 177.425 100.360 178.415 ;
        RECT 98.315 176.875 98.485 177.255 ;
        RECT 98.665 176.705 98.995 177.085 ;
        RECT 99.175 176.875 99.435 177.380 ;
        RECT 99.695 177.255 100.360 177.425 ;
        RECT 99.695 176.965 99.865 177.255 ;
        RECT 100.035 176.705 100.365 177.085 ;
        RECT 100.535 176.965 100.720 179.085 ;
        RECT 100.960 178.795 101.225 179.255 ;
        RECT 101.395 178.660 101.645 179.085 ;
        RECT 101.855 178.810 102.960 178.980 ;
        RECT 101.340 178.530 101.645 178.660 ;
        RECT 100.890 177.335 101.170 178.285 ;
        RECT 101.340 177.425 101.510 178.530 ;
        RECT 101.680 177.745 101.920 178.340 ;
        RECT 102.090 178.275 102.620 178.640 ;
        RECT 102.090 177.575 102.260 178.275 ;
        RECT 102.790 178.195 102.960 178.810 ;
        RECT 103.130 178.455 103.300 179.255 ;
        RECT 103.470 178.755 103.720 179.085 ;
        RECT 103.945 178.785 104.830 178.955 ;
        RECT 102.790 178.105 103.300 178.195 ;
        RECT 101.340 177.295 101.565 177.425 ;
        RECT 101.735 177.355 102.260 177.575 ;
        RECT 102.430 177.935 103.300 178.105 ;
        RECT 100.975 176.705 101.225 177.165 ;
        RECT 101.395 177.155 101.565 177.295 ;
        RECT 102.430 177.155 102.600 177.935 ;
        RECT 103.130 177.865 103.300 177.935 ;
        RECT 102.810 177.685 103.010 177.715 ;
        RECT 103.470 177.685 103.640 178.755 ;
        RECT 103.810 177.865 104.000 178.585 ;
        RECT 102.810 177.385 103.640 177.685 ;
        RECT 104.170 177.655 104.490 178.615 ;
        RECT 101.395 176.985 101.730 177.155 ;
        RECT 101.925 176.985 102.600 177.155 ;
        RECT 102.920 176.705 103.290 177.205 ;
        RECT 103.470 177.155 103.640 177.385 ;
        RECT 104.025 177.325 104.490 177.655 ;
        RECT 104.660 177.945 104.830 178.785 ;
        RECT 105.010 178.755 105.325 179.255 ;
        RECT 105.555 178.525 105.895 179.085 ;
        RECT 105.000 178.150 105.895 178.525 ;
        RECT 106.065 178.245 106.235 179.255 ;
        RECT 105.705 177.945 105.895 178.150 ;
        RECT 106.405 178.195 106.735 179.040 ;
        RECT 106.965 178.535 107.425 179.085 ;
        RECT 107.615 178.535 107.945 179.255 ;
        RECT 106.405 178.115 106.795 178.195 ;
        RECT 106.580 178.065 106.795 178.115 ;
        RECT 104.660 177.615 105.535 177.945 ;
        RECT 105.705 177.615 106.455 177.945 ;
        RECT 104.660 177.155 104.830 177.615 ;
        RECT 105.705 177.445 105.905 177.615 ;
        RECT 106.625 177.485 106.795 178.065 ;
        RECT 106.570 177.445 106.795 177.485 ;
        RECT 103.470 176.985 103.875 177.155 ;
        RECT 104.045 176.985 104.830 177.155 ;
        RECT 105.105 176.705 105.315 177.235 ;
        RECT 105.575 176.920 105.905 177.445 ;
        RECT 106.415 177.360 106.795 177.445 ;
        RECT 106.075 176.705 106.245 177.315 ;
        RECT 106.415 176.925 106.745 177.360 ;
        RECT 106.965 177.165 107.215 178.535 ;
        RECT 108.145 178.365 108.445 178.915 ;
        RECT 108.615 178.585 108.895 179.255 ;
        RECT 109.765 178.915 110.905 179.085 ;
        RECT 109.765 178.455 110.065 178.915 ;
        RECT 107.505 178.195 108.445 178.365 ;
        RECT 107.505 177.945 107.675 178.195 ;
        RECT 108.815 177.945 109.080 178.305 ;
        RECT 110.235 178.285 110.565 178.745 ;
        RECT 107.385 177.615 107.675 177.945 ;
        RECT 107.845 177.695 108.185 177.945 ;
        RECT 108.405 177.695 109.080 177.945 ;
        RECT 109.805 178.065 110.565 178.285 ;
        RECT 110.735 178.285 110.905 178.915 ;
        RECT 111.075 178.455 111.405 179.255 ;
        RECT 111.575 178.285 111.850 179.085 ;
        RECT 110.735 178.075 111.850 178.285 ;
        RECT 112.945 178.090 113.235 179.255 ;
        RECT 113.405 178.165 115.075 179.255 ;
        RECT 107.505 177.525 107.675 177.615 ;
        RECT 109.805 177.525 110.020 178.065 ;
        RECT 110.190 177.695 110.960 177.895 ;
        RECT 111.130 177.695 111.850 177.895 ;
        RECT 107.505 177.335 108.895 177.525 ;
        RECT 109.805 177.355 111.405 177.525 ;
        RECT 106.965 176.875 107.525 177.165 ;
        RECT 107.695 176.705 107.945 177.165 ;
        RECT 108.565 176.975 108.895 177.335 ;
        RECT 110.235 177.345 111.405 177.355 ;
        RECT 109.775 176.705 110.065 177.175 ;
        RECT 110.235 176.875 110.565 177.345 ;
        RECT 110.735 176.705 110.905 177.175 ;
        RECT 111.075 176.875 111.405 177.345 ;
        RECT 111.575 176.705 111.850 177.525 ;
        RECT 113.405 177.475 114.155 177.995 ;
        RECT 114.325 177.645 115.075 178.165 ;
        RECT 115.335 178.325 115.505 179.085 ;
        RECT 115.685 178.495 116.015 179.255 ;
        RECT 115.335 178.155 116.000 178.325 ;
        RECT 116.185 178.180 116.455 179.085 ;
        RECT 116.715 178.585 116.885 179.085 ;
        RECT 117.055 178.755 117.385 179.255 ;
        RECT 116.715 178.415 117.380 178.585 ;
        RECT 115.830 178.010 116.000 178.155 ;
        RECT 115.265 177.605 115.595 177.975 ;
        RECT 115.830 177.680 116.115 178.010 ;
        RECT 112.945 176.705 113.235 177.430 ;
        RECT 113.405 176.705 115.075 177.475 ;
        RECT 115.830 177.425 116.000 177.680 ;
        RECT 115.335 177.255 116.000 177.425 ;
        RECT 116.285 177.380 116.455 178.180 ;
        RECT 116.630 177.595 116.980 178.245 ;
        RECT 117.150 177.425 117.380 178.415 ;
        RECT 115.335 176.875 115.505 177.255 ;
        RECT 115.685 176.705 116.015 177.085 ;
        RECT 116.195 176.875 116.455 177.380 ;
        RECT 116.715 177.255 117.380 177.425 ;
        RECT 116.715 176.965 116.885 177.255 ;
        RECT 117.055 176.705 117.385 177.085 ;
        RECT 117.555 176.965 117.740 179.085 ;
        RECT 117.980 178.795 118.245 179.255 ;
        RECT 118.415 178.660 118.665 179.085 ;
        RECT 118.875 178.810 119.980 178.980 ;
        RECT 118.360 178.530 118.665 178.660 ;
        RECT 117.910 177.335 118.190 178.285 ;
        RECT 118.360 177.425 118.530 178.530 ;
        RECT 118.700 177.745 118.940 178.340 ;
        RECT 119.110 178.275 119.640 178.640 ;
        RECT 119.110 177.575 119.280 178.275 ;
        RECT 119.810 178.195 119.980 178.810 ;
        RECT 120.150 178.455 120.320 179.255 ;
        RECT 120.490 178.755 120.740 179.085 ;
        RECT 120.965 178.785 121.850 178.955 ;
        RECT 119.810 178.105 120.320 178.195 ;
        RECT 118.360 177.295 118.585 177.425 ;
        RECT 118.755 177.355 119.280 177.575 ;
        RECT 119.450 177.935 120.320 178.105 ;
        RECT 117.995 176.705 118.245 177.165 ;
        RECT 118.415 177.155 118.585 177.295 ;
        RECT 119.450 177.155 119.620 177.935 ;
        RECT 120.150 177.865 120.320 177.935 ;
        RECT 119.830 177.685 120.030 177.715 ;
        RECT 120.490 177.685 120.660 178.755 ;
        RECT 120.830 177.865 121.020 178.585 ;
        RECT 119.830 177.385 120.660 177.685 ;
        RECT 121.190 177.655 121.510 178.615 ;
        RECT 118.415 176.985 118.750 177.155 ;
        RECT 118.945 176.985 119.620 177.155 ;
        RECT 119.940 176.705 120.310 177.205 ;
        RECT 120.490 177.155 120.660 177.385 ;
        RECT 121.045 177.325 121.510 177.655 ;
        RECT 121.680 177.945 121.850 178.785 ;
        RECT 122.030 178.755 122.345 179.255 ;
        RECT 122.575 178.525 122.915 179.085 ;
        RECT 122.020 178.150 122.915 178.525 ;
        RECT 123.085 178.245 123.255 179.255 ;
        RECT 122.725 177.945 122.915 178.150 ;
        RECT 123.425 178.195 123.755 179.040 ;
        RECT 123.425 178.115 123.815 178.195 ;
        RECT 123.985 178.165 127.495 179.255 ;
        RECT 128.215 178.635 128.385 179.065 ;
        RECT 128.555 178.805 128.885 179.255 ;
        RECT 128.215 178.405 128.890 178.635 ;
        RECT 123.600 178.065 123.815 178.115 ;
        RECT 121.680 177.615 122.555 177.945 ;
        RECT 122.725 177.615 123.475 177.945 ;
        RECT 121.680 177.155 121.850 177.615 ;
        RECT 122.725 177.445 122.925 177.615 ;
        RECT 123.645 177.485 123.815 178.065 ;
        RECT 123.590 177.445 123.815 177.485 ;
        RECT 120.490 176.985 120.895 177.155 ;
        RECT 121.065 176.985 121.850 177.155 ;
        RECT 122.125 176.705 122.335 177.235 ;
        RECT 122.595 176.920 122.925 177.445 ;
        RECT 123.435 177.360 123.815 177.445 ;
        RECT 123.985 177.475 125.635 177.995 ;
        RECT 125.805 177.645 127.495 178.165 ;
        RECT 123.095 176.705 123.265 177.315 ;
        RECT 123.435 176.925 123.765 177.360 ;
        RECT 123.985 176.705 127.495 177.475 ;
        RECT 128.185 177.385 128.485 178.235 ;
        RECT 128.655 177.755 128.890 178.405 ;
        RECT 129.060 178.095 129.345 179.040 ;
        RECT 129.525 178.785 130.210 179.255 ;
        RECT 129.520 178.265 130.215 178.575 ;
        RECT 130.390 178.200 130.695 178.985 ;
        RECT 129.060 177.945 129.920 178.095 ;
        RECT 129.060 177.925 130.345 177.945 ;
        RECT 128.655 177.425 129.190 177.755 ;
        RECT 129.360 177.565 130.345 177.925 ;
        RECT 128.655 177.275 128.875 177.425 ;
        RECT 128.130 176.705 128.465 177.210 ;
        RECT 128.635 176.900 128.875 177.275 ;
        RECT 129.360 177.230 129.530 177.565 ;
        RECT 130.520 177.395 130.695 178.200 ;
        RECT 130.885 178.165 134.395 179.255 ;
        RECT 129.155 177.035 129.530 177.230 ;
        RECT 129.155 176.890 129.325 177.035 ;
        RECT 129.890 176.705 130.285 177.200 ;
        RECT 130.455 176.875 130.695 177.395 ;
        RECT 130.885 177.475 132.535 177.995 ;
        RECT 132.705 177.645 134.395 178.165 ;
        RECT 135.025 178.115 135.285 179.255 ;
        RECT 135.525 178.745 137.140 179.075 ;
        RECT 135.535 177.945 135.705 178.505 ;
        RECT 135.965 178.405 137.140 178.575 ;
        RECT 137.310 178.455 137.590 179.255 ;
        RECT 135.965 178.115 136.295 178.405 ;
        RECT 136.970 178.285 137.140 178.405 ;
        RECT 136.465 177.945 136.710 178.235 ;
        RECT 136.970 178.115 137.630 178.285 ;
        RECT 137.800 178.115 138.075 179.085 ;
        RECT 137.460 177.945 137.630 178.115 ;
        RECT 135.030 177.695 135.365 177.945 ;
        RECT 135.535 177.615 136.250 177.945 ;
        RECT 136.465 177.615 137.290 177.945 ;
        RECT 137.460 177.615 137.735 177.945 ;
        RECT 135.535 177.525 135.785 177.615 ;
        RECT 130.885 176.705 134.395 177.475 ;
        RECT 135.025 176.705 135.285 177.525 ;
        RECT 135.455 177.105 135.785 177.525 ;
        RECT 137.460 177.445 137.630 177.615 ;
        RECT 135.965 177.275 137.630 177.445 ;
        RECT 137.905 177.380 138.075 178.115 ;
        RECT 138.705 178.090 138.995 179.255 ;
        RECT 139.165 178.700 139.770 179.255 ;
        RECT 139.945 178.745 140.425 179.085 ;
        RECT 140.595 178.710 140.850 179.255 ;
        RECT 139.165 178.600 139.780 178.700 ;
        RECT 139.595 178.575 139.780 178.600 ;
        RECT 139.165 177.980 139.425 178.430 ;
        RECT 139.595 178.330 139.925 178.575 ;
        RECT 140.095 178.255 140.850 178.505 ;
        RECT 141.020 178.385 141.295 179.085 ;
        RECT 140.080 178.220 140.850 178.255 ;
        RECT 140.065 178.210 140.850 178.220 ;
        RECT 140.060 178.195 140.955 178.210 ;
        RECT 140.040 178.180 140.955 178.195 ;
        RECT 140.020 178.170 140.955 178.180 ;
        RECT 139.995 178.160 140.955 178.170 ;
        RECT 139.925 178.130 140.955 178.160 ;
        RECT 139.905 178.100 140.955 178.130 ;
        RECT 139.885 178.070 140.955 178.100 ;
        RECT 139.855 178.045 140.955 178.070 ;
        RECT 139.820 178.010 140.955 178.045 ;
        RECT 139.790 178.005 140.955 178.010 ;
        RECT 139.790 178.000 140.180 178.005 ;
        RECT 139.790 177.990 140.155 178.000 ;
        RECT 139.790 177.985 140.140 177.990 ;
        RECT 139.790 177.980 140.125 177.985 ;
        RECT 139.165 177.975 140.125 177.980 ;
        RECT 139.165 177.965 140.115 177.975 ;
        RECT 139.165 177.960 140.105 177.965 ;
        RECT 139.165 177.950 140.095 177.960 ;
        RECT 139.165 177.940 140.090 177.950 ;
        RECT 139.165 177.935 140.085 177.940 ;
        RECT 139.165 177.920 140.075 177.935 ;
        RECT 139.165 177.905 140.070 177.920 ;
        RECT 139.165 177.880 140.060 177.905 ;
        RECT 139.165 177.810 140.055 177.880 ;
        RECT 135.965 176.875 136.225 177.275 ;
        RECT 136.395 176.705 136.725 177.105 ;
        RECT 136.895 176.925 137.065 177.275 ;
        RECT 137.235 176.705 137.610 177.105 ;
        RECT 137.800 177.035 138.075 177.380 ;
        RECT 138.705 176.705 138.995 177.430 ;
        RECT 139.165 177.255 139.715 177.640 ;
        RECT 139.885 177.085 140.055 177.810 ;
        RECT 139.165 176.915 140.055 177.085 ;
        RECT 140.225 177.410 140.555 177.835 ;
        RECT 140.725 177.610 140.955 178.005 ;
        RECT 140.225 176.925 140.445 177.410 ;
        RECT 141.125 177.355 141.295 178.385 ;
        RECT 141.505 178.115 141.735 179.255 ;
        RECT 141.905 178.105 142.235 179.085 ;
        RECT 142.405 178.115 142.615 179.255 ;
        RECT 142.935 178.325 143.105 179.085 ;
        RECT 143.285 178.495 143.615 179.255 ;
        RECT 142.935 178.155 143.600 178.325 ;
        RECT 143.785 178.180 144.055 179.085 ;
        RECT 141.485 177.695 141.815 177.945 ;
        RECT 140.615 176.705 140.865 177.245 ;
        RECT 141.035 176.875 141.295 177.355 ;
        RECT 141.505 176.705 141.735 177.525 ;
        RECT 141.985 177.505 142.235 178.105 ;
        RECT 143.430 178.010 143.600 178.155 ;
        RECT 142.865 177.605 143.195 177.975 ;
        RECT 143.430 177.680 143.715 178.010 ;
        RECT 141.905 176.875 142.235 177.505 ;
        RECT 142.405 176.705 142.615 177.525 ;
        RECT 143.430 177.425 143.600 177.680 ;
        RECT 142.935 177.255 143.600 177.425 ;
        RECT 143.885 177.380 144.055 178.180 ;
        RECT 144.225 178.115 144.505 179.255 ;
        RECT 144.675 178.105 145.005 179.085 ;
        RECT 145.175 178.115 145.435 179.255 ;
        RECT 145.605 178.115 145.885 179.255 ;
        RECT 146.055 178.105 146.385 179.085 ;
        RECT 146.555 178.115 146.815 179.255 ;
        RECT 146.985 178.165 148.195 179.255 ;
        RECT 148.455 178.585 148.625 179.085 ;
        RECT 148.795 178.755 149.125 179.255 ;
        RECT 148.455 178.415 149.120 178.585 ;
        RECT 144.235 177.675 144.570 177.945 ;
        RECT 144.740 177.505 144.910 178.105 ;
        RECT 145.080 177.695 145.415 177.945 ;
        RECT 145.615 177.675 145.950 177.945 ;
        RECT 146.120 177.505 146.290 178.105 ;
        RECT 146.460 177.695 146.795 177.945 ;
        RECT 142.935 176.875 143.105 177.255 ;
        RECT 143.285 176.705 143.615 177.085 ;
        RECT 143.795 176.875 144.055 177.380 ;
        RECT 144.225 176.705 144.535 177.505 ;
        RECT 144.740 176.875 145.435 177.505 ;
        RECT 145.605 176.705 145.915 177.505 ;
        RECT 146.120 176.875 146.815 177.505 ;
        RECT 146.985 177.455 147.505 177.995 ;
        RECT 147.675 177.625 148.195 178.165 ;
        RECT 148.370 177.595 148.720 178.245 ;
        RECT 146.985 176.705 148.195 177.455 ;
        RECT 148.890 177.425 149.120 178.415 ;
        RECT 148.455 177.255 149.120 177.425 ;
        RECT 148.455 176.965 148.625 177.255 ;
        RECT 148.795 176.705 149.125 177.085 ;
        RECT 149.295 176.965 149.480 179.085 ;
        RECT 149.720 178.795 149.985 179.255 ;
        RECT 150.155 178.660 150.405 179.085 ;
        RECT 150.615 178.810 151.720 178.980 ;
        RECT 150.100 178.530 150.405 178.660 ;
        RECT 149.650 177.335 149.930 178.285 ;
        RECT 150.100 177.425 150.270 178.530 ;
        RECT 150.440 177.745 150.680 178.340 ;
        RECT 150.850 178.275 151.380 178.640 ;
        RECT 150.850 177.575 151.020 178.275 ;
        RECT 151.550 178.195 151.720 178.810 ;
        RECT 151.890 178.455 152.060 179.255 ;
        RECT 152.230 178.755 152.480 179.085 ;
        RECT 152.705 178.785 153.590 178.955 ;
        RECT 151.550 178.105 152.060 178.195 ;
        RECT 150.100 177.295 150.325 177.425 ;
        RECT 150.495 177.355 151.020 177.575 ;
        RECT 151.190 177.935 152.060 178.105 ;
        RECT 149.735 176.705 149.985 177.165 ;
        RECT 150.155 177.155 150.325 177.295 ;
        RECT 151.190 177.155 151.360 177.935 ;
        RECT 151.890 177.865 152.060 177.935 ;
        RECT 151.570 177.685 151.770 177.715 ;
        RECT 152.230 177.685 152.400 178.755 ;
        RECT 152.570 177.865 152.760 178.585 ;
        RECT 151.570 177.385 152.400 177.685 ;
        RECT 152.930 177.655 153.250 178.615 ;
        RECT 150.155 176.985 150.490 177.155 ;
        RECT 150.685 176.985 151.360 177.155 ;
        RECT 151.680 176.705 152.050 177.205 ;
        RECT 152.230 177.155 152.400 177.385 ;
        RECT 152.785 177.325 153.250 177.655 ;
        RECT 153.420 177.945 153.590 178.785 ;
        RECT 153.770 178.755 154.085 179.255 ;
        RECT 154.315 178.525 154.655 179.085 ;
        RECT 153.760 178.150 154.655 178.525 ;
        RECT 154.825 178.245 154.995 179.255 ;
        RECT 154.465 177.945 154.655 178.150 ;
        RECT 155.165 178.195 155.495 179.040 ;
        RECT 155.165 178.115 155.555 178.195 ;
        RECT 155.340 178.065 155.555 178.115 ;
        RECT 153.420 177.615 154.295 177.945 ;
        RECT 154.465 177.615 155.215 177.945 ;
        RECT 153.420 177.155 153.590 177.615 ;
        RECT 154.465 177.445 154.665 177.615 ;
        RECT 155.385 177.485 155.555 178.065 ;
        RECT 155.725 178.165 156.935 179.255 ;
        RECT 155.725 177.625 156.245 178.165 ;
        RECT 155.330 177.445 155.555 177.485 ;
        RECT 156.415 177.455 156.935 177.995 ;
        RECT 152.230 176.985 152.635 177.155 ;
        RECT 152.805 176.985 153.590 177.155 ;
        RECT 153.865 176.705 154.075 177.235 ;
        RECT 154.335 176.920 154.665 177.445 ;
        RECT 155.175 177.360 155.555 177.445 ;
        RECT 154.835 176.705 155.005 177.315 ;
        RECT 155.175 176.925 155.505 177.360 ;
        RECT 155.725 176.705 156.935 177.455 ;
        RECT 22.700 176.535 157.020 176.705 ;
        RECT 22.785 175.785 23.995 176.535 ;
        RECT 22.785 175.245 23.305 175.785 ;
        RECT 24.165 175.765 27.675 176.535 ;
        RECT 23.475 175.075 23.995 175.615 ;
        RECT 24.165 175.245 25.815 175.765 ;
        RECT 28.765 175.735 29.460 176.365 ;
        RECT 29.665 175.735 29.975 176.535 ;
        RECT 30.145 176.075 30.705 176.365 ;
        RECT 30.875 176.075 31.125 176.535 ;
        RECT 25.985 175.075 27.675 175.595 ;
        RECT 28.785 175.295 29.120 175.545 ;
        RECT 29.290 175.135 29.460 175.735 ;
        RECT 29.630 175.295 29.965 175.565 ;
        RECT 22.785 173.985 23.995 175.075 ;
        RECT 24.165 173.985 27.675 175.075 ;
        RECT 28.765 173.985 29.025 175.125 ;
        RECT 29.195 174.155 29.525 175.135 ;
        RECT 29.695 173.985 29.975 175.125 ;
        RECT 30.145 174.705 30.395 176.075 ;
        RECT 31.745 175.905 32.075 176.265 ;
        RECT 30.685 175.715 32.075 175.905 ;
        RECT 33.425 175.715 33.635 176.535 ;
        RECT 33.805 175.735 34.135 176.365 ;
        RECT 30.685 175.625 30.855 175.715 ;
        RECT 30.565 175.295 30.855 175.625 ;
        RECT 31.025 175.295 31.365 175.545 ;
        RECT 31.585 175.295 32.260 175.545 ;
        RECT 30.685 175.045 30.855 175.295 ;
        RECT 30.685 174.875 31.625 175.045 ;
        RECT 31.995 174.935 32.260 175.295 ;
        RECT 33.805 175.135 34.055 175.735 ;
        RECT 34.305 175.715 34.535 176.535 ;
        RECT 34.745 175.990 40.090 176.535 ;
        RECT 34.225 175.295 34.555 175.545 ;
        RECT 36.330 175.160 36.670 175.990 ;
        RECT 40.265 175.785 41.475 176.535 ;
        RECT 41.645 175.860 41.915 176.205 ;
        RECT 42.105 176.135 42.485 176.535 ;
        RECT 42.655 175.965 42.825 176.315 ;
        RECT 42.995 176.055 43.730 176.535 ;
        RECT 30.145 174.155 30.605 174.705 ;
        RECT 30.795 173.985 31.125 174.705 ;
        RECT 31.325 174.325 31.625 174.875 ;
        RECT 31.795 173.985 32.075 174.655 ;
        RECT 33.425 173.985 33.635 175.125 ;
        RECT 33.805 174.155 34.135 175.135 ;
        RECT 34.305 173.985 34.535 175.125 ;
        RECT 38.150 174.420 38.500 175.670 ;
        RECT 40.265 175.245 40.785 175.785 ;
        RECT 40.955 175.075 41.475 175.615 ;
        RECT 34.745 173.985 40.090 174.420 ;
        RECT 40.265 173.985 41.475 175.075 ;
        RECT 41.645 175.125 41.815 175.860 ;
        RECT 42.085 175.795 42.825 175.965 ;
        RECT 43.900 175.885 44.210 176.355 ;
        RECT 42.085 175.625 42.255 175.795 ;
        RECT 43.475 175.715 44.210 175.885 ;
        RECT 44.405 175.765 47.915 176.535 ;
        RECT 48.545 175.810 48.835 176.535 ;
        RECT 49.005 175.765 50.675 176.535 ;
        RECT 50.845 176.035 51.105 176.365 ;
        RECT 51.275 176.175 51.605 176.535 ;
        RECT 51.860 176.155 53.160 176.365 ;
        RECT 50.845 176.025 51.075 176.035 ;
        RECT 43.475 175.625 43.725 175.715 ;
        RECT 42.025 175.295 42.255 175.625 ;
        RECT 42.985 175.295 43.725 175.625 ;
        RECT 43.895 175.295 44.230 175.545 ;
        RECT 42.085 175.125 42.255 175.295 ;
        RECT 41.645 174.155 41.915 175.125 ;
        RECT 42.085 174.955 43.330 175.125 ;
        RECT 42.125 173.985 42.405 174.785 ;
        RECT 42.910 174.705 43.330 174.955 ;
        RECT 43.555 174.735 43.725 175.295 ;
        RECT 44.405 175.245 46.055 175.765 ;
        RECT 42.585 174.205 43.780 174.535 ;
        RECT 43.975 173.985 44.230 175.125 ;
        RECT 46.225 175.075 47.915 175.595 ;
        RECT 49.005 175.245 49.755 175.765 ;
        RECT 44.405 173.985 47.915 175.075 ;
        RECT 48.545 173.985 48.835 175.150 ;
        RECT 49.925 175.075 50.675 175.595 ;
        RECT 49.005 173.985 50.675 175.075 ;
        RECT 50.845 174.835 51.015 176.025 ;
        RECT 51.860 176.005 52.030 176.155 ;
        RECT 51.275 175.880 52.030 176.005 ;
        RECT 51.185 175.835 52.030 175.880 ;
        RECT 51.185 175.715 51.455 175.835 ;
        RECT 51.185 175.140 51.355 175.715 ;
        RECT 51.585 175.275 51.995 175.580 ;
        RECT 52.285 175.545 52.495 175.945 ;
        RECT 52.165 175.335 52.495 175.545 ;
        RECT 52.740 175.545 52.960 175.945 ;
        RECT 53.435 175.770 53.890 176.535 ;
        RECT 54.070 175.770 54.525 176.535 ;
        RECT 54.800 176.155 56.100 176.365 ;
        RECT 56.355 176.175 56.685 176.535 ;
        RECT 55.930 176.005 56.100 176.155 ;
        RECT 56.855 176.035 57.115 176.365 ;
        RECT 55.000 175.545 55.220 175.945 ;
        RECT 52.740 175.335 53.215 175.545 ;
        RECT 53.405 175.345 53.895 175.545 ;
        RECT 54.065 175.345 54.555 175.545 ;
        RECT 54.745 175.335 55.220 175.545 ;
        RECT 55.465 175.545 55.675 175.945 ;
        RECT 55.930 175.880 56.685 176.005 ;
        RECT 55.930 175.835 56.775 175.880 ;
        RECT 56.505 175.715 56.775 175.835 ;
        RECT 55.465 175.335 55.795 175.545 ;
        RECT 55.965 175.275 56.375 175.580 ;
        RECT 51.185 175.105 51.385 175.140 ;
        RECT 52.715 175.105 53.890 175.165 ;
        RECT 51.185 174.995 53.890 175.105 ;
        RECT 51.245 174.935 53.045 174.995 ;
        RECT 52.715 174.905 53.045 174.935 ;
        RECT 50.845 174.155 51.105 174.835 ;
        RECT 51.275 173.985 51.525 174.765 ;
        RECT 51.775 174.735 52.610 174.745 ;
        RECT 53.200 174.735 53.385 174.825 ;
        RECT 51.775 174.535 53.385 174.735 ;
        RECT 51.775 174.155 52.025 174.535 ;
        RECT 53.155 174.495 53.385 174.535 ;
        RECT 53.635 174.375 53.890 174.995 ;
        RECT 52.195 173.985 52.550 174.365 ;
        RECT 53.555 174.155 53.890 174.375 ;
        RECT 54.070 175.105 55.245 175.165 ;
        RECT 56.605 175.140 56.775 175.715 ;
        RECT 56.575 175.105 56.775 175.140 ;
        RECT 54.070 174.995 56.775 175.105 ;
        RECT 54.070 174.375 54.325 174.995 ;
        RECT 54.915 174.935 56.715 174.995 ;
        RECT 54.915 174.905 55.245 174.935 ;
        RECT 56.945 174.835 57.115 176.035 ;
        RECT 57.375 175.985 57.545 176.275 ;
        RECT 57.715 176.155 58.045 176.535 ;
        RECT 57.375 175.815 58.040 175.985 ;
        RECT 57.290 174.995 57.640 175.645 ;
        RECT 54.575 174.735 54.760 174.825 ;
        RECT 55.350 174.735 56.185 174.745 ;
        RECT 54.575 174.535 56.185 174.735 ;
        RECT 54.575 174.495 54.805 174.535 ;
        RECT 54.070 174.155 54.405 174.375 ;
        RECT 55.410 173.985 55.765 174.365 ;
        RECT 55.935 174.155 56.185 174.535 ;
        RECT 56.435 173.985 56.685 174.765 ;
        RECT 56.855 174.155 57.115 174.835 ;
        RECT 57.810 174.825 58.040 175.815 ;
        RECT 57.375 174.655 58.040 174.825 ;
        RECT 57.375 174.155 57.545 174.655 ;
        RECT 57.715 173.985 58.045 174.485 ;
        RECT 58.215 174.155 58.400 176.275 ;
        RECT 58.655 176.075 58.905 176.535 ;
        RECT 59.075 176.085 59.410 176.255 ;
        RECT 59.605 176.085 60.280 176.255 ;
        RECT 59.075 175.945 59.245 176.085 ;
        RECT 58.570 174.955 58.850 175.905 ;
        RECT 59.020 175.815 59.245 175.945 ;
        RECT 59.020 174.710 59.190 175.815 ;
        RECT 59.415 175.665 59.940 175.885 ;
        RECT 59.360 174.900 59.600 175.495 ;
        RECT 59.770 174.965 59.940 175.665 ;
        RECT 60.110 175.305 60.280 176.085 ;
        RECT 60.600 176.035 60.970 176.535 ;
        RECT 61.150 176.085 61.555 176.255 ;
        RECT 61.725 176.085 62.510 176.255 ;
        RECT 61.150 175.855 61.320 176.085 ;
        RECT 60.490 175.555 61.320 175.855 ;
        RECT 61.705 175.585 62.170 175.915 ;
        RECT 60.490 175.525 60.690 175.555 ;
        RECT 60.810 175.305 60.980 175.375 ;
        RECT 60.110 175.135 60.980 175.305 ;
        RECT 60.470 175.045 60.980 175.135 ;
        RECT 59.020 174.580 59.325 174.710 ;
        RECT 59.770 174.600 60.300 174.965 ;
        RECT 58.640 173.985 58.905 174.445 ;
        RECT 59.075 174.155 59.325 174.580 ;
        RECT 60.470 174.430 60.640 175.045 ;
        RECT 59.535 174.260 60.640 174.430 ;
        RECT 60.810 173.985 60.980 174.785 ;
        RECT 61.150 174.485 61.320 175.555 ;
        RECT 61.490 174.655 61.680 175.375 ;
        RECT 61.850 174.625 62.170 175.585 ;
        RECT 62.340 175.625 62.510 176.085 ;
        RECT 62.785 176.005 62.995 176.535 ;
        RECT 63.255 175.795 63.585 176.320 ;
        RECT 63.755 175.925 63.925 176.535 ;
        RECT 64.095 175.880 64.425 176.315 ;
        RECT 64.095 175.795 64.475 175.880 ;
        RECT 63.385 175.625 63.585 175.795 ;
        RECT 64.250 175.755 64.475 175.795 ;
        RECT 62.340 175.295 63.215 175.625 ;
        RECT 63.385 175.295 64.135 175.625 ;
        RECT 61.150 174.155 61.400 174.485 ;
        RECT 62.340 174.455 62.510 175.295 ;
        RECT 63.385 175.090 63.575 175.295 ;
        RECT 64.305 175.175 64.475 175.755 ;
        RECT 64.645 175.765 66.315 176.535 ;
        RECT 64.645 175.245 65.395 175.765 ;
        RECT 64.260 175.125 64.475 175.175 ;
        RECT 62.680 174.715 63.575 175.090 ;
        RECT 64.085 175.045 64.475 175.125 ;
        RECT 65.565 175.075 66.315 175.595 ;
        RECT 61.625 174.285 62.510 174.455 ;
        RECT 62.690 173.985 63.005 174.485 ;
        RECT 63.235 174.155 63.575 174.715 ;
        RECT 63.745 173.985 63.915 174.995 ;
        RECT 64.085 174.200 64.415 175.045 ;
        RECT 64.645 173.985 66.315 175.075 ;
        RECT 66.495 174.165 66.755 176.355 ;
        RECT 67.015 176.165 67.685 176.535 ;
        RECT 67.865 175.985 68.175 176.355 ;
        RECT 66.945 175.785 68.175 175.985 ;
        RECT 66.945 175.115 67.235 175.785 ;
        RECT 68.355 175.605 68.585 176.245 ;
        RECT 68.765 175.805 69.055 176.535 ;
        RECT 69.245 175.785 70.455 176.535 ;
        RECT 70.625 175.885 70.885 176.365 ;
        RECT 71.055 175.995 71.305 176.535 ;
        RECT 67.415 175.295 67.880 175.605 ;
        RECT 68.060 175.295 68.585 175.605 ;
        RECT 68.765 175.295 69.065 175.625 ;
        RECT 69.245 175.245 69.765 175.785 ;
        RECT 66.945 174.895 67.715 175.115 ;
        RECT 66.925 173.985 67.265 174.715 ;
        RECT 67.445 174.165 67.715 174.895 ;
        RECT 67.895 174.875 69.055 175.115 ;
        RECT 69.935 175.075 70.455 175.615 ;
        RECT 67.895 174.165 68.125 174.875 ;
        RECT 68.295 173.985 68.625 174.695 ;
        RECT 68.795 174.165 69.055 174.875 ;
        RECT 69.245 173.985 70.455 175.075 ;
        RECT 70.625 174.855 70.795 175.885 ;
        RECT 71.475 175.830 71.695 176.315 ;
        RECT 70.965 175.235 71.195 175.630 ;
        RECT 71.365 175.405 71.695 175.830 ;
        RECT 71.865 176.155 72.755 176.325 ;
        RECT 71.865 175.430 72.035 176.155 ;
        RECT 72.205 175.600 72.755 175.985 ;
        RECT 72.925 175.785 74.135 176.535 ;
        RECT 74.305 175.810 74.595 176.535 ;
        RECT 74.765 175.795 75.150 176.365 ;
        RECT 75.320 176.075 75.645 176.535 ;
        RECT 76.165 175.905 76.445 176.365 ;
        RECT 71.865 175.360 72.755 175.430 ;
        RECT 71.860 175.335 72.755 175.360 ;
        RECT 71.850 175.320 72.755 175.335 ;
        RECT 71.845 175.305 72.755 175.320 ;
        RECT 71.835 175.300 72.755 175.305 ;
        RECT 71.830 175.290 72.755 175.300 ;
        RECT 71.825 175.280 72.755 175.290 ;
        RECT 71.815 175.275 72.755 175.280 ;
        RECT 71.805 175.265 72.755 175.275 ;
        RECT 71.795 175.260 72.755 175.265 ;
        RECT 71.795 175.255 72.130 175.260 ;
        RECT 71.780 175.250 72.130 175.255 ;
        RECT 71.765 175.240 72.130 175.250 ;
        RECT 71.740 175.235 72.130 175.240 ;
        RECT 70.965 175.230 72.130 175.235 ;
        RECT 70.965 175.195 72.100 175.230 ;
        RECT 70.965 175.170 72.065 175.195 ;
        RECT 70.965 175.140 72.035 175.170 ;
        RECT 70.965 175.110 72.015 175.140 ;
        RECT 70.965 175.080 71.995 175.110 ;
        RECT 70.965 175.070 71.925 175.080 ;
        RECT 70.965 175.060 71.900 175.070 ;
        RECT 70.965 175.045 71.880 175.060 ;
        RECT 70.965 175.030 71.860 175.045 ;
        RECT 71.070 175.020 71.855 175.030 ;
        RECT 71.070 174.985 71.840 175.020 ;
        RECT 70.625 174.155 70.900 174.855 ;
        RECT 71.070 174.735 71.825 174.985 ;
        RECT 71.995 174.665 72.325 174.910 ;
        RECT 72.495 174.810 72.755 175.260 ;
        RECT 72.925 175.245 73.445 175.785 ;
        RECT 73.615 175.075 74.135 175.615 ;
        RECT 72.140 174.640 72.325 174.665 ;
        RECT 72.140 174.540 72.755 174.640 ;
        RECT 71.070 173.985 71.325 174.530 ;
        RECT 71.495 174.155 71.975 174.495 ;
        RECT 72.150 173.985 72.755 174.540 ;
        RECT 72.925 173.985 74.135 175.075 ;
        RECT 74.305 173.985 74.595 175.150 ;
        RECT 74.765 175.125 75.045 175.795 ;
        RECT 75.320 175.735 76.445 175.905 ;
        RECT 75.320 175.625 75.770 175.735 ;
        RECT 75.215 175.295 75.770 175.625 ;
        RECT 76.635 175.565 77.035 176.365 ;
        RECT 77.435 176.075 77.705 176.535 ;
        RECT 77.875 175.905 78.160 176.365 ;
        RECT 78.450 176.135 78.785 176.535 ;
        RECT 78.955 175.965 79.160 176.365 ;
        RECT 79.370 176.055 79.645 176.535 ;
        RECT 79.855 176.035 80.115 176.365 ;
        RECT 74.765 174.155 75.150 175.125 ;
        RECT 75.320 174.835 75.770 175.295 ;
        RECT 75.940 175.005 77.035 175.565 ;
        RECT 75.320 174.615 76.445 174.835 ;
        RECT 75.320 173.985 75.645 174.445 ;
        RECT 76.165 174.155 76.445 174.615 ;
        RECT 76.635 174.155 77.035 175.005 ;
        RECT 77.205 175.735 78.160 175.905 ;
        RECT 78.475 175.795 79.160 175.965 ;
        RECT 77.205 174.835 77.415 175.735 ;
        RECT 77.585 175.005 78.275 175.565 ;
        RECT 77.205 174.615 78.160 174.835 ;
        RECT 77.435 173.985 77.705 174.445 ;
        RECT 77.875 174.155 78.160 174.615 ;
        RECT 78.475 174.765 78.815 175.795 ;
        RECT 78.985 175.125 79.235 175.625 ;
        RECT 79.415 175.295 79.775 175.875 ;
        RECT 79.945 175.125 80.115 176.035 ;
        RECT 80.285 175.765 82.875 176.535 ;
        RECT 80.285 175.245 81.495 175.765 ;
        RECT 78.985 174.955 80.115 175.125 ;
        RECT 81.665 175.075 82.875 175.595 ;
        RECT 78.475 174.590 79.140 174.765 ;
        RECT 78.450 173.985 78.785 174.410 ;
        RECT 78.955 174.185 79.140 174.590 ;
        RECT 79.345 173.985 79.675 174.765 ;
        RECT 79.845 174.185 80.115 174.955 ;
        RECT 80.285 173.985 82.875 175.075 ;
        RECT 83.055 174.165 83.315 176.355 ;
        RECT 83.575 176.165 84.245 176.535 ;
        RECT 84.425 175.985 84.735 176.355 ;
        RECT 83.505 175.785 84.735 175.985 ;
        RECT 83.505 175.115 83.795 175.785 ;
        RECT 84.915 175.605 85.145 176.245 ;
        RECT 85.325 175.805 85.615 176.535 ;
        RECT 85.805 175.765 89.315 176.535 ;
        RECT 89.485 175.785 90.695 176.535 ;
        RECT 90.955 175.985 91.125 176.275 ;
        RECT 91.295 176.155 91.625 176.535 ;
        RECT 90.955 175.815 91.620 175.985 ;
        RECT 83.975 175.295 84.440 175.605 ;
        RECT 84.620 175.295 85.145 175.605 ;
        RECT 85.325 175.295 85.625 175.625 ;
        RECT 85.805 175.245 87.455 175.765 ;
        RECT 83.505 174.895 84.275 175.115 ;
        RECT 83.485 173.985 83.825 174.715 ;
        RECT 84.005 174.165 84.275 174.895 ;
        RECT 84.455 174.875 85.615 175.115 ;
        RECT 87.625 175.075 89.315 175.595 ;
        RECT 89.485 175.245 90.005 175.785 ;
        RECT 90.175 175.075 90.695 175.615 ;
        RECT 84.455 174.165 84.685 174.875 ;
        RECT 84.855 173.985 85.185 174.695 ;
        RECT 85.355 174.165 85.615 174.875 ;
        RECT 85.805 173.985 89.315 175.075 ;
        RECT 89.485 173.985 90.695 175.075 ;
        RECT 90.870 174.995 91.220 175.645 ;
        RECT 91.390 174.825 91.620 175.815 ;
        RECT 90.955 174.655 91.620 174.825 ;
        RECT 90.955 174.155 91.125 174.655 ;
        RECT 91.295 173.985 91.625 174.485 ;
        RECT 91.795 174.155 91.980 176.275 ;
        RECT 92.235 176.075 92.485 176.535 ;
        RECT 92.655 176.085 92.990 176.255 ;
        RECT 93.185 176.085 93.860 176.255 ;
        RECT 92.655 175.945 92.825 176.085 ;
        RECT 92.150 174.955 92.430 175.905 ;
        RECT 92.600 175.815 92.825 175.945 ;
        RECT 92.600 174.710 92.770 175.815 ;
        RECT 92.995 175.665 93.520 175.885 ;
        RECT 92.940 174.900 93.180 175.495 ;
        RECT 93.350 174.965 93.520 175.665 ;
        RECT 93.690 175.305 93.860 176.085 ;
        RECT 94.180 176.035 94.550 176.535 ;
        RECT 94.730 176.085 95.135 176.255 ;
        RECT 95.305 176.085 96.090 176.255 ;
        RECT 94.730 175.855 94.900 176.085 ;
        RECT 94.070 175.555 94.900 175.855 ;
        RECT 95.285 175.585 95.750 175.915 ;
        RECT 94.070 175.525 94.270 175.555 ;
        RECT 94.390 175.305 94.560 175.375 ;
        RECT 93.690 175.135 94.560 175.305 ;
        RECT 94.050 175.045 94.560 175.135 ;
        RECT 92.600 174.580 92.905 174.710 ;
        RECT 93.350 174.600 93.880 174.965 ;
        RECT 92.220 173.985 92.485 174.445 ;
        RECT 92.655 174.155 92.905 174.580 ;
        RECT 94.050 174.430 94.220 175.045 ;
        RECT 93.115 174.260 94.220 174.430 ;
        RECT 94.390 173.985 94.560 174.785 ;
        RECT 94.730 174.485 94.900 175.555 ;
        RECT 95.070 174.655 95.260 175.375 ;
        RECT 95.430 174.625 95.750 175.585 ;
        RECT 95.920 175.625 96.090 176.085 ;
        RECT 96.365 176.005 96.575 176.535 ;
        RECT 96.835 175.795 97.165 176.320 ;
        RECT 97.335 175.925 97.505 176.535 ;
        RECT 97.675 175.880 98.005 176.315 ;
        RECT 97.675 175.795 98.055 175.880 ;
        RECT 96.965 175.625 97.165 175.795 ;
        RECT 97.830 175.755 98.055 175.795 ;
        RECT 95.920 175.295 96.795 175.625 ;
        RECT 96.965 175.295 97.715 175.625 ;
        RECT 94.730 174.155 94.980 174.485 ;
        RECT 95.920 174.455 96.090 175.295 ;
        RECT 96.965 175.090 97.155 175.295 ;
        RECT 97.885 175.175 98.055 175.755 ;
        RECT 98.225 175.765 99.895 176.535 ;
        RECT 100.065 175.810 100.355 176.535 ;
        RECT 100.530 175.795 100.785 176.365 ;
        RECT 100.955 176.135 101.285 176.535 ;
        RECT 101.710 176.000 102.240 176.365 ;
        RECT 101.710 175.965 101.885 176.000 ;
        RECT 100.955 175.795 101.885 175.965 ;
        RECT 98.225 175.245 98.975 175.765 ;
        RECT 97.840 175.125 98.055 175.175 ;
        RECT 96.260 174.715 97.155 175.090 ;
        RECT 97.665 175.045 98.055 175.125 ;
        RECT 99.145 175.075 99.895 175.595 ;
        RECT 95.205 174.285 96.090 174.455 ;
        RECT 96.270 173.985 96.585 174.485 ;
        RECT 96.815 174.155 97.155 174.715 ;
        RECT 97.325 173.985 97.495 174.995 ;
        RECT 97.665 174.200 97.995 175.045 ;
        RECT 98.225 173.985 99.895 175.075 ;
        RECT 100.065 173.985 100.355 175.150 ;
        RECT 100.530 175.125 100.700 175.795 ;
        RECT 100.955 175.625 101.125 175.795 ;
        RECT 100.870 175.295 101.125 175.625 ;
        RECT 101.350 175.295 101.545 175.625 ;
        RECT 100.530 174.155 100.865 175.125 ;
        RECT 101.035 173.985 101.205 175.125 ;
        RECT 101.375 174.325 101.545 175.295 ;
        RECT 101.715 174.665 101.885 175.795 ;
        RECT 102.055 175.005 102.225 175.805 ;
        RECT 102.430 175.515 102.705 176.365 ;
        RECT 102.425 175.345 102.705 175.515 ;
        RECT 102.430 175.205 102.705 175.345 ;
        RECT 102.875 175.005 103.065 176.365 ;
        RECT 103.245 176.000 103.755 176.535 ;
        RECT 103.975 175.725 104.220 176.330 ;
        RECT 104.665 175.765 107.255 176.535 ;
        RECT 107.885 176.075 108.445 176.365 ;
        RECT 108.615 176.075 108.865 176.535 ;
        RECT 103.265 175.555 104.495 175.725 ;
        RECT 102.055 174.835 103.065 175.005 ;
        RECT 103.235 174.990 103.985 175.180 ;
        RECT 101.715 174.495 102.840 174.665 ;
        RECT 103.235 174.325 103.405 174.990 ;
        RECT 104.155 174.745 104.495 175.555 ;
        RECT 104.665 175.245 105.875 175.765 ;
        RECT 106.045 175.075 107.255 175.595 ;
        RECT 101.375 174.155 103.405 174.325 ;
        RECT 103.575 173.985 103.745 174.745 ;
        RECT 103.980 174.335 104.495 174.745 ;
        RECT 104.665 173.985 107.255 175.075 ;
        RECT 107.885 174.705 108.135 176.075 ;
        RECT 109.485 175.905 109.815 176.265 ;
        RECT 108.425 175.715 109.815 175.905 ;
        RECT 110.185 175.765 113.695 176.535 ;
        RECT 114.325 176.075 114.885 176.365 ;
        RECT 115.055 176.075 115.305 176.535 ;
        RECT 108.425 175.625 108.595 175.715 ;
        RECT 108.305 175.295 108.595 175.625 ;
        RECT 108.765 175.295 109.105 175.545 ;
        RECT 109.325 175.295 110.000 175.545 ;
        RECT 108.425 175.045 108.595 175.295 ;
        RECT 108.425 174.875 109.365 175.045 ;
        RECT 109.735 174.935 110.000 175.295 ;
        RECT 110.185 175.245 111.835 175.765 ;
        RECT 112.005 175.075 113.695 175.595 ;
        RECT 107.885 174.155 108.345 174.705 ;
        RECT 108.535 173.985 108.865 174.705 ;
        RECT 109.065 174.325 109.365 174.875 ;
        RECT 109.535 173.985 109.815 174.655 ;
        RECT 110.185 173.985 113.695 175.075 ;
        RECT 114.325 174.705 114.575 176.075 ;
        RECT 115.925 175.905 116.255 176.265 ;
        RECT 114.865 175.715 116.255 175.905 ;
        RECT 117.550 175.795 117.805 176.365 ;
        RECT 117.975 176.135 118.305 176.535 ;
        RECT 118.730 176.000 119.260 176.365 ;
        RECT 118.730 175.965 118.905 176.000 ;
        RECT 117.975 175.795 118.905 175.965 ;
        RECT 114.865 175.625 115.035 175.715 ;
        RECT 114.745 175.295 115.035 175.625 ;
        RECT 115.205 175.295 115.545 175.545 ;
        RECT 115.765 175.295 116.440 175.545 ;
        RECT 114.865 175.045 115.035 175.295 ;
        RECT 114.865 174.875 115.805 175.045 ;
        RECT 116.175 174.935 116.440 175.295 ;
        RECT 117.550 175.125 117.720 175.795 ;
        RECT 117.975 175.625 118.145 175.795 ;
        RECT 117.890 175.295 118.145 175.625 ;
        RECT 118.370 175.295 118.565 175.625 ;
        RECT 114.325 174.155 114.785 174.705 ;
        RECT 114.975 173.985 115.305 174.705 ;
        RECT 115.505 174.325 115.805 174.875 ;
        RECT 115.975 173.985 116.255 174.655 ;
        RECT 117.550 174.155 117.885 175.125 ;
        RECT 118.055 173.985 118.225 175.125 ;
        RECT 118.395 174.325 118.565 175.295 ;
        RECT 118.735 174.665 118.905 175.795 ;
        RECT 119.075 175.005 119.245 175.805 ;
        RECT 119.450 175.515 119.725 176.365 ;
        RECT 119.445 175.345 119.725 175.515 ;
        RECT 119.450 175.205 119.725 175.345 ;
        RECT 119.895 175.005 120.085 176.365 ;
        RECT 120.265 176.000 120.775 176.535 ;
        RECT 120.995 175.725 121.240 176.330 ;
        RECT 121.685 176.075 122.245 176.365 ;
        RECT 122.415 176.075 122.665 176.535 ;
        RECT 120.285 175.555 121.515 175.725 ;
        RECT 119.075 174.835 120.085 175.005 ;
        RECT 120.255 174.990 121.005 175.180 ;
        RECT 118.735 174.495 119.860 174.665 ;
        RECT 120.255 174.325 120.425 174.990 ;
        RECT 121.175 174.745 121.515 175.555 ;
        RECT 118.395 174.155 120.425 174.325 ;
        RECT 120.595 173.985 120.765 174.745 ;
        RECT 121.000 174.335 121.515 174.745 ;
        RECT 121.685 174.705 121.935 176.075 ;
        RECT 123.285 175.905 123.615 176.265 ;
        RECT 122.225 175.715 123.615 175.905 ;
        RECT 123.985 175.765 125.655 176.535 ;
        RECT 125.825 175.810 126.115 176.535 ;
        RECT 126.905 175.975 127.235 176.365 ;
        RECT 127.405 176.145 128.590 176.315 ;
        RECT 128.850 176.065 129.020 176.535 ;
        RECT 126.905 175.795 127.415 175.975 ;
        RECT 122.225 175.625 122.395 175.715 ;
        RECT 122.105 175.295 122.395 175.625 ;
        RECT 122.565 175.295 122.905 175.545 ;
        RECT 123.125 175.295 123.800 175.545 ;
        RECT 122.225 175.045 122.395 175.295 ;
        RECT 122.225 174.875 123.165 175.045 ;
        RECT 123.535 174.935 123.800 175.295 ;
        RECT 123.985 175.245 124.735 175.765 ;
        RECT 124.905 175.075 125.655 175.595 ;
        RECT 126.745 175.335 127.075 175.625 ;
        RECT 127.245 175.165 127.415 175.795 ;
        RECT 127.820 175.885 128.205 175.975 ;
        RECT 129.190 175.885 129.520 176.350 ;
        RECT 127.820 175.715 129.520 175.885 ;
        RECT 129.690 175.715 129.860 176.535 ;
        RECT 130.030 175.715 130.715 176.355 ;
        RECT 127.585 175.335 127.915 175.545 ;
        RECT 128.095 175.295 128.475 175.545 ;
        RECT 121.685 174.155 122.145 174.705 ;
        RECT 122.335 173.985 122.665 174.705 ;
        RECT 122.865 174.325 123.165 174.875 ;
        RECT 123.335 173.985 123.615 174.655 ;
        RECT 123.985 173.985 125.655 175.075 ;
        RECT 125.825 173.985 126.115 175.150 ;
        RECT 126.900 174.995 127.985 175.165 ;
        RECT 126.900 174.155 127.200 174.995 ;
        RECT 127.395 173.985 127.645 174.825 ;
        RECT 127.815 174.745 127.985 174.995 ;
        RECT 128.155 174.915 128.475 175.295 ;
        RECT 128.665 175.335 129.150 175.545 ;
        RECT 129.340 175.335 129.790 175.545 ;
        RECT 129.960 175.335 130.295 175.545 ;
        RECT 128.665 175.175 129.040 175.335 ;
        RECT 128.645 175.005 129.040 175.175 ;
        RECT 129.960 175.165 130.130 175.335 ;
        RECT 128.665 174.915 129.040 175.005 ;
        RECT 129.210 174.995 130.130 175.165 ;
        RECT 129.210 174.745 129.380 174.995 ;
        RECT 127.815 174.575 129.380 174.745 ;
        RECT 128.235 174.155 129.040 174.575 ;
        RECT 129.550 173.985 129.880 174.825 ;
        RECT 130.465 174.745 130.715 175.715 ;
        RECT 130.885 175.765 132.555 176.535 ;
        RECT 133.185 175.795 133.570 176.365 ;
        RECT 133.740 176.075 134.065 176.535 ;
        RECT 134.585 175.905 134.865 176.365 ;
        RECT 130.885 175.245 131.635 175.765 ;
        RECT 131.805 175.075 132.555 175.595 ;
        RECT 130.050 174.155 130.715 174.745 ;
        RECT 130.885 173.985 132.555 175.075 ;
        RECT 133.185 175.125 133.465 175.795 ;
        RECT 133.740 175.735 134.865 175.905 ;
        RECT 133.740 175.625 134.190 175.735 ;
        RECT 133.635 175.295 134.190 175.625 ;
        RECT 135.055 175.565 135.455 176.365 ;
        RECT 135.855 176.075 136.125 176.535 ;
        RECT 136.295 175.905 136.580 176.365 ;
        RECT 136.890 176.145 137.220 176.535 ;
        RECT 137.390 175.975 137.615 176.355 ;
        RECT 133.185 174.155 133.570 175.125 ;
        RECT 133.740 174.835 134.190 175.295 ;
        RECT 134.360 175.005 135.455 175.565 ;
        RECT 133.740 174.615 134.865 174.835 ;
        RECT 133.740 173.985 134.065 174.445 ;
        RECT 134.585 174.155 134.865 174.615 ;
        RECT 135.055 174.155 135.455 175.005 ;
        RECT 135.625 175.735 136.580 175.905 ;
        RECT 135.625 174.835 135.835 175.735 ;
        RECT 136.005 175.005 136.695 175.565 ;
        RECT 136.875 175.295 137.115 175.945 ;
        RECT 137.285 175.795 137.615 175.975 ;
        RECT 137.285 175.125 137.460 175.795 ;
        RECT 137.815 175.625 138.045 176.245 ;
        RECT 138.225 175.805 138.525 176.535 ;
        RECT 138.820 175.905 139.105 176.365 ;
        RECT 139.275 176.075 139.545 176.535 ;
        RECT 138.820 175.735 139.775 175.905 ;
        RECT 137.630 175.295 138.045 175.625 ;
        RECT 138.225 175.295 138.520 175.625 ;
        RECT 136.875 174.935 137.460 175.125 ;
        RECT 135.625 174.615 136.580 174.835 ;
        RECT 135.855 173.985 136.125 174.445 ;
        RECT 136.295 174.155 136.580 174.615 ;
        RECT 136.875 174.165 137.150 174.935 ;
        RECT 137.630 174.765 138.525 175.095 ;
        RECT 138.705 175.005 139.395 175.565 ;
        RECT 139.565 174.835 139.775 175.735 ;
        RECT 137.320 174.595 138.525 174.765 ;
        RECT 137.320 174.165 137.650 174.595 ;
        RECT 137.820 173.985 138.015 174.425 ;
        RECT 138.195 174.165 138.525 174.595 ;
        RECT 138.820 174.615 139.775 174.835 ;
        RECT 139.945 175.565 140.345 176.365 ;
        RECT 140.535 175.905 140.815 176.365 ;
        RECT 141.335 176.075 141.660 176.535 ;
        RECT 140.535 175.735 141.660 175.905 ;
        RECT 141.830 175.795 142.215 176.365 ;
        RECT 141.210 175.625 141.660 175.735 ;
        RECT 139.945 175.005 141.040 175.565 ;
        RECT 141.210 175.295 141.765 175.625 ;
        RECT 138.820 174.155 139.105 174.615 ;
        RECT 139.275 173.985 139.545 174.445 ;
        RECT 139.945 174.155 140.345 175.005 ;
        RECT 141.210 174.835 141.660 175.295 ;
        RECT 141.935 175.125 142.215 175.795 ;
        RECT 140.535 174.615 141.660 174.835 ;
        RECT 140.535 174.155 140.815 174.615 ;
        RECT 141.335 173.985 141.660 174.445 ;
        RECT 141.830 174.155 142.215 175.125 ;
        RECT 142.420 175.795 143.035 176.365 ;
        RECT 143.205 176.025 143.420 176.535 ;
        RECT 143.650 176.025 143.930 176.355 ;
        RECT 144.110 176.025 144.350 176.535 ;
        RECT 145.770 176.025 146.010 176.535 ;
        RECT 146.190 176.025 146.470 176.355 ;
        RECT 146.700 176.025 146.915 176.535 ;
        RECT 142.420 174.775 142.735 175.795 ;
        RECT 142.905 175.125 143.075 175.625 ;
        RECT 143.325 175.295 143.590 175.855 ;
        RECT 143.760 175.125 143.930 176.025 ;
        RECT 144.100 175.295 144.455 175.855 ;
        RECT 145.665 175.295 146.020 175.855 ;
        RECT 146.190 175.125 146.360 176.025 ;
        RECT 146.530 175.295 146.795 175.855 ;
        RECT 147.085 175.795 147.700 176.365 ;
        RECT 147.905 176.155 148.795 176.325 ;
        RECT 147.045 175.125 147.215 175.625 ;
        RECT 142.905 174.955 144.330 175.125 ;
        RECT 142.420 174.155 142.955 174.775 ;
        RECT 143.125 173.985 143.455 174.785 ;
        RECT 143.940 174.780 144.330 174.955 ;
        RECT 145.790 174.955 147.215 175.125 ;
        RECT 145.790 174.780 146.180 174.955 ;
        RECT 146.665 173.985 146.995 174.785 ;
        RECT 147.385 174.775 147.700 175.795 ;
        RECT 147.905 175.600 148.455 175.985 ;
        RECT 148.625 175.430 148.795 176.155 ;
        RECT 147.905 175.360 148.795 175.430 ;
        RECT 148.965 175.830 149.185 176.315 ;
        RECT 149.355 175.995 149.605 176.535 ;
        RECT 149.775 175.885 150.035 176.365 ;
        RECT 148.965 175.405 149.295 175.830 ;
        RECT 147.905 175.335 148.800 175.360 ;
        RECT 147.905 175.320 148.810 175.335 ;
        RECT 147.905 175.305 148.815 175.320 ;
        RECT 147.905 175.300 148.825 175.305 ;
        RECT 147.905 175.290 148.830 175.300 ;
        RECT 147.905 175.280 148.835 175.290 ;
        RECT 147.905 175.275 148.845 175.280 ;
        RECT 147.905 175.265 148.855 175.275 ;
        RECT 147.905 175.260 148.865 175.265 ;
        RECT 147.905 174.810 148.165 175.260 ;
        RECT 148.530 175.255 148.865 175.260 ;
        RECT 148.530 175.250 148.880 175.255 ;
        RECT 148.530 175.240 148.895 175.250 ;
        RECT 148.530 175.235 148.920 175.240 ;
        RECT 149.465 175.235 149.695 175.630 ;
        RECT 148.530 175.230 149.695 175.235 ;
        RECT 148.560 175.195 149.695 175.230 ;
        RECT 148.595 175.170 149.695 175.195 ;
        RECT 148.625 175.140 149.695 175.170 ;
        RECT 148.645 175.110 149.695 175.140 ;
        RECT 148.665 175.080 149.695 175.110 ;
        RECT 148.735 175.070 149.695 175.080 ;
        RECT 148.760 175.060 149.695 175.070 ;
        RECT 148.780 175.045 149.695 175.060 ;
        RECT 148.800 175.030 149.695 175.045 ;
        RECT 148.805 175.020 149.590 175.030 ;
        RECT 148.820 174.985 149.590 175.020 ;
        RECT 147.165 174.155 147.700 174.775 ;
        RECT 148.335 174.665 148.665 174.910 ;
        RECT 148.835 174.735 149.590 174.985 ;
        RECT 149.865 174.855 150.035 175.885 ;
        RECT 148.335 174.640 148.520 174.665 ;
        RECT 147.905 174.540 148.520 174.640 ;
        RECT 147.905 173.985 148.510 174.540 ;
        RECT 148.685 174.155 149.165 174.495 ;
        RECT 149.335 173.985 149.590 174.530 ;
        RECT 149.760 174.155 150.035 174.855 ;
        RECT 150.205 175.860 150.465 176.365 ;
        RECT 150.645 176.155 150.975 176.535 ;
        RECT 151.155 175.985 151.325 176.365 ;
        RECT 150.205 175.060 150.375 175.860 ;
        RECT 150.660 175.815 151.325 175.985 ;
        RECT 150.660 175.560 150.830 175.815 ;
        RECT 151.585 175.810 151.875 176.535 ;
        RECT 152.045 175.785 153.255 176.535 ;
        RECT 150.545 175.230 150.830 175.560 ;
        RECT 151.065 175.265 151.395 175.635 ;
        RECT 152.045 175.245 152.565 175.785 ;
        RECT 153.485 175.715 153.695 176.535 ;
        RECT 153.865 175.735 154.195 176.365 ;
        RECT 150.660 175.085 150.830 175.230 ;
        RECT 150.205 174.155 150.475 175.060 ;
        RECT 150.660 174.915 151.325 175.085 ;
        RECT 150.645 173.985 150.975 174.745 ;
        RECT 151.155 174.155 151.325 174.915 ;
        RECT 151.585 173.985 151.875 175.150 ;
        RECT 152.735 175.075 153.255 175.615 ;
        RECT 153.865 175.135 154.115 175.735 ;
        RECT 154.365 175.715 154.595 176.535 ;
        RECT 155.725 175.785 156.935 176.535 ;
        RECT 154.285 175.295 154.615 175.545 ;
        RECT 152.045 173.985 153.255 175.075 ;
        RECT 153.485 173.985 153.695 175.125 ;
        RECT 153.865 174.155 154.195 175.135 ;
        RECT 154.365 173.985 154.595 175.125 ;
        RECT 155.725 175.075 156.245 175.615 ;
        RECT 156.415 175.245 156.935 175.785 ;
        RECT 155.725 173.985 156.935 175.075 ;
        RECT 22.700 173.815 157.020 173.985 ;
        RECT 22.785 172.725 23.995 173.815 ;
        RECT 22.785 172.015 23.305 172.555 ;
        RECT 23.475 172.185 23.995 172.725 ;
        RECT 24.255 172.885 24.425 173.645 ;
        RECT 24.605 173.055 24.935 173.815 ;
        RECT 24.255 172.715 24.920 172.885 ;
        RECT 25.105 172.740 25.375 173.645 ;
        RECT 24.750 172.570 24.920 172.715 ;
        RECT 24.185 172.165 24.515 172.535 ;
        RECT 24.750 172.240 25.035 172.570 ;
        RECT 22.785 171.265 23.995 172.015 ;
        RECT 24.750 171.985 24.920 172.240 ;
        RECT 24.255 171.815 24.920 171.985 ;
        RECT 25.205 171.940 25.375 172.740 ;
        RECT 25.545 172.675 25.825 173.815 ;
        RECT 25.995 172.665 26.325 173.645 ;
        RECT 26.495 172.675 26.755 173.815 ;
        RECT 26.925 172.945 27.200 173.645 ;
        RECT 27.410 173.270 27.625 173.815 ;
        RECT 27.795 173.305 28.270 173.645 ;
        RECT 28.440 173.310 29.055 173.815 ;
        RECT 28.440 173.135 28.635 173.310 ;
        RECT 25.555 172.235 25.890 172.505 ;
        RECT 26.060 172.065 26.230 172.665 ;
        RECT 26.400 172.255 26.735 172.505 ;
        RECT 24.255 171.435 24.425 171.815 ;
        RECT 24.605 171.265 24.935 171.645 ;
        RECT 25.115 171.435 25.375 171.940 ;
        RECT 25.545 171.265 25.855 172.065 ;
        RECT 26.060 171.435 26.755 172.065 ;
        RECT 26.925 171.915 27.095 172.945 ;
        RECT 27.370 172.775 28.085 173.070 ;
        RECT 28.305 172.945 28.635 173.135 ;
        RECT 28.805 172.775 29.055 173.140 ;
        RECT 27.265 172.605 29.055 172.775 ;
        RECT 27.265 172.175 27.495 172.605 ;
        RECT 26.925 171.435 27.185 171.915 ;
        RECT 27.665 171.905 28.075 172.425 ;
        RECT 27.355 171.265 27.685 171.725 ;
        RECT 27.875 171.485 28.075 171.905 ;
        RECT 28.245 171.750 28.500 172.605 ;
        RECT 29.295 172.425 29.465 173.645 ;
        RECT 29.715 173.305 29.975 173.815 ;
        RECT 30.605 173.260 31.210 173.815 ;
        RECT 31.385 173.305 31.865 173.645 ;
        RECT 32.035 173.270 32.290 173.815 ;
        RECT 30.605 173.160 31.220 173.260 ;
        RECT 31.035 173.135 31.220 173.160 ;
        RECT 28.670 172.175 29.465 172.425 ;
        RECT 29.635 172.255 29.975 173.135 ;
        RECT 30.605 172.540 30.865 172.990 ;
        RECT 31.035 172.890 31.365 173.135 ;
        RECT 31.535 172.815 32.290 173.065 ;
        RECT 32.460 172.945 32.735 173.645 ;
        RECT 31.520 172.780 32.290 172.815 ;
        RECT 31.505 172.770 32.290 172.780 ;
        RECT 31.500 172.755 32.395 172.770 ;
        RECT 31.480 172.740 32.395 172.755 ;
        RECT 31.460 172.730 32.395 172.740 ;
        RECT 31.435 172.720 32.395 172.730 ;
        RECT 31.365 172.690 32.395 172.720 ;
        RECT 31.345 172.660 32.395 172.690 ;
        RECT 31.325 172.630 32.395 172.660 ;
        RECT 31.295 172.605 32.395 172.630 ;
        RECT 31.260 172.570 32.395 172.605 ;
        RECT 31.230 172.565 32.395 172.570 ;
        RECT 31.230 172.560 31.620 172.565 ;
        RECT 31.230 172.550 31.595 172.560 ;
        RECT 31.230 172.545 31.580 172.550 ;
        RECT 31.230 172.540 31.565 172.545 ;
        RECT 30.605 172.535 31.565 172.540 ;
        RECT 30.605 172.525 31.555 172.535 ;
        RECT 30.605 172.520 31.545 172.525 ;
        RECT 30.605 172.510 31.535 172.520 ;
        RECT 30.605 172.500 31.530 172.510 ;
        RECT 30.605 172.495 31.525 172.500 ;
        RECT 30.605 172.480 31.515 172.495 ;
        RECT 30.605 172.465 31.510 172.480 ;
        RECT 30.605 172.440 31.500 172.465 ;
        RECT 30.605 172.370 31.495 172.440 ;
        RECT 29.215 172.085 29.465 172.175 ;
        RECT 28.245 171.485 29.035 171.750 ;
        RECT 29.215 171.665 29.545 172.085 ;
        RECT 29.715 171.265 29.975 172.085 ;
        RECT 30.605 171.815 31.155 172.200 ;
        RECT 31.325 171.645 31.495 172.370 ;
        RECT 30.605 171.475 31.495 171.645 ;
        RECT 31.665 171.970 31.995 172.395 ;
        RECT 32.165 172.170 32.395 172.565 ;
        RECT 31.665 171.485 31.885 171.970 ;
        RECT 32.565 171.915 32.735 172.945 ;
        RECT 32.055 171.265 32.305 171.805 ;
        RECT 32.475 171.435 32.735 171.915 ;
        RECT 32.905 172.945 33.180 173.645 ;
        RECT 33.350 173.270 33.605 173.815 ;
        RECT 33.775 173.305 34.255 173.645 ;
        RECT 34.430 173.260 35.035 173.815 ;
        RECT 34.420 173.160 35.035 173.260 ;
        RECT 34.420 173.135 34.605 173.160 ;
        RECT 32.905 171.915 33.075 172.945 ;
        RECT 33.350 172.815 34.105 173.065 ;
        RECT 34.275 172.890 34.605 173.135 ;
        RECT 33.350 172.780 34.120 172.815 ;
        RECT 33.350 172.770 34.135 172.780 ;
        RECT 33.245 172.755 34.140 172.770 ;
        RECT 33.245 172.740 34.160 172.755 ;
        RECT 33.245 172.730 34.180 172.740 ;
        RECT 33.245 172.720 34.205 172.730 ;
        RECT 33.245 172.690 34.275 172.720 ;
        RECT 33.245 172.660 34.295 172.690 ;
        RECT 33.245 172.630 34.315 172.660 ;
        RECT 33.245 172.605 34.345 172.630 ;
        RECT 33.245 172.570 34.380 172.605 ;
        RECT 33.245 172.565 34.410 172.570 ;
        RECT 33.245 172.170 33.475 172.565 ;
        RECT 34.020 172.560 34.410 172.565 ;
        RECT 34.045 172.550 34.410 172.560 ;
        RECT 34.060 172.545 34.410 172.550 ;
        RECT 34.075 172.540 34.410 172.545 ;
        RECT 34.775 172.540 35.035 172.990 ;
        RECT 35.665 172.650 35.955 173.815 ;
        RECT 37.085 172.675 37.315 173.815 ;
        RECT 37.485 172.665 37.815 173.645 ;
        RECT 37.985 172.675 38.195 173.815 ;
        RECT 38.725 173.175 39.055 173.605 ;
        RECT 38.600 173.005 39.055 173.175 ;
        RECT 39.235 173.175 39.485 173.595 ;
        RECT 39.715 173.345 40.045 173.815 ;
        RECT 40.275 173.175 40.525 173.595 ;
        RECT 39.235 173.005 40.525 173.175 ;
        RECT 34.075 172.535 35.035 172.540 ;
        RECT 34.085 172.525 35.035 172.535 ;
        RECT 34.095 172.520 35.035 172.525 ;
        RECT 34.105 172.510 35.035 172.520 ;
        RECT 34.110 172.500 35.035 172.510 ;
        RECT 34.115 172.495 35.035 172.500 ;
        RECT 34.125 172.480 35.035 172.495 ;
        RECT 34.130 172.465 35.035 172.480 ;
        RECT 34.140 172.440 35.035 172.465 ;
        RECT 33.645 171.970 33.975 172.395 ;
        RECT 33.725 171.945 33.975 171.970 ;
        RECT 32.905 171.435 33.165 171.915 ;
        RECT 33.335 171.265 33.585 171.805 ;
        RECT 33.755 171.485 33.975 171.945 ;
        RECT 34.145 172.370 35.035 172.440 ;
        RECT 34.145 171.645 34.315 172.370 ;
        RECT 37.065 172.255 37.395 172.505 ;
        RECT 34.485 171.815 35.035 172.200 ;
        RECT 34.145 171.475 35.035 171.645 ;
        RECT 35.665 171.265 35.955 171.990 ;
        RECT 37.085 171.265 37.315 172.085 ;
        RECT 37.565 172.065 37.815 172.665 ;
        RECT 37.485 171.435 37.815 172.065 ;
        RECT 37.985 171.265 38.195 172.085 ;
        RECT 38.600 172.005 38.770 173.005 ;
        RECT 38.940 172.175 39.185 172.835 ;
        RECT 39.400 172.175 39.665 172.835 ;
        RECT 39.860 172.175 40.145 172.835 ;
        RECT 40.320 172.505 40.535 172.835 ;
        RECT 40.715 172.675 40.965 173.815 ;
        RECT 41.135 172.755 41.465 173.605 ;
        RECT 40.320 172.175 40.625 172.505 ;
        RECT 40.795 172.175 41.105 172.505 ;
        RECT 40.795 172.005 40.965 172.175 ;
        RECT 38.600 171.835 40.965 172.005 ;
        RECT 41.275 171.990 41.465 172.755 ;
        RECT 41.650 173.425 41.985 173.645 ;
        RECT 42.990 173.435 43.345 173.815 ;
        RECT 41.650 172.805 41.905 173.425 ;
        RECT 42.155 173.265 42.385 173.305 ;
        RECT 43.515 173.265 43.765 173.645 ;
        RECT 42.155 173.065 43.765 173.265 ;
        RECT 42.155 172.975 42.340 173.065 ;
        RECT 42.930 173.055 43.765 173.065 ;
        RECT 44.015 173.035 44.265 173.815 ;
        RECT 44.435 172.965 44.695 173.645 ;
        RECT 44.865 173.305 46.055 173.595 ;
        RECT 42.495 172.865 42.825 172.895 ;
        RECT 42.495 172.805 44.295 172.865 ;
        RECT 41.650 172.695 44.355 172.805 ;
        RECT 41.650 172.635 42.825 172.695 ;
        RECT 44.155 172.660 44.355 172.695 ;
        RECT 41.645 172.255 42.135 172.455 ;
        RECT 42.325 172.255 42.800 172.465 ;
        RECT 38.755 171.265 39.085 171.665 ;
        RECT 39.255 171.495 39.585 171.835 ;
        RECT 40.635 171.265 40.965 171.665 ;
        RECT 41.135 171.480 41.465 171.990 ;
        RECT 41.650 171.265 42.105 172.030 ;
        RECT 42.580 171.855 42.800 172.255 ;
        RECT 43.045 172.255 43.375 172.465 ;
        RECT 43.045 171.855 43.255 172.255 ;
        RECT 43.545 172.220 43.955 172.525 ;
        RECT 44.185 172.085 44.355 172.660 ;
        RECT 44.085 171.965 44.355 172.085 ;
        RECT 43.510 171.920 44.355 171.965 ;
        RECT 43.510 171.795 44.265 171.920 ;
        RECT 43.510 171.645 43.680 171.795 ;
        RECT 44.525 171.765 44.695 172.965 ;
        RECT 44.885 172.965 46.055 173.135 ;
        RECT 46.225 173.015 46.505 173.815 ;
        RECT 44.885 172.675 45.210 172.965 ;
        RECT 45.885 172.845 46.055 172.965 ;
        RECT 45.380 172.505 45.575 172.795 ;
        RECT 45.885 172.675 46.545 172.845 ;
        RECT 46.715 172.675 46.990 173.645 ;
        RECT 47.255 173.145 47.425 173.645 ;
        RECT 47.595 173.315 47.925 173.815 ;
        RECT 47.255 172.975 47.920 173.145 ;
        RECT 46.375 172.505 46.545 172.675 ;
        RECT 44.865 172.175 45.210 172.505 ;
        RECT 45.380 172.175 46.205 172.505 ;
        RECT 46.375 172.175 46.650 172.505 ;
        RECT 46.375 172.005 46.545 172.175 ;
        RECT 42.380 171.435 43.680 171.645 ;
        RECT 43.935 171.265 44.265 171.625 ;
        RECT 44.435 171.435 44.695 171.765 ;
        RECT 44.880 171.835 46.545 172.005 ;
        RECT 46.820 171.940 46.990 172.675 ;
        RECT 47.170 172.155 47.520 172.805 ;
        RECT 47.690 171.985 47.920 172.975 ;
        RECT 44.880 171.485 45.135 171.835 ;
        RECT 45.305 171.265 45.635 171.665 ;
        RECT 45.805 171.485 45.975 171.835 ;
        RECT 46.145 171.265 46.525 171.665 ;
        RECT 46.715 171.595 46.990 171.940 ;
        RECT 47.255 171.815 47.920 171.985 ;
        RECT 47.255 171.525 47.425 171.815 ;
        RECT 47.595 171.265 47.925 171.645 ;
        RECT 48.095 171.525 48.280 173.645 ;
        RECT 48.520 173.355 48.785 173.815 ;
        RECT 48.955 173.220 49.205 173.645 ;
        RECT 49.415 173.370 50.520 173.540 ;
        RECT 48.900 173.090 49.205 173.220 ;
        RECT 48.450 171.895 48.730 172.845 ;
        RECT 48.900 171.985 49.070 173.090 ;
        RECT 49.240 172.305 49.480 172.900 ;
        RECT 49.650 172.835 50.180 173.200 ;
        RECT 49.650 172.135 49.820 172.835 ;
        RECT 50.350 172.755 50.520 173.370 ;
        RECT 50.690 173.015 50.860 173.815 ;
        RECT 51.030 173.315 51.280 173.645 ;
        RECT 51.505 173.345 52.390 173.515 ;
        RECT 50.350 172.665 50.860 172.755 ;
        RECT 48.900 171.855 49.125 171.985 ;
        RECT 49.295 171.915 49.820 172.135 ;
        RECT 49.990 172.495 50.860 172.665 ;
        RECT 48.535 171.265 48.785 171.725 ;
        RECT 48.955 171.715 49.125 171.855 ;
        RECT 49.990 171.715 50.160 172.495 ;
        RECT 50.690 172.425 50.860 172.495 ;
        RECT 50.370 172.245 50.570 172.275 ;
        RECT 51.030 172.245 51.200 173.315 ;
        RECT 51.370 172.425 51.560 173.145 ;
        RECT 50.370 171.945 51.200 172.245 ;
        RECT 51.730 172.215 52.050 173.175 ;
        RECT 48.955 171.545 49.290 171.715 ;
        RECT 49.485 171.545 50.160 171.715 ;
        RECT 50.480 171.265 50.850 171.765 ;
        RECT 51.030 171.715 51.200 171.945 ;
        RECT 51.585 171.885 52.050 172.215 ;
        RECT 52.220 172.505 52.390 173.345 ;
        RECT 52.570 173.315 52.885 173.815 ;
        RECT 53.115 173.085 53.455 173.645 ;
        RECT 52.560 172.710 53.455 173.085 ;
        RECT 53.625 172.805 53.795 173.815 ;
        RECT 53.265 172.505 53.455 172.710 ;
        RECT 53.965 172.755 54.295 173.600 ;
        RECT 53.965 172.675 54.355 172.755 ;
        RECT 54.525 172.725 55.735 173.815 ;
        RECT 54.140 172.625 54.355 172.675 ;
        RECT 52.220 172.175 53.095 172.505 ;
        RECT 53.265 172.175 54.015 172.505 ;
        RECT 52.220 171.715 52.390 172.175 ;
        RECT 53.265 172.005 53.465 172.175 ;
        RECT 54.185 172.045 54.355 172.625 ;
        RECT 54.130 172.005 54.355 172.045 ;
        RECT 51.030 171.545 51.435 171.715 ;
        RECT 51.605 171.545 52.390 171.715 ;
        RECT 52.665 171.265 52.875 171.795 ;
        RECT 53.135 171.480 53.465 172.005 ;
        RECT 53.975 171.920 54.355 172.005 ;
        RECT 54.525 172.015 55.045 172.555 ;
        RECT 55.215 172.185 55.735 172.725 ;
        RECT 55.905 172.675 56.290 173.645 ;
        RECT 56.460 173.355 56.785 173.815 ;
        RECT 57.305 173.185 57.585 173.645 ;
        RECT 56.460 172.965 57.585 173.185 ;
        RECT 53.635 171.265 53.805 171.875 ;
        RECT 53.975 171.485 54.305 171.920 ;
        RECT 54.525 171.265 55.735 172.015 ;
        RECT 55.905 172.005 56.185 172.675 ;
        RECT 56.460 172.505 56.910 172.965 ;
        RECT 57.775 172.795 58.175 173.645 ;
        RECT 58.575 173.355 58.845 173.815 ;
        RECT 59.015 173.185 59.300 173.645 ;
        RECT 56.355 172.175 56.910 172.505 ;
        RECT 57.080 172.235 58.175 172.795 ;
        RECT 56.460 172.065 56.910 172.175 ;
        RECT 55.905 171.435 56.290 172.005 ;
        RECT 56.460 171.895 57.585 172.065 ;
        RECT 56.460 171.265 56.785 171.725 ;
        RECT 57.305 171.435 57.585 171.895 ;
        RECT 57.775 171.435 58.175 172.235 ;
        RECT 58.345 172.965 59.300 173.185 ;
        RECT 58.345 172.065 58.555 172.965 ;
        RECT 58.725 172.235 59.415 172.795 ;
        RECT 59.585 172.725 61.255 173.815 ;
        RECT 58.345 171.895 59.300 172.065 ;
        RECT 58.575 171.265 58.845 171.725 ;
        RECT 59.015 171.435 59.300 171.895 ;
        RECT 59.585 172.035 60.335 172.555 ;
        RECT 60.505 172.205 61.255 172.725 ;
        RECT 61.425 172.650 61.715 173.815 ;
        RECT 61.885 172.675 62.270 173.645 ;
        RECT 62.440 173.355 62.765 173.815 ;
        RECT 63.285 173.185 63.565 173.645 ;
        RECT 62.440 172.965 63.565 173.185 ;
        RECT 59.585 171.265 61.255 172.035 ;
        RECT 61.885 172.005 62.165 172.675 ;
        RECT 62.440 172.505 62.890 172.965 ;
        RECT 63.755 172.795 64.155 173.645 ;
        RECT 64.555 173.355 64.825 173.815 ;
        RECT 64.995 173.185 65.280 173.645 ;
        RECT 62.335 172.175 62.890 172.505 ;
        RECT 63.060 172.235 64.155 172.795 ;
        RECT 62.440 172.065 62.890 172.175 ;
        RECT 61.425 171.265 61.715 171.990 ;
        RECT 61.885 171.435 62.270 172.005 ;
        RECT 62.440 171.895 63.565 172.065 ;
        RECT 62.440 171.265 62.765 171.725 ;
        RECT 63.285 171.435 63.565 171.895 ;
        RECT 63.755 171.435 64.155 172.235 ;
        RECT 64.325 172.965 65.280 173.185 ;
        RECT 64.325 172.065 64.535 172.965 ;
        RECT 64.705 172.235 65.395 172.795 ;
        RECT 65.565 172.725 67.235 173.815 ;
        RECT 67.495 173.145 67.665 173.645 ;
        RECT 67.835 173.315 68.165 173.815 ;
        RECT 67.495 172.975 68.160 173.145 ;
        RECT 64.325 171.895 65.280 172.065 ;
        RECT 64.555 171.265 64.825 171.725 ;
        RECT 64.995 171.435 65.280 171.895 ;
        RECT 65.565 172.035 66.315 172.555 ;
        RECT 66.485 172.205 67.235 172.725 ;
        RECT 67.410 172.155 67.760 172.805 ;
        RECT 65.565 171.265 67.235 172.035 ;
        RECT 67.930 171.985 68.160 172.975 ;
        RECT 67.495 171.815 68.160 171.985 ;
        RECT 67.495 171.525 67.665 171.815 ;
        RECT 67.835 171.265 68.165 171.645 ;
        RECT 68.335 171.525 68.520 173.645 ;
        RECT 68.760 173.355 69.025 173.815 ;
        RECT 69.195 173.220 69.445 173.645 ;
        RECT 69.655 173.370 70.760 173.540 ;
        RECT 69.140 173.090 69.445 173.220 ;
        RECT 68.690 171.895 68.970 172.845 ;
        RECT 69.140 171.985 69.310 173.090 ;
        RECT 69.480 172.305 69.720 172.900 ;
        RECT 69.890 172.835 70.420 173.200 ;
        RECT 69.890 172.135 70.060 172.835 ;
        RECT 70.590 172.755 70.760 173.370 ;
        RECT 70.930 173.015 71.100 173.815 ;
        RECT 71.270 173.315 71.520 173.645 ;
        RECT 71.745 173.345 72.630 173.515 ;
        RECT 70.590 172.665 71.100 172.755 ;
        RECT 69.140 171.855 69.365 171.985 ;
        RECT 69.535 171.915 70.060 172.135 ;
        RECT 70.230 172.495 71.100 172.665 ;
        RECT 68.775 171.265 69.025 171.725 ;
        RECT 69.195 171.715 69.365 171.855 ;
        RECT 70.230 171.715 70.400 172.495 ;
        RECT 70.930 172.425 71.100 172.495 ;
        RECT 70.610 172.245 70.810 172.275 ;
        RECT 71.270 172.245 71.440 173.315 ;
        RECT 71.610 172.425 71.800 173.145 ;
        RECT 70.610 171.945 71.440 172.245 ;
        RECT 71.970 172.215 72.290 173.175 ;
        RECT 69.195 171.545 69.530 171.715 ;
        RECT 69.725 171.545 70.400 171.715 ;
        RECT 70.720 171.265 71.090 171.765 ;
        RECT 71.270 171.715 71.440 171.945 ;
        RECT 71.825 171.885 72.290 172.215 ;
        RECT 72.460 172.505 72.630 173.345 ;
        RECT 72.810 173.315 73.125 173.815 ;
        RECT 73.355 173.085 73.695 173.645 ;
        RECT 72.800 172.710 73.695 173.085 ;
        RECT 73.865 172.805 74.035 173.815 ;
        RECT 73.505 172.505 73.695 172.710 ;
        RECT 74.205 172.755 74.535 173.600 ;
        RECT 74.770 173.390 75.105 173.815 ;
        RECT 75.275 173.210 75.460 173.615 ;
        RECT 74.795 173.035 75.460 173.210 ;
        RECT 75.665 173.035 75.995 173.815 ;
        RECT 74.205 172.675 74.595 172.755 ;
        RECT 74.380 172.625 74.595 172.675 ;
        RECT 72.460 172.175 73.335 172.505 ;
        RECT 73.505 172.175 74.255 172.505 ;
        RECT 72.460 171.715 72.630 172.175 ;
        RECT 73.505 172.005 73.705 172.175 ;
        RECT 74.425 172.045 74.595 172.625 ;
        RECT 74.370 172.005 74.595 172.045 ;
        RECT 71.270 171.545 71.675 171.715 ;
        RECT 71.845 171.545 72.630 171.715 ;
        RECT 72.905 171.265 73.115 171.795 ;
        RECT 73.375 171.480 73.705 172.005 ;
        RECT 74.215 171.920 74.595 172.005 ;
        RECT 74.795 172.005 75.135 173.035 ;
        RECT 76.165 172.845 76.435 173.615 ;
        RECT 76.695 173.145 76.865 173.645 ;
        RECT 77.035 173.315 77.365 173.815 ;
        RECT 76.695 172.975 77.360 173.145 ;
        RECT 75.305 172.675 76.435 172.845 ;
        RECT 75.305 172.175 75.555 172.675 ;
        RECT 73.875 171.265 74.045 171.875 ;
        RECT 74.215 171.485 74.545 171.920 ;
        RECT 74.795 171.835 75.480 172.005 ;
        RECT 75.735 171.925 76.095 172.505 ;
        RECT 74.770 171.265 75.105 171.665 ;
        RECT 75.275 171.435 75.480 171.835 ;
        RECT 76.265 171.765 76.435 172.675 ;
        RECT 76.610 172.155 76.960 172.805 ;
        RECT 77.130 171.985 77.360 172.975 ;
        RECT 75.690 171.265 75.965 171.745 ;
        RECT 76.175 171.435 76.435 171.765 ;
        RECT 76.695 171.815 77.360 171.985 ;
        RECT 76.695 171.525 76.865 171.815 ;
        RECT 77.035 171.265 77.365 171.645 ;
        RECT 77.535 171.525 77.720 173.645 ;
        RECT 77.960 173.355 78.225 173.815 ;
        RECT 78.395 173.220 78.645 173.645 ;
        RECT 78.855 173.370 79.960 173.540 ;
        RECT 78.340 173.090 78.645 173.220 ;
        RECT 77.890 171.895 78.170 172.845 ;
        RECT 78.340 171.985 78.510 173.090 ;
        RECT 78.680 172.305 78.920 172.900 ;
        RECT 79.090 172.835 79.620 173.200 ;
        RECT 79.090 172.135 79.260 172.835 ;
        RECT 79.790 172.755 79.960 173.370 ;
        RECT 80.130 173.015 80.300 173.815 ;
        RECT 80.470 173.315 80.720 173.645 ;
        RECT 80.945 173.345 81.830 173.515 ;
        RECT 79.790 172.665 80.300 172.755 ;
        RECT 78.340 171.855 78.565 171.985 ;
        RECT 78.735 171.915 79.260 172.135 ;
        RECT 79.430 172.495 80.300 172.665 ;
        RECT 77.975 171.265 78.225 171.725 ;
        RECT 78.395 171.715 78.565 171.855 ;
        RECT 79.430 171.715 79.600 172.495 ;
        RECT 80.130 172.425 80.300 172.495 ;
        RECT 79.810 172.245 80.010 172.275 ;
        RECT 80.470 172.245 80.640 173.315 ;
        RECT 80.810 172.425 81.000 173.145 ;
        RECT 79.810 171.945 80.640 172.245 ;
        RECT 81.170 172.215 81.490 173.175 ;
        RECT 78.395 171.545 78.730 171.715 ;
        RECT 78.925 171.545 79.600 171.715 ;
        RECT 79.920 171.265 80.290 171.765 ;
        RECT 80.470 171.715 80.640 171.945 ;
        RECT 81.025 171.885 81.490 172.215 ;
        RECT 81.660 172.505 81.830 173.345 ;
        RECT 82.010 173.315 82.325 173.815 ;
        RECT 82.555 173.085 82.895 173.645 ;
        RECT 82.000 172.710 82.895 173.085 ;
        RECT 83.065 172.805 83.235 173.815 ;
        RECT 82.705 172.505 82.895 172.710 ;
        RECT 83.405 172.755 83.735 173.600 ;
        RECT 83.970 172.845 84.245 173.645 ;
        RECT 84.415 173.015 84.745 173.815 ;
        RECT 84.915 173.475 86.055 173.645 ;
        RECT 84.915 172.845 85.085 173.475 ;
        RECT 83.405 172.675 83.795 172.755 ;
        RECT 83.580 172.625 83.795 172.675 ;
        RECT 83.970 172.635 85.085 172.845 ;
        RECT 85.255 172.845 85.585 173.305 ;
        RECT 85.755 173.015 86.055 173.475 ;
        RECT 85.255 172.625 86.015 172.845 ;
        RECT 87.185 172.650 87.475 173.815 ;
        RECT 87.645 172.945 87.920 173.645 ;
        RECT 88.090 173.270 88.345 173.815 ;
        RECT 88.515 173.305 88.995 173.645 ;
        RECT 89.170 173.260 89.775 173.815 ;
        RECT 89.160 173.160 89.775 173.260 ;
        RECT 89.160 173.135 89.345 173.160 ;
        RECT 81.660 172.175 82.535 172.505 ;
        RECT 82.705 172.175 83.455 172.505 ;
        RECT 81.660 171.715 81.830 172.175 ;
        RECT 82.705 172.005 82.905 172.175 ;
        RECT 83.625 172.045 83.795 172.625 ;
        RECT 83.970 172.255 84.690 172.455 ;
        RECT 84.860 172.255 85.630 172.455 ;
        RECT 85.800 172.085 86.015 172.625 ;
        RECT 83.570 172.005 83.795 172.045 ;
        RECT 80.470 171.545 80.875 171.715 ;
        RECT 81.045 171.545 81.830 171.715 ;
        RECT 82.105 171.265 82.315 171.795 ;
        RECT 82.575 171.480 82.905 172.005 ;
        RECT 83.415 171.920 83.795 172.005 ;
        RECT 83.075 171.265 83.245 171.875 ;
        RECT 83.415 171.485 83.745 171.920 ;
        RECT 83.970 171.265 84.245 172.085 ;
        RECT 84.415 171.915 86.015 172.085 ;
        RECT 84.415 171.905 85.585 171.915 ;
        RECT 84.415 171.435 84.745 171.905 ;
        RECT 84.915 171.265 85.085 171.735 ;
        RECT 85.255 171.435 85.585 171.905 ;
        RECT 85.755 171.265 86.045 171.735 ;
        RECT 87.185 171.265 87.475 171.990 ;
        RECT 87.645 171.915 87.815 172.945 ;
        RECT 88.090 172.815 88.845 173.065 ;
        RECT 89.015 172.890 89.345 173.135 ;
        RECT 88.090 172.780 88.860 172.815 ;
        RECT 88.090 172.770 88.875 172.780 ;
        RECT 87.985 172.755 88.880 172.770 ;
        RECT 87.985 172.740 88.900 172.755 ;
        RECT 87.985 172.730 88.920 172.740 ;
        RECT 87.985 172.720 88.945 172.730 ;
        RECT 87.985 172.690 89.015 172.720 ;
        RECT 87.985 172.660 89.035 172.690 ;
        RECT 87.985 172.630 89.055 172.660 ;
        RECT 87.985 172.605 89.085 172.630 ;
        RECT 87.985 172.570 89.120 172.605 ;
        RECT 87.985 172.565 89.150 172.570 ;
        RECT 87.985 172.170 88.215 172.565 ;
        RECT 88.760 172.560 89.150 172.565 ;
        RECT 88.785 172.550 89.150 172.560 ;
        RECT 88.800 172.545 89.150 172.550 ;
        RECT 88.815 172.540 89.150 172.545 ;
        RECT 89.515 172.540 89.775 172.990 ;
        RECT 88.815 172.535 89.775 172.540 ;
        RECT 88.825 172.525 89.775 172.535 ;
        RECT 88.835 172.520 89.775 172.525 ;
        RECT 88.845 172.510 89.775 172.520 ;
        RECT 88.850 172.500 89.775 172.510 ;
        RECT 88.855 172.495 89.775 172.500 ;
        RECT 88.865 172.480 89.775 172.495 ;
        RECT 88.870 172.465 89.775 172.480 ;
        RECT 88.880 172.440 89.775 172.465 ;
        RECT 88.385 171.970 88.715 172.395 ;
        RECT 87.645 171.435 87.905 171.915 ;
        RECT 88.075 171.265 88.325 171.805 ;
        RECT 88.495 171.485 88.715 171.970 ;
        RECT 88.885 172.370 89.775 172.440 ;
        RECT 89.945 172.740 90.215 173.645 ;
        RECT 90.385 173.055 90.715 173.815 ;
        RECT 90.895 172.885 91.065 173.645 ;
        RECT 88.885 171.645 89.055 172.370 ;
        RECT 89.225 171.815 89.775 172.200 ;
        RECT 89.945 171.940 90.115 172.740 ;
        RECT 90.400 172.715 91.065 172.885 ;
        RECT 91.325 172.725 92.995 173.815 ;
        RECT 90.400 172.570 90.570 172.715 ;
        RECT 90.285 172.240 90.570 172.570 ;
        RECT 90.400 171.985 90.570 172.240 ;
        RECT 90.805 172.165 91.135 172.535 ;
        RECT 91.325 172.035 92.075 172.555 ;
        RECT 92.245 172.205 92.995 172.725 ;
        RECT 93.170 172.675 93.505 173.645 ;
        RECT 93.675 172.675 93.845 173.815 ;
        RECT 94.015 173.475 96.045 173.645 ;
        RECT 88.885 171.475 89.775 171.645 ;
        RECT 89.945 171.435 90.205 171.940 ;
        RECT 90.400 171.815 91.065 171.985 ;
        RECT 90.385 171.265 90.715 171.645 ;
        RECT 90.895 171.435 91.065 171.815 ;
        RECT 91.325 171.265 92.995 172.035 ;
        RECT 93.170 172.005 93.340 172.675 ;
        RECT 94.015 172.505 94.185 173.475 ;
        RECT 93.510 172.175 93.765 172.505 ;
        RECT 93.990 172.175 94.185 172.505 ;
        RECT 94.355 173.135 95.480 173.305 ;
        RECT 93.595 172.005 93.765 172.175 ;
        RECT 94.355 172.005 94.525 173.135 ;
        RECT 93.170 171.435 93.425 172.005 ;
        RECT 93.595 171.835 94.525 172.005 ;
        RECT 94.695 172.795 95.705 172.965 ;
        RECT 94.695 171.995 94.865 172.795 ;
        RECT 94.350 171.800 94.525 171.835 ;
        RECT 93.595 171.265 93.925 171.665 ;
        RECT 94.350 171.435 94.880 171.800 ;
        RECT 95.070 171.775 95.345 172.595 ;
        RECT 95.065 171.605 95.345 171.775 ;
        RECT 95.070 171.435 95.345 171.605 ;
        RECT 95.515 171.435 95.705 172.795 ;
        RECT 95.875 172.810 96.045 173.475 ;
        RECT 96.215 173.055 96.385 173.815 ;
        RECT 96.620 173.055 97.135 173.465 ;
        RECT 95.875 172.620 96.625 172.810 ;
        RECT 96.795 172.245 97.135 173.055 ;
        RECT 97.305 172.725 98.975 173.815 ;
        RECT 95.905 172.075 97.135 172.245 ;
        RECT 95.885 171.265 96.395 171.800 ;
        RECT 96.615 171.470 96.860 172.075 ;
        RECT 97.305 172.035 98.055 172.555 ;
        RECT 98.225 172.205 98.975 172.725 ;
        RECT 99.605 172.845 99.915 173.645 ;
        RECT 100.085 173.015 100.395 173.815 ;
        RECT 100.565 173.185 100.825 173.645 ;
        RECT 100.995 173.355 101.250 173.815 ;
        RECT 101.425 173.185 101.685 173.645 ;
        RECT 100.565 173.015 101.685 173.185 ;
        RECT 99.605 172.675 100.635 172.845 ;
        RECT 97.305 171.265 98.975 172.035 ;
        RECT 99.605 171.765 99.775 172.675 ;
        RECT 99.945 171.935 100.295 172.505 ;
        RECT 100.465 172.425 100.635 172.675 ;
        RECT 101.425 172.765 101.685 173.015 ;
        RECT 101.855 172.945 102.140 173.815 ;
        RECT 102.455 172.885 102.625 173.645 ;
        RECT 102.805 173.055 103.135 173.815 ;
        RECT 101.425 172.595 102.180 172.765 ;
        RECT 102.455 172.715 103.120 172.885 ;
        RECT 103.305 172.740 103.575 173.645 ;
        RECT 103.835 173.145 104.005 173.645 ;
        RECT 104.175 173.315 104.505 173.815 ;
        RECT 103.835 172.975 104.500 173.145 ;
        RECT 100.465 172.255 101.605 172.425 ;
        RECT 101.775 172.085 102.180 172.595 ;
        RECT 102.950 172.570 103.120 172.715 ;
        RECT 102.385 172.165 102.715 172.535 ;
        RECT 102.950 172.240 103.235 172.570 ;
        RECT 100.530 171.915 102.180 172.085 ;
        RECT 102.950 171.985 103.120 172.240 ;
        RECT 99.605 171.435 99.905 171.765 ;
        RECT 100.075 171.265 100.350 171.745 ;
        RECT 100.530 171.525 100.825 171.915 ;
        RECT 100.995 171.265 101.250 171.745 ;
        RECT 101.425 171.525 101.685 171.915 ;
        RECT 102.455 171.815 103.120 171.985 ;
        RECT 103.405 171.940 103.575 172.740 ;
        RECT 103.750 172.155 104.100 172.805 ;
        RECT 104.270 171.985 104.500 172.975 ;
        RECT 101.855 171.265 102.135 171.745 ;
        RECT 102.455 171.435 102.625 171.815 ;
        RECT 102.805 171.265 103.135 171.645 ;
        RECT 103.315 171.435 103.575 171.940 ;
        RECT 103.835 171.815 104.500 171.985 ;
        RECT 103.835 171.525 104.005 171.815 ;
        RECT 104.175 171.265 104.505 171.645 ;
        RECT 104.675 171.525 104.860 173.645 ;
        RECT 105.100 173.355 105.365 173.815 ;
        RECT 105.535 173.220 105.785 173.645 ;
        RECT 105.995 173.370 107.100 173.540 ;
        RECT 105.480 173.090 105.785 173.220 ;
        RECT 105.030 171.895 105.310 172.845 ;
        RECT 105.480 171.985 105.650 173.090 ;
        RECT 105.820 172.305 106.060 172.900 ;
        RECT 106.230 172.835 106.760 173.200 ;
        RECT 106.230 172.135 106.400 172.835 ;
        RECT 106.930 172.755 107.100 173.370 ;
        RECT 107.270 173.015 107.440 173.815 ;
        RECT 107.610 173.315 107.860 173.645 ;
        RECT 108.085 173.345 108.970 173.515 ;
        RECT 106.930 172.665 107.440 172.755 ;
        RECT 105.480 171.855 105.705 171.985 ;
        RECT 105.875 171.915 106.400 172.135 ;
        RECT 106.570 172.495 107.440 172.665 ;
        RECT 105.115 171.265 105.365 171.725 ;
        RECT 105.535 171.715 105.705 171.855 ;
        RECT 106.570 171.715 106.740 172.495 ;
        RECT 107.270 172.425 107.440 172.495 ;
        RECT 106.950 172.245 107.150 172.275 ;
        RECT 107.610 172.245 107.780 173.315 ;
        RECT 107.950 172.425 108.140 173.145 ;
        RECT 106.950 171.945 107.780 172.245 ;
        RECT 108.310 172.215 108.630 173.175 ;
        RECT 105.535 171.545 105.870 171.715 ;
        RECT 106.065 171.545 106.740 171.715 ;
        RECT 107.060 171.265 107.430 171.765 ;
        RECT 107.610 171.715 107.780 171.945 ;
        RECT 108.165 171.885 108.630 172.215 ;
        RECT 108.800 172.505 108.970 173.345 ;
        RECT 109.150 173.315 109.465 173.815 ;
        RECT 109.695 173.085 110.035 173.645 ;
        RECT 109.140 172.710 110.035 173.085 ;
        RECT 110.205 172.805 110.375 173.815 ;
        RECT 109.845 172.505 110.035 172.710 ;
        RECT 110.545 172.755 110.875 173.600 ;
        RECT 111.655 172.885 111.825 173.645 ;
        RECT 112.005 173.055 112.335 173.815 ;
        RECT 110.545 172.675 110.935 172.755 ;
        RECT 111.655 172.715 112.320 172.885 ;
        RECT 112.505 172.740 112.775 173.645 ;
        RECT 110.720 172.625 110.935 172.675 ;
        RECT 108.800 172.175 109.675 172.505 ;
        RECT 109.845 172.175 110.595 172.505 ;
        RECT 108.800 171.715 108.970 172.175 ;
        RECT 109.845 172.005 110.045 172.175 ;
        RECT 110.765 172.045 110.935 172.625 ;
        RECT 112.150 172.570 112.320 172.715 ;
        RECT 111.585 172.165 111.915 172.535 ;
        RECT 112.150 172.240 112.435 172.570 ;
        RECT 110.710 172.005 110.935 172.045 ;
        RECT 107.610 171.545 108.015 171.715 ;
        RECT 108.185 171.545 108.970 171.715 ;
        RECT 109.245 171.265 109.455 171.795 ;
        RECT 109.715 171.480 110.045 172.005 ;
        RECT 110.555 171.920 110.935 172.005 ;
        RECT 112.150 171.985 112.320 172.240 ;
        RECT 110.215 171.265 110.385 171.875 ;
        RECT 110.555 171.485 110.885 171.920 ;
        RECT 111.655 171.815 112.320 171.985 ;
        RECT 112.605 171.940 112.775 172.740 ;
        RECT 112.945 172.650 113.235 173.815 ;
        RECT 113.495 173.145 113.665 173.645 ;
        RECT 113.835 173.315 114.165 173.815 ;
        RECT 113.495 172.975 114.160 173.145 ;
        RECT 113.410 172.155 113.760 172.805 ;
        RECT 111.655 171.435 111.825 171.815 ;
        RECT 112.005 171.265 112.335 171.645 ;
        RECT 112.515 171.435 112.775 171.940 ;
        RECT 112.945 171.265 113.235 171.990 ;
        RECT 113.930 171.985 114.160 172.975 ;
        RECT 113.495 171.815 114.160 171.985 ;
        RECT 113.495 171.525 113.665 171.815 ;
        RECT 113.835 171.265 114.165 171.645 ;
        RECT 114.335 171.525 114.520 173.645 ;
        RECT 114.760 173.355 115.025 173.815 ;
        RECT 115.195 173.220 115.445 173.645 ;
        RECT 115.655 173.370 116.760 173.540 ;
        RECT 115.140 173.090 115.445 173.220 ;
        RECT 114.690 171.895 114.970 172.845 ;
        RECT 115.140 171.985 115.310 173.090 ;
        RECT 115.480 172.305 115.720 172.900 ;
        RECT 115.890 172.835 116.420 173.200 ;
        RECT 115.890 172.135 116.060 172.835 ;
        RECT 116.590 172.755 116.760 173.370 ;
        RECT 116.930 173.015 117.100 173.815 ;
        RECT 117.270 173.315 117.520 173.645 ;
        RECT 117.745 173.345 118.630 173.515 ;
        RECT 116.590 172.665 117.100 172.755 ;
        RECT 115.140 171.855 115.365 171.985 ;
        RECT 115.535 171.915 116.060 172.135 ;
        RECT 116.230 172.495 117.100 172.665 ;
        RECT 114.775 171.265 115.025 171.725 ;
        RECT 115.195 171.715 115.365 171.855 ;
        RECT 116.230 171.715 116.400 172.495 ;
        RECT 116.930 172.425 117.100 172.495 ;
        RECT 116.610 172.245 116.810 172.275 ;
        RECT 117.270 172.245 117.440 173.315 ;
        RECT 117.610 172.425 117.800 173.145 ;
        RECT 116.610 171.945 117.440 172.245 ;
        RECT 117.970 172.215 118.290 173.175 ;
        RECT 115.195 171.545 115.530 171.715 ;
        RECT 115.725 171.545 116.400 171.715 ;
        RECT 116.720 171.265 117.090 171.765 ;
        RECT 117.270 171.715 117.440 171.945 ;
        RECT 117.825 171.885 118.290 172.215 ;
        RECT 118.460 172.505 118.630 173.345 ;
        RECT 118.810 173.315 119.125 173.815 ;
        RECT 119.355 173.085 119.695 173.645 ;
        RECT 118.800 172.710 119.695 173.085 ;
        RECT 119.865 172.805 120.035 173.815 ;
        RECT 119.505 172.505 119.695 172.710 ;
        RECT 120.205 172.755 120.535 173.600 ;
        RECT 120.765 173.095 121.225 173.645 ;
        RECT 121.415 173.095 121.745 173.815 ;
        RECT 120.205 172.675 120.595 172.755 ;
        RECT 120.380 172.625 120.595 172.675 ;
        RECT 118.460 172.175 119.335 172.505 ;
        RECT 119.505 172.175 120.255 172.505 ;
        RECT 118.460 171.715 118.630 172.175 ;
        RECT 119.505 172.005 119.705 172.175 ;
        RECT 120.425 172.045 120.595 172.625 ;
        RECT 120.370 172.005 120.595 172.045 ;
        RECT 117.270 171.545 117.675 171.715 ;
        RECT 117.845 171.545 118.630 171.715 ;
        RECT 118.905 171.265 119.115 171.795 ;
        RECT 119.375 171.480 119.705 172.005 ;
        RECT 120.215 171.920 120.595 172.005 ;
        RECT 119.875 171.265 120.045 171.875 ;
        RECT 120.215 171.485 120.545 171.920 ;
        RECT 120.765 171.725 121.015 173.095 ;
        RECT 121.945 172.925 122.245 173.475 ;
        RECT 122.415 173.145 122.695 173.815 ;
        RECT 121.305 172.755 122.245 172.925 ;
        RECT 121.305 172.505 121.475 172.755 ;
        RECT 122.615 172.505 122.880 172.865 ;
        RECT 123.525 172.635 123.845 173.815 ;
        RECT 124.015 172.795 124.215 173.585 ;
        RECT 124.540 172.985 124.925 173.645 ;
        RECT 125.320 173.055 126.105 173.815 ;
        RECT 124.515 172.885 124.925 172.985 ;
        RECT 124.015 172.625 124.345 172.795 ;
        RECT 124.515 172.675 126.125 172.885 ;
        RECT 121.185 172.175 121.475 172.505 ;
        RECT 121.645 172.255 121.985 172.505 ;
        RECT 122.205 172.255 122.880 172.505 ;
        RECT 124.165 172.505 124.345 172.625 ;
        RECT 123.525 172.255 123.990 172.455 ;
        RECT 124.165 172.255 124.495 172.505 ;
        RECT 124.665 172.455 125.130 172.505 ;
        RECT 124.665 172.285 125.135 172.455 ;
        RECT 124.665 172.255 125.130 172.285 ;
        RECT 125.325 172.255 125.680 172.505 ;
        RECT 121.305 172.085 121.475 172.175 ;
        RECT 121.305 171.895 122.695 172.085 ;
        RECT 125.850 172.075 126.125 172.675 ;
        RECT 120.765 171.435 121.325 171.725 ;
        RECT 121.495 171.265 121.745 171.725 ;
        RECT 122.365 171.535 122.695 171.895 ;
        RECT 123.525 171.875 124.705 172.045 ;
        RECT 123.525 171.460 123.865 171.875 ;
        RECT 124.035 171.265 124.205 171.705 ;
        RECT 124.375 171.655 124.705 171.875 ;
        RECT 124.875 171.895 126.125 172.075 ;
        RECT 124.875 171.825 125.240 171.895 ;
        RECT 124.375 171.475 125.625 171.655 ;
        RECT 125.895 171.265 126.065 171.725 ;
        RECT 126.295 171.545 126.575 173.645 ;
        RECT 126.765 172.975 127.020 173.645 ;
        RECT 127.190 173.055 127.520 173.815 ;
        RECT 127.690 173.215 127.940 173.645 ;
        RECT 128.110 173.395 128.465 173.815 ;
        RECT 128.655 173.475 129.825 173.645 ;
        RECT 128.655 173.435 128.985 173.475 ;
        RECT 129.095 173.215 129.325 173.305 ;
        RECT 127.690 172.975 129.325 173.215 ;
        RECT 129.495 172.975 129.825 173.475 ;
        RECT 126.765 172.965 126.975 172.975 ;
        RECT 126.765 171.845 126.935 172.965 ;
        RECT 129.995 172.805 130.165 173.645 ;
        RECT 131.435 173.145 131.605 173.645 ;
        RECT 131.775 173.315 132.105 173.815 ;
        RECT 131.435 172.975 132.100 173.145 ;
        RECT 127.105 172.635 130.165 172.805 ;
        RECT 127.105 172.085 127.275 172.635 ;
        RECT 127.495 172.285 127.870 172.455 ;
        RECT 127.505 172.255 127.870 172.285 ;
        RECT 128.040 172.255 128.370 172.455 ;
        RECT 127.105 171.915 127.905 172.085 ;
        RECT 126.765 171.765 126.950 171.845 ;
        RECT 126.765 171.435 127.020 171.765 ;
        RECT 127.235 171.265 127.565 171.745 ;
        RECT 127.735 171.685 127.905 171.915 ;
        RECT 128.085 171.855 128.370 172.255 ;
        RECT 128.640 172.255 129.115 172.455 ;
        RECT 129.285 172.255 129.730 172.455 ;
        RECT 129.900 172.255 130.250 172.465 ;
        RECT 128.640 171.855 128.920 172.255 ;
        RECT 131.350 172.155 131.700 172.805 ;
        RECT 129.100 171.915 130.165 172.085 ;
        RECT 131.870 171.985 132.100 172.975 ;
        RECT 129.100 171.685 129.270 171.915 ;
        RECT 127.735 171.435 129.270 171.685 ;
        RECT 129.495 171.265 129.825 171.745 ;
        RECT 129.995 171.435 130.165 171.915 ;
        RECT 131.435 171.815 132.100 171.985 ;
        RECT 131.435 171.525 131.605 171.815 ;
        RECT 131.775 171.265 132.105 171.645 ;
        RECT 132.275 171.525 132.460 173.645 ;
        RECT 132.700 173.355 132.965 173.815 ;
        RECT 133.135 173.220 133.385 173.645 ;
        RECT 133.595 173.370 134.700 173.540 ;
        RECT 133.080 173.090 133.385 173.220 ;
        RECT 132.630 171.895 132.910 172.845 ;
        RECT 133.080 171.985 133.250 173.090 ;
        RECT 133.420 172.305 133.660 172.900 ;
        RECT 133.830 172.835 134.360 173.200 ;
        RECT 133.830 172.135 134.000 172.835 ;
        RECT 134.530 172.755 134.700 173.370 ;
        RECT 134.870 173.015 135.040 173.815 ;
        RECT 135.210 173.315 135.460 173.645 ;
        RECT 135.685 173.345 136.570 173.515 ;
        RECT 134.530 172.665 135.040 172.755 ;
        RECT 133.080 171.855 133.305 171.985 ;
        RECT 133.475 171.915 134.000 172.135 ;
        RECT 134.170 172.495 135.040 172.665 ;
        RECT 132.715 171.265 132.965 171.725 ;
        RECT 133.135 171.715 133.305 171.855 ;
        RECT 134.170 171.715 134.340 172.495 ;
        RECT 134.870 172.425 135.040 172.495 ;
        RECT 134.550 172.245 134.750 172.275 ;
        RECT 135.210 172.245 135.380 173.315 ;
        RECT 135.550 172.425 135.740 173.145 ;
        RECT 134.550 171.945 135.380 172.245 ;
        RECT 135.910 172.215 136.230 173.175 ;
        RECT 133.135 171.545 133.470 171.715 ;
        RECT 133.665 171.545 134.340 171.715 ;
        RECT 134.660 171.265 135.030 171.765 ;
        RECT 135.210 171.715 135.380 171.945 ;
        RECT 135.765 171.885 136.230 172.215 ;
        RECT 136.400 172.505 136.570 173.345 ;
        RECT 136.750 173.315 137.065 173.815 ;
        RECT 137.295 173.085 137.635 173.645 ;
        RECT 136.740 172.710 137.635 173.085 ;
        RECT 137.805 172.805 137.975 173.815 ;
        RECT 137.445 172.505 137.635 172.710 ;
        RECT 138.145 172.755 138.475 173.600 ;
        RECT 138.145 172.675 138.535 172.755 ;
        RECT 138.320 172.625 138.535 172.675 ;
        RECT 138.705 172.650 138.995 173.815 ;
        RECT 140.145 172.755 140.475 173.600 ;
        RECT 140.645 172.805 140.815 173.815 ;
        RECT 140.985 173.085 141.325 173.645 ;
        RECT 141.555 173.315 141.870 173.815 ;
        RECT 142.050 173.345 142.935 173.515 ;
        RECT 140.085 172.675 140.475 172.755 ;
        RECT 140.985 172.710 141.880 173.085 ;
        RECT 136.400 172.175 137.275 172.505 ;
        RECT 137.445 172.175 138.195 172.505 ;
        RECT 136.400 171.715 136.570 172.175 ;
        RECT 137.445 172.005 137.645 172.175 ;
        RECT 138.365 172.045 138.535 172.625 ;
        RECT 138.310 172.005 138.535 172.045 ;
        RECT 135.210 171.545 135.615 171.715 ;
        RECT 135.785 171.545 136.570 171.715 ;
        RECT 136.845 171.265 137.055 171.795 ;
        RECT 137.315 171.480 137.645 172.005 ;
        RECT 138.155 171.920 138.535 172.005 ;
        RECT 140.085 172.625 140.300 172.675 ;
        RECT 140.085 172.045 140.255 172.625 ;
        RECT 140.985 172.505 141.175 172.710 ;
        RECT 142.050 172.505 142.220 173.345 ;
        RECT 143.160 173.315 143.410 173.645 ;
        RECT 140.425 172.175 141.175 172.505 ;
        RECT 141.345 172.175 142.220 172.505 ;
        RECT 140.085 172.005 140.310 172.045 ;
        RECT 140.975 172.005 141.175 172.175 ;
        RECT 137.815 171.265 137.985 171.875 ;
        RECT 138.155 171.485 138.485 171.920 ;
        RECT 138.705 171.265 138.995 171.990 ;
        RECT 140.085 171.920 140.465 172.005 ;
        RECT 140.135 171.485 140.465 171.920 ;
        RECT 140.635 171.265 140.805 171.875 ;
        RECT 140.975 171.480 141.305 172.005 ;
        RECT 141.565 171.265 141.775 171.795 ;
        RECT 142.050 171.715 142.220 172.175 ;
        RECT 142.390 172.215 142.710 173.175 ;
        RECT 142.880 172.425 143.070 173.145 ;
        RECT 143.240 172.245 143.410 173.315 ;
        RECT 143.580 173.015 143.750 173.815 ;
        RECT 143.920 173.370 145.025 173.540 ;
        RECT 143.920 172.755 144.090 173.370 ;
        RECT 145.235 173.220 145.485 173.645 ;
        RECT 145.655 173.355 145.920 173.815 ;
        RECT 144.260 172.835 144.790 173.200 ;
        RECT 145.235 173.090 145.540 173.220 ;
        RECT 143.580 172.665 144.090 172.755 ;
        RECT 143.580 172.495 144.450 172.665 ;
        RECT 143.580 172.425 143.750 172.495 ;
        RECT 143.870 172.245 144.070 172.275 ;
        RECT 142.390 171.885 142.855 172.215 ;
        RECT 143.240 171.945 144.070 172.245 ;
        RECT 143.240 171.715 143.410 171.945 ;
        RECT 142.050 171.545 142.835 171.715 ;
        RECT 143.005 171.545 143.410 171.715 ;
        RECT 143.590 171.265 143.960 171.765 ;
        RECT 144.280 171.715 144.450 172.495 ;
        RECT 144.620 172.135 144.790 172.835 ;
        RECT 144.960 172.305 145.200 172.900 ;
        RECT 144.620 171.915 145.145 172.135 ;
        RECT 145.370 171.985 145.540 173.090 ;
        RECT 145.315 171.855 145.540 171.985 ;
        RECT 145.710 171.895 145.990 172.845 ;
        RECT 145.315 171.715 145.485 171.855 ;
        RECT 144.280 171.545 144.955 171.715 ;
        RECT 145.150 171.545 145.485 171.715 ;
        RECT 145.655 171.265 145.905 171.725 ;
        RECT 146.160 171.525 146.345 173.645 ;
        RECT 146.515 173.315 146.845 173.815 ;
        RECT 147.015 173.145 147.185 173.645 ;
        RECT 146.520 172.975 147.185 173.145 ;
        RECT 147.455 173.225 147.715 173.615 ;
        RECT 147.885 173.405 148.215 173.815 ;
        RECT 147.455 173.025 148.215 173.225 ;
        RECT 146.520 171.985 146.750 172.975 ;
        RECT 146.920 172.155 147.270 172.805 ;
        RECT 147.465 172.155 147.695 172.845 ;
        RECT 147.875 172.345 148.215 173.025 ;
        RECT 148.405 172.525 148.735 173.635 ;
        RECT 148.905 172.905 149.095 173.635 ;
        RECT 149.265 173.085 149.595 173.815 ;
        RECT 149.775 172.905 149.945 173.635 ;
        RECT 148.905 172.705 149.945 172.905 ;
        RECT 150.205 172.725 151.875 173.815 ;
        RECT 146.520 171.815 147.185 171.985 ;
        RECT 147.875 171.895 148.105 172.345 ;
        RECT 148.405 172.225 148.940 172.525 ;
        RECT 146.515 171.265 146.845 171.645 ;
        RECT 147.015 171.525 147.185 171.815 ;
        RECT 147.725 171.445 148.105 171.895 ;
        RECT 148.285 171.265 148.515 172.045 ;
        RECT 148.695 171.975 148.940 172.225 ;
        RECT 149.120 172.175 149.515 172.525 ;
        RECT 149.710 172.175 150.000 172.525 ;
        RECT 148.695 171.445 149.125 171.975 ;
        RECT 149.305 171.555 149.515 172.175 ;
        RECT 150.205 172.035 150.955 172.555 ;
        RECT 151.125 172.205 151.875 172.725 ;
        RECT 152.565 172.675 152.775 173.815 ;
        RECT 152.945 172.665 153.275 173.645 ;
        RECT 153.445 172.675 153.675 173.815 ;
        RECT 153.885 172.725 155.555 173.815 ;
        RECT 149.685 171.265 150.015 171.995 ;
        RECT 150.205 171.265 151.875 172.035 ;
        RECT 152.565 171.265 152.775 172.085 ;
        RECT 152.945 172.065 153.195 172.665 ;
        RECT 153.365 172.255 153.695 172.505 ;
        RECT 152.945 171.435 153.275 172.065 ;
        RECT 153.445 171.265 153.675 172.085 ;
        RECT 153.885 172.035 154.635 172.555 ;
        RECT 154.805 172.205 155.555 172.725 ;
        RECT 155.725 172.725 156.935 173.815 ;
        RECT 155.725 172.185 156.245 172.725 ;
        RECT 153.885 171.265 155.555 172.035 ;
        RECT 156.415 172.015 156.935 172.555 ;
        RECT 155.725 171.265 156.935 172.015 ;
        RECT 22.700 171.095 157.020 171.265 ;
        RECT 22.785 170.345 23.995 171.095 ;
        RECT 24.255 170.545 24.425 170.835 ;
        RECT 24.595 170.715 24.925 171.095 ;
        RECT 24.255 170.375 24.920 170.545 ;
        RECT 22.785 169.805 23.305 170.345 ;
        RECT 23.475 169.635 23.995 170.175 ;
        RECT 22.785 168.545 23.995 169.635 ;
        RECT 24.170 169.555 24.520 170.205 ;
        RECT 24.690 169.385 24.920 170.375 ;
        RECT 24.255 169.215 24.920 169.385 ;
        RECT 24.255 168.715 24.425 169.215 ;
        RECT 24.595 168.545 24.925 169.045 ;
        RECT 25.095 168.715 25.280 170.835 ;
        RECT 25.535 170.635 25.785 171.095 ;
        RECT 25.955 170.645 26.290 170.815 ;
        RECT 26.485 170.645 27.160 170.815 ;
        RECT 25.955 170.505 26.125 170.645 ;
        RECT 25.450 169.515 25.730 170.465 ;
        RECT 25.900 170.375 26.125 170.505 ;
        RECT 25.900 169.270 26.070 170.375 ;
        RECT 26.295 170.225 26.820 170.445 ;
        RECT 26.240 169.460 26.480 170.055 ;
        RECT 26.650 169.525 26.820 170.225 ;
        RECT 26.990 169.865 27.160 170.645 ;
        RECT 27.480 170.595 27.850 171.095 ;
        RECT 28.030 170.645 28.435 170.815 ;
        RECT 28.605 170.645 29.390 170.815 ;
        RECT 28.030 170.415 28.200 170.645 ;
        RECT 27.370 170.115 28.200 170.415 ;
        RECT 28.585 170.145 29.050 170.475 ;
        RECT 27.370 170.085 27.570 170.115 ;
        RECT 27.690 169.865 27.860 169.935 ;
        RECT 26.990 169.695 27.860 169.865 ;
        RECT 27.350 169.605 27.860 169.695 ;
        RECT 25.900 169.140 26.205 169.270 ;
        RECT 26.650 169.160 27.180 169.525 ;
        RECT 25.520 168.545 25.785 169.005 ;
        RECT 25.955 168.715 26.205 169.140 ;
        RECT 27.350 168.990 27.520 169.605 ;
        RECT 26.415 168.820 27.520 168.990 ;
        RECT 27.690 168.545 27.860 169.345 ;
        RECT 28.030 169.045 28.200 170.115 ;
        RECT 28.370 169.215 28.560 169.935 ;
        RECT 28.730 169.185 29.050 170.145 ;
        RECT 29.220 170.185 29.390 170.645 ;
        RECT 29.665 170.565 29.875 171.095 ;
        RECT 30.135 170.355 30.465 170.880 ;
        RECT 30.635 170.485 30.805 171.095 ;
        RECT 30.975 170.440 31.305 170.875 ;
        RECT 32.470 170.445 32.780 170.915 ;
        RECT 32.950 170.615 33.685 171.095 ;
        RECT 33.855 170.525 34.025 170.875 ;
        RECT 34.195 170.695 34.575 171.095 ;
        RECT 30.975 170.355 31.355 170.440 ;
        RECT 30.265 170.185 30.465 170.355 ;
        RECT 31.130 170.315 31.355 170.355 ;
        RECT 29.220 169.855 30.095 170.185 ;
        RECT 30.265 169.855 31.015 170.185 ;
        RECT 28.030 168.715 28.280 169.045 ;
        RECT 29.220 169.015 29.390 169.855 ;
        RECT 30.265 169.650 30.455 169.855 ;
        RECT 31.185 169.735 31.355 170.315 ;
        RECT 32.470 170.275 33.205 170.445 ;
        RECT 33.855 170.355 34.595 170.525 ;
        RECT 34.765 170.420 35.035 170.765 ;
        RECT 32.955 170.185 33.205 170.275 ;
        RECT 34.425 170.185 34.595 170.355 ;
        RECT 32.450 169.855 32.785 170.105 ;
        RECT 32.955 169.855 33.695 170.185 ;
        RECT 34.425 169.855 34.655 170.185 ;
        RECT 31.140 169.685 31.355 169.735 ;
        RECT 29.560 169.275 30.455 169.650 ;
        RECT 30.965 169.605 31.355 169.685 ;
        RECT 28.505 168.845 29.390 169.015 ;
        RECT 29.570 168.545 29.885 169.045 ;
        RECT 30.115 168.715 30.455 169.275 ;
        RECT 30.625 168.545 30.795 169.555 ;
        RECT 30.965 168.760 31.295 169.605 ;
        RECT 32.450 168.545 32.705 169.685 ;
        RECT 32.955 169.295 33.125 169.855 ;
        RECT 34.425 169.685 34.595 169.855 ;
        RECT 34.865 169.685 35.035 170.420 ;
        RECT 35.210 170.330 35.665 171.095 ;
        RECT 35.940 170.715 37.240 170.925 ;
        RECT 37.495 170.735 37.825 171.095 ;
        RECT 37.070 170.565 37.240 170.715 ;
        RECT 37.995 170.595 38.255 170.925 ;
        RECT 38.025 170.585 38.255 170.595 ;
        RECT 36.140 170.105 36.360 170.505 ;
        RECT 35.205 169.905 35.695 170.105 ;
        RECT 35.885 169.895 36.360 170.105 ;
        RECT 36.605 170.105 36.815 170.505 ;
        RECT 37.070 170.440 37.825 170.565 ;
        RECT 37.070 170.395 37.915 170.440 ;
        RECT 37.645 170.275 37.915 170.395 ;
        RECT 36.605 169.895 36.935 170.105 ;
        RECT 37.105 169.835 37.515 170.140 ;
        RECT 33.350 169.515 34.595 169.685 ;
        RECT 33.350 169.265 33.770 169.515 ;
        RECT 32.900 168.765 34.095 169.095 ;
        RECT 34.275 168.545 34.555 169.345 ;
        RECT 34.765 168.715 35.035 169.685 ;
        RECT 35.210 169.665 36.385 169.725 ;
        RECT 37.745 169.700 37.915 170.275 ;
        RECT 37.715 169.665 37.915 169.700 ;
        RECT 35.210 169.555 37.915 169.665 ;
        RECT 35.210 168.935 35.465 169.555 ;
        RECT 36.055 169.495 37.855 169.555 ;
        RECT 36.055 169.465 36.385 169.495 ;
        RECT 38.085 169.395 38.255 170.585 ;
        RECT 38.425 170.345 39.635 171.095 ;
        RECT 39.805 170.755 40.410 170.925 ;
        RECT 39.805 170.585 40.495 170.755 ;
        RECT 38.425 169.805 38.945 170.345 ;
        RECT 39.805 170.295 40.410 170.585 ;
        RECT 39.115 169.635 39.635 170.175 ;
        RECT 35.715 169.295 35.900 169.385 ;
        RECT 36.490 169.295 37.325 169.305 ;
        RECT 35.715 169.095 37.325 169.295 ;
        RECT 35.715 169.055 35.945 169.095 ;
        RECT 35.210 168.715 35.545 168.935 ;
        RECT 36.550 168.545 36.905 168.925 ;
        RECT 37.075 168.715 37.325 169.095 ;
        RECT 37.575 168.545 37.825 169.325 ;
        RECT 37.995 168.715 38.255 169.395 ;
        RECT 38.425 168.545 39.635 169.635 ;
        RECT 39.805 169.395 40.035 170.295 ;
        RECT 40.205 169.565 40.535 170.105 ;
        RECT 40.745 169.565 41.075 170.925 ;
        RECT 41.470 170.555 41.815 170.925 ;
        RECT 42.005 170.725 42.335 171.095 ;
        RECT 42.505 170.555 42.835 170.925 ;
        RECT 41.470 170.355 42.835 170.555 ;
        RECT 43.025 170.295 43.720 170.925 ;
        RECT 43.925 170.295 44.235 171.095 ;
        RECT 44.405 170.325 47.915 171.095 ;
        RECT 48.545 170.370 48.835 171.095 ;
        RECT 49.555 170.445 49.725 170.925 ;
        RECT 49.905 170.615 50.145 171.095 ;
        RECT 50.395 170.445 50.565 170.925 ;
        RECT 50.735 170.615 51.065 171.095 ;
        RECT 51.235 170.445 51.405 170.925 ;
        RECT 41.245 169.565 41.535 170.185 ;
        RECT 41.705 169.565 42.335 170.185 ;
        RECT 42.505 169.565 42.835 170.175 ;
        RECT 43.045 169.855 43.380 170.105 ;
        RECT 43.550 169.695 43.720 170.295 ;
        RECT 43.890 169.855 44.225 170.125 ;
        RECT 44.405 169.805 46.055 170.325 ;
        RECT 49.555 170.275 50.190 170.445 ;
        RECT 50.395 170.275 51.405 170.445 ;
        RECT 51.575 170.295 51.905 171.095 ;
        RECT 52.225 170.595 52.485 170.925 ;
        RECT 52.655 170.735 52.985 171.095 ;
        RECT 53.240 170.715 54.540 170.925 ;
        RECT 52.225 170.585 52.455 170.595 ;
        RECT 39.805 169.155 41.815 169.395 ;
        RECT 40.010 168.545 40.340 168.985 ;
        RECT 40.510 168.715 40.745 169.155 ;
        RECT 40.930 168.545 41.260 168.925 ;
        RECT 41.470 168.715 41.815 169.155 ;
        RECT 41.990 168.810 42.335 169.565 ;
        RECT 42.505 168.545 42.835 169.385 ;
        RECT 43.025 168.545 43.285 169.685 ;
        RECT 43.455 168.715 43.785 169.695 ;
        RECT 43.955 168.545 44.235 169.685 ;
        RECT 46.225 169.635 47.915 170.155 ;
        RECT 50.020 170.105 50.190 170.275 ;
        RECT 49.470 169.865 49.850 170.105 ;
        RECT 50.020 169.935 50.520 170.105 ;
        RECT 50.910 170.075 51.405 170.275 ;
        RECT 44.405 168.545 47.915 169.635 ;
        RECT 48.545 168.545 48.835 169.710 ;
        RECT 50.020 169.695 50.190 169.935 ;
        RECT 50.905 169.905 51.405 170.075 ;
        RECT 50.910 169.735 51.405 169.905 ;
        RECT 49.475 169.525 50.190 169.695 ;
        RECT 50.395 169.565 51.405 169.735 ;
        RECT 49.475 168.715 49.805 169.525 ;
        RECT 49.975 168.545 50.215 169.345 ;
        RECT 50.395 168.715 50.565 169.565 ;
        RECT 50.735 168.545 51.065 169.345 ;
        RECT 51.235 168.715 51.405 169.565 ;
        RECT 51.575 168.545 51.905 169.695 ;
        RECT 52.225 169.395 52.395 170.585 ;
        RECT 53.240 170.565 53.410 170.715 ;
        RECT 52.655 170.440 53.410 170.565 ;
        RECT 52.565 170.395 53.410 170.440 ;
        RECT 52.565 170.275 52.835 170.395 ;
        RECT 52.565 169.700 52.735 170.275 ;
        RECT 52.965 169.835 53.375 170.140 ;
        RECT 53.665 170.105 53.875 170.505 ;
        RECT 53.545 169.895 53.875 170.105 ;
        RECT 54.120 170.105 54.340 170.505 ;
        RECT 54.815 170.330 55.270 171.095 ;
        RECT 55.450 170.330 55.905 171.095 ;
        RECT 56.180 170.715 57.480 170.925 ;
        RECT 57.735 170.735 58.065 171.095 ;
        RECT 57.310 170.565 57.480 170.715 ;
        RECT 58.235 170.595 58.495 170.925 ;
        RECT 58.265 170.585 58.495 170.595 ;
        RECT 56.380 170.105 56.600 170.505 ;
        RECT 54.120 169.895 54.595 170.105 ;
        RECT 54.785 169.905 55.275 170.105 ;
        RECT 55.445 169.905 55.935 170.105 ;
        RECT 56.125 169.895 56.600 170.105 ;
        RECT 56.845 170.105 57.055 170.505 ;
        RECT 57.310 170.440 58.065 170.565 ;
        RECT 57.310 170.395 58.155 170.440 ;
        RECT 57.885 170.275 58.155 170.395 ;
        RECT 56.845 169.895 57.175 170.105 ;
        RECT 57.345 169.835 57.755 170.140 ;
        RECT 52.565 169.665 52.765 169.700 ;
        RECT 54.095 169.665 55.270 169.725 ;
        RECT 52.565 169.555 55.270 169.665 ;
        RECT 52.625 169.495 54.425 169.555 ;
        RECT 54.095 169.465 54.425 169.495 ;
        RECT 52.225 168.715 52.485 169.395 ;
        RECT 52.655 168.545 52.905 169.325 ;
        RECT 53.155 169.295 53.990 169.305 ;
        RECT 54.580 169.295 54.765 169.385 ;
        RECT 53.155 169.095 54.765 169.295 ;
        RECT 53.155 168.715 53.405 169.095 ;
        RECT 54.535 169.055 54.765 169.095 ;
        RECT 55.015 168.935 55.270 169.555 ;
        RECT 53.575 168.545 53.930 168.925 ;
        RECT 54.935 168.715 55.270 168.935 ;
        RECT 55.450 169.665 56.625 169.725 ;
        RECT 57.985 169.700 58.155 170.275 ;
        RECT 57.955 169.665 58.155 169.700 ;
        RECT 55.450 169.555 58.155 169.665 ;
        RECT 55.450 168.935 55.705 169.555 ;
        RECT 56.295 169.495 58.095 169.555 ;
        RECT 56.295 169.465 56.625 169.495 ;
        RECT 58.325 169.395 58.495 170.585 ;
        RECT 58.715 170.440 59.045 170.875 ;
        RECT 59.215 170.485 59.385 171.095 ;
        RECT 58.665 170.355 59.045 170.440 ;
        RECT 59.555 170.355 59.885 170.880 ;
        RECT 60.145 170.565 60.355 171.095 ;
        RECT 60.630 170.645 61.415 170.815 ;
        RECT 61.585 170.645 61.990 170.815 ;
        RECT 58.665 170.315 58.890 170.355 ;
        RECT 58.665 169.735 58.835 170.315 ;
        RECT 59.555 170.185 59.755 170.355 ;
        RECT 60.630 170.185 60.800 170.645 ;
        RECT 59.005 169.855 59.755 170.185 ;
        RECT 59.925 169.855 60.800 170.185 ;
        RECT 58.665 169.685 58.880 169.735 ;
        RECT 58.665 169.605 59.055 169.685 ;
        RECT 55.955 169.295 56.140 169.385 ;
        RECT 56.730 169.295 57.565 169.305 ;
        RECT 55.955 169.095 57.565 169.295 ;
        RECT 55.955 169.055 56.185 169.095 ;
        RECT 55.450 168.715 55.785 168.935 ;
        RECT 56.790 168.545 57.145 168.925 ;
        RECT 57.315 168.715 57.565 169.095 ;
        RECT 57.815 168.545 58.065 169.325 ;
        RECT 58.235 168.715 58.495 169.395 ;
        RECT 58.725 168.760 59.055 169.605 ;
        RECT 59.565 169.650 59.755 169.855 ;
        RECT 59.225 168.545 59.395 169.555 ;
        RECT 59.565 169.275 60.460 169.650 ;
        RECT 59.565 168.715 59.905 169.275 ;
        RECT 60.135 168.545 60.450 169.045 ;
        RECT 60.630 169.015 60.800 169.855 ;
        RECT 60.970 170.145 61.435 170.475 ;
        RECT 61.820 170.415 61.990 170.645 ;
        RECT 62.170 170.595 62.540 171.095 ;
        RECT 62.860 170.645 63.535 170.815 ;
        RECT 63.730 170.645 64.065 170.815 ;
        RECT 60.970 169.185 61.290 170.145 ;
        RECT 61.820 170.115 62.650 170.415 ;
        RECT 61.460 169.215 61.650 169.935 ;
        RECT 61.820 169.045 61.990 170.115 ;
        RECT 62.450 170.085 62.650 170.115 ;
        RECT 62.160 169.865 62.330 169.935 ;
        RECT 62.860 169.865 63.030 170.645 ;
        RECT 63.895 170.505 64.065 170.645 ;
        RECT 64.235 170.635 64.485 171.095 ;
        RECT 62.160 169.695 63.030 169.865 ;
        RECT 63.200 170.225 63.725 170.445 ;
        RECT 63.895 170.375 64.120 170.505 ;
        RECT 62.160 169.605 62.670 169.695 ;
        RECT 60.630 168.845 61.515 169.015 ;
        RECT 61.740 168.715 61.990 169.045 ;
        RECT 62.160 168.545 62.330 169.345 ;
        RECT 62.500 168.990 62.670 169.605 ;
        RECT 63.200 169.525 63.370 170.225 ;
        RECT 62.840 169.160 63.370 169.525 ;
        RECT 63.540 169.460 63.780 170.055 ;
        RECT 63.950 169.270 64.120 170.375 ;
        RECT 64.290 169.515 64.570 170.465 ;
        RECT 63.815 169.140 64.120 169.270 ;
        RECT 62.500 168.820 63.605 168.990 ;
        RECT 63.815 168.715 64.065 169.140 ;
        RECT 64.235 168.545 64.500 169.005 ;
        RECT 64.740 168.715 64.925 170.835 ;
        RECT 65.095 170.715 65.425 171.095 ;
        RECT 65.595 170.545 65.765 170.835 ;
        RECT 65.100 170.375 65.765 170.545 ;
        RECT 65.100 169.385 65.330 170.375 ;
        RECT 66.025 170.325 69.535 171.095 ;
        RECT 65.500 169.555 65.850 170.205 ;
        RECT 66.025 169.805 67.675 170.325 ;
        RECT 67.845 169.635 69.535 170.155 ;
        RECT 65.100 169.215 65.765 169.385 ;
        RECT 65.095 168.545 65.425 169.045 ;
        RECT 65.595 168.715 65.765 169.215 ;
        RECT 66.025 168.545 69.535 169.635 ;
        RECT 69.715 168.725 69.975 170.915 ;
        RECT 70.235 170.725 70.905 171.095 ;
        RECT 71.085 170.545 71.395 170.915 ;
        RECT 70.165 170.345 71.395 170.545 ;
        RECT 70.165 169.675 70.455 170.345 ;
        RECT 71.575 170.165 71.805 170.805 ;
        RECT 71.985 170.365 72.275 171.095 ;
        RECT 72.465 170.325 74.135 171.095 ;
        RECT 74.305 170.370 74.595 171.095 ;
        RECT 74.765 170.325 78.275 171.095 ;
        RECT 70.635 169.855 71.100 170.165 ;
        RECT 71.280 169.855 71.805 170.165 ;
        RECT 71.985 169.855 72.285 170.185 ;
        RECT 72.465 169.805 73.215 170.325 ;
        RECT 70.165 169.455 70.935 169.675 ;
        RECT 70.145 168.545 70.485 169.275 ;
        RECT 70.665 168.725 70.935 169.455 ;
        RECT 71.115 169.435 72.275 169.675 ;
        RECT 73.385 169.635 74.135 170.155 ;
        RECT 74.765 169.805 76.415 170.325 ;
        RECT 71.115 168.725 71.345 169.435 ;
        RECT 71.515 168.545 71.845 169.255 ;
        RECT 72.015 168.725 72.275 169.435 ;
        RECT 72.465 168.545 74.135 169.635 ;
        RECT 74.305 168.545 74.595 169.710 ;
        RECT 76.585 169.635 78.275 170.155 ;
        RECT 74.765 168.545 78.275 169.635 ;
        RECT 78.915 168.725 79.175 170.915 ;
        RECT 79.435 170.725 80.105 171.095 ;
        RECT 80.285 170.545 80.595 170.915 ;
        RECT 79.365 170.345 80.595 170.545 ;
        RECT 79.365 169.675 79.655 170.345 ;
        RECT 80.775 170.165 81.005 170.805 ;
        RECT 81.185 170.365 81.475 171.095 ;
        RECT 82.860 170.285 83.105 170.890 ;
        RECT 83.325 170.560 83.835 171.095 ;
        RECT 79.835 169.855 80.300 170.165 ;
        RECT 80.480 169.855 81.005 170.165 ;
        RECT 81.185 169.855 81.485 170.185 ;
        RECT 82.585 170.115 83.815 170.285 ;
        RECT 79.365 169.455 80.135 169.675 ;
        RECT 79.345 168.545 79.685 169.275 ;
        RECT 79.865 168.725 80.135 169.455 ;
        RECT 80.315 169.435 81.475 169.675 ;
        RECT 80.315 168.725 80.545 169.435 ;
        RECT 80.715 168.545 81.045 169.255 ;
        RECT 81.215 168.725 81.475 169.435 ;
        RECT 82.585 169.305 82.925 170.115 ;
        RECT 83.095 169.550 83.845 169.740 ;
        RECT 82.585 168.895 83.100 169.305 ;
        RECT 83.335 168.545 83.505 169.305 ;
        RECT 83.675 168.885 83.845 169.550 ;
        RECT 84.015 169.565 84.205 170.925 ;
        RECT 84.375 170.075 84.650 170.925 ;
        RECT 84.840 170.560 85.370 170.925 ;
        RECT 85.795 170.695 86.125 171.095 ;
        RECT 85.195 170.525 85.370 170.560 ;
        RECT 84.375 169.905 84.655 170.075 ;
        RECT 84.375 169.765 84.650 169.905 ;
        RECT 84.855 169.565 85.025 170.365 ;
        RECT 84.015 169.395 85.025 169.565 ;
        RECT 85.195 170.355 86.125 170.525 ;
        RECT 86.295 170.355 86.550 170.925 ;
        RECT 86.815 170.545 86.985 170.835 ;
        RECT 87.155 170.715 87.485 171.095 ;
        RECT 86.815 170.375 87.480 170.545 ;
        RECT 85.195 169.225 85.365 170.355 ;
        RECT 85.955 170.185 86.125 170.355 ;
        RECT 84.240 169.055 85.365 169.225 ;
        RECT 85.535 169.855 85.730 170.185 ;
        RECT 85.955 169.855 86.210 170.185 ;
        RECT 85.535 168.885 85.705 169.855 ;
        RECT 86.380 169.685 86.550 170.355 ;
        RECT 83.675 168.715 85.705 168.885 ;
        RECT 85.875 168.545 86.045 169.685 ;
        RECT 86.215 168.715 86.550 169.685 ;
        RECT 86.730 169.555 87.080 170.205 ;
        RECT 87.250 169.385 87.480 170.375 ;
        RECT 86.815 169.215 87.480 169.385 ;
        RECT 86.815 168.715 86.985 169.215 ;
        RECT 87.155 168.545 87.485 169.045 ;
        RECT 87.655 168.715 87.840 170.835 ;
        RECT 88.095 170.635 88.345 171.095 ;
        RECT 88.515 170.645 88.850 170.815 ;
        RECT 89.045 170.645 89.720 170.815 ;
        RECT 88.515 170.505 88.685 170.645 ;
        RECT 88.010 169.515 88.290 170.465 ;
        RECT 88.460 170.375 88.685 170.505 ;
        RECT 88.460 169.270 88.630 170.375 ;
        RECT 88.855 170.225 89.380 170.445 ;
        RECT 88.800 169.460 89.040 170.055 ;
        RECT 89.210 169.525 89.380 170.225 ;
        RECT 89.550 169.865 89.720 170.645 ;
        RECT 90.040 170.595 90.410 171.095 ;
        RECT 90.590 170.645 90.995 170.815 ;
        RECT 91.165 170.645 91.950 170.815 ;
        RECT 90.590 170.415 90.760 170.645 ;
        RECT 89.930 170.115 90.760 170.415 ;
        RECT 91.145 170.145 91.610 170.475 ;
        RECT 89.930 170.085 90.130 170.115 ;
        RECT 90.250 169.865 90.420 169.935 ;
        RECT 89.550 169.695 90.420 169.865 ;
        RECT 89.910 169.605 90.420 169.695 ;
        RECT 88.460 169.140 88.765 169.270 ;
        RECT 89.210 169.160 89.740 169.525 ;
        RECT 88.080 168.545 88.345 169.005 ;
        RECT 88.515 168.715 88.765 169.140 ;
        RECT 89.910 168.990 90.080 169.605 ;
        RECT 88.975 168.820 90.080 168.990 ;
        RECT 90.250 168.545 90.420 169.345 ;
        RECT 90.590 169.045 90.760 170.115 ;
        RECT 90.930 169.215 91.120 169.935 ;
        RECT 91.290 169.185 91.610 170.145 ;
        RECT 91.780 170.185 91.950 170.645 ;
        RECT 92.225 170.565 92.435 171.095 ;
        RECT 92.695 170.355 93.025 170.880 ;
        RECT 93.195 170.485 93.365 171.095 ;
        RECT 93.535 170.440 93.865 170.875 ;
        RECT 93.535 170.355 93.915 170.440 ;
        RECT 92.825 170.185 93.025 170.355 ;
        RECT 93.690 170.315 93.915 170.355 ;
        RECT 91.780 169.855 92.655 170.185 ;
        RECT 92.825 169.855 93.575 170.185 ;
        RECT 90.590 168.715 90.840 169.045 ;
        RECT 91.780 169.015 91.950 169.855 ;
        RECT 92.825 169.650 93.015 169.855 ;
        RECT 93.745 169.735 93.915 170.315 ;
        RECT 94.085 170.325 95.755 171.095 ;
        RECT 96.385 170.420 96.645 170.925 ;
        RECT 96.825 170.715 97.155 171.095 ;
        RECT 97.335 170.545 97.505 170.925 ;
        RECT 94.085 169.805 94.835 170.325 ;
        RECT 93.700 169.685 93.915 169.735 ;
        RECT 92.120 169.275 93.015 169.650 ;
        RECT 93.525 169.605 93.915 169.685 ;
        RECT 95.005 169.635 95.755 170.155 ;
        RECT 91.065 168.845 91.950 169.015 ;
        RECT 92.130 168.545 92.445 169.045 ;
        RECT 92.675 168.715 93.015 169.275 ;
        RECT 93.185 168.545 93.355 169.555 ;
        RECT 93.525 168.760 93.855 169.605 ;
        RECT 94.085 168.545 95.755 169.635 ;
        RECT 96.385 169.620 96.555 170.420 ;
        RECT 96.840 170.375 97.505 170.545 ;
        RECT 97.965 170.465 98.295 170.825 ;
        RECT 98.915 170.635 99.165 171.095 ;
        RECT 99.335 170.635 99.895 170.925 ;
        RECT 96.840 170.120 97.010 170.375 ;
        RECT 97.965 170.275 99.355 170.465 ;
        RECT 96.725 169.790 97.010 170.120 ;
        RECT 97.245 169.825 97.575 170.195 ;
        RECT 99.185 170.185 99.355 170.275 ;
        RECT 97.780 169.855 98.455 170.105 ;
        RECT 98.675 169.855 99.015 170.105 ;
        RECT 99.185 169.855 99.475 170.185 ;
        RECT 96.840 169.645 97.010 169.790 ;
        RECT 96.385 168.715 96.655 169.620 ;
        RECT 96.840 169.475 97.505 169.645 ;
        RECT 97.780 169.495 98.045 169.855 ;
        RECT 99.185 169.605 99.355 169.855 ;
        RECT 96.825 168.545 97.155 169.305 ;
        RECT 97.335 168.715 97.505 169.475 ;
        RECT 98.415 169.435 99.355 169.605 ;
        RECT 97.965 168.545 98.245 169.215 ;
        RECT 98.415 168.885 98.715 169.435 ;
        RECT 99.645 169.265 99.895 170.635 ;
        RECT 100.065 170.370 100.355 171.095 ;
        RECT 100.530 170.355 100.785 170.925 ;
        RECT 100.955 170.695 101.285 171.095 ;
        RECT 101.710 170.560 102.240 170.925 ;
        RECT 101.710 170.525 101.885 170.560 ;
        RECT 100.955 170.355 101.885 170.525 ;
        RECT 98.915 168.545 99.245 169.265 ;
        RECT 99.435 168.715 99.895 169.265 ;
        RECT 100.065 168.545 100.355 169.710 ;
        RECT 100.530 169.685 100.700 170.355 ;
        RECT 100.955 170.185 101.125 170.355 ;
        RECT 100.870 169.855 101.125 170.185 ;
        RECT 101.350 169.855 101.545 170.185 ;
        RECT 100.530 168.715 100.865 169.685 ;
        RECT 101.035 168.545 101.205 169.685 ;
        RECT 101.375 168.885 101.545 169.855 ;
        RECT 101.715 169.225 101.885 170.355 ;
        RECT 102.055 169.565 102.225 170.365 ;
        RECT 102.430 170.075 102.705 170.925 ;
        RECT 102.425 169.905 102.705 170.075 ;
        RECT 102.430 169.765 102.705 169.905 ;
        RECT 102.875 169.565 103.065 170.925 ;
        RECT 103.245 170.560 103.755 171.095 ;
        RECT 103.975 170.285 104.220 170.890 ;
        RECT 105.130 170.355 105.385 170.925 ;
        RECT 105.555 170.695 105.885 171.095 ;
        RECT 106.310 170.560 106.840 170.925 ;
        RECT 106.310 170.525 106.485 170.560 ;
        RECT 105.555 170.355 106.485 170.525 ;
        RECT 107.030 170.415 107.305 170.925 ;
        RECT 103.265 170.115 104.495 170.285 ;
        RECT 102.055 169.395 103.065 169.565 ;
        RECT 103.235 169.550 103.985 169.740 ;
        RECT 101.715 169.055 102.840 169.225 ;
        RECT 103.235 168.885 103.405 169.550 ;
        RECT 104.155 169.305 104.495 170.115 ;
        RECT 101.375 168.715 103.405 168.885 ;
        RECT 103.575 168.545 103.745 169.305 ;
        RECT 103.980 168.895 104.495 169.305 ;
        RECT 105.130 169.685 105.300 170.355 ;
        RECT 105.555 170.185 105.725 170.355 ;
        RECT 105.470 169.855 105.725 170.185 ;
        RECT 105.950 169.855 106.145 170.185 ;
        RECT 105.130 168.715 105.465 169.685 ;
        RECT 105.635 168.545 105.805 169.685 ;
        RECT 105.975 168.885 106.145 169.855 ;
        RECT 106.315 169.225 106.485 170.355 ;
        RECT 106.655 169.565 106.825 170.365 ;
        RECT 107.025 170.245 107.305 170.415 ;
        RECT 107.030 169.765 107.305 170.245 ;
        RECT 107.475 169.565 107.665 170.925 ;
        RECT 107.845 170.560 108.355 171.095 ;
        RECT 108.575 170.285 108.820 170.890 ;
        RECT 109.265 170.325 111.855 171.095 ;
        RECT 112.030 170.355 112.285 170.925 ;
        RECT 112.455 170.695 112.785 171.095 ;
        RECT 113.210 170.560 113.740 170.925 ;
        RECT 113.210 170.525 113.385 170.560 ;
        RECT 112.455 170.355 113.385 170.525 ;
        RECT 107.865 170.115 109.095 170.285 ;
        RECT 106.655 169.395 107.665 169.565 ;
        RECT 107.835 169.550 108.585 169.740 ;
        RECT 106.315 169.055 107.440 169.225 ;
        RECT 107.835 168.885 108.005 169.550 ;
        RECT 108.755 169.305 109.095 170.115 ;
        RECT 109.265 169.805 110.475 170.325 ;
        RECT 110.645 169.635 111.855 170.155 ;
        RECT 105.975 168.715 108.005 168.885 ;
        RECT 108.175 168.545 108.345 169.305 ;
        RECT 108.580 168.895 109.095 169.305 ;
        RECT 109.265 168.545 111.855 169.635 ;
        RECT 112.030 169.685 112.200 170.355 ;
        RECT 112.455 170.185 112.625 170.355 ;
        RECT 112.370 169.855 112.625 170.185 ;
        RECT 112.850 169.855 113.045 170.185 ;
        RECT 112.030 168.715 112.365 169.685 ;
        RECT 112.535 168.545 112.705 169.685 ;
        RECT 112.875 168.885 113.045 169.855 ;
        RECT 113.215 169.225 113.385 170.355 ;
        RECT 113.555 169.565 113.725 170.365 ;
        RECT 113.930 170.075 114.205 170.925 ;
        RECT 113.925 169.905 114.205 170.075 ;
        RECT 113.930 169.765 114.205 169.905 ;
        RECT 114.375 169.565 114.565 170.925 ;
        RECT 114.745 170.560 115.255 171.095 ;
        RECT 115.475 170.285 115.720 170.890 ;
        RECT 117.175 170.545 117.345 170.925 ;
        RECT 117.525 170.715 117.855 171.095 ;
        RECT 117.175 170.375 117.840 170.545 ;
        RECT 118.035 170.420 118.295 170.925 ;
        RECT 114.765 170.115 115.995 170.285 ;
        RECT 113.555 169.395 114.565 169.565 ;
        RECT 114.735 169.550 115.485 169.740 ;
        RECT 113.215 169.055 114.340 169.225 ;
        RECT 114.735 168.885 114.905 169.550 ;
        RECT 115.655 169.305 115.995 170.115 ;
        RECT 117.105 169.825 117.435 170.195 ;
        RECT 117.670 170.120 117.840 170.375 ;
        RECT 117.670 169.790 117.955 170.120 ;
        RECT 117.670 169.645 117.840 169.790 ;
        RECT 112.875 168.715 114.905 168.885 ;
        RECT 115.075 168.545 115.245 169.305 ;
        RECT 115.480 168.895 115.995 169.305 ;
        RECT 117.175 169.475 117.840 169.645 ;
        RECT 118.125 169.620 118.295 170.420 ;
        RECT 118.555 170.545 118.725 170.835 ;
        RECT 118.895 170.715 119.225 171.095 ;
        RECT 118.555 170.375 119.220 170.545 ;
        RECT 117.175 168.715 117.345 169.475 ;
        RECT 117.525 168.545 117.855 169.305 ;
        RECT 118.025 168.715 118.295 169.620 ;
        RECT 118.470 169.555 118.820 170.205 ;
        RECT 118.990 169.385 119.220 170.375 ;
        RECT 118.555 169.215 119.220 169.385 ;
        RECT 118.555 168.715 118.725 169.215 ;
        RECT 118.895 168.545 119.225 169.045 ;
        RECT 119.395 168.715 119.580 170.835 ;
        RECT 119.835 170.635 120.085 171.095 ;
        RECT 120.255 170.645 120.590 170.815 ;
        RECT 120.785 170.645 121.460 170.815 ;
        RECT 120.255 170.505 120.425 170.645 ;
        RECT 119.750 169.515 120.030 170.465 ;
        RECT 120.200 170.375 120.425 170.505 ;
        RECT 120.200 169.270 120.370 170.375 ;
        RECT 120.595 170.225 121.120 170.445 ;
        RECT 120.540 169.460 120.780 170.055 ;
        RECT 120.950 169.525 121.120 170.225 ;
        RECT 121.290 169.865 121.460 170.645 ;
        RECT 121.780 170.595 122.150 171.095 ;
        RECT 122.330 170.645 122.735 170.815 ;
        RECT 122.905 170.645 123.690 170.815 ;
        RECT 122.330 170.415 122.500 170.645 ;
        RECT 121.670 170.115 122.500 170.415 ;
        RECT 122.885 170.145 123.350 170.475 ;
        RECT 121.670 170.085 121.870 170.115 ;
        RECT 121.990 169.865 122.160 169.935 ;
        RECT 121.290 169.695 122.160 169.865 ;
        RECT 121.650 169.605 122.160 169.695 ;
        RECT 120.200 169.140 120.505 169.270 ;
        RECT 120.950 169.160 121.480 169.525 ;
        RECT 119.820 168.545 120.085 169.005 ;
        RECT 120.255 168.715 120.505 169.140 ;
        RECT 121.650 168.990 121.820 169.605 ;
        RECT 120.715 168.820 121.820 168.990 ;
        RECT 121.990 168.545 122.160 169.345 ;
        RECT 122.330 169.045 122.500 170.115 ;
        RECT 122.670 169.215 122.860 169.935 ;
        RECT 123.030 169.185 123.350 170.145 ;
        RECT 123.520 170.185 123.690 170.645 ;
        RECT 123.965 170.565 124.175 171.095 ;
        RECT 124.435 170.355 124.765 170.880 ;
        RECT 124.935 170.485 125.105 171.095 ;
        RECT 125.275 170.440 125.605 170.875 ;
        RECT 125.275 170.355 125.655 170.440 ;
        RECT 125.825 170.370 126.115 171.095 ;
        RECT 124.565 170.185 124.765 170.355 ;
        RECT 125.430 170.315 125.655 170.355 ;
        RECT 123.520 169.855 124.395 170.185 ;
        RECT 124.565 169.855 125.315 170.185 ;
        RECT 122.330 168.715 122.580 169.045 ;
        RECT 123.520 169.015 123.690 169.855 ;
        RECT 124.565 169.650 124.755 169.855 ;
        RECT 125.485 169.735 125.655 170.315 ;
        RECT 125.440 169.685 125.655 169.735 ;
        RECT 123.860 169.275 124.755 169.650 ;
        RECT 125.265 169.605 125.655 169.685 ;
        RECT 122.805 168.845 123.690 169.015 ;
        RECT 123.870 168.545 124.185 169.045 ;
        RECT 124.415 168.715 124.755 169.275 ;
        RECT 124.925 168.545 125.095 169.555 ;
        RECT 125.265 168.760 125.595 169.605 ;
        RECT 125.825 168.545 126.115 169.710 ;
        RECT 126.285 168.715 126.565 170.815 ;
        RECT 126.795 170.635 126.965 171.095 ;
        RECT 127.235 170.705 128.485 170.885 ;
        RECT 127.620 170.465 127.985 170.535 ;
        RECT 126.735 170.285 127.985 170.465 ;
        RECT 128.155 170.485 128.485 170.705 ;
        RECT 128.655 170.655 128.825 171.095 ;
        RECT 128.995 170.485 129.335 170.900 ;
        RECT 128.155 170.315 129.335 170.485 ;
        RECT 129.505 170.595 129.765 170.925 ;
        RECT 129.935 170.735 130.265 171.095 ;
        RECT 130.520 170.715 131.820 170.925 ;
        RECT 129.505 170.585 129.735 170.595 ;
        RECT 126.735 169.685 127.010 170.285 ;
        RECT 127.180 169.855 127.535 170.105 ;
        RECT 127.730 170.075 128.195 170.105 ;
        RECT 127.725 169.905 128.195 170.075 ;
        RECT 127.730 169.855 128.195 169.905 ;
        RECT 128.365 169.855 128.695 170.105 ;
        RECT 128.870 169.905 129.335 170.105 ;
        RECT 128.515 169.735 128.695 169.855 ;
        RECT 126.735 169.475 128.345 169.685 ;
        RECT 128.515 169.565 128.845 169.735 ;
        RECT 127.935 169.375 128.345 169.475 ;
        RECT 126.755 168.545 127.540 169.305 ;
        RECT 127.935 168.715 128.320 169.375 ;
        RECT 128.645 168.775 128.845 169.565 ;
        RECT 129.015 168.545 129.335 169.725 ;
        RECT 129.505 169.395 129.675 170.585 ;
        RECT 130.520 170.565 130.690 170.715 ;
        RECT 129.935 170.440 130.690 170.565 ;
        RECT 129.845 170.395 130.690 170.440 ;
        RECT 129.845 170.275 130.115 170.395 ;
        RECT 129.845 169.700 130.015 170.275 ;
        RECT 130.245 169.835 130.655 170.140 ;
        RECT 130.945 170.105 131.155 170.505 ;
        RECT 130.825 169.895 131.155 170.105 ;
        RECT 131.400 170.105 131.620 170.505 ;
        RECT 132.095 170.330 132.550 171.095 ;
        RECT 132.725 170.550 138.070 171.095 ;
        RECT 131.400 169.895 131.875 170.105 ;
        RECT 132.065 169.905 132.555 170.105 ;
        RECT 129.845 169.665 130.045 169.700 ;
        RECT 131.375 169.665 132.550 169.725 ;
        RECT 134.310 169.720 134.650 170.550 ;
        RECT 138.305 170.275 138.515 171.095 ;
        RECT 138.685 170.295 139.015 170.925 ;
        RECT 129.845 169.555 132.550 169.665 ;
        RECT 129.905 169.495 131.705 169.555 ;
        RECT 131.375 169.465 131.705 169.495 ;
        RECT 129.505 168.715 129.765 169.395 ;
        RECT 129.935 168.545 130.185 169.325 ;
        RECT 130.435 169.295 131.270 169.305 ;
        RECT 131.860 169.295 132.045 169.385 ;
        RECT 130.435 169.095 132.045 169.295 ;
        RECT 130.435 168.715 130.685 169.095 ;
        RECT 131.815 169.055 132.045 169.095 ;
        RECT 132.295 168.935 132.550 169.555 ;
        RECT 136.130 168.980 136.480 170.230 ;
        RECT 138.685 169.695 138.935 170.295 ;
        RECT 139.185 170.275 139.415 171.095 ;
        RECT 139.625 170.325 141.295 171.095 ;
        RECT 141.465 170.715 142.355 170.885 ;
        RECT 139.105 169.855 139.435 170.105 ;
        RECT 139.625 169.805 140.375 170.325 ;
        RECT 141.465 170.160 142.015 170.545 ;
        RECT 130.855 168.545 131.210 168.925 ;
        RECT 132.215 168.715 132.550 168.935 ;
        RECT 132.725 168.545 138.070 168.980 ;
        RECT 138.305 168.545 138.515 169.685 ;
        RECT 138.685 168.715 139.015 169.695 ;
        RECT 139.185 168.545 139.415 169.685 ;
        RECT 140.545 169.635 141.295 170.155 ;
        RECT 142.185 169.990 142.355 170.715 ;
        RECT 139.625 168.545 141.295 169.635 ;
        RECT 141.465 169.920 142.355 169.990 ;
        RECT 142.525 170.415 142.745 170.875 ;
        RECT 142.915 170.555 143.165 171.095 ;
        RECT 143.335 170.445 143.595 170.925 ;
        RECT 143.765 170.550 149.110 171.095 ;
        RECT 142.525 170.390 142.775 170.415 ;
        RECT 142.525 169.965 142.855 170.390 ;
        RECT 141.465 169.895 142.360 169.920 ;
        RECT 141.465 169.880 142.370 169.895 ;
        RECT 141.465 169.865 142.375 169.880 ;
        RECT 141.465 169.860 142.385 169.865 ;
        RECT 141.465 169.850 142.390 169.860 ;
        RECT 141.465 169.840 142.395 169.850 ;
        RECT 141.465 169.835 142.405 169.840 ;
        RECT 141.465 169.825 142.415 169.835 ;
        RECT 141.465 169.820 142.425 169.825 ;
        RECT 141.465 169.370 141.725 169.820 ;
        RECT 142.090 169.815 142.425 169.820 ;
        RECT 142.090 169.810 142.440 169.815 ;
        RECT 142.090 169.800 142.455 169.810 ;
        RECT 142.090 169.795 142.480 169.800 ;
        RECT 143.025 169.795 143.255 170.190 ;
        RECT 142.090 169.790 143.255 169.795 ;
        RECT 142.120 169.755 143.255 169.790 ;
        RECT 142.155 169.730 143.255 169.755 ;
        RECT 142.185 169.700 143.255 169.730 ;
        RECT 142.205 169.670 143.255 169.700 ;
        RECT 142.225 169.640 143.255 169.670 ;
        RECT 142.295 169.630 143.255 169.640 ;
        RECT 142.320 169.620 143.255 169.630 ;
        RECT 142.340 169.605 143.255 169.620 ;
        RECT 142.360 169.590 143.255 169.605 ;
        RECT 142.365 169.580 143.150 169.590 ;
        RECT 142.380 169.545 143.150 169.580 ;
        RECT 141.895 169.225 142.225 169.470 ;
        RECT 142.395 169.295 143.150 169.545 ;
        RECT 143.425 169.415 143.595 170.445 ;
        RECT 145.350 169.720 145.690 170.550 ;
        RECT 149.285 170.325 150.955 171.095 ;
        RECT 151.585 170.370 151.875 171.095 ;
        RECT 152.045 170.355 152.430 170.925 ;
        RECT 152.600 170.635 152.925 171.095 ;
        RECT 153.445 170.465 153.725 170.925 ;
        RECT 141.895 169.200 142.080 169.225 ;
        RECT 141.465 169.100 142.080 169.200 ;
        RECT 141.465 168.545 142.070 169.100 ;
        RECT 142.245 168.715 142.725 169.055 ;
        RECT 142.895 168.545 143.150 169.090 ;
        RECT 143.320 168.715 143.595 169.415 ;
        RECT 147.170 168.980 147.520 170.230 ;
        RECT 149.285 169.805 150.035 170.325 ;
        RECT 150.205 169.635 150.955 170.155 ;
        RECT 143.765 168.545 149.110 168.980 ;
        RECT 149.285 168.545 150.955 169.635 ;
        RECT 151.585 168.545 151.875 169.710 ;
        RECT 152.045 169.685 152.325 170.355 ;
        RECT 152.600 170.295 153.725 170.465 ;
        RECT 152.600 170.185 153.050 170.295 ;
        RECT 152.495 169.855 153.050 170.185 ;
        RECT 153.915 170.125 154.315 170.925 ;
        RECT 154.715 170.635 154.985 171.095 ;
        RECT 155.155 170.465 155.440 170.925 ;
        RECT 152.045 168.715 152.430 169.685 ;
        RECT 152.600 169.395 153.050 169.855 ;
        RECT 153.220 169.565 154.315 170.125 ;
        RECT 152.600 169.175 153.725 169.395 ;
        RECT 152.600 168.545 152.925 169.005 ;
        RECT 153.445 168.715 153.725 169.175 ;
        RECT 153.915 168.715 154.315 169.565 ;
        RECT 154.485 170.295 155.440 170.465 ;
        RECT 155.725 170.345 156.935 171.095 ;
        RECT 154.485 169.395 154.695 170.295 ;
        RECT 154.865 169.565 155.555 170.125 ;
        RECT 155.725 169.635 156.245 170.175 ;
        RECT 156.415 169.805 156.935 170.345 ;
        RECT 154.485 169.175 155.440 169.395 ;
        RECT 154.715 168.545 154.985 169.005 ;
        RECT 155.155 168.715 155.440 169.175 ;
        RECT 155.725 168.545 156.935 169.635 ;
        RECT 22.700 168.375 157.020 168.545 ;
        RECT 22.785 167.285 23.995 168.375 ;
        RECT 24.165 167.940 29.510 168.375 ;
        RECT 22.785 166.575 23.305 167.115 ;
        RECT 23.475 166.745 23.995 167.285 ;
        RECT 22.785 165.825 23.995 166.575 ;
        RECT 25.750 166.370 26.090 167.200 ;
        RECT 27.570 166.690 27.920 167.940 ;
        RECT 29.685 167.285 31.355 168.375 ;
        RECT 29.685 166.595 30.435 167.115 ;
        RECT 30.605 166.765 31.355 167.285 ;
        RECT 31.985 167.945 32.325 168.205 ;
        RECT 24.165 165.825 29.510 166.370 ;
        RECT 29.685 165.825 31.355 166.595 ;
        RECT 31.985 166.545 32.245 167.945 ;
        RECT 32.495 167.575 32.825 168.375 ;
        RECT 33.290 167.405 33.540 168.205 ;
        RECT 33.725 167.655 34.055 168.375 ;
        RECT 34.275 167.405 34.525 168.205 ;
        RECT 34.695 167.995 35.030 168.375 ;
        RECT 32.435 167.235 34.625 167.405 ;
        RECT 32.435 167.065 32.750 167.235 ;
        RECT 32.420 166.815 32.750 167.065 ;
        RECT 31.985 166.035 32.325 166.545 ;
        RECT 32.495 165.825 32.765 166.625 ;
        RECT 32.945 166.095 33.225 167.065 ;
        RECT 33.405 166.095 33.705 167.065 ;
        RECT 33.885 166.100 34.235 167.065 ;
        RECT 34.455 166.325 34.625 167.235 ;
        RECT 34.795 166.505 35.035 167.815 ;
        RECT 35.665 167.210 35.955 168.375 ;
        RECT 36.130 167.235 36.385 168.375 ;
        RECT 36.580 167.825 37.775 168.155 ;
        RECT 36.635 167.065 36.805 167.625 ;
        RECT 37.030 167.405 37.450 167.655 ;
        RECT 37.955 167.575 38.235 168.375 ;
        RECT 37.030 167.235 38.275 167.405 ;
        RECT 38.445 167.235 38.715 168.205 ;
        RECT 38.885 167.285 42.395 168.375 ;
        RECT 38.105 167.065 38.275 167.235 ;
        RECT 36.130 166.815 36.465 167.065 ;
        RECT 36.635 166.735 37.375 167.065 ;
        RECT 38.105 166.735 38.335 167.065 ;
        RECT 36.635 166.645 36.885 166.735 ;
        RECT 34.455 165.995 34.950 166.325 ;
        RECT 35.665 165.825 35.955 166.550 ;
        RECT 36.150 166.475 36.885 166.645 ;
        RECT 38.105 166.565 38.275 166.735 ;
        RECT 36.150 166.005 36.460 166.475 ;
        RECT 37.535 166.395 38.275 166.565 ;
        RECT 38.545 166.500 38.715 167.235 ;
        RECT 36.630 165.825 37.365 166.305 ;
        RECT 37.535 166.045 37.705 166.395 ;
        RECT 37.875 165.825 38.255 166.225 ;
        RECT 38.445 166.155 38.715 166.500 ;
        RECT 38.885 166.595 40.535 167.115 ;
        RECT 40.705 166.765 42.395 167.285 ;
        RECT 42.585 167.485 42.845 168.195 ;
        RECT 43.015 167.665 43.345 168.375 ;
        RECT 43.515 167.485 43.745 168.195 ;
        RECT 42.585 167.245 43.745 167.485 ;
        RECT 43.925 167.465 44.195 168.195 ;
        RECT 44.375 167.645 44.715 168.375 ;
        RECT 43.925 167.245 44.695 167.465 ;
        RECT 42.575 166.735 42.875 167.065 ;
        RECT 43.055 166.755 43.580 167.065 ;
        RECT 43.760 166.755 44.225 167.065 ;
        RECT 38.885 165.825 42.395 166.595 ;
        RECT 42.585 165.825 42.875 166.555 ;
        RECT 43.055 166.115 43.285 166.755 ;
        RECT 44.405 166.575 44.695 167.245 ;
        RECT 43.465 166.375 44.695 166.575 ;
        RECT 43.465 166.005 43.775 166.375 ;
        RECT 43.955 165.825 44.625 166.195 ;
        RECT 44.885 166.005 45.145 168.195 ;
        RECT 45.330 167.235 45.605 168.205 ;
        RECT 45.815 167.575 46.095 168.375 ;
        RECT 46.265 167.865 47.455 168.155 ;
        RECT 47.715 167.705 47.885 168.205 ;
        RECT 48.055 167.875 48.385 168.375 ;
        RECT 46.265 167.525 47.435 167.695 ;
        RECT 47.715 167.535 48.380 167.705 ;
        RECT 46.265 167.405 46.435 167.525 ;
        RECT 45.775 167.235 46.435 167.405 ;
        RECT 45.330 166.500 45.500 167.235 ;
        RECT 45.775 167.065 45.945 167.235 ;
        RECT 46.745 167.065 46.940 167.355 ;
        RECT 47.110 167.235 47.435 167.525 ;
        RECT 45.670 166.735 45.945 167.065 ;
        RECT 46.115 166.735 46.940 167.065 ;
        RECT 47.110 166.735 47.455 167.065 ;
        RECT 45.775 166.565 45.945 166.735 ;
        RECT 47.630 166.715 47.980 167.365 ;
        RECT 45.330 166.155 45.605 166.500 ;
        RECT 45.775 166.395 47.440 166.565 ;
        RECT 48.150 166.545 48.380 167.535 ;
        RECT 45.795 165.825 46.175 166.225 ;
        RECT 46.345 166.045 46.515 166.395 ;
        RECT 46.685 165.825 47.015 166.225 ;
        RECT 47.185 166.045 47.440 166.395 ;
        RECT 47.715 166.375 48.380 166.545 ;
        RECT 47.715 166.085 47.885 166.375 ;
        RECT 48.055 165.825 48.385 166.205 ;
        RECT 48.555 166.085 48.740 168.205 ;
        RECT 48.980 167.915 49.245 168.375 ;
        RECT 49.415 167.780 49.665 168.205 ;
        RECT 49.875 167.930 50.980 168.100 ;
        RECT 49.360 167.650 49.665 167.780 ;
        RECT 48.910 166.455 49.190 167.405 ;
        RECT 49.360 166.545 49.530 167.650 ;
        RECT 49.700 166.865 49.940 167.460 ;
        RECT 50.110 167.395 50.640 167.760 ;
        RECT 50.110 166.695 50.280 167.395 ;
        RECT 50.810 167.315 50.980 167.930 ;
        RECT 51.150 167.575 51.320 168.375 ;
        RECT 51.490 167.875 51.740 168.205 ;
        RECT 51.965 167.905 52.850 168.075 ;
        RECT 50.810 167.225 51.320 167.315 ;
        RECT 49.360 166.415 49.585 166.545 ;
        RECT 49.755 166.475 50.280 166.695 ;
        RECT 50.450 167.055 51.320 167.225 ;
        RECT 48.995 165.825 49.245 166.285 ;
        RECT 49.415 166.275 49.585 166.415 ;
        RECT 50.450 166.275 50.620 167.055 ;
        RECT 51.150 166.985 51.320 167.055 ;
        RECT 50.830 166.805 51.030 166.835 ;
        RECT 51.490 166.805 51.660 167.875 ;
        RECT 51.830 166.985 52.020 167.705 ;
        RECT 50.830 166.505 51.660 166.805 ;
        RECT 52.190 166.775 52.510 167.735 ;
        RECT 49.415 166.105 49.750 166.275 ;
        RECT 49.945 166.105 50.620 166.275 ;
        RECT 50.940 165.825 51.310 166.325 ;
        RECT 51.490 166.275 51.660 166.505 ;
        RECT 52.045 166.445 52.510 166.775 ;
        RECT 52.680 167.065 52.850 167.905 ;
        RECT 53.030 167.875 53.345 168.375 ;
        RECT 53.575 167.645 53.915 168.205 ;
        RECT 53.020 167.270 53.915 167.645 ;
        RECT 54.085 167.365 54.255 168.375 ;
        RECT 53.725 167.065 53.915 167.270 ;
        RECT 54.425 167.315 54.755 168.160 ;
        RECT 54.985 167.505 55.260 168.205 ;
        RECT 55.430 167.830 55.685 168.375 ;
        RECT 55.855 167.865 56.335 168.205 ;
        RECT 56.510 167.820 57.115 168.375 ;
        RECT 56.500 167.720 57.115 167.820 ;
        RECT 56.500 167.695 56.685 167.720 ;
        RECT 54.425 167.235 54.815 167.315 ;
        RECT 54.600 167.185 54.815 167.235 ;
        RECT 52.680 166.735 53.555 167.065 ;
        RECT 53.725 166.735 54.475 167.065 ;
        RECT 52.680 166.275 52.850 166.735 ;
        RECT 53.725 166.565 53.925 166.735 ;
        RECT 54.645 166.605 54.815 167.185 ;
        RECT 54.590 166.565 54.815 166.605 ;
        RECT 51.490 166.105 51.895 166.275 ;
        RECT 52.065 166.105 52.850 166.275 ;
        RECT 53.125 165.825 53.335 166.355 ;
        RECT 53.595 166.040 53.925 166.565 ;
        RECT 54.435 166.480 54.815 166.565 ;
        RECT 54.095 165.825 54.265 166.435 ;
        RECT 54.435 166.045 54.765 166.480 ;
        RECT 54.985 166.475 55.155 167.505 ;
        RECT 55.430 167.375 56.185 167.625 ;
        RECT 56.355 167.450 56.685 167.695 ;
        RECT 55.430 167.340 56.200 167.375 ;
        RECT 55.430 167.330 56.215 167.340 ;
        RECT 55.325 167.315 56.220 167.330 ;
        RECT 55.325 167.300 56.240 167.315 ;
        RECT 55.325 167.290 56.260 167.300 ;
        RECT 55.325 167.280 56.285 167.290 ;
        RECT 55.325 167.250 56.355 167.280 ;
        RECT 55.325 167.220 56.375 167.250 ;
        RECT 55.325 167.190 56.395 167.220 ;
        RECT 55.325 167.165 56.425 167.190 ;
        RECT 55.325 167.130 56.460 167.165 ;
        RECT 55.325 167.125 56.490 167.130 ;
        RECT 55.325 166.730 55.555 167.125 ;
        RECT 56.100 167.120 56.490 167.125 ;
        RECT 56.125 167.110 56.490 167.120 ;
        RECT 56.140 167.105 56.490 167.110 ;
        RECT 56.155 167.100 56.490 167.105 ;
        RECT 56.855 167.100 57.115 167.550 ;
        RECT 56.155 167.095 57.115 167.100 ;
        RECT 56.165 167.085 57.115 167.095 ;
        RECT 56.175 167.080 57.115 167.085 ;
        RECT 56.185 167.070 57.115 167.080 ;
        RECT 56.190 167.060 57.115 167.070 ;
        RECT 56.195 167.055 57.115 167.060 ;
        RECT 56.205 167.040 57.115 167.055 ;
        RECT 56.210 167.025 57.115 167.040 ;
        RECT 56.220 167.000 57.115 167.025 ;
        RECT 55.725 166.530 56.055 166.955 ;
        RECT 54.985 165.995 55.245 166.475 ;
        RECT 55.415 165.825 55.665 166.365 ;
        RECT 55.835 166.045 56.055 166.530 ;
        RECT 56.225 166.930 57.115 167.000 ;
        RECT 57.285 167.235 57.670 168.205 ;
        RECT 57.840 167.915 58.165 168.375 ;
        RECT 58.685 167.745 58.965 168.205 ;
        RECT 57.840 167.525 58.965 167.745 ;
        RECT 56.225 166.205 56.395 166.930 ;
        RECT 56.565 166.375 57.115 166.760 ;
        RECT 57.285 166.565 57.565 167.235 ;
        RECT 57.840 167.065 58.290 167.525 ;
        RECT 59.155 167.355 59.555 168.205 ;
        RECT 59.955 167.915 60.225 168.375 ;
        RECT 60.395 167.745 60.680 168.205 ;
        RECT 57.735 166.735 58.290 167.065 ;
        RECT 58.460 166.795 59.555 167.355 ;
        RECT 57.840 166.625 58.290 166.735 ;
        RECT 56.225 166.035 57.115 166.205 ;
        RECT 57.285 165.995 57.670 166.565 ;
        RECT 57.840 166.455 58.965 166.625 ;
        RECT 57.840 165.825 58.165 166.285 ;
        RECT 58.685 165.995 58.965 166.455 ;
        RECT 59.155 165.995 59.555 166.795 ;
        RECT 59.725 167.525 60.680 167.745 ;
        RECT 59.725 166.625 59.935 167.525 ;
        RECT 60.105 166.795 60.795 167.355 ;
        RECT 61.425 167.210 61.715 168.375 ;
        RECT 62.435 167.705 62.605 168.205 ;
        RECT 62.775 167.875 63.105 168.375 ;
        RECT 62.435 167.535 63.100 167.705 ;
        RECT 62.350 166.715 62.700 167.365 ;
        RECT 59.725 166.455 60.680 166.625 ;
        RECT 59.955 165.825 60.225 166.285 ;
        RECT 60.395 165.995 60.680 166.455 ;
        RECT 61.425 165.825 61.715 166.550 ;
        RECT 62.870 166.545 63.100 167.535 ;
        RECT 62.435 166.375 63.100 166.545 ;
        RECT 62.435 166.085 62.605 166.375 ;
        RECT 62.775 165.825 63.105 166.205 ;
        RECT 63.275 166.085 63.460 168.205 ;
        RECT 63.700 167.915 63.965 168.375 ;
        RECT 64.135 167.780 64.385 168.205 ;
        RECT 64.595 167.930 65.700 168.100 ;
        RECT 64.080 167.650 64.385 167.780 ;
        RECT 63.630 166.455 63.910 167.405 ;
        RECT 64.080 166.545 64.250 167.650 ;
        RECT 64.420 166.865 64.660 167.460 ;
        RECT 64.830 167.395 65.360 167.760 ;
        RECT 64.830 166.695 65.000 167.395 ;
        RECT 65.530 167.315 65.700 167.930 ;
        RECT 65.870 167.575 66.040 168.375 ;
        RECT 66.210 167.875 66.460 168.205 ;
        RECT 66.685 167.905 67.570 168.075 ;
        RECT 65.530 167.225 66.040 167.315 ;
        RECT 64.080 166.415 64.305 166.545 ;
        RECT 64.475 166.475 65.000 166.695 ;
        RECT 65.170 167.055 66.040 167.225 ;
        RECT 63.715 165.825 63.965 166.285 ;
        RECT 64.135 166.275 64.305 166.415 ;
        RECT 65.170 166.275 65.340 167.055 ;
        RECT 65.870 166.985 66.040 167.055 ;
        RECT 65.550 166.805 65.750 166.835 ;
        RECT 66.210 166.805 66.380 167.875 ;
        RECT 66.550 166.985 66.740 167.705 ;
        RECT 65.550 166.505 66.380 166.805 ;
        RECT 66.910 166.775 67.230 167.735 ;
        RECT 64.135 166.105 64.470 166.275 ;
        RECT 64.665 166.105 65.340 166.275 ;
        RECT 65.660 165.825 66.030 166.325 ;
        RECT 66.210 166.275 66.380 166.505 ;
        RECT 66.765 166.445 67.230 166.775 ;
        RECT 67.400 167.065 67.570 167.905 ;
        RECT 67.750 167.875 68.065 168.375 ;
        RECT 68.295 167.645 68.635 168.205 ;
        RECT 67.740 167.270 68.635 167.645 ;
        RECT 68.805 167.365 68.975 168.375 ;
        RECT 68.445 167.065 68.635 167.270 ;
        RECT 69.145 167.315 69.475 168.160 ;
        RECT 69.145 167.235 69.535 167.315 ;
        RECT 69.320 167.185 69.535 167.235 ;
        RECT 67.400 166.735 68.275 167.065 ;
        RECT 68.445 166.735 69.195 167.065 ;
        RECT 67.400 166.275 67.570 166.735 ;
        RECT 68.445 166.565 68.645 166.735 ;
        RECT 69.365 166.605 69.535 167.185 ;
        RECT 69.310 166.565 69.535 166.605 ;
        RECT 66.210 166.105 66.615 166.275 ;
        RECT 66.785 166.105 67.570 166.275 ;
        RECT 67.845 165.825 68.055 166.355 ;
        RECT 68.315 166.040 68.645 166.565 ;
        RECT 69.155 166.480 69.535 166.565 ;
        RECT 70.625 167.235 71.010 168.205 ;
        RECT 71.180 167.915 71.505 168.375 ;
        RECT 72.025 167.745 72.305 168.205 ;
        RECT 71.180 167.525 72.305 167.745 ;
        RECT 70.625 166.565 70.905 167.235 ;
        RECT 71.180 167.065 71.630 167.525 ;
        RECT 72.495 167.355 72.895 168.205 ;
        RECT 73.295 167.915 73.565 168.375 ;
        RECT 73.735 167.745 74.020 168.205 ;
        RECT 71.075 166.735 71.630 167.065 ;
        RECT 71.800 166.795 72.895 167.355 ;
        RECT 71.180 166.625 71.630 166.735 ;
        RECT 68.815 165.825 68.985 166.435 ;
        RECT 69.155 166.045 69.485 166.480 ;
        RECT 70.625 165.995 71.010 166.565 ;
        RECT 71.180 166.455 72.305 166.625 ;
        RECT 71.180 165.825 71.505 166.285 ;
        RECT 72.025 165.995 72.305 166.455 ;
        RECT 72.495 165.995 72.895 166.795 ;
        RECT 73.065 167.525 74.020 167.745 ;
        RECT 73.065 166.625 73.275 167.525 ;
        RECT 73.445 166.795 74.135 167.355 ;
        RECT 74.310 167.235 74.645 168.205 ;
        RECT 74.815 167.235 74.985 168.375 ;
        RECT 75.155 168.035 77.185 168.205 ;
        RECT 73.065 166.455 74.020 166.625 ;
        RECT 73.295 165.825 73.565 166.285 ;
        RECT 73.735 165.995 74.020 166.455 ;
        RECT 74.310 166.565 74.480 167.235 ;
        RECT 75.155 167.065 75.325 168.035 ;
        RECT 74.650 166.735 74.905 167.065 ;
        RECT 75.130 166.735 75.325 167.065 ;
        RECT 75.495 167.695 76.620 167.865 ;
        RECT 74.735 166.565 74.905 166.735 ;
        RECT 75.495 166.565 75.665 167.695 ;
        RECT 74.310 165.995 74.565 166.565 ;
        RECT 74.735 166.395 75.665 166.565 ;
        RECT 75.835 167.355 76.845 167.525 ;
        RECT 75.835 166.555 76.005 167.355 ;
        RECT 75.490 166.360 75.665 166.395 ;
        RECT 74.735 165.825 75.065 166.225 ;
        RECT 75.490 165.995 76.020 166.360 ;
        RECT 76.210 166.335 76.485 167.155 ;
        RECT 76.205 166.165 76.485 166.335 ;
        RECT 76.210 165.995 76.485 166.165 ;
        RECT 76.655 165.995 76.845 167.355 ;
        RECT 77.015 167.370 77.185 168.035 ;
        RECT 77.355 167.615 77.525 168.375 ;
        RECT 77.760 167.615 78.275 168.025 ;
        RECT 77.015 167.180 77.765 167.370 ;
        RECT 77.935 166.805 78.275 167.615 ;
        RECT 78.445 167.285 79.655 168.375 ;
        RECT 79.825 167.865 81.025 168.105 ;
        RECT 81.205 167.950 81.535 168.375 ;
        RECT 82.050 167.950 82.410 168.375 ;
        RECT 82.615 167.780 82.875 167.960 ;
        RECT 81.240 167.695 82.875 167.780 ;
        RECT 77.045 166.635 78.275 166.805 ;
        RECT 77.025 165.825 77.535 166.360 ;
        RECT 77.755 166.030 78.000 166.635 ;
        RECT 78.445 166.575 78.965 167.115 ;
        RECT 79.135 166.745 79.655 167.285 ;
        RECT 79.825 167.235 80.130 167.665 ;
        RECT 80.300 167.610 82.875 167.695 ;
        RECT 80.300 167.525 81.410 167.610 ;
        RECT 82.195 167.550 82.875 167.610 ;
        RECT 78.445 165.825 79.655 166.575 ;
        RECT 79.825 166.565 79.995 167.235 ;
        RECT 80.300 167.065 80.470 167.525 ;
        RECT 80.170 166.735 80.470 167.065 ;
        RECT 80.730 166.815 81.265 167.355 ;
        RECT 81.630 167.235 82.025 167.440 ;
        RECT 81.515 166.675 81.685 167.065 ;
        RECT 81.365 166.645 81.685 166.675 ;
        RECT 80.800 166.565 81.685 166.645 ;
        RECT 79.825 166.505 81.685 166.565 ;
        RECT 79.825 166.475 81.535 166.505 ;
        RECT 79.825 166.395 80.970 166.475 ;
        RECT 79.825 166.345 80.130 166.395 ;
        RECT 79.875 166.045 80.130 166.345 ;
        RECT 80.300 165.825 80.630 166.225 ;
        RECT 80.800 166.045 80.970 166.395 ;
        RECT 81.855 166.335 82.025 167.235 ;
        RECT 82.195 166.645 82.365 167.550 ;
        RECT 82.535 166.815 82.875 167.380 ;
        RECT 83.045 167.285 84.715 168.375 ;
        RECT 85.085 167.705 85.365 168.375 ;
        RECT 85.535 167.485 85.835 168.035 ;
        RECT 86.035 167.655 86.365 168.375 ;
        RECT 86.555 167.655 87.015 168.205 ;
        RECT 82.195 166.475 82.875 166.645 ;
        RECT 81.270 165.825 81.440 166.305 ;
        RECT 81.675 166.005 82.025 166.335 ;
        RECT 82.195 165.825 82.365 166.305 ;
        RECT 82.615 166.030 82.875 166.475 ;
        RECT 83.045 166.595 83.795 167.115 ;
        RECT 83.965 166.765 84.715 167.285 ;
        RECT 84.900 167.065 85.165 167.425 ;
        RECT 85.535 167.315 86.475 167.485 ;
        RECT 86.305 167.065 86.475 167.315 ;
        RECT 84.900 166.815 85.575 167.065 ;
        RECT 85.795 166.815 86.135 167.065 ;
        RECT 86.305 166.735 86.595 167.065 ;
        RECT 86.305 166.645 86.475 166.735 ;
        RECT 83.045 165.825 84.715 166.595 ;
        RECT 85.085 166.455 86.475 166.645 ;
        RECT 85.085 166.095 85.415 166.455 ;
        RECT 86.765 166.285 87.015 167.655 ;
        RECT 87.185 167.210 87.475 168.375 ;
        RECT 87.650 167.405 87.925 168.205 ;
        RECT 88.095 167.575 88.425 168.375 ;
        RECT 88.595 168.035 89.735 168.205 ;
        RECT 88.595 167.405 88.765 168.035 ;
        RECT 87.650 167.195 88.765 167.405 ;
        RECT 88.935 167.405 89.265 167.865 ;
        RECT 89.435 167.575 89.735 168.035 ;
        RECT 90.015 167.405 90.375 167.580 ;
        RECT 90.960 167.575 91.130 168.375 ;
        RECT 91.300 167.745 91.630 168.205 ;
        RECT 91.800 167.915 91.970 168.375 ;
        RECT 91.300 167.575 92.075 167.745 ;
        RECT 88.935 167.185 89.695 167.405 ;
        RECT 90.015 167.235 91.475 167.405 ;
        RECT 87.650 166.815 88.370 167.015 ;
        RECT 88.540 166.815 89.310 167.015 ;
        RECT 89.480 166.645 89.695 167.185 ;
        RECT 90.010 166.675 90.205 167.065 ;
        RECT 86.035 165.825 86.285 166.285 ;
        RECT 86.455 165.995 87.015 166.285 ;
        RECT 87.185 165.825 87.475 166.550 ;
        RECT 87.650 165.825 87.925 166.645 ;
        RECT 88.095 166.475 89.695 166.645 ;
        RECT 90.005 166.505 90.205 166.675 ;
        RECT 88.095 166.465 89.265 166.475 ;
        RECT 88.095 165.995 88.425 166.465 ;
        RECT 88.595 165.825 88.765 166.295 ;
        RECT 88.935 165.995 89.265 166.465 ;
        RECT 90.375 166.335 90.555 167.235 ;
        RECT 90.725 166.505 91.135 167.065 ;
        RECT 91.305 166.735 91.475 167.235 ;
        RECT 91.645 166.565 92.075 167.575 ;
        RECT 92.245 167.285 95.755 168.375 ;
        RECT 96.015 167.705 96.185 168.205 ;
        RECT 96.355 167.875 96.685 168.375 ;
        RECT 96.015 167.535 96.680 167.705 ;
        RECT 91.380 166.395 92.075 166.565 ;
        RECT 92.245 166.595 93.895 167.115 ;
        RECT 94.065 166.765 95.755 167.285 ;
        RECT 95.930 166.715 96.280 167.365 ;
        RECT 89.435 165.825 89.725 166.295 ;
        RECT 89.965 165.825 90.205 166.335 ;
        RECT 90.375 165.995 90.665 166.335 ;
        RECT 90.895 165.825 91.210 166.335 ;
        RECT 91.380 166.125 91.550 166.395 ;
        RECT 91.720 165.825 92.050 166.225 ;
        RECT 92.245 165.825 95.755 166.595 ;
        RECT 96.450 166.545 96.680 167.535 ;
        RECT 96.015 166.375 96.680 166.545 ;
        RECT 96.015 166.085 96.185 166.375 ;
        RECT 96.355 165.825 96.685 166.205 ;
        RECT 96.855 166.085 97.040 168.205 ;
        RECT 97.280 167.915 97.545 168.375 ;
        RECT 97.715 167.780 97.965 168.205 ;
        RECT 98.175 167.930 99.280 168.100 ;
        RECT 97.660 167.650 97.965 167.780 ;
        RECT 97.210 166.455 97.490 167.405 ;
        RECT 97.660 166.545 97.830 167.650 ;
        RECT 98.000 166.865 98.240 167.460 ;
        RECT 98.410 167.395 98.940 167.760 ;
        RECT 98.410 166.695 98.580 167.395 ;
        RECT 99.110 167.315 99.280 167.930 ;
        RECT 99.450 167.575 99.620 168.375 ;
        RECT 99.790 167.875 100.040 168.205 ;
        RECT 100.265 167.905 101.150 168.075 ;
        RECT 99.110 167.225 99.620 167.315 ;
        RECT 97.660 166.415 97.885 166.545 ;
        RECT 98.055 166.475 98.580 166.695 ;
        RECT 98.750 167.055 99.620 167.225 ;
        RECT 97.295 165.825 97.545 166.285 ;
        RECT 97.715 166.275 97.885 166.415 ;
        RECT 98.750 166.275 98.920 167.055 ;
        RECT 99.450 166.985 99.620 167.055 ;
        RECT 99.130 166.805 99.330 166.835 ;
        RECT 99.790 166.805 99.960 167.875 ;
        RECT 100.130 166.985 100.320 167.705 ;
        RECT 99.130 166.505 99.960 166.805 ;
        RECT 100.490 166.775 100.810 167.735 ;
        RECT 97.715 166.105 98.050 166.275 ;
        RECT 98.245 166.105 98.920 166.275 ;
        RECT 99.240 165.825 99.610 166.325 ;
        RECT 99.790 166.275 99.960 166.505 ;
        RECT 100.345 166.445 100.810 166.775 ;
        RECT 100.980 167.065 101.150 167.905 ;
        RECT 101.330 167.875 101.645 168.375 ;
        RECT 101.875 167.645 102.215 168.205 ;
        RECT 101.320 167.270 102.215 167.645 ;
        RECT 102.385 167.365 102.555 168.375 ;
        RECT 102.025 167.065 102.215 167.270 ;
        RECT 102.725 167.315 103.055 168.160 ;
        RECT 103.390 167.915 103.560 168.375 ;
        RECT 103.730 167.745 104.060 168.205 ;
        RECT 103.285 167.575 104.060 167.745 ;
        RECT 104.230 167.575 104.400 168.375 ;
        RECT 102.725 167.235 103.115 167.315 ;
        RECT 102.900 167.185 103.115 167.235 ;
        RECT 100.980 166.735 101.855 167.065 ;
        RECT 102.025 166.735 102.775 167.065 ;
        RECT 100.980 166.275 101.150 166.735 ;
        RECT 102.025 166.565 102.225 166.735 ;
        RECT 102.945 166.605 103.115 167.185 ;
        RECT 102.890 166.565 103.115 166.605 ;
        RECT 99.790 166.105 100.195 166.275 ;
        RECT 100.365 166.105 101.150 166.275 ;
        RECT 101.425 165.825 101.635 166.355 ;
        RECT 101.895 166.040 102.225 166.565 ;
        RECT 102.735 166.480 103.115 166.565 ;
        RECT 103.285 166.565 103.715 167.575 ;
        RECT 104.985 167.405 105.345 167.580 ;
        RECT 103.885 167.235 105.345 167.405 ;
        RECT 105.655 167.405 106.015 167.580 ;
        RECT 106.600 167.575 106.770 168.375 ;
        RECT 106.940 167.745 107.270 168.205 ;
        RECT 107.440 167.915 107.610 168.375 ;
        RECT 106.940 167.575 107.715 167.745 ;
        RECT 105.655 167.235 107.115 167.405 ;
        RECT 103.885 166.735 104.055 167.235 ;
        RECT 102.395 165.825 102.565 166.435 ;
        RECT 102.735 166.045 103.065 166.480 ;
        RECT 103.285 166.395 103.980 166.565 ;
        RECT 104.225 166.505 104.635 167.065 ;
        RECT 103.310 165.825 103.640 166.225 ;
        RECT 103.810 166.125 103.980 166.395 ;
        RECT 104.805 166.335 104.985 167.235 ;
        RECT 105.155 166.675 105.350 167.065 ;
        RECT 105.650 167.015 105.845 167.065 ;
        RECT 105.645 166.845 105.845 167.015 ;
        RECT 105.155 166.505 105.355 166.675 ;
        RECT 105.650 166.505 105.845 166.845 ;
        RECT 106.015 166.335 106.195 167.235 ;
        RECT 106.365 166.505 106.775 167.065 ;
        RECT 106.945 166.735 107.115 167.235 ;
        RECT 107.285 166.565 107.715 167.575 ;
        RECT 107.890 167.405 108.165 168.205 ;
        RECT 108.335 167.575 108.665 168.375 ;
        RECT 108.835 168.035 109.975 168.205 ;
        RECT 108.835 167.405 109.005 168.035 ;
        RECT 107.890 167.195 109.005 167.405 ;
        RECT 109.175 167.405 109.505 167.865 ;
        RECT 109.675 167.575 109.975 168.035 ;
        RECT 109.175 167.355 109.935 167.405 ;
        RECT 109.175 167.185 109.955 167.355 ;
        RECT 110.185 167.285 112.775 168.375 ;
        RECT 107.890 166.815 108.610 167.015 ;
        RECT 108.780 166.815 109.550 167.015 ;
        RECT 109.720 166.645 109.935 167.185 ;
        RECT 107.020 166.395 107.715 166.565 ;
        RECT 104.150 165.825 104.465 166.335 ;
        RECT 104.695 165.995 104.985 166.335 ;
        RECT 105.155 165.825 105.395 166.335 ;
        RECT 105.605 165.825 105.845 166.335 ;
        RECT 106.015 165.995 106.305 166.335 ;
        RECT 106.535 165.825 106.850 166.335 ;
        RECT 107.020 166.125 107.190 166.395 ;
        RECT 107.360 165.825 107.690 166.225 ;
        RECT 107.890 165.825 108.165 166.645 ;
        RECT 108.335 166.475 109.935 166.645 ;
        RECT 110.185 166.595 111.395 167.115 ;
        RECT 111.565 166.765 112.775 167.285 ;
        RECT 112.945 167.210 113.235 168.375 ;
        RECT 113.405 167.285 116.915 168.375 ;
        RECT 113.405 166.595 115.055 167.115 ;
        RECT 115.225 166.765 116.915 167.285 ;
        RECT 118.010 167.235 118.345 168.205 ;
        RECT 118.515 167.235 118.685 168.375 ;
        RECT 118.855 168.035 120.885 168.205 ;
        RECT 108.335 166.465 109.505 166.475 ;
        RECT 108.335 165.995 108.665 166.465 ;
        RECT 108.835 165.825 109.005 166.295 ;
        RECT 109.175 165.995 109.505 166.465 ;
        RECT 109.675 165.825 109.965 166.295 ;
        RECT 110.185 165.825 112.775 166.595 ;
        RECT 112.945 165.825 113.235 166.550 ;
        RECT 113.405 165.825 116.915 166.595 ;
        RECT 118.010 166.565 118.180 167.235 ;
        RECT 118.855 167.065 119.025 168.035 ;
        RECT 118.350 166.735 118.605 167.065 ;
        RECT 118.830 166.735 119.025 167.065 ;
        RECT 119.195 167.695 120.320 167.865 ;
        RECT 118.435 166.565 118.605 166.735 ;
        RECT 119.195 166.565 119.365 167.695 ;
        RECT 118.010 165.995 118.265 166.565 ;
        RECT 118.435 166.395 119.365 166.565 ;
        RECT 119.535 167.355 120.545 167.525 ;
        RECT 119.535 166.555 119.705 167.355 ;
        RECT 119.910 166.675 120.185 167.155 ;
        RECT 119.905 166.505 120.185 166.675 ;
        RECT 119.190 166.360 119.365 166.395 ;
        RECT 118.435 165.825 118.765 166.225 ;
        RECT 119.190 165.995 119.720 166.360 ;
        RECT 119.910 165.995 120.185 166.505 ;
        RECT 120.355 165.995 120.545 167.355 ;
        RECT 120.715 167.370 120.885 168.035 ;
        RECT 121.055 167.615 121.225 168.375 ;
        RECT 121.460 167.615 121.975 168.025 ;
        RECT 122.145 167.940 127.490 168.375 ;
        RECT 120.715 167.180 121.465 167.370 ;
        RECT 121.635 166.805 121.975 167.615 ;
        RECT 120.745 166.635 121.975 166.805 ;
        RECT 120.725 165.825 121.235 166.360 ;
        RECT 121.455 166.030 121.700 166.635 ;
        RECT 123.730 166.370 124.070 167.200 ;
        RECT 125.550 166.690 125.900 167.940 ;
        RECT 127.665 167.285 131.175 168.375 ;
        RECT 127.665 166.595 129.315 167.115 ;
        RECT 129.485 166.765 131.175 167.285 ;
        RECT 131.805 167.235 132.065 168.375 ;
        RECT 132.235 167.225 132.565 168.205 ;
        RECT 132.735 167.235 133.015 168.375 ;
        RECT 133.205 167.485 133.465 168.195 ;
        RECT 133.635 167.665 133.965 168.375 ;
        RECT 134.135 167.485 134.365 168.195 ;
        RECT 133.205 167.245 134.365 167.485 ;
        RECT 134.545 167.465 134.815 168.195 ;
        RECT 134.995 167.645 135.335 168.375 ;
        RECT 134.545 167.245 135.315 167.465 ;
        RECT 131.825 166.815 132.160 167.065 ;
        RECT 132.330 166.625 132.500 167.225 ;
        RECT 132.670 166.795 133.005 167.065 ;
        RECT 133.195 166.735 133.495 167.065 ;
        RECT 133.675 166.755 134.200 167.065 ;
        RECT 134.380 166.755 134.845 167.065 ;
        RECT 122.145 165.825 127.490 166.370 ;
        RECT 127.665 165.825 131.175 166.595 ;
        RECT 131.805 165.995 132.500 166.625 ;
        RECT 132.705 165.825 133.015 166.625 ;
        RECT 133.205 165.825 133.495 166.555 ;
        RECT 133.675 166.115 133.905 166.755 ;
        RECT 135.025 166.575 135.315 167.245 ;
        RECT 134.085 166.375 135.315 166.575 ;
        RECT 134.085 166.005 134.395 166.375 ;
        RECT 134.575 165.825 135.245 166.195 ;
        RECT 135.505 166.005 135.765 168.195 ;
        RECT 136.035 167.445 136.205 168.205 ;
        RECT 136.385 167.615 136.715 168.375 ;
        RECT 136.035 167.275 136.700 167.445 ;
        RECT 136.885 167.300 137.155 168.205 ;
        RECT 136.530 167.130 136.700 167.275 ;
        RECT 135.965 166.725 136.295 167.095 ;
        RECT 136.530 166.800 136.815 167.130 ;
        RECT 136.530 166.545 136.700 166.800 ;
        RECT 136.035 166.375 136.700 166.545 ;
        RECT 136.985 166.500 137.155 167.300 ;
        RECT 137.325 167.285 138.535 168.375 ;
        RECT 136.035 165.995 136.205 166.375 ;
        RECT 136.385 165.825 136.715 166.205 ;
        RECT 136.895 165.995 137.155 166.500 ;
        RECT 137.325 166.575 137.845 167.115 ;
        RECT 138.015 166.745 138.535 167.285 ;
        RECT 138.705 167.210 138.995 168.375 ;
        RECT 139.255 167.445 139.425 168.205 ;
        RECT 139.605 167.615 139.935 168.375 ;
        RECT 139.255 167.275 139.920 167.445 ;
        RECT 140.105 167.300 140.375 168.205 ;
        RECT 140.545 167.940 145.890 168.375 ;
        RECT 139.750 167.130 139.920 167.275 ;
        RECT 139.185 166.725 139.515 167.095 ;
        RECT 139.750 166.800 140.035 167.130 ;
        RECT 137.325 165.825 138.535 166.575 ;
        RECT 138.705 165.825 138.995 166.550 ;
        RECT 139.750 166.545 139.920 166.800 ;
        RECT 139.255 166.375 139.920 166.545 ;
        RECT 140.205 166.500 140.375 167.300 ;
        RECT 139.255 165.995 139.425 166.375 ;
        RECT 139.605 165.825 139.935 166.205 ;
        RECT 140.115 165.995 140.375 166.500 ;
        RECT 142.130 166.370 142.470 167.200 ;
        RECT 143.950 166.690 144.300 167.940 ;
        RECT 146.065 167.285 147.275 168.375 ;
        RECT 147.535 167.705 147.705 168.205 ;
        RECT 147.875 167.875 148.205 168.375 ;
        RECT 147.535 167.535 148.200 167.705 ;
        RECT 146.065 166.575 146.585 167.115 ;
        RECT 146.755 166.745 147.275 167.285 ;
        RECT 147.450 166.715 147.800 167.365 ;
        RECT 140.545 165.825 145.890 166.370 ;
        RECT 146.065 165.825 147.275 166.575 ;
        RECT 147.970 166.545 148.200 167.535 ;
        RECT 147.535 166.375 148.200 166.545 ;
        RECT 147.535 166.085 147.705 166.375 ;
        RECT 147.875 165.825 148.205 166.205 ;
        RECT 148.375 166.085 148.560 168.205 ;
        RECT 148.800 167.915 149.065 168.375 ;
        RECT 149.235 167.780 149.485 168.205 ;
        RECT 149.695 167.930 150.800 168.100 ;
        RECT 149.180 167.650 149.485 167.780 ;
        RECT 148.730 166.455 149.010 167.405 ;
        RECT 149.180 166.545 149.350 167.650 ;
        RECT 149.520 166.865 149.760 167.460 ;
        RECT 149.930 167.395 150.460 167.760 ;
        RECT 149.930 166.695 150.100 167.395 ;
        RECT 150.630 167.315 150.800 167.930 ;
        RECT 150.970 167.575 151.140 168.375 ;
        RECT 151.310 167.875 151.560 168.205 ;
        RECT 151.785 167.905 152.670 168.075 ;
        RECT 150.630 167.225 151.140 167.315 ;
        RECT 149.180 166.415 149.405 166.545 ;
        RECT 149.575 166.475 150.100 166.695 ;
        RECT 150.270 167.055 151.140 167.225 ;
        RECT 148.815 165.825 149.065 166.285 ;
        RECT 149.235 166.275 149.405 166.415 ;
        RECT 150.270 166.275 150.440 167.055 ;
        RECT 150.970 166.985 151.140 167.055 ;
        RECT 150.650 166.805 150.850 166.835 ;
        RECT 151.310 166.805 151.480 167.875 ;
        RECT 151.650 166.985 151.840 167.705 ;
        RECT 150.650 166.505 151.480 166.805 ;
        RECT 152.010 166.775 152.330 167.735 ;
        RECT 149.235 166.105 149.570 166.275 ;
        RECT 149.765 166.105 150.440 166.275 ;
        RECT 150.760 165.825 151.130 166.325 ;
        RECT 151.310 166.275 151.480 166.505 ;
        RECT 151.865 166.445 152.330 166.775 ;
        RECT 152.500 167.065 152.670 167.905 ;
        RECT 152.850 167.875 153.165 168.375 ;
        RECT 153.395 167.645 153.735 168.205 ;
        RECT 152.840 167.270 153.735 167.645 ;
        RECT 153.905 167.365 154.075 168.375 ;
        RECT 153.545 167.065 153.735 167.270 ;
        RECT 154.245 167.315 154.575 168.160 ;
        RECT 154.245 167.235 154.635 167.315 ;
        RECT 154.420 167.185 154.635 167.235 ;
        RECT 152.500 166.735 153.375 167.065 ;
        RECT 153.545 166.735 154.295 167.065 ;
        RECT 152.500 166.275 152.670 166.735 ;
        RECT 153.545 166.565 153.745 166.735 ;
        RECT 154.465 166.605 154.635 167.185 ;
        RECT 155.725 167.285 156.935 168.375 ;
        RECT 155.725 166.745 156.245 167.285 ;
        RECT 154.410 166.565 154.635 166.605 ;
        RECT 156.415 166.575 156.935 167.115 ;
        RECT 151.310 166.105 151.715 166.275 ;
        RECT 151.885 166.105 152.670 166.275 ;
        RECT 152.945 165.825 153.155 166.355 ;
        RECT 153.415 166.040 153.745 166.565 ;
        RECT 154.255 166.480 154.635 166.565 ;
        RECT 153.915 165.825 154.085 166.435 ;
        RECT 154.255 166.045 154.585 166.480 ;
        RECT 155.725 165.825 156.935 166.575 ;
        RECT 22.700 165.655 157.020 165.825 ;
        RECT 22.785 164.905 23.995 165.655 ;
        RECT 22.785 164.365 23.305 164.905 ;
        RECT 24.165 164.885 27.675 165.655 ;
        RECT 27.880 164.915 28.495 165.485 ;
        RECT 28.665 165.145 28.880 165.655 ;
        RECT 29.110 165.145 29.390 165.475 ;
        RECT 29.570 165.145 29.810 165.655 ;
        RECT 23.475 164.195 23.995 164.735 ;
        RECT 24.165 164.365 25.815 164.885 ;
        RECT 25.985 164.195 27.675 164.715 ;
        RECT 22.785 163.105 23.995 164.195 ;
        RECT 24.165 163.105 27.675 164.195 ;
        RECT 27.880 163.895 28.195 164.915 ;
        RECT 28.365 164.245 28.535 164.745 ;
        RECT 28.785 164.415 29.050 164.975 ;
        RECT 29.220 164.245 29.390 165.145 ;
        RECT 29.560 164.415 29.915 164.975 ;
        RECT 30.145 164.885 33.655 165.655 ;
        RECT 33.825 164.905 35.035 165.655 ;
        RECT 30.145 164.365 31.795 164.885 ;
        RECT 28.365 164.075 29.790 164.245 ;
        RECT 31.965 164.195 33.655 164.715 ;
        RECT 33.825 164.365 34.345 164.905 ;
        RECT 35.245 164.835 35.475 165.655 ;
        RECT 35.645 164.855 35.975 165.485 ;
        RECT 34.515 164.195 35.035 164.735 ;
        RECT 35.225 164.415 35.555 164.665 ;
        RECT 35.725 164.255 35.975 164.855 ;
        RECT 36.145 164.835 36.355 165.655 ;
        RECT 36.585 165.110 41.930 165.655 ;
        RECT 38.170 164.280 38.510 165.110 ;
        RECT 42.105 164.885 43.775 165.655 ;
        RECT 27.880 163.275 28.415 163.895 ;
        RECT 28.585 163.105 28.915 163.905 ;
        RECT 29.400 163.900 29.790 164.075 ;
        RECT 30.145 163.105 33.655 164.195 ;
        RECT 33.825 163.105 35.035 164.195 ;
        RECT 35.245 163.105 35.475 164.245 ;
        RECT 35.645 163.275 35.975 164.255 ;
        RECT 36.145 163.105 36.355 164.245 ;
        RECT 39.990 163.540 40.340 164.790 ;
        RECT 42.105 164.365 42.855 164.885 ;
        RECT 44.405 164.855 44.715 165.655 ;
        RECT 44.920 164.855 45.615 165.485 ;
        RECT 45.935 164.855 46.265 165.655 ;
        RECT 46.435 165.005 46.605 165.485 ;
        RECT 46.775 165.175 47.105 165.655 ;
        RECT 47.275 165.005 47.445 165.485 ;
        RECT 47.695 165.175 47.935 165.655 ;
        RECT 48.115 165.005 48.285 165.485 ;
        RECT 43.025 164.195 43.775 164.715 ;
        RECT 44.415 164.415 44.750 164.685 ;
        RECT 44.920 164.255 45.090 164.855 ;
        RECT 46.435 164.835 47.445 165.005 ;
        RECT 47.650 164.835 48.285 165.005 ;
        RECT 48.545 164.930 48.835 165.655 ;
        RECT 49.155 164.855 49.485 165.655 ;
        RECT 49.655 165.005 49.825 165.485 ;
        RECT 49.995 165.175 50.325 165.655 ;
        RECT 50.495 165.005 50.665 165.485 ;
        RECT 50.915 165.175 51.155 165.655 ;
        RECT 51.335 165.005 51.505 165.485 ;
        RECT 49.655 164.835 50.665 165.005 ;
        RECT 50.870 164.835 51.505 165.005 ;
        RECT 51.765 164.915 52.150 165.485 ;
        RECT 52.320 165.195 52.645 165.655 ;
        RECT 53.165 165.025 53.445 165.485 ;
        RECT 45.260 164.415 45.595 164.665 ;
        RECT 46.435 164.295 46.930 164.835 ;
        RECT 47.650 164.665 47.820 164.835 ;
        RECT 47.320 164.495 47.820 164.665 ;
        RECT 36.585 163.105 41.930 163.540 ;
        RECT 42.105 163.105 43.775 164.195 ;
        RECT 44.405 163.105 44.685 164.245 ;
        RECT 44.855 163.275 45.185 164.255 ;
        RECT 45.355 163.105 45.615 164.245 ;
        RECT 45.935 163.105 46.265 164.255 ;
        RECT 46.435 164.125 47.445 164.295 ;
        RECT 46.435 163.275 46.605 164.125 ;
        RECT 46.775 163.105 47.105 163.905 ;
        RECT 47.275 163.275 47.445 164.125 ;
        RECT 47.650 164.255 47.820 164.495 ;
        RECT 47.990 164.425 48.370 164.665 ;
        RECT 49.655 164.295 50.150 164.835 ;
        RECT 50.870 164.665 51.040 164.835 ;
        RECT 50.540 164.495 51.040 164.665 ;
        RECT 47.650 164.085 48.365 164.255 ;
        RECT 47.625 163.105 47.865 163.905 ;
        RECT 48.035 163.275 48.365 164.085 ;
        RECT 48.545 163.105 48.835 164.270 ;
        RECT 49.155 163.105 49.485 164.255 ;
        RECT 49.655 164.125 50.665 164.295 ;
        RECT 49.655 163.275 49.825 164.125 ;
        RECT 49.995 163.105 50.325 163.905 ;
        RECT 50.495 163.275 50.665 164.125 ;
        RECT 50.870 164.255 51.040 164.495 ;
        RECT 51.210 164.425 51.590 164.665 ;
        RECT 50.870 164.085 51.585 164.255 ;
        RECT 50.845 163.105 51.085 163.905 ;
        RECT 51.255 163.275 51.585 164.085 ;
        RECT 51.765 164.245 52.045 164.915 ;
        RECT 52.320 164.855 53.445 165.025 ;
        RECT 52.320 164.745 52.770 164.855 ;
        RECT 52.215 164.415 52.770 164.745 ;
        RECT 53.635 164.685 54.035 165.485 ;
        RECT 54.435 165.195 54.705 165.655 ;
        RECT 54.875 165.025 55.160 165.485 ;
        RECT 51.765 163.275 52.150 164.245 ;
        RECT 52.320 163.955 52.770 164.415 ;
        RECT 52.940 164.125 54.035 164.685 ;
        RECT 52.320 163.735 53.445 163.955 ;
        RECT 52.320 163.105 52.645 163.565 ;
        RECT 53.165 163.275 53.445 163.735 ;
        RECT 53.635 163.275 54.035 164.125 ;
        RECT 54.205 164.855 55.160 165.025 ;
        RECT 55.445 164.885 57.115 165.655 ;
        RECT 57.335 165.000 57.665 165.435 ;
        RECT 57.835 165.045 58.005 165.655 ;
        RECT 57.285 164.915 57.665 165.000 ;
        RECT 58.175 164.915 58.505 165.440 ;
        RECT 58.765 165.125 58.975 165.655 ;
        RECT 59.250 165.205 60.035 165.375 ;
        RECT 60.205 165.205 60.610 165.375 ;
        RECT 54.205 163.955 54.415 164.855 ;
        RECT 54.585 164.125 55.275 164.685 ;
        RECT 55.445 164.365 56.195 164.885 ;
        RECT 57.285 164.875 57.510 164.915 ;
        RECT 56.365 164.195 57.115 164.715 ;
        RECT 54.205 163.735 55.160 163.955 ;
        RECT 54.435 163.105 54.705 163.565 ;
        RECT 54.875 163.275 55.160 163.735 ;
        RECT 55.445 163.105 57.115 164.195 ;
        RECT 57.285 164.295 57.455 164.875 ;
        RECT 58.175 164.745 58.375 164.915 ;
        RECT 59.250 164.745 59.420 165.205 ;
        RECT 57.625 164.415 58.375 164.745 ;
        RECT 58.545 164.415 59.420 164.745 ;
        RECT 57.285 164.245 57.500 164.295 ;
        RECT 57.285 164.165 57.675 164.245 ;
        RECT 57.345 163.320 57.675 164.165 ;
        RECT 58.185 164.210 58.375 164.415 ;
        RECT 57.845 163.105 58.015 164.115 ;
        RECT 58.185 163.835 59.080 164.210 ;
        RECT 58.185 163.275 58.525 163.835 ;
        RECT 58.755 163.105 59.070 163.605 ;
        RECT 59.250 163.575 59.420 164.415 ;
        RECT 59.590 164.705 60.055 165.035 ;
        RECT 60.440 164.975 60.610 165.205 ;
        RECT 60.790 165.155 61.160 165.655 ;
        RECT 61.480 165.205 62.155 165.375 ;
        RECT 62.350 165.205 62.685 165.375 ;
        RECT 59.590 163.745 59.910 164.705 ;
        RECT 60.440 164.675 61.270 164.975 ;
        RECT 60.080 163.775 60.270 164.495 ;
        RECT 60.440 163.605 60.610 164.675 ;
        RECT 61.070 164.645 61.270 164.675 ;
        RECT 60.780 164.425 60.950 164.495 ;
        RECT 61.480 164.425 61.650 165.205 ;
        RECT 62.515 165.065 62.685 165.205 ;
        RECT 62.855 165.195 63.105 165.655 ;
        RECT 60.780 164.255 61.650 164.425 ;
        RECT 61.820 164.785 62.345 165.005 ;
        RECT 62.515 164.935 62.740 165.065 ;
        RECT 60.780 164.165 61.290 164.255 ;
        RECT 59.250 163.405 60.135 163.575 ;
        RECT 60.360 163.275 60.610 163.605 ;
        RECT 60.780 163.105 60.950 163.905 ;
        RECT 61.120 163.550 61.290 164.165 ;
        RECT 61.820 164.085 61.990 164.785 ;
        RECT 61.460 163.720 61.990 164.085 ;
        RECT 62.160 164.020 62.400 164.615 ;
        RECT 62.570 163.830 62.740 164.935 ;
        RECT 62.910 164.075 63.190 165.025 ;
        RECT 62.435 163.700 62.740 163.830 ;
        RECT 61.120 163.380 62.225 163.550 ;
        RECT 62.435 163.275 62.685 163.700 ;
        RECT 62.855 163.105 63.120 163.565 ;
        RECT 63.360 163.275 63.545 165.395 ;
        RECT 63.715 165.275 64.045 165.655 ;
        RECT 64.215 165.105 64.385 165.395 ;
        RECT 63.720 164.935 64.385 165.105 ;
        RECT 63.720 163.945 63.950 164.935 ;
        RECT 64.120 164.115 64.470 164.765 ;
        RECT 63.720 163.775 64.385 163.945 ;
        RECT 63.715 163.105 64.045 163.605 ;
        RECT 64.215 163.275 64.385 163.775 ;
        RECT 65.115 163.285 65.375 165.475 ;
        RECT 65.635 165.285 66.305 165.655 ;
        RECT 66.485 165.105 66.795 165.475 ;
        RECT 65.565 164.905 66.795 165.105 ;
        RECT 65.565 164.235 65.855 164.905 ;
        RECT 66.975 164.725 67.205 165.365 ;
        RECT 67.385 164.925 67.675 165.655 ;
        RECT 68.785 165.005 69.045 165.485 ;
        RECT 69.215 165.115 69.465 165.655 ;
        RECT 66.035 164.415 66.500 164.725 ;
        RECT 66.680 164.415 67.205 164.725 ;
        RECT 67.385 164.415 67.685 164.745 ;
        RECT 65.565 164.015 66.335 164.235 ;
        RECT 65.545 163.105 65.885 163.835 ;
        RECT 66.065 163.285 66.335 164.015 ;
        RECT 66.515 163.995 67.675 164.235 ;
        RECT 66.515 163.285 66.745 163.995 ;
        RECT 66.915 163.105 67.245 163.815 ;
        RECT 67.415 163.285 67.675 163.995 ;
        RECT 68.785 163.975 68.955 165.005 ;
        RECT 69.635 164.950 69.855 165.435 ;
        RECT 69.125 164.355 69.355 164.750 ;
        RECT 69.525 164.525 69.855 164.950 ;
        RECT 70.025 165.275 70.915 165.445 ;
        RECT 70.025 164.550 70.195 165.275 ;
        RECT 70.365 164.720 70.915 165.105 ;
        RECT 71.285 165.025 71.615 165.385 ;
        RECT 72.235 165.195 72.485 165.655 ;
        RECT 72.655 165.195 73.215 165.485 ;
        RECT 71.285 164.835 72.675 165.025 ;
        RECT 72.505 164.745 72.675 164.835 ;
        RECT 70.025 164.480 70.915 164.550 ;
        RECT 70.020 164.455 70.915 164.480 ;
        RECT 70.010 164.440 70.915 164.455 ;
        RECT 70.005 164.425 70.915 164.440 ;
        RECT 69.995 164.420 70.915 164.425 ;
        RECT 69.990 164.410 70.915 164.420 ;
        RECT 69.985 164.400 70.915 164.410 ;
        RECT 69.975 164.395 70.915 164.400 ;
        RECT 69.965 164.385 70.915 164.395 ;
        RECT 69.955 164.380 70.915 164.385 ;
        RECT 69.955 164.375 70.290 164.380 ;
        RECT 69.940 164.370 70.290 164.375 ;
        RECT 69.925 164.360 70.290 164.370 ;
        RECT 69.900 164.355 70.290 164.360 ;
        RECT 69.125 164.350 70.290 164.355 ;
        RECT 69.125 164.315 70.260 164.350 ;
        RECT 69.125 164.290 70.225 164.315 ;
        RECT 69.125 164.260 70.195 164.290 ;
        RECT 69.125 164.230 70.175 164.260 ;
        RECT 69.125 164.200 70.155 164.230 ;
        RECT 69.125 164.190 70.085 164.200 ;
        RECT 69.125 164.180 70.060 164.190 ;
        RECT 69.125 164.165 70.040 164.180 ;
        RECT 69.125 164.150 70.020 164.165 ;
        RECT 69.230 164.140 70.015 164.150 ;
        RECT 69.230 164.105 70.000 164.140 ;
        RECT 68.785 163.275 69.060 163.975 ;
        RECT 69.230 163.855 69.985 164.105 ;
        RECT 70.155 163.785 70.485 164.030 ;
        RECT 70.655 163.930 70.915 164.380 ;
        RECT 71.100 164.415 71.775 164.665 ;
        RECT 71.995 164.415 72.335 164.665 ;
        RECT 72.505 164.415 72.795 164.745 ;
        RECT 71.100 164.055 71.365 164.415 ;
        RECT 72.505 164.165 72.675 164.415 ;
        RECT 71.735 163.995 72.675 164.165 ;
        RECT 70.300 163.760 70.485 163.785 ;
        RECT 70.300 163.660 70.915 163.760 ;
        RECT 69.230 163.105 69.485 163.650 ;
        RECT 69.655 163.275 70.135 163.615 ;
        RECT 70.310 163.105 70.915 163.660 ;
        RECT 71.285 163.105 71.565 163.775 ;
        RECT 71.735 163.445 72.035 163.995 ;
        RECT 72.965 163.825 73.215 165.195 ;
        RECT 74.305 164.930 74.595 165.655 ;
        RECT 74.855 165.105 75.025 165.485 ;
        RECT 75.205 165.275 75.535 165.655 ;
        RECT 74.855 164.935 75.520 165.105 ;
        RECT 75.715 164.980 75.975 165.485 ;
        RECT 74.785 164.385 75.115 164.755 ;
        RECT 75.350 164.680 75.520 164.935 ;
        RECT 75.350 164.350 75.635 164.680 ;
        RECT 72.235 163.105 72.565 163.825 ;
        RECT 72.755 163.275 73.215 163.825 ;
        RECT 74.305 163.105 74.595 164.270 ;
        RECT 75.350 164.205 75.520 164.350 ;
        RECT 74.855 164.035 75.520 164.205 ;
        RECT 75.805 164.180 75.975 164.980 ;
        RECT 76.145 164.885 77.815 165.655 ;
        RECT 78.445 165.025 78.785 165.485 ;
        RECT 78.955 165.195 79.205 165.655 ;
        RECT 79.395 165.275 83.085 165.485 ;
        RECT 83.275 165.195 83.525 165.655 ;
        RECT 76.145 164.365 76.895 164.885 ;
        RECT 78.445 164.835 79.645 165.025 ;
        RECT 79.815 164.835 81.325 165.105 ;
        RECT 81.495 165.025 83.085 165.105 ;
        RECT 83.695 165.025 84.025 165.485 ;
        RECT 84.195 165.195 84.365 165.655 ;
        RECT 84.535 165.025 84.865 165.485 ;
        RECT 81.495 164.835 84.865 165.025 ;
        RECT 85.035 164.835 85.365 165.655 ;
        RECT 77.065 164.195 77.815 164.715 ;
        RECT 74.855 163.275 75.025 164.035 ;
        RECT 75.205 163.105 75.535 163.865 ;
        RECT 75.705 163.275 75.975 164.180 ;
        RECT 76.145 163.105 77.815 164.195 ;
        RECT 78.445 164.295 78.620 164.835 ;
        RECT 79.365 164.665 79.645 164.835 ;
        RECT 81.155 164.665 81.325 164.835 ;
        RECT 86.345 164.815 86.600 165.655 ;
        RECT 86.770 164.980 87.000 165.325 ;
        RECT 87.190 165.255 87.570 165.655 ;
        RECT 87.740 165.085 87.910 165.435 ;
        RECT 88.080 165.175 88.810 165.655 ;
        RECT 78.790 164.465 79.140 164.665 ;
        RECT 79.365 164.465 80.985 164.665 ;
        RECT 81.155 164.295 81.460 164.665 ;
        RECT 81.630 164.465 82.840 164.665 ;
        RECT 83.150 164.635 84.860 164.665 ;
        RECT 83.105 164.465 84.860 164.635 ;
        RECT 78.445 163.275 78.785 164.295 ;
        RECT 78.955 163.105 79.645 164.295 ;
        RECT 79.815 164.075 84.865 164.295 ;
        RECT 79.815 163.275 80.145 164.075 ;
        RECT 80.315 163.105 80.485 163.905 ;
        RECT 80.655 163.735 81.825 164.075 ;
        RECT 80.655 163.275 80.985 163.735 ;
        RECT 81.155 163.105 81.325 163.565 ;
        RECT 81.495 163.275 81.825 163.735 ;
        RECT 81.995 163.105 82.165 163.905 ;
        RECT 82.335 163.275 82.665 164.075 ;
        RECT 82.835 163.105 83.525 163.905 ;
        RECT 83.695 163.275 84.025 164.075 ;
        RECT 84.195 163.105 84.365 163.905 ;
        RECT 84.535 163.275 84.865 164.075 ;
        RECT 85.035 163.105 85.365 164.295 ;
        RECT 86.345 163.105 86.600 164.280 ;
        RECT 86.770 164.245 86.940 164.980 ;
        RECT 87.170 164.915 87.910 165.085 ;
        RECT 88.980 165.005 89.295 165.475 ;
        RECT 89.545 165.195 89.790 165.655 ;
        RECT 87.170 164.745 87.340 164.915 ;
        RECT 88.560 164.835 89.295 165.005 ;
        RECT 88.560 164.745 88.805 164.835 ;
        RECT 87.110 164.415 87.340 164.745 ;
        RECT 88.070 164.415 88.805 164.745 ;
        RECT 88.975 164.415 89.315 164.665 ;
        RECT 89.485 164.415 89.800 165.025 ;
        RECT 89.970 164.665 90.220 165.475 ;
        RECT 90.390 165.130 90.650 165.655 ;
        RECT 90.820 165.005 91.080 165.460 ;
        RECT 91.250 165.175 91.510 165.655 ;
        RECT 91.680 165.005 91.940 165.460 ;
        RECT 92.110 165.175 92.370 165.655 ;
        RECT 92.540 165.005 92.800 165.460 ;
        RECT 92.970 165.175 93.230 165.655 ;
        RECT 93.400 165.005 93.660 165.460 ;
        RECT 93.830 165.175 94.130 165.655 ;
        RECT 90.820 164.835 94.130 165.005 ;
        RECT 89.970 164.415 92.990 164.665 ;
        RECT 87.170 164.245 87.340 164.415 ;
        RECT 86.770 163.275 87.000 164.245 ;
        RECT 87.170 164.075 88.415 164.245 ;
        RECT 87.210 163.105 87.490 163.905 ;
        RECT 87.995 163.825 88.415 164.075 ;
        RECT 88.635 163.855 88.805 164.415 ;
        RECT 87.670 163.325 88.860 163.655 ;
        RECT 89.055 163.105 89.315 164.245 ;
        RECT 89.495 163.105 89.790 164.215 ;
        RECT 89.970 163.280 90.220 164.415 ;
        RECT 93.160 164.245 94.130 164.835 ;
        RECT 90.390 163.105 90.650 164.215 ;
        RECT 90.820 164.005 94.130 164.245 ;
        RECT 94.570 164.900 94.805 165.230 ;
        RECT 94.975 164.915 95.305 165.655 ;
        RECT 95.540 165.275 96.735 165.485 ;
        RECT 94.570 164.245 94.740 164.900 ;
        RECT 95.540 164.835 95.815 165.275 ;
        RECT 95.985 164.935 96.315 165.105 ;
        RECT 95.990 164.835 96.315 164.935 ;
        RECT 96.485 165.045 96.735 165.275 ;
        RECT 96.905 165.215 97.075 165.655 ;
        RECT 97.245 165.045 97.595 165.485 ;
        RECT 97.930 165.145 98.170 165.655 ;
        RECT 98.350 165.145 98.630 165.475 ;
        RECT 98.860 165.145 99.075 165.655 ;
        RECT 96.485 164.835 97.595 165.045 ;
        RECT 94.915 164.415 95.260 164.745 ;
        RECT 95.490 164.245 95.820 164.665 ;
        RECT 94.570 164.075 95.820 164.245 ;
        RECT 90.820 163.280 91.080 164.005 ;
        RECT 91.250 163.105 91.510 163.835 ;
        RECT 91.680 163.280 91.940 164.005 ;
        RECT 92.110 163.105 92.370 163.835 ;
        RECT 92.540 163.280 92.800 164.005 ;
        RECT 92.970 163.105 93.230 163.835 ;
        RECT 93.400 163.280 93.660 164.005 ;
        RECT 94.570 163.880 94.870 164.075 ;
        RECT 95.990 163.905 96.270 164.835 ;
        RECT 96.450 164.465 97.595 164.665 ;
        RECT 96.450 164.295 96.640 164.465 ;
        RECT 97.825 164.415 98.180 164.975 ;
        RECT 96.445 164.125 96.640 164.295 ;
        RECT 98.350 164.245 98.520 165.145 ;
        RECT 98.690 164.415 98.955 164.975 ;
        RECT 99.245 164.915 99.860 165.485 ;
        RECT 100.065 164.930 100.355 165.655 ;
        RECT 100.615 165.105 100.785 165.485 ;
        RECT 101.000 165.275 101.330 165.655 ;
        RECT 100.615 164.935 101.330 165.105 ;
        RECT 99.205 164.245 99.375 164.745 ;
        RECT 96.450 164.085 96.640 164.125 ;
        RECT 96.820 163.905 97.095 164.245 ;
        RECT 93.830 163.105 94.125 163.835 ;
        RECT 95.040 163.105 95.295 163.905 ;
        RECT 95.495 163.735 97.095 163.905 ;
        RECT 95.495 163.275 95.825 163.735 ;
        RECT 95.995 163.105 96.570 163.565 ;
        RECT 96.740 163.275 97.095 163.735 ;
        RECT 97.265 163.105 97.595 164.245 ;
        RECT 97.950 164.075 99.375 164.245 ;
        RECT 97.950 163.900 98.340 164.075 ;
        RECT 98.825 163.105 99.155 163.905 ;
        RECT 99.545 163.895 99.860 164.915 ;
        RECT 100.525 164.385 100.880 164.755 ;
        RECT 101.160 164.745 101.330 164.935 ;
        RECT 101.500 164.910 101.755 165.485 ;
        RECT 101.160 164.415 101.415 164.745 ;
        RECT 99.325 163.275 99.860 163.895 ;
        RECT 100.065 163.105 100.355 164.270 ;
        RECT 101.160 164.205 101.330 164.415 ;
        RECT 100.615 164.035 101.330 164.205 ;
        RECT 101.585 164.180 101.755 164.910 ;
        RECT 101.930 164.815 102.190 165.655 ;
        RECT 102.365 164.885 104.955 165.655 ;
        RECT 105.675 165.105 105.845 165.485 ;
        RECT 106.060 165.275 106.390 165.655 ;
        RECT 105.675 164.935 106.390 165.105 ;
        RECT 102.365 164.365 103.575 164.885 ;
        RECT 100.615 163.275 100.785 164.035 ;
        RECT 101.000 163.105 101.330 163.865 ;
        RECT 101.500 163.275 101.755 164.180 ;
        RECT 101.930 163.105 102.190 164.255 ;
        RECT 103.745 164.195 104.955 164.715 ;
        RECT 105.585 164.385 105.940 164.755 ;
        RECT 106.220 164.745 106.390 164.935 ;
        RECT 106.560 164.910 106.815 165.485 ;
        RECT 106.220 164.415 106.475 164.745 ;
        RECT 106.220 164.205 106.390 164.415 ;
        RECT 102.365 163.105 104.955 164.195 ;
        RECT 105.675 164.035 106.390 164.205 ;
        RECT 106.645 164.180 106.815 164.910 ;
        RECT 106.990 164.815 107.250 165.655 ;
        RECT 108.405 164.835 108.615 165.655 ;
        RECT 108.785 164.855 109.115 165.485 ;
        RECT 108.785 164.255 109.035 164.855 ;
        RECT 109.285 164.835 109.515 165.655 ;
        RECT 109.725 164.885 113.235 165.655 ;
        RECT 113.955 165.105 114.125 165.395 ;
        RECT 114.295 165.275 114.625 165.655 ;
        RECT 113.955 164.935 114.620 165.105 ;
        RECT 109.205 164.415 109.535 164.665 ;
        RECT 109.725 164.365 111.375 164.885 ;
        RECT 105.675 163.275 105.845 164.035 ;
        RECT 106.060 163.105 106.390 163.865 ;
        RECT 106.560 163.275 106.815 164.180 ;
        RECT 106.990 163.105 107.250 164.255 ;
        RECT 108.405 163.105 108.615 164.245 ;
        RECT 108.785 163.275 109.115 164.255 ;
        RECT 109.285 163.105 109.515 164.245 ;
        RECT 111.545 164.195 113.235 164.715 ;
        RECT 109.725 163.105 113.235 164.195 ;
        RECT 113.870 164.115 114.220 164.765 ;
        RECT 114.390 163.945 114.620 164.935 ;
        RECT 113.955 163.775 114.620 163.945 ;
        RECT 113.955 163.275 114.125 163.775 ;
        RECT 114.295 163.105 114.625 163.605 ;
        RECT 114.795 163.275 114.980 165.395 ;
        RECT 115.235 165.195 115.485 165.655 ;
        RECT 115.655 165.205 115.990 165.375 ;
        RECT 116.185 165.205 116.860 165.375 ;
        RECT 115.655 165.065 115.825 165.205 ;
        RECT 115.150 164.075 115.430 165.025 ;
        RECT 115.600 164.935 115.825 165.065 ;
        RECT 115.600 163.830 115.770 164.935 ;
        RECT 115.995 164.785 116.520 165.005 ;
        RECT 115.940 164.020 116.180 164.615 ;
        RECT 116.350 164.085 116.520 164.785 ;
        RECT 116.690 164.425 116.860 165.205 ;
        RECT 117.180 165.155 117.550 165.655 ;
        RECT 117.730 165.205 118.135 165.375 ;
        RECT 118.305 165.205 119.090 165.375 ;
        RECT 117.730 164.975 117.900 165.205 ;
        RECT 117.070 164.675 117.900 164.975 ;
        RECT 118.285 164.705 118.750 165.035 ;
        RECT 117.070 164.645 117.270 164.675 ;
        RECT 117.390 164.425 117.560 164.495 ;
        RECT 116.690 164.255 117.560 164.425 ;
        RECT 117.050 164.165 117.560 164.255 ;
        RECT 115.600 163.700 115.905 163.830 ;
        RECT 116.350 163.720 116.880 164.085 ;
        RECT 115.220 163.105 115.485 163.565 ;
        RECT 115.655 163.275 115.905 163.700 ;
        RECT 117.050 163.550 117.220 164.165 ;
        RECT 116.115 163.380 117.220 163.550 ;
        RECT 117.390 163.105 117.560 163.905 ;
        RECT 117.730 163.605 117.900 164.675 ;
        RECT 118.070 163.775 118.260 164.495 ;
        RECT 118.430 163.745 118.750 164.705 ;
        RECT 118.920 164.745 119.090 165.205 ;
        RECT 119.365 165.125 119.575 165.655 ;
        RECT 119.835 164.915 120.165 165.440 ;
        RECT 120.335 165.045 120.505 165.655 ;
        RECT 120.675 165.000 121.005 165.435 ;
        RECT 121.340 165.025 121.625 165.485 ;
        RECT 121.795 165.195 122.065 165.655 ;
        RECT 120.675 164.915 121.055 165.000 ;
        RECT 119.965 164.745 120.165 164.915 ;
        RECT 120.830 164.875 121.055 164.915 ;
        RECT 118.920 164.415 119.795 164.745 ;
        RECT 119.965 164.415 120.715 164.745 ;
        RECT 117.730 163.275 117.980 163.605 ;
        RECT 118.920 163.575 119.090 164.415 ;
        RECT 119.965 164.210 120.155 164.415 ;
        RECT 120.885 164.295 121.055 164.875 ;
        RECT 121.340 164.855 122.295 165.025 ;
        RECT 120.840 164.245 121.055 164.295 ;
        RECT 119.260 163.835 120.155 164.210 ;
        RECT 120.665 164.165 121.055 164.245 ;
        RECT 118.205 163.405 119.090 163.575 ;
        RECT 119.270 163.105 119.585 163.605 ;
        RECT 119.815 163.275 120.155 163.835 ;
        RECT 120.325 163.105 120.495 164.115 ;
        RECT 120.665 163.320 120.995 164.165 ;
        RECT 121.225 164.125 121.915 164.685 ;
        RECT 122.085 163.955 122.295 164.855 ;
        RECT 121.340 163.735 122.295 163.955 ;
        RECT 122.465 164.685 122.865 165.485 ;
        RECT 123.055 165.025 123.335 165.485 ;
        RECT 123.855 165.195 124.180 165.655 ;
        RECT 123.055 164.855 124.180 165.025 ;
        RECT 124.350 164.915 124.735 165.485 ;
        RECT 125.825 164.930 126.115 165.655 ;
        RECT 123.730 164.745 124.180 164.855 ;
        RECT 122.465 164.125 123.560 164.685 ;
        RECT 123.730 164.415 124.285 164.745 ;
        RECT 121.340 163.275 121.625 163.735 ;
        RECT 121.795 163.105 122.065 163.565 ;
        RECT 122.465 163.275 122.865 164.125 ;
        RECT 123.730 163.955 124.180 164.415 ;
        RECT 124.455 164.245 124.735 164.915 ;
        RECT 126.285 164.885 128.875 165.655 ;
        RECT 129.050 165.165 129.305 165.655 ;
        RECT 129.475 165.145 130.705 165.485 ;
        RECT 130.970 165.155 131.465 165.485 ;
        RECT 126.285 164.365 127.495 164.885 ;
        RECT 123.055 163.735 124.180 163.955 ;
        RECT 123.055 163.275 123.335 163.735 ;
        RECT 123.855 163.105 124.180 163.565 ;
        RECT 124.350 163.275 124.735 164.245 ;
        RECT 125.825 163.105 126.115 164.270 ;
        RECT 127.665 164.195 128.875 164.715 ;
        RECT 129.070 164.415 129.290 164.995 ;
        RECT 129.475 164.245 129.655 165.145 ;
        RECT 129.825 164.415 130.200 164.975 ;
        RECT 130.375 164.915 130.705 165.145 ;
        RECT 130.405 164.415 130.715 164.745 ;
        RECT 126.285 163.105 128.875 164.195 ;
        RECT 129.050 163.105 129.305 164.245 ;
        RECT 129.475 164.075 130.705 164.245 ;
        RECT 129.475 163.275 129.805 164.075 ;
        RECT 129.975 163.105 130.205 163.905 ;
        RECT 130.375 163.275 130.705 164.075 ;
        RECT 130.885 163.665 131.125 164.975 ;
        RECT 131.295 164.245 131.465 165.155 ;
        RECT 131.685 164.415 132.035 165.380 ;
        RECT 132.215 164.415 132.515 165.385 ;
        RECT 132.695 164.415 132.975 165.385 ;
        RECT 133.155 164.855 133.425 165.655 ;
        RECT 133.595 164.935 133.935 165.445 ;
        RECT 134.105 165.275 134.995 165.445 ;
        RECT 133.170 164.415 133.500 164.665 ;
        RECT 133.170 164.245 133.485 164.415 ;
        RECT 131.295 164.075 133.485 164.245 ;
        RECT 130.890 163.105 131.225 163.485 ;
        RECT 131.395 163.275 131.645 164.075 ;
        RECT 131.865 163.105 132.195 163.825 ;
        RECT 132.380 163.275 132.630 164.075 ;
        RECT 133.095 163.105 133.425 163.905 ;
        RECT 133.675 163.535 133.935 164.935 ;
        RECT 134.105 164.720 134.655 165.105 ;
        RECT 134.825 164.550 134.995 165.275 ;
        RECT 134.105 164.480 134.995 164.550 ;
        RECT 135.165 164.950 135.385 165.435 ;
        RECT 135.555 165.115 135.805 165.655 ;
        RECT 135.975 165.005 136.235 165.485 ;
        RECT 135.165 164.525 135.495 164.950 ;
        RECT 134.105 164.455 135.000 164.480 ;
        RECT 134.105 164.440 135.010 164.455 ;
        RECT 134.105 164.425 135.015 164.440 ;
        RECT 134.105 164.420 135.025 164.425 ;
        RECT 134.105 164.410 135.030 164.420 ;
        RECT 134.105 164.400 135.035 164.410 ;
        RECT 134.105 164.395 135.045 164.400 ;
        RECT 134.105 164.385 135.055 164.395 ;
        RECT 134.105 164.380 135.065 164.385 ;
        RECT 134.105 163.930 134.365 164.380 ;
        RECT 134.730 164.375 135.065 164.380 ;
        RECT 134.730 164.370 135.080 164.375 ;
        RECT 134.730 164.360 135.095 164.370 ;
        RECT 134.730 164.355 135.120 164.360 ;
        RECT 135.665 164.355 135.895 164.750 ;
        RECT 134.730 164.350 135.895 164.355 ;
        RECT 134.760 164.315 135.895 164.350 ;
        RECT 134.795 164.290 135.895 164.315 ;
        RECT 134.825 164.260 135.895 164.290 ;
        RECT 134.845 164.230 135.895 164.260 ;
        RECT 134.865 164.200 135.895 164.230 ;
        RECT 134.935 164.190 135.895 164.200 ;
        RECT 134.960 164.180 135.895 164.190 ;
        RECT 134.980 164.165 135.895 164.180 ;
        RECT 135.000 164.150 135.895 164.165 ;
        RECT 135.005 164.140 135.790 164.150 ;
        RECT 135.020 164.105 135.790 164.140 ;
        RECT 134.535 163.785 134.865 164.030 ;
        RECT 135.035 163.855 135.790 164.105 ;
        RECT 136.065 163.975 136.235 165.005 ;
        RECT 136.455 165.000 136.785 165.435 ;
        RECT 136.955 165.045 137.125 165.655 ;
        RECT 136.405 164.915 136.785 165.000 ;
        RECT 137.295 164.915 137.625 165.440 ;
        RECT 137.885 165.125 138.095 165.655 ;
        RECT 138.370 165.205 139.155 165.375 ;
        RECT 139.325 165.205 139.730 165.375 ;
        RECT 136.405 164.875 136.630 164.915 ;
        RECT 136.405 164.295 136.575 164.875 ;
        RECT 137.295 164.745 137.495 164.915 ;
        RECT 138.370 164.745 138.540 165.205 ;
        RECT 136.745 164.415 137.495 164.745 ;
        RECT 137.665 164.415 138.540 164.745 ;
        RECT 136.405 164.245 136.620 164.295 ;
        RECT 136.405 164.165 136.795 164.245 ;
        RECT 134.535 163.760 134.720 163.785 ;
        RECT 133.595 163.275 133.935 163.535 ;
        RECT 134.105 163.660 134.720 163.760 ;
        RECT 134.105 163.105 134.710 163.660 ;
        RECT 134.885 163.275 135.365 163.615 ;
        RECT 135.535 163.105 135.790 163.650 ;
        RECT 135.960 163.275 136.235 163.975 ;
        RECT 136.465 163.320 136.795 164.165 ;
        RECT 137.305 164.210 137.495 164.415 ;
        RECT 136.965 163.105 137.135 164.115 ;
        RECT 137.305 163.835 138.200 164.210 ;
        RECT 137.305 163.275 137.645 163.835 ;
        RECT 137.875 163.105 138.190 163.605 ;
        RECT 138.370 163.575 138.540 164.415 ;
        RECT 138.710 164.705 139.175 165.035 ;
        RECT 139.560 164.975 139.730 165.205 ;
        RECT 139.910 165.155 140.280 165.655 ;
        RECT 140.600 165.205 141.275 165.375 ;
        RECT 141.470 165.205 141.805 165.375 ;
        RECT 138.710 163.745 139.030 164.705 ;
        RECT 139.560 164.675 140.390 164.975 ;
        RECT 139.200 163.775 139.390 164.495 ;
        RECT 139.560 163.605 139.730 164.675 ;
        RECT 140.190 164.645 140.390 164.675 ;
        RECT 139.900 164.425 140.070 164.495 ;
        RECT 140.600 164.425 140.770 165.205 ;
        RECT 141.635 165.065 141.805 165.205 ;
        RECT 141.975 165.195 142.225 165.655 ;
        RECT 139.900 164.255 140.770 164.425 ;
        RECT 140.940 164.785 141.465 165.005 ;
        RECT 141.635 164.935 141.860 165.065 ;
        RECT 139.900 164.165 140.410 164.255 ;
        RECT 138.370 163.405 139.255 163.575 ;
        RECT 139.480 163.275 139.730 163.605 ;
        RECT 139.900 163.105 140.070 163.905 ;
        RECT 140.240 163.550 140.410 164.165 ;
        RECT 140.940 164.085 141.110 164.785 ;
        RECT 140.580 163.720 141.110 164.085 ;
        RECT 141.280 164.020 141.520 164.615 ;
        RECT 141.690 163.830 141.860 164.935 ;
        RECT 142.030 164.075 142.310 165.025 ;
        RECT 141.555 163.700 141.860 163.830 ;
        RECT 140.240 163.380 141.345 163.550 ;
        RECT 141.555 163.275 141.805 163.700 ;
        RECT 141.975 163.105 142.240 163.565 ;
        RECT 142.480 163.275 142.665 165.395 ;
        RECT 142.835 165.275 143.165 165.655 ;
        RECT 143.335 165.105 143.505 165.395 ;
        RECT 143.765 165.110 149.110 165.655 ;
        RECT 142.840 164.935 143.505 165.105 ;
        RECT 142.840 163.945 143.070 164.935 ;
        RECT 143.240 164.115 143.590 164.765 ;
        RECT 145.350 164.280 145.690 165.110 ;
        RECT 149.285 164.885 150.955 165.655 ;
        RECT 151.585 164.930 151.875 165.655 ;
        RECT 152.045 164.885 155.555 165.655 ;
        RECT 155.725 164.905 156.935 165.655 ;
        RECT 142.840 163.775 143.505 163.945 ;
        RECT 142.835 163.105 143.165 163.605 ;
        RECT 143.335 163.275 143.505 163.775 ;
        RECT 147.170 163.540 147.520 164.790 ;
        RECT 149.285 164.365 150.035 164.885 ;
        RECT 150.205 164.195 150.955 164.715 ;
        RECT 152.045 164.365 153.695 164.885 ;
        RECT 143.765 163.105 149.110 163.540 ;
        RECT 149.285 163.105 150.955 164.195 ;
        RECT 151.585 163.105 151.875 164.270 ;
        RECT 153.865 164.195 155.555 164.715 ;
        RECT 152.045 163.105 155.555 164.195 ;
        RECT 155.725 164.195 156.245 164.735 ;
        RECT 156.415 164.365 156.935 164.905 ;
        RECT 155.725 163.105 156.935 164.195 ;
        RECT 22.700 162.935 157.020 163.105 ;
        RECT 22.785 161.845 23.995 162.935 ;
        RECT 24.255 162.265 24.425 162.765 ;
        RECT 24.595 162.435 24.925 162.935 ;
        RECT 24.255 162.095 24.920 162.265 ;
        RECT 22.785 161.135 23.305 161.675 ;
        RECT 23.475 161.305 23.995 161.845 ;
        RECT 24.170 161.275 24.520 161.925 ;
        RECT 22.785 160.385 23.995 161.135 ;
        RECT 24.690 161.105 24.920 162.095 ;
        RECT 24.255 160.935 24.920 161.105 ;
        RECT 24.255 160.645 24.425 160.935 ;
        RECT 24.595 160.385 24.925 160.765 ;
        RECT 25.095 160.645 25.280 162.765 ;
        RECT 25.520 162.475 25.785 162.935 ;
        RECT 25.955 162.340 26.205 162.765 ;
        RECT 26.415 162.490 27.520 162.660 ;
        RECT 25.900 162.210 26.205 162.340 ;
        RECT 25.450 161.015 25.730 161.965 ;
        RECT 25.900 161.105 26.070 162.210 ;
        RECT 26.240 161.425 26.480 162.020 ;
        RECT 26.650 161.955 27.180 162.320 ;
        RECT 26.650 161.255 26.820 161.955 ;
        RECT 27.350 161.875 27.520 162.490 ;
        RECT 27.690 162.135 27.860 162.935 ;
        RECT 28.030 162.435 28.280 162.765 ;
        RECT 28.505 162.465 29.390 162.635 ;
        RECT 27.350 161.785 27.860 161.875 ;
        RECT 25.900 160.975 26.125 161.105 ;
        RECT 26.295 161.035 26.820 161.255 ;
        RECT 26.990 161.615 27.860 161.785 ;
        RECT 25.535 160.385 25.785 160.845 ;
        RECT 25.955 160.835 26.125 160.975 ;
        RECT 26.990 160.835 27.160 161.615 ;
        RECT 27.690 161.545 27.860 161.615 ;
        RECT 27.370 161.365 27.570 161.395 ;
        RECT 28.030 161.365 28.200 162.435 ;
        RECT 28.370 161.545 28.560 162.265 ;
        RECT 27.370 161.065 28.200 161.365 ;
        RECT 28.730 161.335 29.050 162.295 ;
        RECT 25.955 160.665 26.290 160.835 ;
        RECT 26.485 160.665 27.160 160.835 ;
        RECT 27.480 160.385 27.850 160.885 ;
        RECT 28.030 160.835 28.200 161.065 ;
        RECT 28.585 161.005 29.050 161.335 ;
        RECT 29.220 161.625 29.390 162.465 ;
        RECT 29.570 162.435 29.885 162.935 ;
        RECT 30.115 162.205 30.455 162.765 ;
        RECT 29.560 161.830 30.455 162.205 ;
        RECT 30.625 161.925 30.795 162.935 ;
        RECT 30.265 161.625 30.455 161.830 ;
        RECT 30.965 161.875 31.295 162.720 ;
        RECT 31.525 162.425 31.785 162.935 ;
        RECT 30.965 161.795 31.355 161.875 ;
        RECT 31.140 161.745 31.355 161.795 ;
        RECT 29.220 161.295 30.095 161.625 ;
        RECT 30.265 161.295 31.015 161.625 ;
        RECT 29.220 160.835 29.390 161.295 ;
        RECT 30.265 161.125 30.465 161.295 ;
        RECT 31.185 161.165 31.355 161.745 ;
        RECT 31.525 161.375 31.865 162.255 ;
        RECT 32.035 161.545 32.205 162.765 ;
        RECT 32.445 162.430 33.060 162.935 ;
        RECT 32.445 161.895 32.695 162.260 ;
        RECT 32.865 162.255 33.060 162.430 ;
        RECT 33.230 162.425 33.705 162.765 ;
        RECT 33.875 162.390 34.090 162.935 ;
        RECT 32.865 162.065 33.195 162.255 ;
        RECT 33.415 161.895 34.130 162.190 ;
        RECT 34.300 162.065 34.575 162.765 ;
        RECT 32.445 161.725 34.235 161.895 ;
        RECT 32.035 161.295 32.830 161.545 ;
        RECT 32.035 161.205 32.285 161.295 ;
        RECT 31.130 161.125 31.355 161.165 ;
        RECT 28.030 160.665 28.435 160.835 ;
        RECT 28.605 160.665 29.390 160.835 ;
        RECT 29.665 160.385 29.875 160.915 ;
        RECT 30.135 160.600 30.465 161.125 ;
        RECT 30.975 161.040 31.355 161.125 ;
        RECT 30.635 160.385 30.805 160.995 ;
        RECT 30.975 160.605 31.305 161.040 ;
        RECT 31.525 160.385 31.785 161.205 ;
        RECT 31.955 160.785 32.285 161.205 ;
        RECT 33.000 160.870 33.255 161.725 ;
        RECT 32.465 160.605 33.255 160.870 ;
        RECT 33.425 161.025 33.835 161.545 ;
        RECT 34.005 161.295 34.235 161.725 ;
        RECT 34.405 161.035 34.575 162.065 ;
        RECT 35.665 161.770 35.955 162.935 ;
        RECT 36.215 162.265 36.385 162.765 ;
        RECT 36.555 162.435 36.885 162.935 ;
        RECT 36.215 162.095 36.880 162.265 ;
        RECT 36.130 161.275 36.480 161.925 ;
        RECT 33.425 160.605 33.625 161.025 ;
        RECT 33.815 160.385 34.145 160.845 ;
        RECT 34.315 160.555 34.575 161.035 ;
        RECT 35.665 160.385 35.955 161.110 ;
        RECT 36.650 161.105 36.880 162.095 ;
        RECT 36.215 160.935 36.880 161.105 ;
        RECT 36.215 160.645 36.385 160.935 ;
        RECT 36.555 160.385 36.885 160.765 ;
        RECT 37.055 160.645 37.240 162.765 ;
        RECT 37.480 162.475 37.745 162.935 ;
        RECT 37.915 162.340 38.165 162.765 ;
        RECT 38.375 162.490 39.480 162.660 ;
        RECT 37.860 162.210 38.165 162.340 ;
        RECT 37.410 161.015 37.690 161.965 ;
        RECT 37.860 161.105 38.030 162.210 ;
        RECT 38.200 161.425 38.440 162.020 ;
        RECT 38.610 161.955 39.140 162.320 ;
        RECT 38.610 161.255 38.780 161.955 ;
        RECT 39.310 161.875 39.480 162.490 ;
        RECT 39.650 162.135 39.820 162.935 ;
        RECT 39.990 162.435 40.240 162.765 ;
        RECT 40.465 162.465 41.350 162.635 ;
        RECT 39.310 161.785 39.820 161.875 ;
        RECT 37.860 160.975 38.085 161.105 ;
        RECT 38.255 161.035 38.780 161.255 ;
        RECT 38.950 161.615 39.820 161.785 ;
        RECT 37.495 160.385 37.745 160.845 ;
        RECT 37.915 160.835 38.085 160.975 ;
        RECT 38.950 160.835 39.120 161.615 ;
        RECT 39.650 161.545 39.820 161.615 ;
        RECT 39.330 161.365 39.530 161.395 ;
        RECT 39.990 161.365 40.160 162.435 ;
        RECT 40.330 161.545 40.520 162.265 ;
        RECT 39.330 161.065 40.160 161.365 ;
        RECT 40.690 161.335 41.010 162.295 ;
        RECT 37.915 160.665 38.250 160.835 ;
        RECT 38.445 160.665 39.120 160.835 ;
        RECT 39.440 160.385 39.810 160.885 ;
        RECT 39.990 160.835 40.160 161.065 ;
        RECT 40.545 161.005 41.010 161.335 ;
        RECT 41.180 161.625 41.350 162.465 ;
        RECT 41.530 162.435 41.845 162.935 ;
        RECT 42.075 162.205 42.415 162.765 ;
        RECT 41.520 161.830 42.415 162.205 ;
        RECT 42.585 161.925 42.755 162.935 ;
        RECT 42.225 161.625 42.415 161.830 ;
        RECT 42.925 161.875 43.255 162.720 ;
        RECT 43.485 162.065 43.760 162.765 ;
        RECT 43.930 162.390 44.185 162.935 ;
        RECT 44.355 162.425 44.835 162.765 ;
        RECT 45.010 162.380 45.615 162.935 ;
        RECT 45.000 162.280 45.615 162.380 ;
        RECT 45.000 162.255 45.185 162.280 ;
        RECT 42.925 161.795 43.315 161.875 ;
        RECT 43.100 161.745 43.315 161.795 ;
        RECT 41.180 161.295 42.055 161.625 ;
        RECT 42.225 161.295 42.975 161.625 ;
        RECT 41.180 160.835 41.350 161.295 ;
        RECT 42.225 161.125 42.425 161.295 ;
        RECT 43.145 161.165 43.315 161.745 ;
        RECT 43.090 161.125 43.315 161.165 ;
        RECT 39.990 160.665 40.395 160.835 ;
        RECT 40.565 160.665 41.350 160.835 ;
        RECT 41.625 160.385 41.835 160.915 ;
        RECT 42.095 160.600 42.425 161.125 ;
        RECT 42.935 161.040 43.315 161.125 ;
        RECT 42.595 160.385 42.765 160.995 ;
        RECT 42.935 160.605 43.265 161.040 ;
        RECT 43.485 161.035 43.655 162.065 ;
        RECT 43.930 161.935 44.685 162.185 ;
        RECT 44.855 162.010 45.185 162.255 ;
        RECT 43.930 161.900 44.700 161.935 ;
        RECT 43.930 161.890 44.715 161.900 ;
        RECT 43.825 161.875 44.720 161.890 ;
        RECT 43.825 161.860 44.740 161.875 ;
        RECT 43.825 161.850 44.760 161.860 ;
        RECT 43.825 161.840 44.785 161.850 ;
        RECT 43.825 161.810 44.855 161.840 ;
        RECT 43.825 161.780 44.875 161.810 ;
        RECT 43.825 161.750 44.895 161.780 ;
        RECT 43.825 161.725 44.925 161.750 ;
        RECT 43.825 161.690 44.960 161.725 ;
        RECT 43.825 161.685 44.990 161.690 ;
        RECT 43.825 161.290 44.055 161.685 ;
        RECT 44.600 161.680 44.990 161.685 ;
        RECT 44.625 161.670 44.990 161.680 ;
        RECT 44.640 161.665 44.990 161.670 ;
        RECT 44.655 161.660 44.990 161.665 ;
        RECT 45.355 161.660 45.615 162.110 ;
        RECT 44.655 161.655 45.615 161.660 ;
        RECT 44.665 161.645 45.615 161.655 ;
        RECT 44.675 161.640 45.615 161.645 ;
        RECT 44.685 161.630 45.615 161.640 ;
        RECT 44.690 161.620 45.615 161.630 ;
        RECT 44.695 161.615 45.615 161.620 ;
        RECT 44.705 161.600 45.615 161.615 ;
        RECT 44.710 161.585 45.615 161.600 ;
        RECT 44.720 161.560 45.615 161.585 ;
        RECT 44.225 161.090 44.555 161.515 ;
        RECT 43.485 160.555 43.745 161.035 ;
        RECT 43.915 160.385 44.165 160.925 ;
        RECT 44.335 160.605 44.555 161.090 ;
        RECT 44.725 161.490 45.615 161.560 ;
        RECT 44.725 160.765 44.895 161.490 ;
        RECT 45.065 160.935 45.615 161.320 ;
        RECT 44.725 160.595 45.615 160.765 ;
        RECT 46.715 160.565 46.975 162.755 ;
        RECT 47.145 162.205 47.485 162.935 ;
        RECT 47.665 162.025 47.935 162.755 ;
        RECT 47.165 161.805 47.935 162.025 ;
        RECT 48.115 162.045 48.345 162.755 ;
        RECT 48.515 162.225 48.845 162.935 ;
        RECT 49.015 162.045 49.275 162.755 ;
        RECT 48.115 161.805 49.275 162.045 ;
        RECT 49.465 162.085 49.725 162.765 ;
        RECT 49.895 162.155 50.145 162.935 ;
        RECT 50.395 162.385 50.645 162.765 ;
        RECT 50.815 162.555 51.170 162.935 ;
        RECT 52.175 162.545 52.510 162.765 ;
        RECT 51.775 162.385 52.005 162.425 ;
        RECT 50.395 162.185 52.005 162.385 ;
        RECT 50.395 162.175 51.230 162.185 ;
        RECT 51.820 162.095 52.005 162.185 ;
        RECT 47.165 161.135 47.455 161.805 ;
        RECT 47.635 161.315 48.100 161.625 ;
        RECT 48.280 161.315 48.805 161.625 ;
        RECT 47.165 160.935 48.395 161.135 ;
        RECT 47.235 160.385 47.905 160.755 ;
        RECT 48.085 160.565 48.395 160.935 ;
        RECT 48.575 160.675 48.805 161.315 ;
        RECT 48.985 161.295 49.285 161.625 ;
        RECT 48.985 160.385 49.275 161.115 ;
        RECT 49.465 160.885 49.635 162.085 ;
        RECT 51.335 161.985 51.665 162.015 ;
        RECT 49.865 161.925 51.665 161.985 ;
        RECT 52.255 161.925 52.510 162.545 ;
        RECT 52.800 162.305 53.085 162.765 ;
        RECT 53.255 162.475 53.525 162.935 ;
        RECT 52.800 162.085 53.755 162.305 ;
        RECT 49.805 161.815 52.510 161.925 ;
        RECT 49.805 161.780 50.005 161.815 ;
        RECT 49.805 161.205 49.975 161.780 ;
        RECT 51.335 161.755 52.510 161.815 ;
        RECT 50.205 161.340 50.615 161.645 ;
        RECT 50.785 161.375 51.115 161.585 ;
        RECT 49.805 161.085 50.075 161.205 ;
        RECT 49.805 161.040 50.650 161.085 ;
        RECT 49.895 160.915 50.650 161.040 ;
        RECT 50.905 160.975 51.115 161.375 ;
        RECT 51.360 161.375 51.835 161.585 ;
        RECT 52.025 161.375 52.515 161.575 ;
        RECT 51.360 160.975 51.580 161.375 ;
        RECT 52.685 161.355 53.375 161.915 ;
        RECT 53.545 161.185 53.755 162.085 ;
        RECT 49.465 160.555 49.725 160.885 ;
        RECT 50.480 160.765 50.650 160.915 ;
        RECT 49.895 160.385 50.225 160.745 ;
        RECT 50.480 160.555 51.780 160.765 ;
        RECT 52.055 160.385 52.510 161.150 ;
        RECT 52.800 161.015 53.755 161.185 ;
        RECT 53.925 161.915 54.325 162.765 ;
        RECT 54.515 162.305 54.795 162.765 ;
        RECT 55.315 162.475 55.640 162.935 ;
        RECT 54.515 162.085 55.640 162.305 ;
        RECT 53.925 161.355 55.020 161.915 ;
        RECT 55.190 161.625 55.640 162.085 ;
        RECT 55.810 161.795 56.195 162.765 ;
        RECT 56.480 162.305 56.765 162.765 ;
        RECT 56.935 162.475 57.205 162.935 ;
        RECT 56.480 162.085 57.435 162.305 ;
        RECT 52.800 160.555 53.085 161.015 ;
        RECT 53.255 160.385 53.525 160.845 ;
        RECT 53.925 160.555 54.325 161.355 ;
        RECT 55.190 161.295 55.745 161.625 ;
        RECT 55.190 161.185 55.640 161.295 ;
        RECT 54.515 161.015 55.640 161.185 ;
        RECT 55.915 161.125 56.195 161.795 ;
        RECT 56.365 161.355 57.055 161.915 ;
        RECT 57.225 161.185 57.435 162.085 ;
        RECT 54.515 160.555 54.795 161.015 ;
        RECT 55.315 160.385 55.640 160.845 ;
        RECT 55.810 160.555 56.195 161.125 ;
        RECT 56.480 161.015 57.435 161.185 ;
        RECT 57.605 161.915 58.005 162.765 ;
        RECT 58.195 162.305 58.475 162.765 ;
        RECT 58.995 162.475 59.320 162.935 ;
        RECT 58.195 162.085 59.320 162.305 ;
        RECT 57.605 161.355 58.700 161.915 ;
        RECT 58.870 161.625 59.320 162.085 ;
        RECT 59.490 161.795 59.875 162.765 ;
        RECT 60.045 161.845 61.255 162.935 ;
        RECT 56.480 160.555 56.765 161.015 ;
        RECT 56.935 160.385 57.205 160.845 ;
        RECT 57.605 160.555 58.005 161.355 ;
        RECT 58.870 161.295 59.425 161.625 ;
        RECT 58.870 161.185 59.320 161.295 ;
        RECT 58.195 161.015 59.320 161.185 ;
        RECT 59.595 161.125 59.875 161.795 ;
        RECT 58.195 160.555 58.475 161.015 ;
        RECT 58.995 160.385 59.320 160.845 ;
        RECT 59.490 160.555 59.875 161.125 ;
        RECT 60.045 161.135 60.565 161.675 ;
        RECT 60.735 161.305 61.255 161.845 ;
        RECT 61.425 161.770 61.715 162.935 ;
        RECT 61.885 162.065 62.160 162.765 ;
        RECT 62.330 162.390 62.585 162.935 ;
        RECT 62.755 162.425 63.235 162.765 ;
        RECT 63.410 162.380 64.015 162.935 ;
        RECT 64.185 162.500 69.530 162.935 ;
        RECT 63.400 162.280 64.015 162.380 ;
        RECT 63.400 162.255 63.585 162.280 ;
        RECT 60.045 160.385 61.255 161.135 ;
        RECT 61.425 160.385 61.715 161.110 ;
        RECT 61.885 161.035 62.055 162.065 ;
        RECT 62.330 161.935 63.085 162.185 ;
        RECT 63.255 162.010 63.585 162.255 ;
        RECT 62.330 161.900 63.100 161.935 ;
        RECT 62.330 161.890 63.115 161.900 ;
        RECT 62.225 161.875 63.120 161.890 ;
        RECT 62.225 161.860 63.140 161.875 ;
        RECT 62.225 161.850 63.160 161.860 ;
        RECT 62.225 161.840 63.185 161.850 ;
        RECT 62.225 161.810 63.255 161.840 ;
        RECT 62.225 161.780 63.275 161.810 ;
        RECT 62.225 161.750 63.295 161.780 ;
        RECT 62.225 161.725 63.325 161.750 ;
        RECT 62.225 161.690 63.360 161.725 ;
        RECT 62.225 161.685 63.390 161.690 ;
        RECT 62.225 161.290 62.455 161.685 ;
        RECT 63.000 161.680 63.390 161.685 ;
        RECT 63.025 161.670 63.390 161.680 ;
        RECT 63.040 161.665 63.390 161.670 ;
        RECT 63.055 161.660 63.390 161.665 ;
        RECT 63.755 161.660 64.015 162.110 ;
        RECT 63.055 161.655 64.015 161.660 ;
        RECT 63.065 161.645 64.015 161.655 ;
        RECT 63.075 161.640 64.015 161.645 ;
        RECT 63.085 161.630 64.015 161.640 ;
        RECT 63.090 161.620 64.015 161.630 ;
        RECT 63.095 161.615 64.015 161.620 ;
        RECT 63.105 161.600 64.015 161.615 ;
        RECT 63.110 161.585 64.015 161.600 ;
        RECT 63.120 161.560 64.015 161.585 ;
        RECT 62.625 161.090 62.955 161.515 ;
        RECT 61.885 160.555 62.145 161.035 ;
        RECT 62.315 160.385 62.565 160.925 ;
        RECT 62.735 160.605 62.955 161.090 ;
        RECT 63.125 161.490 64.015 161.560 ;
        RECT 63.125 160.765 63.295 161.490 ;
        RECT 63.465 160.935 64.015 161.320 ;
        RECT 65.770 160.930 66.110 161.760 ;
        RECT 67.590 161.250 67.940 162.500 ;
        RECT 70.685 161.875 71.015 162.720 ;
        RECT 71.185 161.925 71.355 162.935 ;
        RECT 71.525 162.205 71.865 162.765 ;
        RECT 72.095 162.435 72.410 162.935 ;
        RECT 72.590 162.465 73.475 162.635 ;
        RECT 70.625 161.795 71.015 161.875 ;
        RECT 71.525 161.830 72.420 162.205 ;
        RECT 70.625 161.745 70.840 161.795 ;
        RECT 70.625 161.165 70.795 161.745 ;
        RECT 71.525 161.625 71.715 161.830 ;
        RECT 72.590 161.625 72.760 162.465 ;
        RECT 73.700 162.435 73.950 162.765 ;
        RECT 70.965 161.295 71.715 161.625 ;
        RECT 71.885 161.295 72.760 161.625 ;
        RECT 70.625 161.125 70.850 161.165 ;
        RECT 71.515 161.125 71.715 161.295 ;
        RECT 70.625 161.040 71.005 161.125 ;
        RECT 63.125 160.595 64.015 160.765 ;
        RECT 64.185 160.385 69.530 160.930 ;
        RECT 70.675 160.605 71.005 161.040 ;
        RECT 71.175 160.385 71.345 160.995 ;
        RECT 71.515 160.600 71.845 161.125 ;
        RECT 72.105 160.385 72.315 160.915 ;
        RECT 72.590 160.835 72.760 161.295 ;
        RECT 72.930 161.335 73.250 162.295 ;
        RECT 73.420 161.545 73.610 162.265 ;
        RECT 73.780 161.365 73.950 162.435 ;
        RECT 74.120 162.135 74.290 162.935 ;
        RECT 74.460 162.490 75.565 162.660 ;
        RECT 74.460 161.875 74.630 162.490 ;
        RECT 75.775 162.340 76.025 162.765 ;
        RECT 76.195 162.475 76.460 162.935 ;
        RECT 74.800 161.955 75.330 162.320 ;
        RECT 75.775 162.210 76.080 162.340 ;
        RECT 74.120 161.785 74.630 161.875 ;
        RECT 74.120 161.615 74.990 161.785 ;
        RECT 74.120 161.545 74.290 161.615 ;
        RECT 74.410 161.365 74.610 161.395 ;
        RECT 72.930 161.005 73.395 161.335 ;
        RECT 73.780 161.065 74.610 161.365 ;
        RECT 73.780 160.835 73.950 161.065 ;
        RECT 72.590 160.665 73.375 160.835 ;
        RECT 73.545 160.665 73.950 160.835 ;
        RECT 74.130 160.385 74.500 160.885 ;
        RECT 74.820 160.835 74.990 161.615 ;
        RECT 75.160 161.255 75.330 161.955 ;
        RECT 75.500 161.425 75.740 162.020 ;
        RECT 75.160 161.035 75.685 161.255 ;
        RECT 75.910 161.105 76.080 162.210 ;
        RECT 75.855 160.975 76.080 161.105 ;
        RECT 76.250 161.015 76.530 161.965 ;
        RECT 75.855 160.835 76.025 160.975 ;
        RECT 74.820 160.665 75.495 160.835 ;
        RECT 75.690 160.665 76.025 160.835 ;
        RECT 76.195 160.385 76.445 160.845 ;
        RECT 76.700 160.645 76.885 162.765 ;
        RECT 77.055 162.435 77.385 162.935 ;
        RECT 77.555 162.265 77.725 162.765 ;
        RECT 77.060 162.095 77.725 162.265 ;
        RECT 77.060 161.105 77.290 162.095 ;
        RECT 77.460 161.275 77.810 161.925 ;
        RECT 77.985 161.845 79.655 162.935 ;
        RECT 77.985 161.155 78.735 161.675 ;
        RECT 78.905 161.325 79.655 161.845 ;
        RECT 80.095 161.745 80.425 162.935 ;
        RECT 80.595 161.965 80.925 162.765 ;
        RECT 81.095 162.135 81.265 162.935 ;
        RECT 81.435 161.965 81.765 162.765 ;
        RECT 81.935 162.135 82.625 162.935 ;
        RECT 82.795 161.965 83.125 162.765 ;
        RECT 83.295 162.135 83.465 162.935 ;
        RECT 83.635 162.305 83.965 162.765 ;
        RECT 84.135 162.475 84.305 162.935 ;
        RECT 84.475 162.305 84.805 162.765 ;
        RECT 83.635 161.965 84.805 162.305 ;
        RECT 84.975 162.135 85.145 162.935 ;
        RECT 85.315 161.965 85.645 162.765 ;
        RECT 80.595 161.745 85.645 161.965 ;
        RECT 85.815 161.745 86.505 162.935 ;
        RECT 86.675 161.745 87.015 162.765 ;
        RECT 87.185 161.770 87.475 162.935 ;
        RECT 87.650 161.795 87.985 162.765 ;
        RECT 88.155 161.795 88.325 162.935 ;
        RECT 88.495 162.595 90.525 162.765 ;
        RECT 80.600 161.375 82.310 161.575 ;
        RECT 82.620 161.375 83.830 161.575 ;
        RECT 84.000 161.375 84.305 161.745 ;
        RECT 84.475 161.375 86.095 161.575 ;
        RECT 86.320 161.375 86.670 161.575 ;
        RECT 84.135 161.205 84.305 161.375 ;
        RECT 85.815 161.205 86.095 161.375 ;
        RECT 86.840 161.205 87.015 161.745 ;
        RECT 77.060 160.935 77.725 161.105 ;
        RECT 77.055 160.385 77.385 160.765 ;
        RECT 77.555 160.645 77.725 160.935 ;
        RECT 77.985 160.385 79.655 161.155 ;
        RECT 80.095 160.385 80.425 161.205 ;
        RECT 80.595 161.015 83.965 161.205 ;
        RECT 80.595 160.555 80.925 161.015 ;
        RECT 81.095 160.385 81.265 160.845 ;
        RECT 81.435 160.555 81.765 161.015 ;
        RECT 82.375 160.935 83.965 161.015 ;
        RECT 84.135 160.935 85.645 161.205 ;
        RECT 85.815 161.015 87.015 161.205 ;
        RECT 87.650 161.125 87.820 161.795 ;
        RECT 88.495 161.625 88.665 162.595 ;
        RECT 87.990 161.295 88.245 161.625 ;
        RECT 88.470 161.295 88.665 161.625 ;
        RECT 88.835 162.255 89.960 162.425 ;
        RECT 88.075 161.125 88.245 161.295 ;
        RECT 88.835 161.125 89.005 162.255 ;
        RECT 81.935 160.385 82.185 160.845 ;
        RECT 82.375 160.555 86.065 160.765 ;
        RECT 86.255 160.385 86.505 160.845 ;
        RECT 86.675 160.555 87.015 161.015 ;
        RECT 87.185 160.385 87.475 161.110 ;
        RECT 87.650 160.555 87.905 161.125 ;
        RECT 88.075 160.955 89.005 161.125 ;
        RECT 89.175 161.915 90.185 162.085 ;
        RECT 89.175 161.115 89.345 161.915 ;
        RECT 89.550 161.575 89.825 161.715 ;
        RECT 89.545 161.405 89.825 161.575 ;
        RECT 88.830 160.920 89.005 160.955 ;
        RECT 88.075 160.385 88.405 160.785 ;
        RECT 88.830 160.555 89.360 160.920 ;
        RECT 89.550 160.555 89.825 161.405 ;
        RECT 89.995 160.555 90.185 161.915 ;
        RECT 90.355 161.930 90.525 162.595 ;
        RECT 90.695 162.175 90.865 162.935 ;
        RECT 91.100 162.175 91.615 162.585 ;
        RECT 90.355 161.740 91.105 161.930 ;
        RECT 91.275 161.365 91.615 162.175 ;
        RECT 92.350 162.135 92.605 162.935 ;
        RECT 92.775 161.965 93.105 162.765 ;
        RECT 93.275 162.135 93.445 162.935 ;
        RECT 93.615 161.965 93.945 162.765 ;
        RECT 90.385 161.195 91.615 161.365 ;
        RECT 92.245 161.795 93.945 161.965 ;
        RECT 94.115 161.795 94.375 162.935 ;
        RECT 94.545 162.500 99.890 162.935 ;
        RECT 92.245 161.205 92.525 161.795 ;
        RECT 92.695 161.375 93.445 161.625 ;
        RECT 93.615 161.375 94.375 161.625 ;
        RECT 90.365 160.385 90.875 160.920 ;
        RECT 91.095 160.590 91.340 161.195 ;
        RECT 92.245 160.955 93.105 161.205 ;
        RECT 93.275 161.015 94.375 161.185 ;
        RECT 92.355 160.765 92.685 160.785 ;
        RECT 93.275 160.765 93.525 161.015 ;
        RECT 92.355 160.555 93.525 160.765 ;
        RECT 93.695 160.385 93.865 160.845 ;
        RECT 94.035 160.555 94.375 161.015 ;
        RECT 96.130 160.930 96.470 161.760 ;
        RECT 97.950 161.250 98.300 162.500 ;
        RECT 100.615 162.005 100.785 162.765 ;
        RECT 101.000 162.175 101.330 162.935 ;
        RECT 100.615 161.835 101.330 162.005 ;
        RECT 101.500 161.860 101.755 162.765 ;
        RECT 100.525 161.285 100.880 161.655 ;
        RECT 101.160 161.625 101.330 161.835 ;
        RECT 101.160 161.295 101.415 161.625 ;
        RECT 101.160 161.105 101.330 161.295 ;
        RECT 101.585 161.130 101.755 161.860 ;
        RECT 101.930 161.785 102.190 162.935 ;
        RECT 102.365 161.965 102.675 162.765 ;
        RECT 102.845 162.135 103.155 162.935 ;
        RECT 103.325 162.305 103.585 162.765 ;
        RECT 103.755 162.475 104.010 162.935 ;
        RECT 104.185 162.305 104.445 162.765 ;
        RECT 103.325 162.135 104.445 162.305 ;
        RECT 102.365 161.795 103.395 161.965 ;
        RECT 100.615 160.935 101.330 161.105 ;
        RECT 94.545 160.385 99.890 160.930 ;
        RECT 100.615 160.555 100.785 160.935 ;
        RECT 101.000 160.385 101.330 160.765 ;
        RECT 101.500 160.555 101.755 161.130 ;
        RECT 101.930 160.385 102.190 161.225 ;
        RECT 102.365 160.885 102.535 161.795 ;
        RECT 102.705 161.055 103.055 161.625 ;
        RECT 103.225 161.545 103.395 161.795 ;
        RECT 104.185 161.885 104.445 162.135 ;
        RECT 104.615 162.065 104.900 162.935 ;
        RECT 105.675 162.265 105.845 162.765 ;
        RECT 106.015 162.435 106.345 162.935 ;
        RECT 105.675 162.095 106.340 162.265 ;
        RECT 104.185 161.715 104.940 161.885 ;
        RECT 103.225 161.375 104.365 161.545 ;
        RECT 104.535 161.205 104.940 161.715 ;
        RECT 105.590 161.275 105.940 161.925 ;
        RECT 103.290 161.035 104.940 161.205 ;
        RECT 106.110 161.105 106.340 162.095 ;
        RECT 102.365 160.555 102.665 160.885 ;
        RECT 102.835 160.385 103.110 160.865 ;
        RECT 103.290 160.645 103.585 161.035 ;
        RECT 103.755 160.385 104.010 160.865 ;
        RECT 104.185 160.645 104.445 161.035 ;
        RECT 105.675 160.935 106.340 161.105 ;
        RECT 104.615 160.385 104.895 160.865 ;
        RECT 105.675 160.645 105.845 160.935 ;
        RECT 106.015 160.385 106.345 160.765 ;
        RECT 106.515 160.645 106.700 162.765 ;
        RECT 106.940 162.475 107.205 162.935 ;
        RECT 107.375 162.340 107.625 162.765 ;
        RECT 107.835 162.490 108.940 162.660 ;
        RECT 107.320 162.210 107.625 162.340 ;
        RECT 106.870 161.015 107.150 161.965 ;
        RECT 107.320 161.105 107.490 162.210 ;
        RECT 107.660 161.425 107.900 162.020 ;
        RECT 108.070 161.955 108.600 162.320 ;
        RECT 108.070 161.255 108.240 161.955 ;
        RECT 108.770 161.875 108.940 162.490 ;
        RECT 109.110 162.135 109.280 162.935 ;
        RECT 109.450 162.435 109.700 162.765 ;
        RECT 109.925 162.465 110.810 162.635 ;
        RECT 108.770 161.785 109.280 161.875 ;
        RECT 107.320 160.975 107.545 161.105 ;
        RECT 107.715 161.035 108.240 161.255 ;
        RECT 108.410 161.615 109.280 161.785 ;
        RECT 106.955 160.385 107.205 160.845 ;
        RECT 107.375 160.835 107.545 160.975 ;
        RECT 108.410 160.835 108.580 161.615 ;
        RECT 109.110 161.545 109.280 161.615 ;
        RECT 108.790 161.365 108.990 161.395 ;
        RECT 109.450 161.365 109.620 162.435 ;
        RECT 109.790 161.545 109.980 162.265 ;
        RECT 108.790 161.065 109.620 161.365 ;
        RECT 110.150 161.335 110.470 162.295 ;
        RECT 107.375 160.665 107.710 160.835 ;
        RECT 107.905 160.665 108.580 160.835 ;
        RECT 108.900 160.385 109.270 160.885 ;
        RECT 109.450 160.835 109.620 161.065 ;
        RECT 110.005 161.005 110.470 161.335 ;
        RECT 110.640 161.625 110.810 162.465 ;
        RECT 110.990 162.435 111.305 162.935 ;
        RECT 111.535 162.205 111.875 162.765 ;
        RECT 110.980 161.830 111.875 162.205 ;
        RECT 112.045 161.925 112.215 162.935 ;
        RECT 111.685 161.625 111.875 161.830 ;
        RECT 112.385 161.875 112.715 162.720 ;
        RECT 112.385 161.795 112.775 161.875 ;
        RECT 112.560 161.745 112.775 161.795 ;
        RECT 112.945 161.770 113.235 162.935 ;
        RECT 113.405 161.795 113.790 162.765 ;
        RECT 113.960 162.475 114.285 162.935 ;
        RECT 114.805 162.305 115.085 162.765 ;
        RECT 113.960 162.085 115.085 162.305 ;
        RECT 110.640 161.295 111.515 161.625 ;
        RECT 111.685 161.295 112.435 161.625 ;
        RECT 110.640 160.835 110.810 161.295 ;
        RECT 111.685 161.125 111.885 161.295 ;
        RECT 112.605 161.165 112.775 161.745 ;
        RECT 112.550 161.125 112.775 161.165 ;
        RECT 109.450 160.665 109.855 160.835 ;
        RECT 110.025 160.665 110.810 160.835 ;
        RECT 111.085 160.385 111.295 160.915 ;
        RECT 111.555 160.600 111.885 161.125 ;
        RECT 112.395 161.040 112.775 161.125 ;
        RECT 113.405 161.125 113.685 161.795 ;
        RECT 113.960 161.625 114.410 162.085 ;
        RECT 115.275 161.915 115.675 162.765 ;
        RECT 116.075 162.475 116.345 162.935 ;
        RECT 116.515 162.305 116.800 162.765 ;
        RECT 113.855 161.295 114.410 161.625 ;
        RECT 114.580 161.355 115.675 161.915 ;
        RECT 113.960 161.185 114.410 161.295 ;
        RECT 112.055 160.385 112.225 160.995 ;
        RECT 112.395 160.605 112.725 161.040 ;
        RECT 112.945 160.385 113.235 161.110 ;
        RECT 113.405 160.555 113.790 161.125 ;
        RECT 113.960 161.015 115.085 161.185 ;
        RECT 113.960 160.385 114.285 160.845 ;
        RECT 114.805 160.555 115.085 161.015 ;
        RECT 115.275 160.555 115.675 161.355 ;
        RECT 115.845 162.085 116.800 162.305 ;
        RECT 115.845 161.185 116.055 162.085 ;
        RECT 116.225 161.355 116.915 161.915 ;
        RECT 117.545 161.795 117.930 162.765 ;
        RECT 118.100 162.475 118.425 162.935 ;
        RECT 118.945 162.305 119.225 162.765 ;
        RECT 118.100 162.085 119.225 162.305 ;
        RECT 115.845 161.015 116.800 161.185 ;
        RECT 116.075 160.385 116.345 160.845 ;
        RECT 116.515 160.555 116.800 161.015 ;
        RECT 117.545 161.125 117.825 161.795 ;
        RECT 118.100 161.625 118.550 162.085 ;
        RECT 119.415 161.915 119.815 162.765 ;
        RECT 120.215 162.475 120.485 162.935 ;
        RECT 120.655 162.305 120.940 162.765 ;
        RECT 117.995 161.295 118.550 161.625 ;
        RECT 118.720 161.355 119.815 161.915 ;
        RECT 118.100 161.185 118.550 161.295 ;
        RECT 117.545 160.555 117.930 161.125 ;
        RECT 118.100 161.015 119.225 161.185 ;
        RECT 118.100 160.385 118.425 160.845 ;
        RECT 118.945 160.555 119.225 161.015 ;
        RECT 119.415 160.555 119.815 161.355 ;
        RECT 119.985 162.085 120.940 162.305 ;
        RECT 121.225 162.085 121.485 162.765 ;
        RECT 121.655 162.155 121.905 162.935 ;
        RECT 122.155 162.385 122.405 162.765 ;
        RECT 122.575 162.555 122.930 162.935 ;
        RECT 123.935 162.545 124.270 162.765 ;
        RECT 123.535 162.385 123.765 162.425 ;
        RECT 122.155 162.185 123.765 162.385 ;
        RECT 122.155 162.175 122.990 162.185 ;
        RECT 123.580 162.095 123.765 162.185 ;
        RECT 119.985 161.185 120.195 162.085 ;
        RECT 120.365 161.355 121.055 161.915 ;
        RECT 119.985 161.015 120.940 161.185 ;
        RECT 120.215 160.385 120.485 160.845 ;
        RECT 120.655 160.555 120.940 161.015 ;
        RECT 121.225 160.885 121.395 162.085 ;
        RECT 123.095 161.985 123.425 162.015 ;
        RECT 121.625 161.925 123.425 161.985 ;
        RECT 124.015 161.925 124.270 162.545 ;
        RECT 121.565 161.815 124.270 161.925 ;
        RECT 121.565 161.780 121.765 161.815 ;
        RECT 121.565 161.205 121.735 161.780 ;
        RECT 123.095 161.755 124.270 161.815 ;
        RECT 125.455 161.925 125.625 162.765 ;
        RECT 125.795 162.595 126.965 162.765 ;
        RECT 125.795 162.095 126.125 162.595 ;
        RECT 126.635 162.555 126.965 162.595 ;
        RECT 127.155 162.515 127.510 162.935 ;
        RECT 126.295 162.335 126.525 162.425 ;
        RECT 127.680 162.335 127.930 162.765 ;
        RECT 126.295 162.095 127.930 162.335 ;
        RECT 128.100 162.175 128.430 162.935 ;
        RECT 128.600 162.095 128.855 162.765 ;
        RECT 125.455 161.755 128.515 161.925 ;
        RECT 121.965 161.340 122.375 161.645 ;
        RECT 122.545 161.375 122.875 161.585 ;
        RECT 121.565 161.085 121.835 161.205 ;
        RECT 121.565 161.040 122.410 161.085 ;
        RECT 121.655 160.915 122.410 161.040 ;
        RECT 122.665 160.975 122.875 161.375 ;
        RECT 123.120 161.375 123.595 161.585 ;
        RECT 123.785 161.375 124.275 161.575 ;
        RECT 125.370 161.375 125.720 161.585 ;
        RECT 125.890 161.375 126.335 161.575 ;
        RECT 126.505 161.375 126.980 161.575 ;
        RECT 123.120 160.975 123.340 161.375 ;
        RECT 121.225 160.555 121.485 160.885 ;
        RECT 122.240 160.765 122.410 160.915 ;
        RECT 121.655 160.385 121.985 160.745 ;
        RECT 122.240 160.555 123.540 160.765 ;
        RECT 123.815 160.385 124.270 161.150 ;
        RECT 125.455 161.035 126.520 161.205 ;
        RECT 125.455 160.555 125.625 161.035 ;
        RECT 125.795 160.385 126.125 160.865 ;
        RECT 126.350 160.805 126.520 161.035 ;
        RECT 126.700 160.975 126.980 161.375 ;
        RECT 127.250 161.375 127.580 161.575 ;
        RECT 127.750 161.405 128.125 161.575 ;
        RECT 127.750 161.375 128.115 161.405 ;
        RECT 127.250 160.975 127.535 161.375 ;
        RECT 128.345 161.205 128.515 161.755 ;
        RECT 127.715 161.035 128.515 161.205 ;
        RECT 127.715 160.805 127.885 161.035 ;
        RECT 128.685 160.965 128.855 162.095 ;
        RECT 129.045 161.845 130.715 162.935 ;
        RECT 128.670 160.895 128.855 160.965 ;
        RECT 128.645 160.885 128.855 160.895 ;
        RECT 126.350 160.555 127.885 160.805 ;
        RECT 128.055 160.385 128.385 160.865 ;
        RECT 128.600 160.555 128.855 160.885 ;
        RECT 129.045 161.155 129.795 161.675 ;
        RECT 129.965 161.325 130.715 161.845 ;
        RECT 130.925 161.795 131.155 162.935 ;
        RECT 131.325 161.785 131.655 162.765 ;
        RECT 131.825 161.795 132.035 162.935 ;
        RECT 132.265 161.845 133.475 162.935 ;
        RECT 133.645 162.425 133.905 162.935 ;
        RECT 130.905 161.375 131.235 161.625 ;
        RECT 129.045 160.385 130.715 161.155 ;
        RECT 130.925 160.385 131.155 161.205 ;
        RECT 131.405 161.185 131.655 161.785 ;
        RECT 131.325 160.555 131.655 161.185 ;
        RECT 131.825 160.385 132.035 161.205 ;
        RECT 132.265 161.135 132.785 161.675 ;
        RECT 132.955 161.305 133.475 161.845 ;
        RECT 133.645 161.375 133.985 162.255 ;
        RECT 134.155 161.545 134.325 162.765 ;
        RECT 134.565 162.430 135.180 162.935 ;
        RECT 134.565 161.895 134.815 162.260 ;
        RECT 134.985 162.255 135.180 162.430 ;
        RECT 135.350 162.425 135.825 162.765 ;
        RECT 135.995 162.390 136.210 162.935 ;
        RECT 134.985 162.065 135.315 162.255 ;
        RECT 135.535 161.895 136.250 162.190 ;
        RECT 136.420 162.065 136.695 162.765 ;
        RECT 134.565 161.725 136.355 161.895 ;
        RECT 134.155 161.295 134.950 161.545 ;
        RECT 134.155 161.205 134.405 161.295 ;
        RECT 132.265 160.385 133.475 161.135 ;
        RECT 133.645 160.385 133.905 161.205 ;
        RECT 134.075 160.785 134.405 161.205 ;
        RECT 135.120 160.870 135.375 161.725 ;
        RECT 134.585 160.605 135.375 160.870 ;
        RECT 135.545 161.025 135.955 161.545 ;
        RECT 136.125 161.295 136.355 161.725 ;
        RECT 136.525 161.035 136.695 162.065 ;
        RECT 136.865 161.845 138.535 162.935 ;
        RECT 135.545 160.605 135.745 161.025 ;
        RECT 135.935 160.385 136.265 160.845 ;
        RECT 136.435 160.555 136.695 161.035 ;
        RECT 136.865 161.155 137.615 161.675 ;
        RECT 137.785 161.325 138.535 161.845 ;
        RECT 138.705 161.770 138.995 162.935 ;
        RECT 139.225 161.875 139.555 162.720 ;
        RECT 139.725 161.925 139.895 162.935 ;
        RECT 140.065 162.205 140.405 162.765 ;
        RECT 140.635 162.435 140.950 162.935 ;
        RECT 141.130 162.465 142.015 162.635 ;
        RECT 139.165 161.795 139.555 161.875 ;
        RECT 140.065 161.830 140.960 162.205 ;
        RECT 139.165 161.745 139.380 161.795 ;
        RECT 139.165 161.165 139.335 161.745 ;
        RECT 140.065 161.625 140.255 161.830 ;
        RECT 141.130 161.625 141.300 162.465 ;
        RECT 142.240 162.435 142.490 162.765 ;
        RECT 139.505 161.295 140.255 161.625 ;
        RECT 140.425 161.295 141.300 161.625 ;
        RECT 136.865 160.385 138.535 161.155 ;
        RECT 139.165 161.125 139.390 161.165 ;
        RECT 140.055 161.125 140.255 161.295 ;
        RECT 138.705 160.385 138.995 161.110 ;
        RECT 139.165 161.040 139.545 161.125 ;
        RECT 139.215 160.605 139.545 161.040 ;
        RECT 139.715 160.385 139.885 160.995 ;
        RECT 140.055 160.600 140.385 161.125 ;
        RECT 140.645 160.385 140.855 160.915 ;
        RECT 141.130 160.835 141.300 161.295 ;
        RECT 141.470 161.335 141.790 162.295 ;
        RECT 141.960 161.545 142.150 162.265 ;
        RECT 142.320 161.365 142.490 162.435 ;
        RECT 142.660 162.135 142.830 162.935 ;
        RECT 143.000 162.490 144.105 162.660 ;
        RECT 143.000 161.875 143.170 162.490 ;
        RECT 144.315 162.340 144.565 162.765 ;
        RECT 144.735 162.475 145.000 162.935 ;
        RECT 143.340 161.955 143.870 162.320 ;
        RECT 144.315 162.210 144.620 162.340 ;
        RECT 142.660 161.785 143.170 161.875 ;
        RECT 142.660 161.615 143.530 161.785 ;
        RECT 142.660 161.545 142.830 161.615 ;
        RECT 142.950 161.365 143.150 161.395 ;
        RECT 141.470 161.005 141.935 161.335 ;
        RECT 142.320 161.065 143.150 161.365 ;
        RECT 142.320 160.835 142.490 161.065 ;
        RECT 141.130 160.665 141.915 160.835 ;
        RECT 142.085 160.665 142.490 160.835 ;
        RECT 142.670 160.385 143.040 160.885 ;
        RECT 143.360 160.835 143.530 161.615 ;
        RECT 143.700 161.255 143.870 161.955 ;
        RECT 144.040 161.425 144.280 162.020 ;
        RECT 143.700 161.035 144.225 161.255 ;
        RECT 144.450 161.105 144.620 162.210 ;
        RECT 144.395 160.975 144.620 161.105 ;
        RECT 144.790 161.015 145.070 161.965 ;
        RECT 144.395 160.835 144.565 160.975 ;
        RECT 143.360 160.665 144.035 160.835 ;
        RECT 144.230 160.665 144.565 160.835 ;
        RECT 144.735 160.385 144.985 160.845 ;
        RECT 145.240 160.645 145.425 162.765 ;
        RECT 145.595 162.435 145.925 162.935 ;
        RECT 146.095 162.265 146.265 162.765 ;
        RECT 145.600 162.095 146.265 162.265 ;
        RECT 146.615 162.265 146.785 162.765 ;
        RECT 146.955 162.435 147.285 162.935 ;
        RECT 146.615 162.095 147.280 162.265 ;
        RECT 145.600 161.105 145.830 162.095 ;
        RECT 146.000 161.275 146.350 161.925 ;
        RECT 146.530 161.275 146.880 161.925 ;
        RECT 147.050 161.105 147.280 162.095 ;
        RECT 145.600 160.935 146.265 161.105 ;
        RECT 145.595 160.385 145.925 160.765 ;
        RECT 146.095 160.645 146.265 160.935 ;
        RECT 146.615 160.935 147.280 161.105 ;
        RECT 146.615 160.645 146.785 160.935 ;
        RECT 146.955 160.385 147.285 160.765 ;
        RECT 147.455 160.645 147.640 162.765 ;
        RECT 147.880 162.475 148.145 162.935 ;
        RECT 148.315 162.340 148.565 162.765 ;
        RECT 148.775 162.490 149.880 162.660 ;
        RECT 148.260 162.210 148.565 162.340 ;
        RECT 147.810 161.015 148.090 161.965 ;
        RECT 148.260 161.105 148.430 162.210 ;
        RECT 148.600 161.425 148.840 162.020 ;
        RECT 149.010 161.955 149.540 162.320 ;
        RECT 149.010 161.255 149.180 161.955 ;
        RECT 149.710 161.875 149.880 162.490 ;
        RECT 150.050 162.135 150.220 162.935 ;
        RECT 150.390 162.435 150.640 162.765 ;
        RECT 150.865 162.465 151.750 162.635 ;
        RECT 149.710 161.785 150.220 161.875 ;
        RECT 148.260 160.975 148.485 161.105 ;
        RECT 148.655 161.035 149.180 161.255 ;
        RECT 149.350 161.615 150.220 161.785 ;
        RECT 147.895 160.385 148.145 160.845 ;
        RECT 148.315 160.835 148.485 160.975 ;
        RECT 149.350 160.835 149.520 161.615 ;
        RECT 150.050 161.545 150.220 161.615 ;
        RECT 149.730 161.365 149.930 161.395 ;
        RECT 150.390 161.365 150.560 162.435 ;
        RECT 150.730 161.545 150.920 162.265 ;
        RECT 149.730 161.065 150.560 161.365 ;
        RECT 151.090 161.335 151.410 162.295 ;
        RECT 148.315 160.665 148.650 160.835 ;
        RECT 148.845 160.665 149.520 160.835 ;
        RECT 149.840 160.385 150.210 160.885 ;
        RECT 150.390 160.835 150.560 161.065 ;
        RECT 150.945 161.005 151.410 161.335 ;
        RECT 151.580 161.625 151.750 162.465 ;
        RECT 151.930 162.435 152.245 162.935 ;
        RECT 152.475 162.205 152.815 162.765 ;
        RECT 151.920 161.830 152.815 162.205 ;
        RECT 152.985 161.925 153.155 162.935 ;
        RECT 152.625 161.625 152.815 161.830 ;
        RECT 153.325 161.875 153.655 162.720 ;
        RECT 153.325 161.795 153.715 161.875 ;
        RECT 153.885 161.845 155.555 162.935 ;
        RECT 153.500 161.745 153.715 161.795 ;
        RECT 151.580 161.295 152.455 161.625 ;
        RECT 152.625 161.295 153.375 161.625 ;
        RECT 151.580 160.835 151.750 161.295 ;
        RECT 152.625 161.125 152.825 161.295 ;
        RECT 153.545 161.165 153.715 161.745 ;
        RECT 153.490 161.125 153.715 161.165 ;
        RECT 150.390 160.665 150.795 160.835 ;
        RECT 150.965 160.665 151.750 160.835 ;
        RECT 152.025 160.385 152.235 160.915 ;
        RECT 152.495 160.600 152.825 161.125 ;
        RECT 153.335 161.040 153.715 161.125 ;
        RECT 153.885 161.155 154.635 161.675 ;
        RECT 154.805 161.325 155.555 161.845 ;
        RECT 155.725 161.845 156.935 162.935 ;
        RECT 155.725 161.305 156.245 161.845 ;
        RECT 152.995 160.385 153.165 160.995 ;
        RECT 153.335 160.605 153.665 161.040 ;
        RECT 153.885 160.385 155.555 161.155 ;
        RECT 156.415 161.135 156.935 161.675 ;
        RECT 155.725 160.385 156.935 161.135 ;
        RECT 22.700 160.215 157.020 160.385 ;
        RECT 22.785 159.465 23.995 160.215 ;
        RECT 24.625 159.540 24.885 160.045 ;
        RECT 25.065 159.835 25.395 160.215 ;
        RECT 25.575 159.665 25.745 160.045 ;
        RECT 22.785 158.925 23.305 159.465 ;
        RECT 23.475 158.755 23.995 159.295 ;
        RECT 22.785 157.665 23.995 158.755 ;
        RECT 24.625 158.740 24.795 159.540 ;
        RECT 25.080 159.495 25.745 159.665 ;
        RECT 26.005 159.565 26.265 160.045 ;
        RECT 26.435 159.675 26.685 160.215 ;
        RECT 25.080 159.240 25.250 159.495 ;
        RECT 24.965 158.910 25.250 159.240 ;
        RECT 25.485 158.945 25.815 159.315 ;
        RECT 25.080 158.765 25.250 158.910 ;
        RECT 24.625 157.835 24.895 158.740 ;
        RECT 25.080 158.595 25.745 158.765 ;
        RECT 25.065 157.665 25.395 158.425 ;
        RECT 25.575 157.835 25.745 158.595 ;
        RECT 26.005 158.535 26.175 159.565 ;
        RECT 26.855 159.510 27.075 159.995 ;
        RECT 26.345 158.915 26.575 159.310 ;
        RECT 26.745 159.085 27.075 159.510 ;
        RECT 27.245 159.835 28.135 160.005 ;
        RECT 27.245 159.110 27.415 159.835 ;
        RECT 28.550 159.735 28.850 160.215 ;
        RECT 27.585 159.280 28.135 159.665 ;
        RECT 29.020 159.565 29.280 160.020 ;
        RECT 29.450 159.735 29.710 160.215 ;
        RECT 29.880 159.565 30.140 160.020 ;
        RECT 30.310 159.735 30.570 160.215 ;
        RECT 30.740 159.565 31.000 160.020 ;
        RECT 31.170 159.735 31.430 160.215 ;
        RECT 31.600 159.565 31.860 160.020 ;
        RECT 32.030 159.690 32.290 160.215 ;
        RECT 28.550 159.395 31.860 159.565 ;
        RECT 27.245 159.040 28.135 159.110 ;
        RECT 27.240 159.015 28.135 159.040 ;
        RECT 27.230 159.000 28.135 159.015 ;
        RECT 27.225 158.985 28.135 159.000 ;
        RECT 27.215 158.980 28.135 158.985 ;
        RECT 27.210 158.970 28.135 158.980 ;
        RECT 27.205 158.960 28.135 158.970 ;
        RECT 27.195 158.955 28.135 158.960 ;
        RECT 27.185 158.945 28.135 158.955 ;
        RECT 27.175 158.940 28.135 158.945 ;
        RECT 27.175 158.935 27.510 158.940 ;
        RECT 27.160 158.930 27.510 158.935 ;
        RECT 27.145 158.920 27.510 158.930 ;
        RECT 27.120 158.915 27.510 158.920 ;
        RECT 26.345 158.910 27.510 158.915 ;
        RECT 26.345 158.875 27.480 158.910 ;
        RECT 26.345 158.850 27.445 158.875 ;
        RECT 26.345 158.820 27.415 158.850 ;
        RECT 26.345 158.790 27.395 158.820 ;
        RECT 26.345 158.760 27.375 158.790 ;
        RECT 26.345 158.750 27.305 158.760 ;
        RECT 26.345 158.740 27.280 158.750 ;
        RECT 26.345 158.725 27.260 158.740 ;
        RECT 26.345 158.710 27.240 158.725 ;
        RECT 26.450 158.700 27.235 158.710 ;
        RECT 26.450 158.665 27.220 158.700 ;
        RECT 26.005 157.835 26.280 158.535 ;
        RECT 26.450 158.415 27.205 158.665 ;
        RECT 27.375 158.345 27.705 158.590 ;
        RECT 27.875 158.490 28.135 158.940 ;
        RECT 28.550 158.805 29.520 159.395 ;
        RECT 32.460 159.225 32.710 160.035 ;
        RECT 32.890 159.755 33.135 160.215 ;
        RECT 33.455 159.665 33.625 160.045 ;
        RECT 33.805 159.835 34.135 160.215 ;
        RECT 29.690 158.975 32.710 159.225 ;
        RECT 32.880 158.975 33.195 159.585 ;
        RECT 33.455 159.495 34.120 159.665 ;
        RECT 34.315 159.540 34.575 160.045 ;
        RECT 28.550 158.565 31.860 158.805 ;
        RECT 27.520 158.320 27.705 158.345 ;
        RECT 27.520 158.220 28.135 158.320 ;
        RECT 26.450 157.665 26.705 158.210 ;
        RECT 26.875 157.835 27.355 158.175 ;
        RECT 27.530 157.665 28.135 158.220 ;
        RECT 28.555 157.665 28.850 158.395 ;
        RECT 29.020 157.840 29.280 158.565 ;
        RECT 29.450 157.665 29.710 158.395 ;
        RECT 29.880 157.840 30.140 158.565 ;
        RECT 30.310 157.665 30.570 158.395 ;
        RECT 30.740 157.840 31.000 158.565 ;
        RECT 31.170 157.665 31.430 158.395 ;
        RECT 31.600 157.840 31.860 158.565 ;
        RECT 32.030 157.665 32.290 158.775 ;
        RECT 32.460 157.840 32.710 158.975 ;
        RECT 33.385 158.945 33.715 159.315 ;
        RECT 33.950 159.240 34.120 159.495 ;
        RECT 33.950 158.910 34.235 159.240 ;
        RECT 32.890 157.665 33.185 158.775 ;
        RECT 33.950 158.765 34.120 158.910 ;
        RECT 33.455 158.595 34.120 158.765 ;
        RECT 34.405 158.740 34.575 159.540 ;
        RECT 35.265 159.395 35.475 160.215 ;
        RECT 35.645 159.415 35.975 160.045 ;
        RECT 35.645 158.815 35.895 159.415 ;
        RECT 36.145 159.395 36.375 160.215 ;
        RECT 36.585 159.445 38.255 160.215 ;
        RECT 38.450 159.565 38.760 160.035 ;
        RECT 38.930 159.735 39.665 160.215 ;
        RECT 39.835 159.645 40.005 159.995 ;
        RECT 40.175 159.815 40.555 160.215 ;
        RECT 36.065 158.975 36.395 159.225 ;
        RECT 36.585 158.925 37.335 159.445 ;
        RECT 38.450 159.395 39.185 159.565 ;
        RECT 39.835 159.475 40.575 159.645 ;
        RECT 40.745 159.540 41.015 159.885 ;
        RECT 41.490 159.645 41.660 159.895 ;
        RECT 38.935 159.305 39.185 159.395 ;
        RECT 40.405 159.305 40.575 159.475 ;
        RECT 33.455 157.835 33.625 158.595 ;
        RECT 33.805 157.665 34.135 158.425 ;
        RECT 34.305 157.835 34.575 158.740 ;
        RECT 35.265 157.665 35.475 158.805 ;
        RECT 35.645 157.835 35.975 158.815 ;
        RECT 36.145 157.665 36.375 158.805 ;
        RECT 37.505 158.755 38.255 159.275 ;
        RECT 38.430 158.975 38.765 159.225 ;
        RECT 38.935 158.975 39.675 159.305 ;
        RECT 40.405 158.975 40.635 159.305 ;
        RECT 36.585 157.665 38.255 158.755 ;
        RECT 38.430 157.665 38.685 158.805 ;
        RECT 38.935 158.415 39.105 158.975 ;
        RECT 40.405 158.805 40.575 158.975 ;
        RECT 40.845 158.855 41.015 159.540 ;
        RECT 40.785 158.805 41.015 158.855 ;
        RECT 39.330 158.635 40.575 158.805 ;
        RECT 39.330 158.385 39.750 158.635 ;
        RECT 38.880 157.885 40.075 158.215 ;
        RECT 40.255 157.665 40.535 158.465 ;
        RECT 40.745 157.835 41.015 158.805 ;
        RECT 41.185 159.475 41.660 159.645 ;
        RECT 41.895 159.475 42.225 160.215 ;
        RECT 42.395 159.645 42.595 159.990 ;
        RECT 42.765 159.815 43.095 160.215 ;
        RECT 43.265 159.645 43.465 160.000 ;
        RECT 43.635 159.820 43.965 160.215 ;
        RECT 44.405 159.715 44.665 160.045 ;
        RECT 44.835 159.855 45.165 160.215 ;
        RECT 45.420 159.835 46.720 160.045 ;
        RECT 42.395 159.475 44.235 159.645 ;
        RECT 41.185 158.505 41.355 159.475 ;
        RECT 41.525 158.685 41.875 159.305 ;
        RECT 42.045 158.685 42.365 159.305 ;
        RECT 42.535 158.685 42.865 159.305 ;
        RECT 43.035 158.685 43.335 159.305 ;
        RECT 43.575 158.505 43.795 159.305 ;
        RECT 41.185 158.295 43.795 158.505 ;
        RECT 41.895 157.665 42.225 158.115 ;
        RECT 43.975 157.850 44.235 159.475 ;
        RECT 44.405 158.515 44.575 159.715 ;
        RECT 45.420 159.685 45.590 159.835 ;
        RECT 44.835 159.560 45.590 159.685 ;
        RECT 44.745 159.515 45.590 159.560 ;
        RECT 44.745 159.395 45.015 159.515 ;
        RECT 44.745 158.820 44.915 159.395 ;
        RECT 45.145 158.955 45.555 159.260 ;
        RECT 45.845 159.225 46.055 159.625 ;
        RECT 45.725 159.015 46.055 159.225 ;
        RECT 46.300 159.225 46.520 159.625 ;
        RECT 46.995 159.450 47.450 160.215 ;
        RECT 48.545 159.490 48.835 160.215 ;
        RECT 50.170 159.735 50.470 160.215 ;
        RECT 50.640 159.565 50.900 160.020 ;
        RECT 51.070 159.735 51.330 160.215 ;
        RECT 51.500 159.565 51.760 160.020 ;
        RECT 51.930 159.735 52.190 160.215 ;
        RECT 52.360 159.565 52.620 160.020 ;
        RECT 52.790 159.735 53.050 160.215 ;
        RECT 53.220 159.565 53.480 160.020 ;
        RECT 53.650 159.690 53.910 160.215 ;
        RECT 50.170 159.395 53.480 159.565 ;
        RECT 46.300 159.015 46.775 159.225 ;
        RECT 46.965 159.025 47.455 159.225 ;
        RECT 44.745 158.785 44.945 158.820 ;
        RECT 46.275 158.785 47.450 158.845 ;
        RECT 44.745 158.675 47.450 158.785 ;
        RECT 44.805 158.615 46.605 158.675 ;
        RECT 46.275 158.585 46.605 158.615 ;
        RECT 44.405 157.835 44.665 158.515 ;
        RECT 44.835 157.665 45.085 158.445 ;
        RECT 45.335 158.415 46.170 158.425 ;
        RECT 46.760 158.415 46.945 158.505 ;
        RECT 45.335 158.215 46.945 158.415 ;
        RECT 45.335 157.835 45.585 158.215 ;
        RECT 46.715 158.175 46.945 158.215 ;
        RECT 47.195 158.055 47.450 158.675 ;
        RECT 45.755 157.665 46.110 158.045 ;
        RECT 47.115 157.835 47.450 158.055 ;
        RECT 48.545 157.665 48.835 158.830 ;
        RECT 50.170 158.805 51.140 159.395 ;
        RECT 54.080 159.225 54.330 160.035 ;
        RECT 54.510 159.755 54.755 160.215 ;
        RECT 51.310 158.975 54.330 159.225 ;
        RECT 54.500 158.975 54.815 159.585 ;
        RECT 55.035 159.560 55.365 159.995 ;
        RECT 55.535 159.605 55.705 160.215 ;
        RECT 54.985 159.475 55.365 159.560 ;
        RECT 55.875 159.475 56.205 160.000 ;
        RECT 56.465 159.685 56.675 160.215 ;
        RECT 56.950 159.765 57.735 159.935 ;
        RECT 57.905 159.765 58.310 159.935 ;
        RECT 54.985 159.435 55.210 159.475 ;
        RECT 50.170 158.565 53.480 158.805 ;
        RECT 50.175 157.665 50.470 158.395 ;
        RECT 50.640 157.840 50.900 158.565 ;
        RECT 51.070 157.665 51.330 158.395 ;
        RECT 51.500 157.840 51.760 158.565 ;
        RECT 51.930 157.665 52.190 158.395 ;
        RECT 52.360 157.840 52.620 158.565 ;
        RECT 52.790 157.665 53.050 158.395 ;
        RECT 53.220 157.840 53.480 158.565 ;
        RECT 53.650 157.665 53.910 158.775 ;
        RECT 54.080 157.840 54.330 158.975 ;
        RECT 54.985 158.855 55.155 159.435 ;
        RECT 55.875 159.305 56.075 159.475 ;
        RECT 56.950 159.305 57.120 159.765 ;
        RECT 55.325 158.975 56.075 159.305 ;
        RECT 56.245 158.975 57.120 159.305 ;
        RECT 54.985 158.805 55.200 158.855 ;
        RECT 54.510 157.665 54.805 158.775 ;
        RECT 54.985 158.725 55.375 158.805 ;
        RECT 55.045 157.880 55.375 158.725 ;
        RECT 55.885 158.770 56.075 158.975 ;
        RECT 55.545 157.665 55.715 158.675 ;
        RECT 55.885 158.395 56.780 158.770 ;
        RECT 55.885 157.835 56.225 158.395 ;
        RECT 56.455 157.665 56.770 158.165 ;
        RECT 56.950 158.135 57.120 158.975 ;
        RECT 57.290 159.265 57.755 159.595 ;
        RECT 58.140 159.535 58.310 159.765 ;
        RECT 58.490 159.715 58.860 160.215 ;
        RECT 59.180 159.765 59.855 159.935 ;
        RECT 60.050 159.765 60.385 159.935 ;
        RECT 57.290 158.305 57.610 159.265 ;
        RECT 58.140 159.235 58.970 159.535 ;
        RECT 57.780 158.335 57.970 159.055 ;
        RECT 58.140 158.165 58.310 159.235 ;
        RECT 58.770 159.205 58.970 159.235 ;
        RECT 58.480 158.985 58.650 159.055 ;
        RECT 59.180 158.985 59.350 159.765 ;
        RECT 60.215 159.625 60.385 159.765 ;
        RECT 60.555 159.755 60.805 160.215 ;
        RECT 58.480 158.815 59.350 158.985 ;
        RECT 59.520 159.345 60.045 159.565 ;
        RECT 60.215 159.495 60.440 159.625 ;
        RECT 58.480 158.725 58.990 158.815 ;
        RECT 56.950 157.965 57.835 158.135 ;
        RECT 58.060 157.835 58.310 158.165 ;
        RECT 58.480 157.665 58.650 158.465 ;
        RECT 58.820 158.110 58.990 158.725 ;
        RECT 59.520 158.645 59.690 159.345 ;
        RECT 59.160 158.280 59.690 158.645 ;
        RECT 59.860 158.580 60.100 159.175 ;
        RECT 60.270 158.390 60.440 159.495 ;
        RECT 60.610 158.635 60.890 159.585 ;
        RECT 60.135 158.260 60.440 158.390 ;
        RECT 58.820 157.940 59.925 158.110 ;
        RECT 60.135 157.835 60.385 158.260 ;
        RECT 60.555 157.665 60.820 158.125 ;
        RECT 61.060 157.835 61.245 159.955 ;
        RECT 61.415 159.835 61.745 160.215 ;
        RECT 61.915 159.665 62.085 159.955 ;
        RECT 62.345 159.835 63.235 160.005 ;
        RECT 61.420 159.495 62.085 159.665 ;
        RECT 61.420 158.505 61.650 159.495 ;
        RECT 61.820 158.675 62.170 159.325 ;
        RECT 62.345 159.280 62.895 159.665 ;
        RECT 63.065 159.110 63.235 159.835 ;
        RECT 62.345 159.040 63.235 159.110 ;
        RECT 63.405 159.510 63.625 159.995 ;
        RECT 63.795 159.675 64.045 160.215 ;
        RECT 64.215 159.565 64.475 160.045 ;
        RECT 63.405 159.085 63.735 159.510 ;
        RECT 62.345 159.015 63.240 159.040 ;
        RECT 62.345 159.000 63.250 159.015 ;
        RECT 62.345 158.985 63.255 159.000 ;
        RECT 62.345 158.980 63.265 158.985 ;
        RECT 62.345 158.970 63.270 158.980 ;
        RECT 62.345 158.960 63.275 158.970 ;
        RECT 62.345 158.955 63.285 158.960 ;
        RECT 62.345 158.945 63.295 158.955 ;
        RECT 62.345 158.940 63.305 158.945 ;
        RECT 61.420 158.335 62.085 158.505 ;
        RECT 62.345 158.490 62.605 158.940 ;
        RECT 62.970 158.935 63.305 158.940 ;
        RECT 62.970 158.930 63.320 158.935 ;
        RECT 62.970 158.920 63.335 158.930 ;
        RECT 62.970 158.915 63.360 158.920 ;
        RECT 63.905 158.915 64.135 159.310 ;
        RECT 62.970 158.910 64.135 158.915 ;
        RECT 63.000 158.875 64.135 158.910 ;
        RECT 63.035 158.850 64.135 158.875 ;
        RECT 63.065 158.820 64.135 158.850 ;
        RECT 63.085 158.790 64.135 158.820 ;
        RECT 63.105 158.760 64.135 158.790 ;
        RECT 63.175 158.750 64.135 158.760 ;
        RECT 63.200 158.740 64.135 158.750 ;
        RECT 63.220 158.725 64.135 158.740 ;
        RECT 63.240 158.710 64.135 158.725 ;
        RECT 63.245 158.700 64.030 158.710 ;
        RECT 63.260 158.665 64.030 158.700 ;
        RECT 61.415 157.665 61.745 158.165 ;
        RECT 61.915 157.835 62.085 158.335 ;
        RECT 62.775 158.345 63.105 158.590 ;
        RECT 63.275 158.415 64.030 158.665 ;
        RECT 64.305 158.535 64.475 159.565 ;
        RECT 64.645 159.445 66.315 160.215 ;
        RECT 66.510 159.815 66.840 160.215 ;
        RECT 67.010 159.645 67.180 159.915 ;
        RECT 67.350 159.705 67.665 160.215 ;
        RECT 67.895 159.705 68.185 160.045 ;
        RECT 68.355 159.705 68.595 160.215 ;
        RECT 66.485 159.475 67.180 159.645 ;
        RECT 64.645 158.925 65.395 159.445 ;
        RECT 65.565 158.755 66.315 159.275 ;
        RECT 62.775 158.320 62.960 158.345 ;
        RECT 62.345 158.220 62.960 158.320 ;
        RECT 62.345 157.665 62.950 158.220 ;
        RECT 63.125 157.835 63.605 158.175 ;
        RECT 63.775 157.665 64.030 158.210 ;
        RECT 64.200 157.835 64.475 158.535 ;
        RECT 64.645 157.665 66.315 158.755 ;
        RECT 66.485 158.465 66.915 159.475 ;
        RECT 67.085 158.805 67.255 159.305 ;
        RECT 67.425 158.975 67.835 159.535 ;
        RECT 68.005 158.805 68.185 159.705 ;
        RECT 68.355 159.195 68.550 159.535 ;
        RECT 68.785 159.445 70.455 160.215 ;
        RECT 70.825 159.585 71.155 159.945 ;
        RECT 71.775 159.755 72.025 160.215 ;
        RECT 72.195 159.755 72.755 160.045 ;
        RECT 68.355 159.025 68.555 159.195 ;
        RECT 68.355 158.975 68.550 159.025 ;
        RECT 68.785 158.925 69.535 159.445 ;
        RECT 70.825 159.395 72.215 159.585 ;
        RECT 72.045 159.305 72.215 159.395 ;
        RECT 67.085 158.635 68.545 158.805 ;
        RECT 69.705 158.755 70.455 159.275 ;
        RECT 66.485 158.295 67.260 158.465 ;
        RECT 66.590 157.665 66.760 158.125 ;
        RECT 66.930 157.835 67.260 158.295 ;
        RECT 67.430 157.665 67.600 158.465 ;
        RECT 68.185 158.460 68.545 158.635 ;
        RECT 68.785 157.665 70.455 158.755 ;
        RECT 70.640 158.975 71.315 159.225 ;
        RECT 71.535 158.975 71.875 159.225 ;
        RECT 72.045 158.975 72.335 159.305 ;
        RECT 70.640 158.615 70.905 158.975 ;
        RECT 72.045 158.725 72.215 158.975 ;
        RECT 71.275 158.555 72.215 158.725 ;
        RECT 70.825 157.665 71.105 158.335 ;
        RECT 71.275 158.005 71.575 158.555 ;
        RECT 72.505 158.385 72.755 159.755 ;
        RECT 71.775 157.665 72.105 158.385 ;
        RECT 72.295 157.835 72.755 158.385 ;
        RECT 72.925 159.540 73.185 160.045 ;
        RECT 73.365 159.835 73.695 160.215 ;
        RECT 73.875 159.665 74.045 160.045 ;
        RECT 72.925 158.740 73.095 159.540 ;
        RECT 73.380 159.495 74.045 159.665 ;
        RECT 73.380 159.240 73.550 159.495 ;
        RECT 74.305 159.490 74.595 160.215 ;
        RECT 75.230 159.475 75.485 160.045 ;
        RECT 75.655 159.815 75.985 160.215 ;
        RECT 76.410 159.680 76.940 160.045 ;
        RECT 76.410 159.645 76.585 159.680 ;
        RECT 75.655 159.475 76.585 159.645 ;
        RECT 73.265 158.910 73.550 159.240 ;
        RECT 73.785 158.945 74.115 159.315 ;
        RECT 73.380 158.765 73.550 158.910 ;
        RECT 72.925 157.835 73.195 158.740 ;
        RECT 73.380 158.595 74.045 158.765 ;
        RECT 73.365 157.665 73.695 158.425 ;
        RECT 73.875 157.835 74.045 158.595 ;
        RECT 74.305 157.665 74.595 158.830 ;
        RECT 75.230 158.805 75.400 159.475 ;
        RECT 75.655 159.305 75.825 159.475 ;
        RECT 75.570 158.975 75.825 159.305 ;
        RECT 76.050 158.975 76.245 159.305 ;
        RECT 75.230 157.835 75.565 158.805 ;
        RECT 75.735 157.665 75.905 158.805 ;
        RECT 76.075 158.005 76.245 158.975 ;
        RECT 76.415 158.345 76.585 159.475 ;
        RECT 76.755 158.685 76.925 159.485 ;
        RECT 77.130 159.195 77.405 160.045 ;
        RECT 77.125 159.025 77.405 159.195 ;
        RECT 77.130 158.885 77.405 159.025 ;
        RECT 77.575 158.685 77.765 160.045 ;
        RECT 77.945 159.680 78.455 160.215 ;
        RECT 78.675 159.405 78.920 160.010 ;
        RECT 79.365 159.835 80.255 160.005 ;
        RECT 77.965 159.235 79.195 159.405 ;
        RECT 79.365 159.280 79.915 159.665 ;
        RECT 76.755 158.515 77.765 158.685 ;
        RECT 77.935 158.670 78.685 158.860 ;
        RECT 76.415 158.175 77.540 158.345 ;
        RECT 77.935 158.005 78.105 158.670 ;
        RECT 78.855 158.425 79.195 159.235 ;
        RECT 80.085 159.110 80.255 159.835 ;
        RECT 79.365 159.040 80.255 159.110 ;
        RECT 80.425 159.510 80.645 159.995 ;
        RECT 80.815 159.675 81.065 160.215 ;
        RECT 81.235 159.565 81.495 160.045 ;
        RECT 80.425 159.085 80.755 159.510 ;
        RECT 79.365 159.015 80.260 159.040 ;
        RECT 79.365 159.000 80.270 159.015 ;
        RECT 79.365 158.985 80.275 159.000 ;
        RECT 79.365 158.980 80.285 158.985 ;
        RECT 79.365 158.970 80.290 158.980 ;
        RECT 79.365 158.960 80.295 158.970 ;
        RECT 79.365 158.955 80.305 158.960 ;
        RECT 79.365 158.945 80.315 158.955 ;
        RECT 79.365 158.940 80.325 158.945 ;
        RECT 79.365 158.490 79.625 158.940 ;
        RECT 79.990 158.935 80.325 158.940 ;
        RECT 79.990 158.930 80.340 158.935 ;
        RECT 79.990 158.920 80.355 158.930 ;
        RECT 79.990 158.915 80.380 158.920 ;
        RECT 80.925 158.915 81.155 159.310 ;
        RECT 79.990 158.910 81.155 158.915 ;
        RECT 80.020 158.875 81.155 158.910 ;
        RECT 80.055 158.850 81.155 158.875 ;
        RECT 80.085 158.820 81.155 158.850 ;
        RECT 80.105 158.790 81.155 158.820 ;
        RECT 80.125 158.760 81.155 158.790 ;
        RECT 80.195 158.750 81.155 158.760 ;
        RECT 80.220 158.740 81.155 158.750 ;
        RECT 80.240 158.725 81.155 158.740 ;
        RECT 80.260 158.710 81.155 158.725 ;
        RECT 80.265 158.700 81.050 158.710 ;
        RECT 80.280 158.665 81.050 158.700 ;
        RECT 76.075 157.835 78.105 158.005 ;
        RECT 78.275 157.665 78.445 158.425 ;
        RECT 78.680 158.015 79.195 158.425 ;
        RECT 79.795 158.345 80.125 158.590 ;
        RECT 80.295 158.415 81.050 158.665 ;
        RECT 81.325 158.535 81.495 159.565 ;
        RECT 81.705 159.395 81.935 160.215 ;
        RECT 82.105 159.415 82.435 160.045 ;
        RECT 81.685 158.975 82.015 159.225 ;
        RECT 82.185 158.815 82.435 159.415 ;
        RECT 82.605 159.395 82.815 160.215 ;
        RECT 83.045 159.465 84.255 160.215 ;
        RECT 84.625 159.585 84.955 159.945 ;
        RECT 85.575 159.755 85.825 160.215 ;
        RECT 85.995 159.755 86.555 160.045 ;
        RECT 83.045 158.925 83.565 159.465 ;
        RECT 84.625 159.395 86.015 159.585 ;
        RECT 85.845 159.305 86.015 159.395 ;
        RECT 79.795 158.320 79.980 158.345 ;
        RECT 79.365 158.220 79.980 158.320 ;
        RECT 79.365 157.665 79.970 158.220 ;
        RECT 80.145 157.835 80.625 158.175 ;
        RECT 80.795 157.665 81.050 158.210 ;
        RECT 81.220 157.835 81.495 158.535 ;
        RECT 81.705 157.665 81.935 158.805 ;
        RECT 82.105 157.835 82.435 158.815 ;
        RECT 82.605 157.665 82.815 158.805 ;
        RECT 83.735 158.755 84.255 159.295 ;
        RECT 83.045 157.665 84.255 158.755 ;
        RECT 84.440 158.975 85.115 159.225 ;
        RECT 85.335 158.975 85.675 159.225 ;
        RECT 85.845 158.975 86.135 159.305 ;
        RECT 84.440 158.615 84.705 158.975 ;
        RECT 85.845 158.725 86.015 158.975 ;
        RECT 85.075 158.555 86.015 158.725 ;
        RECT 84.625 157.665 84.905 158.335 ;
        RECT 85.075 158.005 85.375 158.555 ;
        RECT 86.305 158.385 86.555 159.755 ;
        RECT 86.815 159.665 86.985 159.955 ;
        RECT 87.155 159.835 87.485 160.215 ;
        RECT 86.815 159.495 87.480 159.665 ;
        RECT 86.730 158.675 87.080 159.325 ;
        RECT 87.250 158.505 87.480 159.495 ;
        RECT 85.575 157.665 85.905 158.385 ;
        RECT 86.095 157.835 86.555 158.385 ;
        RECT 86.815 158.335 87.480 158.505 ;
        RECT 86.815 157.835 86.985 158.335 ;
        RECT 87.155 157.665 87.485 158.165 ;
        RECT 87.655 157.835 87.840 159.955 ;
        RECT 88.095 159.755 88.345 160.215 ;
        RECT 88.515 159.765 88.850 159.935 ;
        RECT 89.045 159.765 89.720 159.935 ;
        RECT 88.515 159.625 88.685 159.765 ;
        RECT 88.010 158.635 88.290 159.585 ;
        RECT 88.460 159.495 88.685 159.625 ;
        RECT 88.460 158.390 88.630 159.495 ;
        RECT 88.855 159.345 89.380 159.565 ;
        RECT 88.800 158.580 89.040 159.175 ;
        RECT 89.210 158.645 89.380 159.345 ;
        RECT 89.550 158.985 89.720 159.765 ;
        RECT 90.040 159.715 90.410 160.215 ;
        RECT 90.590 159.765 90.995 159.935 ;
        RECT 91.165 159.765 91.950 159.935 ;
        RECT 90.590 159.535 90.760 159.765 ;
        RECT 89.930 159.235 90.760 159.535 ;
        RECT 91.145 159.265 91.610 159.595 ;
        RECT 89.930 159.205 90.130 159.235 ;
        RECT 90.250 158.985 90.420 159.055 ;
        RECT 89.550 158.815 90.420 158.985 ;
        RECT 89.910 158.725 90.420 158.815 ;
        RECT 88.460 158.260 88.765 158.390 ;
        RECT 89.210 158.280 89.740 158.645 ;
        RECT 88.080 157.665 88.345 158.125 ;
        RECT 88.515 157.835 88.765 158.260 ;
        RECT 89.910 158.110 90.080 158.725 ;
        RECT 88.975 157.940 90.080 158.110 ;
        RECT 90.250 157.665 90.420 158.465 ;
        RECT 90.590 158.165 90.760 159.235 ;
        RECT 90.930 158.335 91.120 159.055 ;
        RECT 91.290 158.305 91.610 159.265 ;
        RECT 91.780 159.305 91.950 159.765 ;
        RECT 92.225 159.685 92.435 160.215 ;
        RECT 92.695 159.475 93.025 160.000 ;
        RECT 93.195 159.605 93.365 160.215 ;
        RECT 93.535 159.560 93.865 159.995 ;
        RECT 93.535 159.475 93.915 159.560 ;
        RECT 92.825 159.305 93.025 159.475 ;
        RECT 93.690 159.435 93.915 159.475 ;
        RECT 91.780 158.975 92.655 159.305 ;
        RECT 92.825 158.975 93.575 159.305 ;
        RECT 90.590 157.835 90.840 158.165 ;
        RECT 91.780 158.135 91.950 158.975 ;
        RECT 92.825 158.770 93.015 158.975 ;
        RECT 93.745 158.855 93.915 159.435 ;
        RECT 93.700 158.805 93.915 158.855 ;
        RECT 92.120 158.395 93.015 158.770 ;
        RECT 93.525 158.725 93.915 158.805 ;
        RECT 91.065 157.965 91.950 158.135 ;
        RECT 92.130 157.665 92.445 158.165 ;
        RECT 92.675 157.835 93.015 158.395 ;
        RECT 93.185 157.665 93.355 158.675 ;
        RECT 93.525 157.880 93.855 158.725 ;
        RECT 95.015 157.845 95.275 160.035 ;
        RECT 95.535 159.845 96.205 160.215 ;
        RECT 96.385 159.665 96.695 160.035 ;
        RECT 95.465 159.465 96.695 159.665 ;
        RECT 95.465 158.795 95.755 159.465 ;
        RECT 96.875 159.285 97.105 159.925 ;
        RECT 97.285 159.485 97.575 160.215 ;
        RECT 97.765 159.445 99.435 160.215 ;
        RECT 100.065 159.490 100.355 160.215 ;
        RECT 95.935 158.975 96.400 159.285 ;
        RECT 96.580 158.975 97.105 159.285 ;
        RECT 97.285 158.975 97.585 159.305 ;
        RECT 97.765 158.925 98.515 159.445 ;
        RECT 100.985 159.415 101.295 160.215 ;
        RECT 101.500 159.415 102.195 160.045 ;
        RECT 102.365 159.445 104.035 160.215 ;
        RECT 95.465 158.575 96.235 158.795 ;
        RECT 95.445 157.665 95.785 158.395 ;
        RECT 95.965 157.845 96.235 158.575 ;
        RECT 96.415 158.555 97.575 158.795 ;
        RECT 98.685 158.755 99.435 159.275 ;
        RECT 100.995 158.975 101.330 159.245 ;
        RECT 96.415 157.845 96.645 158.555 ;
        RECT 96.815 157.665 97.145 158.375 ;
        RECT 97.315 157.845 97.575 158.555 ;
        RECT 97.765 157.665 99.435 158.755 ;
        RECT 100.065 157.665 100.355 158.830 ;
        RECT 101.500 158.815 101.670 159.415 ;
        RECT 101.840 158.975 102.175 159.225 ;
        RECT 102.365 158.925 103.115 159.445 ;
        RECT 104.670 159.395 104.945 160.215 ;
        RECT 105.115 159.575 105.445 160.045 ;
        RECT 105.615 159.745 105.785 160.215 ;
        RECT 105.955 159.575 106.285 160.045 ;
        RECT 106.455 159.745 106.745 160.215 ;
        RECT 105.115 159.565 106.285 159.575 ;
        RECT 106.965 159.715 107.225 160.045 ;
        RECT 107.395 159.855 107.725 160.215 ;
        RECT 107.980 159.835 109.280 160.045 ;
        RECT 106.965 159.705 107.195 159.715 ;
        RECT 105.115 159.395 106.715 159.565 ;
        RECT 100.985 157.665 101.265 158.805 ;
        RECT 101.435 157.835 101.765 158.815 ;
        RECT 101.935 157.665 102.195 158.805 ;
        RECT 103.285 158.755 104.035 159.275 ;
        RECT 104.670 159.025 105.390 159.225 ;
        RECT 105.560 159.025 106.330 159.225 ;
        RECT 106.500 158.855 106.715 159.395 ;
        RECT 102.365 157.665 104.035 158.755 ;
        RECT 104.670 158.635 105.785 158.845 ;
        RECT 104.670 157.835 104.945 158.635 ;
        RECT 105.115 157.665 105.445 158.465 ;
        RECT 105.615 158.005 105.785 158.635 ;
        RECT 105.955 158.685 106.735 158.855 ;
        RECT 105.955 158.635 106.715 158.685 ;
        RECT 105.955 158.175 106.285 158.635 ;
        RECT 106.965 158.515 107.135 159.705 ;
        RECT 107.980 159.685 108.150 159.835 ;
        RECT 107.395 159.560 108.150 159.685 ;
        RECT 107.305 159.515 108.150 159.560 ;
        RECT 107.305 159.395 107.575 159.515 ;
        RECT 107.305 158.820 107.475 159.395 ;
        RECT 107.705 158.955 108.115 159.260 ;
        RECT 108.405 159.225 108.615 159.625 ;
        RECT 108.285 159.015 108.615 159.225 ;
        RECT 108.860 159.225 109.080 159.625 ;
        RECT 109.555 159.450 110.010 160.215 ;
        RECT 110.185 159.445 111.855 160.215 ;
        RECT 112.030 159.450 112.485 160.215 ;
        RECT 112.760 159.835 114.060 160.045 ;
        RECT 114.315 159.855 114.645 160.215 ;
        RECT 113.890 159.685 114.060 159.835 ;
        RECT 114.815 159.715 115.075 160.045 ;
        RECT 114.845 159.705 115.075 159.715 ;
        RECT 108.860 159.015 109.335 159.225 ;
        RECT 109.525 159.025 110.015 159.225 ;
        RECT 110.185 158.925 110.935 159.445 ;
        RECT 107.305 158.785 107.505 158.820 ;
        RECT 108.835 158.785 110.010 158.845 ;
        RECT 107.305 158.675 110.010 158.785 ;
        RECT 111.105 158.755 111.855 159.275 ;
        RECT 112.960 159.225 113.180 159.625 ;
        RECT 112.025 159.025 112.515 159.225 ;
        RECT 112.705 159.015 113.180 159.225 ;
        RECT 113.425 159.225 113.635 159.625 ;
        RECT 113.890 159.560 114.645 159.685 ;
        RECT 113.890 159.515 114.735 159.560 ;
        RECT 114.465 159.395 114.735 159.515 ;
        RECT 113.425 159.015 113.755 159.225 ;
        RECT 113.925 158.955 114.335 159.260 ;
        RECT 107.365 158.615 109.165 158.675 ;
        RECT 108.835 158.585 109.165 158.615 ;
        RECT 106.455 158.005 106.755 158.465 ;
        RECT 105.615 157.835 106.755 158.005 ;
        RECT 106.965 157.835 107.225 158.515 ;
        RECT 107.395 157.665 107.645 158.445 ;
        RECT 107.895 158.415 108.730 158.425 ;
        RECT 109.320 158.415 109.505 158.505 ;
        RECT 107.895 158.215 109.505 158.415 ;
        RECT 107.895 157.835 108.145 158.215 ;
        RECT 109.275 158.175 109.505 158.215 ;
        RECT 109.755 158.055 110.010 158.675 ;
        RECT 108.315 157.665 108.670 158.045 ;
        RECT 109.675 157.835 110.010 158.055 ;
        RECT 110.185 157.665 111.855 158.755 ;
        RECT 112.030 158.785 113.205 158.845 ;
        RECT 114.565 158.820 114.735 159.395 ;
        RECT 114.535 158.785 114.735 158.820 ;
        RECT 112.030 158.675 114.735 158.785 ;
        RECT 112.030 158.055 112.285 158.675 ;
        RECT 112.875 158.615 114.675 158.675 ;
        RECT 112.875 158.585 113.205 158.615 ;
        RECT 114.905 158.515 115.075 159.705 ;
        RECT 115.335 159.665 115.505 159.955 ;
        RECT 115.675 159.835 116.005 160.215 ;
        RECT 115.335 159.495 116.000 159.665 ;
        RECT 115.250 158.675 115.600 159.325 ;
        RECT 112.535 158.415 112.720 158.505 ;
        RECT 113.310 158.415 114.145 158.425 ;
        RECT 112.535 158.215 114.145 158.415 ;
        RECT 112.535 158.175 112.765 158.215 ;
        RECT 112.030 157.835 112.365 158.055 ;
        RECT 113.370 157.665 113.725 158.045 ;
        RECT 113.895 157.835 114.145 158.215 ;
        RECT 114.395 157.665 114.645 158.445 ;
        RECT 114.815 157.835 115.075 158.515 ;
        RECT 115.770 158.505 116.000 159.495 ;
        RECT 115.335 158.335 116.000 158.505 ;
        RECT 115.335 157.835 115.505 158.335 ;
        RECT 115.675 157.665 116.005 158.165 ;
        RECT 116.175 157.835 116.360 159.955 ;
        RECT 116.615 159.755 116.865 160.215 ;
        RECT 117.035 159.765 117.370 159.935 ;
        RECT 117.565 159.765 118.240 159.935 ;
        RECT 117.035 159.625 117.205 159.765 ;
        RECT 116.530 158.635 116.810 159.585 ;
        RECT 116.980 159.495 117.205 159.625 ;
        RECT 116.980 158.390 117.150 159.495 ;
        RECT 117.375 159.345 117.900 159.565 ;
        RECT 117.320 158.580 117.560 159.175 ;
        RECT 117.730 158.645 117.900 159.345 ;
        RECT 118.070 158.985 118.240 159.765 ;
        RECT 118.560 159.715 118.930 160.215 ;
        RECT 119.110 159.765 119.515 159.935 ;
        RECT 119.685 159.765 120.470 159.935 ;
        RECT 119.110 159.535 119.280 159.765 ;
        RECT 118.450 159.235 119.280 159.535 ;
        RECT 119.665 159.265 120.130 159.595 ;
        RECT 118.450 159.205 118.650 159.235 ;
        RECT 118.770 158.985 118.940 159.055 ;
        RECT 118.070 158.815 118.940 158.985 ;
        RECT 118.430 158.725 118.940 158.815 ;
        RECT 116.980 158.260 117.285 158.390 ;
        RECT 117.730 158.280 118.260 158.645 ;
        RECT 116.600 157.665 116.865 158.125 ;
        RECT 117.035 157.835 117.285 158.260 ;
        RECT 118.430 158.110 118.600 158.725 ;
        RECT 117.495 157.940 118.600 158.110 ;
        RECT 118.770 157.665 118.940 158.465 ;
        RECT 119.110 158.165 119.280 159.235 ;
        RECT 119.450 158.335 119.640 159.055 ;
        RECT 119.810 158.305 120.130 159.265 ;
        RECT 120.300 159.305 120.470 159.765 ;
        RECT 120.745 159.685 120.955 160.215 ;
        RECT 121.215 159.475 121.545 160.000 ;
        RECT 121.715 159.605 121.885 160.215 ;
        RECT 122.055 159.560 122.385 159.995 ;
        RECT 122.630 159.565 122.940 160.035 ;
        RECT 123.110 159.735 123.845 160.215 ;
        RECT 124.015 159.645 124.185 159.995 ;
        RECT 124.355 159.815 124.735 160.215 ;
        RECT 122.055 159.475 122.435 159.560 ;
        RECT 121.345 159.305 121.545 159.475 ;
        RECT 122.210 159.435 122.435 159.475 ;
        RECT 120.300 158.975 121.175 159.305 ;
        RECT 121.345 158.975 122.095 159.305 ;
        RECT 119.110 157.835 119.360 158.165 ;
        RECT 120.300 158.135 120.470 158.975 ;
        RECT 121.345 158.770 121.535 158.975 ;
        RECT 122.265 158.855 122.435 159.435 ;
        RECT 122.630 159.395 123.365 159.565 ;
        RECT 124.015 159.475 124.755 159.645 ;
        RECT 124.925 159.540 125.195 159.885 ;
        RECT 123.115 159.305 123.365 159.395 ;
        RECT 124.585 159.305 124.755 159.475 ;
        RECT 122.610 158.975 122.945 159.225 ;
        RECT 123.115 158.975 123.855 159.305 ;
        RECT 124.585 158.975 124.815 159.305 ;
        RECT 122.220 158.805 122.435 158.855 ;
        RECT 120.640 158.395 121.535 158.770 ;
        RECT 122.045 158.725 122.435 158.805 ;
        RECT 119.585 157.965 120.470 158.135 ;
        RECT 120.650 157.665 120.965 158.165 ;
        RECT 121.195 157.835 121.535 158.395 ;
        RECT 121.705 157.665 121.875 158.675 ;
        RECT 122.045 157.880 122.375 158.725 ;
        RECT 122.610 157.665 122.865 158.805 ;
        RECT 123.115 158.415 123.285 158.975 ;
        RECT 124.585 158.805 124.755 158.975 ;
        RECT 125.025 158.805 125.195 159.540 ;
        RECT 125.825 159.490 126.115 160.215 ;
        RECT 126.305 159.525 126.545 160.045 ;
        RECT 126.715 159.720 127.110 160.215 ;
        RECT 127.675 159.885 127.845 160.030 ;
        RECT 127.470 159.690 127.845 159.885 ;
        RECT 123.510 158.635 124.755 158.805 ;
        RECT 123.510 158.385 123.930 158.635 ;
        RECT 123.060 157.885 124.255 158.215 ;
        RECT 124.435 157.665 124.715 158.465 ;
        RECT 124.925 157.835 125.195 158.805 ;
        RECT 125.825 157.665 126.115 158.830 ;
        RECT 126.305 158.720 126.480 159.525 ;
        RECT 127.470 159.355 127.640 159.690 ;
        RECT 128.125 159.645 128.365 160.020 ;
        RECT 128.535 159.710 128.870 160.215 ;
        RECT 128.125 159.495 128.345 159.645 ;
        RECT 126.655 158.995 127.640 159.355 ;
        RECT 127.810 159.165 128.345 159.495 ;
        RECT 126.655 158.975 127.940 158.995 ;
        RECT 127.080 158.825 127.940 158.975 ;
        RECT 126.305 157.935 126.610 158.720 ;
        RECT 126.785 158.345 127.480 158.655 ;
        RECT 126.790 157.665 127.475 158.135 ;
        RECT 127.655 157.880 127.940 158.825 ;
        RECT 128.110 158.515 128.345 159.165 ;
        RECT 128.515 158.685 128.815 159.535 ;
        RECT 129.065 159.525 129.305 160.045 ;
        RECT 129.475 159.720 129.870 160.215 ;
        RECT 130.435 159.885 130.605 160.030 ;
        RECT 130.230 159.690 130.605 159.885 ;
        RECT 129.065 158.720 129.240 159.525 ;
        RECT 130.230 159.355 130.400 159.690 ;
        RECT 130.885 159.645 131.125 160.020 ;
        RECT 131.295 159.710 131.630 160.215 ;
        RECT 130.885 159.495 131.105 159.645 ;
        RECT 129.415 158.995 130.400 159.355 ;
        RECT 130.570 159.165 131.105 159.495 ;
        RECT 129.415 158.975 130.700 158.995 ;
        RECT 129.840 158.825 130.700 158.975 ;
        RECT 128.110 158.285 128.785 158.515 ;
        RECT 128.115 157.665 128.445 158.115 ;
        RECT 128.615 157.855 128.785 158.285 ;
        RECT 129.065 157.935 129.370 158.720 ;
        RECT 129.545 158.345 130.240 158.655 ;
        RECT 129.550 157.665 130.235 158.135 ;
        RECT 130.415 157.880 130.700 158.825 ;
        RECT 130.870 158.515 131.105 159.165 ;
        RECT 131.275 158.685 131.575 159.535 ;
        RECT 131.865 159.395 132.075 160.215 ;
        RECT 132.245 159.415 132.575 160.045 ;
        RECT 132.245 158.815 132.495 159.415 ;
        RECT 132.745 159.395 132.975 160.215 ;
        RECT 133.185 159.445 135.775 160.215 ;
        RECT 136.405 159.835 137.295 160.005 ;
        RECT 132.665 158.975 132.995 159.225 ;
        RECT 133.185 158.925 134.395 159.445 ;
        RECT 136.405 159.280 136.955 159.665 ;
        RECT 130.870 158.285 131.545 158.515 ;
        RECT 130.875 157.665 131.205 158.115 ;
        RECT 131.375 157.855 131.545 158.285 ;
        RECT 131.865 157.665 132.075 158.805 ;
        RECT 132.245 157.835 132.575 158.815 ;
        RECT 132.745 157.665 132.975 158.805 ;
        RECT 134.565 158.755 135.775 159.275 ;
        RECT 137.125 159.110 137.295 159.835 ;
        RECT 133.185 157.665 135.775 158.755 ;
        RECT 136.405 159.040 137.295 159.110 ;
        RECT 137.465 159.510 137.685 159.995 ;
        RECT 137.855 159.675 138.105 160.215 ;
        RECT 138.275 159.565 138.535 160.045 ;
        RECT 137.465 159.085 137.795 159.510 ;
        RECT 136.405 159.015 137.300 159.040 ;
        RECT 136.405 159.000 137.310 159.015 ;
        RECT 136.405 158.985 137.315 159.000 ;
        RECT 136.405 158.980 137.325 158.985 ;
        RECT 136.405 158.970 137.330 158.980 ;
        RECT 136.405 158.960 137.335 158.970 ;
        RECT 136.405 158.955 137.345 158.960 ;
        RECT 136.405 158.945 137.355 158.955 ;
        RECT 136.405 158.940 137.365 158.945 ;
        RECT 136.405 158.490 136.665 158.940 ;
        RECT 137.030 158.935 137.365 158.940 ;
        RECT 137.030 158.930 137.380 158.935 ;
        RECT 137.030 158.920 137.395 158.930 ;
        RECT 137.030 158.915 137.420 158.920 ;
        RECT 137.965 158.915 138.195 159.310 ;
        RECT 137.030 158.910 138.195 158.915 ;
        RECT 137.060 158.875 138.195 158.910 ;
        RECT 137.095 158.850 138.195 158.875 ;
        RECT 137.125 158.820 138.195 158.850 ;
        RECT 137.145 158.790 138.195 158.820 ;
        RECT 137.165 158.760 138.195 158.790 ;
        RECT 137.235 158.750 138.195 158.760 ;
        RECT 137.260 158.740 138.195 158.750 ;
        RECT 137.280 158.725 138.195 158.740 ;
        RECT 137.300 158.710 138.195 158.725 ;
        RECT 137.305 158.700 138.090 158.710 ;
        RECT 137.320 158.665 138.090 158.700 ;
        RECT 136.835 158.345 137.165 158.590 ;
        RECT 137.335 158.415 138.090 158.665 ;
        RECT 138.365 158.535 138.535 159.565 ;
        RECT 138.705 159.445 142.215 160.215 ;
        RECT 143.305 159.475 143.770 160.020 ;
        RECT 138.705 158.925 140.355 159.445 ;
        RECT 140.525 158.755 142.215 159.275 ;
        RECT 136.835 158.320 137.020 158.345 ;
        RECT 136.405 158.220 137.020 158.320 ;
        RECT 136.405 157.665 137.010 158.220 ;
        RECT 137.185 157.835 137.665 158.175 ;
        RECT 137.835 157.665 138.090 158.210 ;
        RECT 138.260 157.835 138.535 158.535 ;
        RECT 138.705 157.665 142.215 158.755 ;
        RECT 143.305 158.515 143.475 159.475 ;
        RECT 144.275 159.395 144.445 160.215 ;
        RECT 144.615 159.565 144.945 160.045 ;
        RECT 145.115 159.825 145.465 160.215 ;
        RECT 145.635 159.645 145.865 160.045 ;
        RECT 145.355 159.565 145.865 159.645 ;
        RECT 144.615 159.475 145.865 159.565 ;
        RECT 146.035 159.475 146.355 159.955 ;
        RECT 144.615 159.395 145.525 159.475 ;
        RECT 143.645 158.855 143.890 159.305 ;
        RECT 144.150 159.025 144.845 159.225 ;
        RECT 145.015 159.055 145.615 159.225 ;
        RECT 145.015 158.855 145.185 159.055 ;
        RECT 145.845 158.885 146.015 159.305 ;
        RECT 143.645 158.685 145.185 158.855 ;
        RECT 145.355 158.715 146.015 158.885 ;
        RECT 145.355 158.515 145.525 158.715 ;
        RECT 146.185 158.545 146.355 159.475 ;
        RECT 146.985 159.415 147.295 160.215 ;
        RECT 147.500 159.415 148.195 160.045 ;
        RECT 148.365 159.445 150.955 160.215 ;
        RECT 151.585 159.490 151.875 160.215 ;
        RECT 152.045 159.475 152.430 160.045 ;
        RECT 152.600 159.755 152.925 160.215 ;
        RECT 153.445 159.585 153.725 160.045 ;
        RECT 146.995 158.975 147.330 159.245 ;
        RECT 147.500 158.815 147.670 159.415 ;
        RECT 147.840 158.975 148.175 159.225 ;
        RECT 148.365 158.925 149.575 159.445 ;
        RECT 143.305 158.345 145.525 158.515 ;
        RECT 145.695 158.345 146.355 158.545 ;
        RECT 143.305 157.665 143.605 158.175 ;
        RECT 143.775 157.835 144.105 158.345 ;
        RECT 145.695 158.175 145.865 158.345 ;
        RECT 144.275 157.665 144.905 158.175 ;
        RECT 145.485 158.005 145.865 158.175 ;
        RECT 146.035 157.665 146.335 158.175 ;
        RECT 146.985 157.665 147.265 158.805 ;
        RECT 147.435 157.835 147.765 158.815 ;
        RECT 147.935 157.665 148.195 158.805 ;
        RECT 149.745 158.755 150.955 159.275 ;
        RECT 148.365 157.665 150.955 158.755 ;
        RECT 151.585 157.665 151.875 158.830 ;
        RECT 152.045 158.805 152.325 159.475 ;
        RECT 152.600 159.415 153.725 159.585 ;
        RECT 152.600 159.305 153.050 159.415 ;
        RECT 152.495 158.975 153.050 159.305 ;
        RECT 153.915 159.245 154.315 160.045 ;
        RECT 154.715 159.755 154.985 160.215 ;
        RECT 155.155 159.585 155.440 160.045 ;
        RECT 152.045 157.835 152.430 158.805 ;
        RECT 152.600 158.515 153.050 158.975 ;
        RECT 153.220 158.685 154.315 159.245 ;
        RECT 152.600 158.295 153.725 158.515 ;
        RECT 152.600 157.665 152.925 158.125 ;
        RECT 153.445 157.835 153.725 158.295 ;
        RECT 153.915 157.835 154.315 158.685 ;
        RECT 154.485 159.415 155.440 159.585 ;
        RECT 155.725 159.465 156.935 160.215 ;
        RECT 154.485 158.515 154.695 159.415 ;
        RECT 154.865 158.685 155.555 159.245 ;
        RECT 155.725 158.755 156.245 159.295 ;
        RECT 156.415 158.925 156.935 159.465 ;
        RECT 154.485 158.295 155.440 158.515 ;
        RECT 154.715 157.665 154.985 158.125 ;
        RECT 155.155 157.835 155.440 158.295 ;
        RECT 155.725 157.665 156.935 158.755 ;
        RECT 22.700 157.495 157.020 157.665 ;
        RECT 22.785 156.405 23.995 157.495 ;
        RECT 24.165 156.405 27.675 157.495 ;
        RECT 22.785 155.695 23.305 156.235 ;
        RECT 23.475 155.865 23.995 156.405 ;
        RECT 24.165 155.715 25.815 156.235 ;
        RECT 25.985 155.885 27.675 156.405 ;
        RECT 28.305 156.625 28.580 157.325 ;
        RECT 28.750 156.950 29.005 157.495 ;
        RECT 29.175 156.985 29.655 157.325 ;
        RECT 29.830 156.940 30.435 157.495 ;
        RECT 29.820 156.840 30.435 156.940 ;
        RECT 29.820 156.815 30.005 156.840 ;
        RECT 22.785 154.945 23.995 155.695 ;
        RECT 24.165 154.945 27.675 155.715 ;
        RECT 28.305 155.595 28.475 156.625 ;
        RECT 28.750 156.495 29.505 156.745 ;
        RECT 29.675 156.570 30.005 156.815 ;
        RECT 28.750 156.460 29.520 156.495 ;
        RECT 28.750 156.450 29.535 156.460 ;
        RECT 28.645 156.435 29.540 156.450 ;
        RECT 28.645 156.420 29.560 156.435 ;
        RECT 28.645 156.410 29.580 156.420 ;
        RECT 28.645 156.400 29.605 156.410 ;
        RECT 28.645 156.370 29.675 156.400 ;
        RECT 28.645 156.340 29.695 156.370 ;
        RECT 28.645 156.310 29.715 156.340 ;
        RECT 28.645 156.285 29.745 156.310 ;
        RECT 28.645 156.250 29.780 156.285 ;
        RECT 28.645 156.245 29.810 156.250 ;
        RECT 28.645 155.850 28.875 156.245 ;
        RECT 29.420 156.240 29.810 156.245 ;
        RECT 29.445 156.230 29.810 156.240 ;
        RECT 29.460 156.225 29.810 156.230 ;
        RECT 29.475 156.220 29.810 156.225 ;
        RECT 30.175 156.220 30.435 156.670 ;
        RECT 30.605 156.355 30.865 157.495 ;
        RECT 31.035 156.345 31.365 157.325 ;
        RECT 31.535 156.355 31.815 157.495 ;
        RECT 31.985 156.355 32.265 157.495 ;
        RECT 32.435 156.345 32.765 157.325 ;
        RECT 32.935 156.355 33.195 157.495 ;
        RECT 33.365 156.355 33.625 157.495 ;
        RECT 33.795 156.345 34.125 157.325 ;
        RECT 34.295 156.355 34.575 157.495 ;
        RECT 29.475 156.215 30.435 156.220 ;
        RECT 29.485 156.205 30.435 156.215 ;
        RECT 29.495 156.200 30.435 156.205 ;
        RECT 29.505 156.190 30.435 156.200 ;
        RECT 29.510 156.180 30.435 156.190 ;
        RECT 29.515 156.175 30.435 156.180 ;
        RECT 29.525 156.160 30.435 156.175 ;
        RECT 29.530 156.145 30.435 156.160 ;
        RECT 29.540 156.120 30.435 156.145 ;
        RECT 29.045 155.650 29.375 156.075 ;
        RECT 28.305 155.115 28.565 155.595 ;
        RECT 28.735 154.945 28.985 155.485 ;
        RECT 29.155 155.165 29.375 155.650 ;
        RECT 29.545 156.050 30.435 156.120 ;
        RECT 29.545 155.325 29.715 156.050 ;
        RECT 30.625 155.935 30.960 156.185 ;
        RECT 29.885 155.495 30.435 155.880 ;
        RECT 31.130 155.745 31.300 156.345 ;
        RECT 31.470 155.915 31.805 156.185 ;
        RECT 31.995 155.915 32.330 156.185 ;
        RECT 32.500 155.745 32.670 156.345 ;
        RECT 33.885 156.305 34.060 156.345 ;
        RECT 35.665 156.330 35.955 157.495 ;
        RECT 36.125 156.405 37.795 157.495 ;
        RECT 32.840 155.935 33.175 156.185 ;
        RECT 33.385 155.935 33.720 156.185 ;
        RECT 33.890 155.745 34.060 156.305 ;
        RECT 34.230 155.915 34.565 156.185 ;
        RECT 29.545 155.155 30.435 155.325 ;
        RECT 30.605 155.115 31.300 155.745 ;
        RECT 31.505 154.945 31.815 155.745 ;
        RECT 31.985 154.945 32.295 155.745 ;
        RECT 32.500 155.115 33.195 155.745 ;
        RECT 33.365 155.115 34.060 155.745 ;
        RECT 34.265 154.945 34.575 155.745 ;
        RECT 36.125 155.715 36.875 156.235 ;
        RECT 37.045 155.885 37.795 156.405 ;
        RECT 37.970 156.355 38.225 157.495 ;
        RECT 38.420 156.945 39.615 157.275 ;
        RECT 38.475 156.185 38.645 156.745 ;
        RECT 38.870 156.525 39.290 156.775 ;
        RECT 39.795 156.695 40.075 157.495 ;
        RECT 38.870 156.355 40.115 156.525 ;
        RECT 40.285 156.355 40.555 157.325 ;
        RECT 41.645 156.355 41.925 157.495 ;
        RECT 39.945 156.185 40.115 156.355 ;
        RECT 40.325 156.305 40.555 156.355 ;
        RECT 42.095 156.345 42.425 157.325 ;
        RECT 42.595 156.355 42.855 157.495 ;
        RECT 37.970 155.935 38.305 156.185 ;
        RECT 38.475 155.855 39.215 156.185 ;
        RECT 39.945 155.855 40.175 156.185 ;
        RECT 38.475 155.765 38.725 155.855 ;
        RECT 35.665 154.945 35.955 155.670 ;
        RECT 36.125 154.945 37.795 155.715 ;
        RECT 37.990 155.595 38.725 155.765 ;
        RECT 39.945 155.685 40.115 155.855 ;
        RECT 37.990 155.125 38.300 155.595 ;
        RECT 39.375 155.515 40.115 155.685 ;
        RECT 40.385 155.620 40.555 156.305 ;
        RECT 41.655 155.915 41.990 156.185 ;
        RECT 42.160 155.745 42.330 156.345 ;
        RECT 42.500 155.935 42.835 156.185 ;
        RECT 43.485 155.890 43.765 157.325 ;
        RECT 43.935 156.720 44.645 157.495 ;
        RECT 44.815 156.550 45.145 157.325 ;
        RECT 43.995 156.335 45.145 156.550 ;
        RECT 38.470 154.945 39.205 155.425 ;
        RECT 39.375 155.165 39.545 155.515 ;
        RECT 39.715 154.945 40.095 155.345 ;
        RECT 40.285 155.275 40.555 155.620 ;
        RECT 41.645 154.945 41.955 155.745 ;
        RECT 42.160 155.115 42.855 155.745 ;
        RECT 43.485 155.115 43.825 155.890 ;
        RECT 43.995 155.765 44.280 156.335 ;
        RECT 44.465 155.935 44.935 156.165 ;
        RECT 45.340 156.135 45.555 157.250 ;
        RECT 45.735 156.775 46.065 157.495 ;
        RECT 45.845 156.135 46.075 156.475 ;
        RECT 46.245 156.405 47.915 157.495 ;
        RECT 48.175 156.825 48.345 157.325 ;
        RECT 48.515 156.995 48.845 157.495 ;
        RECT 48.175 156.655 48.840 156.825 ;
        RECT 45.105 155.955 45.555 156.135 ;
        RECT 45.105 155.935 45.435 155.955 ;
        RECT 45.745 155.935 46.075 156.135 ;
        RECT 43.995 155.575 44.705 155.765 ;
        RECT 44.405 155.435 44.705 155.575 ;
        RECT 44.895 155.575 46.075 155.765 ;
        RECT 44.895 155.495 45.225 155.575 ;
        RECT 44.405 155.425 44.720 155.435 ;
        RECT 44.405 155.415 44.730 155.425 ;
        RECT 44.405 155.410 44.740 155.415 ;
        RECT 43.995 154.945 44.165 155.405 ;
        RECT 44.405 155.400 44.745 155.410 ;
        RECT 44.405 155.395 44.750 155.400 ;
        RECT 44.405 155.385 44.755 155.395 ;
        RECT 44.405 155.380 44.760 155.385 ;
        RECT 44.405 155.115 44.765 155.380 ;
        RECT 45.395 154.945 45.565 155.405 ;
        RECT 45.735 155.115 46.075 155.575 ;
        RECT 46.245 155.715 46.995 156.235 ;
        RECT 47.165 155.885 47.915 156.405 ;
        RECT 48.090 155.835 48.440 156.485 ;
        RECT 46.245 154.945 47.915 155.715 ;
        RECT 48.610 155.665 48.840 156.655 ;
        RECT 48.175 155.495 48.840 155.665 ;
        RECT 48.175 155.205 48.345 155.495 ;
        RECT 48.515 154.945 48.845 155.325 ;
        RECT 49.015 155.205 49.200 157.325 ;
        RECT 49.440 157.035 49.705 157.495 ;
        RECT 49.875 156.900 50.125 157.325 ;
        RECT 50.335 157.050 51.440 157.220 ;
        RECT 49.820 156.770 50.125 156.900 ;
        RECT 49.370 155.575 49.650 156.525 ;
        RECT 49.820 155.665 49.990 156.770 ;
        RECT 50.160 155.985 50.400 156.580 ;
        RECT 50.570 156.515 51.100 156.880 ;
        RECT 50.570 155.815 50.740 156.515 ;
        RECT 51.270 156.435 51.440 157.050 ;
        RECT 51.610 156.695 51.780 157.495 ;
        RECT 51.950 156.995 52.200 157.325 ;
        RECT 52.425 157.025 53.310 157.195 ;
        RECT 51.270 156.345 51.780 156.435 ;
        RECT 49.820 155.535 50.045 155.665 ;
        RECT 50.215 155.595 50.740 155.815 ;
        RECT 50.910 156.175 51.780 156.345 ;
        RECT 49.455 154.945 49.705 155.405 ;
        RECT 49.875 155.395 50.045 155.535 ;
        RECT 50.910 155.395 51.080 156.175 ;
        RECT 51.610 156.105 51.780 156.175 ;
        RECT 51.290 155.925 51.490 155.955 ;
        RECT 51.950 155.925 52.120 156.995 ;
        RECT 52.290 156.105 52.480 156.825 ;
        RECT 51.290 155.625 52.120 155.925 ;
        RECT 52.650 155.895 52.970 156.855 ;
        RECT 49.875 155.225 50.210 155.395 ;
        RECT 50.405 155.225 51.080 155.395 ;
        RECT 51.400 154.945 51.770 155.445 ;
        RECT 51.950 155.395 52.120 155.625 ;
        RECT 52.505 155.565 52.970 155.895 ;
        RECT 53.140 156.185 53.310 157.025 ;
        RECT 53.490 156.995 53.805 157.495 ;
        RECT 54.035 156.765 54.375 157.325 ;
        RECT 53.480 156.390 54.375 156.765 ;
        RECT 54.545 156.485 54.715 157.495 ;
        RECT 54.185 156.185 54.375 156.390 ;
        RECT 54.885 156.435 55.215 157.280 ;
        RECT 54.885 156.355 55.275 156.435 ;
        RECT 55.445 156.405 57.115 157.495 ;
        RECT 55.060 156.305 55.275 156.355 ;
        RECT 53.140 155.855 54.015 156.185 ;
        RECT 54.185 155.855 54.935 156.185 ;
        RECT 53.140 155.395 53.310 155.855 ;
        RECT 54.185 155.685 54.385 155.855 ;
        RECT 55.105 155.725 55.275 156.305 ;
        RECT 55.050 155.685 55.275 155.725 ;
        RECT 51.950 155.225 52.355 155.395 ;
        RECT 52.525 155.225 53.310 155.395 ;
        RECT 53.585 154.945 53.795 155.475 ;
        RECT 54.055 155.160 54.385 155.685 ;
        RECT 54.895 155.600 55.275 155.685 ;
        RECT 55.445 155.715 56.195 156.235 ;
        RECT 56.365 155.885 57.115 156.405 ;
        RECT 57.305 156.605 57.565 157.315 ;
        RECT 57.735 156.785 58.065 157.495 ;
        RECT 58.235 156.605 58.465 157.315 ;
        RECT 57.305 156.365 58.465 156.605 ;
        RECT 58.645 156.585 58.915 157.315 ;
        RECT 59.095 156.765 59.435 157.495 ;
        RECT 58.645 156.365 59.415 156.585 ;
        RECT 57.295 155.855 57.595 156.185 ;
        RECT 57.775 155.875 58.300 156.185 ;
        RECT 58.480 155.875 58.945 156.185 ;
        RECT 54.555 154.945 54.725 155.555 ;
        RECT 54.895 155.165 55.225 155.600 ;
        RECT 55.445 154.945 57.115 155.715 ;
        RECT 57.305 154.945 57.595 155.675 ;
        RECT 57.775 155.235 58.005 155.875 ;
        RECT 59.125 155.695 59.415 156.365 ;
        RECT 58.185 155.495 59.415 155.695 ;
        RECT 58.185 155.125 58.495 155.495 ;
        RECT 58.675 154.945 59.345 155.315 ;
        RECT 59.605 155.125 59.865 157.315 ;
        RECT 60.045 156.405 61.255 157.495 ;
        RECT 60.045 155.695 60.565 156.235 ;
        RECT 60.735 155.865 61.255 156.405 ;
        RECT 61.425 156.330 61.715 157.495 ;
        RECT 61.945 156.435 62.275 157.280 ;
        RECT 62.445 156.485 62.615 157.495 ;
        RECT 62.785 156.765 63.125 157.325 ;
        RECT 63.355 156.995 63.670 157.495 ;
        RECT 63.850 157.025 64.735 157.195 ;
        RECT 61.885 156.355 62.275 156.435 ;
        RECT 62.785 156.390 63.680 156.765 ;
        RECT 61.885 156.305 62.100 156.355 ;
        RECT 61.885 155.725 62.055 156.305 ;
        RECT 62.785 156.185 62.975 156.390 ;
        RECT 63.850 156.185 64.020 157.025 ;
        RECT 64.960 156.995 65.210 157.325 ;
        RECT 62.225 155.855 62.975 156.185 ;
        RECT 63.145 155.855 64.020 156.185 ;
        RECT 60.045 154.945 61.255 155.695 ;
        RECT 61.885 155.685 62.110 155.725 ;
        RECT 62.775 155.685 62.975 155.855 ;
        RECT 61.425 154.945 61.715 155.670 ;
        RECT 61.885 155.600 62.265 155.685 ;
        RECT 61.935 155.165 62.265 155.600 ;
        RECT 62.435 154.945 62.605 155.555 ;
        RECT 62.775 155.160 63.105 155.685 ;
        RECT 63.365 154.945 63.575 155.475 ;
        RECT 63.850 155.395 64.020 155.855 ;
        RECT 64.190 155.895 64.510 156.855 ;
        RECT 64.680 156.105 64.870 156.825 ;
        RECT 65.040 155.925 65.210 156.995 ;
        RECT 65.380 156.695 65.550 157.495 ;
        RECT 65.720 157.050 66.825 157.220 ;
        RECT 65.720 156.435 65.890 157.050 ;
        RECT 67.035 156.900 67.285 157.325 ;
        RECT 67.455 157.035 67.720 157.495 ;
        RECT 66.060 156.515 66.590 156.880 ;
        RECT 67.035 156.770 67.340 156.900 ;
        RECT 65.380 156.345 65.890 156.435 ;
        RECT 65.380 156.175 66.250 156.345 ;
        RECT 65.380 156.105 65.550 156.175 ;
        RECT 65.670 155.925 65.870 155.955 ;
        RECT 64.190 155.565 64.655 155.895 ;
        RECT 65.040 155.625 65.870 155.925 ;
        RECT 65.040 155.395 65.210 155.625 ;
        RECT 63.850 155.225 64.635 155.395 ;
        RECT 64.805 155.225 65.210 155.395 ;
        RECT 65.390 154.945 65.760 155.445 ;
        RECT 66.080 155.395 66.250 156.175 ;
        RECT 66.420 155.815 66.590 156.515 ;
        RECT 66.760 155.985 67.000 156.580 ;
        RECT 66.420 155.595 66.945 155.815 ;
        RECT 67.170 155.665 67.340 156.770 ;
        RECT 67.115 155.535 67.340 155.665 ;
        RECT 67.510 155.575 67.790 156.525 ;
        RECT 67.115 155.395 67.285 155.535 ;
        RECT 66.080 155.225 66.755 155.395 ;
        RECT 66.950 155.225 67.285 155.395 ;
        RECT 67.455 154.945 67.705 155.405 ;
        RECT 67.960 155.205 68.145 157.325 ;
        RECT 68.315 156.995 68.645 157.495 ;
        RECT 68.815 156.825 68.985 157.325 ;
        RECT 68.320 156.655 68.985 156.825 ;
        RECT 69.795 156.825 69.965 157.325 ;
        RECT 70.135 156.995 70.465 157.495 ;
        RECT 69.795 156.655 70.460 156.825 ;
        RECT 68.320 155.665 68.550 156.655 ;
        RECT 68.720 155.835 69.070 156.485 ;
        RECT 69.710 155.835 70.060 156.485 ;
        RECT 70.230 155.665 70.460 156.655 ;
        RECT 68.320 155.495 68.985 155.665 ;
        RECT 68.315 154.945 68.645 155.325 ;
        RECT 68.815 155.205 68.985 155.495 ;
        RECT 69.795 155.495 70.460 155.665 ;
        RECT 69.795 155.205 69.965 155.495 ;
        RECT 70.135 154.945 70.465 155.325 ;
        RECT 70.635 155.205 70.820 157.325 ;
        RECT 71.060 157.035 71.325 157.495 ;
        RECT 71.495 156.900 71.745 157.325 ;
        RECT 71.955 157.050 73.060 157.220 ;
        RECT 71.440 156.770 71.745 156.900 ;
        RECT 70.990 155.575 71.270 156.525 ;
        RECT 71.440 155.665 71.610 156.770 ;
        RECT 71.780 155.985 72.020 156.580 ;
        RECT 72.190 156.515 72.720 156.880 ;
        RECT 72.190 155.815 72.360 156.515 ;
        RECT 72.890 156.435 73.060 157.050 ;
        RECT 73.230 156.695 73.400 157.495 ;
        RECT 73.570 156.995 73.820 157.325 ;
        RECT 74.045 157.025 74.930 157.195 ;
        RECT 72.890 156.345 73.400 156.435 ;
        RECT 71.440 155.535 71.665 155.665 ;
        RECT 71.835 155.595 72.360 155.815 ;
        RECT 72.530 156.175 73.400 156.345 ;
        RECT 71.075 154.945 71.325 155.405 ;
        RECT 71.495 155.395 71.665 155.535 ;
        RECT 72.530 155.395 72.700 156.175 ;
        RECT 73.230 156.105 73.400 156.175 ;
        RECT 72.910 155.925 73.110 155.955 ;
        RECT 73.570 155.925 73.740 156.995 ;
        RECT 73.910 156.105 74.100 156.825 ;
        RECT 72.910 155.625 73.740 155.925 ;
        RECT 74.270 155.895 74.590 156.855 ;
        RECT 71.495 155.225 71.830 155.395 ;
        RECT 72.025 155.225 72.700 155.395 ;
        RECT 73.020 154.945 73.390 155.445 ;
        RECT 73.570 155.395 73.740 155.625 ;
        RECT 74.125 155.565 74.590 155.895 ;
        RECT 74.760 156.185 74.930 157.025 ;
        RECT 75.110 156.995 75.425 157.495 ;
        RECT 75.655 156.765 75.995 157.325 ;
        RECT 75.100 156.390 75.995 156.765 ;
        RECT 76.165 156.485 76.335 157.495 ;
        RECT 75.805 156.185 75.995 156.390 ;
        RECT 76.505 156.435 76.835 157.280 ;
        RECT 77.065 157.060 82.410 157.495 ;
        RECT 76.505 156.355 76.895 156.435 ;
        RECT 76.680 156.305 76.895 156.355 ;
        RECT 74.760 155.855 75.635 156.185 ;
        RECT 75.805 155.855 76.555 156.185 ;
        RECT 74.760 155.395 74.930 155.855 ;
        RECT 75.805 155.685 76.005 155.855 ;
        RECT 76.725 155.725 76.895 156.305 ;
        RECT 76.670 155.685 76.895 155.725 ;
        RECT 73.570 155.225 73.975 155.395 ;
        RECT 74.145 155.225 74.930 155.395 ;
        RECT 75.205 154.945 75.415 155.475 ;
        RECT 75.675 155.160 76.005 155.685 ;
        RECT 76.515 155.600 76.895 155.685 ;
        RECT 76.175 154.945 76.345 155.555 ;
        RECT 76.515 155.165 76.845 155.600 ;
        RECT 78.650 155.490 78.990 156.320 ;
        RECT 80.470 155.810 80.820 157.060 ;
        RECT 82.585 156.405 86.095 157.495 ;
        RECT 82.585 155.715 84.235 156.235 ;
        RECT 84.405 155.885 86.095 156.405 ;
        RECT 87.185 156.330 87.475 157.495 ;
        RECT 87.735 156.565 87.905 157.325 ;
        RECT 88.085 156.735 88.415 157.495 ;
        RECT 87.735 156.395 88.400 156.565 ;
        RECT 88.585 156.420 88.855 157.325 ;
        RECT 88.230 156.250 88.400 156.395 ;
        RECT 87.665 155.845 87.995 156.215 ;
        RECT 88.230 155.920 88.515 156.250 ;
        RECT 77.065 154.945 82.410 155.490 ;
        RECT 82.585 154.945 86.095 155.715 ;
        RECT 87.185 154.945 87.475 155.670 ;
        RECT 88.230 155.665 88.400 155.920 ;
        RECT 87.735 155.495 88.400 155.665 ;
        RECT 88.685 155.620 88.855 156.420 ;
        RECT 90.035 156.565 90.205 157.325 ;
        RECT 90.385 156.735 90.715 157.495 ;
        RECT 90.035 156.395 90.700 156.565 ;
        RECT 90.885 156.420 91.155 157.325 ;
        RECT 91.415 156.825 91.585 157.325 ;
        RECT 91.755 156.995 92.085 157.495 ;
        RECT 91.415 156.655 92.080 156.825 ;
        RECT 90.530 156.250 90.700 156.395 ;
        RECT 89.965 155.845 90.295 156.215 ;
        RECT 90.530 155.920 90.815 156.250 ;
        RECT 90.530 155.665 90.700 155.920 ;
        RECT 87.735 155.115 87.905 155.495 ;
        RECT 88.085 154.945 88.415 155.325 ;
        RECT 88.595 155.115 88.855 155.620 ;
        RECT 90.035 155.495 90.700 155.665 ;
        RECT 90.985 155.620 91.155 156.420 ;
        RECT 91.330 155.835 91.680 156.485 ;
        RECT 91.850 155.665 92.080 156.655 ;
        RECT 90.035 155.115 90.205 155.495 ;
        RECT 90.385 154.945 90.715 155.325 ;
        RECT 90.895 155.115 91.155 155.620 ;
        RECT 91.415 155.495 92.080 155.665 ;
        RECT 91.415 155.205 91.585 155.495 ;
        RECT 91.755 154.945 92.085 155.325 ;
        RECT 92.255 155.205 92.440 157.325 ;
        RECT 92.680 157.035 92.945 157.495 ;
        RECT 93.115 156.900 93.365 157.325 ;
        RECT 93.575 157.050 94.680 157.220 ;
        RECT 93.060 156.770 93.365 156.900 ;
        RECT 92.610 155.575 92.890 156.525 ;
        RECT 93.060 155.665 93.230 156.770 ;
        RECT 93.400 155.985 93.640 156.580 ;
        RECT 93.810 156.515 94.340 156.880 ;
        RECT 93.810 155.815 93.980 156.515 ;
        RECT 94.510 156.435 94.680 157.050 ;
        RECT 94.850 156.695 95.020 157.495 ;
        RECT 95.190 156.995 95.440 157.325 ;
        RECT 95.665 157.025 96.550 157.195 ;
        RECT 94.510 156.345 95.020 156.435 ;
        RECT 93.060 155.535 93.285 155.665 ;
        RECT 93.455 155.595 93.980 155.815 ;
        RECT 94.150 156.175 95.020 156.345 ;
        RECT 92.695 154.945 92.945 155.405 ;
        RECT 93.115 155.395 93.285 155.535 ;
        RECT 94.150 155.395 94.320 156.175 ;
        RECT 94.850 156.105 95.020 156.175 ;
        RECT 94.530 155.925 94.730 155.955 ;
        RECT 95.190 155.925 95.360 156.995 ;
        RECT 95.530 156.105 95.720 156.825 ;
        RECT 94.530 155.625 95.360 155.925 ;
        RECT 95.890 155.895 96.210 156.855 ;
        RECT 93.115 155.225 93.450 155.395 ;
        RECT 93.645 155.225 94.320 155.395 ;
        RECT 94.640 154.945 95.010 155.445 ;
        RECT 95.190 155.395 95.360 155.625 ;
        RECT 95.745 155.565 96.210 155.895 ;
        RECT 96.380 156.185 96.550 157.025 ;
        RECT 96.730 156.995 97.045 157.495 ;
        RECT 97.275 156.765 97.615 157.325 ;
        RECT 96.720 156.390 97.615 156.765 ;
        RECT 97.785 156.485 97.955 157.495 ;
        RECT 97.425 156.185 97.615 156.390 ;
        RECT 98.125 156.435 98.455 157.280 ;
        RECT 99.665 156.435 99.995 157.280 ;
        RECT 100.165 156.485 100.335 157.495 ;
        RECT 100.505 156.765 100.845 157.325 ;
        RECT 101.075 156.995 101.390 157.495 ;
        RECT 101.570 157.025 102.455 157.195 ;
        RECT 98.125 156.355 98.515 156.435 ;
        RECT 98.300 156.305 98.515 156.355 ;
        RECT 96.380 155.855 97.255 156.185 ;
        RECT 97.425 155.855 98.175 156.185 ;
        RECT 96.380 155.395 96.550 155.855 ;
        RECT 97.425 155.685 97.625 155.855 ;
        RECT 98.345 155.725 98.515 156.305 ;
        RECT 98.290 155.685 98.515 155.725 ;
        RECT 95.190 155.225 95.595 155.395 ;
        RECT 95.765 155.225 96.550 155.395 ;
        RECT 96.825 154.945 97.035 155.475 ;
        RECT 97.295 155.160 97.625 155.685 ;
        RECT 98.135 155.600 98.515 155.685 ;
        RECT 99.605 156.355 99.995 156.435 ;
        RECT 100.505 156.390 101.400 156.765 ;
        RECT 99.605 156.305 99.820 156.355 ;
        RECT 99.605 155.725 99.775 156.305 ;
        RECT 100.505 156.185 100.695 156.390 ;
        RECT 101.570 156.185 101.740 157.025 ;
        RECT 102.680 156.995 102.930 157.325 ;
        RECT 99.945 155.855 100.695 156.185 ;
        RECT 100.865 155.855 101.740 156.185 ;
        RECT 99.605 155.685 99.830 155.725 ;
        RECT 100.495 155.685 100.695 155.855 ;
        RECT 99.605 155.600 99.985 155.685 ;
        RECT 97.795 154.945 97.965 155.555 ;
        RECT 98.135 155.165 98.465 155.600 ;
        RECT 99.655 155.165 99.985 155.600 ;
        RECT 100.155 154.945 100.325 155.555 ;
        RECT 100.495 155.160 100.825 155.685 ;
        RECT 101.085 154.945 101.295 155.475 ;
        RECT 101.570 155.395 101.740 155.855 ;
        RECT 101.910 155.895 102.230 156.855 ;
        RECT 102.400 156.105 102.590 156.825 ;
        RECT 102.760 155.925 102.930 156.995 ;
        RECT 103.100 156.695 103.270 157.495 ;
        RECT 103.440 157.050 104.545 157.220 ;
        RECT 103.440 156.435 103.610 157.050 ;
        RECT 104.755 156.900 105.005 157.325 ;
        RECT 105.175 157.035 105.440 157.495 ;
        RECT 103.780 156.515 104.310 156.880 ;
        RECT 104.755 156.770 105.060 156.900 ;
        RECT 103.100 156.345 103.610 156.435 ;
        RECT 103.100 156.175 103.970 156.345 ;
        RECT 103.100 156.105 103.270 156.175 ;
        RECT 103.390 155.925 103.590 155.955 ;
        RECT 101.910 155.565 102.375 155.895 ;
        RECT 102.760 155.625 103.590 155.925 ;
        RECT 102.760 155.395 102.930 155.625 ;
        RECT 101.570 155.225 102.355 155.395 ;
        RECT 102.525 155.225 102.930 155.395 ;
        RECT 103.110 154.945 103.480 155.445 ;
        RECT 103.800 155.395 103.970 156.175 ;
        RECT 104.140 155.815 104.310 156.515 ;
        RECT 104.480 155.985 104.720 156.580 ;
        RECT 104.140 155.595 104.665 155.815 ;
        RECT 104.890 155.665 105.060 156.770 ;
        RECT 104.835 155.535 105.060 155.665 ;
        RECT 105.230 155.575 105.510 156.525 ;
        RECT 104.835 155.395 105.005 155.535 ;
        RECT 103.800 155.225 104.475 155.395 ;
        RECT 104.670 155.225 105.005 155.395 ;
        RECT 105.175 154.945 105.425 155.405 ;
        RECT 105.680 155.205 105.865 157.325 ;
        RECT 106.035 156.995 106.365 157.495 ;
        RECT 106.535 156.825 106.705 157.325 ;
        RECT 106.040 156.655 106.705 156.825 ;
        RECT 106.040 155.665 106.270 156.655 ;
        RECT 107.890 156.525 108.165 157.325 ;
        RECT 108.335 156.695 108.665 157.495 ;
        RECT 108.835 157.155 109.975 157.325 ;
        RECT 108.835 156.525 109.005 157.155 ;
        RECT 106.440 155.835 106.790 156.485 ;
        RECT 107.890 156.315 109.005 156.525 ;
        RECT 109.175 156.525 109.505 156.985 ;
        RECT 109.675 156.695 109.975 157.155 ;
        RECT 109.175 156.305 109.935 156.525 ;
        RECT 110.185 156.405 112.775 157.495 ;
        RECT 107.890 155.935 108.610 156.135 ;
        RECT 108.780 155.935 109.550 156.135 ;
        RECT 109.720 155.765 109.935 156.305 ;
        RECT 106.040 155.495 106.705 155.665 ;
        RECT 106.035 154.945 106.365 155.325 ;
        RECT 106.535 155.205 106.705 155.495 ;
        RECT 107.890 154.945 108.165 155.765 ;
        RECT 108.335 155.595 109.935 155.765 ;
        RECT 110.185 155.715 111.395 156.235 ;
        RECT 111.565 155.885 112.775 156.405 ;
        RECT 112.945 156.330 113.235 157.495 ;
        RECT 113.405 156.355 113.790 157.325 ;
        RECT 113.960 157.035 114.285 157.495 ;
        RECT 114.805 156.865 115.085 157.325 ;
        RECT 113.960 156.645 115.085 156.865 ;
        RECT 108.335 155.585 109.505 155.595 ;
        RECT 108.335 155.115 108.665 155.585 ;
        RECT 108.835 154.945 109.005 155.415 ;
        RECT 109.175 155.115 109.505 155.585 ;
        RECT 109.675 154.945 109.965 155.415 ;
        RECT 110.185 154.945 112.775 155.715 ;
        RECT 113.405 155.685 113.685 156.355 ;
        RECT 113.960 156.185 114.410 156.645 ;
        RECT 115.275 156.475 115.675 157.325 ;
        RECT 116.075 157.035 116.345 157.495 ;
        RECT 116.515 156.865 116.800 157.325 ;
        RECT 113.855 155.855 114.410 156.185 ;
        RECT 114.580 155.915 115.675 156.475 ;
        RECT 113.960 155.745 114.410 155.855 ;
        RECT 112.945 154.945 113.235 155.670 ;
        RECT 113.405 155.115 113.790 155.685 ;
        RECT 113.960 155.575 115.085 155.745 ;
        RECT 113.960 154.945 114.285 155.405 ;
        RECT 114.805 155.115 115.085 155.575 ;
        RECT 115.275 155.115 115.675 155.915 ;
        RECT 115.845 156.645 116.800 156.865 ;
        RECT 117.085 156.645 117.345 157.325 ;
        RECT 117.515 156.715 117.765 157.495 ;
        RECT 118.015 156.945 118.265 157.325 ;
        RECT 118.435 157.115 118.790 157.495 ;
        RECT 119.795 157.105 120.130 157.325 ;
        RECT 119.395 156.945 119.625 156.985 ;
        RECT 118.015 156.745 119.625 156.945 ;
        RECT 118.015 156.735 118.850 156.745 ;
        RECT 119.440 156.655 119.625 156.745 ;
        RECT 115.845 155.745 116.055 156.645 ;
        RECT 116.225 155.915 116.915 156.475 ;
        RECT 115.845 155.575 116.800 155.745 ;
        RECT 116.075 154.945 116.345 155.405 ;
        RECT 116.515 155.115 116.800 155.575 ;
        RECT 117.085 155.455 117.255 156.645 ;
        RECT 118.955 156.545 119.285 156.575 ;
        RECT 117.485 156.485 119.285 156.545 ;
        RECT 119.875 156.485 120.130 157.105 ;
        RECT 121.340 156.865 121.625 157.325 ;
        RECT 121.795 157.035 122.065 157.495 ;
        RECT 121.340 156.645 122.295 156.865 ;
        RECT 117.425 156.375 120.130 156.485 ;
        RECT 117.425 156.340 117.625 156.375 ;
        RECT 117.425 155.765 117.595 156.340 ;
        RECT 118.955 156.315 120.130 156.375 ;
        RECT 117.825 155.900 118.235 156.205 ;
        RECT 118.405 155.935 118.735 156.145 ;
        RECT 117.425 155.645 117.695 155.765 ;
        RECT 117.425 155.600 118.270 155.645 ;
        RECT 117.515 155.475 118.270 155.600 ;
        RECT 118.525 155.535 118.735 155.935 ;
        RECT 118.980 155.935 119.455 156.145 ;
        RECT 119.645 155.935 120.135 156.135 ;
        RECT 118.980 155.535 119.200 155.935 ;
        RECT 121.225 155.915 121.915 156.475 ;
        RECT 122.085 155.745 122.295 156.645 ;
        RECT 117.085 155.445 117.315 155.455 ;
        RECT 117.085 155.115 117.345 155.445 ;
        RECT 118.100 155.325 118.270 155.475 ;
        RECT 117.515 154.945 117.845 155.305 ;
        RECT 118.100 155.115 119.400 155.325 ;
        RECT 119.675 154.945 120.130 155.710 ;
        RECT 121.340 155.575 122.295 155.745 ;
        RECT 122.465 156.475 122.865 157.325 ;
        RECT 123.055 156.865 123.335 157.325 ;
        RECT 123.855 157.035 124.180 157.495 ;
        RECT 123.055 156.645 124.180 156.865 ;
        RECT 122.465 155.915 123.560 156.475 ;
        RECT 123.730 156.185 124.180 156.645 ;
        RECT 124.350 156.355 124.735 157.325 ;
        RECT 121.340 155.115 121.625 155.575 ;
        RECT 121.795 154.945 122.065 155.405 ;
        RECT 122.465 155.115 122.865 155.915 ;
        RECT 123.730 155.855 124.285 156.185 ;
        RECT 123.730 155.745 124.180 155.855 ;
        RECT 123.055 155.575 124.180 155.745 ;
        RECT 124.455 155.685 124.735 156.355 ;
        RECT 123.055 155.115 123.335 155.575 ;
        RECT 123.855 154.945 124.180 155.405 ;
        RECT 124.350 155.115 124.735 155.685 ;
        RECT 124.905 156.645 125.165 157.325 ;
        RECT 125.335 156.715 125.585 157.495 ;
        RECT 125.835 156.945 126.085 157.325 ;
        RECT 126.255 157.115 126.610 157.495 ;
        RECT 127.615 157.105 127.950 157.325 ;
        RECT 127.215 156.945 127.445 156.985 ;
        RECT 125.835 156.745 127.445 156.945 ;
        RECT 125.835 156.735 126.670 156.745 ;
        RECT 127.260 156.655 127.445 156.745 ;
        RECT 124.905 155.455 125.075 156.645 ;
        RECT 126.775 156.545 127.105 156.575 ;
        RECT 125.305 156.485 127.105 156.545 ;
        RECT 127.695 156.485 127.950 157.105 ;
        RECT 125.245 156.375 127.950 156.485 ;
        RECT 125.245 156.340 125.445 156.375 ;
        RECT 125.245 155.765 125.415 156.340 ;
        RECT 126.775 156.315 127.950 156.375 ;
        RECT 128.125 156.315 128.445 157.495 ;
        RECT 128.615 156.475 128.815 157.265 ;
        RECT 129.140 156.665 129.525 157.325 ;
        RECT 129.920 156.735 130.705 157.495 ;
        RECT 129.115 156.565 129.525 156.665 ;
        RECT 128.615 156.305 128.945 156.475 ;
        RECT 129.115 156.355 130.725 156.565 ;
        RECT 125.645 155.900 126.055 156.205 ;
        RECT 128.765 156.185 128.945 156.305 ;
        RECT 126.225 155.935 126.555 156.145 ;
        RECT 125.245 155.645 125.515 155.765 ;
        RECT 125.245 155.600 126.090 155.645 ;
        RECT 125.335 155.475 126.090 155.600 ;
        RECT 126.345 155.535 126.555 155.935 ;
        RECT 126.800 155.935 127.275 156.145 ;
        RECT 127.465 155.935 127.955 156.135 ;
        RECT 128.125 155.935 128.590 156.135 ;
        RECT 128.765 155.935 129.095 156.185 ;
        RECT 129.265 156.135 129.730 156.185 ;
        RECT 129.265 155.965 129.735 156.135 ;
        RECT 129.265 155.935 129.730 155.965 ;
        RECT 129.925 155.935 130.280 156.185 ;
        RECT 126.800 155.535 127.020 155.935 ;
        RECT 130.450 155.755 130.725 156.355 ;
        RECT 124.905 155.445 125.135 155.455 ;
        RECT 124.905 155.115 125.165 155.445 ;
        RECT 125.920 155.325 126.090 155.475 ;
        RECT 125.335 154.945 125.665 155.305 ;
        RECT 125.920 155.115 127.220 155.325 ;
        RECT 127.495 154.945 127.950 155.710 ;
        RECT 128.125 155.555 129.305 155.725 ;
        RECT 128.125 155.140 128.465 155.555 ;
        RECT 128.635 154.945 128.805 155.385 ;
        RECT 128.975 155.335 129.305 155.555 ;
        RECT 129.475 155.575 130.725 155.755 ;
        RECT 129.475 155.505 129.840 155.575 ;
        RECT 128.975 155.155 130.225 155.335 ;
        RECT 130.495 154.945 130.665 155.405 ;
        RECT 130.895 155.225 131.175 157.325 ;
        RECT 131.365 156.605 131.625 157.315 ;
        RECT 131.795 156.785 132.125 157.495 ;
        RECT 132.295 156.605 132.525 157.315 ;
        RECT 131.365 156.365 132.525 156.605 ;
        RECT 132.705 156.585 132.975 157.315 ;
        RECT 133.155 156.765 133.495 157.495 ;
        RECT 132.705 156.365 133.475 156.585 ;
        RECT 131.355 155.855 131.655 156.185 ;
        RECT 131.835 155.875 132.360 156.185 ;
        RECT 132.540 155.875 133.005 156.185 ;
        RECT 131.365 154.945 131.655 155.675 ;
        RECT 131.835 155.235 132.065 155.875 ;
        RECT 133.185 155.695 133.475 156.365 ;
        RECT 132.245 155.495 133.475 155.695 ;
        RECT 132.245 155.125 132.555 155.495 ;
        RECT 132.735 154.945 133.405 155.315 ;
        RECT 133.665 155.125 133.925 157.315 ;
        RECT 135.210 156.525 135.600 156.700 ;
        RECT 136.085 156.695 136.415 157.495 ;
        RECT 136.585 156.705 137.120 157.325 ;
        RECT 135.210 156.355 136.635 156.525 ;
        RECT 135.085 155.625 135.440 156.185 ;
        RECT 135.610 155.455 135.780 156.355 ;
        RECT 135.950 155.625 136.215 156.185 ;
        RECT 136.465 155.855 136.635 156.355 ;
        RECT 136.805 155.685 137.120 156.705 ;
        RECT 137.325 156.355 137.605 157.495 ;
        RECT 137.775 156.345 138.105 157.325 ;
        RECT 138.275 156.355 138.535 157.495 ;
        RECT 137.335 155.915 137.670 156.185 ;
        RECT 137.840 155.745 138.010 156.345 ;
        RECT 138.705 156.330 138.995 157.495 ;
        RECT 139.715 156.565 139.885 157.325 ;
        RECT 140.065 156.735 140.395 157.495 ;
        RECT 139.715 156.395 140.380 156.565 ;
        RECT 140.565 156.420 140.835 157.325 ;
        RECT 141.065 156.435 141.395 157.280 ;
        RECT 141.565 156.485 141.735 157.495 ;
        RECT 141.905 156.765 142.245 157.325 ;
        RECT 142.475 156.995 142.790 157.495 ;
        RECT 142.970 157.025 143.855 157.195 ;
        RECT 140.210 156.250 140.380 156.395 ;
        RECT 138.180 155.935 138.515 156.185 ;
        RECT 139.645 155.845 139.975 156.215 ;
        RECT 140.210 155.920 140.495 156.250 ;
        RECT 135.190 154.945 135.430 155.455 ;
        RECT 135.610 155.125 135.890 155.455 ;
        RECT 136.120 154.945 136.335 155.455 ;
        RECT 136.505 155.115 137.120 155.685 ;
        RECT 137.325 154.945 137.635 155.745 ;
        RECT 137.840 155.115 138.535 155.745 ;
        RECT 138.705 154.945 138.995 155.670 ;
        RECT 140.210 155.665 140.380 155.920 ;
        RECT 139.715 155.495 140.380 155.665 ;
        RECT 140.665 155.620 140.835 156.420 ;
        RECT 139.715 155.115 139.885 155.495 ;
        RECT 140.065 154.945 140.395 155.325 ;
        RECT 140.575 155.115 140.835 155.620 ;
        RECT 141.005 156.355 141.395 156.435 ;
        RECT 141.905 156.390 142.800 156.765 ;
        RECT 141.005 156.305 141.220 156.355 ;
        RECT 141.005 155.725 141.175 156.305 ;
        RECT 141.905 156.185 142.095 156.390 ;
        RECT 142.970 156.185 143.140 157.025 ;
        RECT 144.080 156.995 144.330 157.325 ;
        RECT 141.345 155.855 142.095 156.185 ;
        RECT 142.265 155.855 143.140 156.185 ;
        RECT 141.005 155.685 141.230 155.725 ;
        RECT 141.895 155.685 142.095 155.855 ;
        RECT 141.005 155.600 141.385 155.685 ;
        RECT 141.055 155.165 141.385 155.600 ;
        RECT 141.555 154.945 141.725 155.555 ;
        RECT 141.895 155.160 142.225 155.685 ;
        RECT 142.485 154.945 142.695 155.475 ;
        RECT 142.970 155.395 143.140 155.855 ;
        RECT 143.310 155.895 143.630 156.855 ;
        RECT 143.800 156.105 143.990 156.825 ;
        RECT 144.160 155.925 144.330 156.995 ;
        RECT 144.500 156.695 144.670 157.495 ;
        RECT 144.840 157.050 145.945 157.220 ;
        RECT 144.840 156.435 145.010 157.050 ;
        RECT 146.155 156.900 146.405 157.325 ;
        RECT 146.575 157.035 146.840 157.495 ;
        RECT 145.180 156.515 145.710 156.880 ;
        RECT 146.155 156.770 146.460 156.900 ;
        RECT 144.500 156.345 145.010 156.435 ;
        RECT 144.500 156.175 145.370 156.345 ;
        RECT 144.500 156.105 144.670 156.175 ;
        RECT 144.790 155.925 144.990 155.955 ;
        RECT 143.310 155.565 143.775 155.895 ;
        RECT 144.160 155.625 144.990 155.925 ;
        RECT 144.160 155.395 144.330 155.625 ;
        RECT 142.970 155.225 143.755 155.395 ;
        RECT 143.925 155.225 144.330 155.395 ;
        RECT 144.510 154.945 144.880 155.445 ;
        RECT 145.200 155.395 145.370 156.175 ;
        RECT 145.540 155.815 145.710 156.515 ;
        RECT 145.880 155.985 146.120 156.580 ;
        RECT 145.540 155.595 146.065 155.815 ;
        RECT 146.290 155.665 146.460 156.770 ;
        RECT 146.235 155.535 146.460 155.665 ;
        RECT 146.630 155.575 146.910 156.525 ;
        RECT 146.235 155.395 146.405 155.535 ;
        RECT 145.200 155.225 145.875 155.395 ;
        RECT 146.070 155.225 146.405 155.395 ;
        RECT 146.575 154.945 146.825 155.405 ;
        RECT 147.080 155.205 147.265 157.325 ;
        RECT 147.435 156.995 147.765 157.495 ;
        RECT 147.935 156.825 148.105 157.325 ;
        RECT 147.440 156.655 148.105 156.825 ;
        RECT 147.440 155.665 147.670 156.655 ;
        RECT 147.840 155.835 148.190 156.485 ;
        RECT 148.365 156.405 149.575 157.495 ;
        RECT 148.365 155.695 148.885 156.235 ;
        RECT 149.055 155.865 149.575 156.405 ;
        RECT 149.755 156.385 150.050 157.495 ;
        RECT 150.230 156.185 150.480 157.320 ;
        RECT 150.650 156.385 150.910 157.495 ;
        RECT 151.080 156.595 151.340 157.320 ;
        RECT 151.510 156.765 151.770 157.495 ;
        RECT 151.940 156.595 152.200 157.320 ;
        RECT 152.370 156.765 152.630 157.495 ;
        RECT 152.800 156.595 153.060 157.320 ;
        RECT 153.230 156.765 153.490 157.495 ;
        RECT 153.660 156.595 153.920 157.320 ;
        RECT 154.090 156.765 154.385 157.495 ;
        RECT 151.080 156.355 154.390 156.595 ;
        RECT 147.440 155.495 148.105 155.665 ;
        RECT 147.435 154.945 147.765 155.325 ;
        RECT 147.935 155.205 148.105 155.495 ;
        RECT 148.365 154.945 149.575 155.695 ;
        RECT 149.745 155.575 150.060 156.185 ;
        RECT 150.230 155.935 153.250 156.185 ;
        RECT 149.805 154.945 150.050 155.405 ;
        RECT 150.230 155.125 150.480 155.935 ;
        RECT 153.420 155.765 154.390 156.355 ;
        RECT 155.725 156.405 156.935 157.495 ;
        RECT 155.725 155.865 156.245 156.405 ;
        RECT 151.080 155.595 154.390 155.765 ;
        RECT 156.415 155.695 156.935 156.235 ;
        RECT 150.650 154.945 150.910 155.470 ;
        RECT 151.080 155.140 151.340 155.595 ;
        RECT 151.510 154.945 151.770 155.425 ;
        RECT 151.940 155.140 152.200 155.595 ;
        RECT 152.370 154.945 152.630 155.425 ;
        RECT 152.800 155.140 153.060 155.595 ;
        RECT 153.230 154.945 153.490 155.425 ;
        RECT 153.660 155.140 153.920 155.595 ;
        RECT 154.090 154.945 154.390 155.425 ;
        RECT 155.725 154.945 156.935 155.695 ;
        RECT 22.700 154.775 157.020 154.945 ;
        RECT 22.785 154.025 23.995 154.775 ;
        RECT 24.255 154.225 24.425 154.515 ;
        RECT 24.595 154.395 24.925 154.775 ;
        RECT 24.255 154.055 24.920 154.225 ;
        RECT 22.785 153.485 23.305 154.025 ;
        RECT 23.475 153.315 23.995 153.855 ;
        RECT 22.785 152.225 23.995 153.315 ;
        RECT 24.170 153.235 24.520 153.885 ;
        RECT 24.690 153.065 24.920 154.055 ;
        RECT 24.255 152.895 24.920 153.065 ;
        RECT 24.255 152.395 24.425 152.895 ;
        RECT 24.595 152.225 24.925 152.725 ;
        RECT 25.095 152.395 25.280 154.515 ;
        RECT 25.535 154.315 25.785 154.775 ;
        RECT 25.955 154.325 26.290 154.495 ;
        RECT 26.485 154.325 27.160 154.495 ;
        RECT 25.955 154.185 26.125 154.325 ;
        RECT 25.450 153.195 25.730 154.145 ;
        RECT 25.900 154.055 26.125 154.185 ;
        RECT 25.900 152.950 26.070 154.055 ;
        RECT 26.295 153.905 26.820 154.125 ;
        RECT 26.240 153.140 26.480 153.735 ;
        RECT 26.650 153.205 26.820 153.905 ;
        RECT 26.990 153.545 27.160 154.325 ;
        RECT 27.480 154.275 27.850 154.775 ;
        RECT 28.030 154.325 28.435 154.495 ;
        RECT 28.605 154.325 29.390 154.495 ;
        RECT 28.030 154.095 28.200 154.325 ;
        RECT 27.370 153.795 28.200 154.095 ;
        RECT 28.585 153.825 29.050 154.155 ;
        RECT 27.370 153.765 27.570 153.795 ;
        RECT 27.690 153.545 27.860 153.615 ;
        RECT 26.990 153.375 27.860 153.545 ;
        RECT 27.350 153.285 27.860 153.375 ;
        RECT 25.900 152.820 26.205 152.950 ;
        RECT 26.650 152.840 27.180 153.205 ;
        RECT 25.520 152.225 25.785 152.685 ;
        RECT 25.955 152.395 26.205 152.820 ;
        RECT 27.350 152.670 27.520 153.285 ;
        RECT 26.415 152.500 27.520 152.670 ;
        RECT 27.690 152.225 27.860 153.025 ;
        RECT 28.030 152.725 28.200 153.795 ;
        RECT 28.370 152.895 28.560 153.615 ;
        RECT 28.730 152.865 29.050 153.825 ;
        RECT 29.220 153.865 29.390 154.325 ;
        RECT 29.665 154.245 29.875 154.775 ;
        RECT 30.135 154.035 30.465 154.560 ;
        RECT 30.635 154.165 30.805 154.775 ;
        RECT 30.975 154.120 31.305 154.555 ;
        RECT 30.975 154.035 31.355 154.120 ;
        RECT 30.265 153.865 30.465 154.035 ;
        RECT 31.130 153.995 31.355 154.035 ;
        RECT 29.220 153.535 30.095 153.865 ;
        RECT 30.265 153.535 31.015 153.865 ;
        RECT 28.030 152.395 28.280 152.725 ;
        RECT 29.220 152.695 29.390 153.535 ;
        RECT 30.265 153.330 30.455 153.535 ;
        RECT 31.185 153.415 31.355 153.995 ;
        RECT 31.140 153.365 31.355 153.415 ;
        RECT 29.560 152.955 30.455 153.330 ;
        RECT 30.965 153.285 31.355 153.365 ;
        RECT 31.560 154.035 32.175 154.605 ;
        RECT 32.345 154.265 32.560 154.775 ;
        RECT 32.790 154.265 33.070 154.595 ;
        RECT 33.250 154.265 33.490 154.775 ;
        RECT 28.505 152.525 29.390 152.695 ;
        RECT 29.570 152.225 29.885 152.725 ;
        RECT 30.115 152.395 30.455 152.955 ;
        RECT 30.625 152.225 30.795 153.235 ;
        RECT 30.965 152.440 31.295 153.285 ;
        RECT 31.560 153.015 31.875 154.035 ;
        RECT 32.045 153.365 32.215 153.865 ;
        RECT 32.465 153.535 32.730 154.095 ;
        RECT 32.900 153.365 33.070 154.265 ;
        RECT 33.915 154.225 34.085 154.605 ;
        RECT 34.265 154.395 34.595 154.775 ;
        RECT 33.240 153.535 33.595 154.095 ;
        RECT 33.915 154.055 34.580 154.225 ;
        RECT 34.775 154.100 35.035 154.605 ;
        RECT 33.845 153.505 34.175 153.875 ;
        RECT 34.410 153.800 34.580 154.055 ;
        RECT 34.410 153.470 34.695 153.800 ;
        RECT 32.045 153.195 33.470 153.365 ;
        RECT 34.410 153.325 34.580 153.470 ;
        RECT 31.560 152.395 32.095 153.015 ;
        RECT 32.265 152.225 32.595 153.025 ;
        RECT 33.080 153.020 33.470 153.195 ;
        RECT 33.915 153.155 34.580 153.325 ;
        RECT 34.865 153.300 35.035 154.100 ;
        RECT 35.205 154.025 36.415 154.775 ;
        RECT 35.205 153.485 35.725 154.025 ;
        RECT 36.625 153.955 36.855 154.775 ;
        RECT 37.025 153.975 37.355 154.605 ;
        RECT 35.895 153.315 36.415 153.855 ;
        RECT 36.605 153.535 36.935 153.785 ;
        RECT 37.105 153.375 37.355 153.975 ;
        RECT 37.525 153.955 37.735 154.775 ;
        RECT 37.970 154.010 38.425 154.775 ;
        RECT 38.700 154.395 40.000 154.605 ;
        RECT 40.255 154.415 40.585 154.775 ;
        RECT 39.830 154.245 40.000 154.395 ;
        RECT 40.755 154.275 41.015 154.605 ;
        RECT 40.785 154.265 41.015 154.275 ;
        RECT 38.900 153.785 39.120 154.185 ;
        RECT 37.965 153.585 38.455 153.785 ;
        RECT 38.645 153.575 39.120 153.785 ;
        RECT 39.365 153.785 39.575 154.185 ;
        RECT 39.830 154.120 40.585 154.245 ;
        RECT 39.830 154.075 40.675 154.120 ;
        RECT 40.405 153.955 40.675 154.075 ;
        RECT 39.365 153.575 39.695 153.785 ;
        RECT 39.865 153.515 40.275 153.820 ;
        RECT 33.915 152.395 34.085 153.155 ;
        RECT 34.265 152.225 34.595 152.985 ;
        RECT 34.765 152.395 35.035 153.300 ;
        RECT 35.205 152.225 36.415 153.315 ;
        RECT 36.625 152.225 36.855 153.365 ;
        RECT 37.025 152.395 37.355 153.375 ;
        RECT 37.525 152.225 37.735 153.365 ;
        RECT 37.970 153.345 39.145 153.405 ;
        RECT 40.505 153.380 40.675 153.955 ;
        RECT 40.475 153.345 40.675 153.380 ;
        RECT 37.970 153.235 40.675 153.345 ;
        RECT 37.970 152.615 38.225 153.235 ;
        RECT 38.815 153.175 40.615 153.235 ;
        RECT 38.815 153.145 39.145 153.175 ;
        RECT 40.845 153.075 41.015 154.265 ;
        RECT 41.185 154.005 42.855 154.775 ;
        RECT 43.035 154.245 43.365 154.605 ;
        RECT 43.535 154.415 43.865 154.775 ;
        RECT 44.065 154.245 44.395 154.605 ;
        RECT 43.035 154.035 44.395 154.245 ;
        RECT 44.905 154.015 45.615 154.605 ;
        RECT 41.185 153.485 41.935 154.005 ;
        RECT 42.105 153.315 42.855 153.835 ;
        RECT 43.025 153.535 43.335 153.865 ;
        RECT 43.545 153.535 43.920 153.865 ;
        RECT 44.240 153.535 44.735 153.865 ;
        RECT 38.475 152.975 38.660 153.065 ;
        RECT 39.250 152.975 40.085 152.985 ;
        RECT 38.475 152.775 40.085 152.975 ;
        RECT 38.475 152.735 38.705 152.775 ;
        RECT 37.970 152.395 38.305 152.615 ;
        RECT 39.310 152.225 39.665 152.605 ;
        RECT 39.835 152.395 40.085 152.775 ;
        RECT 40.335 152.225 40.585 153.005 ;
        RECT 40.755 152.395 41.015 153.075 ;
        RECT 41.185 152.225 42.855 153.315 ;
        RECT 43.035 152.225 43.365 153.285 ;
        RECT 43.545 152.610 43.715 153.535 ;
        RECT 43.885 153.045 44.215 153.265 ;
        RECT 44.410 153.245 44.735 153.535 ;
        RECT 44.910 153.245 45.240 153.785 ;
        RECT 45.410 153.045 45.615 154.015 ;
        RECT 45.785 154.005 48.375 154.775 ;
        RECT 48.545 154.050 48.835 154.775 ;
        RECT 49.555 154.225 49.725 154.515 ;
        RECT 49.895 154.395 50.225 154.775 ;
        RECT 49.555 154.055 50.220 154.225 ;
        RECT 45.785 153.485 46.995 154.005 ;
        RECT 47.165 153.315 48.375 153.835 ;
        RECT 43.885 152.815 45.615 153.045 ;
        RECT 43.885 152.415 44.215 152.815 ;
        RECT 44.385 152.225 44.715 152.585 ;
        RECT 44.915 152.395 45.615 152.815 ;
        RECT 45.785 152.225 48.375 153.315 ;
        RECT 48.545 152.225 48.835 153.390 ;
        RECT 49.470 153.235 49.820 153.885 ;
        RECT 49.990 153.065 50.220 154.055 ;
        RECT 49.555 152.895 50.220 153.065 ;
        RECT 49.555 152.395 49.725 152.895 ;
        RECT 49.895 152.225 50.225 152.725 ;
        RECT 50.395 152.395 50.580 154.515 ;
        RECT 50.835 154.315 51.085 154.775 ;
        RECT 51.255 154.325 51.590 154.495 ;
        RECT 51.785 154.325 52.460 154.495 ;
        RECT 51.255 154.185 51.425 154.325 ;
        RECT 50.750 153.195 51.030 154.145 ;
        RECT 51.200 154.055 51.425 154.185 ;
        RECT 51.200 152.950 51.370 154.055 ;
        RECT 51.595 153.905 52.120 154.125 ;
        RECT 51.540 153.140 51.780 153.735 ;
        RECT 51.950 153.205 52.120 153.905 ;
        RECT 52.290 153.545 52.460 154.325 ;
        RECT 52.780 154.275 53.150 154.775 ;
        RECT 53.330 154.325 53.735 154.495 ;
        RECT 53.905 154.325 54.690 154.495 ;
        RECT 53.330 154.095 53.500 154.325 ;
        RECT 52.670 153.795 53.500 154.095 ;
        RECT 53.885 153.825 54.350 154.155 ;
        RECT 52.670 153.765 52.870 153.795 ;
        RECT 52.990 153.545 53.160 153.615 ;
        RECT 52.290 153.375 53.160 153.545 ;
        RECT 52.650 153.285 53.160 153.375 ;
        RECT 51.200 152.820 51.505 152.950 ;
        RECT 51.950 152.840 52.480 153.205 ;
        RECT 50.820 152.225 51.085 152.685 ;
        RECT 51.255 152.395 51.505 152.820 ;
        RECT 52.650 152.670 52.820 153.285 ;
        RECT 51.715 152.500 52.820 152.670 ;
        RECT 52.990 152.225 53.160 153.025 ;
        RECT 53.330 152.725 53.500 153.795 ;
        RECT 53.670 152.895 53.860 153.615 ;
        RECT 54.030 152.865 54.350 153.825 ;
        RECT 54.520 153.865 54.690 154.325 ;
        RECT 54.965 154.245 55.175 154.775 ;
        RECT 55.435 154.035 55.765 154.560 ;
        RECT 55.935 154.165 56.105 154.775 ;
        RECT 56.275 154.120 56.605 154.555 ;
        RECT 56.275 154.035 56.655 154.120 ;
        RECT 55.565 153.865 55.765 154.035 ;
        RECT 56.430 153.995 56.655 154.035 ;
        RECT 54.520 153.535 55.395 153.865 ;
        RECT 55.565 153.535 56.315 153.865 ;
        RECT 53.330 152.395 53.580 152.725 ;
        RECT 54.520 152.695 54.690 153.535 ;
        RECT 55.565 153.330 55.755 153.535 ;
        RECT 56.485 153.415 56.655 153.995 ;
        RECT 56.825 154.005 58.495 154.775 ;
        RECT 58.780 154.145 59.065 154.605 ;
        RECT 59.235 154.315 59.505 154.775 ;
        RECT 56.825 153.485 57.575 154.005 ;
        RECT 58.780 153.975 59.735 154.145 ;
        RECT 56.440 153.365 56.655 153.415 ;
        RECT 54.860 152.955 55.755 153.330 ;
        RECT 56.265 153.285 56.655 153.365 ;
        RECT 57.745 153.315 58.495 153.835 ;
        RECT 53.805 152.525 54.690 152.695 ;
        RECT 54.870 152.225 55.185 152.725 ;
        RECT 55.415 152.395 55.755 152.955 ;
        RECT 55.925 152.225 56.095 153.235 ;
        RECT 56.265 152.440 56.595 153.285 ;
        RECT 56.825 152.225 58.495 153.315 ;
        RECT 58.665 153.245 59.355 153.805 ;
        RECT 59.525 153.075 59.735 153.975 ;
        RECT 58.780 152.855 59.735 153.075 ;
        RECT 59.905 153.805 60.305 154.605 ;
        RECT 60.495 154.145 60.775 154.605 ;
        RECT 61.295 154.315 61.620 154.775 ;
        RECT 60.495 153.975 61.620 154.145 ;
        RECT 61.790 154.035 62.175 154.605 ;
        RECT 62.825 154.045 63.115 154.775 ;
        RECT 61.170 153.865 61.620 153.975 ;
        RECT 59.905 153.245 61.000 153.805 ;
        RECT 61.170 153.535 61.725 153.865 ;
        RECT 58.780 152.395 59.065 152.855 ;
        RECT 59.235 152.225 59.505 152.685 ;
        RECT 59.905 152.395 60.305 153.245 ;
        RECT 61.170 153.075 61.620 153.535 ;
        RECT 61.895 153.365 62.175 154.035 ;
        RECT 62.815 153.535 63.115 153.865 ;
        RECT 63.295 153.845 63.525 154.485 ;
        RECT 63.705 154.225 64.015 154.595 ;
        RECT 64.195 154.405 64.865 154.775 ;
        RECT 63.705 154.025 64.935 154.225 ;
        RECT 63.295 153.535 63.820 153.845 ;
        RECT 64.000 153.535 64.465 153.845 ;
        RECT 60.495 152.855 61.620 153.075 ;
        RECT 60.495 152.395 60.775 152.855 ;
        RECT 61.295 152.225 61.620 152.685 ;
        RECT 61.790 152.395 62.175 153.365 ;
        RECT 64.645 153.355 64.935 154.025 ;
        RECT 62.825 153.115 63.985 153.355 ;
        RECT 62.825 152.405 63.085 153.115 ;
        RECT 63.255 152.225 63.585 152.935 ;
        RECT 63.755 152.405 63.985 153.115 ;
        RECT 64.165 153.135 64.935 153.355 ;
        RECT 64.165 152.405 64.435 153.135 ;
        RECT 64.615 152.225 64.955 152.955 ;
        RECT 65.125 152.405 65.385 154.595 ;
        RECT 66.535 154.305 66.825 154.775 ;
        RECT 66.995 154.135 67.325 154.605 ;
        RECT 67.495 154.305 67.665 154.775 ;
        RECT 67.835 154.135 68.165 154.605 ;
        RECT 66.995 154.125 68.165 154.135 ;
        RECT 66.565 153.955 68.165 154.125 ;
        RECT 68.335 153.955 68.610 154.775 ;
        RECT 68.785 154.230 74.130 154.775 ;
        RECT 66.565 153.415 66.780 153.955 ;
        RECT 66.950 153.585 67.720 153.785 ;
        RECT 67.890 153.585 68.610 153.785 ;
        RECT 66.545 153.245 67.325 153.415 ;
        RECT 66.565 153.195 67.325 153.245 ;
        RECT 66.525 152.565 66.825 153.025 ;
        RECT 66.995 152.735 67.325 153.195 ;
        RECT 67.495 153.195 68.610 153.405 ;
        RECT 70.370 153.400 70.710 154.230 ;
        RECT 74.305 154.050 74.595 154.775 ;
        RECT 75.040 153.965 75.285 154.570 ;
        RECT 75.505 154.240 76.015 154.775 ;
        RECT 67.495 152.565 67.665 153.195 ;
        RECT 66.525 152.395 67.665 152.565 ;
        RECT 67.835 152.225 68.165 153.025 ;
        RECT 68.335 152.395 68.610 153.195 ;
        RECT 72.190 152.660 72.540 153.910 ;
        RECT 74.765 153.795 75.995 153.965 ;
        RECT 68.785 152.225 74.130 152.660 ;
        RECT 74.305 152.225 74.595 153.390 ;
        RECT 74.765 152.985 75.105 153.795 ;
        RECT 75.275 153.230 76.025 153.420 ;
        RECT 74.765 152.575 75.280 152.985 ;
        RECT 75.515 152.225 75.685 152.985 ;
        RECT 75.855 152.565 76.025 153.230 ;
        RECT 76.195 153.245 76.385 154.605 ;
        RECT 76.555 153.755 76.830 154.605 ;
        RECT 77.020 154.240 77.550 154.605 ;
        RECT 77.975 154.375 78.305 154.775 ;
        RECT 77.375 154.205 77.550 154.240 ;
        RECT 76.555 153.585 76.835 153.755 ;
        RECT 76.555 153.445 76.830 153.585 ;
        RECT 77.035 153.245 77.205 154.045 ;
        RECT 76.195 153.075 77.205 153.245 ;
        RECT 77.375 154.035 78.305 154.205 ;
        RECT 78.475 154.035 78.730 154.605 ;
        RECT 77.375 152.905 77.545 154.035 ;
        RECT 78.135 153.865 78.305 154.035 ;
        RECT 76.420 152.735 77.545 152.905 ;
        RECT 77.715 153.535 77.910 153.865 ;
        RECT 78.135 153.535 78.390 153.865 ;
        RECT 77.715 152.565 77.885 153.535 ;
        RECT 78.560 153.365 78.730 154.035 ;
        RECT 78.910 153.955 79.185 154.775 ;
        RECT 79.355 154.135 79.685 154.605 ;
        RECT 79.855 154.305 80.025 154.775 ;
        RECT 80.195 154.135 80.525 154.605 ;
        RECT 80.695 154.305 80.985 154.775 ;
        RECT 79.355 154.125 80.525 154.135 ;
        RECT 79.355 153.955 80.955 154.125 ;
        RECT 78.910 153.585 79.630 153.785 ;
        RECT 79.800 153.585 80.570 153.785 ;
        RECT 80.740 153.415 80.955 153.955 ;
        RECT 81.205 154.025 82.415 154.775 ;
        RECT 82.585 154.125 82.845 154.605 ;
        RECT 83.015 154.235 83.265 154.775 ;
        RECT 81.205 153.485 81.725 154.025 ;
        RECT 75.855 152.395 77.885 152.565 ;
        RECT 78.055 152.225 78.225 153.365 ;
        RECT 78.395 152.395 78.730 153.365 ;
        RECT 78.910 153.195 80.025 153.405 ;
        RECT 78.910 152.395 79.185 153.195 ;
        RECT 79.355 152.225 79.685 153.025 ;
        RECT 79.855 152.565 80.025 153.195 ;
        RECT 80.195 153.195 80.955 153.415 ;
        RECT 81.895 153.315 82.415 153.855 ;
        RECT 80.195 152.735 80.525 153.195 ;
        RECT 80.695 152.565 80.995 153.025 ;
        RECT 79.855 152.395 80.995 152.565 ;
        RECT 81.205 152.225 82.415 153.315 ;
        RECT 82.585 153.095 82.755 154.125 ;
        RECT 83.435 154.070 83.655 154.555 ;
        RECT 82.925 153.475 83.155 153.870 ;
        RECT 83.325 153.645 83.655 154.070 ;
        RECT 83.825 154.395 84.715 154.565 ;
        RECT 83.825 153.670 83.995 154.395 ;
        RECT 84.165 153.840 84.715 154.225 ;
        RECT 84.885 154.035 85.270 154.605 ;
        RECT 85.440 154.315 85.765 154.775 ;
        RECT 86.285 154.145 86.565 154.605 ;
        RECT 83.825 153.600 84.715 153.670 ;
        RECT 83.820 153.575 84.715 153.600 ;
        RECT 83.810 153.560 84.715 153.575 ;
        RECT 83.805 153.545 84.715 153.560 ;
        RECT 83.795 153.540 84.715 153.545 ;
        RECT 83.790 153.530 84.715 153.540 ;
        RECT 83.785 153.520 84.715 153.530 ;
        RECT 83.775 153.515 84.715 153.520 ;
        RECT 83.765 153.505 84.715 153.515 ;
        RECT 83.755 153.500 84.715 153.505 ;
        RECT 83.755 153.495 84.090 153.500 ;
        RECT 83.740 153.490 84.090 153.495 ;
        RECT 83.725 153.480 84.090 153.490 ;
        RECT 83.700 153.475 84.090 153.480 ;
        RECT 82.925 153.470 84.090 153.475 ;
        RECT 82.925 153.435 84.060 153.470 ;
        RECT 82.925 153.410 84.025 153.435 ;
        RECT 82.925 153.380 83.995 153.410 ;
        RECT 82.925 153.350 83.975 153.380 ;
        RECT 82.925 153.320 83.955 153.350 ;
        RECT 82.925 153.310 83.885 153.320 ;
        RECT 82.925 153.300 83.860 153.310 ;
        RECT 82.925 153.285 83.840 153.300 ;
        RECT 82.925 153.270 83.820 153.285 ;
        RECT 83.030 153.260 83.815 153.270 ;
        RECT 83.030 153.225 83.800 153.260 ;
        RECT 82.585 152.395 82.860 153.095 ;
        RECT 83.030 152.975 83.785 153.225 ;
        RECT 83.955 152.905 84.285 153.150 ;
        RECT 84.455 153.050 84.715 153.500 ;
        RECT 84.885 153.365 85.165 154.035 ;
        RECT 85.440 153.975 86.565 154.145 ;
        RECT 85.440 153.865 85.890 153.975 ;
        RECT 85.335 153.535 85.890 153.865 ;
        RECT 86.755 153.805 87.155 154.605 ;
        RECT 87.555 154.315 87.825 154.775 ;
        RECT 87.995 154.145 88.280 154.605 ;
        RECT 84.100 152.880 84.285 152.905 ;
        RECT 84.100 152.780 84.715 152.880 ;
        RECT 83.030 152.225 83.285 152.770 ;
        RECT 83.455 152.395 83.935 152.735 ;
        RECT 84.110 152.225 84.715 152.780 ;
        RECT 84.885 152.395 85.270 153.365 ;
        RECT 85.440 153.075 85.890 153.535 ;
        RECT 86.060 153.245 87.155 153.805 ;
        RECT 85.440 152.855 86.565 153.075 ;
        RECT 85.440 152.225 85.765 152.685 ;
        RECT 86.285 152.395 86.565 152.855 ;
        RECT 86.755 152.395 87.155 153.245 ;
        RECT 87.325 153.975 88.280 154.145 ;
        RECT 87.325 153.075 87.535 153.975 ;
        RECT 88.625 153.955 88.835 154.775 ;
        RECT 89.005 153.975 89.335 154.605 ;
        RECT 87.705 153.245 88.395 153.805 ;
        RECT 89.005 153.375 89.255 153.975 ;
        RECT 89.505 153.955 89.735 154.775 ;
        RECT 89.945 154.035 90.330 154.605 ;
        RECT 90.500 154.315 90.825 154.775 ;
        RECT 91.345 154.145 91.625 154.605 ;
        RECT 89.425 153.535 89.755 153.785 ;
        RECT 87.325 152.855 88.280 153.075 ;
        RECT 87.555 152.225 87.825 152.685 ;
        RECT 87.995 152.395 88.280 152.855 ;
        RECT 88.625 152.225 88.835 153.365 ;
        RECT 89.005 152.395 89.335 153.375 ;
        RECT 89.945 153.365 90.225 154.035 ;
        RECT 90.500 153.975 91.625 154.145 ;
        RECT 90.500 153.865 90.950 153.975 ;
        RECT 90.395 153.535 90.950 153.865 ;
        RECT 91.815 153.805 92.215 154.605 ;
        RECT 92.615 154.315 92.885 154.775 ;
        RECT 93.055 154.145 93.340 154.605 ;
        RECT 89.505 152.225 89.735 153.365 ;
        RECT 89.945 152.395 90.330 153.365 ;
        RECT 90.500 153.075 90.950 153.535 ;
        RECT 91.120 153.245 92.215 153.805 ;
        RECT 90.500 152.855 91.625 153.075 ;
        RECT 90.500 152.225 90.825 152.685 ;
        RECT 91.345 152.395 91.625 152.855 ;
        RECT 91.815 152.395 92.215 153.245 ;
        RECT 92.385 153.975 93.340 154.145 ;
        RECT 94.085 154.125 94.345 154.605 ;
        RECT 94.515 154.315 94.845 154.775 ;
        RECT 95.035 154.135 95.235 154.555 ;
        RECT 92.385 153.075 92.595 153.975 ;
        RECT 92.765 153.245 93.455 153.805 ;
        RECT 94.085 153.095 94.255 154.125 ;
        RECT 94.425 153.435 94.655 153.865 ;
        RECT 94.825 153.615 95.235 154.135 ;
        RECT 95.405 154.290 96.195 154.555 ;
        RECT 95.405 153.435 95.660 154.290 ;
        RECT 96.375 153.955 96.705 154.375 ;
        RECT 96.875 153.955 97.135 154.775 ;
        RECT 97.765 154.395 98.655 154.565 ;
        RECT 96.375 153.865 96.625 153.955 ;
        RECT 95.830 153.615 96.625 153.865 ;
        RECT 97.765 153.840 98.315 154.225 ;
        RECT 94.425 153.265 96.215 153.435 ;
        RECT 92.385 152.855 93.340 153.075 ;
        RECT 92.615 152.225 92.885 152.685 ;
        RECT 93.055 152.395 93.340 152.855 ;
        RECT 94.085 152.395 94.360 153.095 ;
        RECT 94.530 152.970 95.245 153.265 ;
        RECT 95.465 152.905 95.795 153.095 ;
        RECT 94.570 152.225 94.785 152.770 ;
        RECT 94.955 152.395 95.430 152.735 ;
        RECT 95.600 152.730 95.795 152.905 ;
        RECT 95.965 152.900 96.215 153.265 ;
        RECT 95.600 152.225 96.215 152.730 ;
        RECT 96.455 152.395 96.625 153.615 ;
        RECT 96.795 152.905 97.135 153.785 ;
        RECT 98.485 153.670 98.655 154.395 ;
        RECT 97.765 153.600 98.655 153.670 ;
        RECT 98.825 154.070 99.045 154.555 ;
        RECT 99.215 154.235 99.465 154.775 ;
        RECT 99.635 154.125 99.895 154.605 ;
        RECT 98.825 153.645 99.155 154.070 ;
        RECT 97.765 153.575 98.660 153.600 ;
        RECT 97.765 153.560 98.670 153.575 ;
        RECT 97.765 153.545 98.675 153.560 ;
        RECT 97.765 153.540 98.685 153.545 ;
        RECT 97.765 153.530 98.690 153.540 ;
        RECT 97.765 153.520 98.695 153.530 ;
        RECT 97.765 153.515 98.705 153.520 ;
        RECT 97.765 153.505 98.715 153.515 ;
        RECT 97.765 153.500 98.725 153.505 ;
        RECT 97.765 153.050 98.025 153.500 ;
        RECT 98.390 153.495 98.725 153.500 ;
        RECT 98.390 153.490 98.740 153.495 ;
        RECT 98.390 153.480 98.755 153.490 ;
        RECT 98.390 153.475 98.780 153.480 ;
        RECT 99.325 153.475 99.555 153.870 ;
        RECT 98.390 153.470 99.555 153.475 ;
        RECT 98.420 153.435 99.555 153.470 ;
        RECT 98.455 153.410 99.555 153.435 ;
        RECT 98.485 153.380 99.555 153.410 ;
        RECT 98.505 153.350 99.555 153.380 ;
        RECT 98.525 153.320 99.555 153.350 ;
        RECT 98.595 153.310 99.555 153.320 ;
        RECT 98.620 153.300 99.555 153.310 ;
        RECT 98.640 153.285 99.555 153.300 ;
        RECT 98.660 153.270 99.555 153.285 ;
        RECT 98.665 153.260 99.450 153.270 ;
        RECT 98.680 153.225 99.450 153.260 ;
        RECT 98.195 152.905 98.525 153.150 ;
        RECT 98.695 152.975 99.450 153.225 ;
        RECT 99.725 153.095 99.895 154.125 ;
        RECT 100.065 154.050 100.355 154.775 ;
        RECT 101.100 154.145 101.385 154.605 ;
        RECT 101.555 154.315 101.825 154.775 ;
        RECT 101.100 153.975 102.055 154.145 ;
        RECT 98.195 152.880 98.380 152.905 ;
        RECT 97.765 152.780 98.380 152.880 ;
        RECT 96.875 152.225 97.135 152.735 ;
        RECT 97.765 152.225 98.370 152.780 ;
        RECT 98.545 152.395 99.025 152.735 ;
        RECT 99.195 152.225 99.450 152.770 ;
        RECT 99.620 152.395 99.895 153.095 ;
        RECT 100.065 152.225 100.355 153.390 ;
        RECT 100.985 153.245 101.675 153.805 ;
        RECT 101.845 153.075 102.055 153.975 ;
        RECT 101.100 152.855 102.055 153.075 ;
        RECT 102.225 153.805 102.625 154.605 ;
        RECT 102.815 154.145 103.095 154.605 ;
        RECT 103.615 154.315 103.940 154.775 ;
        RECT 102.815 153.975 103.940 154.145 ;
        RECT 104.110 154.035 104.495 154.605 ;
        RECT 103.490 153.865 103.940 153.975 ;
        RECT 102.225 153.245 103.320 153.805 ;
        RECT 103.490 153.535 104.045 153.865 ;
        RECT 101.100 152.395 101.385 152.855 ;
        RECT 101.555 152.225 101.825 152.685 ;
        RECT 102.225 152.395 102.625 153.245 ;
        RECT 103.490 153.075 103.940 153.535 ;
        RECT 104.215 153.365 104.495 154.035 ;
        RECT 104.665 154.005 106.335 154.775 ;
        RECT 106.595 154.225 106.765 154.515 ;
        RECT 106.935 154.395 107.265 154.775 ;
        RECT 106.595 154.055 107.260 154.225 ;
        RECT 104.665 153.485 105.415 154.005 ;
        RECT 102.815 152.855 103.940 153.075 ;
        RECT 102.815 152.395 103.095 152.855 ;
        RECT 103.615 152.225 103.940 152.685 ;
        RECT 104.110 152.395 104.495 153.365 ;
        RECT 105.585 153.315 106.335 153.835 ;
        RECT 104.665 152.225 106.335 153.315 ;
        RECT 106.510 153.235 106.860 153.885 ;
        RECT 107.030 153.065 107.260 154.055 ;
        RECT 106.595 152.895 107.260 153.065 ;
        RECT 106.595 152.395 106.765 152.895 ;
        RECT 106.935 152.225 107.265 152.725 ;
        RECT 107.435 152.395 107.620 154.515 ;
        RECT 107.875 154.315 108.125 154.775 ;
        RECT 108.295 154.325 108.630 154.495 ;
        RECT 108.825 154.325 109.500 154.495 ;
        RECT 108.295 154.185 108.465 154.325 ;
        RECT 107.790 153.195 108.070 154.145 ;
        RECT 108.240 154.055 108.465 154.185 ;
        RECT 108.240 152.950 108.410 154.055 ;
        RECT 108.635 153.905 109.160 154.125 ;
        RECT 108.580 153.140 108.820 153.735 ;
        RECT 108.990 153.205 109.160 153.905 ;
        RECT 109.330 153.545 109.500 154.325 ;
        RECT 109.820 154.275 110.190 154.775 ;
        RECT 110.370 154.325 110.775 154.495 ;
        RECT 110.945 154.325 111.730 154.495 ;
        RECT 110.370 154.095 110.540 154.325 ;
        RECT 109.710 153.795 110.540 154.095 ;
        RECT 110.925 153.825 111.390 154.155 ;
        RECT 109.710 153.765 109.910 153.795 ;
        RECT 110.030 153.545 110.200 153.615 ;
        RECT 109.330 153.375 110.200 153.545 ;
        RECT 109.690 153.285 110.200 153.375 ;
        RECT 108.240 152.820 108.545 152.950 ;
        RECT 108.990 152.840 109.520 153.205 ;
        RECT 107.860 152.225 108.125 152.685 ;
        RECT 108.295 152.395 108.545 152.820 ;
        RECT 109.690 152.670 109.860 153.285 ;
        RECT 108.755 152.500 109.860 152.670 ;
        RECT 110.030 152.225 110.200 153.025 ;
        RECT 110.370 152.725 110.540 153.795 ;
        RECT 110.710 152.895 110.900 153.615 ;
        RECT 111.070 152.865 111.390 153.825 ;
        RECT 111.560 153.865 111.730 154.325 ;
        RECT 112.005 154.245 112.215 154.775 ;
        RECT 112.475 154.035 112.805 154.560 ;
        RECT 112.975 154.165 113.145 154.775 ;
        RECT 113.315 154.120 113.645 154.555 ;
        RECT 113.315 154.035 113.695 154.120 ;
        RECT 112.605 153.865 112.805 154.035 ;
        RECT 113.470 153.995 113.695 154.035 ;
        RECT 111.560 153.535 112.435 153.865 ;
        RECT 112.605 153.535 113.355 153.865 ;
        RECT 110.370 152.395 110.620 152.725 ;
        RECT 111.560 152.695 111.730 153.535 ;
        RECT 112.605 153.330 112.795 153.535 ;
        RECT 113.525 153.415 113.695 153.995 ;
        RECT 113.865 154.005 115.535 154.775 ;
        RECT 115.795 154.225 115.965 154.515 ;
        RECT 116.135 154.395 116.465 154.775 ;
        RECT 115.795 154.055 116.460 154.225 ;
        RECT 113.865 153.485 114.615 154.005 ;
        RECT 113.480 153.365 113.695 153.415 ;
        RECT 111.900 152.955 112.795 153.330 ;
        RECT 113.305 153.285 113.695 153.365 ;
        RECT 114.785 153.315 115.535 153.835 ;
        RECT 110.845 152.525 111.730 152.695 ;
        RECT 111.910 152.225 112.225 152.725 ;
        RECT 112.455 152.395 112.795 152.955 ;
        RECT 112.965 152.225 113.135 153.235 ;
        RECT 113.305 152.440 113.635 153.285 ;
        RECT 113.865 152.225 115.535 153.315 ;
        RECT 115.710 153.235 116.060 153.885 ;
        RECT 116.230 153.065 116.460 154.055 ;
        RECT 115.795 152.895 116.460 153.065 ;
        RECT 115.795 152.395 115.965 152.895 ;
        RECT 116.135 152.225 116.465 152.725 ;
        RECT 116.635 152.395 116.820 154.515 ;
        RECT 117.075 154.315 117.325 154.775 ;
        RECT 117.495 154.325 117.830 154.495 ;
        RECT 118.025 154.325 118.700 154.495 ;
        RECT 117.495 154.185 117.665 154.325 ;
        RECT 116.990 153.195 117.270 154.145 ;
        RECT 117.440 154.055 117.665 154.185 ;
        RECT 117.440 152.950 117.610 154.055 ;
        RECT 117.835 153.905 118.360 154.125 ;
        RECT 117.780 153.140 118.020 153.735 ;
        RECT 118.190 153.205 118.360 153.905 ;
        RECT 118.530 153.545 118.700 154.325 ;
        RECT 119.020 154.275 119.390 154.775 ;
        RECT 119.570 154.325 119.975 154.495 ;
        RECT 120.145 154.325 120.930 154.495 ;
        RECT 119.570 154.095 119.740 154.325 ;
        RECT 118.910 153.795 119.740 154.095 ;
        RECT 120.125 153.825 120.590 154.155 ;
        RECT 118.910 153.765 119.110 153.795 ;
        RECT 119.230 153.545 119.400 153.615 ;
        RECT 118.530 153.375 119.400 153.545 ;
        RECT 118.890 153.285 119.400 153.375 ;
        RECT 117.440 152.820 117.745 152.950 ;
        RECT 118.190 152.840 118.720 153.205 ;
        RECT 117.060 152.225 117.325 152.685 ;
        RECT 117.495 152.395 117.745 152.820 ;
        RECT 118.890 152.670 119.060 153.285 ;
        RECT 117.955 152.500 119.060 152.670 ;
        RECT 119.230 152.225 119.400 153.025 ;
        RECT 119.570 152.725 119.740 153.795 ;
        RECT 119.910 152.895 120.100 153.615 ;
        RECT 120.270 152.865 120.590 153.825 ;
        RECT 120.760 153.865 120.930 154.325 ;
        RECT 121.205 154.245 121.415 154.775 ;
        RECT 121.675 154.035 122.005 154.560 ;
        RECT 122.175 154.165 122.345 154.775 ;
        RECT 122.515 154.120 122.845 154.555 ;
        RECT 122.515 154.035 122.895 154.120 ;
        RECT 121.805 153.865 122.005 154.035 ;
        RECT 122.670 153.995 122.895 154.035 ;
        RECT 120.760 153.535 121.635 153.865 ;
        RECT 121.805 153.535 122.555 153.865 ;
        RECT 119.570 152.395 119.820 152.725 ;
        RECT 120.760 152.695 120.930 153.535 ;
        RECT 121.805 153.330 121.995 153.535 ;
        RECT 122.725 153.415 122.895 153.995 ;
        RECT 123.065 154.005 125.655 154.775 ;
        RECT 125.825 154.050 126.115 154.775 ;
        RECT 126.290 154.010 126.745 154.775 ;
        RECT 127.020 154.395 128.320 154.605 ;
        RECT 128.575 154.415 128.905 154.775 ;
        RECT 128.150 154.245 128.320 154.395 ;
        RECT 129.075 154.275 129.335 154.605 ;
        RECT 129.105 154.265 129.335 154.275 ;
        RECT 123.065 153.485 124.275 154.005 ;
        RECT 122.680 153.365 122.895 153.415 ;
        RECT 121.100 152.955 121.995 153.330 ;
        RECT 122.505 153.285 122.895 153.365 ;
        RECT 124.445 153.315 125.655 153.835 ;
        RECT 127.220 153.785 127.440 154.185 ;
        RECT 126.285 153.585 126.775 153.785 ;
        RECT 126.965 153.575 127.440 153.785 ;
        RECT 127.685 153.785 127.895 154.185 ;
        RECT 128.150 154.120 128.905 154.245 ;
        RECT 128.150 154.075 128.995 154.120 ;
        RECT 128.725 153.955 128.995 154.075 ;
        RECT 127.685 153.575 128.015 153.785 ;
        RECT 128.185 153.515 128.595 153.820 ;
        RECT 120.045 152.525 120.930 152.695 ;
        RECT 121.110 152.225 121.425 152.725 ;
        RECT 121.655 152.395 121.995 152.955 ;
        RECT 122.165 152.225 122.335 153.235 ;
        RECT 122.505 152.440 122.835 153.285 ;
        RECT 123.065 152.225 125.655 153.315 ;
        RECT 125.825 152.225 126.115 153.390 ;
        RECT 126.290 153.345 127.465 153.405 ;
        RECT 128.825 153.380 128.995 153.955 ;
        RECT 128.795 153.345 128.995 153.380 ;
        RECT 126.290 153.235 128.995 153.345 ;
        RECT 126.290 152.615 126.545 153.235 ;
        RECT 127.135 153.175 128.935 153.235 ;
        RECT 127.135 153.145 127.465 153.175 ;
        RECT 129.165 153.075 129.335 154.265 ;
        RECT 129.505 154.005 131.175 154.775 ;
        RECT 129.505 153.485 130.255 154.005 ;
        RECT 131.345 153.975 132.040 154.605 ;
        RECT 132.245 153.975 132.555 154.775 ;
        RECT 132.725 154.125 132.985 154.605 ;
        RECT 133.155 154.235 133.405 154.775 ;
        RECT 130.425 153.315 131.175 153.835 ;
        RECT 131.365 153.535 131.700 153.785 ;
        RECT 131.870 153.375 132.040 153.975 ;
        RECT 132.210 153.535 132.545 153.805 ;
        RECT 126.795 152.975 126.980 153.065 ;
        RECT 127.570 152.975 128.405 152.985 ;
        RECT 126.795 152.775 128.405 152.975 ;
        RECT 126.795 152.735 127.025 152.775 ;
        RECT 126.290 152.395 126.625 152.615 ;
        RECT 127.630 152.225 127.985 152.605 ;
        RECT 128.155 152.395 128.405 152.775 ;
        RECT 128.655 152.225 128.905 153.005 ;
        RECT 129.075 152.395 129.335 153.075 ;
        RECT 129.505 152.225 131.175 153.315 ;
        RECT 131.345 152.225 131.605 153.365 ;
        RECT 131.775 152.395 132.105 153.375 ;
        RECT 132.275 152.225 132.555 153.365 ;
        RECT 132.725 153.095 132.895 154.125 ;
        RECT 133.575 154.095 133.795 154.555 ;
        RECT 133.545 154.070 133.795 154.095 ;
        RECT 133.065 153.475 133.295 153.870 ;
        RECT 133.465 153.645 133.795 154.070 ;
        RECT 133.965 154.395 134.855 154.565 ;
        RECT 133.965 153.670 134.135 154.395 ;
        RECT 134.305 153.840 134.855 154.225 ;
        RECT 135.025 153.955 135.285 154.775 ;
        RECT 135.455 153.955 135.785 154.375 ;
        RECT 135.965 154.290 136.755 154.555 ;
        RECT 135.535 153.865 135.785 153.955 ;
        RECT 133.965 153.600 134.855 153.670 ;
        RECT 133.960 153.575 134.855 153.600 ;
        RECT 133.950 153.560 134.855 153.575 ;
        RECT 133.945 153.545 134.855 153.560 ;
        RECT 133.935 153.540 134.855 153.545 ;
        RECT 133.930 153.530 134.855 153.540 ;
        RECT 133.925 153.520 134.855 153.530 ;
        RECT 133.915 153.515 134.855 153.520 ;
        RECT 133.905 153.505 134.855 153.515 ;
        RECT 133.895 153.500 134.855 153.505 ;
        RECT 133.895 153.495 134.230 153.500 ;
        RECT 133.880 153.490 134.230 153.495 ;
        RECT 133.865 153.480 134.230 153.490 ;
        RECT 133.840 153.475 134.230 153.480 ;
        RECT 133.065 153.470 134.230 153.475 ;
        RECT 133.065 153.435 134.200 153.470 ;
        RECT 133.065 153.410 134.165 153.435 ;
        RECT 133.065 153.380 134.135 153.410 ;
        RECT 133.065 153.350 134.115 153.380 ;
        RECT 133.065 153.320 134.095 153.350 ;
        RECT 133.065 153.310 134.025 153.320 ;
        RECT 133.065 153.300 134.000 153.310 ;
        RECT 133.065 153.285 133.980 153.300 ;
        RECT 133.065 153.270 133.960 153.285 ;
        RECT 133.170 153.260 133.955 153.270 ;
        RECT 133.170 153.225 133.940 153.260 ;
        RECT 132.725 152.395 133.000 153.095 ;
        RECT 133.170 152.975 133.925 153.225 ;
        RECT 134.095 152.905 134.425 153.150 ;
        RECT 134.595 153.050 134.855 153.500 ;
        RECT 135.025 152.905 135.365 153.785 ;
        RECT 135.535 153.615 136.330 153.865 ;
        RECT 134.240 152.880 134.425 152.905 ;
        RECT 134.240 152.780 134.855 152.880 ;
        RECT 133.170 152.225 133.425 152.770 ;
        RECT 133.595 152.395 134.075 152.735 ;
        RECT 134.250 152.225 134.855 152.780 ;
        RECT 135.025 152.225 135.285 152.735 ;
        RECT 135.535 152.395 135.705 153.615 ;
        RECT 136.500 153.435 136.755 154.290 ;
        RECT 136.925 154.135 137.125 154.555 ;
        RECT 137.315 154.315 137.645 154.775 ;
        RECT 136.925 153.615 137.335 154.135 ;
        RECT 137.815 154.125 138.075 154.605 ;
        RECT 137.505 153.435 137.735 153.865 ;
        RECT 135.945 153.265 137.735 153.435 ;
        RECT 135.945 152.900 136.195 153.265 ;
        RECT 136.365 152.905 136.695 153.095 ;
        RECT 136.915 152.970 137.630 153.265 ;
        RECT 137.905 153.095 138.075 154.125 ;
        RECT 138.305 153.955 138.515 154.775 ;
        RECT 138.685 153.975 139.015 154.605 ;
        RECT 138.685 153.375 138.935 153.975 ;
        RECT 139.185 153.955 139.415 154.775 ;
        RECT 139.715 154.225 139.885 154.605 ;
        RECT 140.065 154.395 140.395 154.775 ;
        RECT 139.715 154.055 140.380 154.225 ;
        RECT 140.575 154.100 140.835 154.605 ;
        RECT 141.055 154.120 141.385 154.555 ;
        RECT 141.555 154.165 141.725 154.775 ;
        RECT 139.105 153.535 139.435 153.785 ;
        RECT 139.645 153.505 139.975 153.875 ;
        RECT 140.210 153.800 140.380 154.055 ;
        RECT 140.210 153.470 140.495 153.800 ;
        RECT 136.365 152.730 136.560 152.905 ;
        RECT 135.945 152.225 136.560 152.730 ;
        RECT 136.730 152.395 137.205 152.735 ;
        RECT 137.375 152.225 137.590 152.770 ;
        RECT 137.800 152.395 138.075 153.095 ;
        RECT 138.305 152.225 138.515 153.365 ;
        RECT 138.685 152.395 139.015 153.375 ;
        RECT 139.185 152.225 139.415 153.365 ;
        RECT 140.210 153.325 140.380 153.470 ;
        RECT 139.715 153.155 140.380 153.325 ;
        RECT 140.665 153.300 140.835 154.100 ;
        RECT 139.715 152.395 139.885 153.155 ;
        RECT 140.065 152.225 140.395 152.985 ;
        RECT 140.565 152.395 140.835 153.300 ;
        RECT 141.005 154.035 141.385 154.120 ;
        RECT 141.895 154.035 142.225 154.560 ;
        RECT 142.485 154.245 142.695 154.775 ;
        RECT 142.970 154.325 143.755 154.495 ;
        RECT 143.925 154.325 144.330 154.495 ;
        RECT 141.005 153.995 141.230 154.035 ;
        RECT 141.005 153.415 141.175 153.995 ;
        RECT 141.895 153.865 142.095 154.035 ;
        RECT 142.970 153.865 143.140 154.325 ;
        RECT 141.345 153.535 142.095 153.865 ;
        RECT 142.265 153.535 143.140 153.865 ;
        RECT 141.005 153.365 141.220 153.415 ;
        RECT 141.005 153.285 141.395 153.365 ;
        RECT 141.065 152.440 141.395 153.285 ;
        RECT 141.905 153.330 142.095 153.535 ;
        RECT 141.565 152.225 141.735 153.235 ;
        RECT 141.905 152.955 142.800 153.330 ;
        RECT 141.905 152.395 142.245 152.955 ;
        RECT 142.475 152.225 142.790 152.725 ;
        RECT 142.970 152.695 143.140 153.535 ;
        RECT 143.310 153.825 143.775 154.155 ;
        RECT 144.160 154.095 144.330 154.325 ;
        RECT 144.510 154.275 144.880 154.775 ;
        RECT 145.200 154.325 145.875 154.495 ;
        RECT 146.070 154.325 146.405 154.495 ;
        RECT 143.310 152.865 143.630 153.825 ;
        RECT 144.160 153.795 144.990 154.095 ;
        RECT 143.800 152.895 143.990 153.615 ;
        RECT 144.160 152.725 144.330 153.795 ;
        RECT 144.790 153.765 144.990 153.795 ;
        RECT 144.500 153.545 144.670 153.615 ;
        RECT 145.200 153.545 145.370 154.325 ;
        RECT 146.235 154.185 146.405 154.325 ;
        RECT 146.575 154.315 146.825 154.775 ;
        RECT 144.500 153.375 145.370 153.545 ;
        RECT 145.540 153.905 146.065 154.125 ;
        RECT 146.235 154.055 146.460 154.185 ;
        RECT 144.500 153.285 145.010 153.375 ;
        RECT 142.970 152.525 143.855 152.695 ;
        RECT 144.080 152.395 144.330 152.725 ;
        RECT 144.500 152.225 144.670 153.025 ;
        RECT 144.840 152.670 145.010 153.285 ;
        RECT 145.540 153.205 145.710 153.905 ;
        RECT 145.180 152.840 145.710 153.205 ;
        RECT 145.880 153.140 146.120 153.735 ;
        RECT 146.290 152.950 146.460 154.055 ;
        RECT 146.630 153.195 146.910 154.145 ;
        RECT 146.155 152.820 146.460 152.950 ;
        RECT 144.840 152.500 145.945 152.670 ;
        RECT 146.155 152.395 146.405 152.820 ;
        RECT 146.575 152.225 146.840 152.685 ;
        RECT 147.080 152.395 147.265 154.515 ;
        RECT 147.435 154.395 147.765 154.775 ;
        RECT 147.935 154.225 148.105 154.515 ;
        RECT 147.440 154.055 148.105 154.225 ;
        RECT 147.440 153.065 147.670 154.055 ;
        RECT 148.365 154.005 150.955 154.775 ;
        RECT 151.585 154.050 151.875 154.775 ;
        RECT 152.045 154.005 155.555 154.775 ;
        RECT 155.725 154.025 156.935 154.775 ;
        RECT 147.840 153.235 148.190 153.885 ;
        RECT 148.365 153.485 149.575 154.005 ;
        RECT 149.745 153.315 150.955 153.835 ;
        RECT 152.045 153.485 153.695 154.005 ;
        RECT 147.440 152.895 148.105 153.065 ;
        RECT 147.435 152.225 147.765 152.725 ;
        RECT 147.935 152.395 148.105 152.895 ;
        RECT 148.365 152.225 150.955 153.315 ;
        RECT 151.585 152.225 151.875 153.390 ;
        RECT 153.865 153.315 155.555 153.835 ;
        RECT 152.045 152.225 155.555 153.315 ;
        RECT 155.725 153.315 156.245 153.855 ;
        RECT 156.415 153.485 156.935 154.025 ;
        RECT 155.725 152.225 156.935 153.315 ;
        RECT 22.700 152.055 157.020 152.225 ;
        RECT 22.785 150.965 23.995 152.055 ;
        RECT 22.785 150.255 23.305 150.795 ;
        RECT 23.475 150.425 23.995 150.965 ;
        RECT 25.085 150.980 25.355 151.885 ;
        RECT 25.525 151.295 25.855 152.055 ;
        RECT 26.035 151.125 26.205 151.885 ;
        RECT 22.785 149.505 23.995 150.255 ;
        RECT 25.085 150.180 25.255 150.980 ;
        RECT 25.540 150.955 26.205 151.125 ;
        RECT 26.465 150.965 28.135 152.055 ;
        RECT 25.540 150.810 25.710 150.955 ;
        RECT 25.425 150.480 25.710 150.810 ;
        RECT 25.540 150.225 25.710 150.480 ;
        RECT 25.945 150.405 26.275 150.775 ;
        RECT 26.465 150.275 27.215 150.795 ;
        RECT 27.385 150.445 28.135 150.965 ;
        RECT 28.765 150.915 29.045 152.055 ;
        RECT 29.215 150.905 29.545 151.885 ;
        RECT 29.715 150.915 29.975 152.055 ;
        RECT 30.145 151.545 30.405 152.055 ;
        RECT 28.775 150.475 29.110 150.745 ;
        RECT 29.280 150.305 29.450 150.905 ;
        RECT 29.620 150.495 29.955 150.745 ;
        RECT 30.145 150.495 30.485 151.375 ;
        RECT 30.655 150.665 30.825 151.885 ;
        RECT 31.065 151.550 31.680 152.055 ;
        RECT 31.065 151.015 31.315 151.380 ;
        RECT 31.485 151.375 31.680 151.550 ;
        RECT 31.850 151.545 32.325 151.885 ;
        RECT 32.495 151.510 32.710 152.055 ;
        RECT 31.485 151.185 31.815 151.375 ;
        RECT 32.035 151.015 32.750 151.310 ;
        RECT 32.920 151.185 33.195 151.885 ;
        RECT 31.065 150.845 32.855 151.015 ;
        RECT 30.655 150.415 31.450 150.665 ;
        RECT 30.655 150.325 30.905 150.415 ;
        RECT 25.085 149.675 25.345 150.180 ;
        RECT 25.540 150.055 26.205 150.225 ;
        RECT 25.525 149.505 25.855 149.885 ;
        RECT 26.035 149.675 26.205 150.055 ;
        RECT 26.465 149.505 28.135 150.275 ;
        RECT 28.765 149.505 29.075 150.305 ;
        RECT 29.280 149.675 29.975 150.305 ;
        RECT 30.145 149.505 30.405 150.325 ;
        RECT 30.575 149.905 30.905 150.325 ;
        RECT 31.620 149.990 31.875 150.845 ;
        RECT 31.085 149.725 31.875 149.990 ;
        RECT 32.045 150.145 32.455 150.665 ;
        RECT 32.625 150.415 32.855 150.845 ;
        RECT 33.025 150.155 33.195 151.185 ;
        RECT 32.045 149.725 32.245 150.145 ;
        RECT 32.435 149.505 32.765 149.965 ;
        RECT 32.935 149.675 33.195 150.155 ;
        RECT 33.365 151.185 33.640 151.885 ;
        RECT 33.810 151.510 34.065 152.055 ;
        RECT 34.235 151.545 34.715 151.885 ;
        RECT 34.890 151.500 35.495 152.055 ;
        RECT 34.880 151.400 35.495 151.500 ;
        RECT 34.880 151.375 35.065 151.400 ;
        RECT 33.365 150.155 33.535 151.185 ;
        RECT 33.810 151.055 34.565 151.305 ;
        RECT 34.735 151.130 35.065 151.375 ;
        RECT 33.810 151.020 34.580 151.055 ;
        RECT 33.810 151.010 34.595 151.020 ;
        RECT 33.705 150.995 34.600 151.010 ;
        RECT 33.705 150.980 34.620 150.995 ;
        RECT 33.705 150.970 34.640 150.980 ;
        RECT 33.705 150.960 34.665 150.970 ;
        RECT 33.705 150.930 34.735 150.960 ;
        RECT 33.705 150.900 34.755 150.930 ;
        RECT 33.705 150.870 34.775 150.900 ;
        RECT 33.705 150.845 34.805 150.870 ;
        RECT 33.705 150.810 34.840 150.845 ;
        RECT 33.705 150.805 34.870 150.810 ;
        RECT 33.705 150.410 33.935 150.805 ;
        RECT 34.480 150.800 34.870 150.805 ;
        RECT 34.505 150.790 34.870 150.800 ;
        RECT 34.520 150.785 34.870 150.790 ;
        RECT 34.535 150.780 34.870 150.785 ;
        RECT 35.235 150.780 35.495 151.230 ;
        RECT 35.665 150.890 35.955 152.055 ;
        RECT 36.185 150.915 36.395 152.055 ;
        RECT 36.565 150.905 36.895 151.885 ;
        RECT 37.065 150.915 37.295 152.055 ;
        RECT 37.505 150.965 39.175 152.055 ;
        RECT 34.535 150.775 35.495 150.780 ;
        RECT 34.545 150.765 35.495 150.775 ;
        RECT 34.555 150.760 35.495 150.765 ;
        RECT 34.565 150.750 35.495 150.760 ;
        RECT 34.570 150.740 35.495 150.750 ;
        RECT 34.575 150.735 35.495 150.740 ;
        RECT 34.585 150.720 35.495 150.735 ;
        RECT 34.590 150.705 35.495 150.720 ;
        RECT 34.600 150.680 35.495 150.705 ;
        RECT 34.105 150.210 34.435 150.635 ;
        RECT 33.365 149.675 33.625 150.155 ;
        RECT 33.795 149.505 34.045 150.045 ;
        RECT 34.215 149.725 34.435 150.210 ;
        RECT 34.605 150.610 35.495 150.680 ;
        RECT 34.605 149.885 34.775 150.610 ;
        RECT 34.945 150.055 35.495 150.440 ;
        RECT 34.605 149.715 35.495 149.885 ;
        RECT 35.665 149.505 35.955 150.230 ;
        RECT 36.185 149.505 36.395 150.325 ;
        RECT 36.565 150.305 36.815 150.905 ;
        RECT 36.985 150.495 37.315 150.745 ;
        RECT 36.565 149.675 36.895 150.305 ;
        RECT 37.065 149.505 37.295 150.325 ;
        RECT 37.505 150.275 38.255 150.795 ;
        RECT 38.425 150.445 39.175 150.965 ;
        RECT 39.810 150.915 40.065 152.055 ;
        RECT 40.260 151.505 41.455 151.835 ;
        RECT 40.315 150.745 40.485 151.305 ;
        RECT 40.710 151.085 41.130 151.335 ;
        RECT 41.635 151.255 41.915 152.055 ;
        RECT 40.710 150.915 41.955 151.085 ;
        RECT 42.125 150.915 42.395 151.885 ;
        RECT 41.785 150.745 41.955 150.915 ;
        RECT 39.810 150.495 40.145 150.745 ;
        RECT 40.315 150.415 41.055 150.745 ;
        RECT 41.785 150.415 42.015 150.745 ;
        RECT 40.315 150.325 40.565 150.415 ;
        RECT 37.505 149.505 39.175 150.275 ;
        RECT 39.830 150.155 40.565 150.325 ;
        RECT 41.785 150.245 41.955 150.415 ;
        RECT 39.830 149.685 40.140 150.155 ;
        RECT 41.215 150.075 41.955 150.245 ;
        RECT 42.225 150.180 42.395 150.915 ;
        RECT 40.310 149.505 41.045 149.985 ;
        RECT 41.215 149.725 41.385 150.075 ;
        RECT 41.555 149.505 41.935 149.905 ;
        RECT 42.125 149.835 42.395 150.180 ;
        RECT 43.500 149.685 43.780 151.875 ;
        RECT 43.970 150.915 44.255 152.055 ;
        RECT 44.520 151.405 44.690 151.875 ;
        RECT 44.865 151.575 45.195 152.055 ;
        RECT 45.365 151.405 45.545 151.875 ;
        RECT 44.520 151.205 45.545 151.405 ;
        RECT 43.980 150.235 44.240 150.745 ;
        RECT 44.450 150.415 44.710 151.035 ;
        RECT 44.905 150.415 45.330 151.035 ;
        RECT 45.715 150.765 46.045 151.875 ;
        RECT 46.215 151.645 46.565 152.055 ;
        RECT 46.735 151.465 46.975 151.855 ;
        RECT 45.500 150.465 46.045 150.765 ;
        RECT 46.225 151.265 46.975 151.465 ;
        RECT 47.165 151.465 47.865 151.885 ;
        RECT 48.065 151.695 48.395 152.055 ;
        RECT 48.565 151.465 48.895 151.865 ;
        RECT 46.225 150.585 46.565 151.265 ;
        RECT 47.165 151.235 48.895 151.465 ;
        RECT 45.500 150.235 45.720 150.465 ;
        RECT 43.980 150.045 45.720 150.235 ;
        RECT 43.980 149.505 44.710 149.875 ;
        RECT 45.290 149.685 45.720 150.045 ;
        RECT 45.890 149.505 46.135 150.285 ;
        RECT 46.335 149.685 46.565 150.585 ;
        RECT 46.745 149.745 46.975 151.085 ;
        RECT 47.165 150.355 47.370 151.235 ;
        RECT 47.540 150.495 47.870 151.035 ;
        RECT 48.045 150.745 48.370 151.035 ;
        RECT 48.565 151.015 48.895 151.235 ;
        RECT 49.065 150.745 49.235 151.670 ;
        RECT 49.415 150.995 49.745 152.055 ;
        RECT 49.925 150.965 53.435 152.055 ;
        RECT 48.045 150.415 48.540 150.745 ;
        RECT 48.860 150.415 49.235 150.745 ;
        RECT 49.445 150.415 49.755 150.745 ;
        RECT 47.165 150.265 47.395 150.355 ;
        RECT 49.925 150.275 51.575 150.795 ;
        RECT 51.745 150.445 53.435 150.965 ;
        RECT 47.165 149.675 47.875 150.265 ;
        RECT 48.385 150.035 49.745 150.245 ;
        RECT 48.385 149.675 48.715 150.035 ;
        RECT 48.915 149.505 49.245 149.865 ;
        RECT 49.415 149.675 49.745 150.035 ;
        RECT 49.925 149.505 53.435 150.275 ;
        RECT 53.615 149.685 53.875 151.875 ;
        RECT 54.045 151.325 54.385 152.055 ;
        RECT 54.565 151.145 54.835 151.875 ;
        RECT 54.065 150.925 54.835 151.145 ;
        RECT 55.015 151.165 55.245 151.875 ;
        RECT 55.415 151.345 55.745 152.055 ;
        RECT 55.915 151.165 56.175 151.875 ;
        RECT 56.365 151.500 56.970 152.055 ;
        RECT 57.145 151.545 57.625 151.885 ;
        RECT 57.795 151.510 58.050 152.055 ;
        RECT 56.365 151.400 56.980 151.500 ;
        RECT 56.795 151.375 56.980 151.400 ;
        RECT 55.015 150.925 56.175 151.165 ;
        RECT 54.065 150.255 54.355 150.925 ;
        RECT 56.365 150.780 56.625 151.230 ;
        RECT 56.795 151.130 57.125 151.375 ;
        RECT 57.295 151.055 58.050 151.305 ;
        RECT 58.220 151.185 58.495 151.885 ;
        RECT 57.280 151.020 58.050 151.055 ;
        RECT 57.265 151.010 58.050 151.020 ;
        RECT 57.260 150.995 58.155 151.010 ;
        RECT 57.240 150.980 58.155 150.995 ;
        RECT 57.220 150.970 58.155 150.980 ;
        RECT 57.195 150.960 58.155 150.970 ;
        RECT 57.125 150.930 58.155 150.960 ;
        RECT 57.105 150.900 58.155 150.930 ;
        RECT 57.085 150.870 58.155 150.900 ;
        RECT 57.055 150.845 58.155 150.870 ;
        RECT 57.020 150.810 58.155 150.845 ;
        RECT 56.990 150.805 58.155 150.810 ;
        RECT 56.990 150.800 57.380 150.805 ;
        RECT 56.990 150.790 57.355 150.800 ;
        RECT 56.990 150.785 57.340 150.790 ;
        RECT 56.990 150.780 57.325 150.785 ;
        RECT 56.365 150.775 57.325 150.780 ;
        RECT 56.365 150.765 57.315 150.775 ;
        RECT 56.365 150.760 57.305 150.765 ;
        RECT 56.365 150.750 57.295 150.760 ;
        RECT 54.535 150.435 55.000 150.745 ;
        RECT 55.180 150.435 55.705 150.745 ;
        RECT 54.065 150.055 55.295 150.255 ;
        RECT 54.135 149.505 54.805 149.875 ;
        RECT 54.985 149.685 55.295 150.055 ;
        RECT 55.475 149.795 55.705 150.435 ;
        RECT 55.885 150.415 56.185 150.745 ;
        RECT 56.365 150.740 57.290 150.750 ;
        RECT 56.365 150.735 57.285 150.740 ;
        RECT 56.365 150.720 57.275 150.735 ;
        RECT 56.365 150.705 57.270 150.720 ;
        RECT 56.365 150.680 57.260 150.705 ;
        RECT 56.365 150.610 57.255 150.680 ;
        RECT 55.885 149.505 56.175 150.235 ;
        RECT 56.365 150.055 56.915 150.440 ;
        RECT 57.085 149.885 57.255 150.610 ;
        RECT 56.365 149.715 57.255 149.885 ;
        RECT 57.425 150.210 57.755 150.635 ;
        RECT 57.925 150.410 58.155 150.805 ;
        RECT 57.425 149.725 57.645 150.210 ;
        RECT 58.325 150.155 58.495 151.185 ;
        RECT 57.815 149.505 58.065 150.045 ;
        RECT 58.235 149.675 58.495 150.155 ;
        RECT 58.665 151.185 58.940 151.885 ;
        RECT 59.110 151.510 59.365 152.055 ;
        RECT 59.535 151.545 60.015 151.885 ;
        RECT 60.190 151.500 60.795 152.055 ;
        RECT 60.180 151.400 60.795 151.500 ;
        RECT 60.180 151.375 60.365 151.400 ;
        RECT 58.665 150.155 58.835 151.185 ;
        RECT 59.110 151.055 59.865 151.305 ;
        RECT 60.035 151.130 60.365 151.375 ;
        RECT 59.110 151.020 59.880 151.055 ;
        RECT 59.110 151.010 59.895 151.020 ;
        RECT 59.005 150.995 59.900 151.010 ;
        RECT 59.005 150.980 59.920 150.995 ;
        RECT 59.005 150.970 59.940 150.980 ;
        RECT 59.005 150.960 59.965 150.970 ;
        RECT 59.005 150.930 60.035 150.960 ;
        RECT 59.005 150.900 60.055 150.930 ;
        RECT 59.005 150.870 60.075 150.900 ;
        RECT 59.005 150.845 60.105 150.870 ;
        RECT 59.005 150.810 60.140 150.845 ;
        RECT 59.005 150.805 60.170 150.810 ;
        RECT 59.005 150.410 59.235 150.805 ;
        RECT 59.780 150.800 60.170 150.805 ;
        RECT 59.805 150.790 60.170 150.800 ;
        RECT 59.820 150.785 60.170 150.790 ;
        RECT 59.835 150.780 60.170 150.785 ;
        RECT 60.535 150.780 60.795 151.230 ;
        RECT 61.425 150.890 61.715 152.055 ;
        RECT 62.805 151.500 63.410 152.055 ;
        RECT 63.585 151.545 64.065 151.885 ;
        RECT 64.235 151.510 64.490 152.055 ;
        RECT 62.805 151.400 63.420 151.500 ;
        RECT 63.235 151.375 63.420 151.400 ;
        RECT 59.835 150.775 60.795 150.780 ;
        RECT 59.845 150.765 60.795 150.775 ;
        RECT 59.855 150.760 60.795 150.765 ;
        RECT 59.865 150.750 60.795 150.760 ;
        RECT 59.870 150.740 60.795 150.750 ;
        RECT 59.875 150.735 60.795 150.740 ;
        RECT 59.885 150.720 60.795 150.735 ;
        RECT 59.890 150.705 60.795 150.720 ;
        RECT 59.900 150.680 60.795 150.705 ;
        RECT 59.405 150.210 59.735 150.635 ;
        RECT 59.485 150.185 59.735 150.210 ;
        RECT 58.665 149.675 58.925 150.155 ;
        RECT 59.095 149.505 59.345 150.045 ;
        RECT 59.515 149.725 59.735 150.185 ;
        RECT 59.905 150.610 60.795 150.680 ;
        RECT 62.805 150.780 63.065 151.230 ;
        RECT 63.235 151.130 63.565 151.375 ;
        RECT 63.735 151.055 64.490 151.305 ;
        RECT 64.660 151.185 64.935 151.885 ;
        RECT 63.720 151.020 64.490 151.055 ;
        RECT 63.705 151.010 64.490 151.020 ;
        RECT 63.700 150.995 64.595 151.010 ;
        RECT 63.680 150.980 64.595 150.995 ;
        RECT 63.660 150.970 64.595 150.980 ;
        RECT 63.635 150.960 64.595 150.970 ;
        RECT 63.565 150.930 64.595 150.960 ;
        RECT 63.545 150.900 64.595 150.930 ;
        RECT 63.525 150.870 64.595 150.900 ;
        RECT 63.495 150.845 64.595 150.870 ;
        RECT 63.460 150.810 64.595 150.845 ;
        RECT 63.430 150.805 64.595 150.810 ;
        RECT 63.430 150.800 63.820 150.805 ;
        RECT 63.430 150.790 63.795 150.800 ;
        RECT 63.430 150.785 63.780 150.790 ;
        RECT 63.430 150.780 63.765 150.785 ;
        RECT 62.805 150.775 63.765 150.780 ;
        RECT 62.805 150.765 63.755 150.775 ;
        RECT 62.805 150.760 63.745 150.765 ;
        RECT 62.805 150.750 63.735 150.760 ;
        RECT 62.805 150.740 63.730 150.750 ;
        RECT 62.805 150.735 63.725 150.740 ;
        RECT 62.805 150.720 63.715 150.735 ;
        RECT 62.805 150.705 63.710 150.720 ;
        RECT 62.805 150.680 63.700 150.705 ;
        RECT 62.805 150.610 63.695 150.680 ;
        RECT 59.905 149.885 60.075 150.610 ;
        RECT 60.245 150.055 60.795 150.440 ;
        RECT 59.905 149.715 60.795 149.885 ;
        RECT 61.425 149.505 61.715 150.230 ;
        RECT 62.805 150.055 63.355 150.440 ;
        RECT 63.525 149.885 63.695 150.610 ;
        RECT 62.805 149.715 63.695 149.885 ;
        RECT 63.865 150.210 64.195 150.635 ;
        RECT 64.365 150.410 64.595 150.805 ;
        RECT 63.865 149.725 64.085 150.210 ;
        RECT 64.765 150.155 64.935 151.185 ;
        RECT 65.105 150.965 66.315 152.055 ;
        RECT 66.575 151.310 66.845 152.055 ;
        RECT 67.475 152.050 73.750 152.055 ;
        RECT 67.015 151.140 67.305 151.880 ;
        RECT 67.475 151.325 67.730 152.050 ;
        RECT 67.915 151.155 68.175 151.880 ;
        RECT 68.345 151.325 68.590 152.050 ;
        RECT 68.775 151.155 69.035 151.880 ;
        RECT 69.205 151.325 69.450 152.050 ;
        RECT 69.635 151.155 69.895 151.880 ;
        RECT 70.065 151.325 70.310 152.050 ;
        RECT 70.480 151.155 70.740 151.880 ;
        RECT 70.910 151.325 71.170 152.050 ;
        RECT 71.340 151.155 71.600 151.880 ;
        RECT 71.770 151.325 72.030 152.050 ;
        RECT 72.200 151.155 72.460 151.880 ;
        RECT 72.630 151.325 72.890 152.050 ;
        RECT 73.060 151.155 73.320 151.880 ;
        RECT 73.490 151.255 73.750 152.050 ;
        RECT 67.915 151.140 73.320 151.155 ;
        RECT 64.255 149.505 64.505 150.045 ;
        RECT 64.675 149.675 64.935 150.155 ;
        RECT 65.105 150.255 65.625 150.795 ;
        RECT 65.795 150.425 66.315 150.965 ;
        RECT 66.575 150.915 73.320 151.140 ;
        RECT 66.575 150.325 67.740 150.915 ;
        RECT 73.920 150.745 74.170 151.880 ;
        RECT 74.350 151.245 74.610 152.055 ;
        RECT 74.785 150.745 75.030 151.885 ;
        RECT 75.210 151.245 75.505 152.055 ;
        RECT 75.685 150.965 77.355 152.055 ;
        RECT 77.615 151.385 77.785 151.885 ;
        RECT 77.955 151.555 78.285 152.055 ;
        RECT 77.615 151.215 78.280 151.385 ;
        RECT 67.910 150.495 75.030 150.745 ;
        RECT 65.105 149.505 66.315 150.255 ;
        RECT 66.575 150.155 73.320 150.325 ;
        RECT 66.575 149.505 66.875 149.985 ;
        RECT 67.045 149.700 67.305 150.155 ;
        RECT 67.475 149.505 67.735 149.985 ;
        RECT 67.915 149.700 68.175 150.155 ;
        RECT 68.345 149.505 68.595 149.985 ;
        RECT 68.775 149.700 69.035 150.155 ;
        RECT 69.205 149.505 69.455 149.985 ;
        RECT 69.635 149.700 69.895 150.155 ;
        RECT 70.065 149.505 70.310 149.985 ;
        RECT 70.480 149.700 70.755 150.155 ;
        RECT 70.925 149.505 71.170 149.985 ;
        RECT 71.340 149.700 71.600 150.155 ;
        RECT 71.770 149.505 72.030 149.985 ;
        RECT 72.200 149.700 72.460 150.155 ;
        RECT 72.630 149.505 72.890 149.985 ;
        RECT 73.060 149.700 73.320 150.155 ;
        RECT 73.490 149.505 73.750 150.065 ;
        RECT 73.920 149.685 74.170 150.495 ;
        RECT 74.350 149.505 74.610 150.030 ;
        RECT 74.780 149.685 75.030 150.495 ;
        RECT 75.200 150.185 75.515 150.745 ;
        RECT 75.685 150.275 76.435 150.795 ;
        RECT 76.605 150.445 77.355 150.965 ;
        RECT 77.530 150.395 77.880 151.045 ;
        RECT 75.210 149.505 75.515 150.015 ;
        RECT 75.685 149.505 77.355 150.275 ;
        RECT 78.050 150.225 78.280 151.215 ;
        RECT 77.615 150.055 78.280 150.225 ;
        RECT 77.615 149.765 77.785 150.055 ;
        RECT 77.955 149.505 78.285 149.885 ;
        RECT 78.455 149.765 78.640 151.885 ;
        RECT 78.880 151.595 79.145 152.055 ;
        RECT 79.315 151.460 79.565 151.885 ;
        RECT 79.775 151.610 80.880 151.780 ;
        RECT 79.260 151.330 79.565 151.460 ;
        RECT 78.810 150.135 79.090 151.085 ;
        RECT 79.260 150.225 79.430 151.330 ;
        RECT 79.600 150.545 79.840 151.140 ;
        RECT 80.010 151.075 80.540 151.440 ;
        RECT 80.010 150.375 80.180 151.075 ;
        RECT 80.710 150.995 80.880 151.610 ;
        RECT 81.050 151.255 81.220 152.055 ;
        RECT 81.390 151.555 81.640 151.885 ;
        RECT 81.865 151.585 82.750 151.755 ;
        RECT 80.710 150.905 81.220 150.995 ;
        RECT 79.260 150.095 79.485 150.225 ;
        RECT 79.655 150.155 80.180 150.375 ;
        RECT 80.350 150.735 81.220 150.905 ;
        RECT 78.895 149.505 79.145 149.965 ;
        RECT 79.315 149.955 79.485 150.095 ;
        RECT 80.350 149.955 80.520 150.735 ;
        RECT 81.050 150.665 81.220 150.735 ;
        RECT 80.730 150.485 80.930 150.515 ;
        RECT 81.390 150.485 81.560 151.555 ;
        RECT 81.730 150.665 81.920 151.385 ;
        RECT 80.730 150.185 81.560 150.485 ;
        RECT 82.090 150.455 82.410 151.415 ;
        RECT 79.315 149.785 79.650 149.955 ;
        RECT 79.845 149.785 80.520 149.955 ;
        RECT 80.840 149.505 81.210 150.005 ;
        RECT 81.390 149.955 81.560 150.185 ;
        RECT 81.945 150.125 82.410 150.455 ;
        RECT 82.580 150.745 82.750 151.585 ;
        RECT 82.930 151.555 83.245 152.055 ;
        RECT 83.475 151.325 83.815 151.885 ;
        RECT 82.920 150.950 83.815 151.325 ;
        RECT 83.985 151.045 84.155 152.055 ;
        RECT 83.625 150.745 83.815 150.950 ;
        RECT 84.325 150.995 84.655 151.840 ;
        RECT 84.885 151.500 85.490 152.055 ;
        RECT 85.665 151.545 86.145 151.885 ;
        RECT 86.315 151.510 86.570 152.055 ;
        RECT 84.885 151.400 85.500 151.500 ;
        RECT 85.315 151.375 85.500 151.400 ;
        RECT 84.325 150.915 84.715 150.995 ;
        RECT 84.500 150.865 84.715 150.915 ;
        RECT 82.580 150.415 83.455 150.745 ;
        RECT 83.625 150.415 84.375 150.745 ;
        RECT 82.580 149.955 82.750 150.415 ;
        RECT 83.625 150.245 83.825 150.415 ;
        RECT 84.545 150.285 84.715 150.865 ;
        RECT 84.885 150.780 85.145 151.230 ;
        RECT 85.315 151.130 85.645 151.375 ;
        RECT 85.815 151.055 86.570 151.305 ;
        RECT 86.740 151.185 87.015 151.885 ;
        RECT 85.800 151.020 86.570 151.055 ;
        RECT 85.785 151.010 86.570 151.020 ;
        RECT 85.780 150.995 86.675 151.010 ;
        RECT 85.760 150.980 86.675 150.995 ;
        RECT 85.740 150.970 86.675 150.980 ;
        RECT 85.715 150.960 86.675 150.970 ;
        RECT 85.645 150.930 86.675 150.960 ;
        RECT 85.625 150.900 86.675 150.930 ;
        RECT 85.605 150.870 86.675 150.900 ;
        RECT 85.575 150.845 86.675 150.870 ;
        RECT 85.540 150.810 86.675 150.845 ;
        RECT 85.510 150.805 86.675 150.810 ;
        RECT 85.510 150.800 85.900 150.805 ;
        RECT 85.510 150.790 85.875 150.800 ;
        RECT 85.510 150.785 85.860 150.790 ;
        RECT 85.510 150.780 85.845 150.785 ;
        RECT 84.885 150.775 85.845 150.780 ;
        RECT 84.885 150.765 85.835 150.775 ;
        RECT 84.885 150.760 85.825 150.765 ;
        RECT 84.885 150.750 85.815 150.760 ;
        RECT 84.885 150.740 85.810 150.750 ;
        RECT 84.885 150.735 85.805 150.740 ;
        RECT 84.885 150.720 85.795 150.735 ;
        RECT 84.885 150.705 85.790 150.720 ;
        RECT 84.885 150.680 85.780 150.705 ;
        RECT 84.885 150.610 85.775 150.680 ;
        RECT 84.490 150.245 84.715 150.285 ;
        RECT 81.390 149.785 81.795 149.955 ;
        RECT 81.965 149.785 82.750 149.955 ;
        RECT 83.025 149.505 83.235 150.035 ;
        RECT 83.495 149.720 83.825 150.245 ;
        RECT 84.335 150.160 84.715 150.245 ;
        RECT 83.995 149.505 84.165 150.115 ;
        RECT 84.335 149.725 84.665 150.160 ;
        RECT 84.885 150.055 85.435 150.440 ;
        RECT 85.605 149.885 85.775 150.610 ;
        RECT 84.885 149.715 85.775 149.885 ;
        RECT 85.945 150.210 86.275 150.635 ;
        RECT 86.445 150.410 86.675 150.805 ;
        RECT 85.945 149.725 86.165 150.210 ;
        RECT 86.845 150.155 87.015 151.185 ;
        RECT 87.185 150.890 87.475 152.055 ;
        RECT 87.735 151.385 87.905 151.885 ;
        RECT 88.075 151.555 88.405 152.055 ;
        RECT 87.735 151.215 88.400 151.385 ;
        RECT 87.650 150.395 88.000 151.045 ;
        RECT 86.335 149.505 86.585 150.045 ;
        RECT 86.755 149.675 87.015 150.155 ;
        RECT 87.185 149.505 87.475 150.230 ;
        RECT 88.170 150.225 88.400 151.215 ;
        RECT 87.735 150.055 88.400 150.225 ;
        RECT 87.735 149.765 87.905 150.055 ;
        RECT 88.075 149.505 88.405 149.885 ;
        RECT 88.575 149.765 88.760 151.885 ;
        RECT 89.000 151.595 89.265 152.055 ;
        RECT 89.435 151.460 89.685 151.885 ;
        RECT 89.895 151.610 91.000 151.780 ;
        RECT 89.380 151.330 89.685 151.460 ;
        RECT 88.930 150.135 89.210 151.085 ;
        RECT 89.380 150.225 89.550 151.330 ;
        RECT 89.720 150.545 89.960 151.140 ;
        RECT 90.130 151.075 90.660 151.440 ;
        RECT 90.130 150.375 90.300 151.075 ;
        RECT 90.830 150.995 91.000 151.610 ;
        RECT 91.170 151.255 91.340 152.055 ;
        RECT 91.510 151.555 91.760 151.885 ;
        RECT 91.985 151.585 92.870 151.755 ;
        RECT 90.830 150.905 91.340 150.995 ;
        RECT 89.380 150.095 89.605 150.225 ;
        RECT 89.775 150.155 90.300 150.375 ;
        RECT 90.470 150.735 91.340 150.905 ;
        RECT 89.015 149.505 89.265 149.965 ;
        RECT 89.435 149.955 89.605 150.095 ;
        RECT 90.470 149.955 90.640 150.735 ;
        RECT 91.170 150.665 91.340 150.735 ;
        RECT 90.850 150.485 91.050 150.515 ;
        RECT 91.510 150.485 91.680 151.555 ;
        RECT 91.850 150.665 92.040 151.385 ;
        RECT 90.850 150.185 91.680 150.485 ;
        RECT 92.210 150.455 92.530 151.415 ;
        RECT 89.435 149.785 89.770 149.955 ;
        RECT 89.965 149.785 90.640 149.955 ;
        RECT 90.960 149.505 91.330 150.005 ;
        RECT 91.510 149.955 91.680 150.185 ;
        RECT 92.065 150.125 92.530 150.455 ;
        RECT 92.700 150.745 92.870 151.585 ;
        RECT 93.050 151.555 93.365 152.055 ;
        RECT 93.595 151.325 93.935 151.885 ;
        RECT 93.040 150.950 93.935 151.325 ;
        RECT 94.105 151.045 94.275 152.055 ;
        RECT 93.745 150.745 93.935 150.950 ;
        RECT 94.445 150.995 94.775 151.840 ;
        RECT 94.445 150.915 94.835 150.995 ;
        RECT 94.620 150.865 94.835 150.915 ;
        RECT 92.700 150.415 93.575 150.745 ;
        RECT 93.745 150.415 94.495 150.745 ;
        RECT 92.700 149.955 92.870 150.415 ;
        RECT 93.745 150.245 93.945 150.415 ;
        RECT 94.665 150.285 94.835 150.865 ;
        RECT 94.610 150.245 94.835 150.285 ;
        RECT 91.510 149.785 91.915 149.955 ;
        RECT 92.085 149.785 92.870 149.955 ;
        RECT 93.145 149.505 93.355 150.035 ;
        RECT 93.615 149.720 93.945 150.245 ;
        RECT 94.455 150.160 94.835 150.245 ;
        RECT 94.115 149.505 94.285 150.115 ;
        RECT 94.455 149.725 94.785 150.160 ;
        RECT 95.005 149.785 95.285 151.885 ;
        RECT 95.475 151.295 96.260 152.055 ;
        RECT 96.655 151.225 97.040 151.885 ;
        RECT 96.655 151.125 97.065 151.225 ;
        RECT 95.455 150.915 97.065 151.125 ;
        RECT 97.365 151.035 97.565 151.825 ;
        RECT 95.455 150.315 95.730 150.915 ;
        RECT 97.235 150.865 97.565 151.035 ;
        RECT 97.735 150.875 98.055 152.055 ;
        RECT 98.225 151.335 98.685 151.885 ;
        RECT 98.875 151.335 99.205 152.055 ;
        RECT 97.235 150.745 97.415 150.865 ;
        RECT 95.900 150.495 96.255 150.745 ;
        RECT 96.450 150.695 96.915 150.745 ;
        RECT 96.445 150.525 96.915 150.695 ;
        RECT 96.450 150.495 96.915 150.525 ;
        RECT 97.085 150.495 97.415 150.745 ;
        RECT 97.590 150.495 98.055 150.695 ;
        RECT 95.455 150.135 96.705 150.315 ;
        RECT 96.340 150.065 96.705 150.135 ;
        RECT 96.875 150.115 98.055 150.285 ;
        RECT 95.515 149.505 95.685 149.965 ;
        RECT 96.875 149.895 97.205 150.115 ;
        RECT 95.955 149.715 97.205 149.895 ;
        RECT 97.375 149.505 97.545 149.945 ;
        RECT 97.715 149.700 98.055 150.115 ;
        RECT 98.225 149.965 98.475 151.335 ;
        RECT 99.405 151.165 99.705 151.715 ;
        RECT 99.875 151.385 100.155 152.055 ;
        RECT 100.545 151.545 100.845 152.055 ;
        RECT 101.015 151.545 101.395 151.715 ;
        RECT 101.975 151.545 102.605 152.055 ;
        RECT 101.015 151.375 101.185 151.545 ;
        RECT 102.775 151.375 103.105 151.885 ;
        RECT 103.275 151.545 103.575 152.055 ;
        RECT 98.765 150.995 99.705 151.165 ;
        RECT 100.525 151.175 101.185 151.375 ;
        RECT 101.355 151.205 103.575 151.375 ;
        RECT 98.765 150.745 98.935 150.995 ;
        RECT 100.075 150.745 100.340 151.105 ;
        RECT 98.645 150.415 98.935 150.745 ;
        RECT 99.105 150.495 99.445 150.745 ;
        RECT 99.665 150.495 100.340 150.745 ;
        RECT 98.765 150.325 98.935 150.415 ;
        RECT 98.765 150.135 100.155 150.325 ;
        RECT 98.225 149.675 98.785 149.965 ;
        RECT 98.955 149.505 99.205 149.965 ;
        RECT 99.825 149.775 100.155 150.135 ;
        RECT 100.525 150.245 100.695 151.175 ;
        RECT 101.355 151.005 101.525 151.205 ;
        RECT 100.865 150.835 101.525 151.005 ;
        RECT 101.695 150.865 103.235 151.035 ;
        RECT 100.865 150.415 101.035 150.835 ;
        RECT 101.695 150.665 101.865 150.865 ;
        RECT 101.265 150.495 101.865 150.665 ;
        RECT 102.035 150.495 102.730 150.695 ;
        RECT 102.990 150.415 103.235 150.865 ;
        RECT 101.355 150.245 102.265 150.325 ;
        RECT 100.525 149.765 100.845 150.245 ;
        RECT 101.015 150.155 102.265 150.245 ;
        RECT 101.015 150.075 101.525 150.155 ;
        RECT 101.015 149.675 101.245 150.075 ;
        RECT 101.415 149.505 101.765 149.895 ;
        RECT 101.935 149.675 102.265 150.155 ;
        RECT 102.435 149.505 102.605 150.325 ;
        RECT 103.405 150.245 103.575 151.205 ;
        RECT 103.110 149.700 103.575 150.245 ;
        RECT 104.665 151.205 104.925 151.885 ;
        RECT 105.095 151.275 105.345 152.055 ;
        RECT 105.595 151.505 105.845 151.885 ;
        RECT 106.015 151.675 106.370 152.055 ;
        RECT 107.375 151.665 107.710 151.885 ;
        RECT 106.975 151.505 107.205 151.545 ;
        RECT 105.595 151.305 107.205 151.505 ;
        RECT 105.595 151.295 106.430 151.305 ;
        RECT 107.020 151.215 107.205 151.305 ;
        RECT 104.665 150.005 104.835 151.205 ;
        RECT 106.535 151.105 106.865 151.135 ;
        RECT 105.065 151.045 106.865 151.105 ;
        RECT 107.455 151.045 107.710 151.665 ;
        RECT 105.005 150.935 107.710 151.045 ;
        RECT 107.895 150.945 108.190 152.055 ;
        RECT 105.005 150.900 105.205 150.935 ;
        RECT 105.005 150.325 105.175 150.900 ;
        RECT 106.535 150.875 107.710 150.935 ;
        RECT 105.405 150.460 105.815 150.765 ;
        RECT 108.370 150.745 108.620 151.880 ;
        RECT 108.790 150.945 109.050 152.055 ;
        RECT 109.220 151.155 109.480 151.880 ;
        RECT 109.650 151.325 109.910 152.055 ;
        RECT 110.080 151.155 110.340 151.880 ;
        RECT 110.510 151.325 110.770 152.055 ;
        RECT 110.940 151.155 111.200 151.880 ;
        RECT 111.370 151.325 111.630 152.055 ;
        RECT 111.800 151.155 112.060 151.880 ;
        RECT 112.230 151.325 112.525 152.055 ;
        RECT 109.220 150.915 112.530 151.155 ;
        RECT 105.985 150.495 106.315 150.705 ;
        RECT 105.005 150.205 105.275 150.325 ;
        RECT 105.005 150.160 105.850 150.205 ;
        RECT 105.095 150.035 105.850 150.160 ;
        RECT 106.105 150.095 106.315 150.495 ;
        RECT 106.560 150.495 107.035 150.705 ;
        RECT 107.225 150.495 107.715 150.695 ;
        RECT 106.560 150.095 106.780 150.495 ;
        RECT 104.665 149.675 104.925 150.005 ;
        RECT 105.680 149.885 105.850 150.035 ;
        RECT 105.095 149.505 105.425 149.865 ;
        RECT 105.680 149.675 106.980 149.885 ;
        RECT 107.255 149.505 107.710 150.270 ;
        RECT 107.885 150.135 108.200 150.745 ;
        RECT 108.370 150.495 111.390 150.745 ;
        RECT 107.945 149.505 108.190 149.965 ;
        RECT 108.370 149.685 108.620 150.495 ;
        RECT 111.560 150.325 112.530 150.915 ;
        RECT 112.945 150.890 113.235 152.055 ;
        RECT 113.405 150.965 115.075 152.055 ;
        RECT 115.795 151.385 115.965 151.885 ;
        RECT 116.135 151.555 116.465 152.055 ;
        RECT 115.795 151.215 116.460 151.385 ;
        RECT 109.220 150.155 112.530 150.325 ;
        RECT 113.405 150.275 114.155 150.795 ;
        RECT 114.325 150.445 115.075 150.965 ;
        RECT 115.710 150.395 116.060 151.045 ;
        RECT 108.790 149.505 109.050 150.030 ;
        RECT 109.220 149.700 109.480 150.155 ;
        RECT 109.650 149.505 109.910 149.985 ;
        RECT 110.080 149.700 110.340 150.155 ;
        RECT 110.510 149.505 110.770 149.985 ;
        RECT 110.940 149.700 111.200 150.155 ;
        RECT 111.370 149.505 111.630 149.985 ;
        RECT 111.800 149.700 112.060 150.155 ;
        RECT 112.230 149.505 112.530 149.985 ;
        RECT 112.945 149.505 113.235 150.230 ;
        RECT 113.405 149.505 115.075 150.275 ;
        RECT 116.230 150.225 116.460 151.215 ;
        RECT 115.795 150.055 116.460 150.225 ;
        RECT 115.795 149.765 115.965 150.055 ;
        RECT 116.135 149.505 116.465 149.885 ;
        RECT 116.635 149.765 116.820 151.885 ;
        RECT 117.060 151.595 117.325 152.055 ;
        RECT 117.495 151.460 117.745 151.885 ;
        RECT 117.955 151.610 119.060 151.780 ;
        RECT 117.440 151.330 117.745 151.460 ;
        RECT 116.990 150.135 117.270 151.085 ;
        RECT 117.440 150.225 117.610 151.330 ;
        RECT 117.780 150.545 118.020 151.140 ;
        RECT 118.190 151.075 118.720 151.440 ;
        RECT 118.190 150.375 118.360 151.075 ;
        RECT 118.890 150.995 119.060 151.610 ;
        RECT 119.230 151.255 119.400 152.055 ;
        RECT 119.570 151.555 119.820 151.885 ;
        RECT 120.045 151.585 120.930 151.755 ;
        RECT 118.890 150.905 119.400 150.995 ;
        RECT 117.440 150.095 117.665 150.225 ;
        RECT 117.835 150.155 118.360 150.375 ;
        RECT 118.530 150.735 119.400 150.905 ;
        RECT 117.075 149.505 117.325 149.965 ;
        RECT 117.495 149.955 117.665 150.095 ;
        RECT 118.530 149.955 118.700 150.735 ;
        RECT 119.230 150.665 119.400 150.735 ;
        RECT 118.910 150.485 119.110 150.515 ;
        RECT 119.570 150.485 119.740 151.555 ;
        RECT 119.910 150.665 120.100 151.385 ;
        RECT 118.910 150.185 119.740 150.485 ;
        RECT 120.270 150.455 120.590 151.415 ;
        RECT 117.495 149.785 117.830 149.955 ;
        RECT 118.025 149.785 118.700 149.955 ;
        RECT 119.020 149.505 119.390 150.005 ;
        RECT 119.570 149.955 119.740 150.185 ;
        RECT 120.125 150.125 120.590 150.455 ;
        RECT 120.760 150.745 120.930 151.585 ;
        RECT 121.110 151.555 121.425 152.055 ;
        RECT 121.655 151.325 121.995 151.885 ;
        RECT 121.100 150.950 121.995 151.325 ;
        RECT 122.165 151.045 122.335 152.055 ;
        RECT 121.805 150.745 121.995 150.950 ;
        RECT 122.505 150.995 122.835 151.840 ;
        RECT 122.505 150.915 122.895 150.995 ;
        RECT 122.680 150.865 122.895 150.915 ;
        RECT 120.760 150.415 121.635 150.745 ;
        RECT 121.805 150.415 122.555 150.745 ;
        RECT 120.760 149.955 120.930 150.415 ;
        RECT 121.805 150.245 122.005 150.415 ;
        RECT 122.725 150.285 122.895 150.865 ;
        RECT 122.670 150.245 122.895 150.285 ;
        RECT 119.570 149.785 119.975 149.955 ;
        RECT 120.145 149.785 120.930 149.955 ;
        RECT 121.205 149.505 121.415 150.035 ;
        RECT 121.675 149.720 122.005 150.245 ;
        RECT 122.515 150.160 122.895 150.245 ;
        RECT 123.065 150.915 123.450 151.885 ;
        RECT 123.620 151.595 123.945 152.055 ;
        RECT 124.465 151.425 124.745 151.885 ;
        RECT 123.620 151.205 124.745 151.425 ;
        RECT 123.065 150.245 123.345 150.915 ;
        RECT 123.620 150.745 124.070 151.205 ;
        RECT 124.935 151.035 125.335 151.885 ;
        RECT 125.735 151.595 126.005 152.055 ;
        RECT 126.175 151.425 126.460 151.885 ;
        RECT 123.515 150.415 124.070 150.745 ;
        RECT 124.240 150.475 125.335 151.035 ;
        RECT 123.620 150.305 124.070 150.415 ;
        RECT 122.175 149.505 122.345 150.115 ;
        RECT 122.515 149.725 122.845 150.160 ;
        RECT 123.065 149.675 123.450 150.245 ;
        RECT 123.620 150.135 124.745 150.305 ;
        RECT 123.620 149.505 123.945 149.965 ;
        RECT 124.465 149.675 124.745 150.135 ;
        RECT 124.935 149.675 125.335 150.475 ;
        RECT 125.505 151.205 126.460 151.425 ;
        RECT 126.860 151.425 127.145 151.885 ;
        RECT 127.315 151.595 127.585 152.055 ;
        RECT 126.860 151.205 127.815 151.425 ;
        RECT 125.505 150.305 125.715 151.205 ;
        RECT 125.885 150.475 126.575 151.035 ;
        RECT 126.745 150.475 127.435 151.035 ;
        RECT 127.605 150.305 127.815 151.205 ;
        RECT 125.505 150.135 126.460 150.305 ;
        RECT 125.735 149.505 126.005 149.965 ;
        RECT 126.175 149.675 126.460 150.135 ;
        RECT 126.860 150.135 127.815 150.305 ;
        RECT 127.985 151.035 128.385 151.885 ;
        RECT 128.575 151.425 128.855 151.885 ;
        RECT 129.375 151.595 129.700 152.055 ;
        RECT 128.575 151.205 129.700 151.425 ;
        RECT 127.985 150.475 129.080 151.035 ;
        RECT 129.250 150.745 129.700 151.205 ;
        RECT 129.870 150.915 130.255 151.885 ;
        RECT 126.860 149.675 127.145 150.135 ;
        RECT 127.315 149.505 127.585 149.965 ;
        RECT 127.985 149.675 128.385 150.475 ;
        RECT 129.250 150.415 129.805 150.745 ;
        RECT 129.250 150.305 129.700 150.415 ;
        RECT 128.575 150.135 129.700 150.305 ;
        RECT 129.975 150.245 130.255 150.915 ;
        RECT 130.425 150.875 130.745 152.055 ;
        RECT 130.915 151.035 131.115 151.825 ;
        RECT 131.440 151.225 131.825 151.885 ;
        RECT 132.220 151.295 133.005 152.055 ;
        RECT 131.415 151.125 131.825 151.225 ;
        RECT 130.915 150.865 131.245 151.035 ;
        RECT 131.415 150.915 133.025 151.125 ;
        RECT 131.065 150.745 131.245 150.865 ;
        RECT 130.425 150.495 130.890 150.695 ;
        RECT 131.065 150.495 131.395 150.745 ;
        RECT 131.565 150.695 132.030 150.745 ;
        RECT 131.565 150.525 132.035 150.695 ;
        RECT 131.565 150.495 132.030 150.525 ;
        RECT 132.225 150.495 132.580 150.745 ;
        RECT 132.750 150.315 133.025 150.915 ;
        RECT 128.575 149.675 128.855 150.135 ;
        RECT 129.375 149.505 129.700 149.965 ;
        RECT 129.870 149.675 130.255 150.245 ;
        RECT 130.425 150.115 131.605 150.285 ;
        RECT 130.425 149.700 130.765 150.115 ;
        RECT 130.935 149.505 131.105 149.945 ;
        RECT 131.275 149.895 131.605 150.115 ;
        RECT 131.775 150.135 133.025 150.315 ;
        RECT 131.775 150.065 132.140 150.135 ;
        RECT 131.275 149.715 132.525 149.895 ;
        RECT 132.795 149.505 132.965 149.965 ;
        RECT 133.195 149.785 133.475 151.885 ;
        RECT 133.665 151.165 133.925 151.875 ;
        RECT 134.095 151.345 134.425 152.055 ;
        RECT 134.595 151.165 134.825 151.875 ;
        RECT 133.665 150.925 134.825 151.165 ;
        RECT 135.005 151.145 135.275 151.875 ;
        RECT 135.455 151.325 135.795 152.055 ;
        RECT 135.005 150.925 135.775 151.145 ;
        RECT 133.655 150.415 133.955 150.745 ;
        RECT 134.135 150.435 134.660 150.745 ;
        RECT 134.840 150.435 135.305 150.745 ;
        RECT 133.665 149.505 133.955 150.235 ;
        RECT 134.135 149.795 134.365 150.435 ;
        RECT 135.485 150.255 135.775 150.925 ;
        RECT 134.545 150.055 135.775 150.255 ;
        RECT 134.545 149.685 134.855 150.055 ;
        RECT 135.035 149.505 135.705 149.875 ;
        RECT 135.965 149.685 136.225 151.875 ;
        RECT 136.405 151.085 136.675 151.855 ;
        RECT 136.845 151.275 137.175 152.055 ;
        RECT 137.380 151.450 137.565 151.855 ;
        RECT 137.735 151.630 138.070 152.055 ;
        RECT 137.380 151.275 138.045 151.450 ;
        RECT 136.405 150.915 137.535 151.085 ;
        RECT 136.405 150.005 136.575 150.915 ;
        RECT 136.745 150.165 137.105 150.745 ;
        RECT 137.285 150.415 137.535 150.915 ;
        RECT 137.705 150.245 138.045 151.275 ;
        RECT 138.705 150.890 138.995 152.055 ;
        RECT 139.165 151.620 144.510 152.055 ;
        RECT 137.360 150.075 138.045 150.245 ;
        RECT 136.405 149.675 136.665 150.005 ;
        RECT 136.875 149.505 137.150 149.985 ;
        RECT 137.360 149.675 137.565 150.075 ;
        RECT 137.735 149.505 138.070 149.905 ;
        RECT 138.705 149.505 138.995 150.230 ;
        RECT 140.750 150.050 141.090 150.880 ;
        RECT 142.570 150.370 142.920 151.620 ;
        RECT 144.685 150.965 147.275 152.055 ;
        RECT 147.965 150.995 148.295 151.840 ;
        RECT 148.465 151.045 148.635 152.055 ;
        RECT 148.805 151.325 149.145 151.885 ;
        RECT 149.375 151.555 149.690 152.055 ;
        RECT 149.870 151.585 150.755 151.755 ;
        RECT 144.685 150.275 145.895 150.795 ;
        RECT 146.065 150.445 147.275 150.965 ;
        RECT 147.905 150.915 148.295 150.995 ;
        RECT 148.805 150.950 149.700 151.325 ;
        RECT 147.905 150.865 148.120 150.915 ;
        RECT 147.905 150.285 148.075 150.865 ;
        RECT 148.805 150.745 148.995 150.950 ;
        RECT 149.870 150.745 150.040 151.585 ;
        RECT 150.980 151.555 151.230 151.885 ;
        RECT 148.245 150.415 148.995 150.745 ;
        RECT 149.165 150.415 150.040 150.745 ;
        RECT 139.165 149.505 144.510 150.050 ;
        RECT 144.685 149.505 147.275 150.275 ;
        RECT 147.905 150.245 148.130 150.285 ;
        RECT 148.795 150.245 148.995 150.415 ;
        RECT 147.905 150.160 148.285 150.245 ;
        RECT 147.955 149.725 148.285 150.160 ;
        RECT 148.455 149.505 148.625 150.115 ;
        RECT 148.795 149.720 149.125 150.245 ;
        RECT 149.385 149.505 149.595 150.035 ;
        RECT 149.870 149.955 150.040 150.415 ;
        RECT 150.210 150.455 150.530 151.415 ;
        RECT 150.700 150.665 150.890 151.385 ;
        RECT 151.060 150.485 151.230 151.555 ;
        RECT 151.400 151.255 151.570 152.055 ;
        RECT 151.740 151.610 152.845 151.780 ;
        RECT 151.740 150.995 151.910 151.610 ;
        RECT 153.055 151.460 153.305 151.885 ;
        RECT 153.475 151.595 153.740 152.055 ;
        RECT 152.080 151.075 152.610 151.440 ;
        RECT 153.055 151.330 153.360 151.460 ;
        RECT 151.400 150.905 151.910 150.995 ;
        RECT 151.400 150.735 152.270 150.905 ;
        RECT 151.400 150.665 151.570 150.735 ;
        RECT 151.690 150.485 151.890 150.515 ;
        RECT 150.210 150.125 150.675 150.455 ;
        RECT 151.060 150.185 151.890 150.485 ;
        RECT 151.060 149.955 151.230 150.185 ;
        RECT 149.870 149.785 150.655 149.955 ;
        RECT 150.825 149.785 151.230 149.955 ;
        RECT 151.410 149.505 151.780 150.005 ;
        RECT 152.100 149.955 152.270 150.735 ;
        RECT 152.440 150.375 152.610 151.075 ;
        RECT 152.780 150.545 153.020 151.140 ;
        RECT 152.440 150.155 152.965 150.375 ;
        RECT 153.190 150.225 153.360 151.330 ;
        RECT 153.135 150.095 153.360 150.225 ;
        RECT 153.530 150.135 153.810 151.085 ;
        RECT 153.135 149.955 153.305 150.095 ;
        RECT 152.100 149.785 152.775 149.955 ;
        RECT 152.970 149.785 153.305 149.955 ;
        RECT 153.475 149.505 153.725 149.965 ;
        RECT 153.980 149.765 154.165 151.885 ;
        RECT 154.335 151.555 154.665 152.055 ;
        RECT 154.835 151.385 155.005 151.885 ;
        RECT 154.340 151.215 155.005 151.385 ;
        RECT 154.340 150.225 154.570 151.215 ;
        RECT 154.740 150.395 155.090 151.045 ;
        RECT 155.725 150.965 156.935 152.055 ;
        RECT 155.725 150.425 156.245 150.965 ;
        RECT 156.415 150.255 156.935 150.795 ;
        RECT 154.340 150.055 155.005 150.225 ;
        RECT 154.335 149.505 154.665 149.885 ;
        RECT 154.835 149.765 155.005 150.055 ;
        RECT 155.725 149.505 156.935 150.255 ;
        RECT 22.700 149.335 157.020 149.505 ;
        RECT 22.785 148.585 23.995 149.335 ;
        RECT 24.165 148.790 29.510 149.335 ;
        RECT 22.785 148.045 23.305 148.585 ;
        RECT 23.475 147.875 23.995 148.415 ;
        RECT 25.750 147.960 26.090 148.790 ;
        RECT 29.685 148.565 32.275 149.335 ;
        RECT 32.495 148.680 32.825 149.115 ;
        RECT 32.995 148.725 33.165 149.335 ;
        RECT 32.445 148.595 32.825 148.680 ;
        RECT 33.335 148.595 33.665 149.120 ;
        RECT 33.925 148.805 34.135 149.335 ;
        RECT 34.410 148.885 35.195 149.055 ;
        RECT 35.365 148.885 35.770 149.055 ;
        RECT 22.785 146.785 23.995 147.875 ;
        RECT 27.570 147.220 27.920 148.470 ;
        RECT 29.685 148.045 30.895 148.565 ;
        RECT 32.445 148.555 32.670 148.595 ;
        RECT 31.065 147.875 32.275 148.395 ;
        RECT 24.165 146.785 29.510 147.220 ;
        RECT 29.685 146.785 32.275 147.875 ;
        RECT 32.445 147.975 32.615 148.555 ;
        RECT 33.335 148.425 33.535 148.595 ;
        RECT 34.410 148.425 34.580 148.885 ;
        RECT 32.785 148.095 33.535 148.425 ;
        RECT 33.705 148.095 34.580 148.425 ;
        RECT 32.445 147.925 32.660 147.975 ;
        RECT 32.445 147.845 32.835 147.925 ;
        RECT 32.505 147.000 32.835 147.845 ;
        RECT 33.345 147.890 33.535 148.095 ;
        RECT 33.005 146.785 33.175 147.795 ;
        RECT 33.345 147.515 34.240 147.890 ;
        RECT 33.345 146.955 33.685 147.515 ;
        RECT 33.915 146.785 34.230 147.285 ;
        RECT 34.410 147.255 34.580 148.095 ;
        RECT 34.750 148.385 35.215 148.715 ;
        RECT 35.600 148.655 35.770 148.885 ;
        RECT 35.950 148.835 36.320 149.335 ;
        RECT 36.640 148.885 37.315 149.055 ;
        RECT 37.510 148.885 37.845 149.055 ;
        RECT 34.750 147.425 35.070 148.385 ;
        RECT 35.600 148.355 36.430 148.655 ;
        RECT 35.240 147.455 35.430 148.175 ;
        RECT 35.600 147.285 35.770 148.355 ;
        RECT 36.230 148.325 36.430 148.355 ;
        RECT 35.940 148.105 36.110 148.175 ;
        RECT 36.640 148.105 36.810 148.885 ;
        RECT 37.675 148.745 37.845 148.885 ;
        RECT 38.015 148.875 38.265 149.335 ;
        RECT 35.940 147.935 36.810 148.105 ;
        RECT 36.980 148.465 37.505 148.685 ;
        RECT 37.675 148.615 37.900 148.745 ;
        RECT 35.940 147.845 36.450 147.935 ;
        RECT 34.410 147.085 35.295 147.255 ;
        RECT 35.520 146.955 35.770 147.285 ;
        RECT 35.940 146.785 36.110 147.585 ;
        RECT 36.280 147.230 36.450 147.845 ;
        RECT 36.980 147.765 37.150 148.465 ;
        RECT 36.620 147.400 37.150 147.765 ;
        RECT 37.320 147.700 37.560 148.295 ;
        RECT 37.730 147.510 37.900 148.615 ;
        RECT 38.070 147.755 38.350 148.705 ;
        RECT 37.595 147.380 37.900 147.510 ;
        RECT 36.280 147.060 37.385 147.230 ;
        RECT 37.595 146.955 37.845 147.380 ;
        RECT 38.015 146.785 38.280 147.245 ;
        RECT 38.520 146.955 38.705 149.075 ;
        RECT 38.875 148.955 39.205 149.335 ;
        RECT 39.375 148.785 39.545 149.075 ;
        RECT 39.805 148.790 45.150 149.335 ;
        RECT 38.880 148.615 39.545 148.785 ;
        RECT 38.880 147.625 39.110 148.615 ;
        RECT 39.280 147.795 39.630 148.445 ;
        RECT 41.390 147.960 41.730 148.790 ;
        RECT 45.325 148.565 47.915 149.335 ;
        RECT 48.545 148.610 48.835 149.335 ;
        RECT 38.880 147.455 39.545 147.625 ;
        RECT 38.875 146.785 39.205 147.285 ;
        RECT 39.375 146.955 39.545 147.455 ;
        RECT 43.210 147.220 43.560 148.470 ;
        RECT 45.325 148.045 46.535 148.565 ;
        RECT 49.005 148.535 49.700 149.165 ;
        RECT 49.905 148.535 50.215 149.335 ;
        RECT 50.385 148.535 51.080 149.165 ;
        RECT 51.285 148.535 51.595 149.335 ;
        RECT 52.275 148.680 52.605 149.115 ;
        RECT 52.775 148.725 52.945 149.335 ;
        RECT 52.225 148.595 52.605 148.680 ;
        RECT 53.115 148.595 53.445 149.120 ;
        RECT 53.705 148.805 53.915 149.335 ;
        RECT 54.190 148.885 54.975 149.055 ;
        RECT 55.145 148.885 55.550 149.055 ;
        RECT 52.225 148.555 52.450 148.595 ;
        RECT 46.705 147.875 47.915 148.395 ;
        RECT 49.025 148.095 49.360 148.345 ;
        RECT 39.805 146.785 45.150 147.220 ;
        RECT 45.325 146.785 47.915 147.875 ;
        RECT 48.545 146.785 48.835 147.950 ;
        RECT 49.530 147.935 49.700 148.535 ;
        RECT 49.870 148.095 50.205 148.365 ;
        RECT 50.405 148.095 50.740 148.345 ;
        RECT 50.910 147.935 51.080 148.535 ;
        RECT 51.250 148.095 51.585 148.365 ;
        RECT 52.225 147.975 52.395 148.555 ;
        RECT 53.115 148.425 53.315 148.595 ;
        RECT 54.190 148.425 54.360 148.885 ;
        RECT 52.565 148.095 53.315 148.425 ;
        RECT 53.485 148.095 54.360 148.425 ;
        RECT 49.005 146.785 49.265 147.925 ;
        RECT 49.435 146.955 49.765 147.935 ;
        RECT 49.935 146.785 50.215 147.925 ;
        RECT 50.385 146.785 50.645 147.925 ;
        RECT 50.815 146.955 51.145 147.935 ;
        RECT 52.225 147.925 52.440 147.975 ;
        RECT 51.315 146.785 51.595 147.925 ;
        RECT 52.225 147.845 52.615 147.925 ;
        RECT 52.285 147.000 52.615 147.845 ;
        RECT 53.125 147.890 53.315 148.095 ;
        RECT 52.785 146.785 52.955 147.795 ;
        RECT 53.125 147.515 54.020 147.890 ;
        RECT 53.125 146.955 53.465 147.515 ;
        RECT 53.695 146.785 54.010 147.285 ;
        RECT 54.190 147.255 54.360 148.095 ;
        RECT 54.530 148.385 54.995 148.715 ;
        RECT 55.380 148.655 55.550 148.885 ;
        RECT 55.730 148.835 56.100 149.335 ;
        RECT 56.420 148.885 57.095 149.055 ;
        RECT 57.290 148.885 57.625 149.055 ;
        RECT 54.530 147.425 54.850 148.385 ;
        RECT 55.380 148.355 56.210 148.655 ;
        RECT 55.020 147.455 55.210 148.175 ;
        RECT 55.380 147.285 55.550 148.355 ;
        RECT 56.010 148.325 56.210 148.355 ;
        RECT 55.720 148.105 55.890 148.175 ;
        RECT 56.420 148.105 56.590 148.885 ;
        RECT 57.455 148.745 57.625 148.885 ;
        RECT 57.795 148.875 58.045 149.335 ;
        RECT 55.720 147.935 56.590 148.105 ;
        RECT 56.760 148.465 57.285 148.685 ;
        RECT 57.455 148.615 57.680 148.745 ;
        RECT 55.720 147.845 56.230 147.935 ;
        RECT 54.190 147.085 55.075 147.255 ;
        RECT 55.300 146.955 55.550 147.285 ;
        RECT 55.720 146.785 55.890 147.585 ;
        RECT 56.060 147.230 56.230 147.845 ;
        RECT 56.760 147.765 56.930 148.465 ;
        RECT 56.400 147.400 56.930 147.765 ;
        RECT 57.100 147.700 57.340 148.295 ;
        RECT 57.510 147.510 57.680 148.615 ;
        RECT 57.850 147.755 58.130 148.705 ;
        RECT 57.375 147.380 57.680 147.510 ;
        RECT 56.060 147.060 57.165 147.230 ;
        RECT 57.375 146.955 57.625 147.380 ;
        RECT 57.795 146.785 58.060 147.245 ;
        RECT 58.300 146.955 58.485 149.075 ;
        RECT 58.655 148.955 58.985 149.335 ;
        RECT 59.155 148.785 59.325 149.075 ;
        RECT 58.660 148.615 59.325 148.785 ;
        RECT 59.635 148.680 59.965 149.115 ;
        RECT 60.135 148.725 60.305 149.335 ;
        RECT 58.660 147.625 58.890 148.615 ;
        RECT 59.585 148.595 59.965 148.680 ;
        RECT 60.475 148.595 60.805 149.120 ;
        RECT 61.065 148.805 61.275 149.335 ;
        RECT 61.550 148.885 62.335 149.055 ;
        RECT 62.505 148.885 62.910 149.055 ;
        RECT 59.585 148.555 59.810 148.595 ;
        RECT 59.060 147.795 59.410 148.445 ;
        RECT 59.585 147.975 59.755 148.555 ;
        RECT 60.475 148.425 60.675 148.595 ;
        RECT 61.550 148.425 61.720 148.885 ;
        RECT 59.925 148.095 60.675 148.425 ;
        RECT 60.845 148.095 61.720 148.425 ;
        RECT 59.585 147.925 59.800 147.975 ;
        RECT 59.585 147.845 59.975 147.925 ;
        RECT 58.660 147.455 59.325 147.625 ;
        RECT 58.655 146.785 58.985 147.285 ;
        RECT 59.155 146.955 59.325 147.455 ;
        RECT 59.645 147.000 59.975 147.845 ;
        RECT 60.485 147.890 60.675 148.095 ;
        RECT 60.145 146.785 60.315 147.795 ;
        RECT 60.485 147.515 61.380 147.890 ;
        RECT 60.485 146.955 60.825 147.515 ;
        RECT 61.055 146.785 61.370 147.285 ;
        RECT 61.550 147.255 61.720 148.095 ;
        RECT 61.890 148.385 62.355 148.715 ;
        RECT 62.740 148.655 62.910 148.885 ;
        RECT 63.090 148.835 63.460 149.335 ;
        RECT 63.780 148.885 64.455 149.055 ;
        RECT 64.650 148.885 64.985 149.055 ;
        RECT 61.890 147.425 62.210 148.385 ;
        RECT 62.740 148.355 63.570 148.655 ;
        RECT 62.380 147.455 62.570 148.175 ;
        RECT 62.740 147.285 62.910 148.355 ;
        RECT 63.370 148.325 63.570 148.355 ;
        RECT 63.080 148.105 63.250 148.175 ;
        RECT 63.780 148.105 63.950 148.885 ;
        RECT 64.815 148.745 64.985 148.885 ;
        RECT 65.155 148.875 65.405 149.335 ;
        RECT 63.080 147.935 63.950 148.105 ;
        RECT 64.120 148.465 64.645 148.685 ;
        RECT 64.815 148.615 65.040 148.745 ;
        RECT 63.080 147.845 63.590 147.935 ;
        RECT 61.550 147.085 62.435 147.255 ;
        RECT 62.660 146.955 62.910 147.285 ;
        RECT 63.080 146.785 63.250 147.585 ;
        RECT 63.420 147.230 63.590 147.845 ;
        RECT 64.120 147.765 64.290 148.465 ;
        RECT 63.760 147.400 64.290 147.765 ;
        RECT 64.460 147.700 64.700 148.295 ;
        RECT 64.870 147.510 65.040 148.615 ;
        RECT 65.210 147.755 65.490 148.705 ;
        RECT 64.735 147.380 65.040 147.510 ;
        RECT 63.420 147.060 64.525 147.230 ;
        RECT 64.735 146.955 64.985 147.380 ;
        RECT 65.155 146.785 65.420 147.245 ;
        RECT 65.660 146.955 65.845 149.075 ;
        RECT 66.015 148.955 66.345 149.335 ;
        RECT 66.515 148.785 66.685 149.075 ;
        RECT 66.020 148.615 66.685 148.785 ;
        RECT 66.995 148.680 67.325 149.115 ;
        RECT 67.495 148.725 67.665 149.335 ;
        RECT 66.020 147.625 66.250 148.615 ;
        RECT 66.945 148.595 67.325 148.680 ;
        RECT 67.835 148.595 68.165 149.120 ;
        RECT 68.425 148.805 68.635 149.335 ;
        RECT 68.910 148.885 69.695 149.055 ;
        RECT 69.865 148.885 70.270 149.055 ;
        RECT 66.945 148.555 67.170 148.595 ;
        RECT 66.420 147.795 66.770 148.445 ;
        RECT 66.945 147.975 67.115 148.555 ;
        RECT 67.835 148.425 68.035 148.595 ;
        RECT 68.910 148.425 69.080 148.885 ;
        RECT 67.285 148.095 68.035 148.425 ;
        RECT 68.205 148.095 69.080 148.425 ;
        RECT 66.945 147.925 67.160 147.975 ;
        RECT 66.945 147.845 67.335 147.925 ;
        RECT 66.020 147.455 66.685 147.625 ;
        RECT 66.015 146.785 66.345 147.285 ;
        RECT 66.515 146.955 66.685 147.455 ;
        RECT 67.005 147.000 67.335 147.845 ;
        RECT 67.845 147.890 68.035 148.095 ;
        RECT 67.505 146.785 67.675 147.795 ;
        RECT 67.845 147.515 68.740 147.890 ;
        RECT 67.845 146.955 68.185 147.515 ;
        RECT 68.415 146.785 68.730 147.285 ;
        RECT 68.910 147.255 69.080 148.095 ;
        RECT 69.250 148.385 69.715 148.715 ;
        RECT 70.100 148.655 70.270 148.885 ;
        RECT 70.450 148.835 70.820 149.335 ;
        RECT 71.140 148.885 71.815 149.055 ;
        RECT 72.010 148.885 72.345 149.055 ;
        RECT 69.250 147.425 69.570 148.385 ;
        RECT 70.100 148.355 70.930 148.655 ;
        RECT 69.740 147.455 69.930 148.175 ;
        RECT 70.100 147.285 70.270 148.355 ;
        RECT 70.730 148.325 70.930 148.355 ;
        RECT 70.440 148.105 70.610 148.175 ;
        RECT 71.140 148.105 71.310 148.885 ;
        RECT 72.175 148.745 72.345 148.885 ;
        RECT 72.515 148.875 72.765 149.335 ;
        RECT 70.440 147.935 71.310 148.105 ;
        RECT 71.480 148.465 72.005 148.685 ;
        RECT 72.175 148.615 72.400 148.745 ;
        RECT 70.440 147.845 70.950 147.935 ;
        RECT 68.910 147.085 69.795 147.255 ;
        RECT 70.020 146.955 70.270 147.285 ;
        RECT 70.440 146.785 70.610 147.585 ;
        RECT 70.780 147.230 70.950 147.845 ;
        RECT 71.480 147.765 71.650 148.465 ;
        RECT 71.120 147.400 71.650 147.765 ;
        RECT 71.820 147.700 72.060 148.295 ;
        RECT 72.230 147.510 72.400 148.615 ;
        RECT 72.570 147.755 72.850 148.705 ;
        RECT 72.095 147.380 72.400 147.510 ;
        RECT 70.780 147.060 71.885 147.230 ;
        RECT 72.095 146.955 72.345 147.380 ;
        RECT 72.515 146.785 72.780 147.245 ;
        RECT 73.020 146.955 73.205 149.075 ;
        RECT 73.375 148.955 73.705 149.335 ;
        RECT 73.875 148.785 74.045 149.075 ;
        RECT 73.380 148.615 74.045 148.785 ;
        RECT 73.380 147.625 73.610 148.615 ;
        RECT 74.305 148.610 74.595 149.335 ;
        RECT 75.425 148.705 75.755 149.065 ;
        RECT 76.375 148.875 76.625 149.335 ;
        RECT 76.795 148.875 77.355 149.165 ;
        RECT 75.425 148.515 76.815 148.705 ;
        RECT 73.780 147.795 74.130 148.445 ;
        RECT 76.645 148.425 76.815 148.515 ;
        RECT 75.240 148.095 75.915 148.345 ;
        RECT 76.135 148.095 76.475 148.345 ;
        RECT 76.645 148.095 76.935 148.425 ;
        RECT 73.380 147.455 74.045 147.625 ;
        RECT 73.375 146.785 73.705 147.285 ;
        RECT 73.875 146.955 74.045 147.455 ;
        RECT 74.305 146.785 74.595 147.950 ;
        RECT 75.240 147.735 75.505 148.095 ;
        RECT 76.645 147.845 76.815 148.095 ;
        RECT 75.875 147.675 76.815 147.845 ;
        RECT 75.425 146.785 75.705 147.455 ;
        RECT 75.875 147.125 76.175 147.675 ;
        RECT 77.105 147.505 77.355 148.875 ;
        RECT 76.375 146.785 76.705 147.505 ;
        RECT 76.895 146.955 77.355 147.505 ;
        RECT 77.525 148.660 77.785 149.165 ;
        RECT 77.965 148.955 78.295 149.335 ;
        RECT 78.475 148.785 78.645 149.165 ;
        RECT 77.525 147.860 77.695 148.660 ;
        RECT 77.980 148.615 78.645 148.785 ;
        RECT 77.980 148.360 78.150 148.615 ;
        RECT 78.905 148.565 80.575 149.335 ;
        RECT 77.865 148.030 78.150 148.360 ;
        RECT 78.385 148.065 78.715 148.435 ;
        RECT 78.905 148.045 79.655 148.565 ;
        RECT 77.980 147.885 78.150 148.030 ;
        RECT 77.525 146.955 77.795 147.860 ;
        RECT 77.980 147.715 78.645 147.885 ;
        RECT 79.825 147.875 80.575 148.395 ;
        RECT 77.965 146.785 78.295 147.545 ;
        RECT 78.475 146.955 78.645 147.715 ;
        RECT 78.905 146.785 80.575 147.875 ;
        RECT 81.215 146.965 81.475 149.155 ;
        RECT 81.735 148.965 82.405 149.335 ;
        RECT 82.585 148.785 82.895 149.155 ;
        RECT 81.665 148.585 82.895 148.785 ;
        RECT 81.665 147.915 81.955 148.585 ;
        RECT 83.075 148.405 83.305 149.045 ;
        RECT 83.485 148.605 83.775 149.335 ;
        RECT 83.965 148.585 85.175 149.335 ;
        RECT 85.365 148.605 85.655 149.335 ;
        RECT 82.135 148.095 82.600 148.405 ;
        RECT 82.780 148.095 83.305 148.405 ;
        RECT 83.485 148.095 83.785 148.425 ;
        RECT 83.965 148.045 84.485 148.585 ;
        RECT 81.665 147.695 82.435 147.915 ;
        RECT 81.645 146.785 81.985 147.515 ;
        RECT 82.165 146.965 82.435 147.695 ;
        RECT 82.615 147.675 83.775 147.915 ;
        RECT 84.655 147.875 85.175 148.415 ;
        RECT 85.355 148.095 85.655 148.425 ;
        RECT 85.835 148.405 86.065 149.045 ;
        RECT 86.245 148.785 86.555 149.155 ;
        RECT 86.735 148.965 87.405 149.335 ;
        RECT 86.245 148.585 87.475 148.785 ;
        RECT 85.835 148.095 86.360 148.405 ;
        RECT 86.540 148.095 87.005 148.405 ;
        RECT 87.185 147.915 87.475 148.585 ;
        RECT 82.615 146.965 82.845 147.675 ;
        RECT 83.015 146.785 83.345 147.495 ;
        RECT 83.515 146.965 83.775 147.675 ;
        RECT 83.965 146.785 85.175 147.875 ;
        RECT 85.365 147.675 86.525 147.915 ;
        RECT 85.365 146.965 85.625 147.675 ;
        RECT 85.795 146.785 86.125 147.495 ;
        RECT 86.295 146.965 86.525 147.675 ;
        RECT 86.705 147.695 87.475 147.915 ;
        RECT 86.705 146.965 86.975 147.695 ;
        RECT 87.155 146.785 87.495 147.515 ;
        RECT 87.665 146.965 87.925 149.155 ;
        RECT 88.145 148.515 88.375 149.335 ;
        RECT 88.545 148.535 88.875 149.165 ;
        RECT 88.125 148.095 88.455 148.345 ;
        RECT 88.625 147.935 88.875 148.535 ;
        RECT 89.045 148.515 89.255 149.335 ;
        RECT 89.575 148.855 89.875 149.335 ;
        RECT 90.045 148.685 90.305 149.140 ;
        RECT 90.475 148.855 90.735 149.335 ;
        RECT 90.915 148.685 91.175 149.140 ;
        RECT 91.345 148.855 91.595 149.335 ;
        RECT 91.775 148.685 92.035 149.140 ;
        RECT 92.205 148.855 92.455 149.335 ;
        RECT 92.635 148.685 92.895 149.140 ;
        RECT 93.065 148.855 93.310 149.335 ;
        RECT 93.480 148.685 93.755 149.140 ;
        RECT 93.925 148.855 94.170 149.335 ;
        RECT 94.340 148.685 94.600 149.140 ;
        RECT 94.770 148.855 95.030 149.335 ;
        RECT 95.200 148.685 95.460 149.140 ;
        RECT 95.630 148.855 95.890 149.335 ;
        RECT 96.060 148.685 96.320 149.140 ;
        RECT 96.490 148.775 96.750 149.335 ;
        RECT 89.575 148.515 96.320 148.685 ;
        RECT 88.145 146.785 88.375 147.925 ;
        RECT 88.545 146.955 88.875 147.935 ;
        RECT 89.575 147.925 90.740 148.515 ;
        RECT 96.920 148.345 97.170 149.155 ;
        RECT 97.350 148.810 97.610 149.335 ;
        RECT 97.780 148.345 98.030 149.155 ;
        RECT 98.210 148.825 98.515 149.335 ;
        RECT 90.910 148.095 98.030 148.345 ;
        RECT 98.200 148.095 98.515 148.655 ;
        RECT 98.685 148.585 99.895 149.335 ;
        RECT 100.065 148.610 100.355 149.335 ;
        RECT 100.575 148.680 100.905 149.115 ;
        RECT 101.075 148.725 101.245 149.335 ;
        RECT 100.525 148.595 100.905 148.680 ;
        RECT 101.415 148.595 101.745 149.120 ;
        RECT 102.005 148.805 102.215 149.335 ;
        RECT 102.490 148.885 103.275 149.055 ;
        RECT 103.445 148.885 103.850 149.055 ;
        RECT 89.045 146.785 89.255 147.925 ;
        RECT 89.575 147.700 96.320 147.925 ;
        RECT 89.575 146.785 89.845 147.530 ;
        RECT 90.015 146.960 90.305 147.700 ;
        RECT 90.915 147.685 96.320 147.700 ;
        RECT 90.475 146.790 90.730 147.515 ;
        RECT 90.915 146.960 91.175 147.685 ;
        RECT 91.345 146.790 91.590 147.515 ;
        RECT 91.775 146.960 92.035 147.685 ;
        RECT 92.205 146.790 92.450 147.515 ;
        RECT 92.635 146.960 92.895 147.685 ;
        RECT 93.065 146.790 93.310 147.515 ;
        RECT 93.480 146.960 93.740 147.685 ;
        RECT 93.910 146.790 94.170 147.515 ;
        RECT 94.340 146.960 94.600 147.685 ;
        RECT 94.770 146.790 95.030 147.515 ;
        RECT 95.200 146.960 95.460 147.685 ;
        RECT 95.630 146.790 95.890 147.515 ;
        RECT 96.060 146.960 96.320 147.685 ;
        RECT 96.490 146.790 96.750 147.585 ;
        RECT 96.920 146.960 97.170 148.095 ;
        RECT 90.475 146.785 96.750 146.790 ;
        RECT 97.350 146.785 97.610 147.595 ;
        RECT 97.785 146.955 98.030 148.095 ;
        RECT 98.685 148.045 99.205 148.585 ;
        RECT 100.525 148.555 100.750 148.595 ;
        RECT 99.375 147.875 99.895 148.415 ;
        RECT 100.525 147.975 100.695 148.555 ;
        RECT 101.415 148.425 101.615 148.595 ;
        RECT 102.490 148.425 102.660 148.885 ;
        RECT 100.865 148.095 101.615 148.425 ;
        RECT 101.785 148.095 102.660 148.425 ;
        RECT 98.210 146.785 98.505 147.595 ;
        RECT 98.685 146.785 99.895 147.875 ;
        RECT 100.065 146.785 100.355 147.950 ;
        RECT 100.525 147.925 100.740 147.975 ;
        RECT 100.525 147.845 100.915 147.925 ;
        RECT 100.585 147.000 100.915 147.845 ;
        RECT 101.425 147.890 101.615 148.095 ;
        RECT 101.085 146.785 101.255 147.795 ;
        RECT 101.425 147.515 102.320 147.890 ;
        RECT 101.425 146.955 101.765 147.515 ;
        RECT 101.995 146.785 102.310 147.285 ;
        RECT 102.490 147.255 102.660 148.095 ;
        RECT 102.830 148.385 103.295 148.715 ;
        RECT 103.680 148.655 103.850 148.885 ;
        RECT 104.030 148.835 104.400 149.335 ;
        RECT 104.720 148.885 105.395 149.055 ;
        RECT 105.590 148.885 105.925 149.055 ;
        RECT 102.830 147.425 103.150 148.385 ;
        RECT 103.680 148.355 104.510 148.655 ;
        RECT 103.320 147.455 103.510 148.175 ;
        RECT 103.680 147.285 103.850 148.355 ;
        RECT 104.310 148.325 104.510 148.355 ;
        RECT 104.020 148.105 104.190 148.175 ;
        RECT 104.720 148.105 104.890 148.885 ;
        RECT 105.755 148.745 105.925 148.885 ;
        RECT 106.095 148.875 106.345 149.335 ;
        RECT 104.020 147.935 104.890 148.105 ;
        RECT 105.060 148.465 105.585 148.685 ;
        RECT 105.755 148.615 105.980 148.745 ;
        RECT 104.020 147.845 104.530 147.935 ;
        RECT 102.490 147.085 103.375 147.255 ;
        RECT 103.600 146.955 103.850 147.285 ;
        RECT 104.020 146.785 104.190 147.585 ;
        RECT 104.360 147.230 104.530 147.845 ;
        RECT 105.060 147.765 105.230 148.465 ;
        RECT 104.700 147.400 105.230 147.765 ;
        RECT 105.400 147.700 105.640 148.295 ;
        RECT 105.810 147.510 105.980 148.615 ;
        RECT 106.150 147.755 106.430 148.705 ;
        RECT 105.675 147.380 105.980 147.510 ;
        RECT 104.360 147.060 105.465 147.230 ;
        RECT 105.675 146.955 105.925 147.380 ;
        RECT 106.095 146.785 106.360 147.245 ;
        RECT 106.600 146.955 106.785 149.075 ;
        RECT 106.955 148.955 107.285 149.335 ;
        RECT 107.455 148.785 107.625 149.075 ;
        RECT 106.960 148.615 107.625 148.785 ;
        RECT 107.975 148.785 108.145 149.075 ;
        RECT 108.315 148.955 108.645 149.335 ;
        RECT 107.975 148.615 108.640 148.785 ;
        RECT 106.960 147.625 107.190 148.615 ;
        RECT 107.360 147.795 107.710 148.445 ;
        RECT 107.890 147.795 108.240 148.445 ;
        RECT 108.410 147.625 108.640 148.615 ;
        RECT 106.960 147.455 107.625 147.625 ;
        RECT 106.955 146.785 107.285 147.285 ;
        RECT 107.455 146.955 107.625 147.455 ;
        RECT 107.975 147.455 108.640 147.625 ;
        RECT 107.975 146.955 108.145 147.455 ;
        RECT 108.315 146.785 108.645 147.285 ;
        RECT 108.815 146.955 109.000 149.075 ;
        RECT 109.255 148.875 109.505 149.335 ;
        RECT 109.675 148.885 110.010 149.055 ;
        RECT 110.205 148.885 110.880 149.055 ;
        RECT 109.675 148.745 109.845 148.885 ;
        RECT 109.170 147.755 109.450 148.705 ;
        RECT 109.620 148.615 109.845 148.745 ;
        RECT 109.620 147.510 109.790 148.615 ;
        RECT 110.015 148.465 110.540 148.685 ;
        RECT 109.960 147.700 110.200 148.295 ;
        RECT 110.370 147.765 110.540 148.465 ;
        RECT 110.710 148.105 110.880 148.885 ;
        RECT 111.200 148.835 111.570 149.335 ;
        RECT 111.750 148.885 112.155 149.055 ;
        RECT 112.325 148.885 113.110 149.055 ;
        RECT 111.750 148.655 111.920 148.885 ;
        RECT 111.090 148.355 111.920 148.655 ;
        RECT 112.305 148.385 112.770 148.715 ;
        RECT 111.090 148.325 111.290 148.355 ;
        RECT 111.410 148.105 111.580 148.175 ;
        RECT 110.710 147.935 111.580 148.105 ;
        RECT 111.070 147.845 111.580 147.935 ;
        RECT 109.620 147.380 109.925 147.510 ;
        RECT 110.370 147.400 110.900 147.765 ;
        RECT 109.240 146.785 109.505 147.245 ;
        RECT 109.675 146.955 109.925 147.380 ;
        RECT 111.070 147.230 111.240 147.845 ;
        RECT 110.135 147.060 111.240 147.230 ;
        RECT 111.410 146.785 111.580 147.585 ;
        RECT 111.750 147.285 111.920 148.355 ;
        RECT 112.090 147.455 112.280 148.175 ;
        RECT 112.450 147.425 112.770 148.385 ;
        RECT 112.940 148.425 113.110 148.885 ;
        RECT 113.385 148.805 113.595 149.335 ;
        RECT 113.855 148.595 114.185 149.120 ;
        RECT 114.355 148.725 114.525 149.335 ;
        RECT 114.695 148.680 115.025 149.115 ;
        RECT 116.165 148.825 116.470 149.335 ;
        RECT 114.695 148.595 115.075 148.680 ;
        RECT 113.985 148.425 114.185 148.595 ;
        RECT 114.850 148.555 115.075 148.595 ;
        RECT 112.940 148.095 113.815 148.425 ;
        RECT 113.985 148.095 114.735 148.425 ;
        RECT 111.750 146.955 112.000 147.285 ;
        RECT 112.940 147.255 113.110 148.095 ;
        RECT 113.985 147.890 114.175 148.095 ;
        RECT 114.905 147.975 115.075 148.555 ;
        RECT 116.165 148.095 116.480 148.655 ;
        RECT 116.650 148.345 116.900 149.155 ;
        RECT 117.070 148.810 117.330 149.335 ;
        RECT 117.510 148.345 117.760 149.155 ;
        RECT 117.930 148.775 118.190 149.335 ;
        RECT 118.360 148.685 118.620 149.140 ;
        RECT 118.790 148.855 119.050 149.335 ;
        RECT 119.220 148.685 119.480 149.140 ;
        RECT 119.650 148.855 119.910 149.335 ;
        RECT 120.080 148.685 120.340 149.140 ;
        RECT 120.510 148.855 120.755 149.335 ;
        RECT 120.925 148.685 121.200 149.140 ;
        RECT 121.370 148.855 121.615 149.335 ;
        RECT 121.785 148.685 122.045 149.140 ;
        RECT 122.225 148.855 122.475 149.335 ;
        RECT 122.645 148.685 122.905 149.140 ;
        RECT 123.085 148.855 123.335 149.335 ;
        RECT 123.505 148.685 123.765 149.140 ;
        RECT 123.945 148.855 124.205 149.335 ;
        RECT 124.375 148.685 124.635 149.140 ;
        RECT 124.805 148.855 125.105 149.335 ;
        RECT 118.360 148.515 125.105 148.685 ;
        RECT 125.825 148.610 126.115 149.335 ;
        RECT 126.285 148.835 126.545 149.165 ;
        RECT 126.715 148.975 127.045 149.335 ;
        RECT 127.300 148.955 128.600 149.165 ;
        RECT 116.650 148.095 123.770 148.345 ;
        RECT 114.860 147.925 115.075 147.975 ;
        RECT 113.280 147.515 114.175 147.890 ;
        RECT 114.685 147.845 115.075 147.925 ;
        RECT 112.225 147.085 113.110 147.255 ;
        RECT 113.290 146.785 113.605 147.285 ;
        RECT 113.835 146.955 114.175 147.515 ;
        RECT 114.345 146.785 114.515 147.795 ;
        RECT 114.685 147.000 115.015 147.845 ;
        RECT 116.175 146.785 116.470 147.595 ;
        RECT 116.650 146.955 116.895 148.095 ;
        RECT 117.070 146.785 117.330 147.595 ;
        RECT 117.510 146.960 117.760 148.095 ;
        RECT 123.940 147.925 125.105 148.515 ;
        RECT 118.360 147.700 125.105 147.925 ;
        RECT 118.360 147.685 123.765 147.700 ;
        RECT 117.930 146.790 118.190 147.585 ;
        RECT 118.360 146.960 118.620 147.685 ;
        RECT 118.790 146.790 119.050 147.515 ;
        RECT 119.220 146.960 119.480 147.685 ;
        RECT 119.650 146.790 119.910 147.515 ;
        RECT 120.080 146.960 120.340 147.685 ;
        RECT 120.510 146.790 120.770 147.515 ;
        RECT 120.940 146.960 121.200 147.685 ;
        RECT 121.370 146.790 121.615 147.515 ;
        RECT 121.785 146.960 122.045 147.685 ;
        RECT 122.230 146.790 122.475 147.515 ;
        RECT 122.645 146.960 122.905 147.685 ;
        RECT 123.090 146.790 123.335 147.515 ;
        RECT 123.505 146.960 123.765 147.685 ;
        RECT 123.950 146.790 124.205 147.515 ;
        RECT 124.375 146.960 124.665 147.700 ;
        RECT 117.930 146.785 124.205 146.790 ;
        RECT 124.835 146.785 125.105 147.530 ;
        RECT 125.825 146.785 126.115 147.950 ;
        RECT 126.285 147.635 126.455 148.835 ;
        RECT 127.300 148.805 127.470 148.955 ;
        RECT 126.715 148.680 127.470 148.805 ;
        RECT 126.625 148.635 127.470 148.680 ;
        RECT 126.625 148.515 126.895 148.635 ;
        RECT 126.625 147.940 126.795 148.515 ;
        RECT 127.025 148.075 127.435 148.380 ;
        RECT 127.725 148.345 127.935 148.745 ;
        RECT 127.605 148.135 127.935 148.345 ;
        RECT 128.180 148.345 128.400 148.745 ;
        RECT 128.875 148.570 129.330 149.335 ;
        RECT 129.505 148.835 129.765 149.165 ;
        RECT 129.935 148.975 130.265 149.335 ;
        RECT 130.520 148.955 131.820 149.165 ;
        RECT 129.505 148.825 129.735 148.835 ;
        RECT 128.180 148.135 128.655 148.345 ;
        RECT 128.845 148.145 129.335 148.345 ;
        RECT 126.625 147.905 126.825 147.940 ;
        RECT 128.155 147.905 129.330 147.965 ;
        RECT 126.625 147.795 129.330 147.905 ;
        RECT 126.685 147.735 128.485 147.795 ;
        RECT 128.155 147.705 128.485 147.735 ;
        RECT 126.285 146.955 126.545 147.635 ;
        RECT 126.715 146.785 126.965 147.565 ;
        RECT 127.215 147.535 128.050 147.545 ;
        RECT 128.640 147.535 128.825 147.625 ;
        RECT 127.215 147.335 128.825 147.535 ;
        RECT 127.215 146.955 127.465 147.335 ;
        RECT 128.595 147.295 128.825 147.335 ;
        RECT 129.075 147.175 129.330 147.795 ;
        RECT 127.635 146.785 127.990 147.165 ;
        RECT 128.995 146.955 129.330 147.175 ;
        RECT 129.505 147.635 129.675 148.825 ;
        RECT 130.520 148.805 130.690 148.955 ;
        RECT 129.935 148.680 130.690 148.805 ;
        RECT 129.845 148.635 130.690 148.680 ;
        RECT 129.845 148.515 130.115 148.635 ;
        RECT 129.845 147.940 130.015 148.515 ;
        RECT 130.245 148.075 130.655 148.380 ;
        RECT 130.945 148.345 131.155 148.745 ;
        RECT 130.825 148.135 131.155 148.345 ;
        RECT 131.400 148.345 131.620 148.745 ;
        RECT 132.095 148.570 132.550 149.335 ;
        RECT 132.925 148.705 133.255 149.065 ;
        RECT 133.875 148.875 134.125 149.335 ;
        RECT 134.295 148.875 134.855 149.165 ;
        RECT 132.925 148.515 134.315 148.705 ;
        RECT 134.145 148.425 134.315 148.515 ;
        RECT 131.400 148.135 131.875 148.345 ;
        RECT 132.065 148.145 132.555 148.345 ;
        RECT 132.740 148.095 133.415 148.345 ;
        RECT 133.635 148.095 133.975 148.345 ;
        RECT 134.145 148.095 134.435 148.425 ;
        RECT 129.845 147.905 130.045 147.940 ;
        RECT 131.375 147.905 132.550 147.965 ;
        RECT 129.845 147.795 132.550 147.905 ;
        RECT 129.905 147.735 131.705 147.795 ;
        RECT 131.375 147.705 131.705 147.735 ;
        RECT 129.505 146.955 129.765 147.635 ;
        RECT 129.935 146.785 130.185 147.565 ;
        RECT 130.435 147.535 131.270 147.545 ;
        RECT 131.860 147.535 132.045 147.625 ;
        RECT 130.435 147.335 132.045 147.535 ;
        RECT 130.435 146.955 130.685 147.335 ;
        RECT 131.815 147.295 132.045 147.335 ;
        RECT 132.295 147.175 132.550 147.795 ;
        RECT 132.740 147.735 133.005 148.095 ;
        RECT 134.145 147.845 134.315 148.095 ;
        RECT 133.375 147.675 134.315 147.845 ;
        RECT 130.855 146.785 131.210 147.165 ;
        RECT 132.215 146.955 132.550 147.175 ;
        RECT 132.925 146.785 133.205 147.455 ;
        RECT 133.375 147.125 133.675 147.675 ;
        RECT 134.605 147.505 134.855 148.875 ;
        RECT 135.085 148.515 135.295 149.335 ;
        RECT 135.465 148.535 135.795 149.165 ;
        RECT 135.465 147.935 135.715 148.535 ;
        RECT 135.965 148.515 136.195 149.335 ;
        RECT 136.405 148.790 141.750 149.335 ;
        RECT 141.925 148.790 147.270 149.335 ;
        RECT 135.885 148.095 136.215 148.345 ;
        RECT 137.990 147.960 138.330 148.790 ;
        RECT 133.875 146.785 134.205 147.505 ;
        RECT 134.395 146.955 134.855 147.505 ;
        RECT 135.085 146.785 135.295 147.925 ;
        RECT 135.465 146.955 135.795 147.935 ;
        RECT 135.965 146.785 136.195 147.925 ;
        RECT 139.810 147.220 140.160 148.470 ;
        RECT 143.510 147.960 143.850 148.790 ;
        RECT 147.995 148.785 148.165 149.165 ;
        RECT 148.345 148.955 148.675 149.335 ;
        RECT 147.995 148.615 148.660 148.785 ;
        RECT 148.855 148.660 149.115 149.165 ;
        RECT 145.330 147.220 145.680 148.470 ;
        RECT 147.925 148.065 148.255 148.435 ;
        RECT 148.490 148.360 148.660 148.615 ;
        RECT 148.490 148.030 148.775 148.360 ;
        RECT 148.490 147.885 148.660 148.030 ;
        RECT 147.995 147.715 148.660 147.885 ;
        RECT 148.945 147.860 149.115 148.660 ;
        RECT 149.285 148.565 150.955 149.335 ;
        RECT 151.585 148.610 151.875 149.335 ;
        RECT 152.045 148.565 155.555 149.335 ;
        RECT 155.725 148.585 156.935 149.335 ;
        RECT 149.285 148.045 150.035 148.565 ;
        RECT 150.205 147.875 150.955 148.395 ;
        RECT 152.045 148.045 153.695 148.565 ;
        RECT 136.405 146.785 141.750 147.220 ;
        RECT 141.925 146.785 147.270 147.220 ;
        RECT 147.995 146.955 148.165 147.715 ;
        RECT 148.345 146.785 148.675 147.545 ;
        RECT 148.845 146.955 149.115 147.860 ;
        RECT 149.285 146.785 150.955 147.875 ;
        RECT 151.585 146.785 151.875 147.950 ;
        RECT 153.865 147.875 155.555 148.395 ;
        RECT 152.045 146.785 155.555 147.875 ;
        RECT 155.725 147.875 156.245 148.415 ;
        RECT 156.415 148.045 156.935 148.585 ;
        RECT 155.725 146.785 156.935 147.875 ;
        RECT 22.700 146.615 157.020 146.785 ;
        RECT 22.785 145.525 23.995 146.615 ;
        RECT 24.165 145.525 25.375 146.615 ;
        RECT 22.785 144.815 23.305 145.355 ;
        RECT 23.475 144.985 23.995 145.525 ;
        RECT 24.165 144.815 24.685 145.355 ;
        RECT 24.855 144.985 25.375 145.525 ;
        RECT 25.545 145.540 25.815 146.445 ;
        RECT 25.985 145.855 26.315 146.615 ;
        RECT 26.495 145.685 26.665 146.445 ;
        RECT 22.785 144.065 23.995 144.815 ;
        RECT 24.165 144.065 25.375 144.815 ;
        RECT 25.545 144.740 25.715 145.540 ;
        RECT 26.000 145.515 26.665 145.685 ;
        RECT 26.925 145.525 28.595 146.615 ;
        RECT 26.000 145.370 26.170 145.515 ;
        RECT 25.885 145.040 26.170 145.370 ;
        RECT 26.000 144.785 26.170 145.040 ;
        RECT 26.405 144.965 26.735 145.335 ;
        RECT 26.925 144.835 27.675 145.355 ;
        RECT 27.845 145.005 28.595 145.525 ;
        RECT 29.225 145.895 29.685 146.445 ;
        RECT 29.875 145.895 30.205 146.615 ;
        RECT 25.545 144.235 25.805 144.740 ;
        RECT 26.000 144.615 26.665 144.785 ;
        RECT 25.985 144.065 26.315 144.445 ;
        RECT 26.495 144.235 26.665 144.615 ;
        RECT 26.925 144.065 28.595 144.835 ;
        RECT 29.225 144.525 29.475 145.895 ;
        RECT 30.405 145.725 30.705 146.275 ;
        RECT 30.875 145.945 31.155 146.615 ;
        RECT 29.765 145.555 30.705 145.725 ;
        RECT 31.560 145.825 32.095 146.445 ;
        RECT 29.765 145.305 29.935 145.555 ;
        RECT 31.075 145.305 31.340 145.665 ;
        RECT 29.645 144.975 29.935 145.305 ;
        RECT 30.105 145.055 30.445 145.305 ;
        RECT 30.665 145.055 31.340 145.305 ;
        RECT 29.765 144.885 29.935 144.975 ;
        RECT 29.765 144.695 31.155 144.885 ;
        RECT 29.225 144.235 29.785 144.525 ;
        RECT 29.955 144.065 30.205 144.525 ;
        RECT 30.825 144.335 31.155 144.695 ;
        RECT 31.560 144.805 31.875 145.825 ;
        RECT 32.265 145.815 32.595 146.615 ;
        RECT 33.080 145.645 33.470 145.820 ;
        RECT 32.045 145.475 33.470 145.645 ;
        RECT 33.825 145.525 35.495 146.615 ;
        RECT 32.045 144.975 32.215 145.475 ;
        RECT 31.560 144.235 32.175 144.805 ;
        RECT 32.465 144.745 32.730 145.305 ;
        RECT 32.900 144.575 33.070 145.475 ;
        RECT 33.240 144.745 33.595 145.305 ;
        RECT 33.825 144.835 34.575 145.355 ;
        RECT 34.745 145.005 35.495 145.525 ;
        RECT 35.665 145.450 35.955 146.615 ;
        RECT 36.125 146.180 41.470 146.615 ;
        RECT 32.345 144.065 32.560 144.575 ;
        RECT 32.790 144.245 33.070 144.575 ;
        RECT 33.250 144.065 33.490 144.575 ;
        RECT 33.825 144.065 35.495 144.835 ;
        RECT 35.665 144.065 35.955 144.790 ;
        RECT 37.710 144.610 38.050 145.440 ;
        RECT 39.530 144.930 39.880 146.180 ;
        RECT 42.565 145.815 42.890 146.615 ;
        RECT 42.585 145.055 42.915 145.640 ;
        RECT 43.085 145.305 43.270 146.395 ;
        RECT 43.440 145.645 43.690 146.445 ;
        RECT 43.860 145.815 44.600 146.615 ;
        RECT 44.785 145.645 45.115 146.445 ;
        RECT 45.285 145.815 46.095 146.615 ;
        RECT 43.440 145.475 45.925 145.645 ;
        RECT 45.755 145.305 45.925 145.475 ;
        RECT 43.085 145.055 43.570 145.305 ;
        RECT 43.915 144.975 44.175 145.305 ;
        RECT 42.565 144.685 43.750 144.855 ;
        RECT 36.125 144.065 41.470 144.610 ;
        RECT 42.565 144.235 42.830 144.685 ;
        RECT 43.000 144.065 43.290 144.515 ;
        RECT 43.460 144.235 43.750 144.685 ;
        RECT 43.930 144.370 44.175 144.975 ;
        RECT 44.425 144.370 44.695 145.305 ;
        RECT 44.875 145.055 45.355 145.305 ;
        RECT 44.875 144.370 45.085 145.055 ;
        RECT 45.755 144.975 46.095 145.305 ;
        RECT 45.755 144.885 45.925 144.975 ;
        RECT 45.255 144.715 45.925 144.885 ;
        RECT 45.255 144.235 45.595 144.715 ;
        RECT 45.775 144.065 46.085 144.545 ;
        RECT 46.265 144.235 46.525 146.445 ;
        RECT 47.255 145.605 47.425 146.445 ;
        RECT 47.595 146.275 48.765 146.445 ;
        RECT 47.595 145.775 47.925 146.275 ;
        RECT 48.435 146.235 48.765 146.275 ;
        RECT 48.955 146.195 49.310 146.615 ;
        RECT 48.095 146.015 48.325 146.105 ;
        RECT 49.480 146.015 49.730 146.445 ;
        RECT 48.095 145.775 49.730 146.015 ;
        RECT 49.900 145.855 50.230 146.615 ;
        RECT 50.400 145.775 50.655 146.445 ;
        RECT 47.255 145.435 50.315 145.605 ;
        RECT 47.170 145.055 47.520 145.265 ;
        RECT 47.690 145.055 48.135 145.255 ;
        RECT 48.305 145.055 48.780 145.255 ;
        RECT 47.255 144.715 48.320 144.885 ;
        RECT 47.255 144.235 47.425 144.715 ;
        RECT 47.595 144.065 47.925 144.545 ;
        RECT 48.150 144.485 48.320 144.715 ;
        RECT 48.500 144.655 48.780 145.055 ;
        RECT 49.050 145.055 49.380 145.255 ;
        RECT 49.550 145.085 49.925 145.255 ;
        RECT 49.550 145.055 49.915 145.085 ;
        RECT 49.050 144.655 49.335 145.055 ;
        RECT 50.145 144.885 50.315 145.435 ;
        RECT 49.515 144.715 50.315 144.885 ;
        RECT 49.515 144.485 49.685 144.715 ;
        RECT 50.485 144.645 50.655 145.775 ;
        RECT 50.905 145.475 51.115 146.615 ;
        RECT 51.285 145.465 51.615 146.445 ;
        RECT 51.785 145.475 52.015 146.615 ;
        RECT 52.265 145.475 52.495 146.615 ;
        RECT 52.665 145.465 52.995 146.445 ;
        RECT 53.165 145.475 53.375 146.615 ;
        RECT 53.605 145.525 56.195 146.615 ;
        RECT 50.470 144.565 50.655 144.645 ;
        RECT 48.150 144.235 49.685 144.485 ;
        RECT 49.855 144.065 50.185 144.545 ;
        RECT 50.400 144.235 50.655 144.565 ;
        RECT 50.905 144.065 51.115 144.885 ;
        RECT 51.285 144.865 51.535 145.465 ;
        RECT 51.705 145.055 52.035 145.305 ;
        RECT 52.245 145.055 52.575 145.305 ;
        RECT 51.285 144.235 51.615 144.865 ;
        RECT 51.785 144.065 52.015 144.885 ;
        RECT 52.265 144.065 52.495 144.885 ;
        RECT 52.745 144.865 52.995 145.465 ;
        RECT 52.665 144.235 52.995 144.865 ;
        RECT 53.165 144.065 53.375 144.885 ;
        RECT 53.605 144.835 54.815 145.355 ;
        RECT 54.985 145.005 56.195 145.525 ;
        RECT 53.605 144.065 56.195 144.835 ;
        RECT 56.375 144.245 56.635 146.435 ;
        RECT 56.805 145.885 57.145 146.615 ;
        RECT 57.325 145.705 57.595 146.435 ;
        RECT 56.825 145.485 57.595 145.705 ;
        RECT 57.775 145.725 58.005 146.435 ;
        RECT 58.175 145.905 58.505 146.615 ;
        RECT 58.675 145.725 58.935 146.435 ;
        RECT 57.775 145.485 58.935 145.725 ;
        RECT 59.125 145.525 60.795 146.615 ;
        RECT 56.825 144.815 57.115 145.485 ;
        RECT 57.295 144.995 57.760 145.305 ;
        RECT 57.940 144.995 58.465 145.305 ;
        RECT 56.825 144.615 58.055 144.815 ;
        RECT 56.895 144.065 57.565 144.435 ;
        RECT 57.745 144.245 58.055 144.615 ;
        RECT 58.235 144.355 58.465 144.995 ;
        RECT 58.645 144.975 58.945 145.305 ;
        RECT 59.125 144.835 59.875 145.355 ;
        RECT 60.045 145.005 60.795 145.525 ;
        RECT 61.425 145.450 61.715 146.615 ;
        RECT 58.645 144.065 58.935 144.795 ;
        RECT 59.125 144.065 60.795 144.835 ;
        RECT 61.425 144.065 61.715 144.790 ;
        RECT 62.815 144.245 63.075 146.435 ;
        RECT 63.245 145.885 63.585 146.615 ;
        RECT 63.765 145.705 64.035 146.435 ;
        RECT 63.265 145.485 64.035 145.705 ;
        RECT 64.215 145.725 64.445 146.435 ;
        RECT 64.615 145.905 64.945 146.615 ;
        RECT 65.115 145.725 65.375 146.435 ;
        RECT 64.215 145.485 65.375 145.725 ;
        RECT 66.035 145.505 66.330 146.615 ;
        RECT 63.265 144.815 63.555 145.485 ;
        RECT 66.510 145.305 66.760 146.440 ;
        RECT 66.930 145.505 67.190 146.615 ;
        RECT 67.360 145.715 67.620 146.440 ;
        RECT 67.790 145.885 68.050 146.615 ;
        RECT 68.220 145.715 68.480 146.440 ;
        RECT 68.650 145.885 68.910 146.615 ;
        RECT 69.080 145.715 69.340 146.440 ;
        RECT 69.510 145.885 69.770 146.615 ;
        RECT 69.940 145.715 70.200 146.440 ;
        RECT 70.370 145.885 70.665 146.615 ;
        RECT 71.175 145.945 71.345 146.445 ;
        RECT 71.515 146.115 71.845 146.615 ;
        RECT 71.175 145.775 71.840 145.945 ;
        RECT 67.360 145.475 70.670 145.715 ;
        RECT 63.735 144.995 64.200 145.305 ;
        RECT 64.380 144.995 64.905 145.305 ;
        RECT 63.265 144.615 64.495 144.815 ;
        RECT 63.335 144.065 64.005 144.435 ;
        RECT 64.185 144.245 64.495 144.615 ;
        RECT 64.675 144.355 64.905 144.995 ;
        RECT 65.085 144.975 65.385 145.305 ;
        RECT 65.085 144.065 65.375 144.795 ;
        RECT 66.025 144.695 66.340 145.305 ;
        RECT 66.510 145.055 69.530 145.305 ;
        RECT 66.085 144.065 66.330 144.525 ;
        RECT 66.510 144.245 66.760 145.055 ;
        RECT 69.700 144.885 70.670 145.475 ;
        RECT 71.090 144.955 71.440 145.605 ;
        RECT 67.360 144.715 70.670 144.885 ;
        RECT 71.610 144.785 71.840 145.775 ;
        RECT 66.930 144.065 67.190 144.590 ;
        RECT 67.360 144.260 67.620 144.715 ;
        RECT 67.790 144.065 68.050 144.545 ;
        RECT 68.220 144.260 68.480 144.715 ;
        RECT 68.650 144.065 68.910 144.545 ;
        RECT 69.080 144.260 69.340 144.715 ;
        RECT 69.510 144.065 69.770 144.545 ;
        RECT 69.940 144.260 70.200 144.715 ;
        RECT 71.175 144.615 71.840 144.785 ;
        RECT 70.370 144.065 70.670 144.545 ;
        RECT 71.175 144.325 71.345 144.615 ;
        RECT 71.515 144.065 71.845 144.445 ;
        RECT 72.015 144.325 72.200 146.445 ;
        RECT 72.440 146.155 72.705 146.615 ;
        RECT 72.875 146.020 73.125 146.445 ;
        RECT 73.335 146.170 74.440 146.340 ;
        RECT 72.820 145.890 73.125 146.020 ;
        RECT 72.370 144.695 72.650 145.645 ;
        RECT 72.820 144.785 72.990 145.890 ;
        RECT 73.160 145.105 73.400 145.700 ;
        RECT 73.570 145.635 74.100 146.000 ;
        RECT 73.570 144.935 73.740 145.635 ;
        RECT 74.270 145.555 74.440 146.170 ;
        RECT 74.610 145.815 74.780 146.615 ;
        RECT 74.950 146.115 75.200 146.445 ;
        RECT 75.425 146.145 76.310 146.315 ;
        RECT 74.270 145.465 74.780 145.555 ;
        RECT 72.820 144.655 73.045 144.785 ;
        RECT 73.215 144.715 73.740 144.935 ;
        RECT 73.910 145.295 74.780 145.465 ;
        RECT 72.455 144.065 72.705 144.525 ;
        RECT 72.875 144.515 73.045 144.655 ;
        RECT 73.910 144.515 74.080 145.295 ;
        RECT 74.610 145.225 74.780 145.295 ;
        RECT 74.290 145.045 74.490 145.075 ;
        RECT 74.950 145.045 75.120 146.115 ;
        RECT 75.290 145.225 75.480 145.945 ;
        RECT 74.290 144.745 75.120 145.045 ;
        RECT 75.650 145.015 75.970 145.975 ;
        RECT 72.875 144.345 73.210 144.515 ;
        RECT 73.405 144.345 74.080 144.515 ;
        RECT 74.400 144.065 74.770 144.565 ;
        RECT 74.950 144.515 75.120 144.745 ;
        RECT 75.505 144.685 75.970 145.015 ;
        RECT 76.140 145.305 76.310 146.145 ;
        RECT 76.490 146.115 76.805 146.615 ;
        RECT 77.035 145.885 77.375 146.445 ;
        RECT 76.480 145.510 77.375 145.885 ;
        RECT 77.545 145.605 77.715 146.615 ;
        RECT 77.185 145.305 77.375 145.510 ;
        RECT 77.885 145.555 78.215 146.400 ;
        RECT 77.885 145.475 78.275 145.555 ;
        RECT 78.060 145.425 78.275 145.475 ;
        RECT 76.140 144.975 77.015 145.305 ;
        RECT 77.185 144.975 77.935 145.305 ;
        RECT 76.140 144.515 76.310 144.975 ;
        RECT 77.185 144.805 77.385 144.975 ;
        RECT 78.105 144.845 78.275 145.425 ;
        RECT 78.050 144.805 78.275 144.845 ;
        RECT 74.950 144.345 75.355 144.515 ;
        RECT 75.525 144.345 76.310 144.515 ;
        RECT 76.585 144.065 76.795 144.595 ;
        RECT 77.055 144.280 77.385 144.805 ;
        RECT 77.895 144.720 78.275 144.805 ;
        RECT 78.450 145.475 78.785 146.445 ;
        RECT 78.955 145.475 79.125 146.615 ;
        RECT 79.295 146.275 81.325 146.445 ;
        RECT 78.450 144.805 78.620 145.475 ;
        RECT 79.295 145.305 79.465 146.275 ;
        RECT 78.790 144.975 79.045 145.305 ;
        RECT 79.270 144.975 79.465 145.305 ;
        RECT 79.635 145.935 80.760 146.105 ;
        RECT 78.875 144.805 79.045 144.975 ;
        RECT 79.635 144.805 79.805 145.935 ;
        RECT 77.555 144.065 77.725 144.675 ;
        RECT 77.895 144.285 78.225 144.720 ;
        RECT 78.450 144.235 78.705 144.805 ;
        RECT 78.875 144.635 79.805 144.805 ;
        RECT 79.975 145.595 80.985 145.765 ;
        RECT 79.975 144.795 80.145 145.595 ;
        RECT 79.630 144.600 79.805 144.635 ;
        RECT 78.875 144.065 79.205 144.465 ;
        RECT 79.630 144.235 80.160 144.600 ;
        RECT 80.350 144.575 80.625 145.395 ;
        RECT 80.345 144.405 80.625 144.575 ;
        RECT 80.350 144.235 80.625 144.405 ;
        RECT 80.795 144.235 80.985 145.595 ;
        RECT 81.155 145.610 81.325 146.275 ;
        RECT 81.495 145.855 81.665 146.615 ;
        RECT 81.900 145.855 82.415 146.265 ;
        RECT 81.155 145.420 81.905 145.610 ;
        RECT 82.075 145.045 82.415 145.855 ;
        RECT 82.585 145.525 85.175 146.615 ;
        RECT 81.185 144.875 82.415 145.045 ;
        RECT 81.165 144.065 81.675 144.600 ;
        RECT 81.895 144.270 82.140 144.875 ;
        RECT 82.585 144.835 83.795 145.355 ;
        RECT 83.965 145.005 85.175 145.525 ;
        RECT 85.865 145.475 86.075 146.615 ;
        RECT 86.245 145.465 86.575 146.445 ;
        RECT 86.745 145.475 86.975 146.615 ;
        RECT 82.585 144.065 85.175 144.835 ;
        RECT 85.865 144.065 86.075 144.885 ;
        RECT 86.245 144.865 86.495 145.465 ;
        RECT 87.185 145.450 87.475 146.615 ;
        RECT 88.105 145.745 88.380 146.445 ;
        RECT 88.550 146.070 88.805 146.615 ;
        RECT 88.975 146.105 89.455 146.445 ;
        RECT 89.630 146.060 90.235 146.615 ;
        RECT 89.620 145.960 90.235 146.060 ;
        RECT 89.620 145.935 89.805 145.960 ;
        RECT 86.665 145.055 86.995 145.305 ;
        RECT 86.245 144.235 86.575 144.865 ;
        RECT 86.745 144.065 86.975 144.885 ;
        RECT 87.185 144.065 87.475 144.790 ;
        RECT 88.105 144.715 88.275 145.745 ;
        RECT 88.550 145.615 89.305 145.865 ;
        RECT 89.475 145.690 89.805 145.935 ;
        RECT 88.550 145.580 89.320 145.615 ;
        RECT 88.550 145.570 89.335 145.580 ;
        RECT 88.445 145.555 89.340 145.570 ;
        RECT 88.445 145.540 89.360 145.555 ;
        RECT 88.445 145.530 89.380 145.540 ;
        RECT 88.445 145.520 89.405 145.530 ;
        RECT 88.445 145.490 89.475 145.520 ;
        RECT 88.445 145.460 89.495 145.490 ;
        RECT 88.445 145.430 89.515 145.460 ;
        RECT 88.445 145.405 89.545 145.430 ;
        RECT 88.445 145.370 89.580 145.405 ;
        RECT 88.445 145.365 89.610 145.370 ;
        RECT 88.445 144.970 88.675 145.365 ;
        RECT 89.220 145.360 89.610 145.365 ;
        RECT 89.245 145.350 89.610 145.360 ;
        RECT 89.260 145.345 89.610 145.350 ;
        RECT 89.275 145.340 89.610 145.345 ;
        RECT 89.975 145.340 90.235 145.790 ;
        RECT 89.275 145.335 90.235 145.340 ;
        RECT 89.285 145.325 90.235 145.335 ;
        RECT 89.295 145.320 90.235 145.325 ;
        RECT 89.305 145.310 90.235 145.320 ;
        RECT 89.310 145.300 90.235 145.310 ;
        RECT 89.315 145.295 90.235 145.300 ;
        RECT 89.325 145.280 90.235 145.295 ;
        RECT 89.330 145.265 90.235 145.280 ;
        RECT 89.340 145.240 90.235 145.265 ;
        RECT 88.845 144.770 89.175 145.195 ;
        RECT 88.925 144.745 89.175 144.770 ;
        RECT 88.105 144.235 88.365 144.715 ;
        RECT 88.535 144.065 88.785 144.605 ;
        RECT 88.955 144.285 89.175 144.745 ;
        RECT 89.345 145.170 90.235 145.240 ;
        RECT 90.885 145.775 91.140 146.445 ;
        RECT 91.310 145.855 91.640 146.615 ;
        RECT 91.810 146.015 92.060 146.445 ;
        RECT 92.230 146.195 92.585 146.615 ;
        RECT 92.775 146.275 93.945 146.445 ;
        RECT 92.775 146.235 93.105 146.275 ;
        RECT 93.215 146.015 93.445 146.105 ;
        RECT 91.810 145.775 93.445 146.015 ;
        RECT 93.615 145.775 93.945 146.275 ;
        RECT 89.345 144.445 89.515 145.170 ;
        RECT 89.685 144.615 90.235 145.000 ;
        RECT 90.885 144.645 91.055 145.775 ;
        RECT 94.115 145.605 94.285 146.445 ;
        RECT 91.225 145.435 94.285 145.605 ;
        RECT 94.730 145.645 95.120 145.820 ;
        RECT 95.605 145.815 95.935 146.615 ;
        RECT 96.105 145.825 96.640 146.445 ;
        RECT 96.845 146.105 97.105 146.615 ;
        RECT 94.730 145.475 96.155 145.645 ;
        RECT 91.225 144.885 91.395 145.435 ;
        RECT 91.625 145.055 91.990 145.255 ;
        RECT 92.160 145.055 92.490 145.255 ;
        RECT 91.225 144.715 92.025 144.885 ;
        RECT 90.885 144.575 91.070 144.645 ;
        RECT 90.885 144.565 91.095 144.575 ;
        RECT 89.345 144.275 90.235 144.445 ;
        RECT 90.885 144.235 91.140 144.565 ;
        RECT 91.355 144.065 91.685 144.545 ;
        RECT 91.855 144.485 92.025 144.715 ;
        RECT 92.205 144.655 92.490 145.055 ;
        RECT 92.760 145.055 93.235 145.255 ;
        RECT 93.405 145.055 93.850 145.255 ;
        RECT 94.020 145.055 94.370 145.265 ;
        RECT 92.760 144.655 93.040 145.055 ;
        RECT 93.220 144.715 94.285 144.885 ;
        RECT 94.605 144.745 94.960 145.305 ;
        RECT 93.220 144.485 93.390 144.715 ;
        RECT 91.855 144.235 93.390 144.485 ;
        RECT 93.615 144.065 93.945 144.545 ;
        RECT 94.115 144.235 94.285 144.715 ;
        RECT 95.130 144.575 95.300 145.475 ;
        RECT 95.470 144.745 95.735 145.305 ;
        RECT 95.985 144.975 96.155 145.475 ;
        RECT 96.325 144.805 96.640 145.825 ;
        RECT 96.845 145.055 97.185 145.935 ;
        RECT 97.355 145.225 97.525 146.445 ;
        RECT 97.765 146.110 98.380 146.615 ;
        RECT 97.765 145.575 98.015 145.940 ;
        RECT 98.185 145.935 98.380 146.110 ;
        RECT 98.550 146.105 99.025 146.445 ;
        RECT 99.195 146.070 99.410 146.615 ;
        RECT 98.185 145.745 98.515 145.935 ;
        RECT 98.735 145.575 99.450 145.870 ;
        RECT 99.620 145.745 99.895 146.445 ;
        RECT 97.765 145.405 99.555 145.575 ;
        RECT 97.355 144.975 98.150 145.225 ;
        RECT 97.355 144.885 97.605 144.975 ;
        RECT 94.710 144.065 94.950 144.575 ;
        RECT 95.130 144.245 95.410 144.575 ;
        RECT 95.640 144.065 95.855 144.575 ;
        RECT 96.025 144.235 96.640 144.805 ;
        RECT 96.845 144.065 97.105 144.885 ;
        RECT 97.275 144.465 97.605 144.885 ;
        RECT 98.320 144.550 98.575 145.405 ;
        RECT 97.785 144.285 98.575 144.550 ;
        RECT 98.745 144.705 99.155 145.225 ;
        RECT 99.325 144.975 99.555 145.405 ;
        RECT 99.725 144.715 99.895 145.745 ;
        RECT 100.250 145.645 100.640 145.820 ;
        RECT 101.125 145.815 101.455 146.615 ;
        RECT 101.625 145.825 102.160 146.445 ;
        RECT 100.250 145.475 101.675 145.645 ;
        RECT 100.125 144.745 100.480 145.305 ;
        RECT 98.745 144.285 98.945 144.705 ;
        RECT 99.135 144.065 99.465 144.525 ;
        RECT 99.635 144.235 99.895 144.715 ;
        RECT 100.650 144.575 100.820 145.475 ;
        RECT 100.990 144.745 101.255 145.305 ;
        RECT 101.505 144.975 101.675 145.475 ;
        RECT 101.845 144.805 102.160 145.825 ;
        RECT 102.455 145.685 102.625 146.445 ;
        RECT 102.805 145.855 103.135 146.615 ;
        RECT 102.455 145.515 103.120 145.685 ;
        RECT 103.305 145.540 103.575 146.445 ;
        RECT 104.260 145.745 104.545 146.615 ;
        RECT 104.715 145.985 104.975 146.445 ;
        RECT 105.150 146.155 105.405 146.615 ;
        RECT 105.575 145.985 105.835 146.445 ;
        RECT 104.715 145.815 105.835 145.985 ;
        RECT 106.005 145.815 106.315 146.615 ;
        RECT 104.715 145.565 104.975 145.815 ;
        RECT 106.485 145.645 106.795 146.445 ;
        RECT 102.950 145.370 103.120 145.515 ;
        RECT 102.385 144.965 102.715 145.335 ;
        RECT 102.950 145.040 103.235 145.370 ;
        RECT 100.230 144.065 100.470 144.575 ;
        RECT 100.650 144.245 100.930 144.575 ;
        RECT 101.160 144.065 101.375 144.575 ;
        RECT 101.545 144.235 102.160 144.805 ;
        RECT 102.950 144.785 103.120 145.040 ;
        RECT 102.455 144.615 103.120 144.785 ;
        RECT 103.405 144.740 103.575 145.540 ;
        RECT 102.455 144.235 102.625 144.615 ;
        RECT 102.805 144.065 103.135 144.445 ;
        RECT 103.315 144.235 103.575 144.740 ;
        RECT 104.220 145.395 104.975 145.565 ;
        RECT 105.765 145.475 106.795 145.645 ;
        RECT 104.220 144.885 104.625 145.395 ;
        RECT 105.765 145.225 105.935 145.475 ;
        RECT 104.795 145.055 105.935 145.225 ;
        RECT 104.220 144.715 105.870 144.885 ;
        RECT 106.105 144.735 106.455 145.305 ;
        RECT 104.265 144.065 104.545 144.545 ;
        RECT 104.715 144.325 104.975 144.715 ;
        RECT 105.150 144.065 105.405 144.545 ;
        RECT 105.575 144.325 105.870 144.715 ;
        RECT 106.625 144.565 106.795 145.475 ;
        RECT 106.050 144.065 106.325 144.545 ;
        RECT 106.495 144.235 106.795 144.565 ;
        RECT 106.965 145.765 107.225 146.445 ;
        RECT 107.395 145.835 107.645 146.615 ;
        RECT 107.895 146.065 108.145 146.445 ;
        RECT 108.315 146.235 108.670 146.615 ;
        RECT 109.675 146.225 110.010 146.445 ;
        RECT 109.275 146.065 109.505 146.105 ;
        RECT 107.895 145.865 109.505 146.065 ;
        RECT 107.895 145.855 108.730 145.865 ;
        RECT 109.320 145.775 109.505 145.865 ;
        RECT 106.965 144.565 107.135 145.765 ;
        RECT 108.835 145.665 109.165 145.695 ;
        RECT 107.365 145.605 109.165 145.665 ;
        RECT 109.755 145.605 110.010 146.225 ;
        RECT 107.305 145.495 110.010 145.605 ;
        RECT 107.305 145.460 107.505 145.495 ;
        RECT 107.305 144.885 107.475 145.460 ;
        RECT 108.835 145.435 110.010 145.495 ;
        RECT 110.185 145.645 110.495 146.445 ;
        RECT 110.665 145.815 110.975 146.615 ;
        RECT 111.145 145.985 111.405 146.445 ;
        RECT 111.575 146.155 111.830 146.615 ;
        RECT 112.005 145.985 112.265 146.445 ;
        RECT 111.145 145.815 112.265 145.985 ;
        RECT 110.185 145.475 111.215 145.645 ;
        RECT 107.705 145.020 108.115 145.325 ;
        RECT 108.285 145.055 108.615 145.265 ;
        RECT 107.305 144.765 107.575 144.885 ;
        RECT 107.305 144.720 108.150 144.765 ;
        RECT 107.395 144.595 108.150 144.720 ;
        RECT 108.405 144.655 108.615 145.055 ;
        RECT 108.860 145.055 109.335 145.265 ;
        RECT 109.525 145.055 110.015 145.255 ;
        RECT 108.860 144.655 109.080 145.055 ;
        RECT 106.965 144.235 107.225 144.565 ;
        RECT 107.980 144.445 108.150 144.595 ;
        RECT 107.395 144.065 107.725 144.425 ;
        RECT 107.980 144.235 109.280 144.445 ;
        RECT 109.555 144.065 110.010 144.830 ;
        RECT 110.185 144.565 110.355 145.475 ;
        RECT 110.525 144.735 110.875 145.305 ;
        RECT 111.045 145.225 111.215 145.475 ;
        RECT 112.005 145.565 112.265 145.815 ;
        RECT 112.435 145.745 112.720 146.615 ;
        RECT 112.005 145.395 112.760 145.565 ;
        RECT 112.945 145.450 113.235 146.615 ;
        RECT 113.405 145.525 114.615 146.615 ;
        RECT 114.875 145.945 115.045 146.445 ;
        RECT 115.215 146.115 115.545 146.615 ;
        RECT 114.875 145.775 115.540 145.945 ;
        RECT 111.045 145.055 112.185 145.225 ;
        RECT 112.355 144.885 112.760 145.395 ;
        RECT 111.110 144.715 112.760 144.885 ;
        RECT 113.405 144.815 113.925 145.355 ;
        RECT 114.095 144.985 114.615 145.525 ;
        RECT 114.790 144.955 115.140 145.605 ;
        RECT 110.185 144.235 110.485 144.565 ;
        RECT 110.655 144.065 110.930 144.545 ;
        RECT 111.110 144.325 111.405 144.715 ;
        RECT 111.575 144.065 111.830 144.545 ;
        RECT 112.005 144.325 112.265 144.715 ;
        RECT 112.435 144.065 112.715 144.545 ;
        RECT 112.945 144.065 113.235 144.790 ;
        RECT 113.405 144.065 114.615 144.815 ;
        RECT 115.310 144.785 115.540 145.775 ;
        RECT 114.875 144.615 115.540 144.785 ;
        RECT 114.875 144.325 115.045 144.615 ;
        RECT 115.215 144.065 115.545 144.445 ;
        RECT 115.715 144.325 115.900 146.445 ;
        RECT 116.140 146.155 116.405 146.615 ;
        RECT 116.575 146.020 116.825 146.445 ;
        RECT 117.035 146.170 118.140 146.340 ;
        RECT 116.520 145.890 116.825 146.020 ;
        RECT 116.070 144.695 116.350 145.645 ;
        RECT 116.520 144.785 116.690 145.890 ;
        RECT 116.860 145.105 117.100 145.700 ;
        RECT 117.270 145.635 117.800 146.000 ;
        RECT 117.270 144.935 117.440 145.635 ;
        RECT 117.970 145.555 118.140 146.170 ;
        RECT 118.310 145.815 118.480 146.615 ;
        RECT 118.650 146.115 118.900 146.445 ;
        RECT 119.125 146.145 120.010 146.315 ;
        RECT 117.970 145.465 118.480 145.555 ;
        RECT 116.520 144.655 116.745 144.785 ;
        RECT 116.915 144.715 117.440 144.935 ;
        RECT 117.610 145.295 118.480 145.465 ;
        RECT 116.155 144.065 116.405 144.525 ;
        RECT 116.575 144.515 116.745 144.655 ;
        RECT 117.610 144.515 117.780 145.295 ;
        RECT 118.310 145.225 118.480 145.295 ;
        RECT 117.990 145.045 118.190 145.075 ;
        RECT 118.650 145.045 118.820 146.115 ;
        RECT 118.990 145.225 119.180 145.945 ;
        RECT 117.990 144.745 118.820 145.045 ;
        RECT 119.350 145.015 119.670 145.975 ;
        RECT 116.575 144.345 116.910 144.515 ;
        RECT 117.105 144.345 117.780 144.515 ;
        RECT 118.100 144.065 118.470 144.565 ;
        RECT 118.650 144.515 118.820 144.745 ;
        RECT 119.205 144.685 119.670 145.015 ;
        RECT 119.840 145.305 120.010 146.145 ;
        RECT 120.190 146.115 120.505 146.615 ;
        RECT 120.735 145.885 121.075 146.445 ;
        RECT 120.180 145.510 121.075 145.885 ;
        RECT 121.245 145.605 121.415 146.615 ;
        RECT 120.885 145.305 121.075 145.510 ;
        RECT 121.585 145.555 121.915 146.400 ;
        RECT 121.585 145.475 121.975 145.555 ;
        RECT 122.145 145.525 123.355 146.615 ;
        RECT 121.760 145.425 121.975 145.475 ;
        RECT 119.840 144.975 120.715 145.305 ;
        RECT 120.885 144.975 121.635 145.305 ;
        RECT 119.840 144.515 120.010 144.975 ;
        RECT 120.885 144.805 121.085 144.975 ;
        RECT 121.805 144.845 121.975 145.425 ;
        RECT 121.750 144.805 121.975 144.845 ;
        RECT 118.650 144.345 119.055 144.515 ;
        RECT 119.225 144.345 120.010 144.515 ;
        RECT 120.285 144.065 120.495 144.595 ;
        RECT 120.755 144.280 121.085 144.805 ;
        RECT 121.595 144.720 121.975 144.805 ;
        RECT 122.145 144.815 122.665 145.355 ;
        RECT 122.835 144.985 123.355 145.525 ;
        RECT 121.255 144.065 121.425 144.675 ;
        RECT 121.595 144.285 121.925 144.720 ;
        RECT 122.145 144.065 123.355 144.815 ;
        RECT 123.525 144.345 123.805 146.445 ;
        RECT 123.995 145.855 124.780 146.615 ;
        RECT 125.175 145.785 125.560 146.445 ;
        RECT 125.175 145.685 125.585 145.785 ;
        RECT 123.975 145.475 125.585 145.685 ;
        RECT 125.885 145.595 126.085 146.385 ;
        RECT 123.975 144.875 124.250 145.475 ;
        RECT 125.755 145.425 126.085 145.595 ;
        RECT 126.255 145.435 126.575 146.615 ;
        RECT 126.755 145.665 127.030 146.435 ;
        RECT 127.200 146.005 127.530 146.435 ;
        RECT 127.700 146.175 127.895 146.615 ;
        RECT 128.075 146.005 128.405 146.435 ;
        RECT 127.200 145.835 128.405 146.005 ;
        RECT 126.755 145.475 127.340 145.665 ;
        RECT 127.510 145.505 128.405 145.835 ;
        RECT 128.585 145.525 129.795 146.615 ;
        RECT 125.755 145.305 125.935 145.425 ;
        RECT 124.420 145.055 124.775 145.305 ;
        RECT 124.970 145.255 125.435 145.305 ;
        RECT 124.965 145.085 125.435 145.255 ;
        RECT 124.970 145.055 125.435 145.085 ;
        RECT 125.605 145.055 125.935 145.305 ;
        RECT 126.110 145.055 126.575 145.255 ;
        RECT 123.975 144.695 125.225 144.875 ;
        RECT 124.860 144.625 125.225 144.695 ;
        RECT 125.395 144.675 126.575 144.845 ;
        RECT 124.035 144.065 124.205 144.525 ;
        RECT 125.395 144.455 125.725 144.675 ;
        RECT 124.475 144.275 125.725 144.455 ;
        RECT 125.895 144.065 126.065 144.505 ;
        RECT 126.235 144.260 126.575 144.675 ;
        RECT 126.755 144.655 126.995 145.305 ;
        RECT 127.165 144.805 127.340 145.475 ;
        RECT 127.510 144.975 127.925 145.305 ;
        RECT 128.105 144.975 128.400 145.305 ;
        RECT 127.165 144.625 127.495 144.805 ;
        RECT 126.770 144.065 127.100 144.455 ;
        RECT 127.270 144.245 127.495 144.625 ;
        RECT 127.695 144.355 127.925 144.975 ;
        RECT 128.585 144.815 129.105 145.355 ;
        RECT 129.275 144.985 129.795 145.525 ;
        RECT 129.985 145.725 130.245 146.435 ;
        RECT 130.415 145.905 130.745 146.615 ;
        RECT 130.915 145.725 131.145 146.435 ;
        RECT 129.985 145.485 131.145 145.725 ;
        RECT 131.325 145.705 131.595 146.435 ;
        RECT 131.775 145.885 132.115 146.615 ;
        RECT 131.325 145.485 132.095 145.705 ;
        RECT 129.975 144.975 130.275 145.305 ;
        RECT 130.455 144.995 130.980 145.305 ;
        RECT 131.160 144.995 131.625 145.305 ;
        RECT 128.105 144.065 128.405 144.795 ;
        RECT 128.585 144.065 129.795 144.815 ;
        RECT 129.985 144.065 130.275 144.795 ;
        RECT 130.455 144.355 130.685 144.995 ;
        RECT 131.805 144.815 132.095 145.485 ;
        RECT 130.865 144.615 132.095 144.815 ;
        RECT 130.865 144.245 131.175 144.615 ;
        RECT 131.355 144.065 132.025 144.435 ;
        RECT 132.285 144.245 132.545 146.435 ;
        RECT 132.725 145.745 133.000 146.445 ;
        RECT 133.210 146.070 133.425 146.615 ;
        RECT 133.595 146.105 134.070 146.445 ;
        RECT 134.240 146.110 134.855 146.615 ;
        RECT 134.240 145.935 134.435 146.110 ;
        RECT 132.725 144.715 132.895 145.745 ;
        RECT 133.170 145.575 133.885 145.870 ;
        RECT 134.105 145.745 134.435 145.935 ;
        RECT 134.605 145.575 134.855 145.940 ;
        RECT 133.065 145.405 134.855 145.575 ;
        RECT 133.065 144.975 133.295 145.405 ;
        RECT 132.725 144.235 132.985 144.715 ;
        RECT 133.465 144.705 133.875 145.225 ;
        RECT 133.155 144.065 133.485 144.525 ;
        RECT 133.675 144.285 133.875 144.705 ;
        RECT 134.045 144.550 134.300 145.405 ;
        RECT 135.095 145.225 135.265 146.445 ;
        RECT 135.515 146.105 135.775 146.615 ;
        RECT 136.145 145.945 136.425 146.615 ;
        RECT 134.470 144.975 135.265 145.225 ;
        RECT 135.435 145.055 135.775 145.935 ;
        RECT 136.595 145.725 136.895 146.275 ;
        RECT 137.095 145.895 137.425 146.615 ;
        RECT 137.615 145.895 138.075 146.445 ;
        RECT 135.960 145.305 136.225 145.665 ;
        RECT 136.595 145.555 137.535 145.725 ;
        RECT 137.365 145.305 137.535 145.555 ;
        RECT 135.960 145.055 136.635 145.305 ;
        RECT 136.855 145.055 137.195 145.305 ;
        RECT 135.015 144.885 135.265 144.975 ;
        RECT 137.365 144.975 137.655 145.305 ;
        RECT 137.365 144.885 137.535 144.975 ;
        RECT 134.045 144.285 134.835 144.550 ;
        RECT 135.015 144.465 135.345 144.885 ;
        RECT 135.515 144.065 135.775 144.885 ;
        RECT 136.145 144.695 137.535 144.885 ;
        RECT 136.145 144.335 136.475 144.695 ;
        RECT 137.825 144.525 138.075 145.895 ;
        RECT 138.705 145.450 138.995 146.615 ;
        RECT 139.255 145.685 139.425 146.445 ;
        RECT 139.605 145.855 139.935 146.615 ;
        RECT 139.255 145.515 139.920 145.685 ;
        RECT 140.105 145.540 140.375 146.445 ;
        RECT 139.750 145.370 139.920 145.515 ;
        RECT 139.185 144.965 139.515 145.335 ;
        RECT 139.750 145.040 140.035 145.370 ;
        RECT 137.095 144.065 137.345 144.525 ;
        RECT 137.515 144.235 138.075 144.525 ;
        RECT 138.705 144.065 138.995 144.790 ;
        RECT 139.750 144.785 139.920 145.040 ;
        RECT 139.255 144.615 139.920 144.785 ;
        RECT 140.205 144.740 140.375 145.540 ;
        RECT 140.605 145.475 140.815 146.615 ;
        RECT 140.985 145.465 141.315 146.445 ;
        RECT 141.485 145.475 141.715 146.615 ;
        RECT 141.925 145.475 142.205 146.615 ;
        RECT 142.375 145.465 142.705 146.445 ;
        RECT 142.875 145.475 143.135 146.615 ;
        RECT 143.490 145.645 143.880 145.820 ;
        RECT 144.365 145.815 144.695 146.615 ;
        RECT 144.865 145.825 145.400 146.445 ;
        RECT 145.605 146.060 146.210 146.615 ;
        RECT 146.385 146.105 146.865 146.445 ;
        RECT 147.035 146.070 147.290 146.615 ;
        RECT 145.605 145.960 146.220 146.060 ;
        RECT 143.490 145.475 144.915 145.645 ;
        RECT 139.255 144.235 139.425 144.615 ;
        RECT 139.605 144.065 139.935 144.445 ;
        RECT 140.115 144.235 140.375 144.740 ;
        RECT 140.605 144.065 140.815 144.885 ;
        RECT 140.985 144.865 141.235 145.465 ;
        RECT 141.405 145.055 141.735 145.305 ;
        RECT 141.935 145.035 142.270 145.305 ;
        RECT 140.985 144.235 141.315 144.865 ;
        RECT 141.485 144.065 141.715 144.885 ;
        RECT 142.440 144.865 142.610 145.465 ;
        RECT 142.780 145.055 143.115 145.305 ;
        RECT 141.925 144.065 142.235 144.865 ;
        RECT 142.440 144.235 143.135 144.865 ;
        RECT 143.365 144.745 143.720 145.305 ;
        RECT 143.890 144.575 144.060 145.475 ;
        RECT 144.230 144.745 144.495 145.305 ;
        RECT 144.745 144.975 144.915 145.475 ;
        RECT 145.085 144.805 145.400 145.825 ;
        RECT 146.035 145.935 146.220 145.960 ;
        RECT 145.605 145.340 145.865 145.790 ;
        RECT 146.035 145.690 146.365 145.935 ;
        RECT 146.535 145.615 147.290 145.865 ;
        RECT 147.460 145.745 147.735 146.445 ;
        RECT 146.520 145.580 147.290 145.615 ;
        RECT 146.505 145.570 147.290 145.580 ;
        RECT 146.500 145.555 147.395 145.570 ;
        RECT 146.480 145.540 147.395 145.555 ;
        RECT 146.460 145.530 147.395 145.540 ;
        RECT 146.435 145.520 147.395 145.530 ;
        RECT 146.365 145.490 147.395 145.520 ;
        RECT 146.345 145.460 147.395 145.490 ;
        RECT 146.325 145.430 147.395 145.460 ;
        RECT 146.295 145.405 147.395 145.430 ;
        RECT 146.260 145.370 147.395 145.405 ;
        RECT 146.230 145.365 147.395 145.370 ;
        RECT 146.230 145.360 146.620 145.365 ;
        RECT 146.230 145.350 146.595 145.360 ;
        RECT 146.230 145.345 146.580 145.350 ;
        RECT 146.230 145.340 146.565 145.345 ;
        RECT 145.605 145.335 146.565 145.340 ;
        RECT 145.605 145.325 146.555 145.335 ;
        RECT 145.605 145.320 146.545 145.325 ;
        RECT 145.605 145.310 146.535 145.320 ;
        RECT 145.605 145.300 146.530 145.310 ;
        RECT 145.605 145.295 146.525 145.300 ;
        RECT 145.605 145.280 146.515 145.295 ;
        RECT 145.605 145.265 146.510 145.280 ;
        RECT 145.605 145.240 146.500 145.265 ;
        RECT 145.605 145.170 146.495 145.240 ;
        RECT 143.470 144.065 143.710 144.575 ;
        RECT 143.890 144.245 144.170 144.575 ;
        RECT 144.400 144.065 144.615 144.575 ;
        RECT 144.785 144.235 145.400 144.805 ;
        RECT 145.605 144.615 146.155 145.000 ;
        RECT 146.325 144.445 146.495 145.170 ;
        RECT 145.605 144.275 146.495 144.445 ;
        RECT 146.665 144.770 146.995 145.195 ;
        RECT 147.165 144.970 147.395 145.365 ;
        RECT 146.665 144.285 146.885 144.770 ;
        RECT 147.565 144.715 147.735 145.745 ;
        RECT 148.425 145.555 148.755 146.400 ;
        RECT 148.925 145.605 149.095 146.615 ;
        RECT 149.265 145.885 149.605 146.445 ;
        RECT 149.835 146.115 150.150 146.615 ;
        RECT 150.330 146.145 151.215 146.315 ;
        RECT 148.365 145.475 148.755 145.555 ;
        RECT 149.265 145.510 150.160 145.885 ;
        RECT 148.365 145.425 148.580 145.475 ;
        RECT 148.365 144.845 148.535 145.425 ;
        RECT 149.265 145.305 149.455 145.510 ;
        RECT 150.330 145.305 150.500 146.145 ;
        RECT 151.440 146.115 151.690 146.445 ;
        RECT 148.705 144.975 149.455 145.305 ;
        RECT 149.625 144.975 150.500 145.305 ;
        RECT 148.365 144.805 148.590 144.845 ;
        RECT 149.255 144.805 149.455 144.975 ;
        RECT 148.365 144.720 148.745 144.805 ;
        RECT 147.055 144.065 147.305 144.605 ;
        RECT 147.475 144.235 147.735 144.715 ;
        RECT 148.415 144.285 148.745 144.720 ;
        RECT 148.915 144.065 149.085 144.675 ;
        RECT 149.255 144.280 149.585 144.805 ;
        RECT 149.845 144.065 150.055 144.595 ;
        RECT 150.330 144.515 150.500 144.975 ;
        RECT 150.670 145.015 150.990 145.975 ;
        RECT 151.160 145.225 151.350 145.945 ;
        RECT 151.520 145.045 151.690 146.115 ;
        RECT 151.860 145.815 152.030 146.615 ;
        RECT 152.200 146.170 153.305 146.340 ;
        RECT 152.200 145.555 152.370 146.170 ;
        RECT 153.515 146.020 153.765 146.445 ;
        RECT 153.935 146.155 154.200 146.615 ;
        RECT 152.540 145.635 153.070 146.000 ;
        RECT 153.515 145.890 153.820 146.020 ;
        RECT 151.860 145.465 152.370 145.555 ;
        RECT 151.860 145.295 152.730 145.465 ;
        RECT 151.860 145.225 152.030 145.295 ;
        RECT 152.150 145.045 152.350 145.075 ;
        RECT 150.670 144.685 151.135 145.015 ;
        RECT 151.520 144.745 152.350 145.045 ;
        RECT 151.520 144.515 151.690 144.745 ;
        RECT 150.330 144.345 151.115 144.515 ;
        RECT 151.285 144.345 151.690 144.515 ;
        RECT 151.870 144.065 152.240 144.565 ;
        RECT 152.560 144.515 152.730 145.295 ;
        RECT 152.900 144.935 153.070 145.635 ;
        RECT 153.240 145.105 153.480 145.700 ;
        RECT 152.900 144.715 153.425 144.935 ;
        RECT 153.650 144.785 153.820 145.890 ;
        RECT 153.595 144.655 153.820 144.785 ;
        RECT 153.990 144.695 154.270 145.645 ;
        RECT 153.595 144.515 153.765 144.655 ;
        RECT 152.560 144.345 153.235 144.515 ;
        RECT 153.430 144.345 153.765 144.515 ;
        RECT 153.935 144.065 154.185 144.525 ;
        RECT 154.440 144.325 154.625 146.445 ;
        RECT 154.795 146.115 155.125 146.615 ;
        RECT 155.295 145.945 155.465 146.445 ;
        RECT 154.800 145.775 155.465 145.945 ;
        RECT 154.800 144.785 155.030 145.775 ;
        RECT 155.200 144.955 155.550 145.605 ;
        RECT 155.725 145.525 156.935 146.615 ;
        RECT 155.725 144.985 156.245 145.525 ;
        RECT 156.415 144.815 156.935 145.355 ;
        RECT 154.800 144.615 155.465 144.785 ;
        RECT 154.795 144.065 155.125 144.445 ;
        RECT 155.295 144.325 155.465 144.615 ;
        RECT 155.725 144.065 156.935 144.815 ;
        RECT 22.700 143.895 157.020 144.065 ;
        RECT 22.785 143.145 23.995 143.895 ;
        RECT 24.255 143.345 24.425 143.635 ;
        RECT 24.595 143.515 24.925 143.895 ;
        RECT 24.255 143.175 24.920 143.345 ;
        RECT 22.785 142.605 23.305 143.145 ;
        RECT 23.475 142.435 23.995 142.975 ;
        RECT 22.785 141.345 23.995 142.435 ;
        RECT 24.170 142.355 24.520 143.005 ;
        RECT 24.690 142.185 24.920 143.175 ;
        RECT 24.255 142.015 24.920 142.185 ;
        RECT 24.255 141.515 24.425 142.015 ;
        RECT 24.595 141.345 24.925 141.845 ;
        RECT 25.095 141.515 25.280 143.635 ;
        RECT 25.535 143.435 25.785 143.895 ;
        RECT 25.955 143.445 26.290 143.615 ;
        RECT 26.485 143.445 27.160 143.615 ;
        RECT 25.955 143.305 26.125 143.445 ;
        RECT 25.450 142.315 25.730 143.265 ;
        RECT 25.900 143.175 26.125 143.305 ;
        RECT 25.900 142.070 26.070 143.175 ;
        RECT 26.295 143.025 26.820 143.245 ;
        RECT 26.240 142.260 26.480 142.855 ;
        RECT 26.650 142.325 26.820 143.025 ;
        RECT 26.990 142.665 27.160 143.445 ;
        RECT 27.480 143.395 27.850 143.895 ;
        RECT 28.030 143.445 28.435 143.615 ;
        RECT 28.605 143.445 29.390 143.615 ;
        RECT 28.030 143.215 28.200 143.445 ;
        RECT 27.370 142.915 28.200 143.215 ;
        RECT 28.585 142.945 29.050 143.275 ;
        RECT 27.370 142.885 27.570 142.915 ;
        RECT 27.690 142.665 27.860 142.735 ;
        RECT 26.990 142.495 27.860 142.665 ;
        RECT 27.350 142.405 27.860 142.495 ;
        RECT 25.900 141.940 26.205 142.070 ;
        RECT 26.650 141.960 27.180 142.325 ;
        RECT 25.520 141.345 25.785 141.805 ;
        RECT 25.955 141.515 26.205 141.940 ;
        RECT 27.350 141.790 27.520 142.405 ;
        RECT 26.415 141.620 27.520 141.790 ;
        RECT 27.690 141.345 27.860 142.145 ;
        RECT 28.030 141.845 28.200 142.915 ;
        RECT 28.370 142.015 28.560 142.735 ;
        RECT 28.730 141.985 29.050 142.945 ;
        RECT 29.220 142.985 29.390 143.445 ;
        RECT 29.665 143.365 29.875 143.895 ;
        RECT 30.135 143.155 30.465 143.680 ;
        RECT 30.635 143.285 30.805 143.895 ;
        RECT 30.975 143.240 31.305 143.675 ;
        RECT 31.855 143.495 32.185 143.895 ;
        RECT 32.355 143.325 32.685 143.665 ;
        RECT 33.735 143.495 34.065 143.895 ;
        RECT 30.975 143.155 31.355 143.240 ;
        RECT 30.265 142.985 30.465 143.155 ;
        RECT 31.130 143.115 31.355 143.155 ;
        RECT 29.220 142.655 30.095 142.985 ;
        RECT 30.265 142.655 31.015 142.985 ;
        RECT 28.030 141.515 28.280 141.845 ;
        RECT 29.220 141.815 29.390 142.655 ;
        RECT 30.265 142.450 30.455 142.655 ;
        RECT 31.185 142.535 31.355 143.115 ;
        RECT 31.140 142.485 31.355 142.535 ;
        RECT 29.560 142.075 30.455 142.450 ;
        RECT 30.965 142.405 31.355 142.485 ;
        RECT 31.700 143.155 34.065 143.325 ;
        RECT 34.235 143.170 34.565 143.680 ;
        RECT 28.505 141.645 29.390 141.815 ;
        RECT 29.570 141.345 29.885 141.845 ;
        RECT 30.115 141.515 30.455 142.075 ;
        RECT 30.625 141.345 30.795 142.355 ;
        RECT 30.965 141.560 31.295 142.405 ;
        RECT 31.700 142.155 31.870 143.155 ;
        RECT 33.895 142.985 34.065 143.155 ;
        RECT 32.040 142.325 32.285 142.985 ;
        RECT 32.500 142.325 32.765 142.985 ;
        RECT 32.960 142.325 33.245 142.985 ;
        RECT 33.420 142.655 33.725 142.985 ;
        RECT 33.895 142.655 34.205 142.985 ;
        RECT 33.420 142.325 33.635 142.655 ;
        RECT 31.700 141.985 32.155 142.155 ;
        RECT 31.825 141.555 32.155 141.985 ;
        RECT 32.335 141.985 33.625 142.155 ;
        RECT 32.335 141.565 32.585 141.985 ;
        RECT 32.815 141.345 33.145 141.815 ;
        RECT 33.375 141.565 33.625 141.985 ;
        RECT 33.815 141.345 34.065 142.485 ;
        RECT 34.375 142.405 34.565 143.170 ;
        RECT 34.745 143.125 36.415 143.895 ;
        RECT 36.585 143.155 36.970 143.725 ;
        RECT 37.140 143.435 37.465 143.895 ;
        RECT 37.985 143.265 38.265 143.725 ;
        RECT 34.745 142.605 35.495 143.125 ;
        RECT 35.665 142.435 36.415 142.955 ;
        RECT 34.235 141.555 34.565 142.405 ;
        RECT 34.745 141.345 36.415 142.435 ;
        RECT 36.585 142.485 36.865 143.155 ;
        RECT 37.140 143.095 38.265 143.265 ;
        RECT 37.140 142.985 37.590 143.095 ;
        RECT 37.035 142.655 37.590 142.985 ;
        RECT 38.455 142.925 38.855 143.725 ;
        RECT 39.255 143.435 39.525 143.895 ;
        RECT 39.695 143.265 39.980 143.725 ;
        RECT 36.585 141.515 36.970 142.485 ;
        RECT 37.140 142.195 37.590 142.655 ;
        RECT 37.760 142.365 38.855 142.925 ;
        RECT 37.140 141.975 38.265 142.195 ;
        RECT 37.140 141.345 37.465 141.805 ;
        RECT 37.985 141.515 38.265 141.975 ;
        RECT 38.455 141.515 38.855 142.365 ;
        RECT 39.025 143.095 39.980 143.265 ;
        RECT 40.355 143.345 40.525 143.725 ;
        RECT 40.705 143.515 41.035 143.895 ;
        RECT 40.355 143.175 41.020 143.345 ;
        RECT 41.215 143.220 41.475 143.725 ;
        RECT 39.025 142.195 39.235 143.095 ;
        RECT 39.405 142.365 40.095 142.925 ;
        RECT 40.285 142.625 40.615 142.995 ;
        RECT 40.850 142.920 41.020 143.175 ;
        RECT 40.850 142.590 41.135 142.920 ;
        RECT 40.850 142.445 41.020 142.590 ;
        RECT 40.355 142.275 41.020 142.445 ;
        RECT 41.305 142.420 41.475 143.220 ;
        RECT 41.685 143.075 41.915 143.895 ;
        RECT 42.085 143.095 42.415 143.725 ;
        RECT 41.665 142.655 41.995 142.905 ;
        RECT 42.165 142.495 42.415 143.095 ;
        RECT 42.585 143.075 42.795 143.895 ;
        RECT 43.065 143.075 43.295 143.895 ;
        RECT 43.465 143.095 43.795 143.725 ;
        RECT 43.045 142.655 43.375 142.905 ;
        RECT 43.545 142.495 43.795 143.095 ;
        RECT 43.965 143.075 44.175 143.895 ;
        RECT 39.025 141.975 39.980 142.195 ;
        RECT 39.255 141.345 39.525 141.805 ;
        RECT 39.695 141.515 39.980 141.975 ;
        RECT 40.355 141.515 40.525 142.275 ;
        RECT 40.705 141.345 41.035 142.105 ;
        RECT 41.205 141.515 41.475 142.420 ;
        RECT 41.685 141.345 41.915 142.485 ;
        RECT 42.085 141.515 42.415 142.495 ;
        RECT 42.585 141.345 42.795 142.485 ;
        RECT 43.065 141.345 43.295 142.485 ;
        RECT 43.465 141.515 43.795 142.495 ;
        RECT 43.965 141.345 44.175 142.485 ;
        RECT 44.405 141.515 44.685 143.615 ;
        RECT 44.915 143.435 45.085 143.895 ;
        RECT 45.355 143.505 46.605 143.685 ;
        RECT 45.740 143.265 46.105 143.335 ;
        RECT 44.855 143.085 46.105 143.265 ;
        RECT 46.275 143.285 46.605 143.505 ;
        RECT 46.775 143.455 46.945 143.895 ;
        RECT 47.115 143.285 47.455 143.700 ;
        RECT 46.275 143.115 47.455 143.285 ;
        RECT 48.545 143.170 48.835 143.895 ;
        RECT 49.005 143.220 49.275 143.565 ;
        RECT 49.465 143.495 49.845 143.895 ;
        RECT 50.015 143.325 50.185 143.675 ;
        RECT 50.355 143.415 51.090 143.895 ;
        RECT 44.855 142.485 45.130 143.085 ;
        RECT 45.300 142.655 45.655 142.905 ;
        RECT 45.850 142.875 46.315 142.905 ;
        RECT 45.845 142.705 46.315 142.875 ;
        RECT 45.850 142.655 46.315 142.705 ;
        RECT 46.485 142.655 46.815 142.905 ;
        RECT 46.990 142.705 47.455 142.905 ;
        RECT 46.635 142.535 46.815 142.655 ;
        RECT 44.855 142.275 46.465 142.485 ;
        RECT 46.635 142.365 46.965 142.535 ;
        RECT 46.055 142.175 46.465 142.275 ;
        RECT 44.875 141.345 45.660 142.105 ;
        RECT 46.055 141.515 46.440 142.175 ;
        RECT 46.765 141.575 46.965 142.365 ;
        RECT 47.135 141.345 47.455 142.525 ;
        RECT 48.545 141.345 48.835 142.510 ;
        RECT 49.005 142.485 49.175 143.220 ;
        RECT 49.445 143.155 50.185 143.325 ;
        RECT 51.260 143.245 51.570 143.715 ;
        RECT 49.445 142.985 49.615 143.155 ;
        RECT 50.835 143.075 51.570 143.245 ;
        RECT 52.225 143.245 52.485 143.725 ;
        RECT 52.655 143.355 52.905 143.895 ;
        RECT 50.835 142.985 51.085 143.075 ;
        RECT 49.385 142.655 49.615 142.985 ;
        RECT 50.345 142.655 51.085 142.985 ;
        RECT 51.255 142.655 51.590 142.905 ;
        RECT 49.445 142.485 49.615 142.655 ;
        RECT 49.005 141.515 49.275 142.485 ;
        RECT 49.445 142.315 50.690 142.485 ;
        RECT 49.485 141.345 49.765 142.145 ;
        RECT 50.270 142.065 50.690 142.315 ;
        RECT 50.915 142.095 51.085 142.655 ;
        RECT 49.945 141.565 51.140 141.895 ;
        RECT 51.335 141.345 51.590 142.485 ;
        RECT 52.225 142.215 52.395 143.245 ;
        RECT 53.075 143.190 53.295 143.675 ;
        RECT 52.565 142.595 52.795 142.990 ;
        RECT 52.965 142.765 53.295 143.190 ;
        RECT 53.465 143.515 54.355 143.685 ;
        RECT 54.525 143.515 55.415 143.685 ;
        RECT 53.465 142.790 53.635 143.515 ;
        RECT 53.805 142.960 54.355 143.345 ;
        RECT 54.525 142.960 55.075 143.345 ;
        RECT 55.245 142.790 55.415 143.515 ;
        RECT 53.465 142.720 54.355 142.790 ;
        RECT 53.460 142.695 54.355 142.720 ;
        RECT 53.450 142.680 54.355 142.695 ;
        RECT 53.445 142.665 54.355 142.680 ;
        RECT 53.435 142.660 54.355 142.665 ;
        RECT 53.430 142.650 54.355 142.660 ;
        RECT 53.425 142.640 54.355 142.650 ;
        RECT 53.415 142.635 54.355 142.640 ;
        RECT 53.405 142.625 54.355 142.635 ;
        RECT 53.395 142.620 54.355 142.625 ;
        RECT 53.395 142.615 53.730 142.620 ;
        RECT 53.380 142.610 53.730 142.615 ;
        RECT 53.365 142.600 53.730 142.610 ;
        RECT 53.340 142.595 53.730 142.600 ;
        RECT 52.565 142.590 53.730 142.595 ;
        RECT 52.565 142.555 53.700 142.590 ;
        RECT 52.565 142.530 53.665 142.555 ;
        RECT 52.565 142.500 53.635 142.530 ;
        RECT 52.565 142.470 53.615 142.500 ;
        RECT 52.565 142.440 53.595 142.470 ;
        RECT 52.565 142.430 53.525 142.440 ;
        RECT 52.565 142.420 53.500 142.430 ;
        RECT 52.565 142.405 53.480 142.420 ;
        RECT 52.565 142.390 53.460 142.405 ;
        RECT 52.670 142.380 53.455 142.390 ;
        RECT 52.670 142.345 53.440 142.380 ;
        RECT 52.225 141.515 52.500 142.215 ;
        RECT 52.670 142.095 53.425 142.345 ;
        RECT 53.595 142.025 53.925 142.270 ;
        RECT 54.095 142.170 54.355 142.620 ;
        RECT 54.525 142.720 55.415 142.790 ;
        RECT 55.585 143.190 55.805 143.675 ;
        RECT 55.975 143.355 56.225 143.895 ;
        RECT 56.395 143.245 56.655 143.725 ;
        RECT 55.585 142.765 55.915 143.190 ;
        RECT 54.525 142.695 55.420 142.720 ;
        RECT 54.525 142.680 55.430 142.695 ;
        RECT 54.525 142.665 55.435 142.680 ;
        RECT 54.525 142.660 55.445 142.665 ;
        RECT 54.525 142.650 55.450 142.660 ;
        RECT 54.525 142.640 55.455 142.650 ;
        RECT 54.525 142.635 55.465 142.640 ;
        RECT 54.525 142.625 55.475 142.635 ;
        RECT 54.525 142.620 55.485 142.625 ;
        RECT 54.525 142.170 54.785 142.620 ;
        RECT 55.150 142.615 55.485 142.620 ;
        RECT 55.150 142.610 55.500 142.615 ;
        RECT 55.150 142.600 55.515 142.610 ;
        RECT 55.150 142.595 55.540 142.600 ;
        RECT 56.085 142.595 56.315 142.990 ;
        RECT 55.150 142.590 56.315 142.595 ;
        RECT 55.180 142.555 56.315 142.590 ;
        RECT 55.215 142.530 56.315 142.555 ;
        RECT 55.245 142.500 56.315 142.530 ;
        RECT 55.265 142.470 56.315 142.500 ;
        RECT 55.285 142.440 56.315 142.470 ;
        RECT 55.355 142.430 56.315 142.440 ;
        RECT 55.380 142.420 56.315 142.430 ;
        RECT 55.400 142.405 56.315 142.420 ;
        RECT 55.420 142.390 56.315 142.405 ;
        RECT 55.425 142.380 56.210 142.390 ;
        RECT 55.440 142.345 56.210 142.380 ;
        RECT 53.740 142.000 53.925 142.025 ;
        RECT 54.955 142.025 55.285 142.270 ;
        RECT 55.455 142.095 56.210 142.345 ;
        RECT 56.485 142.215 56.655 143.245 ;
        RECT 54.955 142.000 55.140 142.025 ;
        RECT 53.740 141.900 54.355 142.000 ;
        RECT 52.670 141.345 52.925 141.890 ;
        RECT 53.095 141.515 53.575 141.855 ;
        RECT 53.750 141.345 54.355 141.900 ;
        RECT 54.525 141.900 55.140 142.000 ;
        RECT 54.525 141.345 55.130 141.900 ;
        RECT 55.305 141.515 55.785 141.855 ;
        RECT 55.955 141.345 56.210 141.890 ;
        RECT 56.380 141.515 56.655 142.215 ;
        RECT 56.825 143.155 57.210 143.725 ;
        RECT 57.380 143.435 57.705 143.895 ;
        RECT 58.225 143.265 58.505 143.725 ;
        RECT 56.825 142.485 57.105 143.155 ;
        RECT 57.380 143.095 58.505 143.265 ;
        RECT 57.380 142.985 57.830 143.095 ;
        RECT 57.275 142.655 57.830 142.985 ;
        RECT 58.695 142.925 59.095 143.725 ;
        RECT 59.495 143.435 59.765 143.895 ;
        RECT 59.935 143.265 60.220 143.725 ;
        RECT 56.825 141.515 57.210 142.485 ;
        RECT 57.380 142.195 57.830 142.655 ;
        RECT 58.000 142.365 59.095 142.925 ;
        RECT 57.380 141.975 58.505 142.195 ;
        RECT 57.380 141.345 57.705 141.805 ;
        RECT 58.225 141.515 58.505 141.975 ;
        RECT 58.695 141.515 59.095 142.365 ;
        RECT 59.265 143.095 60.220 143.265 ;
        RECT 60.505 143.155 60.890 143.725 ;
        RECT 61.060 143.435 61.385 143.895 ;
        RECT 61.905 143.265 62.185 143.725 ;
        RECT 59.265 142.195 59.475 143.095 ;
        RECT 59.645 142.365 60.335 142.925 ;
        RECT 60.505 142.485 60.785 143.155 ;
        RECT 61.060 143.095 62.185 143.265 ;
        RECT 61.060 142.985 61.510 143.095 ;
        RECT 60.955 142.655 61.510 142.985 ;
        RECT 62.375 142.925 62.775 143.725 ;
        RECT 63.175 143.435 63.445 143.895 ;
        RECT 63.615 143.265 63.900 143.725 ;
        RECT 59.265 141.975 60.220 142.195 ;
        RECT 59.495 141.345 59.765 141.805 ;
        RECT 59.935 141.515 60.220 141.975 ;
        RECT 60.505 141.515 60.890 142.485 ;
        RECT 61.060 142.195 61.510 142.655 ;
        RECT 61.680 142.365 62.775 142.925 ;
        RECT 61.060 141.975 62.185 142.195 ;
        RECT 61.060 141.345 61.385 141.805 ;
        RECT 61.905 141.515 62.185 141.975 ;
        RECT 62.375 141.515 62.775 142.365 ;
        RECT 62.945 143.095 63.900 143.265 ;
        RECT 64.185 143.125 65.855 143.895 ;
        RECT 66.025 143.220 66.285 143.725 ;
        RECT 66.465 143.515 66.795 143.895 ;
        RECT 66.975 143.345 67.145 143.725 ;
        RECT 62.945 142.195 63.155 143.095 ;
        RECT 63.325 142.365 64.015 142.925 ;
        RECT 64.185 142.605 64.935 143.125 ;
        RECT 65.105 142.435 65.855 142.955 ;
        RECT 62.945 141.975 63.900 142.195 ;
        RECT 63.175 141.345 63.445 141.805 ;
        RECT 63.615 141.515 63.900 141.975 ;
        RECT 64.185 141.345 65.855 142.435 ;
        RECT 66.025 142.420 66.195 143.220 ;
        RECT 66.480 143.175 67.145 143.345 ;
        RECT 66.480 142.920 66.650 143.175 ;
        RECT 67.870 143.155 68.125 143.725 ;
        RECT 68.295 143.495 68.625 143.895 ;
        RECT 69.050 143.360 69.580 143.725 ;
        RECT 69.050 143.325 69.225 143.360 ;
        RECT 68.295 143.155 69.225 143.325 ;
        RECT 66.365 142.590 66.650 142.920 ;
        RECT 66.885 142.625 67.215 142.995 ;
        RECT 66.480 142.445 66.650 142.590 ;
        RECT 67.870 142.485 68.040 143.155 ;
        RECT 68.295 142.985 68.465 143.155 ;
        RECT 68.210 142.655 68.465 142.985 ;
        RECT 68.690 142.655 68.885 142.985 ;
        RECT 66.025 141.515 66.295 142.420 ;
        RECT 66.480 142.275 67.145 142.445 ;
        RECT 66.465 141.345 66.795 142.105 ;
        RECT 66.975 141.515 67.145 142.275 ;
        RECT 67.870 141.515 68.205 142.485 ;
        RECT 68.375 141.345 68.545 142.485 ;
        RECT 68.715 141.685 68.885 142.655 ;
        RECT 69.055 142.025 69.225 143.155 ;
        RECT 69.395 142.365 69.565 143.165 ;
        RECT 69.770 142.875 70.045 143.725 ;
        RECT 69.765 142.705 70.045 142.875 ;
        RECT 69.770 142.565 70.045 142.705 ;
        RECT 70.215 142.365 70.405 143.725 ;
        RECT 70.585 143.360 71.095 143.895 ;
        RECT 71.315 143.085 71.560 143.690 ;
        RECT 72.005 143.125 73.675 143.895 ;
        RECT 74.305 143.170 74.595 143.895 ;
        RECT 74.765 143.220 75.025 143.725 ;
        RECT 75.205 143.515 75.535 143.895 ;
        RECT 75.715 143.345 75.885 143.725 ;
        RECT 70.605 142.915 71.835 143.085 ;
        RECT 69.395 142.195 70.405 142.365 ;
        RECT 70.575 142.350 71.325 142.540 ;
        RECT 69.055 141.855 70.180 142.025 ;
        RECT 70.575 141.685 70.745 142.350 ;
        RECT 71.495 142.105 71.835 142.915 ;
        RECT 72.005 142.605 72.755 143.125 ;
        RECT 72.925 142.435 73.675 142.955 ;
        RECT 68.715 141.515 70.745 141.685 ;
        RECT 70.915 141.345 71.085 142.105 ;
        RECT 71.320 141.695 71.835 142.105 ;
        RECT 72.005 141.345 73.675 142.435 ;
        RECT 74.305 141.345 74.595 142.510 ;
        RECT 74.765 142.420 74.935 143.220 ;
        RECT 75.220 143.175 75.885 143.345 ;
        RECT 76.805 143.265 77.135 143.625 ;
        RECT 77.755 143.435 78.005 143.895 ;
        RECT 78.175 143.435 78.735 143.725 ;
        RECT 75.220 142.920 75.390 143.175 ;
        RECT 76.805 143.075 78.195 143.265 ;
        RECT 75.105 142.590 75.390 142.920 ;
        RECT 75.625 142.625 75.955 142.995 ;
        RECT 78.025 142.985 78.195 143.075 ;
        RECT 76.620 142.655 77.295 142.905 ;
        RECT 77.515 142.655 77.855 142.905 ;
        RECT 78.025 142.655 78.315 142.985 ;
        RECT 75.220 142.445 75.390 142.590 ;
        RECT 74.765 141.515 75.035 142.420 ;
        RECT 75.220 142.275 75.885 142.445 ;
        RECT 76.620 142.295 76.885 142.655 ;
        RECT 78.025 142.405 78.195 142.655 ;
        RECT 75.205 141.345 75.535 142.105 ;
        RECT 75.715 141.515 75.885 142.275 ;
        RECT 77.255 142.235 78.195 142.405 ;
        RECT 76.805 141.345 77.085 142.015 ;
        RECT 77.255 141.685 77.555 142.235 ;
        RECT 78.485 142.065 78.735 143.435 ;
        RECT 78.905 143.125 80.575 143.895 ;
        RECT 80.835 143.345 81.005 143.635 ;
        RECT 81.175 143.515 81.505 143.895 ;
        RECT 80.835 143.175 81.500 143.345 ;
        RECT 78.905 142.605 79.655 143.125 ;
        RECT 79.825 142.435 80.575 142.955 ;
        RECT 77.755 141.345 78.085 142.065 ;
        RECT 78.275 141.515 78.735 142.065 ;
        RECT 78.905 141.345 80.575 142.435 ;
        RECT 80.750 142.355 81.100 143.005 ;
        RECT 81.270 142.185 81.500 143.175 ;
        RECT 80.835 142.015 81.500 142.185 ;
        RECT 80.835 141.515 81.005 142.015 ;
        RECT 81.175 141.345 81.505 141.845 ;
        RECT 81.675 141.515 81.860 143.635 ;
        RECT 82.115 143.435 82.365 143.895 ;
        RECT 82.535 143.445 82.870 143.615 ;
        RECT 83.065 143.445 83.740 143.615 ;
        RECT 82.535 143.305 82.705 143.445 ;
        RECT 82.030 142.315 82.310 143.265 ;
        RECT 82.480 143.175 82.705 143.305 ;
        RECT 82.480 142.070 82.650 143.175 ;
        RECT 82.875 143.025 83.400 143.245 ;
        RECT 82.820 142.260 83.060 142.855 ;
        RECT 83.230 142.325 83.400 143.025 ;
        RECT 83.570 142.665 83.740 143.445 ;
        RECT 84.060 143.395 84.430 143.895 ;
        RECT 84.610 143.445 85.015 143.615 ;
        RECT 85.185 143.445 85.970 143.615 ;
        RECT 84.610 143.215 84.780 143.445 ;
        RECT 83.950 142.915 84.780 143.215 ;
        RECT 85.165 142.945 85.630 143.275 ;
        RECT 83.950 142.885 84.150 142.915 ;
        RECT 84.270 142.665 84.440 142.735 ;
        RECT 83.570 142.495 84.440 142.665 ;
        RECT 83.930 142.405 84.440 142.495 ;
        RECT 82.480 141.940 82.785 142.070 ;
        RECT 83.230 141.960 83.760 142.325 ;
        RECT 82.100 141.345 82.365 141.805 ;
        RECT 82.535 141.515 82.785 141.940 ;
        RECT 83.930 141.790 84.100 142.405 ;
        RECT 82.995 141.620 84.100 141.790 ;
        RECT 84.270 141.345 84.440 142.145 ;
        RECT 84.610 141.845 84.780 142.915 ;
        RECT 84.950 142.015 85.140 142.735 ;
        RECT 85.310 141.985 85.630 142.945 ;
        RECT 85.800 142.985 85.970 143.445 ;
        RECT 86.245 143.365 86.455 143.895 ;
        RECT 86.715 143.155 87.045 143.680 ;
        RECT 87.215 143.285 87.385 143.895 ;
        RECT 87.555 143.240 87.885 143.675 ;
        RECT 89.140 143.265 89.425 143.725 ;
        RECT 89.595 143.435 89.865 143.895 ;
        RECT 87.555 143.155 87.935 143.240 ;
        RECT 86.845 142.985 87.045 143.155 ;
        RECT 87.710 143.115 87.935 143.155 ;
        RECT 85.800 142.655 86.675 142.985 ;
        RECT 86.845 142.655 87.595 142.985 ;
        RECT 84.610 141.515 84.860 141.845 ;
        RECT 85.800 141.815 85.970 142.655 ;
        RECT 86.845 142.450 87.035 142.655 ;
        RECT 87.765 142.535 87.935 143.115 ;
        RECT 89.140 143.095 90.095 143.265 ;
        RECT 87.720 142.485 87.935 142.535 ;
        RECT 86.140 142.075 87.035 142.450 ;
        RECT 87.545 142.405 87.935 142.485 ;
        RECT 85.085 141.645 85.970 141.815 ;
        RECT 86.150 141.345 86.465 141.845 ;
        RECT 86.695 141.515 87.035 142.075 ;
        RECT 87.205 141.345 87.375 142.355 ;
        RECT 87.545 141.560 87.875 142.405 ;
        RECT 89.025 142.365 89.715 142.925 ;
        RECT 89.885 142.195 90.095 143.095 ;
        RECT 89.140 141.975 90.095 142.195 ;
        RECT 90.265 142.925 90.665 143.725 ;
        RECT 90.855 143.265 91.135 143.725 ;
        RECT 91.655 143.435 91.980 143.895 ;
        RECT 90.855 143.095 91.980 143.265 ;
        RECT 92.150 143.155 92.535 143.725 ;
        RECT 91.530 142.985 91.980 143.095 ;
        RECT 90.265 142.365 91.360 142.925 ;
        RECT 91.530 142.655 92.085 142.985 ;
        RECT 89.140 141.515 89.425 141.975 ;
        RECT 89.595 141.345 89.865 141.805 ;
        RECT 90.265 141.515 90.665 142.365 ;
        RECT 91.530 142.195 91.980 142.655 ;
        RECT 92.255 142.485 92.535 143.155 ;
        RECT 92.710 143.130 93.165 143.895 ;
        RECT 93.440 143.515 94.740 143.725 ;
        RECT 94.995 143.535 95.325 143.895 ;
        RECT 94.570 143.365 94.740 143.515 ;
        RECT 95.495 143.395 95.755 143.725 ;
        RECT 93.640 142.905 93.860 143.305 ;
        RECT 92.705 142.705 93.195 142.905 ;
        RECT 93.385 142.695 93.860 142.905 ;
        RECT 94.105 142.905 94.315 143.305 ;
        RECT 94.570 143.240 95.325 143.365 ;
        RECT 94.570 143.195 95.415 143.240 ;
        RECT 95.145 143.075 95.415 143.195 ;
        RECT 94.105 142.695 94.435 142.905 ;
        RECT 94.605 142.635 95.015 142.940 ;
        RECT 90.855 141.975 91.980 142.195 ;
        RECT 90.855 141.515 91.135 141.975 ;
        RECT 91.655 141.345 91.980 141.805 ;
        RECT 92.150 141.515 92.535 142.485 ;
        RECT 92.710 142.465 93.885 142.525 ;
        RECT 95.245 142.500 95.415 143.075 ;
        RECT 95.215 142.465 95.415 142.500 ;
        RECT 92.710 142.355 95.415 142.465 ;
        RECT 92.710 141.735 92.965 142.355 ;
        RECT 93.555 142.295 95.355 142.355 ;
        RECT 93.555 142.265 93.885 142.295 ;
        RECT 95.585 142.195 95.755 143.395 ;
        RECT 96.205 143.265 96.585 143.715 ;
        RECT 95.945 142.315 96.175 143.005 ;
        RECT 96.355 142.815 96.585 143.265 ;
        RECT 96.765 143.115 96.995 143.895 ;
        RECT 97.175 143.185 97.605 143.715 ;
        RECT 97.175 142.935 97.420 143.185 ;
        RECT 97.785 142.985 97.995 143.605 ;
        RECT 98.165 143.165 98.495 143.895 ;
        RECT 98.685 143.095 98.995 143.895 ;
        RECT 99.200 143.095 99.895 143.725 ;
        RECT 100.065 143.170 100.355 143.895 ;
        RECT 101.445 143.155 101.830 143.725 ;
        RECT 102.000 143.435 102.325 143.895 ;
        RECT 102.845 143.265 103.125 143.725 ;
        RECT 93.215 142.095 93.400 142.185 ;
        RECT 93.990 142.095 94.825 142.105 ;
        RECT 93.215 141.895 94.825 142.095 ;
        RECT 93.215 141.855 93.445 141.895 ;
        RECT 92.710 141.515 93.045 141.735 ;
        RECT 94.050 141.345 94.405 141.725 ;
        RECT 94.575 141.515 94.825 141.895 ;
        RECT 95.075 141.345 95.325 142.125 ;
        RECT 95.495 141.515 95.755 142.195 ;
        RECT 96.355 142.135 96.695 142.815 ;
        RECT 95.935 141.935 96.695 142.135 ;
        RECT 96.885 142.635 97.420 142.935 ;
        RECT 97.600 142.635 97.995 142.985 ;
        RECT 98.190 142.635 98.480 142.985 ;
        RECT 98.695 142.655 99.030 142.925 ;
        RECT 95.935 141.545 96.195 141.935 ;
        RECT 96.365 141.345 96.695 141.755 ;
        RECT 96.885 141.525 97.215 142.635 ;
        RECT 99.200 142.495 99.370 143.095 ;
        RECT 99.540 142.655 99.875 142.905 ;
        RECT 97.385 142.255 98.425 142.455 ;
        RECT 97.385 141.525 97.575 142.255 ;
        RECT 97.745 141.345 98.075 142.075 ;
        RECT 98.255 141.525 98.425 142.255 ;
        RECT 98.685 141.345 98.965 142.485 ;
        RECT 99.135 141.515 99.465 142.495 ;
        RECT 99.635 141.345 99.895 142.485 ;
        RECT 100.065 141.345 100.355 142.510 ;
        RECT 101.445 142.485 101.725 143.155 ;
        RECT 102.000 143.095 103.125 143.265 ;
        RECT 102.000 142.985 102.450 143.095 ;
        RECT 101.895 142.655 102.450 142.985 ;
        RECT 103.315 142.925 103.715 143.725 ;
        RECT 104.115 143.435 104.385 143.895 ;
        RECT 104.555 143.265 104.840 143.725 ;
        RECT 101.445 141.515 101.830 142.485 ;
        RECT 102.000 142.195 102.450 142.655 ;
        RECT 102.620 142.365 103.715 142.925 ;
        RECT 102.000 141.975 103.125 142.195 ;
        RECT 102.000 141.345 102.325 141.805 ;
        RECT 102.845 141.515 103.125 141.975 ;
        RECT 103.315 141.515 103.715 142.365 ;
        RECT 103.885 143.095 104.840 143.265 ;
        RECT 105.215 143.345 105.385 143.725 ;
        RECT 105.565 143.515 105.895 143.895 ;
        RECT 105.215 143.175 105.880 143.345 ;
        RECT 106.075 143.220 106.335 143.725 ;
        RECT 103.885 142.195 104.095 143.095 ;
        RECT 104.265 142.365 104.955 142.925 ;
        RECT 105.145 142.625 105.475 142.995 ;
        RECT 105.710 142.920 105.880 143.175 ;
        RECT 105.710 142.590 105.995 142.920 ;
        RECT 105.710 142.445 105.880 142.590 ;
        RECT 105.215 142.275 105.880 142.445 ;
        RECT 106.165 142.420 106.335 143.220 ;
        RECT 106.505 143.125 108.175 143.895 ;
        RECT 106.505 142.605 107.255 143.125 ;
        RECT 108.825 143.085 109.065 143.895 ;
        RECT 109.235 143.085 109.565 143.725 ;
        RECT 109.735 143.085 110.005 143.895 ;
        RECT 110.185 143.125 111.855 143.895 ;
        RECT 112.485 143.155 112.870 143.725 ;
        RECT 113.040 143.435 113.365 143.895 ;
        RECT 113.885 143.265 114.165 143.725 ;
        RECT 107.425 142.435 108.175 142.955 ;
        RECT 108.805 142.655 109.155 142.905 ;
        RECT 109.325 142.485 109.495 143.085 ;
        RECT 109.665 142.655 110.015 142.905 ;
        RECT 110.185 142.605 110.935 143.125 ;
        RECT 103.885 141.975 104.840 142.195 ;
        RECT 104.115 141.345 104.385 141.805 ;
        RECT 104.555 141.515 104.840 141.975 ;
        RECT 105.215 141.515 105.385 142.275 ;
        RECT 105.565 141.345 105.895 142.105 ;
        RECT 106.065 141.515 106.335 142.420 ;
        RECT 106.505 141.345 108.175 142.435 ;
        RECT 108.815 142.315 109.495 142.485 ;
        RECT 108.815 141.530 109.145 142.315 ;
        RECT 109.675 141.345 110.005 142.485 ;
        RECT 111.105 142.435 111.855 142.955 ;
        RECT 110.185 141.345 111.855 142.435 ;
        RECT 112.485 142.485 112.765 143.155 ;
        RECT 113.040 143.095 114.165 143.265 ;
        RECT 113.040 142.985 113.490 143.095 ;
        RECT 112.935 142.655 113.490 142.985 ;
        RECT 114.355 142.925 114.755 143.725 ;
        RECT 115.155 143.435 115.425 143.895 ;
        RECT 115.595 143.265 115.880 143.725 ;
        RECT 112.485 141.515 112.870 142.485 ;
        RECT 113.040 142.195 113.490 142.655 ;
        RECT 113.660 142.365 114.755 142.925 ;
        RECT 113.040 141.975 114.165 142.195 ;
        RECT 113.040 141.345 113.365 141.805 ;
        RECT 113.885 141.515 114.165 141.975 ;
        RECT 114.355 141.515 114.755 142.365 ;
        RECT 114.925 143.095 115.880 143.265 ;
        RECT 117.085 143.395 117.345 143.725 ;
        RECT 117.515 143.535 117.845 143.895 ;
        RECT 118.100 143.515 119.400 143.725 ;
        RECT 114.925 142.195 115.135 143.095 ;
        RECT 115.305 142.365 115.995 142.925 ;
        RECT 117.085 142.195 117.255 143.395 ;
        RECT 118.100 143.365 118.270 143.515 ;
        RECT 117.515 143.240 118.270 143.365 ;
        RECT 117.425 143.195 118.270 143.240 ;
        RECT 117.425 143.075 117.695 143.195 ;
        RECT 117.425 142.500 117.595 143.075 ;
        RECT 117.825 142.635 118.235 142.940 ;
        RECT 118.525 142.905 118.735 143.305 ;
        RECT 118.405 142.695 118.735 142.905 ;
        RECT 118.980 142.905 119.200 143.305 ;
        RECT 119.675 143.130 120.130 143.895 ;
        RECT 120.305 143.350 125.650 143.895 ;
        RECT 118.980 142.695 119.455 142.905 ;
        RECT 119.645 142.705 120.135 142.905 ;
        RECT 117.425 142.465 117.625 142.500 ;
        RECT 118.955 142.465 120.130 142.525 ;
        RECT 121.890 142.520 122.230 143.350 ;
        RECT 125.825 143.170 126.115 143.895 ;
        RECT 126.305 143.395 126.560 143.725 ;
        RECT 126.775 143.415 127.105 143.895 ;
        RECT 127.275 143.475 128.810 143.725 ;
        RECT 126.305 143.385 126.515 143.395 ;
        RECT 126.305 143.315 126.490 143.385 ;
        RECT 117.425 142.355 120.130 142.465 ;
        RECT 117.485 142.295 119.285 142.355 ;
        RECT 118.955 142.265 119.285 142.295 ;
        RECT 114.925 141.975 115.880 142.195 ;
        RECT 115.155 141.345 115.425 141.805 ;
        RECT 115.595 141.515 115.880 141.975 ;
        RECT 117.085 141.515 117.345 142.195 ;
        RECT 117.515 141.345 117.765 142.125 ;
        RECT 118.015 142.095 118.850 142.105 ;
        RECT 119.440 142.095 119.625 142.185 ;
        RECT 118.015 141.895 119.625 142.095 ;
        RECT 118.015 141.515 118.265 141.895 ;
        RECT 119.395 141.855 119.625 141.895 ;
        RECT 119.875 141.735 120.130 142.355 ;
        RECT 123.710 141.780 124.060 143.030 ;
        RECT 118.435 141.345 118.790 141.725 ;
        RECT 119.795 141.515 120.130 141.735 ;
        RECT 120.305 141.345 125.650 141.780 ;
        RECT 125.825 141.345 126.115 142.510 ;
        RECT 126.305 142.185 126.475 143.315 ;
        RECT 127.275 143.245 127.445 143.475 ;
        RECT 126.645 143.075 127.445 143.245 ;
        RECT 126.645 142.525 126.815 143.075 ;
        RECT 127.625 142.905 127.910 143.305 ;
        RECT 127.045 142.875 127.410 142.905 ;
        RECT 127.035 142.705 127.410 142.875 ;
        RECT 127.580 142.705 127.910 142.905 ;
        RECT 128.180 142.905 128.460 143.305 ;
        RECT 128.640 143.245 128.810 143.475 ;
        RECT 129.035 143.415 129.365 143.895 ;
        RECT 129.535 143.245 129.705 143.725 ;
        RECT 128.640 143.075 129.705 143.245 ;
        RECT 129.970 143.245 130.240 143.455 ;
        RECT 130.460 143.435 130.790 143.895 ;
        RECT 131.300 143.435 132.050 143.725 ;
        RECT 129.970 143.075 131.305 143.245 ;
        RECT 131.135 142.905 131.305 143.075 ;
        RECT 128.180 142.705 128.655 142.905 ;
        RECT 128.825 142.705 129.270 142.905 ;
        RECT 129.440 142.695 129.790 142.905 ;
        RECT 129.970 142.665 130.320 142.905 ;
        RECT 130.490 142.665 130.965 142.905 ;
        RECT 131.135 142.655 131.510 142.905 ;
        RECT 126.645 142.355 129.705 142.525 ;
        RECT 131.135 142.485 131.305 142.655 ;
        RECT 126.305 141.515 126.560 142.185 ;
        RECT 126.730 141.345 127.060 142.105 ;
        RECT 127.230 141.945 128.865 142.185 ;
        RECT 127.230 141.515 127.480 141.945 ;
        RECT 128.635 141.855 128.865 141.945 ;
        RECT 127.650 141.345 128.005 141.765 ;
        RECT 128.195 141.685 128.525 141.725 ;
        RECT 129.035 141.685 129.365 142.185 ;
        RECT 128.195 141.515 129.365 141.685 ;
        RECT 129.535 141.515 129.705 142.355 ;
        RECT 129.970 142.315 131.305 142.485 ;
        RECT 129.970 142.155 130.250 142.315 ;
        RECT 131.680 142.145 132.050 143.435 ;
        RECT 132.265 143.125 133.935 143.895 ;
        RECT 134.155 143.240 134.485 143.675 ;
        RECT 134.655 143.285 134.825 143.895 ;
        RECT 134.105 143.155 134.485 143.240 ;
        RECT 134.995 143.155 135.325 143.680 ;
        RECT 135.585 143.365 135.795 143.895 ;
        RECT 136.070 143.445 136.855 143.615 ;
        RECT 137.025 143.445 137.430 143.615 ;
        RECT 132.265 142.605 133.015 143.125 ;
        RECT 134.105 143.115 134.330 143.155 ;
        RECT 133.185 142.435 133.935 142.955 ;
        RECT 130.460 141.345 130.710 142.145 ;
        RECT 130.880 141.975 132.050 142.145 ;
        RECT 130.880 141.515 131.210 141.975 ;
        RECT 131.380 141.345 131.595 141.805 ;
        RECT 132.265 141.345 133.935 142.435 ;
        RECT 134.105 142.535 134.275 143.115 ;
        RECT 134.995 142.985 135.195 143.155 ;
        RECT 136.070 142.985 136.240 143.445 ;
        RECT 134.445 142.655 135.195 142.985 ;
        RECT 135.365 142.655 136.240 142.985 ;
        RECT 134.105 142.485 134.320 142.535 ;
        RECT 134.105 142.405 134.495 142.485 ;
        RECT 134.165 141.560 134.495 142.405 ;
        RECT 135.005 142.450 135.195 142.655 ;
        RECT 134.665 141.345 134.835 142.355 ;
        RECT 135.005 142.075 135.900 142.450 ;
        RECT 135.005 141.515 135.345 142.075 ;
        RECT 135.575 141.345 135.890 141.845 ;
        RECT 136.070 141.815 136.240 142.655 ;
        RECT 136.410 142.945 136.875 143.275 ;
        RECT 137.260 143.215 137.430 143.445 ;
        RECT 137.610 143.395 137.980 143.895 ;
        RECT 138.300 143.445 138.975 143.615 ;
        RECT 139.170 143.445 139.505 143.615 ;
        RECT 136.410 141.985 136.730 142.945 ;
        RECT 137.260 142.915 138.090 143.215 ;
        RECT 136.900 142.015 137.090 142.735 ;
        RECT 137.260 141.845 137.430 142.915 ;
        RECT 137.890 142.885 138.090 142.915 ;
        RECT 137.600 142.665 137.770 142.735 ;
        RECT 138.300 142.665 138.470 143.445 ;
        RECT 139.335 143.305 139.505 143.445 ;
        RECT 139.675 143.435 139.925 143.895 ;
        RECT 137.600 142.495 138.470 142.665 ;
        RECT 138.640 143.025 139.165 143.245 ;
        RECT 139.335 143.175 139.560 143.305 ;
        RECT 137.600 142.405 138.110 142.495 ;
        RECT 136.070 141.645 136.955 141.815 ;
        RECT 137.180 141.515 137.430 141.845 ;
        RECT 137.600 141.345 137.770 142.145 ;
        RECT 137.940 141.790 138.110 142.405 ;
        RECT 138.640 142.325 138.810 143.025 ;
        RECT 138.280 141.960 138.810 142.325 ;
        RECT 138.980 142.260 139.220 142.855 ;
        RECT 139.390 142.070 139.560 143.175 ;
        RECT 139.730 142.315 140.010 143.265 ;
        RECT 139.255 141.940 139.560 142.070 ;
        RECT 137.940 141.620 139.045 141.790 ;
        RECT 139.255 141.515 139.505 141.940 ;
        RECT 139.675 141.345 139.940 141.805 ;
        RECT 140.180 141.515 140.365 143.635 ;
        RECT 140.535 143.515 140.865 143.895 ;
        RECT 141.035 143.345 141.205 143.635 ;
        RECT 140.540 143.175 141.205 143.345 ;
        RECT 141.465 143.175 141.805 143.685 ;
        RECT 140.540 142.185 140.770 143.175 ;
        RECT 140.940 142.355 141.290 143.005 ;
        RECT 140.540 142.015 141.205 142.185 ;
        RECT 140.535 141.345 140.865 141.845 ;
        RECT 141.035 141.515 141.205 142.015 ;
        RECT 141.465 141.775 141.725 143.175 ;
        RECT 141.975 143.095 142.245 143.895 ;
        RECT 141.900 142.655 142.230 142.905 ;
        RECT 142.425 142.655 142.705 143.625 ;
        RECT 142.885 142.655 143.185 143.625 ;
        RECT 143.365 142.655 143.715 143.620 ;
        RECT 143.935 143.395 144.430 143.725 ;
        RECT 141.915 142.485 142.230 142.655 ;
        RECT 143.935 142.485 144.105 143.395 ;
        RECT 141.915 142.315 144.105 142.485 ;
        RECT 141.465 141.515 141.805 141.775 ;
        RECT 141.975 141.345 142.305 142.145 ;
        RECT 142.770 141.515 143.020 142.315 ;
        RECT 143.205 141.345 143.535 142.065 ;
        RECT 143.755 141.515 144.005 142.315 ;
        RECT 144.275 141.905 144.515 143.215 ;
        RECT 145.605 143.075 145.865 143.895 ;
        RECT 146.035 143.075 146.365 143.495 ;
        RECT 146.545 143.410 147.335 143.675 ;
        RECT 146.115 142.985 146.365 143.075 ;
        RECT 145.605 142.025 145.945 142.905 ;
        RECT 146.115 142.735 146.910 142.985 ;
        RECT 144.175 141.345 144.510 141.725 ;
        RECT 145.605 141.345 145.865 141.855 ;
        RECT 146.115 141.515 146.285 142.735 ;
        RECT 147.080 142.555 147.335 143.410 ;
        RECT 147.505 143.255 147.705 143.675 ;
        RECT 147.895 143.435 148.225 143.895 ;
        RECT 147.505 142.735 147.915 143.255 ;
        RECT 148.395 143.245 148.655 143.725 ;
        RECT 148.085 142.555 148.315 142.985 ;
        RECT 146.525 142.385 148.315 142.555 ;
        RECT 146.525 142.020 146.775 142.385 ;
        RECT 146.945 142.025 147.275 142.215 ;
        RECT 147.495 142.090 148.210 142.385 ;
        RECT 148.485 142.215 148.655 143.245 ;
        RECT 148.845 143.085 149.085 143.895 ;
        RECT 149.255 143.085 149.585 143.725 ;
        RECT 149.755 143.085 150.025 143.895 ;
        RECT 150.205 143.095 150.900 143.725 ;
        RECT 151.105 143.095 151.415 143.895 ;
        RECT 151.585 143.170 151.875 143.895 ;
        RECT 152.135 143.345 152.305 143.725 ;
        RECT 152.485 143.515 152.815 143.895 ;
        RECT 152.135 143.175 152.800 143.345 ;
        RECT 152.995 143.220 153.255 143.725 ;
        RECT 148.825 142.655 149.175 142.905 ;
        RECT 149.345 142.485 149.515 143.085 ;
        RECT 149.685 142.655 150.035 142.905 ;
        RECT 150.225 142.655 150.560 142.905 ;
        RECT 150.730 142.495 150.900 143.095 ;
        RECT 151.070 142.655 151.405 142.925 ;
        RECT 152.065 142.625 152.395 142.995 ;
        RECT 152.630 142.920 152.800 143.175 ;
        RECT 152.630 142.590 152.915 142.920 ;
        RECT 146.945 141.850 147.140 142.025 ;
        RECT 146.525 141.345 147.140 141.850 ;
        RECT 147.310 141.515 147.785 141.855 ;
        RECT 147.955 141.345 148.170 141.890 ;
        RECT 148.380 141.515 148.655 142.215 ;
        RECT 148.835 142.315 149.515 142.485 ;
        RECT 148.835 141.530 149.165 142.315 ;
        RECT 149.695 141.345 150.025 142.485 ;
        RECT 150.205 141.345 150.465 142.485 ;
        RECT 150.635 141.515 150.965 142.495 ;
        RECT 151.135 141.345 151.415 142.485 ;
        RECT 151.585 141.345 151.875 142.510 ;
        RECT 152.630 142.445 152.800 142.590 ;
        RECT 152.135 142.275 152.800 142.445 ;
        RECT 153.085 142.420 153.255 143.220 ;
        RECT 153.425 143.125 155.095 143.895 ;
        RECT 155.725 143.145 156.935 143.895 ;
        RECT 153.425 142.605 154.175 143.125 ;
        RECT 154.345 142.435 155.095 142.955 ;
        RECT 152.135 141.515 152.305 142.275 ;
        RECT 152.485 141.345 152.815 142.105 ;
        RECT 152.985 141.515 153.255 142.420 ;
        RECT 153.425 141.345 155.095 142.435 ;
        RECT 155.725 142.435 156.245 142.975 ;
        RECT 156.415 142.605 156.935 143.145 ;
        RECT 155.725 141.345 156.935 142.435 ;
        RECT 22.700 141.175 157.020 141.345 ;
        RECT 22.785 140.085 23.995 141.175 ;
        RECT 24.165 140.085 25.835 141.175 ;
        RECT 22.785 139.375 23.305 139.915 ;
        RECT 23.475 139.545 23.995 140.085 ;
        RECT 24.165 139.395 24.915 139.915 ;
        RECT 25.085 139.565 25.835 140.085 ;
        RECT 26.465 140.305 26.740 141.005 ;
        RECT 26.950 140.630 27.165 141.175 ;
        RECT 27.335 140.665 27.810 141.005 ;
        RECT 27.980 140.670 28.595 141.175 ;
        RECT 27.980 140.495 28.175 140.670 ;
        RECT 22.785 138.625 23.995 139.375 ;
        RECT 24.165 138.625 25.835 139.395 ;
        RECT 26.465 139.275 26.635 140.305 ;
        RECT 26.910 140.135 27.625 140.430 ;
        RECT 27.845 140.305 28.175 140.495 ;
        RECT 28.345 140.135 28.595 140.500 ;
        RECT 26.805 139.965 28.595 140.135 ;
        RECT 26.805 139.535 27.035 139.965 ;
        RECT 26.465 138.795 26.725 139.275 ;
        RECT 27.205 139.265 27.615 139.785 ;
        RECT 26.895 138.625 27.225 139.085 ;
        RECT 27.415 138.845 27.615 139.265 ;
        RECT 27.785 139.110 28.040 139.965 ;
        RECT 28.835 139.785 29.005 141.005 ;
        RECT 29.255 140.665 29.515 141.175 ;
        RECT 30.145 140.620 30.750 141.175 ;
        RECT 30.925 140.665 31.405 141.005 ;
        RECT 31.575 140.630 31.830 141.175 ;
        RECT 30.145 140.520 30.760 140.620 ;
        RECT 30.575 140.495 30.760 140.520 ;
        RECT 28.210 139.535 29.005 139.785 ;
        RECT 29.175 139.615 29.515 140.495 ;
        RECT 30.145 139.900 30.405 140.350 ;
        RECT 30.575 140.250 30.905 140.495 ;
        RECT 31.075 140.175 31.830 140.425 ;
        RECT 32.000 140.305 32.275 141.005 ;
        RECT 32.445 140.665 32.705 141.175 ;
        RECT 31.060 140.140 31.830 140.175 ;
        RECT 31.045 140.130 31.830 140.140 ;
        RECT 31.040 140.115 31.935 140.130 ;
        RECT 31.020 140.100 31.935 140.115 ;
        RECT 31.000 140.090 31.935 140.100 ;
        RECT 30.975 140.080 31.935 140.090 ;
        RECT 30.905 140.050 31.935 140.080 ;
        RECT 30.885 140.020 31.935 140.050 ;
        RECT 30.865 139.990 31.935 140.020 ;
        RECT 30.835 139.965 31.935 139.990 ;
        RECT 30.800 139.930 31.935 139.965 ;
        RECT 30.770 139.925 31.935 139.930 ;
        RECT 30.770 139.920 31.160 139.925 ;
        RECT 30.770 139.910 31.135 139.920 ;
        RECT 30.770 139.905 31.120 139.910 ;
        RECT 30.770 139.900 31.105 139.905 ;
        RECT 30.145 139.895 31.105 139.900 ;
        RECT 30.145 139.885 31.095 139.895 ;
        RECT 30.145 139.880 31.085 139.885 ;
        RECT 30.145 139.870 31.075 139.880 ;
        RECT 30.145 139.860 31.070 139.870 ;
        RECT 30.145 139.855 31.065 139.860 ;
        RECT 30.145 139.840 31.055 139.855 ;
        RECT 30.145 139.825 31.050 139.840 ;
        RECT 30.145 139.800 31.040 139.825 ;
        RECT 30.145 139.730 31.035 139.800 ;
        RECT 28.755 139.445 29.005 139.535 ;
        RECT 27.785 138.845 28.575 139.110 ;
        RECT 28.755 139.025 29.085 139.445 ;
        RECT 29.255 138.625 29.515 139.445 ;
        RECT 30.145 139.175 30.695 139.560 ;
        RECT 30.865 139.005 31.035 139.730 ;
        RECT 30.145 138.835 31.035 139.005 ;
        RECT 31.205 139.330 31.535 139.755 ;
        RECT 31.705 139.530 31.935 139.925 ;
        RECT 31.205 138.845 31.425 139.330 ;
        RECT 32.105 139.275 32.275 140.305 ;
        RECT 32.445 139.615 32.785 140.495 ;
        RECT 32.955 139.785 33.125 141.005 ;
        RECT 33.365 140.670 33.980 141.175 ;
        RECT 33.365 140.135 33.615 140.500 ;
        RECT 33.785 140.495 33.980 140.670 ;
        RECT 34.150 140.665 34.625 141.005 ;
        RECT 34.795 140.630 35.010 141.175 ;
        RECT 33.785 140.305 34.115 140.495 ;
        RECT 34.335 140.135 35.050 140.430 ;
        RECT 35.220 140.305 35.495 141.005 ;
        RECT 33.365 139.965 35.155 140.135 ;
        RECT 32.955 139.535 33.750 139.785 ;
        RECT 32.955 139.445 33.205 139.535 ;
        RECT 31.595 138.625 31.845 139.165 ;
        RECT 32.015 138.795 32.275 139.275 ;
        RECT 32.445 138.625 32.705 139.445 ;
        RECT 32.875 139.025 33.205 139.445 ;
        RECT 33.920 139.110 34.175 139.965 ;
        RECT 33.385 138.845 34.175 139.110 ;
        RECT 34.345 139.265 34.755 139.785 ;
        RECT 34.925 139.535 35.155 139.965 ;
        RECT 35.325 139.275 35.495 140.305 ;
        RECT 35.665 140.010 35.955 141.175 ;
        RECT 36.185 140.115 36.515 140.960 ;
        RECT 36.685 140.165 36.855 141.175 ;
        RECT 37.025 140.445 37.365 141.005 ;
        RECT 37.595 140.675 37.910 141.175 ;
        RECT 38.090 140.705 38.975 140.875 ;
        RECT 36.125 140.035 36.515 140.115 ;
        RECT 37.025 140.070 37.920 140.445 ;
        RECT 36.125 139.985 36.340 140.035 ;
        RECT 36.125 139.405 36.295 139.985 ;
        RECT 37.025 139.865 37.215 140.070 ;
        RECT 38.090 139.865 38.260 140.705 ;
        RECT 39.200 140.675 39.450 141.005 ;
        RECT 36.465 139.535 37.215 139.865 ;
        RECT 37.385 139.535 38.260 139.865 ;
        RECT 36.125 139.365 36.350 139.405 ;
        RECT 37.015 139.365 37.215 139.535 ;
        RECT 34.345 138.845 34.545 139.265 ;
        RECT 34.735 138.625 35.065 139.085 ;
        RECT 35.235 138.795 35.495 139.275 ;
        RECT 35.665 138.625 35.955 139.350 ;
        RECT 36.125 139.280 36.505 139.365 ;
        RECT 36.175 138.845 36.505 139.280 ;
        RECT 36.675 138.625 36.845 139.235 ;
        RECT 37.015 138.840 37.345 139.365 ;
        RECT 37.605 138.625 37.815 139.155 ;
        RECT 38.090 139.075 38.260 139.535 ;
        RECT 38.430 139.575 38.750 140.535 ;
        RECT 38.920 139.785 39.110 140.505 ;
        RECT 39.280 139.605 39.450 140.675 ;
        RECT 39.620 140.375 39.790 141.175 ;
        RECT 39.960 140.730 41.065 140.900 ;
        RECT 39.960 140.115 40.130 140.730 ;
        RECT 41.275 140.580 41.525 141.005 ;
        RECT 41.695 140.715 41.960 141.175 ;
        RECT 40.300 140.195 40.830 140.560 ;
        RECT 41.275 140.450 41.580 140.580 ;
        RECT 39.620 140.025 40.130 140.115 ;
        RECT 39.620 139.855 40.490 140.025 ;
        RECT 39.620 139.785 39.790 139.855 ;
        RECT 39.910 139.605 40.110 139.635 ;
        RECT 38.430 139.245 38.895 139.575 ;
        RECT 39.280 139.305 40.110 139.605 ;
        RECT 39.280 139.075 39.450 139.305 ;
        RECT 38.090 138.905 38.875 139.075 ;
        RECT 39.045 138.905 39.450 139.075 ;
        RECT 39.630 138.625 40.000 139.125 ;
        RECT 40.320 139.075 40.490 139.855 ;
        RECT 40.660 139.495 40.830 140.195 ;
        RECT 41.000 139.665 41.240 140.260 ;
        RECT 40.660 139.275 41.185 139.495 ;
        RECT 41.410 139.345 41.580 140.450 ;
        RECT 41.355 139.215 41.580 139.345 ;
        RECT 41.750 139.255 42.030 140.205 ;
        RECT 41.355 139.075 41.525 139.215 ;
        RECT 40.320 138.905 40.995 139.075 ;
        RECT 41.190 138.905 41.525 139.075 ;
        RECT 41.695 138.625 41.945 139.085 ;
        RECT 42.200 138.885 42.385 141.005 ;
        RECT 42.555 140.675 42.885 141.175 ;
        RECT 43.055 140.505 43.225 141.005 ;
        RECT 42.560 140.335 43.225 140.505 ;
        RECT 42.560 139.345 42.790 140.335 ;
        RECT 42.960 139.515 43.310 140.165 ;
        RECT 44.445 140.035 44.675 141.175 ;
        RECT 44.845 140.025 45.175 141.005 ;
        RECT 45.345 140.035 45.555 141.175 ;
        RECT 44.425 139.615 44.755 139.865 ;
        RECT 42.560 139.175 43.225 139.345 ;
        RECT 42.555 138.625 42.885 139.005 ;
        RECT 43.055 138.885 43.225 139.175 ;
        RECT 44.445 138.625 44.675 139.445 ;
        RECT 44.925 139.425 45.175 140.025 ;
        RECT 44.845 138.795 45.175 139.425 ;
        RECT 45.345 138.625 45.555 139.445 ;
        RECT 45.795 138.795 46.055 141.005 ;
        RECT 46.225 140.375 47.035 141.175 ;
        RECT 47.205 140.205 47.535 141.005 ;
        RECT 47.720 140.375 48.460 141.175 ;
        RECT 48.630 140.205 48.880 141.005 ;
        RECT 46.395 140.035 48.880 140.205 ;
        RECT 46.395 139.865 46.565 140.035 ;
        RECT 49.050 139.865 49.235 140.955 ;
        RECT 49.430 140.375 49.755 141.175 ;
        RECT 46.225 139.535 46.565 139.865 ;
        RECT 46.965 139.615 47.445 139.865 ;
        RECT 46.395 139.445 46.565 139.535 ;
        RECT 46.395 139.275 47.065 139.445 ;
        RECT 46.235 138.625 46.545 139.105 ;
        RECT 46.725 138.795 47.065 139.275 ;
        RECT 47.235 138.930 47.445 139.615 ;
        RECT 47.625 138.930 47.895 139.865 ;
        RECT 48.145 139.535 48.405 139.865 ;
        RECT 48.750 139.615 49.235 139.865 ;
        RECT 49.405 139.615 49.735 140.200 ;
        RECT 49.925 140.085 51.135 141.175 ;
        RECT 48.145 138.930 48.390 139.535 ;
        RECT 48.570 139.245 49.755 139.415 ;
        RECT 48.570 138.795 48.860 139.245 ;
        RECT 49.030 138.625 49.320 139.075 ;
        RECT 49.490 138.795 49.755 139.245 ;
        RECT 49.925 139.375 50.445 139.915 ;
        RECT 50.615 139.545 51.135 140.085 ;
        RECT 49.925 138.625 51.135 139.375 ;
        RECT 51.315 138.805 51.575 140.995 ;
        RECT 51.745 140.445 52.085 141.175 ;
        RECT 52.265 140.265 52.535 140.995 ;
        RECT 51.765 140.045 52.535 140.265 ;
        RECT 52.715 140.285 52.945 140.995 ;
        RECT 53.115 140.465 53.445 141.175 ;
        RECT 53.615 140.285 53.875 140.995 ;
        RECT 52.715 140.045 53.875 140.285 ;
        RECT 54.125 140.115 54.455 140.960 ;
        RECT 54.625 140.165 54.795 141.175 ;
        RECT 54.965 140.445 55.305 141.005 ;
        RECT 55.535 140.675 55.850 141.175 ;
        RECT 56.030 140.705 56.915 140.875 ;
        RECT 51.765 139.375 52.055 140.045 ;
        RECT 54.065 140.035 54.455 140.115 ;
        RECT 54.965 140.070 55.860 140.445 ;
        RECT 54.065 139.985 54.280 140.035 ;
        RECT 52.235 139.555 52.700 139.865 ;
        RECT 52.880 139.555 53.405 139.865 ;
        RECT 51.765 139.175 52.995 139.375 ;
        RECT 51.835 138.625 52.505 138.995 ;
        RECT 52.685 138.805 52.995 139.175 ;
        RECT 53.175 138.915 53.405 139.555 ;
        RECT 53.585 139.535 53.885 139.865 ;
        RECT 54.065 139.405 54.235 139.985 ;
        RECT 54.965 139.865 55.155 140.070 ;
        RECT 56.030 139.865 56.200 140.705 ;
        RECT 57.140 140.675 57.390 141.005 ;
        RECT 54.405 139.535 55.155 139.865 ;
        RECT 55.325 139.535 56.200 139.865 ;
        RECT 54.065 139.365 54.290 139.405 ;
        RECT 54.955 139.365 55.155 139.535 ;
        RECT 53.585 138.625 53.875 139.355 ;
        RECT 54.065 139.280 54.445 139.365 ;
        RECT 54.115 138.845 54.445 139.280 ;
        RECT 54.615 138.625 54.785 139.235 ;
        RECT 54.955 138.840 55.285 139.365 ;
        RECT 55.545 138.625 55.755 139.155 ;
        RECT 56.030 139.075 56.200 139.535 ;
        RECT 56.370 139.575 56.690 140.535 ;
        RECT 56.860 139.785 57.050 140.505 ;
        RECT 57.220 139.605 57.390 140.675 ;
        RECT 57.560 140.375 57.730 141.175 ;
        RECT 57.900 140.730 59.005 140.900 ;
        RECT 57.900 140.115 58.070 140.730 ;
        RECT 59.215 140.580 59.465 141.005 ;
        RECT 59.635 140.715 59.900 141.175 ;
        RECT 58.240 140.195 58.770 140.560 ;
        RECT 59.215 140.450 59.520 140.580 ;
        RECT 57.560 140.025 58.070 140.115 ;
        RECT 57.560 139.855 58.430 140.025 ;
        RECT 57.560 139.785 57.730 139.855 ;
        RECT 57.850 139.605 58.050 139.635 ;
        RECT 56.370 139.245 56.835 139.575 ;
        RECT 57.220 139.305 58.050 139.605 ;
        RECT 57.220 139.075 57.390 139.305 ;
        RECT 56.030 138.905 56.815 139.075 ;
        RECT 56.985 138.905 57.390 139.075 ;
        RECT 57.570 138.625 57.940 139.125 ;
        RECT 58.260 139.075 58.430 139.855 ;
        RECT 58.600 139.495 58.770 140.195 ;
        RECT 58.940 139.665 59.180 140.260 ;
        RECT 58.600 139.275 59.125 139.495 ;
        RECT 59.350 139.345 59.520 140.450 ;
        RECT 59.295 139.215 59.520 139.345 ;
        RECT 59.690 139.255 59.970 140.205 ;
        RECT 59.295 139.075 59.465 139.215 ;
        RECT 58.260 138.905 58.935 139.075 ;
        RECT 59.130 138.905 59.465 139.075 ;
        RECT 59.635 138.625 59.885 139.085 ;
        RECT 60.140 138.885 60.325 141.005 ;
        RECT 60.495 140.675 60.825 141.175 ;
        RECT 60.995 140.505 61.165 141.005 ;
        RECT 60.500 140.335 61.165 140.505 ;
        RECT 60.500 139.345 60.730 140.335 ;
        RECT 60.900 139.515 61.250 140.165 ;
        RECT 61.425 140.010 61.715 141.175 ;
        RECT 61.885 140.085 63.555 141.175 ;
        RECT 63.815 140.505 63.985 141.005 ;
        RECT 64.155 140.675 64.485 141.175 ;
        RECT 63.815 140.335 64.480 140.505 ;
        RECT 61.885 139.395 62.635 139.915 ;
        RECT 62.805 139.565 63.555 140.085 ;
        RECT 63.730 139.515 64.080 140.165 ;
        RECT 60.500 139.175 61.165 139.345 ;
        RECT 60.495 138.625 60.825 139.005 ;
        RECT 60.995 138.885 61.165 139.175 ;
        RECT 61.425 138.625 61.715 139.350 ;
        RECT 61.885 138.625 63.555 139.395 ;
        RECT 64.250 139.345 64.480 140.335 ;
        RECT 63.815 139.175 64.480 139.345 ;
        RECT 63.815 138.885 63.985 139.175 ;
        RECT 64.155 138.625 64.485 139.005 ;
        RECT 64.655 138.885 64.840 141.005 ;
        RECT 65.080 140.715 65.345 141.175 ;
        RECT 65.515 140.580 65.765 141.005 ;
        RECT 65.975 140.730 67.080 140.900 ;
        RECT 65.460 140.450 65.765 140.580 ;
        RECT 65.010 139.255 65.290 140.205 ;
        RECT 65.460 139.345 65.630 140.450 ;
        RECT 65.800 139.665 66.040 140.260 ;
        RECT 66.210 140.195 66.740 140.560 ;
        RECT 66.210 139.495 66.380 140.195 ;
        RECT 66.910 140.115 67.080 140.730 ;
        RECT 67.250 140.375 67.420 141.175 ;
        RECT 67.590 140.675 67.840 141.005 ;
        RECT 68.065 140.705 68.950 140.875 ;
        RECT 66.910 140.025 67.420 140.115 ;
        RECT 65.460 139.215 65.685 139.345 ;
        RECT 65.855 139.275 66.380 139.495 ;
        RECT 66.550 139.855 67.420 140.025 ;
        RECT 65.095 138.625 65.345 139.085 ;
        RECT 65.515 139.075 65.685 139.215 ;
        RECT 66.550 139.075 66.720 139.855 ;
        RECT 67.250 139.785 67.420 139.855 ;
        RECT 66.930 139.605 67.130 139.635 ;
        RECT 67.590 139.605 67.760 140.675 ;
        RECT 67.930 139.785 68.120 140.505 ;
        RECT 66.930 139.305 67.760 139.605 ;
        RECT 68.290 139.575 68.610 140.535 ;
        RECT 65.515 138.905 65.850 139.075 ;
        RECT 66.045 138.905 66.720 139.075 ;
        RECT 67.040 138.625 67.410 139.125 ;
        RECT 67.590 139.075 67.760 139.305 ;
        RECT 68.145 139.245 68.610 139.575 ;
        RECT 68.780 139.865 68.950 140.705 ;
        RECT 69.130 140.675 69.445 141.175 ;
        RECT 69.675 140.445 70.015 141.005 ;
        RECT 69.120 140.070 70.015 140.445 ;
        RECT 70.185 140.165 70.355 141.175 ;
        RECT 69.825 139.865 70.015 140.070 ;
        RECT 70.525 140.115 70.855 140.960 ;
        RECT 70.525 140.035 70.915 140.115 ;
        RECT 71.125 140.035 71.355 141.175 ;
        RECT 70.700 139.985 70.915 140.035 ;
        RECT 71.525 140.025 71.855 141.005 ;
        RECT 72.025 140.035 72.235 141.175 ;
        RECT 73.405 140.665 73.705 141.175 ;
        RECT 73.875 140.665 74.255 140.835 ;
        RECT 74.835 140.665 75.465 141.175 ;
        RECT 73.875 140.495 74.045 140.665 ;
        RECT 75.635 140.495 75.965 141.005 ;
        RECT 76.135 140.665 76.435 141.175 ;
        RECT 76.605 140.740 81.950 141.175 ;
        RECT 73.385 140.295 74.045 140.495 ;
        RECT 74.215 140.325 76.435 140.495 ;
        RECT 68.780 139.535 69.655 139.865 ;
        RECT 69.825 139.535 70.575 139.865 ;
        RECT 68.780 139.075 68.950 139.535 ;
        RECT 69.825 139.365 70.025 139.535 ;
        RECT 70.745 139.405 70.915 139.985 ;
        RECT 71.105 139.615 71.435 139.865 ;
        RECT 70.690 139.365 70.915 139.405 ;
        RECT 67.590 138.905 67.995 139.075 ;
        RECT 68.165 138.905 68.950 139.075 ;
        RECT 69.225 138.625 69.435 139.155 ;
        RECT 69.695 138.840 70.025 139.365 ;
        RECT 70.535 139.280 70.915 139.365 ;
        RECT 70.195 138.625 70.365 139.235 ;
        RECT 70.535 138.845 70.865 139.280 ;
        RECT 71.125 138.625 71.355 139.445 ;
        RECT 71.605 139.425 71.855 140.025 ;
        RECT 71.525 138.795 71.855 139.425 ;
        RECT 72.025 138.625 72.235 139.445 ;
        RECT 73.385 139.365 73.555 140.295 ;
        RECT 74.215 140.125 74.385 140.325 ;
        RECT 73.725 139.955 74.385 140.125 ;
        RECT 74.555 139.985 76.095 140.155 ;
        RECT 73.725 139.535 73.895 139.955 ;
        RECT 74.555 139.785 74.725 139.985 ;
        RECT 74.125 139.615 74.725 139.785 ;
        RECT 74.895 139.615 75.590 139.815 ;
        RECT 75.850 139.535 76.095 139.985 ;
        RECT 74.215 139.365 75.125 139.445 ;
        RECT 73.385 138.885 73.705 139.365 ;
        RECT 73.875 139.275 75.125 139.365 ;
        RECT 73.875 139.195 74.385 139.275 ;
        RECT 73.875 138.795 74.105 139.195 ;
        RECT 74.275 138.625 74.625 139.015 ;
        RECT 74.795 138.795 75.125 139.275 ;
        RECT 75.295 138.625 75.465 139.445 ;
        RECT 76.265 139.365 76.435 140.325 ;
        RECT 75.970 138.820 76.435 139.365 ;
        RECT 78.190 139.170 78.530 140.000 ;
        RECT 80.010 139.490 80.360 140.740 ;
        RECT 76.605 138.625 81.950 139.170 ;
        RECT 83.055 138.805 83.315 140.995 ;
        RECT 83.485 140.445 83.825 141.175 ;
        RECT 84.005 140.265 84.275 140.995 ;
        RECT 83.505 140.045 84.275 140.265 ;
        RECT 84.455 140.285 84.685 140.995 ;
        RECT 84.855 140.465 85.185 141.175 ;
        RECT 85.355 140.285 85.615 140.995 ;
        RECT 84.455 140.045 85.615 140.285 ;
        RECT 85.805 140.085 87.015 141.175 ;
        RECT 83.505 139.375 83.795 140.045 ;
        RECT 83.975 139.555 84.440 139.865 ;
        RECT 84.620 139.555 85.145 139.865 ;
        RECT 83.505 139.175 84.735 139.375 ;
        RECT 83.575 138.625 84.245 138.995 ;
        RECT 84.425 138.805 84.735 139.175 ;
        RECT 84.915 138.915 85.145 139.555 ;
        RECT 85.325 139.535 85.625 139.865 ;
        RECT 85.805 139.375 86.325 139.915 ;
        RECT 86.495 139.545 87.015 140.085 ;
        RECT 87.185 140.010 87.475 141.175 ;
        RECT 88.655 140.505 88.825 141.005 ;
        RECT 88.995 140.675 89.325 141.175 ;
        RECT 88.655 140.335 89.320 140.505 ;
        RECT 88.570 139.515 88.920 140.165 ;
        RECT 85.325 138.625 85.615 139.355 ;
        RECT 85.805 138.625 87.015 139.375 ;
        RECT 87.185 138.625 87.475 139.350 ;
        RECT 89.090 139.345 89.320 140.335 ;
        RECT 88.655 139.175 89.320 139.345 ;
        RECT 88.655 138.885 88.825 139.175 ;
        RECT 88.995 138.625 89.325 139.005 ;
        RECT 89.495 138.885 89.680 141.005 ;
        RECT 89.920 140.715 90.185 141.175 ;
        RECT 90.355 140.580 90.605 141.005 ;
        RECT 90.815 140.730 91.920 140.900 ;
        RECT 90.300 140.450 90.605 140.580 ;
        RECT 89.850 139.255 90.130 140.205 ;
        RECT 90.300 139.345 90.470 140.450 ;
        RECT 90.640 139.665 90.880 140.260 ;
        RECT 91.050 140.195 91.580 140.560 ;
        RECT 91.050 139.495 91.220 140.195 ;
        RECT 91.750 140.115 91.920 140.730 ;
        RECT 92.090 140.375 92.260 141.175 ;
        RECT 92.430 140.675 92.680 141.005 ;
        RECT 92.905 140.705 93.790 140.875 ;
        RECT 91.750 140.025 92.260 140.115 ;
        RECT 90.300 139.215 90.525 139.345 ;
        RECT 90.695 139.275 91.220 139.495 ;
        RECT 91.390 139.855 92.260 140.025 ;
        RECT 89.935 138.625 90.185 139.085 ;
        RECT 90.355 139.075 90.525 139.215 ;
        RECT 91.390 139.075 91.560 139.855 ;
        RECT 92.090 139.785 92.260 139.855 ;
        RECT 91.770 139.605 91.970 139.635 ;
        RECT 92.430 139.605 92.600 140.675 ;
        RECT 92.770 139.785 92.960 140.505 ;
        RECT 91.770 139.305 92.600 139.605 ;
        RECT 93.130 139.575 93.450 140.535 ;
        RECT 90.355 138.905 90.690 139.075 ;
        RECT 90.885 138.905 91.560 139.075 ;
        RECT 91.880 138.625 92.250 139.125 ;
        RECT 92.430 139.075 92.600 139.305 ;
        RECT 92.985 139.245 93.450 139.575 ;
        RECT 93.620 139.865 93.790 140.705 ;
        RECT 93.970 140.675 94.285 141.175 ;
        RECT 94.515 140.445 94.855 141.005 ;
        RECT 93.960 140.070 94.855 140.445 ;
        RECT 95.025 140.165 95.195 141.175 ;
        RECT 94.665 139.865 94.855 140.070 ;
        RECT 95.365 140.115 95.695 140.960 ;
        RECT 95.365 140.035 95.755 140.115 ;
        RECT 95.540 139.985 95.755 140.035 ;
        RECT 93.620 139.535 94.495 139.865 ;
        RECT 94.665 139.535 95.415 139.865 ;
        RECT 93.620 139.075 93.790 139.535 ;
        RECT 94.665 139.365 94.865 139.535 ;
        RECT 95.585 139.405 95.755 139.985 ;
        RECT 95.530 139.365 95.755 139.405 ;
        RECT 92.430 138.905 92.835 139.075 ;
        RECT 93.005 138.905 93.790 139.075 ;
        RECT 94.065 138.625 94.275 139.155 ;
        RECT 94.535 138.840 94.865 139.365 ;
        RECT 95.375 139.280 95.755 139.365 ;
        RECT 95.925 140.035 96.310 141.005 ;
        RECT 96.480 140.715 96.805 141.175 ;
        RECT 97.325 140.545 97.605 141.005 ;
        RECT 96.480 140.325 97.605 140.545 ;
        RECT 95.925 139.365 96.205 140.035 ;
        RECT 96.480 139.865 96.930 140.325 ;
        RECT 97.795 140.155 98.195 141.005 ;
        RECT 98.595 140.715 98.865 141.175 ;
        RECT 99.035 140.545 99.320 141.005 ;
        RECT 96.375 139.535 96.930 139.865 ;
        RECT 97.100 139.595 98.195 140.155 ;
        RECT 96.480 139.425 96.930 139.535 ;
        RECT 95.035 138.625 95.205 139.235 ;
        RECT 95.375 138.845 95.705 139.280 ;
        RECT 95.925 138.795 96.310 139.365 ;
        RECT 96.480 139.255 97.605 139.425 ;
        RECT 96.480 138.625 96.805 139.085 ;
        RECT 97.325 138.795 97.605 139.255 ;
        RECT 97.795 138.795 98.195 139.595 ;
        RECT 98.365 140.325 99.320 140.545 ;
        RECT 98.365 139.425 98.575 140.325 ;
        RECT 98.745 139.595 99.435 140.155 ;
        RECT 99.605 140.085 101.275 141.175 ;
        RECT 101.505 140.115 101.835 140.960 ;
        RECT 102.005 140.165 102.175 141.175 ;
        RECT 102.345 140.445 102.685 141.005 ;
        RECT 102.915 140.675 103.230 141.175 ;
        RECT 103.410 140.705 104.295 140.875 ;
        RECT 98.365 139.255 99.320 139.425 ;
        RECT 98.595 138.625 98.865 139.085 ;
        RECT 99.035 138.795 99.320 139.255 ;
        RECT 99.605 139.395 100.355 139.915 ;
        RECT 100.525 139.565 101.275 140.085 ;
        RECT 101.445 140.035 101.835 140.115 ;
        RECT 102.345 140.070 103.240 140.445 ;
        RECT 101.445 139.985 101.660 140.035 ;
        RECT 101.445 139.405 101.615 139.985 ;
        RECT 102.345 139.865 102.535 140.070 ;
        RECT 103.410 139.865 103.580 140.705 ;
        RECT 104.520 140.675 104.770 141.005 ;
        RECT 101.785 139.535 102.535 139.865 ;
        RECT 102.705 139.535 103.580 139.865 ;
        RECT 99.605 138.625 101.275 139.395 ;
        RECT 101.445 139.365 101.670 139.405 ;
        RECT 102.335 139.365 102.535 139.535 ;
        RECT 101.445 139.280 101.825 139.365 ;
        RECT 101.495 138.845 101.825 139.280 ;
        RECT 101.995 138.625 102.165 139.235 ;
        RECT 102.335 138.840 102.665 139.365 ;
        RECT 102.925 138.625 103.135 139.155 ;
        RECT 103.410 139.075 103.580 139.535 ;
        RECT 103.750 139.575 104.070 140.535 ;
        RECT 104.240 139.785 104.430 140.505 ;
        RECT 104.600 139.605 104.770 140.675 ;
        RECT 104.940 140.375 105.110 141.175 ;
        RECT 105.280 140.730 106.385 140.900 ;
        RECT 105.280 140.115 105.450 140.730 ;
        RECT 106.595 140.580 106.845 141.005 ;
        RECT 107.015 140.715 107.280 141.175 ;
        RECT 105.620 140.195 106.150 140.560 ;
        RECT 106.595 140.450 106.900 140.580 ;
        RECT 104.940 140.025 105.450 140.115 ;
        RECT 104.940 139.855 105.810 140.025 ;
        RECT 104.940 139.785 105.110 139.855 ;
        RECT 105.230 139.605 105.430 139.635 ;
        RECT 103.750 139.245 104.215 139.575 ;
        RECT 104.600 139.305 105.430 139.605 ;
        RECT 104.600 139.075 104.770 139.305 ;
        RECT 103.410 138.905 104.195 139.075 ;
        RECT 104.365 138.905 104.770 139.075 ;
        RECT 104.950 138.625 105.320 139.125 ;
        RECT 105.640 139.075 105.810 139.855 ;
        RECT 105.980 139.495 106.150 140.195 ;
        RECT 106.320 139.665 106.560 140.260 ;
        RECT 105.980 139.275 106.505 139.495 ;
        RECT 106.730 139.345 106.900 140.450 ;
        RECT 106.675 139.215 106.900 139.345 ;
        RECT 107.070 139.255 107.350 140.205 ;
        RECT 106.675 139.075 106.845 139.215 ;
        RECT 105.640 138.905 106.315 139.075 ;
        RECT 106.510 138.905 106.845 139.075 ;
        RECT 107.015 138.625 107.265 139.085 ;
        RECT 107.520 138.885 107.705 141.005 ;
        RECT 107.875 140.675 108.205 141.175 ;
        RECT 108.375 140.505 108.545 141.005 ;
        RECT 107.880 140.335 108.545 140.505 ;
        RECT 109.730 140.785 110.065 141.005 ;
        RECT 111.070 140.795 111.425 141.175 ;
        RECT 107.880 139.345 108.110 140.335 ;
        RECT 109.730 140.165 109.985 140.785 ;
        RECT 110.235 140.625 110.465 140.665 ;
        RECT 111.595 140.625 111.845 141.005 ;
        RECT 110.235 140.425 111.845 140.625 ;
        RECT 110.235 140.335 110.420 140.425 ;
        RECT 111.010 140.415 111.845 140.425 ;
        RECT 112.095 140.395 112.345 141.175 ;
        RECT 112.515 140.325 112.775 141.005 ;
        RECT 110.575 140.225 110.905 140.255 ;
        RECT 110.575 140.165 112.375 140.225 ;
        RECT 108.280 139.515 108.630 140.165 ;
        RECT 109.730 140.055 112.435 140.165 ;
        RECT 109.730 139.995 110.905 140.055 ;
        RECT 112.235 140.020 112.435 140.055 ;
        RECT 109.725 139.615 110.215 139.815 ;
        RECT 110.405 139.615 110.880 139.825 ;
        RECT 107.880 139.175 108.545 139.345 ;
        RECT 107.875 138.625 108.205 139.005 ;
        RECT 108.375 138.885 108.545 139.175 ;
        RECT 109.730 138.625 110.185 139.390 ;
        RECT 110.660 139.215 110.880 139.615 ;
        RECT 111.125 139.615 111.455 139.825 ;
        RECT 111.125 139.215 111.335 139.615 ;
        RECT 111.625 139.580 112.035 139.885 ;
        RECT 112.265 139.445 112.435 140.020 ;
        RECT 112.165 139.325 112.435 139.445 ;
        RECT 111.590 139.280 112.435 139.325 ;
        RECT 111.590 139.155 112.345 139.280 ;
        RECT 111.590 139.005 111.760 139.155 ;
        RECT 112.605 139.135 112.775 140.325 ;
        RECT 112.945 140.010 113.235 141.175 ;
        RECT 114.415 140.505 114.585 141.005 ;
        RECT 114.755 140.675 115.085 141.175 ;
        RECT 114.415 140.335 115.080 140.505 ;
        RECT 114.330 139.515 114.680 140.165 ;
        RECT 112.545 139.125 112.775 139.135 ;
        RECT 110.460 138.795 111.760 139.005 ;
        RECT 112.015 138.625 112.345 138.985 ;
        RECT 112.515 138.795 112.775 139.125 ;
        RECT 112.945 138.625 113.235 139.350 ;
        RECT 114.850 139.345 115.080 140.335 ;
        RECT 114.415 139.175 115.080 139.345 ;
        RECT 114.415 138.885 114.585 139.175 ;
        RECT 114.755 138.625 115.085 139.005 ;
        RECT 115.255 138.885 115.440 141.005 ;
        RECT 115.680 140.715 115.945 141.175 ;
        RECT 116.115 140.580 116.365 141.005 ;
        RECT 116.575 140.730 117.680 140.900 ;
        RECT 116.060 140.450 116.365 140.580 ;
        RECT 115.610 139.255 115.890 140.205 ;
        RECT 116.060 139.345 116.230 140.450 ;
        RECT 116.400 139.665 116.640 140.260 ;
        RECT 116.810 140.195 117.340 140.560 ;
        RECT 116.810 139.495 116.980 140.195 ;
        RECT 117.510 140.115 117.680 140.730 ;
        RECT 117.850 140.375 118.020 141.175 ;
        RECT 118.190 140.675 118.440 141.005 ;
        RECT 118.665 140.705 119.550 140.875 ;
        RECT 117.510 140.025 118.020 140.115 ;
        RECT 116.060 139.215 116.285 139.345 ;
        RECT 116.455 139.275 116.980 139.495 ;
        RECT 117.150 139.855 118.020 140.025 ;
        RECT 115.695 138.625 115.945 139.085 ;
        RECT 116.115 139.075 116.285 139.215 ;
        RECT 117.150 139.075 117.320 139.855 ;
        RECT 117.850 139.785 118.020 139.855 ;
        RECT 117.530 139.605 117.730 139.635 ;
        RECT 118.190 139.605 118.360 140.675 ;
        RECT 118.530 139.785 118.720 140.505 ;
        RECT 117.530 139.305 118.360 139.605 ;
        RECT 118.890 139.575 119.210 140.535 ;
        RECT 116.115 138.905 116.450 139.075 ;
        RECT 116.645 138.905 117.320 139.075 ;
        RECT 117.640 138.625 118.010 139.125 ;
        RECT 118.190 139.075 118.360 139.305 ;
        RECT 118.745 139.245 119.210 139.575 ;
        RECT 119.380 139.865 119.550 140.705 ;
        RECT 119.730 140.675 120.045 141.175 ;
        RECT 120.275 140.445 120.615 141.005 ;
        RECT 119.720 140.070 120.615 140.445 ;
        RECT 120.785 140.165 120.955 141.175 ;
        RECT 120.425 139.865 120.615 140.070 ;
        RECT 121.125 140.115 121.455 140.960 ;
        RECT 121.125 140.035 121.515 140.115 ;
        RECT 121.300 139.985 121.515 140.035 ;
        RECT 119.380 139.535 120.255 139.865 ;
        RECT 120.425 139.535 121.175 139.865 ;
        RECT 119.380 139.075 119.550 139.535 ;
        RECT 120.425 139.365 120.625 139.535 ;
        RECT 121.345 139.405 121.515 139.985 ;
        RECT 121.290 139.365 121.515 139.405 ;
        RECT 118.190 138.905 118.595 139.075 ;
        RECT 118.765 138.905 119.550 139.075 ;
        RECT 119.825 138.625 120.035 139.155 ;
        RECT 120.295 138.840 120.625 139.365 ;
        RECT 121.135 139.280 121.515 139.365 ;
        RECT 121.685 140.035 122.070 141.005 ;
        RECT 122.240 140.715 122.565 141.175 ;
        RECT 123.085 140.545 123.365 141.005 ;
        RECT 122.240 140.325 123.365 140.545 ;
        RECT 121.685 139.365 121.965 140.035 ;
        RECT 122.240 139.865 122.690 140.325 ;
        RECT 123.555 140.155 123.955 141.005 ;
        RECT 124.355 140.715 124.625 141.175 ;
        RECT 124.795 140.545 125.080 141.005 ;
        RECT 122.135 139.535 122.690 139.865 ;
        RECT 122.860 139.595 123.955 140.155 ;
        RECT 122.240 139.425 122.690 139.535 ;
        RECT 120.795 138.625 120.965 139.235 ;
        RECT 121.135 138.845 121.465 139.280 ;
        RECT 121.685 138.795 122.070 139.365 ;
        RECT 122.240 139.255 123.365 139.425 ;
        RECT 122.240 138.625 122.565 139.085 ;
        RECT 123.085 138.795 123.365 139.255 ;
        RECT 123.555 138.795 123.955 139.595 ;
        RECT 124.125 140.325 125.080 140.545 ;
        RECT 124.125 139.425 124.335 140.325 ;
        RECT 124.505 139.595 125.195 140.155 ;
        RECT 125.365 140.085 127.035 141.175 ;
        RECT 124.125 139.255 125.080 139.425 ;
        RECT 124.355 138.625 124.625 139.085 ;
        RECT 124.795 138.795 125.080 139.255 ;
        RECT 125.365 139.395 126.115 139.915 ;
        RECT 126.285 139.565 127.035 140.085 ;
        RECT 127.215 140.565 127.545 140.995 ;
        RECT 127.725 140.735 127.920 141.175 ;
        RECT 128.090 140.565 128.420 140.995 ;
        RECT 127.215 140.395 128.420 140.565 ;
        RECT 127.215 140.065 128.110 140.395 ;
        RECT 128.590 140.225 128.865 140.995 ;
        RECT 128.280 140.035 128.865 140.225 ;
        RECT 129.045 140.085 132.555 141.175 ;
        RECT 133.655 140.585 133.915 140.975 ;
        RECT 134.085 140.765 134.415 141.175 ;
        RECT 133.655 140.385 134.415 140.585 ;
        RECT 127.220 139.535 127.515 139.865 ;
        RECT 127.695 139.535 128.110 139.865 ;
        RECT 125.365 138.625 127.035 139.395 ;
        RECT 127.215 138.625 127.515 139.355 ;
        RECT 127.695 138.915 127.925 139.535 ;
        RECT 128.280 139.365 128.455 140.035 ;
        RECT 128.125 139.185 128.455 139.365 ;
        RECT 128.625 139.215 128.865 139.865 ;
        RECT 129.045 139.395 130.695 139.915 ;
        RECT 130.865 139.565 132.555 140.085 ;
        RECT 133.665 139.515 133.895 140.205 ;
        RECT 134.075 139.705 134.415 140.385 ;
        RECT 134.605 139.885 134.935 140.995 ;
        RECT 135.105 140.265 135.295 140.995 ;
        RECT 135.465 140.445 135.795 141.175 ;
        RECT 135.975 140.265 136.145 140.995 ;
        RECT 135.105 140.065 136.145 140.265 ;
        RECT 136.405 140.085 138.075 141.175 ;
        RECT 128.125 138.805 128.350 139.185 ;
        RECT 128.520 138.625 128.850 139.015 ;
        RECT 129.045 138.625 132.555 139.395 ;
        RECT 134.075 139.255 134.305 139.705 ;
        RECT 134.605 139.585 135.140 139.885 ;
        RECT 133.925 138.805 134.305 139.255 ;
        RECT 134.485 138.625 134.715 139.405 ;
        RECT 134.895 139.335 135.140 139.585 ;
        RECT 135.320 139.535 135.715 139.885 ;
        RECT 135.910 139.535 136.200 139.885 ;
        RECT 134.895 138.805 135.325 139.335 ;
        RECT 135.505 138.915 135.715 139.535 ;
        RECT 136.405 139.395 137.155 139.915 ;
        RECT 137.325 139.565 138.075 140.085 ;
        RECT 138.705 140.010 138.995 141.175 ;
        RECT 139.225 140.035 139.435 141.175 ;
        RECT 139.605 140.025 139.935 141.005 ;
        RECT 140.105 140.035 140.335 141.175 ;
        RECT 141.120 140.545 141.405 141.005 ;
        RECT 141.575 140.715 141.845 141.175 ;
        RECT 141.120 140.325 142.075 140.545 ;
        RECT 135.885 138.625 136.215 139.355 ;
        RECT 136.405 138.625 138.075 139.395 ;
        RECT 138.705 138.625 138.995 139.350 ;
        RECT 139.225 138.625 139.435 139.445 ;
        RECT 139.605 139.425 139.855 140.025 ;
        RECT 140.025 139.615 140.355 139.865 ;
        RECT 141.005 139.595 141.695 140.155 ;
        RECT 139.605 138.795 139.935 139.425 ;
        RECT 140.105 138.625 140.335 139.445 ;
        RECT 141.865 139.425 142.075 140.325 ;
        RECT 141.120 139.255 142.075 139.425 ;
        RECT 142.245 140.155 142.645 141.005 ;
        RECT 142.835 140.545 143.115 141.005 ;
        RECT 143.635 140.715 143.960 141.175 ;
        RECT 142.835 140.325 143.960 140.545 ;
        RECT 142.245 139.595 143.340 140.155 ;
        RECT 143.510 139.865 143.960 140.325 ;
        RECT 144.130 140.035 144.515 141.005 ;
        RECT 145.330 140.205 145.720 140.380 ;
        RECT 146.205 140.375 146.535 141.175 ;
        RECT 146.705 140.385 147.240 141.005 ;
        RECT 145.330 140.035 146.755 140.205 ;
        RECT 141.120 138.795 141.405 139.255 ;
        RECT 141.575 138.625 141.845 139.085 ;
        RECT 142.245 138.795 142.645 139.595 ;
        RECT 143.510 139.535 144.065 139.865 ;
        RECT 143.510 139.425 143.960 139.535 ;
        RECT 142.835 139.255 143.960 139.425 ;
        RECT 144.235 139.365 144.515 140.035 ;
        RECT 142.835 138.795 143.115 139.255 ;
        RECT 143.635 138.625 143.960 139.085 ;
        RECT 144.130 138.795 144.515 139.365 ;
        RECT 145.205 139.305 145.560 139.865 ;
        RECT 145.730 139.135 145.900 140.035 ;
        RECT 146.070 139.305 146.335 139.865 ;
        RECT 146.585 139.535 146.755 140.035 ;
        RECT 146.925 139.365 147.240 140.385 ;
        RECT 148.455 140.505 148.625 141.005 ;
        RECT 148.795 140.675 149.125 141.175 ;
        RECT 148.455 140.335 149.120 140.505 ;
        RECT 148.370 139.515 148.720 140.165 ;
        RECT 145.310 138.625 145.550 139.135 ;
        RECT 145.730 138.805 146.010 139.135 ;
        RECT 146.240 138.625 146.455 139.135 ;
        RECT 146.625 138.795 147.240 139.365 ;
        RECT 148.890 139.345 149.120 140.335 ;
        RECT 148.455 139.175 149.120 139.345 ;
        RECT 148.455 138.885 148.625 139.175 ;
        RECT 148.795 138.625 149.125 139.005 ;
        RECT 149.295 138.885 149.480 141.005 ;
        RECT 149.720 140.715 149.985 141.175 ;
        RECT 150.155 140.580 150.405 141.005 ;
        RECT 150.615 140.730 151.720 140.900 ;
        RECT 150.100 140.450 150.405 140.580 ;
        RECT 149.650 139.255 149.930 140.205 ;
        RECT 150.100 139.345 150.270 140.450 ;
        RECT 150.440 139.665 150.680 140.260 ;
        RECT 150.850 140.195 151.380 140.560 ;
        RECT 150.850 139.495 151.020 140.195 ;
        RECT 151.550 140.115 151.720 140.730 ;
        RECT 151.890 140.375 152.060 141.175 ;
        RECT 152.230 140.675 152.480 141.005 ;
        RECT 152.705 140.705 153.590 140.875 ;
        RECT 151.550 140.025 152.060 140.115 ;
        RECT 150.100 139.215 150.325 139.345 ;
        RECT 150.495 139.275 151.020 139.495 ;
        RECT 151.190 139.855 152.060 140.025 ;
        RECT 149.735 138.625 149.985 139.085 ;
        RECT 150.155 139.075 150.325 139.215 ;
        RECT 151.190 139.075 151.360 139.855 ;
        RECT 151.890 139.785 152.060 139.855 ;
        RECT 151.570 139.605 151.770 139.635 ;
        RECT 152.230 139.605 152.400 140.675 ;
        RECT 152.570 139.785 152.760 140.505 ;
        RECT 151.570 139.305 152.400 139.605 ;
        RECT 152.930 139.575 153.250 140.535 ;
        RECT 150.155 138.905 150.490 139.075 ;
        RECT 150.685 138.905 151.360 139.075 ;
        RECT 151.680 138.625 152.050 139.125 ;
        RECT 152.230 139.075 152.400 139.305 ;
        RECT 152.785 139.245 153.250 139.575 ;
        RECT 153.420 139.865 153.590 140.705 ;
        RECT 153.770 140.675 154.085 141.175 ;
        RECT 154.315 140.445 154.655 141.005 ;
        RECT 153.760 140.070 154.655 140.445 ;
        RECT 154.825 140.165 154.995 141.175 ;
        RECT 154.465 139.865 154.655 140.070 ;
        RECT 155.165 140.115 155.495 140.960 ;
        RECT 155.165 140.035 155.555 140.115 ;
        RECT 155.340 139.985 155.555 140.035 ;
        RECT 153.420 139.535 154.295 139.865 ;
        RECT 154.465 139.535 155.215 139.865 ;
        RECT 153.420 139.075 153.590 139.535 ;
        RECT 154.465 139.365 154.665 139.535 ;
        RECT 155.385 139.405 155.555 139.985 ;
        RECT 155.725 140.085 156.935 141.175 ;
        RECT 155.725 139.545 156.245 140.085 ;
        RECT 155.330 139.365 155.555 139.405 ;
        RECT 156.415 139.375 156.935 139.915 ;
        RECT 152.230 138.905 152.635 139.075 ;
        RECT 152.805 138.905 153.590 139.075 ;
        RECT 153.865 138.625 154.075 139.155 ;
        RECT 154.335 138.840 154.665 139.365 ;
        RECT 155.175 139.280 155.555 139.365 ;
        RECT 154.835 138.625 155.005 139.235 ;
        RECT 155.175 138.845 155.505 139.280 ;
        RECT 155.725 138.625 156.935 139.375 ;
        RECT 22.700 138.455 157.020 138.625 ;
        RECT 22.785 137.705 23.995 138.455 ;
        RECT 24.165 137.910 29.510 138.455 ;
        RECT 22.785 137.165 23.305 137.705 ;
        RECT 23.475 136.995 23.995 137.535 ;
        RECT 25.750 137.080 26.090 137.910 ;
        RECT 22.785 135.905 23.995 136.995 ;
        RECT 27.570 136.340 27.920 137.590 ;
        RECT 30.605 137.510 30.945 138.285 ;
        RECT 31.115 137.995 31.285 138.455 ;
        RECT 31.525 138.020 31.885 138.285 ;
        RECT 31.525 138.015 31.880 138.020 ;
        RECT 31.525 138.005 31.875 138.015 ;
        RECT 31.525 138.000 31.870 138.005 ;
        RECT 31.525 137.990 31.865 138.000 ;
        RECT 32.515 137.995 32.685 138.455 ;
        RECT 31.525 137.985 31.860 137.990 ;
        RECT 31.525 137.975 31.850 137.985 ;
        RECT 31.525 137.965 31.840 137.975 ;
        RECT 31.525 137.825 31.825 137.965 ;
        RECT 31.115 137.635 31.825 137.825 ;
        RECT 32.015 137.825 32.345 137.905 ;
        RECT 32.855 137.825 33.195 138.285 ;
        RECT 32.015 137.635 33.195 137.825 ;
        RECT 33.455 137.905 33.625 138.195 ;
        RECT 33.795 138.075 34.125 138.455 ;
        RECT 33.455 137.735 34.120 137.905 ;
        RECT 24.165 135.905 29.510 136.340 ;
        RECT 30.605 136.075 30.885 137.510 ;
        RECT 31.115 137.065 31.400 137.635 ;
        RECT 31.585 137.235 32.055 137.465 ;
        RECT 32.225 137.445 32.555 137.465 ;
        RECT 32.225 137.265 32.675 137.445 ;
        RECT 32.865 137.265 33.195 137.465 ;
        RECT 31.115 136.850 32.265 137.065 ;
        RECT 31.055 135.905 31.765 136.680 ;
        RECT 31.935 136.075 32.265 136.850 ;
        RECT 32.460 136.150 32.675 137.265 ;
        RECT 32.965 136.925 33.195 137.265 ;
        RECT 33.370 136.915 33.720 137.565 ;
        RECT 33.890 136.745 34.120 137.735 ;
        RECT 32.855 135.905 33.185 136.625 ;
        RECT 33.455 136.575 34.120 136.745 ;
        RECT 33.455 136.075 33.625 136.575 ;
        RECT 33.795 135.905 34.125 136.405 ;
        RECT 34.295 136.075 34.480 138.195 ;
        RECT 34.735 137.995 34.985 138.455 ;
        RECT 35.155 138.005 35.490 138.175 ;
        RECT 35.685 138.005 36.360 138.175 ;
        RECT 35.155 137.865 35.325 138.005 ;
        RECT 34.650 136.875 34.930 137.825 ;
        RECT 35.100 137.735 35.325 137.865 ;
        RECT 35.100 136.630 35.270 137.735 ;
        RECT 35.495 137.585 36.020 137.805 ;
        RECT 35.440 136.820 35.680 137.415 ;
        RECT 35.850 136.885 36.020 137.585 ;
        RECT 36.190 137.225 36.360 138.005 ;
        RECT 36.680 137.955 37.050 138.455 ;
        RECT 37.230 138.005 37.635 138.175 ;
        RECT 37.805 138.005 38.590 138.175 ;
        RECT 37.230 137.775 37.400 138.005 ;
        RECT 36.570 137.475 37.400 137.775 ;
        RECT 37.785 137.505 38.250 137.835 ;
        RECT 36.570 137.445 36.770 137.475 ;
        RECT 36.890 137.225 37.060 137.295 ;
        RECT 36.190 137.055 37.060 137.225 ;
        RECT 36.550 136.965 37.060 137.055 ;
        RECT 35.100 136.500 35.405 136.630 ;
        RECT 35.850 136.520 36.380 136.885 ;
        RECT 34.720 135.905 34.985 136.365 ;
        RECT 35.155 136.075 35.405 136.500 ;
        RECT 36.550 136.350 36.720 136.965 ;
        RECT 35.615 136.180 36.720 136.350 ;
        RECT 36.890 135.905 37.060 136.705 ;
        RECT 37.230 136.405 37.400 137.475 ;
        RECT 37.570 136.575 37.760 137.295 ;
        RECT 37.930 136.545 38.250 137.505 ;
        RECT 38.420 137.545 38.590 138.005 ;
        RECT 38.865 137.925 39.075 138.455 ;
        RECT 39.335 137.715 39.665 138.240 ;
        RECT 39.835 137.845 40.005 138.455 ;
        RECT 40.175 137.800 40.505 138.235 ;
        RECT 40.175 137.715 40.555 137.800 ;
        RECT 39.465 137.545 39.665 137.715 ;
        RECT 40.330 137.675 40.555 137.715 ;
        RECT 38.420 137.215 39.295 137.545 ;
        RECT 39.465 137.215 40.215 137.545 ;
        RECT 37.230 136.075 37.480 136.405 ;
        RECT 38.420 136.375 38.590 137.215 ;
        RECT 39.465 137.010 39.655 137.215 ;
        RECT 40.385 137.095 40.555 137.675 ;
        RECT 40.725 137.705 41.935 138.455 ;
        RECT 42.130 137.805 42.440 138.275 ;
        RECT 42.610 137.975 43.345 138.455 ;
        RECT 43.515 137.885 43.685 138.235 ;
        RECT 43.855 138.055 44.235 138.455 ;
        RECT 40.725 137.165 41.245 137.705 ;
        RECT 42.130 137.635 42.865 137.805 ;
        RECT 43.515 137.715 44.255 137.885 ;
        RECT 44.425 137.780 44.695 138.125 ;
        RECT 42.615 137.545 42.865 137.635 ;
        RECT 44.085 137.545 44.255 137.715 ;
        RECT 40.340 137.045 40.555 137.095 ;
        RECT 38.760 136.635 39.655 137.010 ;
        RECT 40.165 136.965 40.555 137.045 ;
        RECT 41.415 136.995 41.935 137.535 ;
        RECT 42.110 137.215 42.445 137.465 ;
        RECT 42.615 137.215 43.355 137.545 ;
        RECT 44.085 137.215 44.315 137.545 ;
        RECT 37.705 136.205 38.590 136.375 ;
        RECT 38.770 135.905 39.085 136.405 ;
        RECT 39.315 136.075 39.655 136.635 ;
        RECT 39.825 135.905 39.995 136.915 ;
        RECT 40.165 136.120 40.495 136.965 ;
        RECT 40.725 135.905 41.935 136.995 ;
        RECT 42.110 135.905 42.365 137.045 ;
        RECT 42.615 136.655 42.785 137.215 ;
        RECT 44.085 137.045 44.255 137.215 ;
        RECT 44.525 137.045 44.695 137.780 ;
        RECT 44.890 137.805 45.200 138.275 ;
        RECT 45.370 137.975 46.105 138.455 ;
        RECT 46.275 137.885 46.445 138.235 ;
        RECT 46.615 138.055 46.995 138.455 ;
        RECT 44.890 137.635 45.625 137.805 ;
        RECT 46.275 137.715 47.015 137.885 ;
        RECT 47.185 137.780 47.455 138.125 ;
        RECT 45.375 137.545 45.625 137.635 ;
        RECT 46.845 137.545 47.015 137.715 ;
        RECT 44.870 137.215 45.205 137.465 ;
        RECT 45.375 137.215 46.115 137.545 ;
        RECT 46.845 137.215 47.075 137.545 ;
        RECT 43.010 136.875 44.255 137.045 ;
        RECT 43.010 136.625 43.430 136.875 ;
        RECT 42.560 136.125 43.755 136.455 ;
        RECT 43.935 135.905 44.215 136.705 ;
        RECT 44.425 136.075 44.695 137.045 ;
        RECT 44.870 135.905 45.125 137.045 ;
        RECT 45.375 136.655 45.545 137.215 ;
        RECT 46.845 137.045 47.015 137.215 ;
        RECT 47.285 137.045 47.455 137.780 ;
        RECT 48.545 137.730 48.835 138.455 ;
        RECT 49.005 137.705 50.215 138.455 ;
        RECT 50.475 137.905 50.645 138.195 ;
        RECT 50.815 138.075 51.145 138.455 ;
        RECT 50.475 137.735 51.140 137.905 ;
        RECT 49.005 137.165 49.525 137.705 ;
        RECT 45.770 136.875 47.015 137.045 ;
        RECT 45.770 136.625 46.190 136.875 ;
        RECT 45.320 136.125 46.515 136.455 ;
        RECT 46.695 135.905 46.975 136.705 ;
        RECT 47.185 136.075 47.455 137.045 ;
        RECT 48.545 135.905 48.835 137.070 ;
        RECT 49.695 136.995 50.215 137.535 ;
        RECT 49.005 135.905 50.215 136.995 ;
        RECT 50.390 136.915 50.740 137.565 ;
        RECT 50.910 136.745 51.140 137.735 ;
        RECT 50.475 136.575 51.140 136.745 ;
        RECT 50.475 136.075 50.645 136.575 ;
        RECT 50.815 135.905 51.145 136.405 ;
        RECT 51.315 136.075 51.500 138.195 ;
        RECT 51.755 137.995 52.005 138.455 ;
        RECT 52.175 138.005 52.510 138.175 ;
        RECT 52.705 138.005 53.380 138.175 ;
        RECT 52.175 137.865 52.345 138.005 ;
        RECT 51.670 136.875 51.950 137.825 ;
        RECT 52.120 137.735 52.345 137.865 ;
        RECT 52.120 136.630 52.290 137.735 ;
        RECT 52.515 137.585 53.040 137.805 ;
        RECT 52.460 136.820 52.700 137.415 ;
        RECT 52.870 136.885 53.040 137.585 ;
        RECT 53.210 137.225 53.380 138.005 ;
        RECT 53.700 137.955 54.070 138.455 ;
        RECT 54.250 138.005 54.655 138.175 ;
        RECT 54.825 138.005 55.610 138.175 ;
        RECT 54.250 137.775 54.420 138.005 ;
        RECT 53.590 137.475 54.420 137.775 ;
        RECT 54.805 137.505 55.270 137.835 ;
        RECT 53.590 137.445 53.790 137.475 ;
        RECT 53.910 137.225 54.080 137.295 ;
        RECT 53.210 137.055 54.080 137.225 ;
        RECT 53.570 136.965 54.080 137.055 ;
        RECT 52.120 136.500 52.425 136.630 ;
        RECT 52.870 136.520 53.400 136.885 ;
        RECT 51.740 135.905 52.005 136.365 ;
        RECT 52.175 136.075 52.425 136.500 ;
        RECT 53.570 136.350 53.740 136.965 ;
        RECT 52.635 136.180 53.740 136.350 ;
        RECT 53.910 135.905 54.080 136.705 ;
        RECT 54.250 136.405 54.420 137.475 ;
        RECT 54.590 136.575 54.780 137.295 ;
        RECT 54.950 136.545 55.270 137.505 ;
        RECT 55.440 137.545 55.610 138.005 ;
        RECT 55.885 137.925 56.095 138.455 ;
        RECT 56.355 137.715 56.685 138.240 ;
        RECT 56.855 137.845 57.025 138.455 ;
        RECT 57.195 137.800 57.525 138.235 ;
        RECT 57.195 137.715 57.575 137.800 ;
        RECT 56.485 137.545 56.685 137.715 ;
        RECT 57.350 137.675 57.575 137.715 ;
        RECT 55.440 137.215 56.315 137.545 ;
        RECT 56.485 137.215 57.235 137.545 ;
        RECT 54.250 136.075 54.500 136.405 ;
        RECT 55.440 136.375 55.610 137.215 ;
        RECT 56.485 137.010 56.675 137.215 ;
        RECT 57.405 137.095 57.575 137.675 ;
        RECT 57.360 137.045 57.575 137.095 ;
        RECT 55.780 136.635 56.675 137.010 ;
        RECT 57.185 136.965 57.575 137.045 ;
        RECT 54.725 136.205 55.610 136.375 ;
        RECT 55.790 135.905 56.105 136.405 ;
        RECT 56.335 136.075 56.675 136.635 ;
        RECT 56.845 135.905 57.015 136.915 ;
        RECT 57.185 136.120 57.515 136.965 ;
        RECT 58.215 136.085 58.475 138.275 ;
        RECT 58.735 138.085 59.405 138.455 ;
        RECT 59.585 137.905 59.895 138.275 ;
        RECT 58.665 137.705 59.895 137.905 ;
        RECT 58.665 137.035 58.955 137.705 ;
        RECT 60.075 137.525 60.305 138.165 ;
        RECT 60.485 137.725 60.775 138.455 ;
        RECT 60.965 137.910 66.310 138.455 ;
        RECT 59.135 137.215 59.600 137.525 ;
        RECT 59.780 137.215 60.305 137.525 ;
        RECT 60.485 137.215 60.785 137.545 ;
        RECT 62.550 137.080 62.890 137.910 ;
        RECT 66.490 137.715 66.745 138.285 ;
        RECT 66.915 138.055 67.245 138.455 ;
        RECT 67.670 137.920 68.200 138.285 ;
        RECT 68.390 138.115 68.665 138.285 ;
        RECT 68.385 137.945 68.665 138.115 ;
        RECT 67.670 137.885 67.845 137.920 ;
        RECT 66.915 137.715 67.845 137.885 ;
        RECT 58.665 136.815 59.435 137.035 ;
        RECT 58.645 135.905 58.985 136.635 ;
        RECT 59.165 136.085 59.435 136.815 ;
        RECT 59.615 136.795 60.775 137.035 ;
        RECT 59.615 136.085 59.845 136.795 ;
        RECT 60.015 135.905 60.345 136.615 ;
        RECT 60.515 136.085 60.775 136.795 ;
        RECT 64.370 136.340 64.720 137.590 ;
        RECT 66.490 137.045 66.660 137.715 ;
        RECT 66.915 137.545 67.085 137.715 ;
        RECT 66.830 137.215 67.085 137.545 ;
        RECT 67.310 137.215 67.505 137.545 ;
        RECT 60.965 135.905 66.310 136.340 ;
        RECT 66.490 136.075 66.825 137.045 ;
        RECT 66.995 135.905 67.165 137.045 ;
        RECT 67.335 136.245 67.505 137.215 ;
        RECT 67.675 136.585 67.845 137.715 ;
        RECT 68.015 136.925 68.185 137.725 ;
        RECT 68.390 137.125 68.665 137.945 ;
        RECT 68.835 136.925 69.025 138.285 ;
        RECT 69.205 137.920 69.715 138.455 ;
        RECT 69.935 137.645 70.180 138.250 ;
        RECT 70.645 137.645 70.885 138.455 ;
        RECT 71.055 137.645 71.385 138.285 ;
        RECT 71.555 137.645 71.825 138.455 ;
        RECT 72.005 137.685 73.675 138.455 ;
        RECT 74.305 137.730 74.595 138.455 ;
        RECT 75.230 137.715 75.485 138.285 ;
        RECT 75.655 138.055 75.985 138.455 ;
        RECT 76.410 137.920 76.940 138.285 ;
        RECT 76.410 137.885 76.585 137.920 ;
        RECT 75.655 137.715 76.585 137.885 ;
        RECT 69.225 137.475 70.455 137.645 ;
        RECT 68.015 136.755 69.025 136.925 ;
        RECT 69.195 136.910 69.945 137.100 ;
        RECT 67.675 136.415 68.800 136.585 ;
        RECT 69.195 136.245 69.365 136.910 ;
        RECT 70.115 136.665 70.455 137.475 ;
        RECT 70.625 137.215 70.975 137.465 ;
        RECT 71.145 137.045 71.315 137.645 ;
        RECT 71.485 137.215 71.835 137.465 ;
        RECT 72.005 137.165 72.755 137.685 ;
        RECT 67.335 136.075 69.365 136.245 ;
        RECT 69.535 135.905 69.705 136.665 ;
        RECT 69.940 136.255 70.455 136.665 ;
        RECT 70.635 136.875 71.315 137.045 ;
        RECT 70.635 136.090 70.965 136.875 ;
        RECT 71.495 135.905 71.825 137.045 ;
        RECT 72.925 136.995 73.675 137.515 ;
        RECT 72.005 135.905 73.675 136.995 ;
        RECT 74.305 135.905 74.595 137.070 ;
        RECT 75.230 137.045 75.400 137.715 ;
        RECT 75.655 137.545 75.825 137.715 ;
        RECT 75.570 137.215 75.825 137.545 ;
        RECT 76.050 137.215 76.245 137.545 ;
        RECT 75.230 136.075 75.565 137.045 ;
        RECT 75.735 135.905 75.905 137.045 ;
        RECT 76.075 136.245 76.245 137.215 ;
        RECT 76.415 136.585 76.585 137.715 ;
        RECT 76.755 136.925 76.925 137.725 ;
        RECT 77.130 137.435 77.405 138.285 ;
        RECT 77.125 137.265 77.405 137.435 ;
        RECT 77.130 137.125 77.405 137.265 ;
        RECT 77.575 136.925 77.765 138.285 ;
        RECT 77.945 137.920 78.455 138.455 ;
        RECT 78.675 137.645 78.920 138.250 ;
        RECT 79.365 137.685 82.875 138.455 ;
        RECT 83.965 137.805 84.225 138.285 ;
        RECT 84.395 137.915 84.645 138.455 ;
        RECT 77.965 137.475 79.195 137.645 ;
        RECT 76.755 136.755 77.765 136.925 ;
        RECT 77.935 136.910 78.685 137.100 ;
        RECT 76.415 136.415 77.540 136.585 ;
        RECT 77.935 136.245 78.105 136.910 ;
        RECT 78.855 136.665 79.195 137.475 ;
        RECT 79.365 137.165 81.015 137.685 ;
        RECT 81.185 136.995 82.875 137.515 ;
        RECT 76.075 136.075 78.105 136.245 ;
        RECT 78.275 135.905 78.445 136.665 ;
        RECT 78.680 136.255 79.195 136.665 ;
        RECT 79.365 135.905 82.875 136.995 ;
        RECT 83.965 136.775 84.135 137.805 ;
        RECT 84.815 137.750 85.035 138.235 ;
        RECT 84.305 137.155 84.535 137.550 ;
        RECT 84.705 137.325 85.035 137.750 ;
        RECT 85.205 138.075 86.095 138.245 ;
        RECT 85.205 137.350 85.375 138.075 ;
        RECT 85.545 137.520 86.095 137.905 ;
        RECT 86.265 137.715 86.650 138.285 ;
        RECT 86.820 137.995 87.145 138.455 ;
        RECT 87.665 137.825 87.945 138.285 ;
        RECT 85.205 137.280 86.095 137.350 ;
        RECT 85.200 137.255 86.095 137.280 ;
        RECT 85.190 137.240 86.095 137.255 ;
        RECT 85.185 137.225 86.095 137.240 ;
        RECT 85.175 137.220 86.095 137.225 ;
        RECT 85.170 137.210 86.095 137.220 ;
        RECT 85.165 137.200 86.095 137.210 ;
        RECT 85.155 137.195 86.095 137.200 ;
        RECT 85.145 137.185 86.095 137.195 ;
        RECT 85.135 137.180 86.095 137.185 ;
        RECT 85.135 137.175 85.470 137.180 ;
        RECT 85.120 137.170 85.470 137.175 ;
        RECT 85.105 137.160 85.470 137.170 ;
        RECT 85.080 137.155 85.470 137.160 ;
        RECT 84.305 137.150 85.470 137.155 ;
        RECT 84.305 137.115 85.440 137.150 ;
        RECT 84.305 137.090 85.405 137.115 ;
        RECT 84.305 137.060 85.375 137.090 ;
        RECT 84.305 137.030 85.355 137.060 ;
        RECT 84.305 137.000 85.335 137.030 ;
        RECT 84.305 136.990 85.265 137.000 ;
        RECT 84.305 136.980 85.240 136.990 ;
        RECT 84.305 136.965 85.220 136.980 ;
        RECT 84.305 136.950 85.200 136.965 ;
        RECT 84.410 136.940 85.195 136.950 ;
        RECT 84.410 136.905 85.180 136.940 ;
        RECT 83.965 136.075 84.240 136.775 ;
        RECT 84.410 136.655 85.165 136.905 ;
        RECT 85.335 136.585 85.665 136.830 ;
        RECT 85.835 136.730 86.095 137.180 ;
        RECT 86.265 137.045 86.545 137.715 ;
        RECT 86.820 137.655 87.945 137.825 ;
        RECT 86.820 137.545 87.270 137.655 ;
        RECT 86.715 137.215 87.270 137.545 ;
        RECT 88.135 137.485 88.535 138.285 ;
        RECT 88.935 137.995 89.205 138.455 ;
        RECT 89.375 137.825 89.660 138.285 ;
        RECT 85.480 136.560 85.665 136.585 ;
        RECT 85.480 136.460 86.095 136.560 ;
        RECT 84.410 135.905 84.665 136.450 ;
        RECT 84.835 136.075 85.315 136.415 ;
        RECT 85.490 135.905 86.095 136.460 ;
        RECT 86.265 136.075 86.650 137.045 ;
        RECT 86.820 136.755 87.270 137.215 ;
        RECT 87.440 136.925 88.535 137.485 ;
        RECT 86.820 136.535 87.945 136.755 ;
        RECT 86.820 135.905 87.145 136.365 ;
        RECT 87.665 136.075 87.945 136.535 ;
        RECT 88.135 136.075 88.535 136.925 ;
        RECT 88.705 137.655 89.660 137.825 ;
        RECT 89.980 137.715 90.595 138.285 ;
        RECT 90.765 137.945 90.980 138.455 ;
        RECT 91.210 137.945 91.490 138.275 ;
        RECT 91.670 137.945 91.910 138.455 ;
        RECT 88.705 136.755 88.915 137.655 ;
        RECT 89.085 136.925 89.775 137.485 ;
        RECT 88.705 136.535 89.660 136.755 ;
        RECT 88.935 135.905 89.205 136.365 ;
        RECT 89.375 136.075 89.660 136.535 ;
        RECT 89.980 136.695 90.295 137.715 ;
        RECT 90.465 137.045 90.635 137.545 ;
        RECT 90.885 137.215 91.150 137.775 ;
        RECT 91.320 137.045 91.490 137.945 ;
        RECT 91.660 137.215 92.015 137.775 ;
        RECT 92.285 137.635 92.515 138.455 ;
        RECT 92.685 137.655 93.015 138.285 ;
        RECT 92.265 137.215 92.595 137.465 ;
        RECT 92.765 137.055 93.015 137.655 ;
        RECT 93.185 137.635 93.395 138.455 ;
        RECT 93.785 137.895 94.115 138.285 ;
        RECT 94.285 138.065 95.470 138.235 ;
        RECT 95.730 137.985 95.900 138.455 ;
        RECT 93.785 137.715 94.295 137.895 ;
        RECT 93.625 137.255 93.955 137.545 ;
        RECT 94.125 137.085 94.295 137.715 ;
        RECT 94.700 137.805 95.085 137.895 ;
        RECT 96.070 137.805 96.400 138.270 ;
        RECT 94.700 137.635 96.400 137.805 ;
        RECT 96.570 137.635 96.740 138.455 ;
        RECT 96.910 137.635 97.595 138.275 ;
        RECT 97.770 137.925 98.060 138.275 ;
        RECT 98.255 138.095 98.585 138.455 ;
        RECT 98.755 137.925 98.985 138.230 ;
        RECT 97.770 137.755 98.985 137.925 ;
        RECT 94.465 137.255 94.795 137.465 ;
        RECT 94.975 137.215 95.355 137.465 ;
        RECT 90.465 136.875 91.890 137.045 ;
        RECT 89.980 136.075 90.515 136.695 ;
        RECT 90.685 135.905 91.015 136.705 ;
        RECT 91.500 136.700 91.890 136.875 ;
        RECT 92.285 135.905 92.515 137.045 ;
        RECT 92.685 136.075 93.015 137.055 ;
        RECT 93.185 135.905 93.395 137.045 ;
        RECT 93.780 136.915 94.865 137.085 ;
        RECT 93.780 136.075 94.080 136.915 ;
        RECT 94.275 135.905 94.525 136.745 ;
        RECT 94.695 136.665 94.865 136.915 ;
        RECT 95.035 136.835 95.355 137.215 ;
        RECT 95.545 137.255 96.030 137.465 ;
        RECT 96.220 137.255 96.670 137.465 ;
        RECT 96.840 137.255 97.175 137.465 ;
        RECT 95.545 137.095 95.920 137.255 ;
        RECT 95.525 136.925 95.920 137.095 ;
        RECT 96.840 137.085 97.010 137.255 ;
        RECT 95.545 136.835 95.920 136.925 ;
        RECT 96.090 136.915 97.010 137.085 ;
        RECT 96.090 136.665 96.260 136.915 ;
        RECT 94.695 136.495 96.260 136.665 ;
        RECT 95.115 136.075 95.920 136.495 ;
        RECT 96.430 135.905 96.760 136.745 ;
        RECT 97.345 136.665 97.595 137.635 ;
        RECT 99.175 137.585 99.345 138.150 ;
        RECT 100.065 137.730 100.355 138.455 ;
        RECT 100.690 137.945 100.930 138.455 ;
        RECT 101.110 137.945 101.390 138.275 ;
        RECT 101.620 137.945 101.835 138.455 ;
        RECT 97.830 137.435 98.090 137.545 ;
        RECT 97.825 137.265 98.090 137.435 ;
        RECT 97.830 137.215 98.090 137.265 ;
        RECT 98.270 137.215 98.655 137.545 ;
        RECT 98.825 137.415 99.345 137.585 ;
        RECT 96.930 136.075 97.595 136.665 ;
        RECT 97.770 135.905 98.090 137.045 ;
        RECT 98.270 136.165 98.465 137.215 ;
        RECT 98.825 137.035 98.995 137.415 ;
        RECT 98.645 136.755 98.995 137.035 ;
        RECT 99.185 136.885 99.430 137.245 ;
        RECT 100.585 137.215 100.940 137.775 ;
        RECT 98.645 136.075 98.975 136.755 ;
        RECT 99.175 135.905 99.430 136.705 ;
        RECT 100.065 135.905 100.355 137.070 ;
        RECT 101.110 137.045 101.280 137.945 ;
        RECT 101.450 137.215 101.715 137.775 ;
        RECT 102.005 137.715 102.620 138.285 ;
        RECT 102.825 138.075 103.715 138.245 ;
        RECT 101.965 137.045 102.135 137.545 ;
        RECT 100.710 136.875 102.135 137.045 ;
        RECT 100.710 136.700 101.100 136.875 ;
        RECT 101.585 135.905 101.915 136.705 ;
        RECT 102.305 136.695 102.620 137.715 ;
        RECT 102.825 137.520 103.375 137.905 ;
        RECT 103.545 137.350 103.715 138.075 ;
        RECT 102.825 137.280 103.715 137.350 ;
        RECT 103.885 137.750 104.105 138.235 ;
        RECT 104.275 137.915 104.525 138.455 ;
        RECT 104.695 137.805 104.955 138.285 ;
        RECT 103.885 137.325 104.215 137.750 ;
        RECT 102.825 137.255 103.720 137.280 ;
        RECT 102.825 137.240 103.730 137.255 ;
        RECT 102.825 137.225 103.735 137.240 ;
        RECT 102.825 137.220 103.745 137.225 ;
        RECT 102.825 137.210 103.750 137.220 ;
        RECT 102.825 137.200 103.755 137.210 ;
        RECT 102.825 137.195 103.765 137.200 ;
        RECT 102.825 137.185 103.775 137.195 ;
        RECT 102.825 137.180 103.785 137.185 ;
        RECT 102.825 136.730 103.085 137.180 ;
        RECT 103.450 137.175 103.785 137.180 ;
        RECT 103.450 137.170 103.800 137.175 ;
        RECT 103.450 137.160 103.815 137.170 ;
        RECT 103.450 137.155 103.840 137.160 ;
        RECT 104.385 137.155 104.615 137.550 ;
        RECT 103.450 137.150 104.615 137.155 ;
        RECT 103.480 137.115 104.615 137.150 ;
        RECT 103.515 137.090 104.615 137.115 ;
        RECT 103.545 137.060 104.615 137.090 ;
        RECT 103.565 137.030 104.615 137.060 ;
        RECT 103.585 137.000 104.615 137.030 ;
        RECT 103.655 136.990 104.615 137.000 ;
        RECT 103.680 136.980 104.615 136.990 ;
        RECT 103.700 136.965 104.615 136.980 ;
        RECT 103.720 136.950 104.615 136.965 ;
        RECT 103.725 136.940 104.510 136.950 ;
        RECT 103.740 136.905 104.510 136.940 ;
        RECT 102.085 136.075 102.620 136.695 ;
        RECT 103.255 136.585 103.585 136.830 ;
        RECT 103.755 136.655 104.510 136.905 ;
        RECT 104.785 136.775 104.955 137.805 ;
        RECT 105.135 137.645 105.405 138.455 ;
        RECT 105.575 137.645 105.905 138.285 ;
        RECT 106.075 137.645 106.315 138.455 ;
        RECT 106.595 137.905 106.765 138.195 ;
        RECT 106.935 138.075 107.265 138.455 ;
        RECT 106.595 137.735 107.260 137.905 ;
        RECT 105.125 137.215 105.475 137.465 ;
        RECT 105.645 137.045 105.815 137.645 ;
        RECT 105.985 137.215 106.335 137.465 ;
        RECT 103.255 136.560 103.440 136.585 ;
        RECT 102.825 136.460 103.440 136.560 ;
        RECT 102.825 135.905 103.430 136.460 ;
        RECT 103.605 136.075 104.085 136.415 ;
        RECT 104.255 135.905 104.510 136.450 ;
        RECT 104.680 136.075 104.955 136.775 ;
        RECT 105.135 135.905 105.465 137.045 ;
        RECT 105.645 136.875 106.325 137.045 ;
        RECT 106.510 136.915 106.860 137.565 ;
        RECT 105.995 136.090 106.325 136.875 ;
        RECT 107.030 136.745 107.260 137.735 ;
        RECT 106.595 136.575 107.260 136.745 ;
        RECT 106.595 136.075 106.765 136.575 ;
        RECT 106.935 135.905 107.265 136.405 ;
        RECT 107.435 136.075 107.620 138.195 ;
        RECT 107.875 137.995 108.125 138.455 ;
        RECT 108.295 138.005 108.630 138.175 ;
        RECT 108.825 138.005 109.500 138.175 ;
        RECT 108.295 137.865 108.465 138.005 ;
        RECT 107.790 136.875 108.070 137.825 ;
        RECT 108.240 137.735 108.465 137.865 ;
        RECT 108.240 136.630 108.410 137.735 ;
        RECT 108.635 137.585 109.160 137.805 ;
        RECT 108.580 136.820 108.820 137.415 ;
        RECT 108.990 136.885 109.160 137.585 ;
        RECT 109.330 137.225 109.500 138.005 ;
        RECT 109.820 137.955 110.190 138.455 ;
        RECT 110.370 138.005 110.775 138.175 ;
        RECT 110.945 138.005 111.730 138.175 ;
        RECT 110.370 137.775 110.540 138.005 ;
        RECT 109.710 137.475 110.540 137.775 ;
        RECT 110.925 137.505 111.390 137.835 ;
        RECT 109.710 137.445 109.910 137.475 ;
        RECT 110.030 137.225 110.200 137.295 ;
        RECT 109.330 137.055 110.200 137.225 ;
        RECT 109.690 136.965 110.200 137.055 ;
        RECT 108.240 136.500 108.545 136.630 ;
        RECT 108.990 136.520 109.520 136.885 ;
        RECT 107.860 135.905 108.125 136.365 ;
        RECT 108.295 136.075 108.545 136.500 ;
        RECT 109.690 136.350 109.860 136.965 ;
        RECT 108.755 136.180 109.860 136.350 ;
        RECT 110.030 135.905 110.200 136.705 ;
        RECT 110.370 136.405 110.540 137.475 ;
        RECT 110.710 136.575 110.900 137.295 ;
        RECT 111.070 136.545 111.390 137.505 ;
        RECT 111.560 137.545 111.730 138.005 ;
        RECT 112.005 137.925 112.215 138.455 ;
        RECT 112.475 137.715 112.805 138.240 ;
        RECT 112.975 137.845 113.145 138.455 ;
        RECT 113.315 137.800 113.645 138.235 ;
        RECT 113.315 137.715 113.695 137.800 ;
        RECT 112.605 137.545 112.805 137.715 ;
        RECT 113.470 137.675 113.695 137.715 ;
        RECT 111.560 137.215 112.435 137.545 ;
        RECT 112.605 137.215 113.355 137.545 ;
        RECT 110.370 136.075 110.620 136.405 ;
        RECT 111.560 136.375 111.730 137.215 ;
        RECT 112.605 137.010 112.795 137.215 ;
        RECT 113.525 137.095 113.695 137.675 ;
        RECT 113.480 137.045 113.695 137.095 ;
        RECT 111.900 136.635 112.795 137.010 ;
        RECT 113.305 136.965 113.695 137.045 ;
        RECT 113.865 137.715 114.250 138.285 ;
        RECT 114.420 137.995 114.745 138.455 ;
        RECT 115.265 137.825 115.545 138.285 ;
        RECT 113.865 137.045 114.145 137.715 ;
        RECT 114.420 137.655 115.545 137.825 ;
        RECT 114.420 137.545 114.870 137.655 ;
        RECT 114.315 137.215 114.870 137.545 ;
        RECT 115.735 137.485 116.135 138.285 ;
        RECT 116.535 137.995 116.805 138.455 ;
        RECT 116.975 137.825 117.260 138.285 ;
        RECT 110.845 136.205 111.730 136.375 ;
        RECT 111.910 135.905 112.225 136.405 ;
        RECT 112.455 136.075 112.795 136.635 ;
        RECT 112.965 135.905 113.135 136.915 ;
        RECT 113.305 136.120 113.635 136.965 ;
        RECT 113.865 136.075 114.250 137.045 ;
        RECT 114.420 136.755 114.870 137.215 ;
        RECT 115.040 136.925 116.135 137.485 ;
        RECT 114.420 136.535 115.545 136.755 ;
        RECT 114.420 135.905 114.745 136.365 ;
        RECT 115.265 136.075 115.545 136.535 ;
        RECT 115.735 136.075 116.135 136.925 ;
        RECT 116.305 137.655 117.260 137.825 ;
        RECT 118.005 137.715 118.390 138.285 ;
        RECT 118.560 137.995 118.885 138.455 ;
        RECT 119.405 137.825 119.685 138.285 ;
        RECT 116.305 136.755 116.515 137.655 ;
        RECT 116.685 136.925 117.375 137.485 ;
        RECT 118.005 137.045 118.285 137.715 ;
        RECT 118.560 137.655 119.685 137.825 ;
        RECT 118.560 137.545 119.010 137.655 ;
        RECT 118.455 137.215 119.010 137.545 ;
        RECT 119.875 137.485 120.275 138.285 ;
        RECT 120.675 137.995 120.945 138.455 ;
        RECT 121.115 137.825 121.400 138.285 ;
        RECT 116.305 136.535 117.260 136.755 ;
        RECT 116.535 135.905 116.805 136.365 ;
        RECT 116.975 136.075 117.260 136.535 ;
        RECT 118.005 136.075 118.390 137.045 ;
        RECT 118.560 136.755 119.010 137.215 ;
        RECT 119.180 136.925 120.275 137.485 ;
        RECT 118.560 136.535 119.685 136.755 ;
        RECT 118.560 135.905 118.885 136.365 ;
        RECT 119.405 136.075 119.685 136.535 ;
        RECT 119.875 136.075 120.275 136.925 ;
        RECT 120.445 137.655 121.400 137.825 ;
        RECT 121.685 137.715 122.070 138.285 ;
        RECT 122.240 137.995 122.565 138.455 ;
        RECT 123.085 137.825 123.365 138.285 ;
        RECT 120.445 136.755 120.655 137.655 ;
        RECT 120.825 136.925 121.515 137.485 ;
        RECT 121.685 137.045 121.965 137.715 ;
        RECT 122.240 137.655 123.365 137.825 ;
        RECT 122.240 137.545 122.690 137.655 ;
        RECT 122.135 137.215 122.690 137.545 ;
        RECT 123.555 137.485 123.955 138.285 ;
        RECT 124.355 137.995 124.625 138.455 ;
        RECT 124.795 137.825 125.080 138.285 ;
        RECT 120.445 136.535 121.400 136.755 ;
        RECT 120.675 135.905 120.945 136.365 ;
        RECT 121.115 136.075 121.400 136.535 ;
        RECT 121.685 136.075 122.070 137.045 ;
        RECT 122.240 136.755 122.690 137.215 ;
        RECT 122.860 136.925 123.955 137.485 ;
        RECT 122.240 136.535 123.365 136.755 ;
        RECT 122.240 135.905 122.565 136.365 ;
        RECT 123.085 136.075 123.365 136.535 ;
        RECT 123.555 136.075 123.955 136.925 ;
        RECT 124.125 137.655 125.080 137.825 ;
        RECT 125.825 137.730 126.115 138.455 ;
        RECT 126.325 137.945 126.725 138.455 ;
        RECT 127.300 137.840 127.470 138.285 ;
        RECT 127.640 138.055 128.360 138.455 ;
        RECT 128.530 137.885 128.700 138.285 ;
        RECT 128.935 138.010 129.365 138.455 ;
        RECT 124.125 136.755 124.335 137.655 ;
        RECT 124.505 136.925 125.195 137.485 ;
        RECT 124.125 136.535 125.080 136.755 ;
        RECT 124.355 135.905 124.625 136.365 ;
        RECT 124.795 136.075 125.080 136.535 ;
        RECT 125.825 135.905 126.115 137.070 ;
        RECT 126.340 136.885 126.600 137.775 ;
        RECT 126.800 137.185 127.060 137.775 ;
        RECT 127.300 137.670 127.650 137.840 ;
        RECT 126.800 136.885 127.280 137.185 ;
        RECT 126.365 136.535 127.305 136.705 ;
        RECT 126.365 136.075 126.545 136.535 ;
        RECT 126.715 135.905 126.965 136.365 ;
        RECT 127.135 136.285 127.305 136.535 ;
        RECT 127.480 136.645 127.650 137.670 ;
        RECT 127.820 137.715 128.700 137.885 ;
        RECT 129.535 137.730 129.795 138.285 ;
        RECT 127.820 136.995 127.990 137.715 ;
        RECT 128.180 137.165 128.470 137.545 ;
        RECT 127.820 136.825 128.340 136.995 ;
        RECT 128.640 136.925 128.970 137.545 ;
        RECT 129.195 137.215 129.450 137.545 ;
        RECT 127.480 136.475 127.890 136.645 ;
        RECT 128.170 136.635 128.340 136.825 ;
        RECT 129.195 136.735 129.365 137.215 ;
        RECT 129.620 137.015 129.795 137.730 ;
        RECT 127.635 136.340 127.890 136.475 ;
        RECT 128.605 136.565 129.365 136.735 ;
        RECT 128.605 136.340 128.775 136.565 ;
        RECT 127.135 136.115 127.465 136.285 ;
        RECT 127.635 136.170 128.775 136.340 ;
        RECT 127.635 136.075 127.890 136.170 ;
        RECT 129.035 135.905 129.365 136.305 ;
        RECT 129.535 136.075 129.795 137.015 ;
        RECT 129.965 137.955 130.225 138.285 ;
        RECT 130.395 138.095 130.725 138.455 ;
        RECT 130.980 138.075 132.280 138.285 ;
        RECT 129.965 137.945 130.195 137.955 ;
        RECT 129.965 136.755 130.135 137.945 ;
        RECT 130.980 137.925 131.150 138.075 ;
        RECT 130.395 137.800 131.150 137.925 ;
        RECT 130.305 137.755 131.150 137.800 ;
        RECT 130.305 137.635 130.575 137.755 ;
        RECT 130.305 137.060 130.475 137.635 ;
        RECT 130.705 137.195 131.115 137.500 ;
        RECT 131.405 137.465 131.615 137.865 ;
        RECT 131.285 137.255 131.615 137.465 ;
        RECT 131.860 137.465 132.080 137.865 ;
        RECT 132.555 137.690 133.010 138.455 ;
        RECT 133.735 137.905 133.905 138.195 ;
        RECT 134.075 138.075 134.405 138.455 ;
        RECT 133.735 137.735 134.400 137.905 ;
        RECT 131.860 137.255 132.335 137.465 ;
        RECT 132.525 137.265 133.015 137.465 ;
        RECT 130.305 137.025 130.505 137.060 ;
        RECT 131.835 137.025 133.010 137.085 ;
        RECT 130.305 136.915 133.010 137.025 ;
        RECT 133.650 136.915 134.000 137.565 ;
        RECT 130.365 136.855 132.165 136.915 ;
        RECT 131.835 136.825 132.165 136.855 ;
        RECT 129.965 136.075 130.225 136.755 ;
        RECT 130.395 135.905 130.645 136.685 ;
        RECT 130.895 136.655 131.730 136.665 ;
        RECT 132.320 136.655 132.505 136.745 ;
        RECT 130.895 136.455 132.505 136.655 ;
        RECT 130.895 136.075 131.145 136.455 ;
        RECT 132.275 136.415 132.505 136.455 ;
        RECT 132.755 136.295 133.010 136.915 ;
        RECT 134.170 136.745 134.400 137.735 ;
        RECT 131.315 135.905 131.670 136.285 ;
        RECT 132.675 136.075 133.010 136.295 ;
        RECT 133.735 136.575 134.400 136.745 ;
        RECT 133.735 136.075 133.905 136.575 ;
        RECT 134.075 135.905 134.405 136.405 ;
        RECT 134.575 136.075 134.760 138.195 ;
        RECT 135.015 137.995 135.265 138.455 ;
        RECT 135.435 138.005 135.770 138.175 ;
        RECT 135.965 138.005 136.640 138.175 ;
        RECT 135.435 137.865 135.605 138.005 ;
        RECT 134.930 136.875 135.210 137.825 ;
        RECT 135.380 137.735 135.605 137.865 ;
        RECT 135.380 136.630 135.550 137.735 ;
        RECT 135.775 137.585 136.300 137.805 ;
        RECT 135.720 136.820 135.960 137.415 ;
        RECT 136.130 136.885 136.300 137.585 ;
        RECT 136.470 137.225 136.640 138.005 ;
        RECT 136.960 137.955 137.330 138.455 ;
        RECT 137.510 138.005 137.915 138.175 ;
        RECT 138.085 138.005 138.870 138.175 ;
        RECT 137.510 137.775 137.680 138.005 ;
        RECT 136.850 137.475 137.680 137.775 ;
        RECT 138.065 137.505 138.530 137.835 ;
        RECT 136.850 137.445 137.050 137.475 ;
        RECT 137.170 137.225 137.340 137.295 ;
        RECT 136.470 137.055 137.340 137.225 ;
        RECT 136.830 136.965 137.340 137.055 ;
        RECT 135.380 136.500 135.685 136.630 ;
        RECT 136.130 136.520 136.660 136.885 ;
        RECT 135.000 135.905 135.265 136.365 ;
        RECT 135.435 136.075 135.685 136.500 ;
        RECT 136.830 136.350 137.000 136.965 ;
        RECT 135.895 136.180 137.000 136.350 ;
        RECT 137.170 135.905 137.340 136.705 ;
        RECT 137.510 136.405 137.680 137.475 ;
        RECT 137.850 136.575 138.040 137.295 ;
        RECT 138.210 136.545 138.530 137.505 ;
        RECT 138.700 137.545 138.870 138.005 ;
        RECT 139.145 137.925 139.355 138.455 ;
        RECT 139.615 137.715 139.945 138.240 ;
        RECT 140.115 137.845 140.285 138.455 ;
        RECT 140.455 137.800 140.785 138.235 ;
        RECT 140.455 137.715 140.835 137.800 ;
        RECT 139.745 137.545 139.945 137.715 ;
        RECT 140.610 137.675 140.835 137.715 ;
        RECT 138.700 137.215 139.575 137.545 ;
        RECT 139.745 137.215 140.495 137.545 ;
        RECT 137.510 136.075 137.760 136.405 ;
        RECT 138.700 136.375 138.870 137.215 ;
        RECT 139.745 137.010 139.935 137.215 ;
        RECT 140.665 137.095 140.835 137.675 ;
        RECT 141.065 137.635 141.275 138.455 ;
        RECT 141.445 137.655 141.775 138.285 ;
        RECT 140.620 137.045 140.835 137.095 ;
        RECT 141.445 137.055 141.695 137.655 ;
        RECT 141.945 137.635 142.175 138.455 ;
        RECT 143.365 137.635 143.575 138.455 ;
        RECT 143.745 137.655 144.075 138.285 ;
        RECT 141.865 137.215 142.195 137.465 ;
        RECT 143.745 137.055 143.995 137.655 ;
        RECT 144.245 137.635 144.475 138.455 ;
        RECT 144.685 137.635 144.945 138.455 ;
        RECT 145.115 137.635 145.445 138.055 ;
        RECT 145.625 137.970 146.415 138.235 ;
        RECT 145.195 137.545 145.445 137.635 ;
        RECT 144.165 137.215 144.495 137.465 ;
        RECT 139.040 136.635 139.935 137.010 ;
        RECT 140.445 136.965 140.835 137.045 ;
        RECT 137.985 136.205 138.870 136.375 ;
        RECT 139.050 135.905 139.365 136.405 ;
        RECT 139.595 136.075 139.935 136.635 ;
        RECT 140.105 135.905 140.275 136.915 ;
        RECT 140.445 136.120 140.775 136.965 ;
        RECT 141.065 135.905 141.275 137.045 ;
        RECT 141.445 136.075 141.775 137.055 ;
        RECT 141.945 135.905 142.175 137.045 ;
        RECT 143.365 135.905 143.575 137.045 ;
        RECT 143.745 136.075 144.075 137.055 ;
        RECT 144.245 135.905 144.475 137.045 ;
        RECT 144.685 136.585 145.025 137.465 ;
        RECT 145.195 137.295 145.990 137.545 ;
        RECT 144.685 135.905 144.945 136.415 ;
        RECT 145.195 136.075 145.365 137.295 ;
        RECT 146.160 137.115 146.415 137.970 ;
        RECT 146.585 137.815 146.785 138.235 ;
        RECT 146.975 137.995 147.305 138.455 ;
        RECT 146.585 137.295 146.995 137.815 ;
        RECT 147.475 137.805 147.735 138.285 ;
        RECT 147.165 137.115 147.395 137.545 ;
        RECT 145.605 136.945 147.395 137.115 ;
        RECT 145.605 136.580 145.855 136.945 ;
        RECT 146.025 136.585 146.355 136.775 ;
        RECT 146.575 136.650 147.290 136.945 ;
        RECT 147.565 136.775 147.735 137.805 ;
        RECT 147.905 137.705 149.115 138.455 ;
        RECT 149.375 137.905 149.545 138.285 ;
        RECT 149.725 138.075 150.055 138.455 ;
        RECT 149.375 137.735 150.040 137.905 ;
        RECT 150.235 137.780 150.495 138.285 ;
        RECT 147.905 137.165 148.425 137.705 ;
        RECT 148.595 136.995 149.115 137.535 ;
        RECT 149.305 137.185 149.635 137.555 ;
        RECT 149.870 137.480 150.040 137.735 ;
        RECT 149.870 137.150 150.155 137.480 ;
        RECT 149.870 137.005 150.040 137.150 ;
        RECT 146.025 136.410 146.220 136.585 ;
        RECT 145.605 135.905 146.220 136.410 ;
        RECT 146.390 136.075 146.865 136.415 ;
        RECT 147.035 135.905 147.250 136.450 ;
        RECT 147.460 136.075 147.735 136.775 ;
        RECT 147.905 135.905 149.115 136.995 ;
        RECT 149.375 136.835 150.040 137.005 ;
        RECT 150.325 136.980 150.495 137.780 ;
        RECT 151.585 137.730 151.875 138.455 ;
        RECT 152.045 137.685 155.555 138.455 ;
        RECT 155.725 137.705 156.935 138.455 ;
        RECT 152.045 137.165 153.695 137.685 ;
        RECT 149.375 136.075 149.545 136.835 ;
        RECT 149.725 135.905 150.055 136.665 ;
        RECT 150.225 136.075 150.495 136.980 ;
        RECT 151.585 135.905 151.875 137.070 ;
        RECT 153.865 136.995 155.555 137.515 ;
        RECT 152.045 135.905 155.555 136.995 ;
        RECT 155.725 136.995 156.245 137.535 ;
        RECT 156.415 137.165 156.935 137.705 ;
        RECT 155.725 135.905 156.935 136.995 ;
        RECT 22.700 135.735 157.020 135.905 ;
        RECT 22.785 134.645 23.995 135.735 ;
        RECT 24.165 134.645 26.755 135.735 ;
        RECT 22.785 133.935 23.305 134.475 ;
        RECT 23.475 134.105 23.995 134.645 ;
        RECT 24.165 133.955 25.375 134.475 ;
        RECT 25.545 134.125 26.755 134.645 ;
        RECT 26.960 134.945 27.495 135.565 ;
        RECT 22.785 133.185 23.995 133.935 ;
        RECT 24.165 133.185 26.755 133.955 ;
        RECT 26.960 133.925 27.275 134.945 ;
        RECT 27.665 134.935 27.995 135.735 ;
        RECT 28.480 134.765 28.870 134.940 ;
        RECT 27.445 134.595 28.870 134.765 ;
        RECT 29.225 134.865 29.500 135.565 ;
        RECT 29.670 135.190 29.925 135.735 ;
        RECT 30.095 135.225 30.575 135.565 ;
        RECT 30.750 135.180 31.355 135.735 ;
        RECT 30.740 135.080 31.355 135.180 ;
        RECT 30.740 135.055 30.925 135.080 ;
        RECT 27.445 134.095 27.615 134.595 ;
        RECT 26.960 133.355 27.575 133.925 ;
        RECT 27.865 133.865 28.130 134.425 ;
        RECT 28.300 133.695 28.470 134.595 ;
        RECT 28.640 133.865 28.995 134.425 ;
        RECT 29.225 133.835 29.395 134.865 ;
        RECT 29.670 134.735 30.425 134.985 ;
        RECT 30.595 134.810 30.925 135.055 ;
        RECT 29.670 134.700 30.440 134.735 ;
        RECT 29.670 134.690 30.455 134.700 ;
        RECT 29.565 134.675 30.460 134.690 ;
        RECT 29.565 134.660 30.480 134.675 ;
        RECT 29.565 134.650 30.500 134.660 ;
        RECT 29.565 134.640 30.525 134.650 ;
        RECT 29.565 134.610 30.595 134.640 ;
        RECT 29.565 134.580 30.615 134.610 ;
        RECT 29.565 134.550 30.635 134.580 ;
        RECT 29.565 134.525 30.665 134.550 ;
        RECT 29.565 134.490 30.700 134.525 ;
        RECT 29.565 134.485 30.730 134.490 ;
        RECT 29.565 134.090 29.795 134.485 ;
        RECT 30.340 134.480 30.730 134.485 ;
        RECT 30.365 134.470 30.730 134.480 ;
        RECT 30.380 134.465 30.730 134.470 ;
        RECT 30.395 134.460 30.730 134.465 ;
        RECT 31.095 134.460 31.355 134.910 ;
        RECT 31.525 134.595 31.805 135.735 ;
        RECT 31.975 134.585 32.305 135.565 ;
        RECT 32.475 134.595 32.735 135.735 ;
        RECT 32.905 134.645 35.495 135.735 ;
        RECT 30.395 134.455 31.355 134.460 ;
        RECT 30.405 134.445 31.355 134.455 ;
        RECT 30.415 134.440 31.355 134.445 ;
        RECT 30.425 134.430 31.355 134.440 ;
        RECT 30.430 134.420 31.355 134.430 ;
        RECT 30.435 134.415 31.355 134.420 ;
        RECT 30.445 134.400 31.355 134.415 ;
        RECT 30.450 134.385 31.355 134.400 ;
        RECT 30.460 134.360 31.355 134.385 ;
        RECT 29.965 133.890 30.295 134.315 ;
        RECT 27.745 133.185 27.960 133.695 ;
        RECT 28.190 133.365 28.470 133.695 ;
        RECT 28.650 133.185 28.890 133.695 ;
        RECT 29.225 133.355 29.485 133.835 ;
        RECT 29.655 133.185 29.905 133.725 ;
        RECT 30.075 133.405 30.295 133.890 ;
        RECT 30.465 134.290 31.355 134.360 ;
        RECT 30.465 133.565 30.635 134.290 ;
        RECT 31.535 134.155 31.870 134.425 ;
        RECT 30.805 133.735 31.355 134.120 ;
        RECT 32.040 133.985 32.210 134.585 ;
        RECT 32.380 134.175 32.715 134.425 ;
        RECT 30.465 133.395 31.355 133.565 ;
        RECT 31.525 133.185 31.835 133.985 ;
        RECT 32.040 133.355 32.735 133.985 ;
        RECT 32.905 133.955 34.115 134.475 ;
        RECT 34.285 134.125 35.495 134.645 ;
        RECT 35.665 134.570 35.955 135.735 ;
        RECT 36.125 134.595 36.510 135.565 ;
        RECT 36.680 135.275 37.005 135.735 ;
        RECT 37.525 135.105 37.805 135.565 ;
        RECT 36.680 134.885 37.805 135.105 ;
        RECT 32.905 133.185 35.495 133.955 ;
        RECT 36.125 133.925 36.405 134.595 ;
        RECT 36.680 134.425 37.130 134.885 ;
        RECT 37.995 134.715 38.395 135.565 ;
        RECT 38.795 135.275 39.065 135.735 ;
        RECT 39.235 135.105 39.520 135.565 ;
        RECT 36.575 134.095 37.130 134.425 ;
        RECT 37.300 134.155 38.395 134.715 ;
        RECT 36.680 133.985 37.130 134.095 ;
        RECT 35.665 133.185 35.955 133.910 ;
        RECT 36.125 133.355 36.510 133.925 ;
        RECT 36.680 133.815 37.805 133.985 ;
        RECT 36.680 133.185 37.005 133.645 ;
        RECT 37.525 133.355 37.805 133.815 ;
        RECT 37.995 133.355 38.395 134.155 ;
        RECT 38.565 134.885 39.520 135.105 ;
        RECT 38.565 133.985 38.775 134.885 ;
        RECT 38.945 134.155 39.635 134.715 ;
        RECT 39.805 134.645 41.015 135.735 ;
        RECT 38.565 133.815 39.520 133.985 ;
        RECT 38.795 133.185 39.065 133.645 ;
        RECT 39.235 133.355 39.520 133.815 ;
        RECT 39.805 133.935 40.325 134.475 ;
        RECT 40.495 134.105 41.015 134.645 ;
        RECT 41.185 134.595 41.475 135.735 ;
        RECT 41.645 135.015 42.095 135.565 ;
        RECT 42.285 135.015 42.615 135.735 ;
        RECT 39.805 133.185 41.015 133.935 ;
        RECT 41.185 133.185 41.475 133.985 ;
        RECT 41.645 133.645 41.895 135.015 ;
        RECT 42.825 134.845 43.125 135.395 ;
        RECT 43.295 135.065 43.575 135.735 ;
        RECT 42.185 134.675 43.125 134.845 ;
        RECT 42.185 134.425 42.355 134.675 ;
        RECT 43.460 134.425 43.775 134.865 ;
        RECT 42.065 134.095 42.355 134.425 ;
        RECT 42.525 134.175 42.855 134.425 ;
        RECT 43.085 134.175 43.775 134.425 ;
        RECT 43.945 134.595 44.330 135.565 ;
        RECT 44.500 135.275 44.825 135.735 ;
        RECT 45.345 135.105 45.625 135.565 ;
        RECT 44.500 134.885 45.625 135.105 ;
        RECT 42.185 134.005 42.355 134.095 ;
        RECT 42.185 133.815 43.575 134.005 ;
        RECT 41.645 133.355 42.195 133.645 ;
        RECT 42.365 133.185 42.615 133.645 ;
        RECT 43.245 133.455 43.575 133.815 ;
        RECT 43.945 133.925 44.225 134.595 ;
        RECT 44.500 134.425 44.950 134.885 ;
        RECT 45.815 134.715 46.215 135.565 ;
        RECT 46.615 135.275 46.885 135.735 ;
        RECT 47.055 135.105 47.340 135.565 ;
        RECT 44.395 134.095 44.950 134.425 ;
        RECT 45.120 134.155 46.215 134.715 ;
        RECT 44.500 133.985 44.950 134.095 ;
        RECT 43.945 133.355 44.330 133.925 ;
        RECT 44.500 133.815 45.625 133.985 ;
        RECT 44.500 133.185 44.825 133.645 ;
        RECT 45.345 133.355 45.625 133.815 ;
        RECT 45.815 133.355 46.215 134.155 ;
        RECT 46.385 134.885 47.340 135.105 ;
        RECT 46.385 133.985 46.595 134.885 ;
        RECT 46.765 134.155 47.455 134.715 ;
        RECT 47.625 134.645 51.135 135.735 ;
        RECT 51.305 134.645 52.515 135.735 ;
        RECT 46.385 133.815 47.340 133.985 ;
        RECT 46.615 133.185 46.885 133.645 ;
        RECT 47.055 133.355 47.340 133.815 ;
        RECT 47.625 133.955 49.275 134.475 ;
        RECT 49.445 134.125 51.135 134.645 ;
        RECT 47.625 133.185 51.135 133.955 ;
        RECT 51.305 133.935 51.825 134.475 ;
        RECT 51.995 134.105 52.515 134.645 ;
        RECT 52.685 134.595 53.070 135.565 ;
        RECT 53.240 135.275 53.565 135.735 ;
        RECT 54.085 135.105 54.365 135.565 ;
        RECT 53.240 134.885 54.365 135.105 ;
        RECT 51.305 133.185 52.515 133.935 ;
        RECT 52.685 133.925 52.965 134.595 ;
        RECT 53.240 134.425 53.690 134.885 ;
        RECT 54.555 134.715 54.955 135.565 ;
        RECT 55.355 135.275 55.625 135.735 ;
        RECT 55.795 135.105 56.080 135.565 ;
        RECT 53.135 134.095 53.690 134.425 ;
        RECT 53.860 134.155 54.955 134.715 ;
        RECT 53.240 133.985 53.690 134.095 ;
        RECT 52.685 133.355 53.070 133.925 ;
        RECT 53.240 133.815 54.365 133.985 ;
        RECT 53.240 133.185 53.565 133.645 ;
        RECT 54.085 133.355 54.365 133.815 ;
        RECT 54.555 133.355 54.955 134.155 ;
        RECT 55.125 134.885 56.080 135.105 ;
        RECT 55.125 133.985 55.335 134.885 ;
        RECT 55.505 134.155 56.195 134.715 ;
        RECT 56.365 134.645 59.875 135.735 ;
        RECT 60.045 134.645 61.255 135.735 ;
        RECT 55.125 133.815 56.080 133.985 ;
        RECT 55.355 133.185 55.625 133.645 ;
        RECT 55.795 133.355 56.080 133.815 ;
        RECT 56.365 133.955 58.015 134.475 ;
        RECT 58.185 134.125 59.875 134.645 ;
        RECT 56.365 133.185 59.875 133.955 ;
        RECT 60.045 133.935 60.565 134.475 ;
        RECT 60.735 134.105 61.255 134.645 ;
        RECT 61.425 134.570 61.715 135.735 ;
        RECT 61.885 135.300 67.230 135.735 ;
        RECT 60.045 133.185 61.255 133.935 ;
        RECT 61.425 133.185 61.715 133.910 ;
        RECT 63.470 133.730 63.810 134.560 ;
        RECT 65.290 134.050 65.640 135.300 ;
        RECT 67.405 134.645 69.995 135.735 ;
        RECT 67.405 133.955 68.615 134.475 ;
        RECT 68.785 134.125 69.995 134.645 ;
        RECT 70.715 134.805 70.885 135.565 ;
        RECT 71.065 134.975 71.395 135.735 ;
        RECT 70.715 134.635 71.380 134.805 ;
        RECT 71.565 134.660 71.835 135.565 ;
        RECT 72.095 135.065 72.265 135.565 ;
        RECT 72.435 135.235 72.765 135.735 ;
        RECT 72.095 134.895 72.760 135.065 ;
        RECT 71.210 134.490 71.380 134.635 ;
        RECT 70.645 134.085 70.975 134.455 ;
        RECT 71.210 134.160 71.495 134.490 ;
        RECT 61.885 133.185 67.230 133.730 ;
        RECT 67.405 133.185 69.995 133.955 ;
        RECT 71.210 133.905 71.380 134.160 ;
        RECT 70.715 133.735 71.380 133.905 ;
        RECT 71.665 133.860 71.835 134.660 ;
        RECT 72.010 134.075 72.360 134.725 ;
        RECT 72.530 133.905 72.760 134.895 ;
        RECT 70.715 133.355 70.885 133.735 ;
        RECT 71.065 133.185 71.395 133.565 ;
        RECT 71.575 133.355 71.835 133.860 ;
        RECT 72.095 133.735 72.760 133.905 ;
        RECT 72.095 133.445 72.265 133.735 ;
        RECT 72.435 133.185 72.765 133.565 ;
        RECT 72.935 133.445 73.120 135.565 ;
        RECT 73.360 135.275 73.625 135.735 ;
        RECT 73.795 135.140 74.045 135.565 ;
        RECT 74.255 135.290 75.360 135.460 ;
        RECT 73.740 135.010 74.045 135.140 ;
        RECT 73.290 133.815 73.570 134.765 ;
        RECT 73.740 133.905 73.910 135.010 ;
        RECT 74.080 134.225 74.320 134.820 ;
        RECT 74.490 134.755 75.020 135.120 ;
        RECT 74.490 134.055 74.660 134.755 ;
        RECT 75.190 134.675 75.360 135.290 ;
        RECT 75.530 134.935 75.700 135.735 ;
        RECT 75.870 135.235 76.120 135.565 ;
        RECT 76.345 135.265 77.230 135.435 ;
        RECT 75.190 134.585 75.700 134.675 ;
        RECT 73.740 133.775 73.965 133.905 ;
        RECT 74.135 133.835 74.660 134.055 ;
        RECT 74.830 134.415 75.700 134.585 ;
        RECT 73.375 133.185 73.625 133.645 ;
        RECT 73.795 133.635 73.965 133.775 ;
        RECT 74.830 133.635 75.000 134.415 ;
        RECT 75.530 134.345 75.700 134.415 ;
        RECT 75.210 134.165 75.410 134.195 ;
        RECT 75.870 134.165 76.040 135.235 ;
        RECT 76.210 134.345 76.400 135.065 ;
        RECT 75.210 133.865 76.040 134.165 ;
        RECT 76.570 134.135 76.890 135.095 ;
        RECT 73.795 133.465 74.130 133.635 ;
        RECT 74.325 133.465 75.000 133.635 ;
        RECT 75.320 133.185 75.690 133.685 ;
        RECT 75.870 133.635 76.040 133.865 ;
        RECT 76.425 133.805 76.890 134.135 ;
        RECT 77.060 134.425 77.230 135.265 ;
        RECT 77.410 135.235 77.725 135.735 ;
        RECT 77.955 135.005 78.295 135.565 ;
        RECT 77.400 134.630 78.295 135.005 ;
        RECT 78.465 134.725 78.635 135.735 ;
        RECT 78.105 134.425 78.295 134.630 ;
        RECT 78.805 134.675 79.135 135.520 ;
        RECT 79.455 135.065 79.625 135.565 ;
        RECT 79.795 135.235 80.125 135.735 ;
        RECT 79.455 134.895 80.120 135.065 ;
        RECT 78.805 134.595 79.195 134.675 ;
        RECT 78.980 134.545 79.195 134.595 ;
        RECT 77.060 134.095 77.935 134.425 ;
        RECT 78.105 134.095 78.855 134.425 ;
        RECT 77.060 133.635 77.230 134.095 ;
        RECT 78.105 133.925 78.305 134.095 ;
        RECT 79.025 133.965 79.195 134.545 ;
        RECT 79.370 134.075 79.720 134.725 ;
        RECT 78.970 133.925 79.195 133.965 ;
        RECT 75.870 133.465 76.275 133.635 ;
        RECT 76.445 133.465 77.230 133.635 ;
        RECT 77.505 133.185 77.715 133.715 ;
        RECT 77.975 133.400 78.305 133.925 ;
        RECT 78.815 133.840 79.195 133.925 ;
        RECT 79.890 133.905 80.120 134.895 ;
        RECT 78.475 133.185 78.645 133.795 ;
        RECT 78.815 133.405 79.145 133.840 ;
        RECT 79.455 133.735 80.120 133.905 ;
        RECT 79.455 133.445 79.625 133.735 ;
        RECT 79.795 133.185 80.125 133.565 ;
        RECT 80.295 133.445 80.480 135.565 ;
        RECT 80.720 135.275 80.985 135.735 ;
        RECT 81.155 135.140 81.405 135.565 ;
        RECT 81.615 135.290 82.720 135.460 ;
        RECT 81.100 135.010 81.405 135.140 ;
        RECT 80.650 133.815 80.930 134.765 ;
        RECT 81.100 133.905 81.270 135.010 ;
        RECT 81.440 134.225 81.680 134.820 ;
        RECT 81.850 134.755 82.380 135.120 ;
        RECT 81.850 134.055 82.020 134.755 ;
        RECT 82.550 134.675 82.720 135.290 ;
        RECT 82.890 134.935 83.060 135.735 ;
        RECT 83.230 135.235 83.480 135.565 ;
        RECT 83.705 135.265 84.590 135.435 ;
        RECT 82.550 134.585 83.060 134.675 ;
        RECT 81.100 133.775 81.325 133.905 ;
        RECT 81.495 133.835 82.020 134.055 ;
        RECT 82.190 134.415 83.060 134.585 ;
        RECT 80.735 133.185 80.985 133.645 ;
        RECT 81.155 133.635 81.325 133.775 ;
        RECT 82.190 133.635 82.360 134.415 ;
        RECT 82.890 134.345 83.060 134.415 ;
        RECT 82.570 134.165 82.770 134.195 ;
        RECT 83.230 134.165 83.400 135.235 ;
        RECT 83.570 134.345 83.760 135.065 ;
        RECT 82.570 133.865 83.400 134.165 ;
        RECT 83.930 134.135 84.250 135.095 ;
        RECT 81.155 133.465 81.490 133.635 ;
        RECT 81.685 133.465 82.360 133.635 ;
        RECT 82.680 133.185 83.050 133.685 ;
        RECT 83.230 133.635 83.400 133.865 ;
        RECT 83.785 133.805 84.250 134.135 ;
        RECT 84.420 134.425 84.590 135.265 ;
        RECT 84.770 135.235 85.085 135.735 ;
        RECT 85.315 135.005 85.655 135.565 ;
        RECT 84.760 134.630 85.655 135.005 ;
        RECT 85.825 134.725 85.995 135.735 ;
        RECT 85.465 134.425 85.655 134.630 ;
        RECT 86.165 134.675 86.495 135.520 ;
        RECT 86.165 134.595 86.555 134.675 ;
        RECT 86.340 134.545 86.555 134.595 ;
        RECT 87.185 134.570 87.475 135.735 ;
        RECT 87.645 134.865 87.920 135.565 ;
        RECT 88.090 135.190 88.345 135.735 ;
        RECT 88.515 135.225 88.995 135.565 ;
        RECT 89.170 135.180 89.775 135.735 ;
        RECT 89.160 135.080 89.775 135.180 ;
        RECT 89.160 135.055 89.345 135.080 ;
        RECT 84.420 134.095 85.295 134.425 ;
        RECT 85.465 134.095 86.215 134.425 ;
        RECT 84.420 133.635 84.590 134.095 ;
        RECT 85.465 133.925 85.665 134.095 ;
        RECT 86.385 133.965 86.555 134.545 ;
        RECT 86.330 133.925 86.555 133.965 ;
        RECT 83.230 133.465 83.635 133.635 ;
        RECT 83.805 133.465 84.590 133.635 ;
        RECT 84.865 133.185 85.075 133.715 ;
        RECT 85.335 133.400 85.665 133.925 ;
        RECT 86.175 133.840 86.555 133.925 ;
        RECT 85.835 133.185 86.005 133.795 ;
        RECT 86.175 133.405 86.505 133.840 ;
        RECT 87.185 133.185 87.475 133.910 ;
        RECT 87.645 133.835 87.815 134.865 ;
        RECT 88.090 134.735 88.845 134.985 ;
        RECT 89.015 134.810 89.345 135.055 ;
        RECT 88.090 134.700 88.860 134.735 ;
        RECT 88.090 134.690 88.875 134.700 ;
        RECT 87.985 134.675 88.880 134.690 ;
        RECT 87.985 134.660 88.900 134.675 ;
        RECT 87.985 134.650 88.920 134.660 ;
        RECT 87.985 134.640 88.945 134.650 ;
        RECT 87.985 134.610 89.015 134.640 ;
        RECT 87.985 134.580 89.035 134.610 ;
        RECT 87.985 134.550 89.055 134.580 ;
        RECT 87.985 134.525 89.085 134.550 ;
        RECT 87.985 134.490 89.120 134.525 ;
        RECT 87.985 134.485 89.150 134.490 ;
        RECT 87.985 134.090 88.215 134.485 ;
        RECT 88.760 134.480 89.150 134.485 ;
        RECT 88.785 134.470 89.150 134.480 ;
        RECT 88.800 134.465 89.150 134.470 ;
        RECT 88.815 134.460 89.150 134.465 ;
        RECT 89.515 134.460 89.775 134.910 ;
        RECT 90.445 134.595 90.675 135.735 ;
        RECT 90.845 134.585 91.175 135.565 ;
        RECT 91.345 134.595 91.555 135.735 ;
        RECT 91.785 134.645 95.295 135.735 ;
        RECT 88.815 134.455 89.775 134.460 ;
        RECT 88.825 134.445 89.775 134.455 ;
        RECT 88.835 134.440 89.775 134.445 ;
        RECT 88.845 134.430 89.775 134.440 ;
        RECT 88.850 134.420 89.775 134.430 ;
        RECT 88.855 134.415 89.775 134.420 ;
        RECT 88.865 134.400 89.775 134.415 ;
        RECT 88.870 134.385 89.775 134.400 ;
        RECT 88.880 134.360 89.775 134.385 ;
        RECT 88.385 133.890 88.715 134.315 ;
        RECT 87.645 133.355 87.905 133.835 ;
        RECT 88.075 133.185 88.325 133.725 ;
        RECT 88.495 133.405 88.715 133.890 ;
        RECT 88.885 134.290 89.775 134.360 ;
        RECT 88.885 133.565 89.055 134.290 ;
        RECT 90.425 134.175 90.755 134.425 ;
        RECT 89.225 133.735 89.775 134.120 ;
        RECT 88.885 133.395 89.775 133.565 ;
        RECT 90.445 133.185 90.675 134.005 ;
        RECT 90.925 133.985 91.175 134.585 ;
        RECT 90.845 133.355 91.175 133.985 ;
        RECT 91.345 133.185 91.555 134.005 ;
        RECT 91.785 133.955 93.435 134.475 ;
        RECT 93.605 134.125 95.295 134.645 ;
        RECT 95.965 134.595 96.195 135.735 ;
        RECT 96.365 134.585 96.695 135.565 ;
        RECT 96.865 134.595 97.075 135.735 ;
        RECT 97.315 134.765 97.645 135.550 ;
        RECT 97.315 134.595 97.995 134.765 ;
        RECT 98.175 134.595 98.505 135.735 ;
        RECT 98.685 135.300 104.030 135.735 ;
        RECT 95.945 134.175 96.275 134.425 ;
        RECT 91.785 133.185 95.295 133.955 ;
        RECT 95.965 133.185 96.195 134.005 ;
        RECT 96.445 133.985 96.695 134.585 ;
        RECT 97.305 134.175 97.655 134.425 ;
        RECT 96.365 133.355 96.695 133.985 ;
        RECT 96.865 133.185 97.075 134.005 ;
        RECT 97.825 133.995 97.995 134.595 ;
        RECT 98.165 134.175 98.515 134.425 ;
        RECT 97.325 133.185 97.565 133.995 ;
        RECT 97.735 133.355 98.065 133.995 ;
        RECT 98.235 133.185 98.505 133.995 ;
        RECT 100.270 133.730 100.610 134.560 ;
        RECT 102.090 134.050 102.440 135.300 ;
        RECT 104.205 134.645 106.795 135.735 ;
        RECT 104.205 133.955 105.415 134.475 ;
        RECT 105.585 134.125 106.795 134.645 ;
        RECT 107.425 134.885 107.685 135.565 ;
        RECT 107.855 134.955 108.105 135.735 ;
        RECT 108.355 135.185 108.605 135.565 ;
        RECT 108.775 135.355 109.130 135.735 ;
        RECT 110.135 135.345 110.470 135.565 ;
        RECT 109.735 135.185 109.965 135.225 ;
        RECT 108.355 134.985 109.965 135.185 ;
        RECT 108.355 134.975 109.190 134.985 ;
        RECT 109.780 134.895 109.965 134.985 ;
        RECT 98.685 133.185 104.030 133.730 ;
        RECT 104.205 133.185 106.795 133.955 ;
        RECT 107.425 133.685 107.595 134.885 ;
        RECT 109.295 134.785 109.625 134.815 ;
        RECT 107.825 134.725 109.625 134.785 ;
        RECT 110.215 134.725 110.470 135.345 ;
        RECT 107.765 134.615 110.470 134.725 ;
        RECT 110.645 134.645 112.315 135.735 ;
        RECT 107.765 134.580 107.965 134.615 ;
        RECT 107.765 134.005 107.935 134.580 ;
        RECT 109.295 134.555 110.470 134.615 ;
        RECT 108.165 134.140 108.575 134.445 ;
        RECT 108.745 134.175 109.075 134.385 ;
        RECT 107.765 133.885 108.035 134.005 ;
        RECT 107.765 133.840 108.610 133.885 ;
        RECT 107.855 133.715 108.610 133.840 ;
        RECT 108.865 133.775 109.075 134.175 ;
        RECT 109.320 134.175 109.795 134.385 ;
        RECT 109.985 134.175 110.475 134.375 ;
        RECT 109.320 133.775 109.540 134.175 ;
        RECT 110.645 133.955 111.395 134.475 ;
        RECT 111.565 134.125 112.315 134.645 ;
        RECT 112.945 134.570 113.235 135.735 ;
        RECT 113.405 134.645 115.995 135.735 ;
        RECT 116.255 135.065 116.425 135.565 ;
        RECT 116.595 135.235 116.925 135.735 ;
        RECT 116.255 134.895 116.920 135.065 ;
        RECT 113.405 133.955 114.615 134.475 ;
        RECT 114.785 134.125 115.995 134.645 ;
        RECT 116.170 134.075 116.520 134.725 ;
        RECT 107.425 133.355 107.685 133.685 ;
        RECT 108.440 133.565 108.610 133.715 ;
        RECT 107.855 133.185 108.185 133.545 ;
        RECT 108.440 133.355 109.740 133.565 ;
        RECT 110.015 133.185 110.470 133.950 ;
        RECT 110.645 133.185 112.315 133.955 ;
        RECT 112.945 133.185 113.235 133.910 ;
        RECT 113.405 133.185 115.995 133.955 ;
        RECT 116.690 133.905 116.920 134.895 ;
        RECT 116.255 133.735 116.920 133.905 ;
        RECT 116.255 133.445 116.425 133.735 ;
        RECT 116.595 133.185 116.925 133.565 ;
        RECT 117.095 133.445 117.280 135.565 ;
        RECT 117.520 135.275 117.785 135.735 ;
        RECT 117.955 135.140 118.205 135.565 ;
        RECT 118.415 135.290 119.520 135.460 ;
        RECT 117.900 135.010 118.205 135.140 ;
        RECT 117.450 133.815 117.730 134.765 ;
        RECT 117.900 133.905 118.070 135.010 ;
        RECT 118.240 134.225 118.480 134.820 ;
        RECT 118.650 134.755 119.180 135.120 ;
        RECT 118.650 134.055 118.820 134.755 ;
        RECT 119.350 134.675 119.520 135.290 ;
        RECT 119.690 134.935 119.860 135.735 ;
        RECT 120.030 135.235 120.280 135.565 ;
        RECT 120.505 135.265 121.390 135.435 ;
        RECT 119.350 134.585 119.860 134.675 ;
        RECT 117.900 133.775 118.125 133.905 ;
        RECT 118.295 133.835 118.820 134.055 ;
        RECT 118.990 134.415 119.860 134.585 ;
        RECT 117.535 133.185 117.785 133.645 ;
        RECT 117.955 133.635 118.125 133.775 ;
        RECT 118.990 133.635 119.160 134.415 ;
        RECT 119.690 134.345 119.860 134.415 ;
        RECT 119.370 134.165 119.570 134.195 ;
        RECT 120.030 134.165 120.200 135.235 ;
        RECT 120.370 134.345 120.560 135.065 ;
        RECT 119.370 133.865 120.200 134.165 ;
        RECT 120.730 134.135 121.050 135.095 ;
        RECT 117.955 133.465 118.290 133.635 ;
        RECT 118.485 133.465 119.160 133.635 ;
        RECT 119.480 133.185 119.850 133.685 ;
        RECT 120.030 133.635 120.200 133.865 ;
        RECT 120.585 133.805 121.050 134.135 ;
        RECT 121.220 134.425 121.390 135.265 ;
        RECT 121.570 135.235 121.885 135.735 ;
        RECT 122.115 135.005 122.455 135.565 ;
        RECT 121.560 134.630 122.455 135.005 ;
        RECT 122.625 134.725 122.795 135.735 ;
        RECT 122.265 134.425 122.455 134.630 ;
        RECT 122.965 134.675 123.295 135.520 ;
        RECT 122.965 134.595 123.355 134.675 ;
        RECT 123.565 134.595 123.795 135.735 ;
        RECT 123.140 134.545 123.355 134.595 ;
        RECT 123.965 134.585 124.295 135.565 ;
        RECT 124.465 134.595 124.675 135.735 ;
        RECT 125.365 134.595 125.645 135.735 ;
        RECT 125.815 134.585 126.145 135.565 ;
        RECT 126.315 134.595 126.575 135.735 ;
        RECT 126.900 134.725 127.200 135.565 ;
        RECT 127.395 134.895 127.645 135.735 ;
        RECT 128.235 135.145 129.040 135.565 ;
        RECT 127.815 134.975 129.380 135.145 ;
        RECT 127.815 134.725 127.985 134.975 ;
        RECT 121.220 134.095 122.095 134.425 ;
        RECT 122.265 134.095 123.015 134.425 ;
        RECT 121.220 133.635 121.390 134.095 ;
        RECT 122.265 133.925 122.465 134.095 ;
        RECT 123.185 133.965 123.355 134.545 ;
        RECT 123.545 134.175 123.875 134.425 ;
        RECT 123.130 133.925 123.355 133.965 ;
        RECT 120.030 133.465 120.435 133.635 ;
        RECT 120.605 133.465 121.390 133.635 ;
        RECT 121.665 133.185 121.875 133.715 ;
        RECT 122.135 133.400 122.465 133.925 ;
        RECT 122.975 133.840 123.355 133.925 ;
        RECT 122.635 133.185 122.805 133.795 ;
        RECT 122.975 133.405 123.305 133.840 ;
        RECT 123.565 133.185 123.795 134.005 ;
        RECT 124.045 133.985 124.295 134.585 ;
        RECT 125.375 134.155 125.710 134.425 ;
        RECT 123.965 133.355 124.295 133.985 ;
        RECT 124.465 133.185 124.675 134.005 ;
        RECT 125.880 133.985 126.050 134.585 ;
        RECT 126.900 134.555 127.985 134.725 ;
        RECT 126.220 134.175 126.555 134.425 ;
        RECT 126.745 134.095 127.075 134.385 ;
        RECT 125.365 133.185 125.675 133.985 ;
        RECT 125.880 133.355 126.575 133.985 ;
        RECT 127.245 133.925 127.415 134.555 ;
        RECT 128.155 134.425 128.475 134.805 ;
        RECT 127.585 134.175 127.915 134.385 ;
        RECT 128.095 134.175 128.475 134.425 ;
        RECT 128.665 134.385 129.040 134.805 ;
        RECT 129.210 134.725 129.380 134.975 ;
        RECT 129.550 134.895 129.880 135.735 ;
        RECT 130.050 134.975 130.715 135.565 ;
        RECT 129.210 134.555 130.130 134.725 ;
        RECT 129.960 134.385 130.130 134.555 ;
        RECT 128.665 134.375 129.150 134.385 ;
        RECT 128.645 134.205 129.150 134.375 ;
        RECT 128.665 134.175 129.150 134.205 ;
        RECT 129.340 134.175 129.790 134.385 ;
        RECT 129.960 134.175 130.295 134.385 ;
        RECT 130.465 134.005 130.715 134.975 ;
        RECT 126.905 133.745 127.415 133.925 ;
        RECT 127.820 133.835 129.520 134.005 ;
        RECT 127.820 133.745 128.205 133.835 ;
        RECT 126.905 133.355 127.235 133.745 ;
        RECT 127.405 133.405 128.590 133.575 ;
        RECT 128.850 133.185 129.020 133.655 ;
        RECT 129.190 133.370 129.520 133.835 ;
        RECT 129.690 133.185 129.860 134.005 ;
        RECT 130.030 133.365 130.715 134.005 ;
        RECT 130.905 134.680 131.210 135.465 ;
        RECT 131.390 135.265 132.075 135.735 ;
        RECT 131.385 134.745 132.080 135.055 ;
        RECT 130.905 133.875 131.080 134.680 ;
        RECT 132.255 134.575 132.540 135.520 ;
        RECT 132.715 135.285 133.045 135.735 ;
        RECT 133.215 135.115 133.385 135.545 ;
        RECT 131.680 134.425 132.540 134.575 ;
        RECT 131.255 134.405 132.540 134.425 ;
        RECT 132.710 134.885 133.385 135.115 ;
        RECT 131.255 134.045 132.240 134.405 ;
        RECT 132.710 134.235 132.945 134.885 ;
        RECT 130.905 133.355 131.145 133.875 ;
        RECT 132.070 133.710 132.240 134.045 ;
        RECT 132.410 133.905 132.945 134.235 ;
        RECT 132.725 133.755 132.945 133.905 ;
        RECT 133.115 133.865 133.415 134.715 ;
        RECT 133.645 134.645 134.855 135.735 ;
        RECT 133.645 133.935 134.165 134.475 ;
        RECT 134.335 134.105 134.855 134.645 ;
        RECT 135.025 134.595 135.410 135.565 ;
        RECT 135.580 135.275 135.905 135.735 ;
        RECT 136.425 135.105 136.705 135.565 ;
        RECT 135.580 134.885 136.705 135.105 ;
        RECT 131.315 133.185 131.710 133.680 ;
        RECT 132.070 133.515 132.445 133.710 ;
        RECT 132.275 133.370 132.445 133.515 ;
        RECT 132.725 133.380 132.965 133.755 ;
        RECT 133.135 133.185 133.470 133.690 ;
        RECT 133.645 133.185 134.855 133.935 ;
        RECT 135.025 133.925 135.305 134.595 ;
        RECT 135.580 134.425 136.030 134.885 ;
        RECT 136.895 134.715 137.295 135.565 ;
        RECT 137.695 135.275 137.965 135.735 ;
        RECT 138.135 135.105 138.420 135.565 ;
        RECT 135.475 134.095 136.030 134.425 ;
        RECT 136.200 134.155 137.295 134.715 ;
        RECT 135.580 133.985 136.030 134.095 ;
        RECT 135.025 133.355 135.410 133.925 ;
        RECT 135.580 133.815 136.705 133.985 ;
        RECT 135.580 133.185 135.905 133.645 ;
        RECT 136.425 133.355 136.705 133.815 ;
        RECT 136.895 133.355 137.295 134.155 ;
        RECT 137.465 134.885 138.420 135.105 ;
        RECT 137.465 133.985 137.675 134.885 ;
        RECT 137.845 134.155 138.535 134.715 ;
        RECT 138.705 134.570 138.995 135.735 ;
        RECT 139.365 135.065 139.645 135.735 ;
        RECT 139.815 134.845 140.115 135.395 ;
        RECT 140.315 135.015 140.645 135.735 ;
        RECT 140.835 135.015 141.295 135.565 ;
        RECT 139.180 134.425 139.445 134.785 ;
        RECT 139.815 134.675 140.755 134.845 ;
        RECT 140.585 134.425 140.755 134.675 ;
        RECT 139.180 134.175 139.855 134.425 ;
        RECT 140.075 134.175 140.415 134.425 ;
        RECT 140.585 134.095 140.875 134.425 ;
        RECT 140.585 134.005 140.755 134.095 ;
        RECT 137.465 133.815 138.420 133.985 ;
        RECT 137.695 133.185 137.965 133.645 ;
        RECT 138.135 133.355 138.420 133.815 ;
        RECT 138.705 133.185 138.995 133.910 ;
        RECT 139.365 133.815 140.755 134.005 ;
        RECT 139.365 133.455 139.695 133.815 ;
        RECT 141.045 133.645 141.295 135.015 ;
        RECT 141.670 134.765 142.000 135.565 ;
        RECT 142.170 134.935 142.500 135.735 ;
        RECT 142.800 134.765 143.130 135.565 ;
        RECT 143.775 134.935 144.025 135.735 ;
        RECT 141.670 134.595 144.105 134.765 ;
        RECT 144.295 134.595 144.465 135.735 ;
        RECT 144.635 134.595 144.975 135.565 ;
        RECT 145.235 135.065 145.405 135.565 ;
        RECT 145.575 135.235 145.905 135.735 ;
        RECT 145.235 134.895 145.900 135.065 ;
        RECT 141.465 134.175 141.815 134.425 ;
        RECT 142.000 133.965 142.170 134.595 ;
        RECT 142.340 134.175 142.670 134.375 ;
        RECT 142.840 134.175 143.170 134.375 ;
        RECT 143.340 134.175 143.760 134.375 ;
        RECT 143.935 134.345 144.105 134.595 ;
        RECT 143.935 134.175 144.630 134.345 ;
        RECT 144.800 134.035 144.975 134.595 ;
        RECT 145.150 134.075 145.500 134.725 ;
        RECT 140.315 133.185 140.565 133.645 ;
        RECT 140.735 133.355 141.295 133.645 ;
        RECT 141.670 133.355 142.170 133.965 ;
        RECT 142.800 133.835 144.025 134.005 ;
        RECT 144.745 133.985 144.975 134.035 ;
        RECT 142.800 133.355 143.130 133.835 ;
        RECT 143.300 133.185 143.525 133.645 ;
        RECT 143.695 133.355 144.025 133.835 ;
        RECT 144.215 133.185 144.465 133.985 ;
        RECT 144.635 133.355 144.975 133.985 ;
        RECT 145.670 133.905 145.900 134.895 ;
        RECT 145.235 133.735 145.900 133.905 ;
        RECT 145.235 133.445 145.405 133.735 ;
        RECT 145.575 133.185 145.905 133.565 ;
        RECT 146.075 133.445 146.260 135.565 ;
        RECT 146.500 135.275 146.765 135.735 ;
        RECT 146.935 135.140 147.185 135.565 ;
        RECT 147.395 135.290 148.500 135.460 ;
        RECT 146.880 135.010 147.185 135.140 ;
        RECT 146.430 133.815 146.710 134.765 ;
        RECT 146.880 133.905 147.050 135.010 ;
        RECT 147.220 134.225 147.460 134.820 ;
        RECT 147.630 134.755 148.160 135.120 ;
        RECT 147.630 134.055 147.800 134.755 ;
        RECT 148.330 134.675 148.500 135.290 ;
        RECT 148.670 134.935 148.840 135.735 ;
        RECT 149.010 135.235 149.260 135.565 ;
        RECT 149.485 135.265 150.370 135.435 ;
        RECT 148.330 134.585 148.840 134.675 ;
        RECT 146.880 133.775 147.105 133.905 ;
        RECT 147.275 133.835 147.800 134.055 ;
        RECT 147.970 134.415 148.840 134.585 ;
        RECT 146.515 133.185 146.765 133.645 ;
        RECT 146.935 133.635 147.105 133.775 ;
        RECT 147.970 133.635 148.140 134.415 ;
        RECT 148.670 134.345 148.840 134.415 ;
        RECT 148.350 134.165 148.550 134.195 ;
        RECT 149.010 134.165 149.180 135.235 ;
        RECT 149.350 134.345 149.540 135.065 ;
        RECT 148.350 133.865 149.180 134.165 ;
        RECT 149.710 134.135 150.030 135.095 ;
        RECT 146.935 133.465 147.270 133.635 ;
        RECT 147.465 133.465 148.140 133.635 ;
        RECT 148.460 133.185 148.830 133.685 ;
        RECT 149.010 133.635 149.180 133.865 ;
        RECT 149.565 133.805 150.030 134.135 ;
        RECT 150.200 134.425 150.370 135.265 ;
        RECT 150.550 135.235 150.865 135.735 ;
        RECT 151.095 135.005 151.435 135.565 ;
        RECT 150.540 134.630 151.435 135.005 ;
        RECT 151.605 134.725 151.775 135.735 ;
        RECT 151.245 134.425 151.435 134.630 ;
        RECT 151.945 134.675 152.275 135.520 ;
        RECT 151.945 134.595 152.335 134.675 ;
        RECT 152.505 134.645 155.095 135.735 ;
        RECT 152.120 134.545 152.335 134.595 ;
        RECT 150.200 134.095 151.075 134.425 ;
        RECT 151.245 134.095 151.995 134.425 ;
        RECT 150.200 133.635 150.370 134.095 ;
        RECT 151.245 133.925 151.445 134.095 ;
        RECT 152.165 133.965 152.335 134.545 ;
        RECT 152.110 133.925 152.335 133.965 ;
        RECT 149.010 133.465 149.415 133.635 ;
        RECT 149.585 133.465 150.370 133.635 ;
        RECT 150.645 133.185 150.855 133.715 ;
        RECT 151.115 133.400 151.445 133.925 ;
        RECT 151.955 133.840 152.335 133.925 ;
        RECT 152.505 133.955 153.715 134.475 ;
        RECT 153.885 134.125 155.095 134.645 ;
        RECT 155.725 134.645 156.935 135.735 ;
        RECT 155.725 134.105 156.245 134.645 ;
        RECT 151.615 133.185 151.785 133.795 ;
        RECT 151.955 133.405 152.285 133.840 ;
        RECT 152.505 133.185 155.095 133.955 ;
        RECT 156.415 133.935 156.935 134.475 ;
        RECT 155.725 133.185 156.935 133.935 ;
        RECT 22.700 133.015 157.020 133.185 ;
        RECT 22.785 132.265 23.995 133.015 ;
        RECT 22.785 131.725 23.305 132.265 ;
        RECT 24.165 132.245 25.835 133.015 ;
        RECT 26.005 132.340 26.265 132.845 ;
        RECT 26.445 132.635 26.775 133.015 ;
        RECT 26.955 132.465 27.125 132.845 ;
        RECT 23.475 131.555 23.995 132.095 ;
        RECT 24.165 131.725 24.915 132.245 ;
        RECT 25.085 131.555 25.835 132.075 ;
        RECT 22.785 130.465 23.995 131.555 ;
        RECT 24.165 130.465 25.835 131.555 ;
        RECT 26.005 131.540 26.175 132.340 ;
        RECT 26.460 132.295 27.125 132.465 ;
        RECT 26.460 132.040 26.630 132.295 ;
        RECT 28.325 132.205 28.565 133.015 ;
        RECT 28.735 132.205 29.065 132.845 ;
        RECT 29.235 132.205 29.505 133.015 ;
        RECT 29.775 132.465 29.945 132.755 ;
        RECT 30.115 132.635 30.445 133.015 ;
        RECT 29.775 132.295 30.440 132.465 ;
        RECT 26.345 131.710 26.630 132.040 ;
        RECT 26.865 131.745 27.195 132.115 ;
        RECT 28.305 131.775 28.655 132.025 ;
        RECT 26.460 131.565 26.630 131.710 ;
        RECT 28.825 131.605 28.995 132.205 ;
        RECT 29.165 131.775 29.515 132.025 ;
        RECT 26.005 130.635 26.275 131.540 ;
        RECT 26.460 131.395 27.125 131.565 ;
        RECT 26.445 130.465 26.775 131.225 ;
        RECT 26.955 130.635 27.125 131.395 ;
        RECT 28.315 131.435 28.995 131.605 ;
        RECT 28.315 130.650 28.645 131.435 ;
        RECT 29.175 130.465 29.505 131.605 ;
        RECT 29.690 131.475 30.040 132.125 ;
        RECT 30.210 131.305 30.440 132.295 ;
        RECT 29.775 131.135 30.440 131.305 ;
        RECT 29.775 130.635 29.945 131.135 ;
        RECT 30.115 130.465 30.445 130.965 ;
        RECT 30.615 130.635 30.800 132.755 ;
        RECT 31.055 132.555 31.305 133.015 ;
        RECT 31.475 132.565 31.810 132.735 ;
        RECT 32.005 132.565 32.680 132.735 ;
        RECT 31.475 132.425 31.645 132.565 ;
        RECT 30.970 131.435 31.250 132.385 ;
        RECT 31.420 132.295 31.645 132.425 ;
        RECT 31.420 131.190 31.590 132.295 ;
        RECT 31.815 132.145 32.340 132.365 ;
        RECT 31.760 131.380 32.000 131.975 ;
        RECT 32.170 131.445 32.340 132.145 ;
        RECT 32.510 131.785 32.680 132.565 ;
        RECT 33.000 132.515 33.370 133.015 ;
        RECT 33.550 132.565 33.955 132.735 ;
        RECT 34.125 132.565 34.910 132.735 ;
        RECT 33.550 132.335 33.720 132.565 ;
        RECT 32.890 132.035 33.720 132.335 ;
        RECT 34.105 132.065 34.570 132.395 ;
        RECT 32.890 132.005 33.090 132.035 ;
        RECT 33.210 131.785 33.380 131.855 ;
        RECT 32.510 131.615 33.380 131.785 ;
        RECT 32.870 131.525 33.380 131.615 ;
        RECT 31.420 131.060 31.725 131.190 ;
        RECT 32.170 131.080 32.700 131.445 ;
        RECT 31.040 130.465 31.305 130.925 ;
        RECT 31.475 130.635 31.725 131.060 ;
        RECT 32.870 130.910 33.040 131.525 ;
        RECT 31.935 130.740 33.040 130.910 ;
        RECT 33.210 130.465 33.380 131.265 ;
        RECT 33.550 130.965 33.720 132.035 ;
        RECT 33.890 131.135 34.080 131.855 ;
        RECT 34.250 131.105 34.570 132.065 ;
        RECT 34.740 132.105 34.910 132.565 ;
        RECT 35.185 132.485 35.395 133.015 ;
        RECT 35.655 132.275 35.985 132.800 ;
        RECT 36.155 132.405 36.325 133.015 ;
        RECT 36.495 132.360 36.825 132.795 ;
        RECT 38.055 132.465 38.225 132.755 ;
        RECT 38.395 132.635 38.725 133.015 ;
        RECT 36.495 132.275 36.875 132.360 ;
        RECT 38.055 132.295 38.720 132.465 ;
        RECT 35.785 132.105 35.985 132.275 ;
        RECT 36.650 132.235 36.875 132.275 ;
        RECT 34.740 131.775 35.615 132.105 ;
        RECT 35.785 131.775 36.535 132.105 ;
        RECT 33.550 130.635 33.800 130.965 ;
        RECT 34.740 130.935 34.910 131.775 ;
        RECT 35.785 131.570 35.975 131.775 ;
        RECT 36.705 131.655 36.875 132.235 ;
        RECT 36.660 131.605 36.875 131.655 ;
        RECT 35.080 131.195 35.975 131.570 ;
        RECT 36.485 131.525 36.875 131.605 ;
        RECT 34.025 130.765 34.910 130.935 ;
        RECT 35.090 130.465 35.405 130.965 ;
        RECT 35.635 130.635 35.975 131.195 ;
        RECT 36.145 130.465 36.315 131.475 ;
        RECT 36.485 130.680 36.815 131.525 ;
        RECT 37.970 131.475 38.320 132.125 ;
        RECT 38.490 131.305 38.720 132.295 ;
        RECT 38.055 131.135 38.720 131.305 ;
        RECT 38.055 130.635 38.225 131.135 ;
        RECT 38.395 130.465 38.725 130.965 ;
        RECT 38.895 130.635 39.080 132.755 ;
        RECT 39.335 132.555 39.585 133.015 ;
        RECT 39.755 132.565 40.090 132.735 ;
        RECT 40.285 132.565 40.960 132.735 ;
        RECT 39.755 132.425 39.925 132.565 ;
        RECT 39.250 131.435 39.530 132.385 ;
        RECT 39.700 132.295 39.925 132.425 ;
        RECT 39.700 131.190 39.870 132.295 ;
        RECT 40.095 132.145 40.620 132.365 ;
        RECT 40.040 131.380 40.280 131.975 ;
        RECT 40.450 131.445 40.620 132.145 ;
        RECT 40.790 131.785 40.960 132.565 ;
        RECT 41.280 132.515 41.650 133.015 ;
        RECT 41.830 132.565 42.235 132.735 ;
        RECT 42.405 132.565 43.190 132.735 ;
        RECT 41.830 132.335 42.000 132.565 ;
        RECT 41.170 132.035 42.000 132.335 ;
        RECT 42.385 132.065 42.850 132.395 ;
        RECT 41.170 132.005 41.370 132.035 ;
        RECT 41.490 131.785 41.660 131.855 ;
        RECT 40.790 131.615 41.660 131.785 ;
        RECT 41.150 131.525 41.660 131.615 ;
        RECT 39.700 131.060 40.005 131.190 ;
        RECT 40.450 131.080 40.980 131.445 ;
        RECT 39.320 130.465 39.585 130.925 ;
        RECT 39.755 130.635 40.005 131.060 ;
        RECT 41.150 130.910 41.320 131.525 ;
        RECT 40.215 130.740 41.320 130.910 ;
        RECT 41.490 130.465 41.660 131.265 ;
        RECT 41.830 130.965 42.000 132.035 ;
        RECT 42.170 131.135 42.360 131.855 ;
        RECT 42.530 131.105 42.850 132.065 ;
        RECT 43.020 132.105 43.190 132.565 ;
        RECT 43.465 132.485 43.675 133.015 ;
        RECT 43.935 132.275 44.265 132.800 ;
        RECT 44.435 132.405 44.605 133.015 ;
        RECT 44.775 132.360 45.105 132.795 ;
        RECT 44.775 132.275 45.155 132.360 ;
        RECT 44.065 132.105 44.265 132.275 ;
        RECT 44.930 132.235 45.155 132.275 ;
        RECT 43.020 131.775 43.895 132.105 ;
        RECT 44.065 131.775 44.815 132.105 ;
        RECT 41.830 130.635 42.080 130.965 ;
        RECT 43.020 130.935 43.190 131.775 ;
        RECT 44.065 131.570 44.255 131.775 ;
        RECT 44.985 131.655 45.155 132.235 ;
        RECT 44.940 131.605 45.155 131.655 ;
        RECT 43.360 131.195 44.255 131.570 ;
        RECT 44.765 131.525 45.155 131.605 ;
        RECT 45.325 132.340 45.585 132.845 ;
        RECT 45.765 132.635 46.095 133.015 ;
        RECT 46.275 132.465 46.445 132.845 ;
        RECT 45.325 131.540 45.495 132.340 ;
        RECT 45.780 132.295 46.445 132.465 ;
        RECT 45.780 132.040 45.950 132.295 ;
        RECT 46.705 132.245 48.375 133.015 ;
        RECT 48.545 132.290 48.835 133.015 ;
        RECT 49.005 132.245 50.675 133.015 ;
        RECT 51.125 132.385 51.505 132.835 ;
        RECT 45.665 131.710 45.950 132.040 ;
        RECT 46.185 131.745 46.515 132.115 ;
        RECT 46.705 131.725 47.455 132.245 ;
        RECT 45.780 131.565 45.950 131.710 ;
        RECT 42.305 130.765 43.190 130.935 ;
        RECT 43.370 130.465 43.685 130.965 ;
        RECT 43.915 130.635 44.255 131.195 ;
        RECT 44.425 130.465 44.595 131.475 ;
        RECT 44.765 130.680 45.095 131.525 ;
        RECT 45.325 130.635 45.595 131.540 ;
        RECT 45.780 131.395 46.445 131.565 ;
        RECT 47.625 131.555 48.375 132.075 ;
        RECT 49.005 131.725 49.755 132.245 ;
        RECT 45.765 130.465 46.095 131.225 ;
        RECT 46.275 130.635 46.445 131.395 ;
        RECT 46.705 130.465 48.375 131.555 ;
        RECT 48.545 130.465 48.835 131.630 ;
        RECT 49.925 131.555 50.675 132.075 ;
        RECT 49.005 130.465 50.675 131.555 ;
        RECT 50.865 131.435 51.095 132.125 ;
        RECT 51.275 131.935 51.505 132.385 ;
        RECT 51.685 132.235 51.915 133.015 ;
        RECT 52.095 132.305 52.525 132.835 ;
        RECT 52.095 132.055 52.340 132.305 ;
        RECT 52.705 132.105 52.915 132.725 ;
        RECT 53.085 132.285 53.415 133.015 ;
        RECT 53.605 132.275 53.920 132.650 ;
        RECT 54.175 132.275 54.345 133.015 ;
        RECT 54.595 132.445 54.765 132.650 ;
        RECT 54.990 132.615 55.365 133.015 ;
        RECT 55.535 132.445 55.705 132.795 ;
        RECT 55.890 132.615 56.220 133.015 ;
        RECT 56.390 132.445 56.560 132.795 ;
        RECT 56.730 132.615 57.110 133.015 ;
        RECT 54.595 132.275 55.095 132.445 ;
        RECT 55.535 132.275 57.130 132.445 ;
        RECT 57.300 132.340 57.575 132.685 ;
        RECT 51.275 131.255 51.615 131.935 ;
        RECT 50.855 131.055 51.615 131.255 ;
        RECT 51.805 131.755 52.340 132.055 ;
        RECT 52.520 131.755 52.915 132.105 ;
        RECT 53.110 131.755 53.400 132.105 ;
        RECT 50.855 130.665 51.115 131.055 ;
        RECT 51.285 130.465 51.615 130.875 ;
        RECT 51.805 130.645 52.135 131.755 ;
        RECT 52.305 131.375 53.345 131.575 ;
        RECT 52.305 130.645 52.495 131.375 ;
        RECT 52.665 130.465 52.995 131.195 ;
        RECT 53.175 130.645 53.345 131.375 ;
        RECT 53.605 131.235 53.775 132.275 ;
        RECT 53.945 131.405 54.295 132.105 ;
        RECT 54.465 131.775 54.755 132.105 ;
        RECT 54.925 132.025 55.095 132.275 ;
        RECT 56.960 132.105 57.130 132.275 ;
        RECT 54.925 131.855 55.350 132.025 ;
        RECT 54.925 131.575 55.095 131.855 ;
        RECT 55.745 131.685 55.915 132.105 ;
        RECT 56.135 131.775 56.790 132.105 ;
        RECT 56.960 131.775 57.235 132.105 ;
        RECT 54.510 131.405 55.095 131.575 ;
        RECT 55.265 131.515 55.915 131.685 ;
        RECT 56.960 131.605 57.130 131.775 ;
        RECT 57.405 131.605 57.575 132.340 ;
        RECT 57.745 132.245 61.255 133.015 ;
        RECT 61.515 132.465 61.685 132.845 ;
        RECT 61.865 132.635 62.195 133.015 ;
        RECT 61.515 132.295 62.180 132.465 ;
        RECT 62.375 132.340 62.635 132.845 ;
        RECT 57.745 131.725 59.395 132.245 ;
        RECT 55.265 131.235 55.435 131.515 ;
        RECT 56.470 131.435 57.130 131.605 ;
        RECT 56.470 131.315 56.640 131.435 ;
        RECT 53.605 131.065 55.435 131.235 ;
        RECT 55.605 131.145 56.640 131.315 ;
        RECT 53.605 130.645 53.865 131.065 ;
        RECT 55.605 130.895 55.775 131.145 ;
        RECT 54.035 130.465 54.365 130.895 ;
        RECT 55.030 130.725 55.775 130.895 ;
        RECT 55.965 130.805 56.640 130.975 ;
        RECT 56.000 130.645 56.640 130.805 ;
        RECT 56.810 130.465 57.090 131.265 ;
        RECT 57.300 130.635 57.575 131.605 ;
        RECT 59.565 131.555 61.255 132.075 ;
        RECT 61.445 131.745 61.775 132.115 ;
        RECT 62.010 132.040 62.180 132.295 ;
        RECT 62.010 131.710 62.295 132.040 ;
        RECT 62.010 131.565 62.180 131.710 ;
        RECT 57.745 130.465 61.255 131.555 ;
        RECT 61.515 131.395 62.180 131.565 ;
        RECT 62.465 131.540 62.635 132.340 ;
        RECT 61.515 130.635 61.685 131.395 ;
        RECT 61.865 130.465 62.195 131.225 ;
        RECT 62.365 130.635 62.635 131.540 ;
        RECT 62.840 132.275 63.455 132.845 ;
        RECT 63.625 132.505 63.840 133.015 ;
        RECT 64.070 132.505 64.350 132.835 ;
        RECT 64.530 132.505 64.770 133.015 ;
        RECT 62.840 131.255 63.155 132.275 ;
        RECT 63.325 131.605 63.495 132.105 ;
        RECT 63.745 131.775 64.010 132.335 ;
        RECT 64.180 131.605 64.350 132.505 ;
        RECT 64.520 131.775 64.875 132.335 ;
        RECT 65.110 132.275 65.365 132.845 ;
        RECT 65.535 132.615 65.865 133.015 ;
        RECT 66.290 132.480 66.820 132.845 ;
        RECT 67.010 132.675 67.285 132.845 ;
        RECT 67.005 132.505 67.285 132.675 ;
        RECT 66.290 132.445 66.465 132.480 ;
        RECT 65.535 132.275 66.465 132.445 ;
        RECT 65.110 131.605 65.280 132.275 ;
        RECT 65.535 132.105 65.705 132.275 ;
        RECT 65.450 131.775 65.705 132.105 ;
        RECT 65.930 131.775 66.125 132.105 ;
        RECT 63.325 131.435 64.750 131.605 ;
        RECT 62.840 130.635 63.375 131.255 ;
        RECT 63.545 130.465 63.875 131.265 ;
        RECT 64.360 131.260 64.750 131.435 ;
        RECT 65.110 130.635 65.445 131.605 ;
        RECT 65.615 130.465 65.785 131.605 ;
        RECT 65.955 130.805 66.125 131.775 ;
        RECT 66.295 131.145 66.465 132.275 ;
        RECT 66.635 131.485 66.805 132.285 ;
        RECT 67.010 131.685 67.285 132.505 ;
        RECT 67.455 131.485 67.645 132.845 ;
        RECT 67.825 132.480 68.335 133.015 ;
        RECT 68.555 132.205 68.800 132.810 ;
        RECT 69.245 132.245 72.755 133.015 ;
        RECT 72.925 132.265 74.135 133.015 ;
        RECT 74.305 132.290 74.595 133.015 ;
        RECT 74.765 132.265 75.975 133.015 ;
        RECT 76.345 132.385 76.675 132.745 ;
        RECT 77.295 132.555 77.545 133.015 ;
        RECT 77.715 132.555 78.275 132.845 ;
        RECT 67.845 132.035 69.075 132.205 ;
        RECT 66.635 131.315 67.645 131.485 ;
        RECT 67.815 131.470 68.565 131.660 ;
        RECT 66.295 130.975 67.420 131.145 ;
        RECT 67.815 130.805 67.985 131.470 ;
        RECT 68.735 131.225 69.075 132.035 ;
        RECT 69.245 131.725 70.895 132.245 ;
        RECT 71.065 131.555 72.755 132.075 ;
        RECT 72.925 131.725 73.445 132.265 ;
        RECT 73.615 131.555 74.135 132.095 ;
        RECT 74.765 131.725 75.285 132.265 ;
        RECT 76.345 132.195 77.735 132.385 ;
        RECT 77.565 132.105 77.735 132.195 ;
        RECT 65.955 130.635 67.985 130.805 ;
        RECT 68.155 130.465 68.325 131.225 ;
        RECT 68.560 130.815 69.075 131.225 ;
        RECT 69.245 130.465 72.755 131.555 ;
        RECT 72.925 130.465 74.135 131.555 ;
        RECT 74.305 130.465 74.595 131.630 ;
        RECT 75.455 131.555 75.975 132.095 ;
        RECT 74.765 130.465 75.975 131.555 ;
        RECT 76.160 131.775 76.835 132.025 ;
        RECT 77.055 131.775 77.395 132.025 ;
        RECT 77.565 131.775 77.855 132.105 ;
        RECT 76.160 131.415 76.425 131.775 ;
        RECT 77.565 131.525 77.735 131.775 ;
        RECT 76.795 131.355 77.735 131.525 ;
        RECT 76.345 130.465 76.625 131.135 ;
        RECT 76.795 130.805 77.095 131.355 ;
        RECT 78.025 131.185 78.275 132.555 ;
        RECT 78.445 132.245 81.955 133.015 ;
        RECT 78.445 131.725 80.095 132.245 ;
        RECT 80.265 131.555 81.955 132.075 ;
        RECT 77.295 130.465 77.625 131.185 ;
        RECT 77.815 130.635 78.275 131.185 ;
        RECT 78.445 130.465 81.955 131.555 ;
        RECT 82.135 130.645 82.395 132.835 ;
        RECT 82.655 132.645 83.325 133.015 ;
        RECT 83.505 132.465 83.815 132.835 ;
        RECT 82.585 132.265 83.815 132.465 ;
        RECT 82.585 131.595 82.875 132.265 ;
        RECT 83.995 132.085 84.225 132.725 ;
        RECT 84.405 132.285 84.695 133.015 ;
        RECT 84.905 132.285 85.195 133.015 ;
        RECT 83.055 131.775 83.520 132.085 ;
        RECT 83.700 131.775 84.225 132.085 ;
        RECT 84.405 131.775 84.705 132.105 ;
        RECT 84.895 131.775 85.195 132.105 ;
        RECT 85.375 132.085 85.605 132.725 ;
        RECT 85.785 132.465 86.095 132.835 ;
        RECT 86.275 132.645 86.945 133.015 ;
        RECT 85.785 132.265 87.015 132.465 ;
        RECT 85.375 131.775 85.900 132.085 ;
        RECT 86.080 131.775 86.545 132.085 ;
        RECT 86.725 131.595 87.015 132.265 ;
        RECT 82.585 131.375 83.355 131.595 ;
        RECT 82.565 130.465 82.905 131.195 ;
        RECT 83.085 130.645 83.355 131.375 ;
        RECT 83.535 131.355 84.695 131.595 ;
        RECT 83.535 130.645 83.765 131.355 ;
        RECT 83.935 130.465 84.265 131.175 ;
        RECT 84.435 130.645 84.695 131.355 ;
        RECT 84.905 131.355 86.065 131.595 ;
        RECT 84.905 130.645 85.165 131.355 ;
        RECT 85.335 130.465 85.665 131.175 ;
        RECT 85.835 130.645 86.065 131.355 ;
        RECT 86.245 131.375 87.015 131.595 ;
        RECT 86.245 130.645 86.515 131.375 ;
        RECT 86.695 130.465 87.035 131.195 ;
        RECT 87.205 130.645 87.465 132.835 ;
        RECT 87.735 132.465 87.905 132.755 ;
        RECT 88.075 132.635 88.405 133.015 ;
        RECT 87.735 132.295 88.400 132.465 ;
        RECT 87.650 131.475 88.000 132.125 ;
        RECT 88.170 131.305 88.400 132.295 ;
        RECT 87.735 131.135 88.400 131.305 ;
        RECT 87.735 130.635 87.905 131.135 ;
        RECT 88.075 130.465 88.405 130.965 ;
        RECT 88.575 130.635 88.760 132.755 ;
        RECT 89.015 132.555 89.265 133.015 ;
        RECT 89.435 132.565 89.770 132.735 ;
        RECT 89.965 132.565 90.640 132.735 ;
        RECT 89.435 132.425 89.605 132.565 ;
        RECT 88.930 131.435 89.210 132.385 ;
        RECT 89.380 132.295 89.605 132.425 ;
        RECT 89.380 131.190 89.550 132.295 ;
        RECT 89.775 132.145 90.300 132.365 ;
        RECT 89.720 131.380 89.960 131.975 ;
        RECT 90.130 131.445 90.300 132.145 ;
        RECT 90.470 131.785 90.640 132.565 ;
        RECT 90.960 132.515 91.330 133.015 ;
        RECT 91.510 132.565 91.915 132.735 ;
        RECT 92.085 132.565 92.870 132.735 ;
        RECT 91.510 132.335 91.680 132.565 ;
        RECT 90.850 132.035 91.680 132.335 ;
        RECT 92.065 132.065 92.530 132.395 ;
        RECT 90.850 132.005 91.050 132.035 ;
        RECT 91.170 131.785 91.340 131.855 ;
        RECT 90.470 131.615 91.340 131.785 ;
        RECT 90.830 131.525 91.340 131.615 ;
        RECT 89.380 131.060 89.685 131.190 ;
        RECT 90.130 131.080 90.660 131.445 ;
        RECT 89.000 130.465 89.265 130.925 ;
        RECT 89.435 130.635 89.685 131.060 ;
        RECT 90.830 130.910 91.000 131.525 ;
        RECT 89.895 130.740 91.000 130.910 ;
        RECT 91.170 130.465 91.340 131.265 ;
        RECT 91.510 130.965 91.680 132.035 ;
        RECT 91.850 131.135 92.040 131.855 ;
        RECT 92.210 131.105 92.530 132.065 ;
        RECT 92.700 132.105 92.870 132.565 ;
        RECT 93.145 132.485 93.355 133.015 ;
        RECT 93.615 132.275 93.945 132.800 ;
        RECT 94.115 132.405 94.285 133.015 ;
        RECT 94.455 132.360 94.785 132.795 ;
        RECT 94.455 132.275 94.835 132.360 ;
        RECT 93.745 132.105 93.945 132.275 ;
        RECT 94.610 132.235 94.835 132.275 ;
        RECT 92.700 131.775 93.575 132.105 ;
        RECT 93.745 131.775 94.495 132.105 ;
        RECT 91.510 130.635 91.760 130.965 ;
        RECT 92.700 130.935 92.870 131.775 ;
        RECT 93.745 131.570 93.935 131.775 ;
        RECT 94.665 131.655 94.835 132.235 ;
        RECT 95.005 132.245 96.675 133.015 ;
        RECT 97.045 132.385 97.375 132.745 ;
        RECT 97.995 132.555 98.245 133.015 ;
        RECT 98.415 132.555 98.975 132.845 ;
        RECT 95.005 131.725 95.755 132.245 ;
        RECT 97.045 132.195 98.435 132.385 ;
        RECT 98.265 132.105 98.435 132.195 ;
        RECT 94.620 131.605 94.835 131.655 ;
        RECT 93.040 131.195 93.935 131.570 ;
        RECT 94.445 131.525 94.835 131.605 ;
        RECT 95.925 131.555 96.675 132.075 ;
        RECT 91.985 130.765 92.870 130.935 ;
        RECT 93.050 130.465 93.365 130.965 ;
        RECT 93.595 130.635 93.935 131.195 ;
        RECT 94.105 130.465 94.275 131.475 ;
        RECT 94.445 130.680 94.775 131.525 ;
        RECT 95.005 130.465 96.675 131.555 ;
        RECT 96.860 131.775 97.535 132.025 ;
        RECT 97.755 131.775 98.095 132.025 ;
        RECT 98.265 131.775 98.555 132.105 ;
        RECT 96.860 131.415 97.125 131.775 ;
        RECT 98.265 131.525 98.435 131.775 ;
        RECT 97.495 131.355 98.435 131.525 ;
        RECT 97.045 130.465 97.325 131.135 ;
        RECT 97.495 130.805 97.795 131.355 ;
        RECT 98.725 131.185 98.975 132.555 ;
        RECT 100.065 132.290 100.355 133.015 ;
        RECT 100.525 132.245 104.035 133.015 ;
        RECT 100.525 131.725 102.175 132.245 ;
        RECT 104.210 132.195 104.485 133.015 ;
        RECT 104.655 132.375 104.985 132.845 ;
        RECT 105.155 132.545 105.325 133.015 ;
        RECT 105.495 132.375 105.825 132.845 ;
        RECT 105.995 132.545 106.285 133.015 ;
        RECT 106.670 132.505 106.910 133.015 ;
        RECT 107.090 132.505 107.370 132.835 ;
        RECT 107.600 132.505 107.815 133.015 ;
        RECT 104.655 132.365 105.825 132.375 ;
        RECT 104.655 132.195 106.255 132.365 ;
        RECT 97.995 130.465 98.325 131.185 ;
        RECT 98.515 130.635 98.975 131.185 ;
        RECT 100.065 130.465 100.355 131.630 ;
        RECT 102.345 131.555 104.035 132.075 ;
        RECT 104.210 131.825 104.930 132.025 ;
        RECT 105.100 131.825 105.870 132.025 ;
        RECT 106.040 131.655 106.255 132.195 ;
        RECT 106.565 131.775 106.920 132.335 ;
        RECT 100.525 130.465 104.035 131.555 ;
        RECT 104.210 131.435 105.325 131.645 ;
        RECT 104.210 130.635 104.485 131.435 ;
        RECT 104.655 130.465 104.985 131.265 ;
        RECT 105.155 130.805 105.325 131.435 ;
        RECT 105.495 131.435 106.255 131.655 ;
        RECT 107.090 131.605 107.260 132.505 ;
        RECT 107.430 131.775 107.695 132.335 ;
        RECT 107.985 132.275 108.600 132.845 ;
        RECT 107.945 131.605 108.115 132.105 ;
        RECT 106.690 131.435 108.115 131.605 ;
        RECT 105.495 130.975 105.825 131.435 ;
        RECT 105.995 130.805 106.295 131.265 ;
        RECT 106.690 131.260 107.080 131.435 ;
        RECT 105.155 130.635 106.295 130.805 ;
        RECT 107.565 130.465 107.895 131.265 ;
        RECT 108.285 131.255 108.600 132.275 ;
        RECT 108.805 132.245 112.315 133.015 ;
        RECT 112.950 132.250 113.405 133.015 ;
        RECT 113.680 132.635 114.980 132.845 ;
        RECT 115.235 132.655 115.565 133.015 ;
        RECT 114.810 132.485 114.980 132.635 ;
        RECT 115.735 132.515 115.995 132.845 ;
        RECT 115.765 132.505 115.995 132.515 ;
        RECT 108.805 131.725 110.455 132.245 ;
        RECT 110.625 131.555 112.315 132.075 ;
        RECT 113.880 132.025 114.100 132.425 ;
        RECT 112.945 131.825 113.435 132.025 ;
        RECT 113.625 131.815 114.100 132.025 ;
        RECT 114.345 132.025 114.555 132.425 ;
        RECT 114.810 132.360 115.565 132.485 ;
        RECT 114.810 132.315 115.655 132.360 ;
        RECT 115.385 132.195 115.655 132.315 ;
        RECT 114.345 131.815 114.675 132.025 ;
        RECT 114.845 131.755 115.255 132.060 ;
        RECT 108.065 130.635 108.600 131.255 ;
        RECT 108.805 130.465 112.315 131.555 ;
        RECT 112.950 131.585 114.125 131.645 ;
        RECT 115.485 131.620 115.655 132.195 ;
        RECT 115.455 131.585 115.655 131.620 ;
        RECT 112.950 131.475 115.655 131.585 ;
        RECT 112.950 130.855 113.205 131.475 ;
        RECT 113.795 131.415 115.595 131.475 ;
        RECT 113.795 131.385 114.125 131.415 ;
        RECT 115.825 131.315 115.995 132.505 ;
        RECT 116.255 132.465 116.425 132.755 ;
        RECT 116.595 132.635 116.925 133.015 ;
        RECT 116.255 132.295 116.920 132.465 ;
        RECT 116.170 131.475 116.520 132.125 ;
        RECT 113.455 131.215 113.640 131.305 ;
        RECT 114.230 131.215 115.065 131.225 ;
        RECT 113.455 131.015 115.065 131.215 ;
        RECT 113.455 130.975 113.685 131.015 ;
        RECT 112.950 130.635 113.285 130.855 ;
        RECT 114.290 130.465 114.645 130.845 ;
        RECT 114.815 130.635 115.065 131.015 ;
        RECT 115.315 130.465 115.565 131.245 ;
        RECT 115.735 130.635 115.995 131.315 ;
        RECT 116.690 131.305 116.920 132.295 ;
        RECT 116.255 131.135 116.920 131.305 ;
        RECT 116.255 130.635 116.425 131.135 ;
        RECT 116.595 130.465 116.925 130.965 ;
        RECT 117.095 130.635 117.280 132.755 ;
        RECT 117.535 132.555 117.785 133.015 ;
        RECT 117.955 132.565 118.290 132.735 ;
        RECT 118.485 132.565 119.160 132.735 ;
        RECT 117.955 132.425 118.125 132.565 ;
        RECT 117.450 131.435 117.730 132.385 ;
        RECT 117.900 132.295 118.125 132.425 ;
        RECT 117.900 131.190 118.070 132.295 ;
        RECT 118.295 132.145 118.820 132.365 ;
        RECT 118.240 131.380 118.480 131.975 ;
        RECT 118.650 131.445 118.820 132.145 ;
        RECT 118.990 131.785 119.160 132.565 ;
        RECT 119.480 132.515 119.850 133.015 ;
        RECT 120.030 132.565 120.435 132.735 ;
        RECT 120.605 132.565 121.390 132.735 ;
        RECT 120.030 132.335 120.200 132.565 ;
        RECT 119.370 132.035 120.200 132.335 ;
        RECT 120.585 132.065 121.050 132.395 ;
        RECT 119.370 132.005 119.570 132.035 ;
        RECT 119.690 131.785 119.860 131.855 ;
        RECT 118.990 131.615 119.860 131.785 ;
        RECT 119.350 131.525 119.860 131.615 ;
        RECT 117.900 131.060 118.205 131.190 ;
        RECT 118.650 131.080 119.180 131.445 ;
        RECT 117.520 130.465 117.785 130.925 ;
        RECT 117.955 130.635 118.205 131.060 ;
        RECT 119.350 130.910 119.520 131.525 ;
        RECT 118.415 130.740 119.520 130.910 ;
        RECT 119.690 130.465 119.860 131.265 ;
        RECT 120.030 130.965 120.200 132.035 ;
        RECT 120.370 131.135 120.560 131.855 ;
        RECT 120.730 131.105 121.050 132.065 ;
        RECT 121.220 132.105 121.390 132.565 ;
        RECT 121.665 132.485 121.875 133.015 ;
        RECT 122.135 132.275 122.465 132.800 ;
        RECT 122.635 132.405 122.805 133.015 ;
        RECT 122.975 132.360 123.305 132.795 ;
        RECT 122.975 132.275 123.355 132.360 ;
        RECT 122.265 132.105 122.465 132.275 ;
        RECT 123.130 132.235 123.355 132.275 ;
        RECT 121.220 131.775 122.095 132.105 ;
        RECT 122.265 131.775 123.015 132.105 ;
        RECT 120.030 130.635 120.280 130.965 ;
        RECT 121.220 130.935 121.390 131.775 ;
        RECT 122.265 131.570 122.455 131.775 ;
        RECT 123.185 131.655 123.355 132.235 ;
        RECT 123.525 132.245 125.195 133.015 ;
        RECT 125.825 132.290 126.115 133.015 ;
        RECT 126.285 132.290 126.545 132.845 ;
        RECT 126.715 132.570 127.145 133.015 ;
        RECT 127.380 132.445 127.550 132.845 ;
        RECT 127.720 132.615 128.440 133.015 ;
        RECT 123.525 131.725 124.275 132.245 ;
        RECT 123.140 131.605 123.355 131.655 ;
        RECT 121.560 131.195 122.455 131.570 ;
        RECT 122.965 131.525 123.355 131.605 ;
        RECT 124.445 131.555 125.195 132.075 ;
        RECT 120.505 130.765 121.390 130.935 ;
        RECT 121.570 130.465 121.885 130.965 ;
        RECT 122.115 130.635 122.455 131.195 ;
        RECT 122.625 130.465 122.795 131.475 ;
        RECT 122.965 130.680 123.295 131.525 ;
        RECT 123.525 130.465 125.195 131.555 ;
        RECT 125.825 130.465 126.115 131.630 ;
        RECT 126.285 131.575 126.460 132.290 ;
        RECT 127.380 132.275 128.260 132.445 ;
        RECT 128.610 132.400 128.780 132.845 ;
        RECT 129.355 132.505 129.755 133.015 ;
        RECT 126.630 131.775 126.885 132.105 ;
        RECT 126.285 130.635 126.545 131.575 ;
        RECT 126.715 131.295 126.885 131.775 ;
        RECT 127.110 131.485 127.440 132.105 ;
        RECT 127.610 131.725 127.900 132.105 ;
        RECT 128.090 131.555 128.260 132.275 ;
        RECT 127.740 131.385 128.260 131.555 ;
        RECT 128.430 132.230 128.780 132.400 ;
        RECT 126.715 131.125 127.475 131.295 ;
        RECT 127.740 131.195 127.910 131.385 ;
        RECT 128.430 131.205 128.600 132.230 ;
        RECT 129.020 131.745 129.280 132.335 ;
        RECT 128.800 131.445 129.280 131.745 ;
        RECT 129.480 131.445 129.740 132.335 ;
        RECT 130.005 132.195 130.235 133.015 ;
        RECT 130.405 132.215 130.735 132.845 ;
        RECT 129.985 131.775 130.315 132.025 ;
        RECT 130.485 131.615 130.735 132.215 ;
        RECT 130.905 132.195 131.115 133.015 ;
        RECT 131.345 132.265 132.555 133.015 ;
        RECT 131.345 131.725 131.865 132.265 ;
        RECT 127.305 130.900 127.475 131.125 ;
        RECT 128.190 131.035 128.600 131.205 ;
        RECT 128.775 131.095 129.715 131.265 ;
        RECT 128.190 130.900 128.445 131.035 ;
        RECT 126.715 130.465 127.045 130.865 ;
        RECT 127.305 130.730 128.445 130.900 ;
        RECT 128.775 130.845 128.945 131.095 ;
        RECT 128.190 130.635 128.445 130.730 ;
        RECT 128.615 130.675 128.945 130.845 ;
        RECT 129.115 130.465 129.365 130.925 ;
        RECT 129.535 130.635 129.715 131.095 ;
        RECT 130.005 130.465 130.235 131.605 ;
        RECT 130.405 130.635 130.735 131.615 ;
        RECT 130.905 130.465 131.115 131.605 ;
        RECT 132.035 131.555 132.555 132.095 ;
        RECT 131.345 130.465 132.555 131.555 ;
        RECT 132.735 130.635 132.995 132.845 ;
        RECT 133.175 132.535 133.485 133.015 ;
        RECT 133.665 132.365 134.005 132.845 ;
        RECT 133.335 132.195 134.005 132.365 ;
        RECT 133.335 132.105 133.505 132.195 ;
        RECT 133.165 131.775 133.505 132.105 ;
        RECT 134.175 132.025 134.385 132.710 ;
        RECT 133.905 131.775 134.385 132.025 ;
        RECT 134.565 131.775 134.835 132.710 ;
        RECT 135.085 132.105 135.330 132.710 ;
        RECT 135.510 132.395 135.800 132.845 ;
        RECT 135.970 132.565 136.260 133.015 ;
        RECT 136.430 132.395 136.695 132.845 ;
        RECT 135.510 132.225 136.695 132.395 ;
        RECT 137.440 132.385 137.725 132.845 ;
        RECT 137.895 132.555 138.165 133.015 ;
        RECT 137.440 132.215 138.395 132.385 ;
        RECT 135.085 131.775 135.345 132.105 ;
        RECT 135.690 131.775 136.175 132.025 ;
        RECT 133.335 131.605 133.505 131.775 ;
        RECT 133.335 131.435 135.820 131.605 ;
        RECT 133.165 130.465 133.975 131.265 ;
        RECT 134.145 130.635 134.475 131.435 ;
        RECT 134.660 130.465 135.400 131.265 ;
        RECT 135.570 130.635 135.820 131.435 ;
        RECT 135.990 130.685 136.175 131.775 ;
        RECT 136.345 131.440 136.675 132.025 ;
        RECT 137.325 131.485 138.015 132.045 ;
        RECT 138.185 131.315 138.395 132.215 ;
        RECT 136.370 130.465 136.695 131.265 ;
        RECT 137.440 131.095 138.395 131.315 ;
        RECT 138.565 132.045 138.965 132.845 ;
        RECT 139.155 132.385 139.435 132.845 ;
        RECT 139.955 132.555 140.280 133.015 ;
        RECT 139.155 132.215 140.280 132.385 ;
        RECT 140.450 132.275 140.835 132.845 ;
        RECT 139.830 132.105 140.280 132.215 ;
        RECT 138.565 131.485 139.660 132.045 ;
        RECT 139.830 131.775 140.385 132.105 ;
        RECT 137.440 130.635 137.725 131.095 ;
        RECT 137.895 130.465 138.165 130.925 ;
        RECT 138.565 130.635 138.965 131.485 ;
        RECT 139.830 131.315 140.280 131.775 ;
        RECT 140.555 131.605 140.835 132.275 ;
        RECT 141.005 132.215 141.700 132.845 ;
        RECT 141.905 132.215 142.215 133.015 ;
        RECT 142.845 132.215 143.155 133.015 ;
        RECT 143.360 132.215 144.055 132.845 ;
        RECT 144.225 132.265 145.435 133.015 ;
        RECT 145.770 132.505 146.010 133.015 ;
        RECT 146.190 132.505 146.470 132.835 ;
        RECT 146.700 132.505 146.915 133.015 ;
        RECT 141.025 131.775 141.360 132.025 ;
        RECT 141.530 131.615 141.700 132.215 ;
        RECT 141.870 131.775 142.205 132.045 ;
        RECT 142.855 131.775 143.190 132.045 ;
        RECT 143.360 131.615 143.530 132.215 ;
        RECT 143.700 131.775 144.035 132.025 ;
        RECT 144.225 131.725 144.745 132.265 ;
        RECT 139.155 131.095 140.280 131.315 ;
        RECT 139.155 130.635 139.435 131.095 ;
        RECT 139.955 130.465 140.280 130.925 ;
        RECT 140.450 130.635 140.835 131.605 ;
        RECT 141.005 130.465 141.265 131.605 ;
        RECT 141.435 130.635 141.765 131.615 ;
        RECT 141.935 130.465 142.215 131.605 ;
        RECT 142.845 130.465 143.125 131.605 ;
        RECT 143.295 130.635 143.625 131.615 ;
        RECT 143.795 130.465 144.055 131.605 ;
        RECT 144.915 131.555 145.435 132.095 ;
        RECT 145.665 131.775 146.020 132.335 ;
        RECT 146.190 131.605 146.360 132.505 ;
        RECT 146.530 131.775 146.795 132.335 ;
        RECT 147.085 132.275 147.700 132.845 ;
        RECT 147.045 131.605 147.215 132.105 ;
        RECT 144.225 130.465 145.435 131.555 ;
        RECT 145.790 131.435 147.215 131.605 ;
        RECT 145.790 131.260 146.180 131.435 ;
        RECT 146.665 130.465 146.995 131.265 ;
        RECT 147.385 131.255 147.700 132.275 ;
        RECT 147.165 130.635 147.700 131.255 ;
        RECT 147.905 132.275 148.290 132.845 ;
        RECT 148.460 132.555 148.785 133.015 ;
        RECT 149.305 132.385 149.585 132.845 ;
        RECT 147.905 131.605 148.185 132.275 ;
        RECT 148.460 132.215 149.585 132.385 ;
        RECT 148.460 132.105 148.910 132.215 ;
        RECT 148.355 131.775 148.910 132.105 ;
        RECT 149.775 132.045 150.175 132.845 ;
        RECT 150.575 132.555 150.845 133.015 ;
        RECT 151.015 132.385 151.300 132.845 ;
        RECT 147.905 130.635 148.290 131.605 ;
        RECT 148.460 131.315 148.910 131.775 ;
        RECT 149.080 131.485 150.175 132.045 ;
        RECT 148.460 131.095 149.585 131.315 ;
        RECT 148.460 130.465 148.785 130.925 ;
        RECT 149.305 130.635 149.585 131.095 ;
        RECT 149.775 130.635 150.175 131.485 ;
        RECT 150.345 132.215 151.300 132.385 ;
        RECT 151.585 132.290 151.875 133.015 ;
        RECT 152.045 132.275 152.430 132.845 ;
        RECT 152.600 132.555 152.925 133.015 ;
        RECT 153.445 132.385 153.725 132.845 ;
        RECT 150.345 131.315 150.555 132.215 ;
        RECT 150.725 131.485 151.415 132.045 ;
        RECT 150.345 131.095 151.300 131.315 ;
        RECT 150.575 130.465 150.845 130.925 ;
        RECT 151.015 130.635 151.300 131.095 ;
        RECT 151.585 130.465 151.875 131.630 ;
        RECT 152.045 131.605 152.325 132.275 ;
        RECT 152.600 132.215 153.725 132.385 ;
        RECT 152.600 132.105 153.050 132.215 ;
        RECT 152.495 131.775 153.050 132.105 ;
        RECT 153.915 132.045 154.315 132.845 ;
        RECT 154.715 132.555 154.985 133.015 ;
        RECT 155.155 132.385 155.440 132.845 ;
        RECT 152.045 130.635 152.430 131.605 ;
        RECT 152.600 131.315 153.050 131.775 ;
        RECT 153.220 131.485 154.315 132.045 ;
        RECT 152.600 131.095 153.725 131.315 ;
        RECT 152.600 130.465 152.925 130.925 ;
        RECT 153.445 130.635 153.725 131.095 ;
        RECT 153.915 130.635 154.315 131.485 ;
        RECT 154.485 132.215 155.440 132.385 ;
        RECT 155.725 132.265 156.935 133.015 ;
        RECT 154.485 131.315 154.695 132.215 ;
        RECT 154.865 131.485 155.555 132.045 ;
        RECT 155.725 131.555 156.245 132.095 ;
        RECT 156.415 131.725 156.935 132.265 ;
        RECT 154.485 131.095 155.440 131.315 ;
        RECT 154.715 130.465 154.985 130.925 ;
        RECT 155.155 130.635 155.440 131.095 ;
        RECT 155.725 130.465 156.935 131.555 ;
        RECT 22.700 130.295 157.020 130.465 ;
        RECT 22.785 129.205 23.995 130.295 ;
        RECT 24.255 129.625 24.425 130.125 ;
        RECT 24.595 129.795 24.925 130.295 ;
        RECT 24.255 129.455 24.920 129.625 ;
        RECT 22.785 128.495 23.305 129.035 ;
        RECT 23.475 128.665 23.995 129.205 ;
        RECT 24.170 128.635 24.520 129.285 ;
        RECT 22.785 127.745 23.995 128.495 ;
        RECT 24.690 128.465 24.920 129.455 ;
        RECT 24.255 128.295 24.920 128.465 ;
        RECT 24.255 128.005 24.425 128.295 ;
        RECT 24.595 127.745 24.925 128.125 ;
        RECT 25.095 128.005 25.280 130.125 ;
        RECT 25.520 129.835 25.785 130.295 ;
        RECT 25.955 129.700 26.205 130.125 ;
        RECT 26.415 129.850 27.520 130.020 ;
        RECT 25.900 129.570 26.205 129.700 ;
        RECT 25.450 128.375 25.730 129.325 ;
        RECT 25.900 128.465 26.070 129.570 ;
        RECT 26.240 128.785 26.480 129.380 ;
        RECT 26.650 129.315 27.180 129.680 ;
        RECT 26.650 128.615 26.820 129.315 ;
        RECT 27.350 129.235 27.520 129.850 ;
        RECT 27.690 129.495 27.860 130.295 ;
        RECT 28.030 129.795 28.280 130.125 ;
        RECT 28.505 129.825 29.390 129.995 ;
        RECT 27.350 129.145 27.860 129.235 ;
        RECT 25.900 128.335 26.125 128.465 ;
        RECT 26.295 128.395 26.820 128.615 ;
        RECT 26.990 128.975 27.860 129.145 ;
        RECT 25.535 127.745 25.785 128.205 ;
        RECT 25.955 128.195 26.125 128.335 ;
        RECT 26.990 128.195 27.160 128.975 ;
        RECT 27.690 128.905 27.860 128.975 ;
        RECT 27.370 128.725 27.570 128.755 ;
        RECT 28.030 128.725 28.200 129.795 ;
        RECT 28.370 128.905 28.560 129.625 ;
        RECT 27.370 128.425 28.200 128.725 ;
        RECT 28.730 128.695 29.050 129.655 ;
        RECT 25.955 128.025 26.290 128.195 ;
        RECT 26.485 128.025 27.160 128.195 ;
        RECT 27.480 127.745 27.850 128.245 ;
        RECT 28.030 128.195 28.200 128.425 ;
        RECT 28.585 128.365 29.050 128.695 ;
        RECT 29.220 128.985 29.390 129.825 ;
        RECT 29.570 129.795 29.885 130.295 ;
        RECT 30.115 129.565 30.455 130.125 ;
        RECT 29.560 129.190 30.455 129.565 ;
        RECT 30.625 129.285 30.795 130.295 ;
        RECT 30.265 128.985 30.455 129.190 ;
        RECT 30.965 129.235 31.295 130.080 ;
        RECT 30.965 129.155 31.355 129.235 ;
        RECT 31.525 129.205 35.035 130.295 ;
        RECT 31.140 129.105 31.355 129.155 ;
        RECT 29.220 128.655 30.095 128.985 ;
        RECT 30.265 128.655 31.015 128.985 ;
        RECT 29.220 128.195 29.390 128.655 ;
        RECT 30.265 128.485 30.465 128.655 ;
        RECT 31.185 128.525 31.355 129.105 ;
        RECT 31.130 128.485 31.355 128.525 ;
        RECT 28.030 128.025 28.435 128.195 ;
        RECT 28.605 128.025 29.390 128.195 ;
        RECT 29.665 127.745 29.875 128.275 ;
        RECT 30.135 127.960 30.465 128.485 ;
        RECT 30.975 128.400 31.355 128.485 ;
        RECT 31.525 128.515 33.175 129.035 ;
        RECT 33.345 128.685 35.035 129.205 ;
        RECT 35.665 129.130 35.955 130.295 ;
        RECT 36.125 129.205 39.635 130.295 ;
        RECT 36.125 128.515 37.775 129.035 ;
        RECT 37.945 128.685 39.635 129.205 ;
        RECT 40.265 129.185 40.525 130.125 ;
        RECT 40.695 129.895 41.025 130.295 ;
        RECT 42.170 130.030 42.425 130.125 ;
        RECT 41.285 129.860 42.425 130.030 ;
        RECT 42.595 129.915 42.925 130.085 ;
        RECT 41.285 129.635 41.455 129.860 ;
        RECT 40.695 129.465 41.455 129.635 ;
        RECT 42.170 129.725 42.425 129.860 ;
        RECT 30.635 127.745 30.805 128.355 ;
        RECT 30.975 127.965 31.305 128.400 ;
        RECT 31.525 127.745 35.035 128.515 ;
        RECT 35.665 127.745 35.955 128.470 ;
        RECT 36.125 127.745 39.635 128.515 ;
        RECT 40.265 128.470 40.440 129.185 ;
        RECT 40.695 128.985 40.865 129.465 ;
        RECT 41.720 129.375 41.890 129.565 ;
        RECT 42.170 129.555 42.580 129.725 ;
        RECT 40.610 128.655 40.865 128.985 ;
        RECT 41.090 128.655 41.420 129.275 ;
        RECT 41.720 129.205 42.240 129.375 ;
        RECT 41.590 128.655 41.880 129.035 ;
        RECT 42.070 128.485 42.240 129.205 ;
        RECT 40.265 127.915 40.525 128.470 ;
        RECT 41.360 128.315 42.240 128.485 ;
        RECT 42.410 128.530 42.580 129.555 ;
        RECT 42.755 129.665 42.925 129.915 ;
        RECT 43.095 129.835 43.345 130.295 ;
        RECT 43.515 129.665 43.695 130.125 ;
        RECT 42.755 129.495 43.695 129.665 ;
        RECT 44.035 129.625 44.205 130.125 ;
        RECT 44.375 129.795 44.705 130.295 ;
        RECT 44.035 129.455 44.700 129.625 ;
        RECT 42.780 129.015 43.260 129.315 ;
        RECT 42.410 128.360 42.760 128.530 ;
        RECT 43.000 128.425 43.260 129.015 ;
        RECT 43.460 128.425 43.720 129.315 ;
        RECT 43.950 128.635 44.300 129.285 ;
        RECT 44.470 128.465 44.700 129.455 ;
        RECT 40.695 127.745 41.125 128.190 ;
        RECT 41.360 127.915 41.530 128.315 ;
        RECT 41.700 127.745 42.420 128.145 ;
        RECT 42.590 127.915 42.760 128.360 ;
        RECT 44.035 128.295 44.700 128.465 ;
        RECT 43.335 127.745 43.735 128.255 ;
        RECT 44.035 128.005 44.205 128.295 ;
        RECT 44.375 127.745 44.705 128.125 ;
        RECT 44.875 128.005 45.060 130.125 ;
        RECT 45.300 129.835 45.565 130.295 ;
        RECT 45.735 129.700 45.985 130.125 ;
        RECT 46.195 129.850 47.300 130.020 ;
        RECT 45.680 129.570 45.985 129.700 ;
        RECT 45.230 128.375 45.510 129.325 ;
        RECT 45.680 128.465 45.850 129.570 ;
        RECT 46.020 128.785 46.260 129.380 ;
        RECT 46.430 129.315 46.960 129.680 ;
        RECT 46.430 128.615 46.600 129.315 ;
        RECT 47.130 129.235 47.300 129.850 ;
        RECT 47.470 129.495 47.640 130.295 ;
        RECT 47.810 129.795 48.060 130.125 ;
        RECT 48.285 129.825 49.170 129.995 ;
        RECT 47.130 129.145 47.640 129.235 ;
        RECT 45.680 128.335 45.905 128.465 ;
        RECT 46.075 128.395 46.600 128.615 ;
        RECT 46.770 128.975 47.640 129.145 ;
        RECT 45.315 127.745 45.565 128.205 ;
        RECT 45.735 128.195 45.905 128.335 ;
        RECT 46.770 128.195 46.940 128.975 ;
        RECT 47.470 128.905 47.640 128.975 ;
        RECT 47.150 128.725 47.350 128.755 ;
        RECT 47.810 128.725 47.980 129.795 ;
        RECT 48.150 128.905 48.340 129.625 ;
        RECT 47.150 128.425 47.980 128.725 ;
        RECT 48.510 128.695 48.830 129.655 ;
        RECT 45.735 128.025 46.070 128.195 ;
        RECT 46.265 128.025 46.940 128.195 ;
        RECT 47.260 127.745 47.630 128.245 ;
        RECT 47.810 128.195 47.980 128.425 ;
        RECT 48.365 128.365 48.830 128.695 ;
        RECT 49.000 128.985 49.170 129.825 ;
        RECT 49.350 129.795 49.665 130.295 ;
        RECT 49.895 129.565 50.235 130.125 ;
        RECT 49.340 129.190 50.235 129.565 ;
        RECT 50.405 129.285 50.575 130.295 ;
        RECT 50.045 128.985 50.235 129.190 ;
        RECT 50.745 129.235 51.075 130.080 ;
        RECT 51.395 129.625 51.565 130.125 ;
        RECT 51.735 129.795 52.065 130.295 ;
        RECT 51.395 129.455 52.060 129.625 ;
        RECT 50.745 129.155 51.135 129.235 ;
        RECT 50.920 129.105 51.135 129.155 ;
        RECT 49.000 128.655 49.875 128.985 ;
        RECT 50.045 128.655 50.795 128.985 ;
        RECT 49.000 128.195 49.170 128.655 ;
        RECT 50.045 128.485 50.245 128.655 ;
        RECT 50.965 128.525 51.135 129.105 ;
        RECT 51.310 128.635 51.660 129.285 ;
        RECT 50.910 128.485 51.135 128.525 ;
        RECT 47.810 128.025 48.215 128.195 ;
        RECT 48.385 128.025 49.170 128.195 ;
        RECT 49.445 127.745 49.655 128.275 ;
        RECT 49.915 127.960 50.245 128.485 ;
        RECT 50.755 128.400 51.135 128.485 ;
        RECT 51.830 128.465 52.060 129.455 ;
        RECT 50.415 127.745 50.585 128.355 ;
        RECT 50.755 127.965 51.085 128.400 ;
        RECT 51.395 128.295 52.060 128.465 ;
        RECT 51.395 128.005 51.565 128.295 ;
        RECT 51.735 127.745 52.065 128.125 ;
        RECT 52.235 128.005 52.420 130.125 ;
        RECT 52.660 129.835 52.925 130.295 ;
        RECT 53.095 129.700 53.345 130.125 ;
        RECT 53.555 129.850 54.660 130.020 ;
        RECT 53.040 129.570 53.345 129.700 ;
        RECT 52.590 128.375 52.870 129.325 ;
        RECT 53.040 128.465 53.210 129.570 ;
        RECT 53.380 128.785 53.620 129.380 ;
        RECT 53.790 129.315 54.320 129.680 ;
        RECT 53.790 128.615 53.960 129.315 ;
        RECT 54.490 129.235 54.660 129.850 ;
        RECT 54.830 129.495 55.000 130.295 ;
        RECT 55.170 129.795 55.420 130.125 ;
        RECT 55.645 129.825 56.530 129.995 ;
        RECT 54.490 129.145 55.000 129.235 ;
        RECT 53.040 128.335 53.265 128.465 ;
        RECT 53.435 128.395 53.960 128.615 ;
        RECT 54.130 128.975 55.000 129.145 ;
        RECT 52.675 127.745 52.925 128.205 ;
        RECT 53.095 128.195 53.265 128.335 ;
        RECT 54.130 128.195 54.300 128.975 ;
        RECT 54.830 128.905 55.000 128.975 ;
        RECT 54.510 128.725 54.710 128.755 ;
        RECT 55.170 128.725 55.340 129.795 ;
        RECT 55.510 128.905 55.700 129.625 ;
        RECT 54.510 128.425 55.340 128.725 ;
        RECT 55.870 128.695 56.190 129.655 ;
        RECT 53.095 128.025 53.430 128.195 ;
        RECT 53.625 128.025 54.300 128.195 ;
        RECT 54.620 127.745 54.990 128.245 ;
        RECT 55.170 128.195 55.340 128.425 ;
        RECT 55.725 128.365 56.190 128.695 ;
        RECT 56.360 128.985 56.530 129.825 ;
        RECT 56.710 129.795 57.025 130.295 ;
        RECT 57.255 129.565 57.595 130.125 ;
        RECT 56.700 129.190 57.595 129.565 ;
        RECT 57.765 129.285 57.935 130.295 ;
        RECT 57.405 128.985 57.595 129.190 ;
        RECT 58.105 129.235 58.435 130.080 ;
        RECT 58.105 129.155 58.495 129.235 ;
        RECT 58.665 129.155 58.945 130.295 ;
        RECT 58.280 129.105 58.495 129.155 ;
        RECT 59.115 129.145 59.445 130.125 ;
        RECT 59.615 129.155 59.875 130.295 ;
        RECT 60.045 129.205 61.255 130.295 ;
        RECT 56.360 128.655 57.235 128.985 ;
        RECT 57.405 128.655 58.155 128.985 ;
        RECT 56.360 128.195 56.530 128.655 ;
        RECT 57.405 128.485 57.605 128.655 ;
        RECT 58.325 128.525 58.495 129.105 ;
        RECT 58.675 128.715 59.010 128.985 ;
        RECT 59.180 128.595 59.350 129.145 ;
        RECT 59.520 128.735 59.855 128.985 ;
        RECT 59.180 128.545 59.355 128.595 ;
        RECT 58.270 128.485 58.495 128.525 ;
        RECT 55.170 128.025 55.575 128.195 ;
        RECT 55.745 128.025 56.530 128.195 ;
        RECT 56.805 127.745 57.015 128.275 ;
        RECT 57.275 127.960 57.605 128.485 ;
        RECT 58.115 128.400 58.495 128.485 ;
        RECT 57.775 127.745 57.945 128.355 ;
        RECT 58.115 127.965 58.445 128.400 ;
        RECT 58.665 127.745 58.975 128.545 ;
        RECT 59.180 127.915 59.875 128.545 ;
        RECT 60.045 128.495 60.565 129.035 ;
        RECT 60.735 128.665 61.255 129.205 ;
        RECT 61.425 129.130 61.715 130.295 ;
        RECT 61.975 129.625 62.145 130.125 ;
        RECT 62.315 129.795 62.645 130.295 ;
        RECT 61.975 129.455 62.640 129.625 ;
        RECT 61.890 128.635 62.240 129.285 ;
        RECT 60.045 127.745 61.255 128.495 ;
        RECT 61.425 127.745 61.715 128.470 ;
        RECT 62.410 128.465 62.640 129.455 ;
        RECT 61.975 128.295 62.640 128.465 ;
        RECT 61.975 128.005 62.145 128.295 ;
        RECT 62.315 127.745 62.645 128.125 ;
        RECT 62.815 128.005 63.000 130.125 ;
        RECT 63.240 129.835 63.505 130.295 ;
        RECT 63.675 129.700 63.925 130.125 ;
        RECT 64.135 129.850 65.240 130.020 ;
        RECT 63.620 129.570 63.925 129.700 ;
        RECT 63.170 128.375 63.450 129.325 ;
        RECT 63.620 128.465 63.790 129.570 ;
        RECT 63.960 128.785 64.200 129.380 ;
        RECT 64.370 129.315 64.900 129.680 ;
        RECT 64.370 128.615 64.540 129.315 ;
        RECT 65.070 129.235 65.240 129.850 ;
        RECT 65.410 129.495 65.580 130.295 ;
        RECT 65.750 129.795 66.000 130.125 ;
        RECT 66.225 129.825 67.110 129.995 ;
        RECT 65.070 129.145 65.580 129.235 ;
        RECT 63.620 128.335 63.845 128.465 ;
        RECT 64.015 128.395 64.540 128.615 ;
        RECT 64.710 128.975 65.580 129.145 ;
        RECT 63.255 127.745 63.505 128.205 ;
        RECT 63.675 128.195 63.845 128.335 ;
        RECT 64.710 128.195 64.880 128.975 ;
        RECT 65.410 128.905 65.580 128.975 ;
        RECT 65.090 128.725 65.290 128.755 ;
        RECT 65.750 128.725 65.920 129.795 ;
        RECT 66.090 128.905 66.280 129.625 ;
        RECT 65.090 128.425 65.920 128.725 ;
        RECT 66.450 128.695 66.770 129.655 ;
        RECT 63.675 128.025 64.010 128.195 ;
        RECT 64.205 128.025 64.880 128.195 ;
        RECT 65.200 127.745 65.570 128.245 ;
        RECT 65.750 128.195 65.920 128.425 ;
        RECT 66.305 128.365 66.770 128.695 ;
        RECT 66.940 128.985 67.110 129.825 ;
        RECT 67.290 129.795 67.605 130.295 ;
        RECT 67.835 129.565 68.175 130.125 ;
        RECT 67.280 129.190 68.175 129.565 ;
        RECT 68.345 129.285 68.515 130.295 ;
        RECT 67.985 128.985 68.175 129.190 ;
        RECT 68.685 129.235 69.015 130.080 ;
        RECT 69.335 129.625 69.505 130.125 ;
        RECT 69.675 129.795 70.005 130.295 ;
        RECT 69.335 129.455 70.000 129.625 ;
        RECT 68.685 129.155 69.075 129.235 ;
        RECT 68.860 129.105 69.075 129.155 ;
        RECT 66.940 128.655 67.815 128.985 ;
        RECT 67.985 128.655 68.735 128.985 ;
        RECT 66.940 128.195 67.110 128.655 ;
        RECT 67.985 128.485 68.185 128.655 ;
        RECT 68.905 128.525 69.075 129.105 ;
        RECT 69.250 128.635 69.600 129.285 ;
        RECT 68.850 128.485 69.075 128.525 ;
        RECT 65.750 128.025 66.155 128.195 ;
        RECT 66.325 128.025 67.110 128.195 ;
        RECT 67.385 127.745 67.595 128.275 ;
        RECT 67.855 127.960 68.185 128.485 ;
        RECT 68.695 128.400 69.075 128.485 ;
        RECT 69.770 128.465 70.000 129.455 ;
        RECT 68.355 127.745 68.525 128.355 ;
        RECT 68.695 127.965 69.025 128.400 ;
        RECT 69.335 128.295 70.000 128.465 ;
        RECT 69.335 128.005 69.505 128.295 ;
        RECT 69.675 127.745 70.005 128.125 ;
        RECT 70.175 128.005 70.360 130.125 ;
        RECT 70.600 129.835 70.865 130.295 ;
        RECT 71.035 129.700 71.285 130.125 ;
        RECT 71.495 129.850 72.600 130.020 ;
        RECT 70.980 129.570 71.285 129.700 ;
        RECT 70.530 128.375 70.810 129.325 ;
        RECT 70.980 128.465 71.150 129.570 ;
        RECT 71.320 128.785 71.560 129.380 ;
        RECT 71.730 129.315 72.260 129.680 ;
        RECT 71.730 128.615 71.900 129.315 ;
        RECT 72.430 129.235 72.600 129.850 ;
        RECT 72.770 129.495 72.940 130.295 ;
        RECT 73.110 129.795 73.360 130.125 ;
        RECT 73.585 129.825 74.470 129.995 ;
        RECT 72.430 129.145 72.940 129.235 ;
        RECT 70.980 128.335 71.205 128.465 ;
        RECT 71.375 128.395 71.900 128.615 ;
        RECT 72.070 128.975 72.940 129.145 ;
        RECT 70.615 127.745 70.865 128.205 ;
        RECT 71.035 128.195 71.205 128.335 ;
        RECT 72.070 128.195 72.240 128.975 ;
        RECT 72.770 128.905 72.940 128.975 ;
        RECT 72.450 128.725 72.650 128.755 ;
        RECT 73.110 128.725 73.280 129.795 ;
        RECT 73.450 128.905 73.640 129.625 ;
        RECT 72.450 128.425 73.280 128.725 ;
        RECT 73.810 128.695 74.130 129.655 ;
        RECT 71.035 128.025 71.370 128.195 ;
        RECT 71.565 128.025 72.240 128.195 ;
        RECT 72.560 127.745 72.930 128.245 ;
        RECT 73.110 128.195 73.280 128.425 ;
        RECT 73.665 128.365 74.130 128.695 ;
        RECT 74.300 128.985 74.470 129.825 ;
        RECT 74.650 129.795 74.965 130.295 ;
        RECT 75.195 129.565 75.535 130.125 ;
        RECT 74.640 129.190 75.535 129.565 ;
        RECT 75.705 129.285 75.875 130.295 ;
        RECT 75.345 128.985 75.535 129.190 ;
        RECT 76.045 129.235 76.375 130.080 ;
        RECT 76.720 129.665 77.005 130.125 ;
        RECT 77.175 129.835 77.445 130.295 ;
        RECT 76.720 129.445 77.675 129.665 ;
        RECT 76.045 129.155 76.435 129.235 ;
        RECT 76.220 129.105 76.435 129.155 ;
        RECT 74.300 128.655 75.175 128.985 ;
        RECT 75.345 128.655 76.095 128.985 ;
        RECT 74.300 128.195 74.470 128.655 ;
        RECT 75.345 128.485 75.545 128.655 ;
        RECT 76.265 128.525 76.435 129.105 ;
        RECT 76.605 128.715 77.295 129.275 ;
        RECT 77.465 128.545 77.675 129.445 ;
        RECT 76.210 128.485 76.435 128.525 ;
        RECT 73.110 128.025 73.515 128.195 ;
        RECT 73.685 128.025 74.470 128.195 ;
        RECT 74.745 127.745 74.955 128.275 ;
        RECT 75.215 127.960 75.545 128.485 ;
        RECT 76.055 128.400 76.435 128.485 ;
        RECT 75.715 127.745 75.885 128.355 ;
        RECT 76.055 127.965 76.385 128.400 ;
        RECT 76.720 128.375 77.675 128.545 ;
        RECT 77.845 129.275 78.245 130.125 ;
        RECT 78.435 129.665 78.715 130.125 ;
        RECT 79.235 129.835 79.560 130.295 ;
        RECT 78.435 129.445 79.560 129.665 ;
        RECT 77.845 128.715 78.940 129.275 ;
        RECT 79.110 128.985 79.560 129.445 ;
        RECT 79.730 129.155 80.115 130.125 ;
        RECT 76.720 127.915 77.005 128.375 ;
        RECT 77.175 127.745 77.445 128.205 ;
        RECT 77.845 127.915 78.245 128.715 ;
        RECT 79.110 128.655 79.665 128.985 ;
        RECT 79.110 128.545 79.560 128.655 ;
        RECT 78.435 128.375 79.560 128.545 ;
        RECT 79.835 128.485 80.115 129.155 ;
        RECT 78.435 127.915 78.715 128.375 ;
        RECT 79.235 127.745 79.560 128.205 ;
        RECT 79.730 127.915 80.115 128.485 ;
        RECT 80.320 129.505 80.855 130.125 ;
        RECT 80.320 128.485 80.635 129.505 ;
        RECT 81.025 129.495 81.355 130.295 ;
        RECT 81.840 129.325 82.230 129.500 ;
        RECT 80.805 129.155 82.230 129.325 ;
        RECT 82.595 129.325 82.925 130.110 ;
        RECT 82.595 129.155 83.275 129.325 ;
        RECT 83.455 129.155 83.785 130.295 ;
        RECT 84.435 129.325 84.765 130.110 ;
        RECT 84.435 129.155 85.115 129.325 ;
        RECT 85.295 129.155 85.625 130.295 ;
        RECT 85.805 129.205 87.015 130.295 ;
        RECT 80.805 128.655 80.975 129.155 ;
        RECT 80.320 127.915 80.935 128.485 ;
        RECT 81.225 128.425 81.490 128.985 ;
        RECT 81.660 128.255 81.830 129.155 ;
        RECT 82.000 128.425 82.355 128.985 ;
        RECT 82.585 128.735 82.935 128.985 ;
        RECT 83.105 128.555 83.275 129.155 ;
        RECT 83.445 128.735 83.795 128.985 ;
        RECT 84.425 128.735 84.775 128.985 ;
        RECT 84.945 128.555 85.115 129.155 ;
        RECT 85.285 128.735 85.635 128.985 ;
        RECT 81.105 127.745 81.320 128.255 ;
        RECT 81.550 127.925 81.830 128.255 ;
        RECT 82.010 127.745 82.250 128.255 ;
        RECT 82.605 127.745 82.845 128.555 ;
        RECT 83.015 127.915 83.345 128.555 ;
        RECT 83.515 127.745 83.785 128.555 ;
        RECT 84.445 127.745 84.685 128.555 ;
        RECT 84.855 127.915 85.185 128.555 ;
        RECT 85.355 127.745 85.625 128.555 ;
        RECT 85.805 128.495 86.325 129.035 ;
        RECT 86.495 128.665 87.015 129.205 ;
        RECT 87.185 129.130 87.475 130.295 ;
        RECT 87.645 129.860 92.990 130.295 ;
        RECT 85.805 127.745 87.015 128.495 ;
        RECT 87.185 127.745 87.475 128.470 ;
        RECT 89.230 128.290 89.570 129.120 ;
        RECT 91.050 128.610 91.400 129.860 ;
        RECT 93.165 129.205 94.835 130.295 ;
        RECT 95.470 129.870 95.805 130.295 ;
        RECT 95.975 129.690 96.160 130.095 ;
        RECT 93.165 128.515 93.915 129.035 ;
        RECT 94.085 128.685 94.835 129.205 ;
        RECT 95.495 129.515 96.160 129.690 ;
        RECT 96.365 129.515 96.695 130.295 ;
        RECT 87.645 127.745 92.990 128.290 ;
        RECT 93.165 127.745 94.835 128.515 ;
        RECT 95.495 128.485 95.835 129.515 ;
        RECT 96.865 129.325 97.135 130.095 ;
        RECT 98.315 129.625 98.485 130.125 ;
        RECT 98.655 129.795 98.985 130.295 ;
        RECT 98.315 129.455 98.980 129.625 ;
        RECT 96.005 129.155 97.135 129.325 ;
        RECT 96.005 128.655 96.255 129.155 ;
        RECT 95.495 128.315 96.180 128.485 ;
        RECT 96.435 128.405 96.795 128.985 ;
        RECT 95.470 127.745 95.805 128.145 ;
        RECT 95.975 127.915 96.180 128.315 ;
        RECT 96.965 128.245 97.135 129.155 ;
        RECT 98.230 128.635 98.580 129.285 ;
        RECT 98.750 128.465 98.980 129.455 ;
        RECT 96.390 127.745 96.665 128.225 ;
        RECT 96.875 127.915 97.135 128.245 ;
        RECT 98.315 128.295 98.980 128.465 ;
        RECT 98.315 128.005 98.485 128.295 ;
        RECT 98.655 127.745 98.985 128.125 ;
        RECT 99.155 128.005 99.340 130.125 ;
        RECT 99.580 129.835 99.845 130.295 ;
        RECT 100.015 129.700 100.265 130.125 ;
        RECT 100.475 129.850 101.580 130.020 ;
        RECT 99.960 129.570 100.265 129.700 ;
        RECT 99.510 128.375 99.790 129.325 ;
        RECT 99.960 128.465 100.130 129.570 ;
        RECT 100.300 128.785 100.540 129.380 ;
        RECT 100.710 129.315 101.240 129.680 ;
        RECT 100.710 128.615 100.880 129.315 ;
        RECT 101.410 129.235 101.580 129.850 ;
        RECT 101.750 129.495 101.920 130.295 ;
        RECT 102.090 129.795 102.340 130.125 ;
        RECT 102.565 129.825 103.450 129.995 ;
        RECT 101.410 129.145 101.920 129.235 ;
        RECT 99.960 128.335 100.185 128.465 ;
        RECT 100.355 128.395 100.880 128.615 ;
        RECT 101.050 128.975 101.920 129.145 ;
        RECT 99.595 127.745 99.845 128.205 ;
        RECT 100.015 128.195 100.185 128.335 ;
        RECT 101.050 128.195 101.220 128.975 ;
        RECT 101.750 128.905 101.920 128.975 ;
        RECT 101.430 128.725 101.630 128.755 ;
        RECT 102.090 128.725 102.260 129.795 ;
        RECT 102.430 128.905 102.620 129.625 ;
        RECT 101.430 128.425 102.260 128.725 ;
        RECT 102.790 128.695 103.110 129.655 ;
        RECT 100.015 128.025 100.350 128.195 ;
        RECT 100.545 128.025 101.220 128.195 ;
        RECT 101.540 127.745 101.910 128.245 ;
        RECT 102.090 128.195 102.260 128.425 ;
        RECT 102.645 128.365 103.110 128.695 ;
        RECT 103.280 128.985 103.450 129.825 ;
        RECT 103.630 129.795 103.945 130.295 ;
        RECT 104.175 129.565 104.515 130.125 ;
        RECT 103.620 129.190 104.515 129.565 ;
        RECT 104.685 129.285 104.855 130.295 ;
        RECT 104.325 128.985 104.515 129.190 ;
        RECT 105.025 129.235 105.355 130.080 ;
        RECT 105.700 129.665 105.985 130.125 ;
        RECT 106.155 129.835 106.425 130.295 ;
        RECT 105.700 129.445 106.655 129.665 ;
        RECT 105.025 129.155 105.415 129.235 ;
        RECT 105.200 129.105 105.415 129.155 ;
        RECT 103.280 128.655 104.155 128.985 ;
        RECT 104.325 128.655 105.075 128.985 ;
        RECT 103.280 128.195 103.450 128.655 ;
        RECT 104.325 128.485 104.525 128.655 ;
        RECT 105.245 128.525 105.415 129.105 ;
        RECT 105.585 128.715 106.275 129.275 ;
        RECT 106.445 128.545 106.655 129.445 ;
        RECT 105.190 128.485 105.415 128.525 ;
        RECT 102.090 128.025 102.495 128.195 ;
        RECT 102.665 128.025 103.450 128.195 ;
        RECT 103.725 127.745 103.935 128.275 ;
        RECT 104.195 127.960 104.525 128.485 ;
        RECT 105.035 128.400 105.415 128.485 ;
        RECT 104.695 127.745 104.865 128.355 ;
        RECT 105.035 127.965 105.365 128.400 ;
        RECT 105.700 128.375 106.655 128.545 ;
        RECT 106.825 129.275 107.225 130.125 ;
        RECT 107.415 129.665 107.695 130.125 ;
        RECT 108.215 129.835 108.540 130.295 ;
        RECT 107.415 129.445 108.540 129.665 ;
        RECT 106.825 128.715 107.920 129.275 ;
        RECT 108.090 128.985 108.540 129.445 ;
        RECT 108.710 129.155 109.095 130.125 ;
        RECT 109.465 129.625 109.745 130.295 ;
        RECT 109.915 129.405 110.215 129.955 ;
        RECT 110.415 129.575 110.745 130.295 ;
        RECT 110.935 129.575 111.395 130.125 ;
        RECT 105.700 127.915 105.985 128.375 ;
        RECT 106.155 127.745 106.425 128.205 ;
        RECT 106.825 127.915 107.225 128.715 ;
        RECT 108.090 128.655 108.645 128.985 ;
        RECT 108.090 128.545 108.540 128.655 ;
        RECT 107.415 128.375 108.540 128.545 ;
        RECT 108.815 128.485 109.095 129.155 ;
        RECT 109.280 128.985 109.545 129.345 ;
        RECT 109.915 129.235 110.855 129.405 ;
        RECT 110.685 128.985 110.855 129.235 ;
        RECT 109.280 128.735 109.955 128.985 ;
        RECT 110.175 128.735 110.515 128.985 ;
        RECT 110.685 128.655 110.975 128.985 ;
        RECT 110.685 128.565 110.855 128.655 ;
        RECT 107.415 127.915 107.695 128.375 ;
        RECT 108.215 127.745 108.540 128.205 ;
        RECT 108.710 127.915 109.095 128.485 ;
        RECT 109.465 128.375 110.855 128.565 ;
        RECT 109.465 128.015 109.795 128.375 ;
        RECT 111.145 128.205 111.395 129.575 ;
        RECT 111.655 129.365 111.825 130.125 ;
        RECT 112.005 129.535 112.335 130.295 ;
        RECT 111.655 129.195 112.320 129.365 ;
        RECT 112.505 129.220 112.775 130.125 ;
        RECT 112.150 129.050 112.320 129.195 ;
        RECT 111.585 128.645 111.915 129.015 ;
        RECT 112.150 128.720 112.435 129.050 ;
        RECT 112.150 128.465 112.320 128.720 ;
        RECT 110.415 127.745 110.665 128.205 ;
        RECT 110.835 127.915 111.395 128.205 ;
        RECT 111.655 128.295 112.320 128.465 ;
        RECT 112.605 128.420 112.775 129.220 ;
        RECT 112.945 129.130 113.235 130.295 ;
        RECT 113.405 129.860 118.750 130.295 ;
        RECT 118.925 129.860 124.270 130.295 ;
        RECT 124.445 129.860 129.790 130.295 ;
        RECT 111.655 127.915 111.825 128.295 ;
        RECT 112.005 127.745 112.335 128.125 ;
        RECT 112.515 127.915 112.775 128.420 ;
        RECT 112.945 127.745 113.235 128.470 ;
        RECT 114.990 128.290 115.330 129.120 ;
        RECT 116.810 128.610 117.160 129.860 ;
        RECT 120.510 128.290 120.850 129.120 ;
        RECT 122.330 128.610 122.680 129.860 ;
        RECT 126.030 128.290 126.370 129.120 ;
        RECT 127.850 128.610 128.200 129.860 ;
        RECT 129.965 129.205 131.175 130.295 ;
        RECT 131.435 129.625 131.605 130.125 ;
        RECT 131.775 129.795 132.105 130.295 ;
        RECT 131.435 129.455 132.100 129.625 ;
        RECT 129.965 128.495 130.485 129.035 ;
        RECT 130.655 128.665 131.175 129.205 ;
        RECT 131.350 128.635 131.700 129.285 ;
        RECT 113.405 127.745 118.750 128.290 ;
        RECT 118.925 127.745 124.270 128.290 ;
        RECT 124.445 127.745 129.790 128.290 ;
        RECT 129.965 127.745 131.175 128.495 ;
        RECT 131.870 128.465 132.100 129.455 ;
        RECT 131.435 128.295 132.100 128.465 ;
        RECT 131.435 128.005 131.605 128.295 ;
        RECT 131.775 127.745 132.105 128.125 ;
        RECT 132.275 128.005 132.460 130.125 ;
        RECT 132.700 129.835 132.965 130.295 ;
        RECT 133.135 129.700 133.385 130.125 ;
        RECT 133.595 129.850 134.700 130.020 ;
        RECT 133.080 129.570 133.385 129.700 ;
        RECT 132.630 128.375 132.910 129.325 ;
        RECT 133.080 128.465 133.250 129.570 ;
        RECT 133.420 128.785 133.660 129.380 ;
        RECT 133.830 129.315 134.360 129.680 ;
        RECT 133.830 128.615 134.000 129.315 ;
        RECT 134.530 129.235 134.700 129.850 ;
        RECT 134.870 129.495 135.040 130.295 ;
        RECT 135.210 129.795 135.460 130.125 ;
        RECT 135.685 129.825 136.570 129.995 ;
        RECT 134.530 129.145 135.040 129.235 ;
        RECT 133.080 128.335 133.305 128.465 ;
        RECT 133.475 128.395 134.000 128.615 ;
        RECT 134.170 128.975 135.040 129.145 ;
        RECT 132.715 127.745 132.965 128.205 ;
        RECT 133.135 128.195 133.305 128.335 ;
        RECT 134.170 128.195 134.340 128.975 ;
        RECT 134.870 128.905 135.040 128.975 ;
        RECT 134.550 128.725 134.750 128.755 ;
        RECT 135.210 128.725 135.380 129.795 ;
        RECT 135.550 128.905 135.740 129.625 ;
        RECT 134.550 128.425 135.380 128.725 ;
        RECT 135.910 128.695 136.230 129.655 ;
        RECT 133.135 128.025 133.470 128.195 ;
        RECT 133.665 128.025 134.340 128.195 ;
        RECT 134.660 127.745 135.030 128.245 ;
        RECT 135.210 128.195 135.380 128.425 ;
        RECT 135.765 128.365 136.230 128.695 ;
        RECT 136.400 128.985 136.570 129.825 ;
        RECT 136.750 129.795 137.065 130.295 ;
        RECT 137.295 129.565 137.635 130.125 ;
        RECT 136.740 129.190 137.635 129.565 ;
        RECT 137.805 129.285 137.975 130.295 ;
        RECT 137.445 128.985 137.635 129.190 ;
        RECT 138.145 129.235 138.475 130.080 ;
        RECT 138.145 129.155 138.535 129.235 ;
        RECT 138.320 129.105 138.535 129.155 ;
        RECT 138.705 129.130 138.995 130.295 ;
        RECT 139.165 129.205 140.835 130.295 ;
        RECT 136.400 128.655 137.275 128.985 ;
        RECT 137.445 128.655 138.195 128.985 ;
        RECT 136.400 128.195 136.570 128.655 ;
        RECT 137.445 128.485 137.645 128.655 ;
        RECT 138.365 128.525 138.535 129.105 ;
        RECT 138.310 128.485 138.535 128.525 ;
        RECT 135.210 128.025 135.615 128.195 ;
        RECT 135.785 128.025 136.570 128.195 ;
        RECT 136.845 127.745 137.055 128.275 ;
        RECT 137.315 127.960 137.645 128.485 ;
        RECT 138.155 128.400 138.535 128.485 ;
        RECT 139.165 128.515 139.915 129.035 ;
        RECT 140.085 128.685 140.835 129.205 ;
        RECT 141.005 129.155 141.390 130.125 ;
        RECT 141.560 129.835 141.885 130.295 ;
        RECT 142.405 129.665 142.685 130.125 ;
        RECT 141.560 129.445 142.685 129.665 ;
        RECT 137.815 127.745 137.985 128.355 ;
        RECT 138.155 127.965 138.485 128.400 ;
        RECT 138.705 127.745 138.995 128.470 ;
        RECT 139.165 127.745 140.835 128.515 ;
        RECT 141.005 128.485 141.285 129.155 ;
        RECT 141.560 128.985 142.010 129.445 ;
        RECT 142.875 129.275 143.275 130.125 ;
        RECT 143.675 129.835 143.945 130.295 ;
        RECT 144.115 129.665 144.400 130.125 ;
        RECT 141.455 128.655 142.010 128.985 ;
        RECT 142.180 128.715 143.275 129.275 ;
        RECT 141.560 128.545 142.010 128.655 ;
        RECT 141.005 127.915 141.390 128.485 ;
        RECT 141.560 128.375 142.685 128.545 ;
        RECT 141.560 127.745 141.885 128.205 ;
        RECT 142.405 127.915 142.685 128.375 ;
        RECT 142.875 127.915 143.275 128.715 ;
        RECT 143.445 129.445 144.400 129.665 ;
        RECT 143.445 128.545 143.655 129.445 ;
        RECT 144.870 129.325 145.260 129.500 ;
        RECT 145.745 129.495 146.075 130.295 ;
        RECT 146.245 129.505 146.780 130.125 ;
        RECT 143.825 128.715 144.515 129.275 ;
        RECT 144.870 129.155 146.295 129.325 ;
        RECT 143.445 128.375 144.400 128.545 ;
        RECT 144.745 128.425 145.100 128.985 ;
        RECT 143.675 127.745 143.945 128.205 ;
        RECT 144.115 127.915 144.400 128.375 ;
        RECT 145.270 128.255 145.440 129.155 ;
        RECT 145.610 128.425 145.875 128.985 ;
        RECT 146.125 128.655 146.295 129.155 ;
        RECT 146.465 128.485 146.780 129.505 ;
        RECT 146.985 129.205 148.195 130.295 ;
        RECT 148.455 129.625 148.625 130.125 ;
        RECT 148.795 129.795 149.125 130.295 ;
        RECT 148.455 129.455 149.120 129.625 ;
        RECT 144.850 127.745 145.090 128.255 ;
        RECT 145.270 127.925 145.550 128.255 ;
        RECT 145.780 127.745 145.995 128.255 ;
        RECT 146.165 127.915 146.780 128.485 ;
        RECT 146.985 128.495 147.505 129.035 ;
        RECT 147.675 128.665 148.195 129.205 ;
        RECT 148.370 128.635 148.720 129.285 ;
        RECT 146.985 127.745 148.195 128.495 ;
        RECT 148.890 128.465 149.120 129.455 ;
        RECT 148.455 128.295 149.120 128.465 ;
        RECT 148.455 128.005 148.625 128.295 ;
        RECT 148.795 127.745 149.125 128.125 ;
        RECT 149.295 128.005 149.480 130.125 ;
        RECT 149.720 129.835 149.985 130.295 ;
        RECT 150.155 129.700 150.405 130.125 ;
        RECT 150.615 129.850 151.720 130.020 ;
        RECT 150.100 129.570 150.405 129.700 ;
        RECT 149.650 128.375 149.930 129.325 ;
        RECT 150.100 128.465 150.270 129.570 ;
        RECT 150.440 128.785 150.680 129.380 ;
        RECT 150.850 129.315 151.380 129.680 ;
        RECT 150.850 128.615 151.020 129.315 ;
        RECT 151.550 129.235 151.720 129.850 ;
        RECT 151.890 129.495 152.060 130.295 ;
        RECT 152.230 129.795 152.480 130.125 ;
        RECT 152.705 129.825 153.590 129.995 ;
        RECT 151.550 129.145 152.060 129.235 ;
        RECT 150.100 128.335 150.325 128.465 ;
        RECT 150.495 128.395 151.020 128.615 ;
        RECT 151.190 128.975 152.060 129.145 ;
        RECT 149.735 127.745 149.985 128.205 ;
        RECT 150.155 128.195 150.325 128.335 ;
        RECT 151.190 128.195 151.360 128.975 ;
        RECT 151.890 128.905 152.060 128.975 ;
        RECT 151.570 128.725 151.770 128.755 ;
        RECT 152.230 128.725 152.400 129.795 ;
        RECT 152.570 128.905 152.760 129.625 ;
        RECT 151.570 128.425 152.400 128.725 ;
        RECT 152.930 128.695 153.250 129.655 ;
        RECT 150.155 128.025 150.490 128.195 ;
        RECT 150.685 128.025 151.360 128.195 ;
        RECT 151.680 127.745 152.050 128.245 ;
        RECT 152.230 128.195 152.400 128.425 ;
        RECT 152.785 128.365 153.250 128.695 ;
        RECT 153.420 128.985 153.590 129.825 ;
        RECT 153.770 129.795 154.085 130.295 ;
        RECT 154.315 129.565 154.655 130.125 ;
        RECT 153.760 129.190 154.655 129.565 ;
        RECT 154.825 129.285 154.995 130.295 ;
        RECT 154.465 128.985 154.655 129.190 ;
        RECT 155.165 129.235 155.495 130.080 ;
        RECT 155.165 129.155 155.555 129.235 ;
        RECT 155.340 129.105 155.555 129.155 ;
        RECT 153.420 128.655 154.295 128.985 ;
        RECT 154.465 128.655 155.215 128.985 ;
        RECT 153.420 128.195 153.590 128.655 ;
        RECT 154.465 128.485 154.665 128.655 ;
        RECT 155.385 128.525 155.555 129.105 ;
        RECT 155.725 129.205 156.935 130.295 ;
        RECT 155.725 128.665 156.245 129.205 ;
        RECT 155.330 128.485 155.555 128.525 ;
        RECT 156.415 128.495 156.935 129.035 ;
        RECT 152.230 128.025 152.635 128.195 ;
        RECT 152.805 128.025 153.590 128.195 ;
        RECT 153.865 127.745 154.075 128.275 ;
        RECT 154.335 127.960 154.665 128.485 ;
        RECT 155.175 128.400 155.555 128.485 ;
        RECT 154.835 127.745 155.005 128.355 ;
        RECT 155.175 127.965 155.505 128.400 ;
        RECT 155.725 127.745 156.935 128.495 ;
        RECT 22.700 127.575 157.020 127.745 ;
        RECT 22.785 126.825 23.995 127.575 ;
        RECT 22.785 126.285 23.305 126.825 ;
        RECT 24.165 126.805 27.675 127.575 ;
        RECT 28.330 127.185 28.660 127.575 ;
        RECT 28.830 127.015 29.055 127.395 ;
        RECT 23.475 126.115 23.995 126.655 ;
        RECT 24.165 126.285 25.815 126.805 ;
        RECT 25.985 126.115 27.675 126.635 ;
        RECT 28.315 126.335 28.555 126.985 ;
        RECT 28.725 126.835 29.055 127.015 ;
        RECT 28.725 126.165 28.900 126.835 ;
        RECT 29.255 126.665 29.485 127.285 ;
        RECT 29.665 126.845 29.965 127.575 ;
        RECT 30.145 126.805 32.735 127.575 ;
        RECT 33.365 127.195 34.255 127.365 ;
        RECT 29.070 126.335 29.485 126.665 ;
        RECT 29.665 126.335 29.960 126.665 ;
        RECT 30.145 126.285 31.355 126.805 ;
        RECT 33.365 126.640 33.915 127.025 ;
        RECT 22.785 125.025 23.995 126.115 ;
        RECT 24.165 125.025 27.675 126.115 ;
        RECT 28.315 125.975 28.900 126.165 ;
        RECT 28.315 125.205 28.590 125.975 ;
        RECT 29.070 125.805 29.965 126.135 ;
        RECT 31.525 126.115 32.735 126.635 ;
        RECT 34.085 126.470 34.255 127.195 ;
        RECT 28.760 125.635 29.965 125.805 ;
        RECT 28.760 125.205 29.090 125.635 ;
        RECT 29.260 125.025 29.455 125.465 ;
        RECT 29.635 125.205 29.965 125.635 ;
        RECT 30.145 125.025 32.735 126.115 ;
        RECT 33.365 126.400 34.255 126.470 ;
        RECT 34.425 126.895 34.645 127.355 ;
        RECT 34.815 127.035 35.065 127.575 ;
        RECT 35.235 126.925 35.495 127.405 ;
        RECT 34.425 126.870 34.675 126.895 ;
        RECT 34.425 126.445 34.755 126.870 ;
        RECT 33.365 126.375 34.260 126.400 ;
        RECT 33.365 126.360 34.270 126.375 ;
        RECT 33.365 126.345 34.275 126.360 ;
        RECT 33.365 126.340 34.285 126.345 ;
        RECT 33.365 126.330 34.290 126.340 ;
        RECT 33.365 126.320 34.295 126.330 ;
        RECT 33.365 126.315 34.305 126.320 ;
        RECT 33.365 126.305 34.315 126.315 ;
        RECT 33.365 126.300 34.325 126.305 ;
        RECT 33.365 125.850 33.625 126.300 ;
        RECT 33.990 126.295 34.325 126.300 ;
        RECT 33.990 126.290 34.340 126.295 ;
        RECT 33.990 126.280 34.355 126.290 ;
        RECT 33.990 126.275 34.380 126.280 ;
        RECT 34.925 126.275 35.155 126.670 ;
        RECT 33.990 126.270 35.155 126.275 ;
        RECT 34.020 126.235 35.155 126.270 ;
        RECT 34.055 126.210 35.155 126.235 ;
        RECT 34.085 126.180 35.155 126.210 ;
        RECT 34.105 126.150 35.155 126.180 ;
        RECT 34.125 126.120 35.155 126.150 ;
        RECT 34.195 126.110 35.155 126.120 ;
        RECT 34.220 126.100 35.155 126.110 ;
        RECT 34.240 126.085 35.155 126.100 ;
        RECT 34.260 126.070 35.155 126.085 ;
        RECT 34.265 126.060 35.050 126.070 ;
        RECT 34.280 126.025 35.050 126.060 ;
        RECT 33.795 125.705 34.125 125.950 ;
        RECT 34.295 125.775 35.050 126.025 ;
        RECT 35.325 125.895 35.495 126.925 ;
        RECT 35.685 127.005 35.940 127.355 ;
        RECT 36.110 127.175 36.440 127.575 ;
        RECT 36.610 127.005 36.780 127.355 ;
        RECT 36.950 127.175 37.330 127.575 ;
        RECT 35.685 126.835 37.350 127.005 ;
        RECT 37.520 126.900 37.795 127.245 ;
        RECT 37.180 126.665 37.350 126.835 ;
        RECT 35.665 126.335 36.015 126.665 ;
        RECT 36.185 126.335 37.010 126.665 ;
        RECT 37.180 126.335 37.455 126.665 ;
        RECT 33.795 125.680 33.980 125.705 ;
        RECT 33.365 125.580 33.980 125.680 ;
        RECT 33.365 125.025 33.970 125.580 ;
        RECT 34.145 125.195 34.625 125.535 ;
        RECT 34.795 125.025 35.050 125.570 ;
        RECT 35.220 125.195 35.495 125.895 ;
        RECT 35.685 125.875 36.015 126.165 ;
        RECT 36.185 126.045 36.410 126.335 ;
        RECT 37.180 126.165 37.350 126.335 ;
        RECT 37.625 126.165 37.795 126.900 ;
        RECT 37.965 126.745 38.255 127.575 ;
        RECT 38.485 127.115 38.730 127.575 ;
        RECT 38.425 126.335 38.740 126.945 ;
        RECT 38.910 126.585 39.160 127.395 ;
        RECT 39.330 127.050 39.590 127.575 ;
        RECT 39.760 126.925 40.020 127.380 ;
        RECT 40.190 127.095 40.450 127.575 ;
        RECT 40.620 126.925 40.880 127.380 ;
        RECT 41.050 127.095 41.310 127.575 ;
        RECT 41.480 126.925 41.740 127.380 ;
        RECT 41.910 127.095 42.170 127.575 ;
        RECT 42.340 126.925 42.600 127.380 ;
        RECT 42.770 127.095 43.070 127.575 ;
        RECT 43.685 126.945 44.015 127.305 ;
        RECT 44.635 127.115 44.885 127.575 ;
        RECT 45.055 127.115 45.615 127.405 ;
        RECT 39.760 126.755 43.070 126.925 ;
        RECT 43.685 126.755 45.075 126.945 ;
        RECT 38.910 126.335 41.930 126.585 ;
        RECT 36.680 125.995 37.350 126.165 ;
        RECT 36.680 125.875 36.850 125.995 ;
        RECT 35.685 125.705 36.850 125.875 ;
        RECT 35.665 125.245 36.860 125.535 ;
        RECT 37.030 125.025 37.310 125.825 ;
        RECT 37.520 125.195 37.795 126.165 ;
        RECT 37.965 125.025 38.255 126.230 ;
        RECT 38.435 125.025 38.730 126.135 ;
        RECT 38.910 125.200 39.160 126.335 ;
        RECT 42.100 126.165 43.070 126.755 ;
        RECT 44.905 126.665 45.075 126.755 ;
        RECT 39.330 125.025 39.590 126.135 ;
        RECT 39.760 125.925 43.070 126.165 ;
        RECT 43.500 126.335 44.175 126.585 ;
        RECT 44.395 126.335 44.735 126.585 ;
        RECT 44.905 126.335 45.195 126.665 ;
        RECT 43.500 125.975 43.765 126.335 ;
        RECT 44.905 126.085 45.075 126.335 ;
        RECT 39.760 125.200 40.020 125.925 ;
        RECT 40.190 125.025 40.450 125.755 ;
        RECT 40.620 125.200 40.880 125.925 ;
        RECT 41.050 125.025 41.310 125.755 ;
        RECT 41.480 125.200 41.740 125.925 ;
        RECT 41.910 125.025 42.170 125.755 ;
        RECT 42.340 125.200 42.600 125.925 ;
        RECT 44.135 125.915 45.075 126.085 ;
        RECT 42.770 125.025 43.065 125.755 ;
        RECT 43.685 125.025 43.965 125.695 ;
        RECT 44.135 125.365 44.435 125.915 ;
        RECT 45.365 125.745 45.615 127.115 ;
        RECT 45.785 126.805 48.375 127.575 ;
        RECT 48.545 126.850 48.835 127.575 ;
        RECT 45.785 126.285 46.995 126.805 ;
        RECT 49.005 126.755 49.265 127.575 ;
        RECT 49.435 126.755 49.765 127.175 ;
        RECT 49.945 127.090 50.735 127.355 ;
        RECT 49.515 126.665 49.765 126.755 ;
        RECT 47.165 126.115 48.375 126.635 ;
        RECT 44.635 125.025 44.965 125.745 ;
        RECT 45.155 125.195 45.615 125.745 ;
        RECT 45.785 125.025 48.375 126.115 ;
        RECT 48.545 125.025 48.835 126.190 ;
        RECT 49.005 125.705 49.345 126.585 ;
        RECT 49.515 126.415 50.310 126.665 ;
        RECT 49.005 125.025 49.265 125.535 ;
        RECT 49.515 125.195 49.685 126.415 ;
        RECT 50.480 126.235 50.735 127.090 ;
        RECT 50.905 126.935 51.105 127.355 ;
        RECT 51.295 127.115 51.625 127.575 ;
        RECT 50.905 126.415 51.315 126.935 ;
        RECT 51.795 126.925 52.055 127.405 ;
        RECT 52.225 127.075 52.565 127.575 ;
        RECT 51.485 126.235 51.715 126.665 ;
        RECT 49.925 126.065 51.715 126.235 ;
        RECT 49.925 125.700 50.175 126.065 ;
        RECT 50.345 125.705 50.675 125.895 ;
        RECT 50.895 125.770 51.610 126.065 ;
        RECT 51.885 125.895 52.055 126.925 ;
        RECT 52.225 126.335 52.565 126.905 ;
        RECT 52.735 126.665 52.980 127.355 ;
        RECT 53.175 127.075 53.505 127.575 ;
        RECT 53.705 127.005 53.875 127.355 ;
        RECT 54.050 127.175 54.380 127.575 ;
        RECT 54.550 127.005 54.720 127.355 ;
        RECT 54.890 127.175 55.270 127.575 ;
        RECT 53.705 126.835 55.290 127.005 ;
        RECT 55.460 126.900 55.735 127.245 ;
        RECT 55.120 126.665 55.290 126.835 ;
        RECT 52.735 126.335 53.390 126.665 ;
        RECT 50.345 125.530 50.540 125.705 ;
        RECT 49.925 125.025 50.540 125.530 ;
        RECT 50.710 125.195 51.185 125.535 ;
        RECT 51.355 125.025 51.570 125.570 ;
        RECT 51.780 125.195 52.055 125.895 ;
        RECT 52.225 125.025 52.565 126.100 ;
        RECT 52.735 125.740 52.975 126.335 ;
        RECT 53.170 125.875 53.490 126.165 ;
        RECT 53.660 126.045 54.400 126.665 ;
        RECT 54.570 126.335 54.950 126.665 ;
        RECT 55.120 126.335 55.395 126.665 ;
        RECT 55.120 126.165 55.290 126.335 ;
        RECT 55.565 126.165 55.735 126.900 ;
        RECT 55.905 126.805 58.495 127.575 ;
        RECT 58.780 126.945 59.065 127.405 ;
        RECT 59.235 127.115 59.505 127.575 ;
        RECT 55.905 126.285 57.115 126.805 ;
        RECT 58.780 126.775 59.735 126.945 ;
        RECT 54.630 125.995 55.290 126.165 ;
        RECT 54.630 125.875 54.800 125.995 ;
        RECT 53.170 125.705 54.800 125.875 ;
        RECT 52.750 125.245 54.800 125.535 ;
        RECT 54.970 125.025 55.250 125.825 ;
        RECT 55.460 125.195 55.735 126.165 ;
        RECT 57.285 126.115 58.495 126.635 ;
        RECT 55.905 125.025 58.495 126.115 ;
        RECT 58.665 126.045 59.355 126.605 ;
        RECT 59.525 125.875 59.735 126.775 ;
        RECT 58.780 125.655 59.735 125.875 ;
        RECT 59.905 126.605 60.305 127.405 ;
        RECT 60.495 126.945 60.775 127.405 ;
        RECT 61.295 127.115 61.620 127.575 ;
        RECT 60.495 126.775 61.620 126.945 ;
        RECT 61.790 126.835 62.175 127.405 ;
        RECT 61.170 126.665 61.620 126.775 ;
        RECT 59.905 126.045 61.000 126.605 ;
        RECT 61.170 126.335 61.725 126.665 ;
        RECT 58.780 125.195 59.065 125.655 ;
        RECT 59.235 125.025 59.505 125.485 ;
        RECT 59.905 125.195 60.305 126.045 ;
        RECT 61.170 125.875 61.620 126.335 ;
        RECT 61.895 126.165 62.175 126.835 ;
        RECT 60.495 125.655 61.620 125.875 ;
        RECT 60.495 125.195 60.775 125.655 ;
        RECT 61.295 125.025 61.620 125.485 ;
        RECT 61.790 125.195 62.175 126.165 ;
        RECT 63.265 126.835 63.730 127.380 ;
        RECT 63.265 125.875 63.435 126.835 ;
        RECT 64.235 126.755 64.405 127.575 ;
        RECT 64.575 126.925 64.905 127.405 ;
        RECT 65.075 127.185 65.425 127.575 ;
        RECT 65.595 127.005 65.825 127.405 ;
        RECT 65.315 126.925 65.825 127.005 ;
        RECT 64.575 126.835 65.825 126.925 ;
        RECT 65.995 126.835 66.315 127.315 ;
        RECT 64.575 126.755 65.485 126.835 ;
        RECT 63.605 126.215 63.850 126.665 ;
        RECT 64.110 126.385 64.805 126.585 ;
        RECT 64.975 126.415 65.575 126.585 ;
        RECT 64.975 126.215 65.145 126.415 ;
        RECT 65.805 126.245 65.975 126.665 ;
        RECT 63.605 126.045 65.145 126.215 ;
        RECT 65.315 126.075 65.975 126.245 ;
        RECT 65.315 125.875 65.485 126.075 ;
        RECT 66.145 125.905 66.315 126.835 ;
        RECT 66.490 126.735 66.750 127.575 ;
        RECT 66.925 126.830 67.180 127.405 ;
        RECT 67.350 127.195 67.680 127.575 ;
        RECT 67.895 127.025 68.065 127.405 ;
        RECT 68.325 127.030 73.670 127.575 ;
        RECT 67.350 126.855 68.065 127.025 ;
        RECT 63.265 125.705 65.485 125.875 ;
        RECT 65.655 125.705 66.315 125.905 ;
        RECT 63.265 125.025 63.565 125.535 ;
        RECT 63.735 125.195 64.065 125.705 ;
        RECT 65.655 125.535 65.825 125.705 ;
        RECT 64.235 125.025 64.865 125.535 ;
        RECT 65.445 125.365 65.825 125.535 ;
        RECT 65.995 125.025 66.295 125.535 ;
        RECT 66.490 125.025 66.750 126.175 ;
        RECT 66.925 126.100 67.095 126.830 ;
        RECT 67.350 126.665 67.520 126.855 ;
        RECT 67.265 126.335 67.520 126.665 ;
        RECT 67.350 126.125 67.520 126.335 ;
        RECT 67.800 126.305 68.155 126.675 ;
        RECT 69.910 126.200 70.250 127.030 ;
        RECT 74.305 126.850 74.595 127.575 ;
        RECT 74.765 126.805 76.435 127.575 ;
        RECT 76.655 127.105 76.945 127.575 ;
        RECT 77.115 126.935 77.445 127.405 ;
        RECT 77.615 127.105 77.785 127.575 ;
        RECT 77.955 126.935 78.285 127.405 ;
        RECT 77.115 126.925 78.285 126.935 ;
        RECT 76.685 126.895 78.285 126.925 ;
        RECT 66.925 125.195 67.180 126.100 ;
        RECT 67.350 125.955 68.065 126.125 ;
        RECT 67.350 125.025 67.680 125.785 ;
        RECT 67.895 125.195 68.065 125.955 ;
        RECT 71.730 125.460 72.080 126.710 ;
        RECT 74.765 126.285 75.515 126.805 ;
        RECT 76.665 126.755 78.285 126.895 ;
        RECT 78.455 126.755 78.730 127.575 ;
        RECT 78.995 127.025 79.165 127.315 ;
        RECT 79.335 127.195 79.665 127.575 ;
        RECT 78.995 126.855 79.660 127.025 ;
        RECT 76.665 126.725 76.900 126.755 ;
        RECT 68.325 125.025 73.670 125.460 ;
        RECT 74.305 125.025 74.595 126.190 ;
        RECT 75.685 126.115 76.435 126.635 ;
        RECT 74.765 125.025 76.435 126.115 ;
        RECT 76.685 126.215 76.900 126.725 ;
        RECT 77.070 126.385 77.840 126.585 ;
        RECT 78.010 126.385 78.730 126.585 ;
        RECT 76.685 125.995 77.445 126.215 ;
        RECT 76.645 125.365 76.945 125.825 ;
        RECT 77.115 125.535 77.445 125.995 ;
        RECT 77.615 125.995 78.730 126.205 ;
        RECT 78.910 126.035 79.260 126.685 ;
        RECT 77.615 125.365 77.785 125.995 ;
        RECT 76.645 125.195 77.785 125.365 ;
        RECT 77.955 125.025 78.285 125.825 ;
        RECT 78.455 125.195 78.730 125.995 ;
        RECT 79.430 125.865 79.660 126.855 ;
        RECT 78.995 125.695 79.660 125.865 ;
        RECT 78.995 125.195 79.165 125.695 ;
        RECT 79.335 125.025 79.665 125.525 ;
        RECT 79.835 125.195 80.020 127.315 ;
        RECT 80.275 127.115 80.525 127.575 ;
        RECT 80.695 127.125 81.030 127.295 ;
        RECT 81.225 127.125 81.900 127.295 ;
        RECT 80.695 126.985 80.865 127.125 ;
        RECT 80.190 125.995 80.470 126.945 ;
        RECT 80.640 126.855 80.865 126.985 ;
        RECT 80.640 125.750 80.810 126.855 ;
        RECT 81.035 126.705 81.560 126.925 ;
        RECT 80.980 125.940 81.220 126.535 ;
        RECT 81.390 126.005 81.560 126.705 ;
        RECT 81.730 126.345 81.900 127.125 ;
        RECT 82.220 127.075 82.590 127.575 ;
        RECT 82.770 127.125 83.175 127.295 ;
        RECT 83.345 127.125 84.130 127.295 ;
        RECT 82.770 126.895 82.940 127.125 ;
        RECT 82.110 126.595 82.940 126.895 ;
        RECT 83.325 126.625 83.790 126.955 ;
        RECT 82.110 126.565 82.310 126.595 ;
        RECT 82.430 126.345 82.600 126.415 ;
        RECT 81.730 126.175 82.600 126.345 ;
        RECT 82.090 126.085 82.600 126.175 ;
        RECT 80.640 125.620 80.945 125.750 ;
        RECT 81.390 125.640 81.920 126.005 ;
        RECT 80.260 125.025 80.525 125.485 ;
        RECT 80.695 125.195 80.945 125.620 ;
        RECT 82.090 125.470 82.260 126.085 ;
        RECT 81.155 125.300 82.260 125.470 ;
        RECT 82.430 125.025 82.600 125.825 ;
        RECT 82.770 125.525 82.940 126.595 ;
        RECT 83.110 125.695 83.300 126.415 ;
        RECT 83.470 125.665 83.790 126.625 ;
        RECT 83.960 126.665 84.130 127.125 ;
        RECT 84.405 127.045 84.615 127.575 ;
        RECT 84.875 126.835 85.205 127.360 ;
        RECT 85.375 126.965 85.545 127.575 ;
        RECT 85.715 126.920 86.045 127.355 ;
        RECT 85.715 126.835 86.095 126.920 ;
        RECT 85.005 126.665 85.205 126.835 ;
        RECT 85.870 126.795 86.095 126.835 ;
        RECT 83.960 126.335 84.835 126.665 ;
        RECT 85.005 126.335 85.755 126.665 ;
        RECT 82.770 125.195 83.020 125.525 ;
        RECT 83.960 125.495 84.130 126.335 ;
        RECT 85.005 126.130 85.195 126.335 ;
        RECT 85.925 126.215 86.095 126.795 ;
        RECT 85.880 126.165 86.095 126.215 ;
        RECT 84.300 125.755 85.195 126.130 ;
        RECT 85.705 126.085 86.095 126.165 ;
        RECT 86.265 126.835 86.650 127.405 ;
        RECT 86.820 127.115 87.145 127.575 ;
        RECT 87.665 126.945 87.945 127.405 ;
        RECT 86.265 126.165 86.545 126.835 ;
        RECT 86.820 126.775 87.945 126.945 ;
        RECT 86.820 126.665 87.270 126.775 ;
        RECT 86.715 126.335 87.270 126.665 ;
        RECT 88.135 126.605 88.535 127.405 ;
        RECT 88.935 127.115 89.205 127.575 ;
        RECT 89.375 126.945 89.660 127.405 ;
        RECT 83.245 125.325 84.130 125.495 ;
        RECT 84.310 125.025 84.625 125.525 ;
        RECT 84.855 125.195 85.195 125.755 ;
        RECT 85.365 125.025 85.535 126.035 ;
        RECT 85.705 125.240 86.035 126.085 ;
        RECT 86.265 125.195 86.650 126.165 ;
        RECT 86.820 125.875 87.270 126.335 ;
        RECT 87.440 126.045 88.535 126.605 ;
        RECT 86.820 125.655 87.945 125.875 ;
        RECT 86.820 125.025 87.145 125.485 ;
        RECT 87.665 125.195 87.945 125.655 ;
        RECT 88.135 125.195 88.535 126.045 ;
        RECT 88.705 126.775 89.660 126.945 ;
        RECT 89.945 126.825 91.155 127.575 ;
        RECT 91.415 127.025 91.585 127.315 ;
        RECT 91.755 127.195 92.085 127.575 ;
        RECT 91.415 126.855 92.080 127.025 ;
        RECT 88.705 125.875 88.915 126.775 ;
        RECT 89.085 126.045 89.775 126.605 ;
        RECT 89.945 126.285 90.465 126.825 ;
        RECT 90.635 126.115 91.155 126.655 ;
        RECT 88.705 125.655 89.660 125.875 ;
        RECT 88.935 125.025 89.205 125.485 ;
        RECT 89.375 125.195 89.660 125.655 ;
        RECT 89.945 125.025 91.155 126.115 ;
        RECT 91.330 126.035 91.680 126.685 ;
        RECT 91.850 125.865 92.080 126.855 ;
        RECT 91.415 125.695 92.080 125.865 ;
        RECT 91.415 125.195 91.585 125.695 ;
        RECT 91.755 125.025 92.085 125.525 ;
        RECT 92.255 125.195 92.440 127.315 ;
        RECT 92.695 127.115 92.945 127.575 ;
        RECT 93.115 127.125 93.450 127.295 ;
        RECT 93.645 127.125 94.320 127.295 ;
        RECT 93.115 126.985 93.285 127.125 ;
        RECT 92.610 125.995 92.890 126.945 ;
        RECT 93.060 126.855 93.285 126.985 ;
        RECT 93.060 125.750 93.230 126.855 ;
        RECT 93.455 126.705 93.980 126.925 ;
        RECT 93.400 125.940 93.640 126.535 ;
        RECT 93.810 126.005 93.980 126.705 ;
        RECT 94.150 126.345 94.320 127.125 ;
        RECT 94.640 127.075 95.010 127.575 ;
        RECT 95.190 127.125 95.595 127.295 ;
        RECT 95.765 127.125 96.550 127.295 ;
        RECT 95.190 126.895 95.360 127.125 ;
        RECT 94.530 126.595 95.360 126.895 ;
        RECT 95.745 126.625 96.210 126.955 ;
        RECT 94.530 126.565 94.730 126.595 ;
        RECT 94.850 126.345 95.020 126.415 ;
        RECT 94.150 126.175 95.020 126.345 ;
        RECT 94.510 126.085 95.020 126.175 ;
        RECT 93.060 125.620 93.365 125.750 ;
        RECT 93.810 125.640 94.340 126.005 ;
        RECT 92.680 125.025 92.945 125.485 ;
        RECT 93.115 125.195 93.365 125.620 ;
        RECT 94.510 125.470 94.680 126.085 ;
        RECT 93.575 125.300 94.680 125.470 ;
        RECT 94.850 125.025 95.020 125.825 ;
        RECT 95.190 125.525 95.360 126.595 ;
        RECT 95.530 125.695 95.720 126.415 ;
        RECT 95.890 125.665 96.210 126.625 ;
        RECT 96.380 126.665 96.550 127.125 ;
        RECT 96.825 127.045 97.035 127.575 ;
        RECT 97.295 126.835 97.625 127.360 ;
        RECT 97.795 126.965 97.965 127.575 ;
        RECT 98.135 126.920 98.465 127.355 ;
        RECT 98.135 126.835 98.515 126.920 ;
        RECT 97.425 126.665 97.625 126.835 ;
        RECT 98.290 126.795 98.515 126.835 ;
        RECT 96.380 126.335 97.255 126.665 ;
        RECT 97.425 126.335 98.175 126.665 ;
        RECT 95.190 125.195 95.440 125.525 ;
        RECT 96.380 125.495 96.550 126.335 ;
        RECT 97.425 126.130 97.615 126.335 ;
        RECT 98.345 126.215 98.515 126.795 ;
        RECT 98.685 126.825 99.895 127.575 ;
        RECT 100.065 126.850 100.355 127.575 ;
        RECT 100.525 126.835 100.910 127.405 ;
        RECT 101.080 127.115 101.405 127.575 ;
        RECT 101.925 126.945 102.205 127.405 ;
        RECT 98.685 126.285 99.205 126.825 ;
        RECT 98.300 126.165 98.515 126.215 ;
        RECT 96.720 125.755 97.615 126.130 ;
        RECT 98.125 126.085 98.515 126.165 ;
        RECT 99.375 126.115 99.895 126.655 ;
        RECT 95.665 125.325 96.550 125.495 ;
        RECT 96.730 125.025 97.045 125.525 ;
        RECT 97.275 125.195 97.615 125.755 ;
        RECT 97.785 125.025 97.955 126.035 ;
        RECT 98.125 125.240 98.455 126.085 ;
        RECT 98.685 125.025 99.895 126.115 ;
        RECT 100.065 125.025 100.355 126.190 ;
        RECT 100.525 126.165 100.805 126.835 ;
        RECT 101.080 126.775 102.205 126.945 ;
        RECT 101.080 126.665 101.530 126.775 ;
        RECT 100.975 126.335 101.530 126.665 ;
        RECT 102.395 126.605 102.795 127.405 ;
        RECT 103.195 127.115 103.465 127.575 ;
        RECT 103.635 126.945 103.920 127.405 ;
        RECT 100.525 125.195 100.910 126.165 ;
        RECT 101.080 125.875 101.530 126.335 ;
        RECT 101.700 126.045 102.795 126.605 ;
        RECT 101.080 125.655 102.205 125.875 ;
        RECT 101.080 125.025 101.405 125.485 ;
        RECT 101.925 125.195 102.205 125.655 ;
        RECT 102.395 125.195 102.795 126.045 ;
        RECT 102.965 126.775 103.920 126.945 ;
        RECT 104.205 126.850 104.465 127.405 ;
        RECT 104.635 127.130 105.065 127.575 ;
        RECT 105.300 127.005 105.470 127.405 ;
        RECT 105.640 127.175 106.360 127.575 ;
        RECT 102.965 125.875 103.175 126.775 ;
        RECT 103.345 126.045 104.035 126.605 ;
        RECT 104.205 126.135 104.380 126.850 ;
        RECT 105.300 126.835 106.180 127.005 ;
        RECT 106.530 126.960 106.700 127.405 ;
        RECT 107.275 127.065 107.675 127.575 ;
        RECT 104.550 126.335 104.805 126.665 ;
        RECT 102.965 125.655 103.920 125.875 ;
        RECT 103.195 125.025 103.465 125.485 ;
        RECT 103.635 125.195 103.920 125.655 ;
        RECT 104.205 125.195 104.465 126.135 ;
        RECT 104.635 125.855 104.805 126.335 ;
        RECT 105.030 126.045 105.360 126.665 ;
        RECT 105.530 126.285 105.820 126.665 ;
        RECT 106.010 126.115 106.180 126.835 ;
        RECT 105.660 125.945 106.180 126.115 ;
        RECT 106.350 126.790 106.700 126.960 ;
        RECT 107.935 126.920 108.265 127.355 ;
        RECT 108.435 126.965 108.605 127.575 ;
        RECT 104.635 125.685 105.395 125.855 ;
        RECT 105.660 125.755 105.830 125.945 ;
        RECT 106.350 125.765 106.520 126.790 ;
        RECT 106.940 126.305 107.200 126.895 ;
        RECT 106.720 126.005 107.200 126.305 ;
        RECT 107.400 126.005 107.660 126.895 ;
        RECT 107.885 126.835 108.265 126.920 ;
        RECT 108.775 126.835 109.105 127.360 ;
        RECT 109.365 127.045 109.575 127.575 ;
        RECT 109.850 127.125 110.635 127.295 ;
        RECT 110.805 127.125 111.210 127.295 ;
        RECT 107.885 126.795 108.110 126.835 ;
        RECT 107.885 126.215 108.055 126.795 ;
        RECT 108.775 126.665 108.975 126.835 ;
        RECT 109.850 126.665 110.020 127.125 ;
        RECT 108.225 126.335 108.975 126.665 ;
        RECT 109.145 126.335 110.020 126.665 ;
        RECT 107.885 126.165 108.100 126.215 ;
        RECT 107.885 126.085 108.275 126.165 ;
        RECT 105.225 125.460 105.395 125.685 ;
        RECT 106.110 125.595 106.520 125.765 ;
        RECT 106.695 125.655 107.635 125.825 ;
        RECT 106.110 125.460 106.365 125.595 ;
        RECT 104.635 125.025 104.965 125.425 ;
        RECT 105.225 125.290 106.365 125.460 ;
        RECT 106.695 125.405 106.865 125.655 ;
        RECT 106.110 125.195 106.365 125.290 ;
        RECT 106.535 125.235 106.865 125.405 ;
        RECT 107.035 125.025 107.285 125.485 ;
        RECT 107.455 125.195 107.635 125.655 ;
        RECT 107.945 125.240 108.275 126.085 ;
        RECT 108.785 126.130 108.975 126.335 ;
        RECT 108.445 125.025 108.615 126.035 ;
        RECT 108.785 125.755 109.680 126.130 ;
        RECT 108.785 125.195 109.125 125.755 ;
        RECT 109.355 125.025 109.670 125.525 ;
        RECT 109.850 125.495 110.020 126.335 ;
        RECT 110.190 126.625 110.655 126.955 ;
        RECT 111.040 126.895 111.210 127.125 ;
        RECT 111.390 127.075 111.760 127.575 ;
        RECT 112.080 127.125 112.755 127.295 ;
        RECT 112.950 127.125 113.285 127.295 ;
        RECT 110.190 125.665 110.510 126.625 ;
        RECT 111.040 126.595 111.870 126.895 ;
        RECT 110.680 125.695 110.870 126.415 ;
        RECT 111.040 125.525 111.210 126.595 ;
        RECT 111.670 126.565 111.870 126.595 ;
        RECT 111.380 126.345 111.550 126.415 ;
        RECT 112.080 126.345 112.250 127.125 ;
        RECT 113.115 126.985 113.285 127.125 ;
        RECT 113.455 127.115 113.705 127.575 ;
        RECT 111.380 126.175 112.250 126.345 ;
        RECT 112.420 126.705 112.945 126.925 ;
        RECT 113.115 126.855 113.340 126.985 ;
        RECT 111.380 126.085 111.890 126.175 ;
        RECT 109.850 125.325 110.735 125.495 ;
        RECT 110.960 125.195 111.210 125.525 ;
        RECT 111.380 125.025 111.550 125.825 ;
        RECT 111.720 125.470 111.890 126.085 ;
        RECT 112.420 126.005 112.590 126.705 ;
        RECT 112.060 125.640 112.590 126.005 ;
        RECT 112.760 125.940 113.000 126.535 ;
        RECT 113.170 125.750 113.340 126.855 ;
        RECT 113.510 125.995 113.790 126.945 ;
        RECT 113.035 125.620 113.340 125.750 ;
        RECT 111.720 125.300 112.825 125.470 ;
        RECT 113.035 125.195 113.285 125.620 ;
        RECT 113.455 125.025 113.720 125.485 ;
        RECT 113.960 125.195 114.145 127.315 ;
        RECT 114.315 127.195 114.645 127.575 ;
        RECT 114.815 127.025 114.985 127.315 ;
        RECT 114.320 126.855 114.985 127.025 ;
        RECT 115.335 127.025 115.505 127.315 ;
        RECT 115.675 127.195 116.005 127.575 ;
        RECT 115.335 126.855 116.000 127.025 ;
        RECT 114.320 125.865 114.550 126.855 ;
        RECT 114.720 126.035 115.070 126.685 ;
        RECT 115.250 126.035 115.600 126.685 ;
        RECT 115.770 125.865 116.000 126.855 ;
        RECT 114.320 125.695 114.985 125.865 ;
        RECT 114.315 125.025 114.645 125.525 ;
        RECT 114.815 125.195 114.985 125.695 ;
        RECT 115.335 125.695 116.000 125.865 ;
        RECT 115.335 125.195 115.505 125.695 ;
        RECT 115.675 125.025 116.005 125.525 ;
        RECT 116.175 125.195 116.360 127.315 ;
        RECT 116.615 127.115 116.865 127.575 ;
        RECT 117.035 127.125 117.370 127.295 ;
        RECT 117.565 127.125 118.240 127.295 ;
        RECT 117.035 126.985 117.205 127.125 ;
        RECT 116.530 125.995 116.810 126.945 ;
        RECT 116.980 126.855 117.205 126.985 ;
        RECT 116.980 125.750 117.150 126.855 ;
        RECT 117.375 126.705 117.900 126.925 ;
        RECT 117.320 125.940 117.560 126.535 ;
        RECT 117.730 126.005 117.900 126.705 ;
        RECT 118.070 126.345 118.240 127.125 ;
        RECT 118.560 127.075 118.930 127.575 ;
        RECT 119.110 127.125 119.515 127.295 ;
        RECT 119.685 127.125 120.470 127.295 ;
        RECT 119.110 126.895 119.280 127.125 ;
        RECT 118.450 126.595 119.280 126.895 ;
        RECT 119.665 126.625 120.130 126.955 ;
        RECT 118.450 126.565 118.650 126.595 ;
        RECT 118.770 126.345 118.940 126.415 ;
        RECT 118.070 126.175 118.940 126.345 ;
        RECT 118.430 126.085 118.940 126.175 ;
        RECT 116.980 125.620 117.285 125.750 ;
        RECT 117.730 125.640 118.260 126.005 ;
        RECT 116.600 125.025 116.865 125.485 ;
        RECT 117.035 125.195 117.285 125.620 ;
        RECT 118.430 125.470 118.600 126.085 ;
        RECT 117.495 125.300 118.600 125.470 ;
        RECT 118.770 125.025 118.940 125.825 ;
        RECT 119.110 125.525 119.280 126.595 ;
        RECT 119.450 125.695 119.640 126.415 ;
        RECT 119.810 125.665 120.130 126.625 ;
        RECT 120.300 126.665 120.470 127.125 ;
        RECT 120.745 127.045 120.955 127.575 ;
        RECT 121.215 126.835 121.545 127.360 ;
        RECT 121.715 126.965 121.885 127.575 ;
        RECT 122.055 126.920 122.385 127.355 ;
        RECT 123.090 126.925 123.400 127.395 ;
        RECT 123.570 127.095 124.305 127.575 ;
        RECT 124.475 127.005 124.645 127.355 ;
        RECT 124.815 127.175 125.195 127.575 ;
        RECT 122.055 126.835 122.435 126.920 ;
        RECT 121.345 126.665 121.545 126.835 ;
        RECT 122.210 126.795 122.435 126.835 ;
        RECT 120.300 126.335 121.175 126.665 ;
        RECT 121.345 126.335 122.095 126.665 ;
        RECT 119.110 125.195 119.360 125.525 ;
        RECT 120.300 125.495 120.470 126.335 ;
        RECT 121.345 126.130 121.535 126.335 ;
        RECT 122.265 126.215 122.435 126.795 ;
        RECT 123.090 126.755 123.825 126.925 ;
        RECT 124.475 126.835 125.215 127.005 ;
        RECT 125.385 126.900 125.655 127.245 ;
        RECT 123.575 126.665 123.825 126.755 ;
        RECT 125.045 126.665 125.215 126.835 ;
        RECT 123.070 126.335 123.405 126.585 ;
        RECT 123.575 126.335 124.315 126.665 ;
        RECT 125.045 126.335 125.275 126.665 ;
        RECT 122.220 126.165 122.435 126.215 ;
        RECT 120.640 125.755 121.535 126.130 ;
        RECT 122.045 126.085 122.435 126.165 ;
        RECT 119.585 125.325 120.470 125.495 ;
        RECT 120.650 125.025 120.965 125.525 ;
        RECT 121.195 125.195 121.535 125.755 ;
        RECT 121.705 125.025 121.875 126.035 ;
        RECT 122.045 125.240 122.375 126.085 ;
        RECT 123.070 125.025 123.325 126.165 ;
        RECT 123.575 125.775 123.745 126.335 ;
        RECT 125.045 126.165 125.215 126.335 ;
        RECT 125.485 126.165 125.655 126.900 ;
        RECT 125.825 126.850 126.115 127.575 ;
        RECT 126.345 127.115 126.590 127.575 ;
        RECT 126.285 126.335 126.600 126.945 ;
        RECT 126.770 126.585 127.020 127.395 ;
        RECT 127.190 127.050 127.450 127.575 ;
        RECT 127.620 126.925 127.880 127.380 ;
        RECT 128.050 127.095 128.310 127.575 ;
        RECT 128.480 126.925 128.740 127.380 ;
        RECT 128.910 127.095 129.170 127.575 ;
        RECT 129.340 126.925 129.600 127.380 ;
        RECT 129.770 127.095 130.030 127.575 ;
        RECT 130.200 126.925 130.460 127.380 ;
        RECT 130.630 127.095 130.930 127.575 ;
        RECT 131.435 127.025 131.605 127.405 ;
        RECT 131.820 127.195 132.150 127.575 ;
        RECT 127.620 126.755 130.930 126.925 ;
        RECT 131.435 126.855 132.150 127.025 ;
        RECT 126.770 126.335 129.790 126.585 ;
        RECT 123.970 125.995 125.215 126.165 ;
        RECT 123.970 125.745 124.390 125.995 ;
        RECT 123.520 125.245 124.715 125.575 ;
        RECT 124.895 125.025 125.175 125.825 ;
        RECT 125.385 125.195 125.655 126.165 ;
        RECT 125.825 125.025 126.115 126.190 ;
        RECT 126.295 125.025 126.590 126.135 ;
        RECT 126.770 125.200 127.020 126.335 ;
        RECT 129.960 126.165 130.930 126.755 ;
        RECT 131.345 126.305 131.700 126.675 ;
        RECT 131.980 126.665 132.150 126.855 ;
        RECT 132.320 126.830 132.575 127.405 ;
        RECT 131.980 126.335 132.235 126.665 ;
        RECT 127.190 125.025 127.450 126.135 ;
        RECT 127.620 125.925 130.930 126.165 ;
        RECT 131.980 126.125 132.150 126.335 ;
        RECT 131.435 125.955 132.150 126.125 ;
        RECT 132.405 126.100 132.575 126.830 ;
        RECT 132.750 126.735 133.010 127.575 ;
        RECT 133.185 126.825 134.395 127.575 ;
        RECT 133.185 126.285 133.705 126.825 ;
        RECT 134.770 126.795 135.270 127.405 ;
        RECT 127.620 125.200 127.880 125.925 ;
        RECT 128.050 125.025 128.310 125.755 ;
        RECT 128.480 125.200 128.740 125.925 ;
        RECT 128.910 125.025 129.170 125.755 ;
        RECT 129.340 125.200 129.600 125.925 ;
        RECT 129.770 125.025 130.030 125.755 ;
        RECT 130.200 125.200 130.460 125.925 ;
        RECT 130.630 125.025 130.925 125.755 ;
        RECT 131.435 125.195 131.605 125.955 ;
        RECT 131.820 125.025 132.150 125.785 ;
        RECT 132.320 125.195 132.575 126.100 ;
        RECT 132.750 125.025 133.010 126.175 ;
        RECT 133.875 126.115 134.395 126.655 ;
        RECT 134.565 126.335 134.915 126.585 ;
        RECT 135.100 126.165 135.270 126.795 ;
        RECT 135.900 126.925 136.230 127.405 ;
        RECT 136.400 127.115 136.625 127.575 ;
        RECT 136.795 126.925 137.125 127.405 ;
        RECT 135.900 126.755 137.125 126.925 ;
        RECT 137.315 126.775 137.565 127.575 ;
        RECT 137.735 126.775 138.075 127.405 ;
        RECT 138.335 127.025 138.505 127.315 ;
        RECT 138.675 127.195 139.005 127.575 ;
        RECT 138.335 126.855 139.000 127.025 ;
        RECT 135.440 126.385 135.770 126.585 ;
        RECT 135.940 126.385 136.270 126.585 ;
        RECT 136.440 126.385 136.860 126.585 ;
        RECT 137.035 126.415 137.730 126.585 ;
        RECT 137.035 126.165 137.205 126.415 ;
        RECT 137.900 126.165 138.075 126.775 ;
        RECT 133.185 125.025 134.395 126.115 ;
        RECT 134.770 125.995 137.205 126.165 ;
        RECT 134.770 125.195 135.100 125.995 ;
        RECT 135.270 125.025 135.600 125.825 ;
        RECT 135.900 125.195 136.230 125.995 ;
        RECT 136.875 125.025 137.125 125.825 ;
        RECT 137.395 125.025 137.565 126.165 ;
        RECT 137.735 125.195 138.075 126.165 ;
        RECT 138.250 126.035 138.600 126.685 ;
        RECT 138.770 125.865 139.000 126.855 ;
        RECT 138.335 125.695 139.000 125.865 ;
        RECT 138.335 125.195 138.505 125.695 ;
        RECT 138.675 125.025 139.005 125.525 ;
        RECT 139.175 125.195 139.360 127.315 ;
        RECT 139.615 127.115 139.865 127.575 ;
        RECT 140.035 127.125 140.370 127.295 ;
        RECT 140.565 127.125 141.240 127.295 ;
        RECT 140.035 126.985 140.205 127.125 ;
        RECT 139.530 125.995 139.810 126.945 ;
        RECT 139.980 126.855 140.205 126.985 ;
        RECT 139.980 125.750 140.150 126.855 ;
        RECT 140.375 126.705 140.900 126.925 ;
        RECT 140.320 125.940 140.560 126.535 ;
        RECT 140.730 126.005 140.900 126.705 ;
        RECT 141.070 126.345 141.240 127.125 ;
        RECT 141.560 127.075 141.930 127.575 ;
        RECT 142.110 127.125 142.515 127.295 ;
        RECT 142.685 127.125 143.470 127.295 ;
        RECT 142.110 126.895 142.280 127.125 ;
        RECT 141.450 126.595 142.280 126.895 ;
        RECT 142.665 126.625 143.130 126.955 ;
        RECT 141.450 126.565 141.650 126.595 ;
        RECT 141.770 126.345 141.940 126.415 ;
        RECT 141.070 126.175 141.940 126.345 ;
        RECT 141.430 126.085 141.940 126.175 ;
        RECT 139.980 125.620 140.285 125.750 ;
        RECT 140.730 125.640 141.260 126.005 ;
        RECT 139.600 125.025 139.865 125.485 ;
        RECT 140.035 125.195 140.285 125.620 ;
        RECT 141.430 125.470 141.600 126.085 ;
        RECT 140.495 125.300 141.600 125.470 ;
        RECT 141.770 125.025 141.940 125.825 ;
        RECT 142.110 125.525 142.280 126.595 ;
        RECT 142.450 125.695 142.640 126.415 ;
        RECT 142.810 125.665 143.130 126.625 ;
        RECT 143.300 126.665 143.470 127.125 ;
        RECT 143.745 127.045 143.955 127.575 ;
        RECT 144.215 126.835 144.545 127.360 ;
        RECT 144.715 126.965 144.885 127.575 ;
        RECT 145.055 126.920 145.385 127.355 ;
        RECT 146.585 127.115 146.830 127.575 ;
        RECT 145.055 126.835 145.435 126.920 ;
        RECT 144.345 126.665 144.545 126.835 ;
        RECT 145.210 126.795 145.435 126.835 ;
        RECT 143.300 126.335 144.175 126.665 ;
        RECT 144.345 126.335 145.095 126.665 ;
        RECT 142.110 125.195 142.360 125.525 ;
        RECT 143.300 125.495 143.470 126.335 ;
        RECT 144.345 126.130 144.535 126.335 ;
        RECT 145.265 126.215 145.435 126.795 ;
        RECT 146.525 126.335 146.840 126.945 ;
        RECT 147.010 126.585 147.260 127.395 ;
        RECT 147.430 127.050 147.690 127.575 ;
        RECT 147.860 126.925 148.120 127.380 ;
        RECT 148.290 127.095 148.550 127.575 ;
        RECT 148.720 126.925 148.980 127.380 ;
        RECT 149.150 127.095 149.410 127.575 ;
        RECT 149.580 126.925 149.840 127.380 ;
        RECT 150.010 127.095 150.270 127.575 ;
        RECT 150.440 126.925 150.700 127.380 ;
        RECT 150.870 127.095 151.170 127.575 ;
        RECT 147.860 126.755 151.170 126.925 ;
        RECT 151.585 126.850 151.875 127.575 ;
        RECT 147.010 126.335 150.030 126.585 ;
        RECT 145.220 126.165 145.435 126.215 ;
        RECT 143.640 125.755 144.535 126.130 ;
        RECT 145.045 126.085 145.435 126.165 ;
        RECT 142.585 125.325 143.470 125.495 ;
        RECT 143.650 125.025 143.965 125.525 ;
        RECT 144.195 125.195 144.535 125.755 ;
        RECT 144.705 125.025 144.875 126.035 ;
        RECT 145.045 125.240 145.375 126.085 ;
        RECT 146.535 125.025 146.830 126.135 ;
        RECT 147.010 125.200 147.260 126.335 ;
        RECT 150.200 126.165 151.170 126.755 ;
        RECT 152.045 126.775 152.385 127.405 ;
        RECT 152.555 126.775 152.805 127.575 ;
        RECT 152.995 126.925 153.325 127.405 ;
        RECT 153.495 127.115 153.720 127.575 ;
        RECT 153.890 126.925 154.220 127.405 ;
        RECT 147.430 125.025 147.690 126.135 ;
        RECT 147.860 125.925 151.170 126.165 ;
        RECT 147.860 125.200 148.120 125.925 ;
        RECT 148.290 125.025 148.550 125.755 ;
        RECT 148.720 125.200 148.980 125.925 ;
        RECT 149.150 125.025 149.410 125.755 ;
        RECT 149.580 125.200 149.840 125.925 ;
        RECT 150.010 125.025 150.270 125.755 ;
        RECT 150.440 125.200 150.700 125.925 ;
        RECT 150.870 125.025 151.165 125.755 ;
        RECT 151.585 125.025 151.875 126.190 ;
        RECT 152.045 126.165 152.220 126.775 ;
        RECT 152.995 126.755 154.220 126.925 ;
        RECT 154.850 126.795 155.350 127.405 ;
        RECT 155.725 126.825 156.935 127.575 ;
        RECT 152.390 126.415 153.085 126.585 ;
        RECT 152.915 126.165 153.085 126.415 ;
        RECT 153.260 126.385 153.680 126.585 ;
        RECT 153.850 126.385 154.180 126.585 ;
        RECT 154.350 126.385 154.680 126.585 ;
        RECT 154.850 126.165 155.020 126.795 ;
        RECT 155.205 126.335 155.555 126.585 ;
        RECT 152.045 125.195 152.385 126.165 ;
        RECT 152.555 125.025 152.725 126.165 ;
        RECT 152.915 125.995 155.350 126.165 ;
        RECT 152.995 125.025 153.245 125.825 ;
        RECT 153.890 125.195 154.220 125.995 ;
        RECT 154.520 125.025 154.850 125.825 ;
        RECT 155.020 125.195 155.350 125.995 ;
        RECT 155.725 126.115 156.245 126.655 ;
        RECT 156.415 126.285 156.935 126.825 ;
        RECT 155.725 125.025 156.935 126.115 ;
        RECT 22.700 124.855 157.020 125.025 ;
        RECT 22.785 123.765 23.995 124.855 ;
        RECT 24.255 124.185 24.425 124.685 ;
        RECT 24.595 124.355 24.925 124.855 ;
        RECT 24.255 124.015 24.920 124.185 ;
        RECT 22.785 123.055 23.305 123.595 ;
        RECT 23.475 123.225 23.995 123.765 ;
        RECT 24.170 123.195 24.520 123.845 ;
        RECT 22.785 122.305 23.995 123.055 ;
        RECT 24.690 123.025 24.920 124.015 ;
        RECT 24.255 122.855 24.920 123.025 ;
        RECT 24.255 122.565 24.425 122.855 ;
        RECT 24.595 122.305 24.925 122.685 ;
        RECT 25.095 122.565 25.280 124.685 ;
        RECT 25.520 124.395 25.785 124.855 ;
        RECT 25.955 124.260 26.205 124.685 ;
        RECT 26.415 124.410 27.520 124.580 ;
        RECT 25.900 124.130 26.205 124.260 ;
        RECT 25.450 122.935 25.730 123.885 ;
        RECT 25.900 123.025 26.070 124.130 ;
        RECT 26.240 123.345 26.480 123.940 ;
        RECT 26.650 123.875 27.180 124.240 ;
        RECT 26.650 123.175 26.820 123.875 ;
        RECT 27.350 123.795 27.520 124.410 ;
        RECT 27.690 124.055 27.860 124.855 ;
        RECT 28.030 124.355 28.280 124.685 ;
        RECT 28.505 124.385 29.390 124.555 ;
        RECT 27.350 123.705 27.860 123.795 ;
        RECT 25.900 122.895 26.125 123.025 ;
        RECT 26.295 122.955 26.820 123.175 ;
        RECT 26.990 123.535 27.860 123.705 ;
        RECT 25.535 122.305 25.785 122.765 ;
        RECT 25.955 122.755 26.125 122.895 ;
        RECT 26.990 122.755 27.160 123.535 ;
        RECT 27.690 123.465 27.860 123.535 ;
        RECT 27.370 123.285 27.570 123.315 ;
        RECT 28.030 123.285 28.200 124.355 ;
        RECT 28.370 123.465 28.560 124.185 ;
        RECT 27.370 122.985 28.200 123.285 ;
        RECT 28.730 123.255 29.050 124.215 ;
        RECT 25.955 122.585 26.290 122.755 ;
        RECT 26.485 122.585 27.160 122.755 ;
        RECT 27.480 122.305 27.850 122.805 ;
        RECT 28.030 122.755 28.200 122.985 ;
        RECT 28.585 122.925 29.050 123.255 ;
        RECT 29.220 123.545 29.390 124.385 ;
        RECT 29.570 124.355 29.885 124.855 ;
        RECT 30.115 124.125 30.455 124.685 ;
        RECT 29.560 123.750 30.455 124.125 ;
        RECT 30.625 123.845 30.795 124.855 ;
        RECT 30.265 123.545 30.455 123.750 ;
        RECT 30.965 123.795 31.295 124.640 ;
        RECT 30.965 123.715 31.355 123.795 ;
        RECT 31.140 123.665 31.355 123.715 ;
        RECT 29.220 123.215 30.095 123.545 ;
        RECT 30.265 123.215 31.015 123.545 ;
        RECT 29.220 122.755 29.390 123.215 ;
        RECT 30.265 123.045 30.465 123.215 ;
        RECT 31.185 123.085 31.355 123.665 ;
        RECT 31.130 123.045 31.355 123.085 ;
        RECT 28.030 122.585 28.435 122.755 ;
        RECT 28.605 122.585 29.390 122.755 ;
        RECT 29.665 122.305 29.875 122.835 ;
        RECT 30.135 122.520 30.465 123.045 ;
        RECT 30.975 122.960 31.355 123.045 ;
        RECT 31.525 123.715 31.910 124.685 ;
        RECT 32.080 124.395 32.405 124.855 ;
        RECT 32.925 124.225 33.205 124.685 ;
        RECT 32.080 124.005 33.205 124.225 ;
        RECT 31.525 123.045 31.805 123.715 ;
        RECT 32.080 123.545 32.530 124.005 ;
        RECT 33.395 123.835 33.795 124.685 ;
        RECT 34.195 124.395 34.465 124.855 ;
        RECT 34.635 124.225 34.920 124.685 ;
        RECT 31.975 123.215 32.530 123.545 ;
        RECT 32.700 123.275 33.795 123.835 ;
        RECT 32.080 123.105 32.530 123.215 ;
        RECT 30.635 122.305 30.805 122.915 ;
        RECT 30.975 122.525 31.305 122.960 ;
        RECT 31.525 122.475 31.910 123.045 ;
        RECT 32.080 122.935 33.205 123.105 ;
        RECT 32.080 122.305 32.405 122.765 ;
        RECT 32.925 122.475 33.205 122.935 ;
        RECT 33.395 122.475 33.795 123.275 ;
        RECT 33.965 124.005 34.920 124.225 ;
        RECT 33.965 123.105 34.175 124.005 ;
        RECT 34.345 123.275 35.035 123.835 ;
        RECT 35.665 123.690 35.955 124.855 ;
        RECT 36.185 123.795 36.515 124.640 ;
        RECT 36.685 123.845 36.855 124.855 ;
        RECT 37.025 124.125 37.365 124.685 ;
        RECT 37.595 124.355 37.910 124.855 ;
        RECT 38.090 124.385 38.975 124.555 ;
        RECT 36.125 123.715 36.515 123.795 ;
        RECT 37.025 123.750 37.920 124.125 ;
        RECT 36.125 123.665 36.340 123.715 ;
        RECT 33.965 122.935 34.920 123.105 ;
        RECT 36.125 123.085 36.295 123.665 ;
        RECT 37.025 123.545 37.215 123.750 ;
        RECT 38.090 123.545 38.260 124.385 ;
        RECT 39.200 124.355 39.450 124.685 ;
        RECT 36.465 123.215 37.215 123.545 ;
        RECT 37.385 123.215 38.260 123.545 ;
        RECT 36.125 123.045 36.350 123.085 ;
        RECT 37.015 123.045 37.215 123.215 ;
        RECT 34.195 122.305 34.465 122.765 ;
        RECT 34.635 122.475 34.920 122.935 ;
        RECT 35.665 122.305 35.955 123.030 ;
        RECT 36.125 122.960 36.505 123.045 ;
        RECT 36.175 122.525 36.505 122.960 ;
        RECT 36.675 122.305 36.845 122.915 ;
        RECT 37.015 122.520 37.345 123.045 ;
        RECT 37.605 122.305 37.815 122.835 ;
        RECT 38.090 122.755 38.260 123.215 ;
        RECT 38.430 123.255 38.750 124.215 ;
        RECT 38.920 123.465 39.110 124.185 ;
        RECT 39.280 123.285 39.450 124.355 ;
        RECT 39.620 124.055 39.790 124.855 ;
        RECT 39.960 124.410 41.065 124.580 ;
        RECT 39.960 123.795 40.130 124.410 ;
        RECT 41.275 124.260 41.525 124.685 ;
        RECT 41.695 124.395 41.960 124.855 ;
        RECT 40.300 123.875 40.830 124.240 ;
        RECT 41.275 124.130 41.580 124.260 ;
        RECT 39.620 123.705 40.130 123.795 ;
        RECT 39.620 123.535 40.490 123.705 ;
        RECT 39.620 123.465 39.790 123.535 ;
        RECT 39.910 123.285 40.110 123.315 ;
        RECT 38.430 122.925 38.895 123.255 ;
        RECT 39.280 122.985 40.110 123.285 ;
        RECT 39.280 122.755 39.450 122.985 ;
        RECT 38.090 122.585 38.875 122.755 ;
        RECT 39.045 122.585 39.450 122.755 ;
        RECT 39.630 122.305 40.000 122.805 ;
        RECT 40.320 122.755 40.490 123.535 ;
        RECT 40.660 123.175 40.830 123.875 ;
        RECT 41.000 123.345 41.240 123.940 ;
        RECT 40.660 122.955 41.185 123.175 ;
        RECT 41.410 123.025 41.580 124.130 ;
        RECT 41.355 122.895 41.580 123.025 ;
        RECT 41.750 122.935 42.030 123.885 ;
        RECT 41.355 122.755 41.525 122.895 ;
        RECT 40.320 122.585 40.995 122.755 ;
        RECT 41.190 122.585 41.525 122.755 ;
        RECT 41.695 122.305 41.945 122.765 ;
        RECT 42.200 122.565 42.385 124.685 ;
        RECT 42.555 124.355 42.885 124.855 ;
        RECT 43.055 124.185 43.225 124.685 ;
        RECT 42.560 124.015 43.225 124.185 ;
        RECT 44.405 124.135 44.865 124.685 ;
        RECT 45.055 124.135 45.385 124.855 ;
        RECT 42.560 123.025 42.790 124.015 ;
        RECT 42.960 123.195 43.310 123.845 ;
        RECT 42.560 122.855 43.225 123.025 ;
        RECT 42.555 122.305 42.885 122.685 ;
        RECT 43.055 122.565 43.225 122.855 ;
        RECT 44.405 122.765 44.655 124.135 ;
        RECT 45.585 123.965 45.885 124.515 ;
        RECT 46.055 124.185 46.335 124.855 ;
        RECT 46.705 124.420 52.050 124.855 ;
        RECT 44.945 123.795 45.885 123.965 ;
        RECT 44.945 123.545 45.115 123.795 ;
        RECT 46.255 123.545 46.520 123.905 ;
        RECT 44.825 123.215 45.115 123.545 ;
        RECT 45.285 123.295 45.625 123.545 ;
        RECT 45.845 123.295 46.520 123.545 ;
        RECT 44.945 123.125 45.115 123.215 ;
        RECT 44.945 122.935 46.335 123.125 ;
        RECT 44.405 122.475 44.965 122.765 ;
        RECT 45.135 122.305 45.385 122.765 ;
        RECT 46.005 122.575 46.335 122.935 ;
        RECT 48.290 122.850 48.630 123.680 ;
        RECT 50.110 123.170 50.460 124.420 ;
        RECT 52.695 123.885 53.025 124.670 ;
        RECT 52.695 123.715 53.375 123.885 ;
        RECT 53.555 123.715 53.885 124.855 ;
        RECT 54.065 124.420 59.410 124.855 ;
        RECT 52.685 123.295 53.035 123.545 ;
        RECT 53.205 123.115 53.375 123.715 ;
        RECT 53.545 123.295 53.895 123.545 ;
        RECT 46.705 122.305 52.050 122.850 ;
        RECT 52.705 122.305 52.945 123.115 ;
        RECT 53.115 122.475 53.445 123.115 ;
        RECT 53.615 122.305 53.885 123.115 ;
        RECT 55.650 122.850 55.990 123.680 ;
        RECT 57.470 123.170 57.820 124.420 ;
        RECT 59.590 123.705 59.850 124.855 ;
        RECT 60.025 123.780 60.280 124.685 ;
        RECT 60.450 124.095 60.780 124.855 ;
        RECT 60.995 123.925 61.165 124.685 ;
        RECT 54.065 122.305 59.410 122.850 ;
        RECT 59.590 122.305 59.850 123.145 ;
        RECT 60.025 123.050 60.195 123.780 ;
        RECT 60.450 123.755 61.165 123.925 ;
        RECT 60.450 123.545 60.620 123.755 ;
        RECT 61.425 123.690 61.715 124.855 ;
        RECT 61.975 123.925 62.145 124.685 ;
        RECT 62.360 124.095 62.690 124.855 ;
        RECT 61.975 123.755 62.690 123.925 ;
        RECT 62.860 123.780 63.115 124.685 ;
        RECT 60.365 123.215 60.620 123.545 ;
        RECT 60.025 122.475 60.280 123.050 ;
        RECT 60.450 123.025 60.620 123.215 ;
        RECT 60.900 123.205 61.255 123.575 ;
        RECT 61.885 123.205 62.240 123.575 ;
        RECT 62.520 123.545 62.690 123.755 ;
        RECT 62.520 123.215 62.775 123.545 ;
        RECT 60.450 122.855 61.165 123.025 ;
        RECT 60.450 122.305 60.780 122.685 ;
        RECT 60.995 122.475 61.165 122.855 ;
        RECT 61.425 122.305 61.715 123.030 ;
        RECT 62.520 123.025 62.690 123.215 ;
        RECT 62.945 123.050 63.115 123.780 ;
        RECT 63.290 123.705 63.550 124.855 ;
        RECT 63.815 123.925 63.985 124.685 ;
        RECT 64.200 124.095 64.530 124.855 ;
        RECT 63.815 123.755 64.530 123.925 ;
        RECT 64.700 123.780 64.955 124.685 ;
        RECT 63.725 123.205 64.080 123.575 ;
        RECT 64.360 123.545 64.530 123.755 ;
        RECT 64.360 123.215 64.615 123.545 ;
        RECT 61.975 122.855 62.690 123.025 ;
        RECT 61.975 122.475 62.145 122.855 ;
        RECT 62.360 122.305 62.690 122.685 ;
        RECT 62.860 122.475 63.115 123.050 ;
        RECT 63.290 122.305 63.550 123.145 ;
        RECT 64.360 123.025 64.530 123.215 ;
        RECT 64.785 123.050 64.955 123.780 ;
        RECT 65.130 123.705 65.390 124.855 ;
        RECT 65.565 123.765 68.155 124.855 ;
        RECT 68.385 123.795 68.715 124.640 ;
        RECT 68.885 123.845 69.055 124.855 ;
        RECT 69.225 124.125 69.565 124.685 ;
        RECT 69.795 124.355 70.110 124.855 ;
        RECT 70.290 124.385 71.175 124.555 ;
        RECT 63.815 122.855 64.530 123.025 ;
        RECT 63.815 122.475 63.985 122.855 ;
        RECT 64.200 122.305 64.530 122.685 ;
        RECT 64.700 122.475 64.955 123.050 ;
        RECT 65.130 122.305 65.390 123.145 ;
        RECT 65.565 123.075 66.775 123.595 ;
        RECT 66.945 123.245 68.155 123.765 ;
        RECT 68.325 123.715 68.715 123.795 ;
        RECT 69.225 123.750 70.120 124.125 ;
        RECT 68.325 123.665 68.540 123.715 ;
        RECT 68.325 123.085 68.495 123.665 ;
        RECT 69.225 123.545 69.415 123.750 ;
        RECT 70.290 123.545 70.460 124.385 ;
        RECT 71.400 124.355 71.650 124.685 ;
        RECT 68.665 123.215 69.415 123.545 ;
        RECT 69.585 123.215 70.460 123.545 ;
        RECT 65.565 122.305 68.155 123.075 ;
        RECT 68.325 123.045 68.550 123.085 ;
        RECT 69.215 123.045 69.415 123.215 ;
        RECT 68.325 122.960 68.705 123.045 ;
        RECT 68.375 122.525 68.705 122.960 ;
        RECT 68.875 122.305 69.045 122.915 ;
        RECT 69.215 122.520 69.545 123.045 ;
        RECT 69.805 122.305 70.015 122.835 ;
        RECT 70.290 122.755 70.460 123.215 ;
        RECT 70.630 123.255 70.950 124.215 ;
        RECT 71.120 123.465 71.310 124.185 ;
        RECT 71.480 123.285 71.650 124.355 ;
        RECT 71.820 124.055 71.990 124.855 ;
        RECT 72.160 124.410 73.265 124.580 ;
        RECT 72.160 123.795 72.330 124.410 ;
        RECT 73.475 124.260 73.725 124.685 ;
        RECT 73.895 124.395 74.160 124.855 ;
        RECT 72.500 123.875 73.030 124.240 ;
        RECT 73.475 124.130 73.780 124.260 ;
        RECT 71.820 123.705 72.330 123.795 ;
        RECT 71.820 123.535 72.690 123.705 ;
        RECT 71.820 123.465 71.990 123.535 ;
        RECT 72.110 123.285 72.310 123.315 ;
        RECT 70.630 122.925 71.095 123.255 ;
        RECT 71.480 122.985 72.310 123.285 ;
        RECT 71.480 122.755 71.650 122.985 ;
        RECT 70.290 122.585 71.075 122.755 ;
        RECT 71.245 122.585 71.650 122.755 ;
        RECT 71.830 122.305 72.200 122.805 ;
        RECT 72.520 122.755 72.690 123.535 ;
        RECT 72.860 123.175 73.030 123.875 ;
        RECT 73.200 123.345 73.440 123.940 ;
        RECT 72.860 122.955 73.385 123.175 ;
        RECT 73.610 123.025 73.780 124.130 ;
        RECT 73.555 122.895 73.780 123.025 ;
        RECT 73.950 122.935 74.230 123.885 ;
        RECT 73.555 122.755 73.725 122.895 ;
        RECT 72.520 122.585 73.195 122.755 ;
        RECT 73.390 122.585 73.725 122.755 ;
        RECT 73.895 122.305 74.145 122.765 ;
        RECT 74.400 122.565 74.585 124.685 ;
        RECT 74.755 124.355 75.085 124.855 ;
        RECT 75.255 124.185 75.425 124.685 ;
        RECT 74.760 124.015 75.425 124.185 ;
        RECT 75.720 124.065 76.255 124.685 ;
        RECT 74.760 123.025 74.990 124.015 ;
        RECT 75.160 123.195 75.510 123.845 ;
        RECT 75.720 123.045 76.035 124.065 ;
        RECT 76.425 124.055 76.755 124.855 ;
        RECT 77.240 123.885 77.630 124.060 ;
        RECT 76.205 123.715 77.630 123.885 ;
        RECT 77.985 123.765 80.575 124.855 ;
        RECT 76.205 123.215 76.375 123.715 ;
        RECT 74.760 122.855 75.425 123.025 ;
        RECT 74.755 122.305 75.085 122.685 ;
        RECT 75.255 122.565 75.425 122.855 ;
        RECT 75.720 122.475 76.335 123.045 ;
        RECT 76.625 122.985 76.890 123.545 ;
        RECT 77.060 122.815 77.230 123.715 ;
        RECT 77.400 122.985 77.755 123.545 ;
        RECT 77.985 123.075 79.195 123.595 ;
        RECT 79.365 123.245 80.575 123.765 ;
        RECT 76.505 122.305 76.720 122.815 ;
        RECT 76.950 122.485 77.230 122.815 ;
        RECT 77.410 122.305 77.650 122.815 ;
        RECT 77.985 122.305 80.575 123.075 ;
        RECT 80.755 122.485 81.015 124.675 ;
        RECT 81.185 124.125 81.525 124.855 ;
        RECT 81.705 123.945 81.975 124.675 ;
        RECT 81.205 123.725 81.975 123.945 ;
        RECT 82.155 123.965 82.385 124.675 ;
        RECT 82.555 124.145 82.885 124.855 ;
        RECT 83.055 123.965 83.315 124.675 ;
        RECT 82.155 123.725 83.315 123.965 ;
        RECT 83.505 123.985 83.780 124.685 ;
        RECT 83.950 124.310 84.205 124.855 ;
        RECT 84.375 124.345 84.855 124.685 ;
        RECT 85.030 124.300 85.635 124.855 ;
        RECT 85.020 124.200 85.635 124.300 ;
        RECT 85.020 124.175 85.205 124.200 ;
        RECT 81.205 123.055 81.495 123.725 ;
        RECT 81.675 123.235 82.140 123.545 ;
        RECT 82.320 123.235 82.845 123.545 ;
        RECT 81.205 122.855 82.435 123.055 ;
        RECT 81.275 122.305 81.945 122.675 ;
        RECT 82.125 122.485 82.435 122.855 ;
        RECT 82.615 122.595 82.845 123.235 ;
        RECT 83.025 123.215 83.325 123.545 ;
        RECT 83.025 122.305 83.315 123.035 ;
        RECT 83.505 122.955 83.675 123.985 ;
        RECT 83.950 123.855 84.705 124.105 ;
        RECT 84.875 123.930 85.205 124.175 ;
        RECT 83.950 123.820 84.720 123.855 ;
        RECT 83.950 123.810 84.735 123.820 ;
        RECT 83.845 123.795 84.740 123.810 ;
        RECT 83.845 123.780 84.760 123.795 ;
        RECT 83.845 123.770 84.780 123.780 ;
        RECT 83.845 123.760 84.805 123.770 ;
        RECT 83.845 123.730 84.875 123.760 ;
        RECT 83.845 123.700 84.895 123.730 ;
        RECT 83.845 123.670 84.915 123.700 ;
        RECT 83.845 123.645 84.945 123.670 ;
        RECT 83.845 123.610 84.980 123.645 ;
        RECT 83.845 123.605 85.010 123.610 ;
        RECT 83.845 123.210 84.075 123.605 ;
        RECT 84.620 123.600 85.010 123.605 ;
        RECT 84.645 123.590 85.010 123.600 ;
        RECT 84.660 123.585 85.010 123.590 ;
        RECT 84.675 123.580 85.010 123.585 ;
        RECT 85.375 123.580 85.635 124.030 ;
        RECT 85.815 123.715 86.145 124.855 ;
        RECT 86.675 123.885 87.005 124.670 ;
        RECT 86.325 123.715 87.005 123.885 ;
        RECT 84.675 123.575 85.635 123.580 ;
        RECT 84.685 123.565 85.635 123.575 ;
        RECT 84.695 123.560 85.635 123.565 ;
        RECT 84.705 123.550 85.635 123.560 ;
        RECT 84.710 123.540 85.635 123.550 ;
        RECT 84.715 123.535 85.635 123.540 ;
        RECT 84.725 123.520 85.635 123.535 ;
        RECT 84.730 123.505 85.635 123.520 ;
        RECT 84.740 123.480 85.635 123.505 ;
        RECT 84.245 123.010 84.575 123.435 ;
        RECT 83.505 122.475 83.765 122.955 ;
        RECT 83.935 122.305 84.185 122.845 ;
        RECT 84.355 122.525 84.575 123.010 ;
        RECT 84.745 123.410 85.635 123.480 ;
        RECT 84.745 122.685 84.915 123.410 ;
        RECT 85.805 123.295 86.155 123.545 ;
        RECT 85.085 122.855 85.635 123.240 ;
        RECT 86.325 123.115 86.495 123.715 ;
        RECT 87.185 123.690 87.475 124.855 ;
        RECT 88.575 123.745 88.870 124.855 ;
        RECT 89.050 123.545 89.300 124.680 ;
        RECT 89.470 123.745 89.730 124.855 ;
        RECT 89.900 123.955 90.160 124.680 ;
        RECT 90.330 124.125 90.590 124.855 ;
        RECT 90.760 123.955 91.020 124.680 ;
        RECT 91.190 124.125 91.450 124.855 ;
        RECT 91.620 123.955 91.880 124.680 ;
        RECT 92.050 124.125 92.310 124.855 ;
        RECT 92.480 123.955 92.740 124.680 ;
        RECT 92.910 124.125 93.205 124.855 ;
        RECT 89.900 123.715 93.210 123.955 ;
        RECT 86.665 123.295 87.015 123.545 ;
        RECT 84.745 122.515 85.635 122.685 ;
        RECT 85.815 122.305 86.085 123.115 ;
        RECT 86.255 122.475 86.585 123.115 ;
        RECT 86.755 122.305 86.995 123.115 ;
        RECT 87.185 122.305 87.475 123.030 ;
        RECT 88.565 122.935 88.880 123.545 ;
        RECT 89.050 123.295 92.070 123.545 ;
        RECT 88.625 122.305 88.870 122.765 ;
        RECT 89.050 122.485 89.300 123.295 ;
        RECT 92.240 123.125 93.210 123.715 ;
        RECT 89.900 122.955 93.210 123.125 ;
        RECT 89.470 122.305 89.730 122.830 ;
        RECT 89.900 122.500 90.160 122.955 ;
        RECT 90.330 122.305 90.590 122.785 ;
        RECT 90.760 122.500 91.020 122.955 ;
        RECT 91.190 122.305 91.450 122.785 ;
        RECT 91.620 122.500 91.880 122.955 ;
        RECT 92.050 122.305 92.310 122.785 ;
        RECT 92.480 122.500 92.740 122.955 ;
        RECT 92.910 122.305 93.210 122.785 ;
        RECT 93.635 122.485 93.895 124.675 ;
        RECT 94.065 124.125 94.405 124.855 ;
        RECT 94.585 123.945 94.855 124.675 ;
        RECT 94.085 123.725 94.855 123.945 ;
        RECT 95.035 123.965 95.265 124.675 ;
        RECT 95.435 124.145 95.765 124.855 ;
        RECT 95.935 123.965 96.195 124.675 ;
        RECT 95.035 123.725 96.195 123.965 ;
        RECT 96.385 123.985 96.660 124.685 ;
        RECT 96.830 124.310 97.085 124.855 ;
        RECT 97.255 124.345 97.735 124.685 ;
        RECT 97.910 124.300 98.515 124.855 ;
        RECT 97.900 124.200 98.515 124.300 ;
        RECT 97.900 124.175 98.085 124.200 ;
        RECT 94.085 123.055 94.375 123.725 ;
        RECT 94.555 123.235 95.020 123.545 ;
        RECT 95.200 123.235 95.725 123.545 ;
        RECT 94.085 122.855 95.315 123.055 ;
        RECT 94.155 122.305 94.825 122.675 ;
        RECT 95.005 122.485 95.315 122.855 ;
        RECT 95.495 122.595 95.725 123.235 ;
        RECT 95.905 123.215 96.205 123.545 ;
        RECT 95.905 122.305 96.195 123.035 ;
        RECT 96.385 122.955 96.555 123.985 ;
        RECT 96.830 123.855 97.585 124.105 ;
        RECT 97.755 123.930 98.085 124.175 ;
        RECT 96.830 123.820 97.600 123.855 ;
        RECT 96.830 123.810 97.615 123.820 ;
        RECT 96.725 123.795 97.620 123.810 ;
        RECT 96.725 123.780 97.640 123.795 ;
        RECT 96.725 123.770 97.660 123.780 ;
        RECT 96.725 123.760 97.685 123.770 ;
        RECT 96.725 123.730 97.755 123.760 ;
        RECT 96.725 123.700 97.775 123.730 ;
        RECT 96.725 123.670 97.795 123.700 ;
        RECT 96.725 123.645 97.825 123.670 ;
        RECT 96.725 123.610 97.860 123.645 ;
        RECT 96.725 123.605 97.890 123.610 ;
        RECT 96.725 123.210 96.955 123.605 ;
        RECT 97.500 123.600 97.890 123.605 ;
        RECT 97.525 123.590 97.890 123.600 ;
        RECT 97.540 123.585 97.890 123.590 ;
        RECT 97.555 123.580 97.890 123.585 ;
        RECT 98.255 123.580 98.515 124.030 ;
        RECT 98.685 123.765 100.355 124.855 ;
        RECT 97.555 123.575 98.515 123.580 ;
        RECT 97.565 123.565 98.515 123.575 ;
        RECT 97.575 123.560 98.515 123.565 ;
        RECT 97.585 123.550 98.515 123.560 ;
        RECT 97.590 123.540 98.515 123.550 ;
        RECT 97.595 123.535 98.515 123.540 ;
        RECT 97.605 123.520 98.515 123.535 ;
        RECT 97.610 123.505 98.515 123.520 ;
        RECT 97.620 123.480 98.515 123.505 ;
        RECT 97.125 123.010 97.455 123.435 ;
        RECT 96.385 122.475 96.645 122.955 ;
        RECT 96.815 122.305 97.065 122.845 ;
        RECT 97.235 122.525 97.455 123.010 ;
        RECT 97.625 123.410 98.515 123.480 ;
        RECT 97.625 122.685 97.795 123.410 ;
        RECT 97.965 122.855 98.515 123.240 ;
        RECT 98.685 123.075 99.435 123.595 ;
        RECT 99.605 123.245 100.355 123.765 ;
        RECT 100.985 123.715 101.370 124.685 ;
        RECT 101.540 124.395 101.865 124.855 ;
        RECT 102.385 124.225 102.665 124.685 ;
        RECT 101.540 124.005 102.665 124.225 ;
        RECT 97.625 122.515 98.515 122.685 ;
        RECT 98.685 122.305 100.355 123.075 ;
        RECT 100.985 123.045 101.265 123.715 ;
        RECT 101.540 123.545 101.990 124.005 ;
        RECT 102.855 123.835 103.255 124.685 ;
        RECT 103.655 124.395 103.925 124.855 ;
        RECT 104.095 124.225 104.380 124.685 ;
        RECT 101.435 123.215 101.990 123.545 ;
        RECT 102.160 123.275 103.255 123.835 ;
        RECT 101.540 123.105 101.990 123.215 ;
        RECT 100.985 122.475 101.370 123.045 ;
        RECT 101.540 122.935 102.665 123.105 ;
        RECT 101.540 122.305 101.865 122.765 ;
        RECT 102.385 122.475 102.665 122.935 ;
        RECT 102.855 122.475 103.255 123.275 ;
        RECT 103.425 124.005 104.380 124.225 ;
        RECT 103.425 123.105 103.635 124.005 ;
        RECT 103.805 123.275 104.495 123.835 ;
        RECT 103.425 122.935 104.380 123.105 ;
        RECT 103.655 122.305 103.925 122.765 ;
        RECT 104.095 122.475 104.380 122.935 ;
        RECT 104.675 122.485 104.935 124.675 ;
        RECT 105.105 124.125 105.445 124.855 ;
        RECT 105.625 123.945 105.895 124.675 ;
        RECT 105.125 123.725 105.895 123.945 ;
        RECT 106.075 123.965 106.305 124.675 ;
        RECT 106.475 124.145 106.805 124.855 ;
        RECT 106.975 123.965 107.235 124.675 ;
        RECT 106.075 123.725 107.235 123.965 ;
        RECT 107.425 123.765 110.015 124.855 ;
        RECT 105.125 123.055 105.415 123.725 ;
        RECT 105.595 123.235 106.060 123.545 ;
        RECT 106.240 123.235 106.765 123.545 ;
        RECT 105.125 122.855 106.355 123.055 ;
        RECT 105.195 122.305 105.865 122.675 ;
        RECT 106.045 122.485 106.355 122.855 ;
        RECT 106.535 122.595 106.765 123.235 ;
        RECT 106.945 123.215 107.245 123.545 ;
        RECT 107.425 123.075 108.635 123.595 ;
        RECT 108.805 123.245 110.015 123.765 ;
        RECT 106.945 122.305 107.235 123.035 ;
        RECT 107.425 122.305 110.015 123.075 ;
        RECT 110.195 122.485 110.455 124.675 ;
        RECT 110.625 124.125 110.965 124.855 ;
        RECT 111.145 123.945 111.415 124.675 ;
        RECT 110.645 123.725 111.415 123.945 ;
        RECT 111.595 123.965 111.825 124.675 ;
        RECT 111.995 124.145 112.325 124.855 ;
        RECT 112.495 123.965 112.755 124.675 ;
        RECT 111.595 123.725 112.755 123.965 ;
        RECT 110.645 123.055 110.935 123.725 ;
        RECT 112.945 123.690 113.235 124.855 ;
        RECT 113.520 124.225 113.805 124.685 ;
        RECT 113.975 124.395 114.245 124.855 ;
        RECT 113.520 124.005 114.475 124.225 ;
        RECT 111.115 123.235 111.580 123.545 ;
        RECT 111.760 123.235 112.285 123.545 ;
        RECT 110.645 122.855 111.875 123.055 ;
        RECT 110.715 122.305 111.385 122.675 ;
        RECT 111.565 122.485 111.875 122.855 ;
        RECT 112.055 122.595 112.285 123.235 ;
        RECT 112.465 123.215 112.765 123.545 ;
        RECT 113.405 123.275 114.095 123.835 ;
        RECT 114.265 123.105 114.475 124.005 ;
        RECT 112.465 122.305 112.755 123.035 ;
        RECT 112.945 122.305 113.235 123.030 ;
        RECT 113.520 122.935 114.475 123.105 ;
        RECT 114.645 123.835 115.045 124.685 ;
        RECT 115.235 124.225 115.515 124.685 ;
        RECT 116.035 124.395 116.360 124.855 ;
        RECT 115.235 124.005 116.360 124.225 ;
        RECT 114.645 123.275 115.740 123.835 ;
        RECT 115.910 123.545 116.360 124.005 ;
        RECT 116.530 123.715 116.915 124.685 ;
        RECT 113.520 122.475 113.805 122.935 ;
        RECT 113.975 122.305 114.245 122.765 ;
        RECT 114.645 122.475 115.045 123.275 ;
        RECT 115.910 123.215 116.465 123.545 ;
        RECT 115.910 123.105 116.360 123.215 ;
        RECT 115.235 122.935 116.360 123.105 ;
        RECT 116.635 123.045 116.915 123.715 ;
        RECT 115.235 122.475 115.515 122.935 ;
        RECT 116.035 122.305 116.360 122.765 ;
        RECT 116.530 122.475 116.915 123.045 ;
        RECT 117.085 123.985 117.360 124.685 ;
        RECT 117.530 124.310 117.785 124.855 ;
        RECT 117.955 124.345 118.435 124.685 ;
        RECT 118.610 124.300 119.215 124.855 ;
        RECT 118.600 124.200 119.215 124.300 ;
        RECT 118.600 124.175 118.785 124.200 ;
        RECT 117.085 122.955 117.255 123.985 ;
        RECT 117.530 123.855 118.285 124.105 ;
        RECT 118.455 123.930 118.785 124.175 ;
        RECT 117.530 123.820 118.300 123.855 ;
        RECT 117.530 123.810 118.315 123.820 ;
        RECT 117.425 123.795 118.320 123.810 ;
        RECT 117.425 123.780 118.340 123.795 ;
        RECT 117.425 123.770 118.360 123.780 ;
        RECT 117.425 123.760 118.385 123.770 ;
        RECT 117.425 123.730 118.455 123.760 ;
        RECT 117.425 123.700 118.475 123.730 ;
        RECT 117.425 123.670 118.495 123.700 ;
        RECT 117.425 123.645 118.525 123.670 ;
        RECT 117.425 123.610 118.560 123.645 ;
        RECT 117.425 123.605 118.590 123.610 ;
        RECT 117.425 123.210 117.655 123.605 ;
        RECT 118.200 123.600 118.590 123.605 ;
        RECT 118.225 123.590 118.590 123.600 ;
        RECT 118.240 123.585 118.590 123.590 ;
        RECT 118.255 123.580 118.590 123.585 ;
        RECT 118.955 123.580 119.215 124.030 ;
        RECT 119.845 123.715 120.105 124.855 ;
        RECT 120.345 124.345 121.960 124.675 ;
        RECT 118.255 123.575 119.215 123.580 ;
        RECT 118.265 123.565 119.215 123.575 ;
        RECT 118.275 123.560 119.215 123.565 ;
        RECT 118.285 123.550 119.215 123.560 ;
        RECT 118.290 123.540 119.215 123.550 ;
        RECT 120.355 123.545 120.525 124.105 ;
        RECT 120.785 124.005 121.960 124.175 ;
        RECT 122.130 124.055 122.410 124.855 ;
        RECT 120.785 123.715 121.115 124.005 ;
        RECT 121.790 123.885 121.960 124.005 ;
        RECT 121.285 123.545 121.530 123.835 ;
        RECT 121.790 123.715 122.450 123.885 ;
        RECT 122.620 123.715 122.895 124.685 ;
        RECT 122.280 123.545 122.450 123.715 ;
        RECT 118.295 123.535 119.215 123.540 ;
        RECT 118.305 123.520 119.215 123.535 ;
        RECT 118.310 123.505 119.215 123.520 ;
        RECT 118.320 123.480 119.215 123.505 ;
        RECT 117.825 123.010 118.155 123.435 ;
        RECT 117.085 122.475 117.345 122.955 ;
        RECT 117.515 122.305 117.765 122.845 ;
        RECT 117.935 122.525 118.155 123.010 ;
        RECT 118.325 123.410 119.215 123.480 ;
        RECT 118.325 122.685 118.495 123.410 ;
        RECT 119.850 123.295 120.185 123.545 ;
        RECT 118.665 122.855 119.215 123.240 ;
        RECT 120.355 123.215 121.070 123.545 ;
        RECT 121.285 123.215 122.110 123.545 ;
        RECT 122.280 123.215 122.555 123.545 ;
        RECT 120.355 123.125 120.605 123.215 ;
        RECT 118.325 122.515 119.215 122.685 ;
        RECT 119.845 122.305 120.105 123.125 ;
        RECT 120.275 122.705 120.605 123.125 ;
        RECT 122.280 123.045 122.450 123.215 ;
        RECT 120.785 122.875 122.450 123.045 ;
        RECT 122.725 122.980 122.895 123.715 ;
        RECT 123.070 123.705 123.330 124.855 ;
        RECT 123.505 123.780 123.760 124.685 ;
        RECT 123.930 124.095 124.260 124.855 ;
        RECT 124.475 123.925 124.645 124.685 ;
        RECT 120.785 122.475 121.045 122.875 ;
        RECT 121.215 122.305 121.545 122.705 ;
        RECT 121.715 122.525 121.885 122.875 ;
        RECT 122.055 122.305 122.430 122.705 ;
        RECT 122.620 122.635 122.895 122.980 ;
        RECT 123.070 122.305 123.330 123.145 ;
        RECT 123.505 123.050 123.675 123.780 ;
        RECT 123.930 123.755 124.645 123.925 ;
        RECT 124.905 123.765 126.115 124.855 ;
        RECT 126.375 124.235 126.545 124.665 ;
        RECT 126.715 124.405 127.045 124.855 ;
        RECT 126.375 124.005 127.050 124.235 ;
        RECT 123.930 123.545 124.100 123.755 ;
        RECT 123.845 123.215 124.100 123.545 ;
        RECT 123.505 122.475 123.760 123.050 ;
        RECT 123.930 123.025 124.100 123.215 ;
        RECT 124.380 123.205 124.735 123.575 ;
        RECT 124.905 123.055 125.425 123.595 ;
        RECT 125.595 123.225 126.115 123.765 ;
        RECT 123.930 122.855 124.645 123.025 ;
        RECT 123.930 122.305 124.260 122.685 ;
        RECT 124.475 122.475 124.645 122.855 ;
        RECT 124.905 122.305 126.115 123.055 ;
        RECT 126.345 122.985 126.645 123.835 ;
        RECT 126.815 123.355 127.050 124.005 ;
        RECT 127.220 123.695 127.505 124.640 ;
        RECT 127.685 124.385 128.370 124.855 ;
        RECT 127.680 123.865 128.375 124.175 ;
        RECT 128.550 123.800 128.855 124.585 ;
        RECT 129.135 124.185 129.305 124.685 ;
        RECT 129.475 124.355 129.805 124.855 ;
        RECT 129.135 124.015 129.800 124.185 ;
        RECT 127.220 123.545 128.080 123.695 ;
        RECT 127.220 123.525 128.505 123.545 ;
        RECT 126.815 123.025 127.350 123.355 ;
        RECT 127.520 123.165 128.505 123.525 ;
        RECT 126.815 122.875 127.035 123.025 ;
        RECT 126.290 122.305 126.625 122.810 ;
        RECT 126.795 122.500 127.035 122.875 ;
        RECT 127.520 122.830 127.690 123.165 ;
        RECT 128.680 122.995 128.855 123.800 ;
        RECT 129.050 123.195 129.400 123.845 ;
        RECT 129.570 123.025 129.800 124.015 ;
        RECT 127.315 122.635 127.690 122.830 ;
        RECT 127.315 122.490 127.485 122.635 ;
        RECT 128.050 122.305 128.445 122.800 ;
        RECT 128.615 122.475 128.855 122.995 ;
        RECT 129.135 122.855 129.800 123.025 ;
        RECT 129.135 122.565 129.305 122.855 ;
        RECT 129.475 122.305 129.805 122.685 ;
        RECT 129.975 122.565 130.160 124.685 ;
        RECT 130.400 124.395 130.665 124.855 ;
        RECT 130.835 124.260 131.085 124.685 ;
        RECT 131.295 124.410 132.400 124.580 ;
        RECT 130.780 124.130 131.085 124.260 ;
        RECT 130.330 122.935 130.610 123.885 ;
        RECT 130.780 123.025 130.950 124.130 ;
        RECT 131.120 123.345 131.360 123.940 ;
        RECT 131.530 123.875 132.060 124.240 ;
        RECT 131.530 123.175 131.700 123.875 ;
        RECT 132.230 123.795 132.400 124.410 ;
        RECT 132.570 124.055 132.740 124.855 ;
        RECT 132.910 124.355 133.160 124.685 ;
        RECT 133.385 124.385 134.270 124.555 ;
        RECT 132.230 123.705 132.740 123.795 ;
        RECT 130.780 122.895 131.005 123.025 ;
        RECT 131.175 122.955 131.700 123.175 ;
        RECT 131.870 123.535 132.740 123.705 ;
        RECT 130.415 122.305 130.665 122.765 ;
        RECT 130.835 122.755 131.005 122.895 ;
        RECT 131.870 122.755 132.040 123.535 ;
        RECT 132.570 123.465 132.740 123.535 ;
        RECT 132.250 123.285 132.450 123.315 ;
        RECT 132.910 123.285 133.080 124.355 ;
        RECT 133.250 123.465 133.440 124.185 ;
        RECT 132.250 122.985 133.080 123.285 ;
        RECT 133.610 123.255 133.930 124.215 ;
        RECT 130.835 122.585 131.170 122.755 ;
        RECT 131.365 122.585 132.040 122.755 ;
        RECT 132.360 122.305 132.730 122.805 ;
        RECT 132.910 122.755 133.080 122.985 ;
        RECT 133.465 122.925 133.930 123.255 ;
        RECT 134.100 123.545 134.270 124.385 ;
        RECT 134.450 124.355 134.765 124.855 ;
        RECT 134.995 124.125 135.335 124.685 ;
        RECT 134.440 123.750 135.335 124.125 ;
        RECT 135.505 123.845 135.675 124.855 ;
        RECT 135.145 123.545 135.335 123.750 ;
        RECT 135.845 123.795 136.175 124.640 ;
        RECT 136.440 124.065 136.975 124.685 ;
        RECT 135.845 123.715 136.235 123.795 ;
        RECT 136.020 123.665 136.235 123.715 ;
        RECT 134.100 123.215 134.975 123.545 ;
        RECT 135.145 123.215 135.895 123.545 ;
        RECT 134.100 122.755 134.270 123.215 ;
        RECT 135.145 123.045 135.345 123.215 ;
        RECT 136.065 123.085 136.235 123.665 ;
        RECT 136.010 123.045 136.235 123.085 ;
        RECT 132.910 122.585 133.315 122.755 ;
        RECT 133.485 122.585 134.270 122.755 ;
        RECT 134.545 122.305 134.755 122.835 ;
        RECT 135.015 122.520 135.345 123.045 ;
        RECT 135.855 122.960 136.235 123.045 ;
        RECT 136.440 123.045 136.755 124.065 ;
        RECT 137.145 124.055 137.475 124.855 ;
        RECT 137.960 123.885 138.350 124.060 ;
        RECT 136.925 123.715 138.350 123.885 ;
        RECT 136.925 123.215 137.095 123.715 ;
        RECT 135.515 122.305 135.685 122.915 ;
        RECT 135.855 122.525 136.185 122.960 ;
        RECT 136.440 122.475 137.055 123.045 ;
        RECT 137.345 122.985 137.610 123.545 ;
        RECT 137.780 122.815 137.950 123.715 ;
        RECT 138.705 123.690 138.995 124.855 ;
        RECT 139.165 123.715 139.550 124.685 ;
        RECT 139.720 124.395 140.045 124.855 ;
        RECT 140.565 124.225 140.845 124.685 ;
        RECT 139.720 124.005 140.845 124.225 ;
        RECT 138.120 122.985 138.475 123.545 ;
        RECT 139.165 123.045 139.445 123.715 ;
        RECT 139.720 123.545 140.170 124.005 ;
        RECT 141.035 123.835 141.435 124.685 ;
        RECT 141.835 124.395 142.105 124.855 ;
        RECT 142.275 124.225 142.560 124.685 ;
        RECT 139.615 123.215 140.170 123.545 ;
        RECT 140.340 123.275 141.435 123.835 ;
        RECT 139.720 123.105 140.170 123.215 ;
        RECT 137.225 122.305 137.440 122.815 ;
        RECT 137.670 122.485 137.950 122.815 ;
        RECT 138.130 122.305 138.370 122.815 ;
        RECT 138.705 122.305 138.995 123.030 ;
        RECT 139.165 122.475 139.550 123.045 ;
        RECT 139.720 122.935 140.845 123.105 ;
        RECT 139.720 122.305 140.045 122.765 ;
        RECT 140.565 122.475 140.845 122.935 ;
        RECT 141.035 122.475 141.435 123.275 ;
        RECT 141.605 124.005 142.560 124.225 ;
        RECT 141.605 123.105 141.815 124.005 ;
        RECT 141.985 123.275 142.675 123.835 ;
        RECT 142.845 123.715 143.115 124.685 ;
        RECT 143.325 124.055 143.605 124.855 ;
        RECT 143.775 124.345 145.430 124.635 ;
        RECT 143.840 124.005 145.430 124.175 ;
        RECT 143.840 123.885 144.010 124.005 ;
        RECT 143.285 123.715 144.010 123.885 ;
        RECT 141.605 122.935 142.560 123.105 ;
        RECT 141.835 122.305 142.105 122.765 ;
        RECT 142.275 122.475 142.560 122.935 ;
        RECT 142.845 122.980 143.015 123.715 ;
        RECT 143.285 123.545 143.455 123.715 ;
        RECT 143.185 123.215 143.455 123.545 ;
        RECT 143.625 123.215 144.030 123.545 ;
        RECT 144.200 123.215 144.910 123.835 ;
        RECT 145.110 123.715 145.430 124.005 ;
        RECT 145.605 123.765 147.275 124.855 ;
        RECT 147.535 124.185 147.705 124.685 ;
        RECT 147.875 124.355 148.205 124.855 ;
        RECT 147.535 124.015 148.200 124.185 ;
        RECT 143.285 123.045 143.455 123.215 ;
        RECT 142.845 122.635 143.115 122.980 ;
        RECT 143.285 122.875 144.895 123.045 ;
        RECT 145.080 122.975 145.430 123.545 ;
        RECT 145.605 123.075 146.355 123.595 ;
        RECT 146.525 123.245 147.275 123.765 ;
        RECT 147.450 123.195 147.800 123.845 ;
        RECT 143.305 122.305 143.685 122.705 ;
        RECT 143.855 122.525 144.025 122.875 ;
        RECT 144.195 122.305 144.525 122.705 ;
        RECT 144.725 122.525 144.895 122.875 ;
        RECT 145.095 122.305 145.425 122.805 ;
        RECT 145.605 122.305 147.275 123.075 ;
        RECT 147.970 123.025 148.200 124.015 ;
        RECT 147.535 122.855 148.200 123.025 ;
        RECT 147.535 122.565 147.705 122.855 ;
        RECT 147.875 122.305 148.205 122.685 ;
        RECT 148.375 122.565 148.560 124.685 ;
        RECT 148.800 124.395 149.065 124.855 ;
        RECT 149.235 124.260 149.485 124.685 ;
        RECT 149.695 124.410 150.800 124.580 ;
        RECT 149.180 124.130 149.485 124.260 ;
        RECT 148.730 122.935 149.010 123.885 ;
        RECT 149.180 123.025 149.350 124.130 ;
        RECT 149.520 123.345 149.760 123.940 ;
        RECT 149.930 123.875 150.460 124.240 ;
        RECT 149.930 123.175 150.100 123.875 ;
        RECT 150.630 123.795 150.800 124.410 ;
        RECT 150.970 124.055 151.140 124.855 ;
        RECT 151.310 124.355 151.560 124.685 ;
        RECT 151.785 124.385 152.670 124.555 ;
        RECT 150.630 123.705 151.140 123.795 ;
        RECT 149.180 122.895 149.405 123.025 ;
        RECT 149.575 122.955 150.100 123.175 ;
        RECT 150.270 123.535 151.140 123.705 ;
        RECT 148.815 122.305 149.065 122.765 ;
        RECT 149.235 122.755 149.405 122.895 ;
        RECT 150.270 122.755 150.440 123.535 ;
        RECT 150.970 123.465 151.140 123.535 ;
        RECT 150.650 123.285 150.850 123.315 ;
        RECT 151.310 123.285 151.480 124.355 ;
        RECT 151.650 123.465 151.840 124.185 ;
        RECT 150.650 122.985 151.480 123.285 ;
        RECT 152.010 123.255 152.330 124.215 ;
        RECT 149.235 122.585 149.570 122.755 ;
        RECT 149.765 122.585 150.440 122.755 ;
        RECT 150.760 122.305 151.130 122.805 ;
        RECT 151.310 122.755 151.480 122.985 ;
        RECT 151.865 122.925 152.330 123.255 ;
        RECT 152.500 123.545 152.670 124.385 ;
        RECT 152.850 124.355 153.165 124.855 ;
        RECT 153.395 124.125 153.735 124.685 ;
        RECT 152.840 123.750 153.735 124.125 ;
        RECT 153.905 123.845 154.075 124.855 ;
        RECT 153.545 123.545 153.735 123.750 ;
        RECT 154.245 123.795 154.575 124.640 ;
        RECT 154.245 123.715 154.635 123.795 ;
        RECT 154.420 123.665 154.635 123.715 ;
        RECT 152.500 123.215 153.375 123.545 ;
        RECT 153.545 123.215 154.295 123.545 ;
        RECT 152.500 122.755 152.670 123.215 ;
        RECT 153.545 123.045 153.745 123.215 ;
        RECT 154.465 123.085 154.635 123.665 ;
        RECT 155.725 123.765 156.935 124.855 ;
        RECT 155.725 123.225 156.245 123.765 ;
        RECT 154.410 123.045 154.635 123.085 ;
        RECT 156.415 123.055 156.935 123.595 ;
        RECT 151.310 122.585 151.715 122.755 ;
        RECT 151.885 122.585 152.670 122.755 ;
        RECT 152.945 122.305 153.155 122.835 ;
        RECT 153.415 122.520 153.745 123.045 ;
        RECT 154.255 122.960 154.635 123.045 ;
        RECT 153.915 122.305 154.085 122.915 ;
        RECT 154.255 122.525 154.585 122.960 ;
        RECT 155.725 122.305 156.935 123.055 ;
        RECT 22.700 122.135 157.020 122.305 ;
        RECT 22.785 121.385 23.995 122.135 ;
        RECT 22.785 120.845 23.305 121.385 ;
        RECT 24.165 121.365 25.835 122.135 ;
        RECT 26.465 121.395 26.850 121.965 ;
        RECT 27.020 121.675 27.345 122.135 ;
        RECT 27.865 121.505 28.145 121.965 ;
        RECT 23.475 120.675 23.995 121.215 ;
        RECT 24.165 120.845 24.915 121.365 ;
        RECT 25.085 120.675 25.835 121.195 ;
        RECT 22.785 119.585 23.995 120.675 ;
        RECT 24.165 119.585 25.835 120.675 ;
        RECT 26.465 120.725 26.745 121.395 ;
        RECT 27.020 121.335 28.145 121.505 ;
        RECT 27.020 121.225 27.470 121.335 ;
        RECT 26.915 120.895 27.470 121.225 ;
        RECT 28.335 121.165 28.735 121.965 ;
        RECT 29.135 121.675 29.405 122.135 ;
        RECT 29.575 121.505 29.860 121.965 ;
        RECT 26.465 119.755 26.850 120.725 ;
        RECT 27.020 120.435 27.470 120.895 ;
        RECT 27.640 120.605 28.735 121.165 ;
        RECT 27.020 120.215 28.145 120.435 ;
        RECT 27.020 119.585 27.345 120.045 ;
        RECT 27.865 119.755 28.145 120.215 ;
        RECT 28.335 119.755 28.735 120.605 ;
        RECT 28.905 121.335 29.860 121.505 ;
        RECT 30.145 121.385 31.355 122.135 ;
        RECT 28.905 120.435 29.115 121.335 ;
        RECT 29.285 120.605 29.975 121.165 ;
        RECT 30.145 120.845 30.665 121.385 ;
        RECT 31.525 121.315 31.785 122.135 ;
        RECT 31.955 121.315 32.285 121.735 ;
        RECT 32.465 121.650 33.255 121.915 ;
        RECT 32.035 121.225 32.285 121.315 ;
        RECT 30.835 120.675 31.355 121.215 ;
        RECT 28.905 120.215 29.860 120.435 ;
        RECT 29.135 119.585 29.405 120.045 ;
        RECT 29.575 119.755 29.860 120.215 ;
        RECT 30.145 119.585 31.355 120.675 ;
        RECT 31.525 120.265 31.865 121.145 ;
        RECT 32.035 120.975 32.830 121.225 ;
        RECT 31.525 119.585 31.785 120.095 ;
        RECT 32.035 119.755 32.205 120.975 ;
        RECT 33.000 120.795 33.255 121.650 ;
        RECT 33.425 121.495 33.625 121.915 ;
        RECT 33.815 121.675 34.145 122.135 ;
        RECT 33.425 120.975 33.835 121.495 ;
        RECT 34.315 121.485 34.575 121.965 ;
        RECT 34.005 120.795 34.235 121.225 ;
        RECT 32.445 120.625 34.235 120.795 ;
        RECT 32.445 120.260 32.695 120.625 ;
        RECT 32.865 120.265 33.195 120.455 ;
        RECT 33.415 120.330 34.130 120.625 ;
        RECT 34.405 120.455 34.575 121.485 ;
        RECT 32.865 120.090 33.060 120.265 ;
        RECT 32.445 119.585 33.060 120.090 ;
        RECT 33.230 119.755 33.705 120.095 ;
        RECT 33.875 119.585 34.090 120.130 ;
        RECT 34.300 119.755 34.575 120.455 ;
        RECT 34.755 119.765 35.015 121.955 ;
        RECT 35.275 121.765 35.945 122.135 ;
        RECT 36.125 121.585 36.435 121.955 ;
        RECT 35.205 121.385 36.435 121.585 ;
        RECT 35.205 120.715 35.495 121.385 ;
        RECT 36.615 121.205 36.845 121.845 ;
        RECT 37.025 121.405 37.315 122.135 ;
        RECT 37.595 121.585 37.765 121.965 ;
        RECT 37.945 121.755 38.275 122.135 ;
        RECT 37.595 121.415 38.260 121.585 ;
        RECT 38.455 121.460 38.715 121.965 ;
        RECT 35.675 120.895 36.140 121.205 ;
        RECT 36.320 120.895 36.845 121.205 ;
        RECT 37.025 120.895 37.325 121.225 ;
        RECT 37.525 120.865 37.855 121.235 ;
        RECT 38.090 121.160 38.260 121.415 ;
        RECT 38.090 120.830 38.375 121.160 ;
        RECT 35.205 120.495 35.975 120.715 ;
        RECT 35.185 119.585 35.525 120.315 ;
        RECT 35.705 119.765 35.975 120.495 ;
        RECT 36.155 120.475 37.315 120.715 ;
        RECT 38.090 120.685 38.260 120.830 ;
        RECT 36.155 119.765 36.385 120.475 ;
        RECT 36.555 119.585 36.885 120.295 ;
        RECT 37.055 119.765 37.315 120.475 ;
        RECT 37.595 120.515 38.260 120.685 ;
        RECT 38.545 120.660 38.715 121.460 ;
        RECT 39.355 121.325 39.625 122.135 ;
        RECT 39.795 121.325 40.125 121.965 ;
        RECT 40.295 121.325 40.535 122.135 ;
        RECT 40.815 121.585 40.985 121.875 ;
        RECT 41.155 121.755 41.485 122.135 ;
        RECT 40.815 121.415 41.480 121.585 ;
        RECT 39.345 120.895 39.695 121.145 ;
        RECT 39.865 120.725 40.035 121.325 ;
        RECT 40.205 120.895 40.555 121.145 ;
        RECT 37.595 119.755 37.765 120.515 ;
        RECT 37.945 119.585 38.275 120.345 ;
        RECT 38.445 119.755 38.715 120.660 ;
        RECT 39.355 119.585 39.685 120.725 ;
        RECT 39.865 120.555 40.545 120.725 ;
        RECT 40.730 120.595 41.080 121.245 ;
        RECT 40.215 119.770 40.545 120.555 ;
        RECT 41.250 120.425 41.480 121.415 ;
        RECT 40.815 120.255 41.480 120.425 ;
        RECT 40.815 119.755 40.985 120.255 ;
        RECT 41.155 119.585 41.485 120.085 ;
        RECT 41.655 119.755 41.840 121.875 ;
        RECT 42.095 121.675 42.345 122.135 ;
        RECT 42.515 121.685 42.850 121.855 ;
        RECT 43.045 121.685 43.720 121.855 ;
        RECT 42.515 121.545 42.685 121.685 ;
        RECT 42.010 120.555 42.290 121.505 ;
        RECT 42.460 121.415 42.685 121.545 ;
        RECT 42.460 120.310 42.630 121.415 ;
        RECT 42.855 121.265 43.380 121.485 ;
        RECT 42.800 120.500 43.040 121.095 ;
        RECT 43.210 120.565 43.380 121.265 ;
        RECT 43.550 120.905 43.720 121.685 ;
        RECT 44.040 121.635 44.410 122.135 ;
        RECT 44.590 121.685 44.995 121.855 ;
        RECT 45.165 121.685 45.950 121.855 ;
        RECT 44.590 121.455 44.760 121.685 ;
        RECT 43.930 121.155 44.760 121.455 ;
        RECT 45.145 121.185 45.610 121.515 ;
        RECT 43.930 121.125 44.130 121.155 ;
        RECT 44.250 120.905 44.420 120.975 ;
        RECT 43.550 120.735 44.420 120.905 ;
        RECT 43.910 120.645 44.420 120.735 ;
        RECT 42.460 120.180 42.765 120.310 ;
        RECT 43.210 120.200 43.740 120.565 ;
        RECT 42.080 119.585 42.345 120.045 ;
        RECT 42.515 119.755 42.765 120.180 ;
        RECT 43.910 120.030 44.080 120.645 ;
        RECT 42.975 119.860 44.080 120.030 ;
        RECT 44.250 119.585 44.420 120.385 ;
        RECT 44.590 120.085 44.760 121.155 ;
        RECT 44.930 120.255 45.120 120.975 ;
        RECT 45.290 120.225 45.610 121.185 ;
        RECT 45.780 121.225 45.950 121.685 ;
        RECT 46.225 121.605 46.435 122.135 ;
        RECT 46.695 121.395 47.025 121.920 ;
        RECT 47.195 121.525 47.365 122.135 ;
        RECT 47.535 121.480 47.865 121.915 ;
        RECT 47.535 121.395 47.915 121.480 ;
        RECT 48.545 121.410 48.835 122.135 ;
        RECT 46.825 121.225 47.025 121.395 ;
        RECT 47.690 121.355 47.915 121.395 ;
        RECT 45.780 120.895 46.655 121.225 ;
        RECT 46.825 120.895 47.575 121.225 ;
        RECT 44.590 119.755 44.840 120.085 ;
        RECT 45.780 120.055 45.950 120.895 ;
        RECT 46.825 120.690 47.015 120.895 ;
        RECT 47.745 120.775 47.915 121.355 ;
        RECT 49.005 121.385 50.215 122.135 ;
        RECT 50.475 121.795 50.645 121.830 ;
        RECT 50.445 121.625 50.645 121.795 ;
        RECT 49.005 120.845 49.525 121.385 ;
        RECT 50.475 121.265 50.645 121.625 ;
        RECT 50.835 121.605 51.065 121.910 ;
        RECT 51.235 121.775 51.565 122.135 ;
        RECT 51.760 121.605 52.050 121.955 ;
        RECT 50.835 121.435 52.050 121.605 ;
        RECT 52.315 121.585 52.485 121.875 ;
        RECT 52.655 121.755 52.985 122.135 ;
        RECT 52.315 121.415 52.980 121.585 ;
        RECT 47.700 120.725 47.915 120.775 ;
        RECT 46.120 120.315 47.015 120.690 ;
        RECT 47.525 120.645 47.915 120.725 ;
        RECT 45.065 119.885 45.950 120.055 ;
        RECT 46.130 119.585 46.445 120.085 ;
        RECT 46.675 119.755 47.015 120.315 ;
        RECT 47.185 119.585 47.355 120.595 ;
        RECT 47.525 119.800 47.855 120.645 ;
        RECT 48.545 119.585 48.835 120.750 ;
        RECT 49.695 120.675 50.215 121.215 ;
        RECT 50.475 121.095 50.995 121.265 ;
        RECT 49.005 119.585 50.215 120.675 ;
        RECT 50.390 120.565 50.635 120.925 ;
        RECT 50.825 120.715 50.995 121.095 ;
        RECT 51.165 120.895 51.550 121.225 ;
        RECT 51.730 121.115 51.990 121.225 ;
        RECT 51.730 120.945 51.995 121.115 ;
        RECT 51.730 120.895 51.990 120.945 ;
        RECT 50.825 120.435 51.175 120.715 ;
        RECT 50.390 119.585 50.645 120.385 ;
        RECT 50.845 119.755 51.175 120.435 ;
        RECT 51.355 119.845 51.550 120.895 ;
        RECT 51.730 119.585 52.050 120.725 ;
        RECT 52.230 120.595 52.580 121.245 ;
        RECT 52.750 120.425 52.980 121.415 ;
        RECT 52.315 120.255 52.980 120.425 ;
        RECT 52.315 119.755 52.485 120.255 ;
        RECT 52.655 119.585 52.985 120.085 ;
        RECT 53.155 119.755 53.340 121.875 ;
        RECT 53.595 121.675 53.845 122.135 ;
        RECT 54.015 121.685 54.350 121.855 ;
        RECT 54.545 121.685 55.220 121.855 ;
        RECT 54.015 121.545 54.185 121.685 ;
        RECT 53.510 120.555 53.790 121.505 ;
        RECT 53.960 121.415 54.185 121.545 ;
        RECT 53.960 120.310 54.130 121.415 ;
        RECT 54.355 121.265 54.880 121.485 ;
        RECT 54.300 120.500 54.540 121.095 ;
        RECT 54.710 120.565 54.880 121.265 ;
        RECT 55.050 120.905 55.220 121.685 ;
        RECT 55.540 121.635 55.910 122.135 ;
        RECT 56.090 121.685 56.495 121.855 ;
        RECT 56.665 121.685 57.450 121.855 ;
        RECT 56.090 121.455 56.260 121.685 ;
        RECT 55.430 121.155 56.260 121.455 ;
        RECT 56.645 121.185 57.110 121.515 ;
        RECT 55.430 121.125 55.630 121.155 ;
        RECT 55.750 120.905 55.920 120.975 ;
        RECT 55.050 120.735 55.920 120.905 ;
        RECT 55.410 120.645 55.920 120.735 ;
        RECT 53.960 120.180 54.265 120.310 ;
        RECT 54.710 120.200 55.240 120.565 ;
        RECT 53.580 119.585 53.845 120.045 ;
        RECT 54.015 119.755 54.265 120.180 ;
        RECT 55.410 120.030 55.580 120.645 ;
        RECT 54.475 119.860 55.580 120.030 ;
        RECT 55.750 119.585 55.920 120.385 ;
        RECT 56.090 120.085 56.260 121.155 ;
        RECT 56.430 120.255 56.620 120.975 ;
        RECT 56.790 120.225 57.110 121.185 ;
        RECT 57.280 121.225 57.450 121.685 ;
        RECT 57.725 121.605 57.935 122.135 ;
        RECT 58.195 121.395 58.525 121.920 ;
        RECT 58.695 121.525 58.865 122.135 ;
        RECT 59.035 121.480 59.365 121.915 ;
        RECT 59.675 121.585 59.845 121.875 ;
        RECT 60.015 121.755 60.345 122.135 ;
        RECT 59.035 121.395 59.415 121.480 ;
        RECT 59.675 121.415 60.340 121.585 ;
        RECT 58.325 121.225 58.525 121.395 ;
        RECT 59.190 121.355 59.415 121.395 ;
        RECT 57.280 120.895 58.155 121.225 ;
        RECT 58.325 120.895 59.075 121.225 ;
        RECT 56.090 119.755 56.340 120.085 ;
        RECT 57.280 120.055 57.450 120.895 ;
        RECT 58.325 120.690 58.515 120.895 ;
        RECT 59.245 120.775 59.415 121.355 ;
        RECT 59.200 120.725 59.415 120.775 ;
        RECT 57.620 120.315 58.515 120.690 ;
        RECT 59.025 120.645 59.415 120.725 ;
        RECT 56.565 119.885 57.450 120.055 ;
        RECT 57.630 119.585 57.945 120.085 ;
        RECT 58.175 119.755 58.515 120.315 ;
        RECT 58.685 119.585 58.855 120.595 ;
        RECT 59.025 119.800 59.355 120.645 ;
        RECT 59.590 120.595 59.940 121.245 ;
        RECT 60.110 120.425 60.340 121.415 ;
        RECT 59.675 120.255 60.340 120.425 ;
        RECT 59.675 119.755 59.845 120.255 ;
        RECT 60.015 119.585 60.345 120.085 ;
        RECT 60.515 119.755 60.700 121.875 ;
        RECT 60.955 121.675 61.205 122.135 ;
        RECT 61.375 121.685 61.710 121.855 ;
        RECT 61.905 121.685 62.580 121.855 ;
        RECT 61.375 121.545 61.545 121.685 ;
        RECT 60.870 120.555 61.150 121.505 ;
        RECT 61.320 121.415 61.545 121.545 ;
        RECT 61.320 120.310 61.490 121.415 ;
        RECT 61.715 121.265 62.240 121.485 ;
        RECT 61.660 120.500 61.900 121.095 ;
        RECT 62.070 120.565 62.240 121.265 ;
        RECT 62.410 120.905 62.580 121.685 ;
        RECT 62.900 121.635 63.270 122.135 ;
        RECT 63.450 121.685 63.855 121.855 ;
        RECT 64.025 121.685 64.810 121.855 ;
        RECT 63.450 121.455 63.620 121.685 ;
        RECT 62.790 121.155 63.620 121.455 ;
        RECT 64.005 121.185 64.470 121.515 ;
        RECT 62.790 121.125 62.990 121.155 ;
        RECT 63.110 120.905 63.280 120.975 ;
        RECT 62.410 120.735 63.280 120.905 ;
        RECT 62.770 120.645 63.280 120.735 ;
        RECT 61.320 120.180 61.625 120.310 ;
        RECT 62.070 120.200 62.600 120.565 ;
        RECT 60.940 119.585 61.205 120.045 ;
        RECT 61.375 119.755 61.625 120.180 ;
        RECT 62.770 120.030 62.940 120.645 ;
        RECT 61.835 119.860 62.940 120.030 ;
        RECT 63.110 119.585 63.280 120.385 ;
        RECT 63.450 120.085 63.620 121.155 ;
        RECT 63.790 120.255 63.980 120.975 ;
        RECT 64.150 120.225 64.470 121.185 ;
        RECT 64.640 121.225 64.810 121.685 ;
        RECT 65.085 121.605 65.295 122.135 ;
        RECT 65.555 121.395 65.885 121.920 ;
        RECT 66.055 121.525 66.225 122.135 ;
        RECT 66.395 121.480 66.725 121.915 ;
        RECT 66.395 121.395 66.775 121.480 ;
        RECT 65.685 121.225 65.885 121.395 ;
        RECT 66.550 121.355 66.775 121.395 ;
        RECT 64.640 120.895 65.515 121.225 ;
        RECT 65.685 120.895 66.435 121.225 ;
        RECT 63.450 119.755 63.700 120.085 ;
        RECT 64.640 120.055 64.810 120.895 ;
        RECT 65.685 120.690 65.875 120.895 ;
        RECT 66.605 120.775 66.775 121.355 ;
        RECT 66.560 120.725 66.775 120.775 ;
        RECT 64.980 120.315 65.875 120.690 ;
        RECT 66.385 120.645 66.775 120.725 ;
        RECT 63.925 119.885 64.810 120.055 ;
        RECT 64.990 119.585 65.305 120.085 ;
        RECT 65.535 119.755 65.875 120.315 ;
        RECT 66.045 119.585 66.215 120.595 ;
        RECT 66.385 119.800 66.715 120.645 ;
        RECT 66.955 119.765 67.215 121.955 ;
        RECT 67.475 121.765 68.145 122.135 ;
        RECT 68.325 121.585 68.635 121.955 ;
        RECT 67.405 121.385 68.635 121.585 ;
        RECT 67.405 120.715 67.695 121.385 ;
        RECT 68.815 121.205 69.045 121.845 ;
        RECT 69.225 121.405 69.515 122.135 ;
        RECT 69.820 121.505 70.105 121.965 ;
        RECT 70.275 121.675 70.545 122.135 ;
        RECT 69.820 121.335 70.775 121.505 ;
        RECT 67.875 120.895 68.340 121.205 ;
        RECT 68.520 120.895 69.045 121.205 ;
        RECT 69.225 120.895 69.525 121.225 ;
        RECT 67.405 120.495 68.175 120.715 ;
        RECT 67.385 119.585 67.725 120.315 ;
        RECT 67.905 119.765 68.175 120.495 ;
        RECT 68.355 120.475 69.515 120.715 ;
        RECT 69.705 120.605 70.395 121.165 ;
        RECT 68.355 119.765 68.585 120.475 ;
        RECT 68.755 119.585 69.085 120.295 ;
        RECT 69.255 119.765 69.515 120.475 ;
        RECT 70.565 120.435 70.775 121.335 ;
        RECT 69.820 120.215 70.775 120.435 ;
        RECT 70.945 121.165 71.345 121.965 ;
        RECT 71.535 121.505 71.815 121.965 ;
        RECT 72.335 121.675 72.660 122.135 ;
        RECT 71.535 121.335 72.660 121.505 ;
        RECT 72.830 121.395 73.215 121.965 ;
        RECT 74.305 121.410 74.595 122.135 ;
        RECT 72.210 121.225 72.660 121.335 ;
        RECT 70.945 120.605 72.040 121.165 ;
        RECT 72.210 120.895 72.765 121.225 ;
        RECT 69.820 119.755 70.105 120.215 ;
        RECT 70.275 119.585 70.545 120.045 ;
        RECT 70.945 119.755 71.345 120.605 ;
        RECT 72.210 120.435 72.660 120.895 ;
        RECT 72.935 120.725 73.215 121.395 ;
        RECT 74.775 121.325 75.045 122.135 ;
        RECT 75.215 121.325 75.545 121.965 ;
        RECT 75.715 121.325 75.955 122.135 ;
        RECT 76.145 121.590 81.490 122.135 ;
        RECT 74.765 120.895 75.115 121.145 ;
        RECT 71.535 120.215 72.660 120.435 ;
        RECT 71.535 119.755 71.815 120.215 ;
        RECT 72.335 119.585 72.660 120.045 ;
        RECT 72.830 119.755 73.215 120.725 ;
        RECT 74.305 119.585 74.595 120.750 ;
        RECT 75.285 120.725 75.455 121.325 ;
        RECT 75.625 120.895 75.975 121.145 ;
        RECT 77.730 120.760 78.070 121.590 ;
        RECT 81.665 121.365 83.335 122.135 ;
        RECT 83.505 121.395 83.890 121.965 ;
        RECT 84.060 121.675 84.385 122.135 ;
        RECT 84.905 121.505 85.185 121.965 ;
        RECT 74.775 119.585 75.105 120.725 ;
        RECT 75.285 120.555 75.965 120.725 ;
        RECT 75.635 119.770 75.965 120.555 ;
        RECT 79.550 120.020 79.900 121.270 ;
        RECT 81.665 120.845 82.415 121.365 ;
        RECT 82.585 120.675 83.335 121.195 ;
        RECT 76.145 119.585 81.490 120.020 ;
        RECT 81.665 119.585 83.335 120.675 ;
        RECT 83.505 120.725 83.785 121.395 ;
        RECT 84.060 121.335 85.185 121.505 ;
        RECT 84.060 121.225 84.510 121.335 ;
        RECT 83.955 120.895 84.510 121.225 ;
        RECT 85.375 121.165 85.775 121.965 ;
        RECT 86.175 121.675 86.445 122.135 ;
        RECT 86.615 121.505 86.900 121.965 ;
        RECT 83.505 119.755 83.890 120.725 ;
        RECT 84.060 120.435 84.510 120.895 ;
        RECT 84.680 120.605 85.775 121.165 ;
        RECT 84.060 120.215 85.185 120.435 ;
        RECT 84.060 119.585 84.385 120.045 ;
        RECT 84.905 119.755 85.185 120.215 ;
        RECT 85.375 119.755 85.775 120.605 ;
        RECT 85.945 121.335 86.900 121.505 ;
        RECT 87.185 121.385 88.395 122.135 ;
        RECT 88.730 121.625 88.970 122.135 ;
        RECT 89.150 121.625 89.430 121.955 ;
        RECT 89.660 121.625 89.875 122.135 ;
        RECT 85.945 120.435 86.155 121.335 ;
        RECT 86.325 120.605 87.015 121.165 ;
        RECT 87.185 120.845 87.705 121.385 ;
        RECT 87.875 120.675 88.395 121.215 ;
        RECT 88.625 120.895 88.980 121.455 ;
        RECT 89.150 120.725 89.320 121.625 ;
        RECT 89.490 120.895 89.755 121.455 ;
        RECT 90.045 121.395 90.660 121.965 ;
        RECT 90.005 120.725 90.175 121.225 ;
        RECT 85.945 120.215 86.900 120.435 ;
        RECT 86.175 119.585 86.445 120.045 ;
        RECT 86.615 119.755 86.900 120.215 ;
        RECT 87.185 119.585 88.395 120.675 ;
        RECT 88.750 120.555 90.175 120.725 ;
        RECT 88.750 120.380 89.140 120.555 ;
        RECT 89.625 119.585 89.955 120.385 ;
        RECT 90.345 120.375 90.660 121.395 ;
        RECT 90.125 119.755 90.660 120.375 ;
        RECT 90.865 121.485 91.125 121.965 ;
        RECT 91.295 121.595 91.545 122.135 ;
        RECT 90.865 120.455 91.035 121.485 ;
        RECT 91.715 121.430 91.935 121.915 ;
        RECT 91.205 120.835 91.435 121.230 ;
        RECT 91.605 121.005 91.935 121.430 ;
        RECT 92.105 121.755 92.995 121.925 ;
        RECT 92.105 121.030 92.275 121.755 ;
        RECT 92.445 121.200 92.995 121.585 ;
        RECT 93.625 121.395 94.010 121.965 ;
        RECT 94.180 121.675 94.505 122.135 ;
        RECT 95.025 121.505 95.305 121.965 ;
        RECT 92.105 120.960 92.995 121.030 ;
        RECT 92.100 120.935 92.995 120.960 ;
        RECT 92.090 120.920 92.995 120.935 ;
        RECT 92.085 120.905 92.995 120.920 ;
        RECT 92.075 120.900 92.995 120.905 ;
        RECT 92.070 120.890 92.995 120.900 ;
        RECT 92.065 120.880 92.995 120.890 ;
        RECT 92.055 120.875 92.995 120.880 ;
        RECT 92.045 120.865 92.995 120.875 ;
        RECT 92.035 120.860 92.995 120.865 ;
        RECT 92.035 120.855 92.370 120.860 ;
        RECT 92.020 120.850 92.370 120.855 ;
        RECT 92.005 120.840 92.370 120.850 ;
        RECT 91.980 120.835 92.370 120.840 ;
        RECT 91.205 120.830 92.370 120.835 ;
        RECT 91.205 120.795 92.340 120.830 ;
        RECT 91.205 120.770 92.305 120.795 ;
        RECT 91.205 120.740 92.275 120.770 ;
        RECT 91.205 120.710 92.255 120.740 ;
        RECT 91.205 120.680 92.235 120.710 ;
        RECT 91.205 120.670 92.165 120.680 ;
        RECT 91.205 120.660 92.140 120.670 ;
        RECT 91.205 120.645 92.120 120.660 ;
        RECT 91.205 120.630 92.100 120.645 ;
        RECT 91.310 120.620 92.095 120.630 ;
        RECT 91.310 120.585 92.080 120.620 ;
        RECT 90.865 119.755 91.140 120.455 ;
        RECT 91.310 120.335 92.065 120.585 ;
        RECT 92.235 120.265 92.565 120.510 ;
        RECT 92.735 120.410 92.995 120.860 ;
        RECT 93.625 120.725 93.905 121.395 ;
        RECT 94.180 121.335 95.305 121.505 ;
        RECT 94.180 121.225 94.630 121.335 ;
        RECT 94.075 120.895 94.630 121.225 ;
        RECT 95.495 121.165 95.895 121.965 ;
        RECT 96.295 121.675 96.565 122.135 ;
        RECT 96.735 121.505 97.020 121.965 ;
        RECT 92.380 120.240 92.565 120.265 ;
        RECT 92.380 120.140 92.995 120.240 ;
        RECT 91.310 119.585 91.565 120.130 ;
        RECT 91.735 119.755 92.215 120.095 ;
        RECT 92.390 119.585 92.995 120.140 ;
        RECT 93.625 119.755 94.010 120.725 ;
        RECT 94.180 120.435 94.630 120.895 ;
        RECT 94.800 120.605 95.895 121.165 ;
        RECT 94.180 120.215 95.305 120.435 ;
        RECT 94.180 119.585 94.505 120.045 ;
        RECT 95.025 119.755 95.305 120.215 ;
        RECT 95.495 119.755 95.895 120.605 ;
        RECT 96.065 121.335 97.020 121.505 ;
        RECT 96.065 120.435 96.275 121.335 ;
        RECT 96.445 120.605 97.135 121.165 ;
        RECT 96.065 120.215 97.020 120.435 ;
        RECT 96.295 119.585 96.565 120.045 ;
        RECT 96.735 119.755 97.020 120.215 ;
        RECT 97.315 119.765 97.575 121.955 ;
        RECT 97.835 121.765 98.505 122.135 ;
        RECT 98.685 121.585 98.995 121.955 ;
        RECT 97.765 121.385 98.995 121.585 ;
        RECT 97.765 120.715 98.055 121.385 ;
        RECT 99.175 121.205 99.405 121.845 ;
        RECT 99.585 121.405 99.875 122.135 ;
        RECT 100.065 121.410 100.355 122.135 ;
        RECT 100.525 121.385 101.735 122.135 ;
        RECT 101.995 121.585 102.165 121.875 ;
        RECT 102.335 121.755 102.665 122.135 ;
        RECT 101.995 121.415 102.660 121.585 ;
        RECT 98.235 120.895 98.700 121.205 ;
        RECT 98.880 120.895 99.405 121.205 ;
        RECT 99.585 120.895 99.885 121.225 ;
        RECT 100.525 120.845 101.045 121.385 ;
        RECT 97.765 120.495 98.535 120.715 ;
        RECT 97.745 119.585 98.085 120.315 ;
        RECT 98.265 119.765 98.535 120.495 ;
        RECT 98.715 120.475 99.875 120.715 ;
        RECT 98.715 119.765 98.945 120.475 ;
        RECT 99.115 119.585 99.445 120.295 ;
        RECT 99.615 119.765 99.875 120.475 ;
        RECT 100.065 119.585 100.355 120.750 ;
        RECT 101.215 120.675 101.735 121.215 ;
        RECT 100.525 119.585 101.735 120.675 ;
        RECT 101.910 120.595 102.260 121.245 ;
        RECT 102.430 120.425 102.660 121.415 ;
        RECT 101.995 120.255 102.660 120.425 ;
        RECT 101.995 119.755 102.165 120.255 ;
        RECT 102.335 119.585 102.665 120.085 ;
        RECT 102.835 119.755 103.020 121.875 ;
        RECT 103.275 121.675 103.525 122.135 ;
        RECT 103.695 121.685 104.030 121.855 ;
        RECT 104.225 121.685 104.900 121.855 ;
        RECT 103.695 121.545 103.865 121.685 ;
        RECT 103.190 120.555 103.470 121.505 ;
        RECT 103.640 121.415 103.865 121.545 ;
        RECT 103.640 120.310 103.810 121.415 ;
        RECT 104.035 121.265 104.560 121.485 ;
        RECT 103.980 120.500 104.220 121.095 ;
        RECT 104.390 120.565 104.560 121.265 ;
        RECT 104.730 120.905 104.900 121.685 ;
        RECT 105.220 121.635 105.590 122.135 ;
        RECT 105.770 121.685 106.175 121.855 ;
        RECT 106.345 121.685 107.130 121.855 ;
        RECT 105.770 121.455 105.940 121.685 ;
        RECT 105.110 121.155 105.940 121.455 ;
        RECT 106.325 121.185 106.790 121.515 ;
        RECT 105.110 121.125 105.310 121.155 ;
        RECT 105.430 120.905 105.600 120.975 ;
        RECT 104.730 120.735 105.600 120.905 ;
        RECT 105.090 120.645 105.600 120.735 ;
        RECT 103.640 120.180 103.945 120.310 ;
        RECT 104.390 120.200 104.920 120.565 ;
        RECT 103.260 119.585 103.525 120.045 ;
        RECT 103.695 119.755 103.945 120.180 ;
        RECT 105.090 120.030 105.260 120.645 ;
        RECT 104.155 119.860 105.260 120.030 ;
        RECT 105.430 119.585 105.600 120.385 ;
        RECT 105.770 120.085 105.940 121.155 ;
        RECT 106.110 120.255 106.300 120.975 ;
        RECT 106.470 120.225 106.790 121.185 ;
        RECT 106.960 121.225 107.130 121.685 ;
        RECT 107.405 121.605 107.615 122.135 ;
        RECT 107.875 121.395 108.205 121.920 ;
        RECT 108.375 121.525 108.545 122.135 ;
        RECT 108.715 121.480 109.045 121.915 ;
        RECT 109.840 121.505 110.125 121.965 ;
        RECT 110.295 121.675 110.565 122.135 ;
        RECT 108.715 121.395 109.095 121.480 ;
        RECT 108.005 121.225 108.205 121.395 ;
        RECT 108.870 121.355 109.095 121.395 ;
        RECT 106.960 120.895 107.835 121.225 ;
        RECT 108.005 120.895 108.755 121.225 ;
        RECT 105.770 119.755 106.020 120.085 ;
        RECT 106.960 120.055 107.130 120.895 ;
        RECT 108.005 120.690 108.195 120.895 ;
        RECT 108.925 120.775 109.095 121.355 ;
        RECT 109.840 121.335 110.795 121.505 ;
        RECT 108.880 120.725 109.095 120.775 ;
        RECT 107.300 120.315 108.195 120.690 ;
        RECT 108.705 120.645 109.095 120.725 ;
        RECT 106.245 119.885 107.130 120.055 ;
        RECT 107.310 119.585 107.625 120.085 ;
        RECT 107.855 119.755 108.195 120.315 ;
        RECT 108.365 119.585 108.535 120.595 ;
        RECT 108.705 119.800 109.035 120.645 ;
        RECT 109.725 120.605 110.415 121.165 ;
        RECT 110.585 120.435 110.795 121.335 ;
        RECT 109.840 120.215 110.795 120.435 ;
        RECT 110.965 121.165 111.365 121.965 ;
        RECT 111.555 121.505 111.835 121.965 ;
        RECT 112.355 121.675 112.680 122.135 ;
        RECT 111.555 121.335 112.680 121.505 ;
        RECT 112.850 121.395 113.235 121.965 ;
        RECT 112.230 121.225 112.680 121.335 ;
        RECT 110.965 120.605 112.060 121.165 ;
        RECT 112.230 120.895 112.785 121.225 ;
        RECT 109.840 119.755 110.125 120.215 ;
        RECT 110.295 119.585 110.565 120.045 ;
        RECT 110.965 119.755 111.365 120.605 ;
        RECT 112.230 120.435 112.680 120.895 ;
        RECT 112.955 120.725 113.235 121.395 ;
        RECT 111.555 120.215 112.680 120.435 ;
        RECT 111.555 119.755 111.835 120.215 ;
        RECT 112.355 119.585 112.680 120.045 ;
        RECT 112.850 119.755 113.235 120.725 ;
        RECT 113.405 121.485 113.665 121.965 ;
        RECT 113.835 121.595 114.085 122.135 ;
        RECT 113.405 120.455 113.575 121.485 ;
        RECT 114.255 121.430 114.475 121.915 ;
        RECT 113.745 120.835 113.975 121.230 ;
        RECT 114.145 121.005 114.475 121.430 ;
        RECT 114.645 121.755 115.535 121.925 ;
        RECT 114.645 121.030 114.815 121.755 ;
        RECT 114.985 121.200 115.535 121.585 ;
        RECT 116.675 121.480 117.005 121.915 ;
        RECT 117.175 121.525 117.345 122.135 ;
        RECT 116.625 121.395 117.005 121.480 ;
        RECT 117.515 121.395 117.845 121.920 ;
        RECT 118.105 121.605 118.315 122.135 ;
        RECT 118.590 121.685 119.375 121.855 ;
        RECT 119.545 121.685 119.950 121.855 ;
        RECT 116.625 121.355 116.850 121.395 ;
        RECT 114.645 120.960 115.535 121.030 ;
        RECT 114.640 120.935 115.535 120.960 ;
        RECT 114.630 120.920 115.535 120.935 ;
        RECT 114.625 120.905 115.535 120.920 ;
        RECT 114.615 120.900 115.535 120.905 ;
        RECT 114.610 120.890 115.535 120.900 ;
        RECT 114.605 120.880 115.535 120.890 ;
        RECT 114.595 120.875 115.535 120.880 ;
        RECT 114.585 120.865 115.535 120.875 ;
        RECT 114.575 120.860 115.535 120.865 ;
        RECT 114.575 120.855 114.910 120.860 ;
        RECT 114.560 120.850 114.910 120.855 ;
        RECT 114.545 120.840 114.910 120.850 ;
        RECT 114.520 120.835 114.910 120.840 ;
        RECT 113.745 120.830 114.910 120.835 ;
        RECT 113.745 120.795 114.880 120.830 ;
        RECT 113.745 120.770 114.845 120.795 ;
        RECT 113.745 120.740 114.815 120.770 ;
        RECT 113.745 120.710 114.795 120.740 ;
        RECT 113.745 120.680 114.775 120.710 ;
        RECT 113.745 120.670 114.705 120.680 ;
        RECT 113.745 120.660 114.680 120.670 ;
        RECT 113.745 120.645 114.660 120.660 ;
        RECT 113.745 120.630 114.640 120.645 ;
        RECT 113.850 120.620 114.635 120.630 ;
        RECT 113.850 120.585 114.620 120.620 ;
        RECT 113.405 119.755 113.680 120.455 ;
        RECT 113.850 120.335 114.605 120.585 ;
        RECT 114.775 120.265 115.105 120.510 ;
        RECT 115.275 120.410 115.535 120.860 ;
        RECT 116.625 120.775 116.795 121.355 ;
        RECT 117.515 121.225 117.715 121.395 ;
        RECT 118.590 121.225 118.760 121.685 ;
        RECT 116.965 120.895 117.715 121.225 ;
        RECT 117.885 120.895 118.760 121.225 ;
        RECT 116.625 120.725 116.840 120.775 ;
        RECT 116.625 120.645 117.015 120.725 ;
        RECT 114.920 120.240 115.105 120.265 ;
        RECT 114.920 120.140 115.535 120.240 ;
        RECT 113.850 119.585 114.105 120.130 ;
        RECT 114.275 119.755 114.755 120.095 ;
        RECT 114.930 119.585 115.535 120.140 ;
        RECT 116.685 119.800 117.015 120.645 ;
        RECT 117.525 120.690 117.715 120.895 ;
        RECT 117.185 119.585 117.355 120.595 ;
        RECT 117.525 120.315 118.420 120.690 ;
        RECT 117.525 119.755 117.865 120.315 ;
        RECT 118.095 119.585 118.410 120.085 ;
        RECT 118.590 120.055 118.760 120.895 ;
        RECT 118.930 121.185 119.395 121.515 ;
        RECT 119.780 121.455 119.950 121.685 ;
        RECT 120.130 121.635 120.500 122.135 ;
        RECT 120.820 121.685 121.495 121.855 ;
        RECT 121.690 121.685 122.025 121.855 ;
        RECT 118.930 120.225 119.250 121.185 ;
        RECT 119.780 121.155 120.610 121.455 ;
        RECT 119.420 120.255 119.610 120.975 ;
        RECT 119.780 120.085 119.950 121.155 ;
        RECT 120.410 121.125 120.610 121.155 ;
        RECT 120.120 120.905 120.290 120.975 ;
        RECT 120.820 120.905 120.990 121.685 ;
        RECT 121.855 121.545 122.025 121.685 ;
        RECT 122.195 121.675 122.445 122.135 ;
        RECT 120.120 120.735 120.990 120.905 ;
        RECT 121.160 121.265 121.685 121.485 ;
        RECT 121.855 121.415 122.080 121.545 ;
        RECT 120.120 120.645 120.630 120.735 ;
        RECT 118.590 119.885 119.475 120.055 ;
        RECT 119.700 119.755 119.950 120.085 ;
        RECT 120.120 119.585 120.290 120.385 ;
        RECT 120.460 120.030 120.630 120.645 ;
        RECT 121.160 120.565 121.330 121.265 ;
        RECT 120.800 120.200 121.330 120.565 ;
        RECT 121.500 120.500 121.740 121.095 ;
        RECT 121.910 120.310 122.080 121.415 ;
        RECT 122.250 120.555 122.530 121.505 ;
        RECT 121.775 120.180 122.080 120.310 ;
        RECT 120.460 119.860 121.565 120.030 ;
        RECT 121.775 119.755 122.025 120.180 ;
        RECT 122.195 119.585 122.460 120.045 ;
        RECT 122.700 119.755 122.885 121.875 ;
        RECT 123.055 121.755 123.385 122.135 ;
        RECT 123.555 121.585 123.725 121.875 ;
        RECT 123.060 121.415 123.725 121.585 ;
        RECT 123.985 121.460 124.245 121.965 ;
        RECT 124.425 121.755 124.755 122.135 ;
        RECT 124.935 121.585 125.105 121.965 ;
        RECT 123.060 120.425 123.290 121.415 ;
        RECT 123.460 120.595 123.810 121.245 ;
        RECT 123.985 120.660 124.155 121.460 ;
        RECT 124.440 121.415 125.105 121.585 ;
        RECT 124.440 121.160 124.610 121.415 ;
        RECT 125.825 121.410 126.115 122.135 ;
        RECT 126.285 121.335 126.980 121.965 ;
        RECT 127.185 121.335 127.495 122.135 ;
        RECT 127.830 121.625 128.070 122.135 ;
        RECT 128.250 121.625 128.530 121.955 ;
        RECT 128.760 121.625 128.975 122.135 ;
        RECT 124.325 120.830 124.610 121.160 ;
        RECT 124.845 120.865 125.175 121.235 ;
        RECT 126.305 120.895 126.640 121.145 ;
        RECT 124.440 120.685 124.610 120.830 ;
        RECT 123.060 120.255 123.725 120.425 ;
        RECT 123.055 119.585 123.385 120.085 ;
        RECT 123.555 119.755 123.725 120.255 ;
        RECT 123.985 119.755 124.255 120.660 ;
        RECT 124.440 120.515 125.105 120.685 ;
        RECT 124.425 119.585 124.755 120.345 ;
        RECT 124.935 119.755 125.105 120.515 ;
        RECT 125.825 119.585 126.115 120.750 ;
        RECT 126.810 120.735 126.980 121.335 ;
        RECT 127.150 120.895 127.485 121.165 ;
        RECT 127.725 120.895 128.080 121.455 ;
        RECT 126.285 119.585 126.545 120.725 ;
        RECT 126.715 119.755 127.045 120.735 ;
        RECT 128.250 120.725 128.420 121.625 ;
        RECT 128.590 120.895 128.855 121.455 ;
        RECT 129.145 121.395 129.760 121.965 ;
        RECT 129.105 120.725 129.275 121.225 ;
        RECT 127.215 119.585 127.495 120.725 ;
        RECT 127.850 120.555 129.275 120.725 ;
        RECT 127.850 120.380 128.240 120.555 ;
        RECT 128.725 119.585 129.055 120.385 ;
        RECT 129.445 120.375 129.760 121.395 ;
        RECT 129.225 119.755 129.760 120.375 ;
        RECT 129.965 121.395 130.350 121.965 ;
        RECT 130.520 121.675 130.845 122.135 ;
        RECT 131.365 121.505 131.645 121.965 ;
        RECT 129.965 120.725 130.245 121.395 ;
        RECT 130.520 121.335 131.645 121.505 ;
        RECT 130.520 121.225 130.970 121.335 ;
        RECT 130.415 120.895 130.970 121.225 ;
        RECT 131.835 121.165 132.235 121.965 ;
        RECT 132.635 121.675 132.905 122.135 ;
        RECT 133.075 121.505 133.360 121.965 ;
        RECT 129.965 119.755 130.350 120.725 ;
        RECT 130.520 120.435 130.970 120.895 ;
        RECT 131.140 120.605 132.235 121.165 ;
        RECT 130.520 120.215 131.645 120.435 ;
        RECT 130.520 119.585 130.845 120.045 ;
        RECT 131.365 119.755 131.645 120.215 ;
        RECT 131.835 119.755 132.235 120.605 ;
        RECT 132.405 121.335 133.360 121.505 ;
        RECT 133.645 121.335 133.985 121.965 ;
        RECT 134.155 121.335 134.405 122.135 ;
        RECT 134.595 121.485 134.925 121.965 ;
        RECT 135.095 121.675 135.320 122.135 ;
        RECT 135.490 121.485 135.820 121.965 ;
        RECT 132.405 120.435 132.615 121.335 ;
        RECT 132.785 120.605 133.475 121.165 ;
        RECT 133.645 120.775 133.820 121.335 ;
        RECT 134.595 121.315 135.820 121.485 ;
        RECT 136.450 121.355 136.950 121.965 ;
        RECT 137.530 121.355 138.030 121.965 ;
        RECT 133.990 120.975 134.685 121.145 ;
        RECT 133.645 120.725 133.875 120.775 ;
        RECT 134.515 120.725 134.685 120.975 ;
        RECT 134.860 120.945 135.280 121.145 ;
        RECT 135.450 120.945 135.780 121.145 ;
        RECT 135.950 120.945 136.280 121.145 ;
        RECT 136.450 120.725 136.620 121.355 ;
        RECT 136.805 120.895 137.155 121.145 ;
        RECT 137.325 120.895 137.675 121.145 ;
        RECT 137.860 120.725 138.030 121.355 ;
        RECT 138.660 121.485 138.990 121.965 ;
        RECT 139.160 121.675 139.385 122.135 ;
        RECT 139.555 121.485 139.885 121.965 ;
        RECT 138.660 121.315 139.885 121.485 ;
        RECT 140.075 121.335 140.325 122.135 ;
        RECT 140.495 121.335 140.835 121.965 ;
        RECT 138.200 120.945 138.530 121.145 ;
        RECT 138.700 120.945 139.030 121.145 ;
        RECT 139.200 120.945 139.620 121.145 ;
        RECT 139.795 120.975 140.490 121.145 ;
        RECT 139.795 120.725 139.965 120.975 ;
        RECT 140.660 120.725 140.835 121.335 ;
        RECT 132.405 120.215 133.360 120.435 ;
        RECT 132.635 119.585 132.905 120.045 ;
        RECT 133.075 119.755 133.360 120.215 ;
        RECT 133.645 119.755 133.985 120.725 ;
        RECT 134.155 119.585 134.325 120.725 ;
        RECT 134.515 120.555 136.950 120.725 ;
        RECT 134.595 119.585 134.845 120.385 ;
        RECT 135.490 119.755 135.820 120.555 ;
        RECT 136.120 119.585 136.450 120.385 ;
        RECT 136.620 119.755 136.950 120.555 ;
        RECT 137.530 120.555 139.965 120.725 ;
        RECT 137.530 119.755 137.860 120.555 ;
        RECT 138.030 119.585 138.360 120.385 ;
        RECT 138.660 119.755 138.990 120.555 ;
        RECT 139.635 119.585 139.885 120.385 ;
        RECT 140.155 119.585 140.325 120.725 ;
        RECT 140.495 119.755 140.835 120.725 ;
        RECT 141.005 121.395 141.390 121.965 ;
        RECT 141.560 121.675 141.885 122.135 ;
        RECT 142.405 121.505 142.685 121.965 ;
        RECT 141.005 120.725 141.285 121.395 ;
        RECT 141.560 121.335 142.685 121.505 ;
        RECT 141.560 121.225 142.010 121.335 ;
        RECT 141.455 120.895 142.010 121.225 ;
        RECT 142.875 121.165 143.275 121.965 ;
        RECT 143.675 121.675 143.945 122.135 ;
        RECT 144.115 121.505 144.400 121.965 ;
        RECT 141.005 119.755 141.390 120.725 ;
        RECT 141.560 120.435 142.010 120.895 ;
        RECT 142.180 120.605 143.275 121.165 ;
        RECT 141.560 120.215 142.685 120.435 ;
        RECT 141.560 119.585 141.885 120.045 ;
        RECT 142.405 119.755 142.685 120.215 ;
        RECT 142.875 119.755 143.275 120.605 ;
        RECT 143.445 121.335 144.400 121.505 ;
        RECT 144.685 121.395 145.070 121.965 ;
        RECT 145.240 121.675 145.565 122.135 ;
        RECT 146.085 121.505 146.365 121.965 ;
        RECT 143.445 120.435 143.655 121.335 ;
        RECT 143.825 120.605 144.515 121.165 ;
        RECT 144.685 120.725 144.965 121.395 ;
        RECT 145.240 121.335 146.365 121.505 ;
        RECT 145.240 121.225 145.690 121.335 ;
        RECT 145.135 120.895 145.690 121.225 ;
        RECT 146.555 121.165 146.955 121.965 ;
        RECT 147.355 121.675 147.625 122.135 ;
        RECT 147.795 121.505 148.080 121.965 ;
        RECT 143.445 120.215 144.400 120.435 ;
        RECT 143.675 119.585 143.945 120.045 ;
        RECT 144.115 119.755 144.400 120.215 ;
        RECT 144.685 119.755 145.070 120.725 ;
        RECT 145.240 120.435 145.690 120.895 ;
        RECT 145.860 120.605 146.955 121.165 ;
        RECT 145.240 120.215 146.365 120.435 ;
        RECT 145.240 119.585 145.565 120.045 ;
        RECT 146.085 119.755 146.365 120.215 ;
        RECT 146.555 119.755 146.955 120.605 ;
        RECT 147.125 121.335 148.080 121.505 ;
        RECT 148.365 121.460 148.635 121.805 ;
        RECT 148.825 121.735 149.205 122.135 ;
        RECT 149.375 121.565 149.545 121.915 ;
        RECT 149.715 121.735 150.045 122.135 ;
        RECT 150.245 121.565 150.415 121.915 ;
        RECT 150.615 121.635 150.945 122.135 ;
        RECT 147.125 120.435 147.335 121.335 ;
        RECT 147.505 120.605 148.195 121.165 ;
        RECT 148.365 120.725 148.535 121.460 ;
        RECT 148.805 121.395 150.415 121.565 ;
        RECT 148.805 121.225 148.975 121.395 ;
        RECT 148.705 120.895 148.975 121.225 ;
        RECT 149.145 120.895 149.550 121.225 ;
        RECT 148.805 120.725 148.975 120.895 ;
        RECT 149.720 120.775 150.430 121.225 ;
        RECT 150.600 120.895 150.950 121.465 ;
        RECT 151.585 121.410 151.875 122.135 ;
        RECT 152.045 121.395 152.430 121.965 ;
        RECT 152.600 121.675 152.925 122.135 ;
        RECT 153.445 121.505 153.725 121.965 ;
        RECT 147.125 120.215 148.080 120.435 ;
        RECT 147.355 119.585 147.625 120.045 ;
        RECT 147.795 119.755 148.080 120.215 ;
        RECT 148.365 119.755 148.635 120.725 ;
        RECT 148.805 120.555 149.530 120.725 ;
        RECT 149.720 120.605 150.435 120.775 ;
        RECT 149.360 120.435 149.530 120.555 ;
        RECT 150.630 120.435 150.950 120.725 ;
        RECT 148.845 119.585 149.125 120.385 ;
        RECT 149.360 120.265 150.950 120.435 ;
        RECT 149.295 119.805 150.950 120.095 ;
        RECT 151.585 119.585 151.875 120.750 ;
        RECT 152.045 120.725 152.325 121.395 ;
        RECT 152.600 121.335 153.725 121.505 ;
        RECT 152.600 121.225 153.050 121.335 ;
        RECT 152.495 120.895 153.050 121.225 ;
        RECT 153.915 121.165 154.315 121.965 ;
        RECT 154.715 121.675 154.985 122.135 ;
        RECT 155.155 121.505 155.440 121.965 ;
        RECT 152.045 119.755 152.430 120.725 ;
        RECT 152.600 120.435 153.050 120.895 ;
        RECT 153.220 120.605 154.315 121.165 ;
        RECT 152.600 120.215 153.725 120.435 ;
        RECT 152.600 119.585 152.925 120.045 ;
        RECT 153.445 119.755 153.725 120.215 ;
        RECT 153.915 119.755 154.315 120.605 ;
        RECT 154.485 121.335 155.440 121.505 ;
        RECT 155.725 121.385 156.935 122.135 ;
        RECT 154.485 120.435 154.695 121.335 ;
        RECT 154.865 120.605 155.555 121.165 ;
        RECT 155.725 120.675 156.245 121.215 ;
        RECT 156.415 120.845 156.935 121.385 ;
        RECT 154.485 120.215 155.440 120.435 ;
        RECT 154.715 119.585 154.985 120.045 ;
        RECT 155.155 119.755 155.440 120.215 ;
        RECT 155.725 119.585 156.935 120.675 ;
        RECT 22.700 119.415 157.020 119.585 ;
        RECT 22.785 118.325 23.995 119.415 ;
        RECT 24.165 118.325 26.755 119.415 ;
        RECT 22.785 117.615 23.305 118.155 ;
        RECT 23.475 117.785 23.995 118.325 ;
        RECT 24.165 117.635 25.375 118.155 ;
        RECT 25.545 117.805 26.755 118.325 ;
        RECT 26.925 117.810 27.205 119.245 ;
        RECT 27.375 118.640 28.085 119.415 ;
        RECT 28.255 118.470 28.585 119.245 ;
        RECT 27.435 118.255 28.585 118.470 ;
        RECT 22.785 116.865 23.995 117.615 ;
        RECT 24.165 116.865 26.755 117.635 ;
        RECT 26.925 117.035 27.265 117.810 ;
        RECT 27.435 117.685 27.720 118.255 ;
        RECT 27.905 117.855 28.375 118.085 ;
        RECT 28.780 118.055 28.995 119.170 ;
        RECT 29.175 118.695 29.505 119.415 ;
        RECT 29.695 118.465 29.970 119.235 ;
        RECT 30.140 118.805 30.470 119.235 ;
        RECT 30.640 118.975 30.835 119.415 ;
        RECT 31.015 118.805 31.345 119.235 ;
        RECT 30.140 118.635 31.345 118.805 ;
        RECT 29.285 118.055 29.515 118.395 ;
        RECT 29.695 118.275 30.280 118.465 ;
        RECT 30.450 118.305 31.345 118.635 ;
        RECT 31.525 118.325 32.735 119.415 ;
        RECT 28.545 117.875 28.995 118.055 ;
        RECT 28.545 117.855 28.875 117.875 ;
        RECT 29.185 117.855 29.515 118.055 ;
        RECT 27.435 117.495 28.145 117.685 ;
        RECT 27.845 117.355 28.145 117.495 ;
        RECT 28.335 117.495 29.515 117.685 ;
        RECT 28.335 117.415 28.665 117.495 ;
        RECT 27.845 117.345 28.160 117.355 ;
        RECT 27.845 117.335 28.170 117.345 ;
        RECT 27.845 117.330 28.180 117.335 ;
        RECT 27.435 116.865 27.605 117.325 ;
        RECT 27.845 117.320 28.185 117.330 ;
        RECT 27.845 117.315 28.190 117.320 ;
        RECT 27.845 117.305 28.195 117.315 ;
        RECT 27.845 117.300 28.200 117.305 ;
        RECT 27.845 117.035 28.205 117.300 ;
        RECT 28.835 116.865 29.005 117.325 ;
        RECT 29.175 117.035 29.515 117.495 ;
        RECT 29.695 117.455 29.935 118.105 ;
        RECT 30.105 117.605 30.280 118.275 ;
        RECT 30.450 117.775 30.865 118.105 ;
        RECT 31.045 117.775 31.340 118.105 ;
        RECT 30.105 117.425 30.435 117.605 ;
        RECT 29.710 116.865 30.040 117.255 ;
        RECT 30.210 117.045 30.435 117.425 ;
        RECT 30.635 117.155 30.865 117.775 ;
        RECT 31.525 117.615 32.045 118.155 ;
        RECT 32.215 117.785 32.735 118.325 ;
        RECT 32.905 118.340 33.175 119.245 ;
        RECT 33.345 118.655 33.675 119.415 ;
        RECT 33.855 118.485 34.025 119.245 ;
        RECT 31.045 116.865 31.345 117.595 ;
        RECT 31.525 116.865 32.735 117.615 ;
        RECT 32.905 117.540 33.075 118.340 ;
        RECT 33.360 118.315 34.025 118.485 ;
        RECT 34.285 118.325 35.495 119.415 ;
        RECT 33.360 118.170 33.530 118.315 ;
        RECT 33.245 117.840 33.530 118.170 ;
        RECT 33.360 117.585 33.530 117.840 ;
        RECT 33.765 117.765 34.095 118.135 ;
        RECT 34.285 117.615 34.805 118.155 ;
        RECT 34.975 117.785 35.495 118.325 ;
        RECT 35.665 118.250 35.955 119.415 ;
        RECT 32.905 117.035 33.165 117.540 ;
        RECT 33.360 117.415 34.025 117.585 ;
        RECT 33.345 116.865 33.675 117.245 ;
        RECT 33.855 117.035 34.025 117.415 ;
        RECT 34.285 116.865 35.495 117.615 ;
        RECT 35.665 116.865 35.955 117.590 ;
        RECT 36.135 117.045 36.395 119.235 ;
        RECT 36.565 118.685 36.905 119.415 ;
        RECT 37.085 118.505 37.355 119.235 ;
        RECT 36.585 118.285 37.355 118.505 ;
        RECT 37.535 118.525 37.765 119.235 ;
        RECT 37.935 118.705 38.265 119.415 ;
        RECT 38.435 118.525 38.695 119.235 ;
        RECT 37.535 118.285 38.695 118.525 ;
        RECT 38.885 118.325 40.555 119.415 ;
        RECT 36.585 117.615 36.875 118.285 ;
        RECT 37.055 117.795 37.520 118.105 ;
        RECT 37.700 117.795 38.225 118.105 ;
        RECT 36.585 117.415 37.815 117.615 ;
        RECT 36.655 116.865 37.325 117.235 ;
        RECT 37.505 117.045 37.815 117.415 ;
        RECT 37.995 117.155 38.225 117.795 ;
        RECT 38.405 117.775 38.705 118.105 ;
        RECT 38.885 117.635 39.635 118.155 ;
        RECT 39.805 117.805 40.555 118.325 ;
        RECT 40.735 118.355 41.065 119.205 ;
        RECT 38.405 116.865 38.695 117.595 ;
        RECT 38.885 116.865 40.555 117.635 ;
        RECT 40.735 117.590 40.925 118.355 ;
        RECT 41.235 118.275 41.485 119.415 ;
        RECT 41.675 118.775 41.925 119.195 ;
        RECT 42.155 118.945 42.485 119.415 ;
        RECT 42.715 118.775 42.965 119.195 ;
        RECT 41.675 118.605 42.965 118.775 ;
        RECT 43.145 118.775 43.475 119.205 ;
        RECT 43.945 118.905 45.605 119.195 ;
        RECT 43.145 118.605 43.600 118.775 ;
        RECT 41.665 118.105 41.880 118.435 ;
        RECT 41.095 117.775 41.405 118.105 ;
        RECT 41.575 117.775 41.880 118.105 ;
        RECT 42.055 117.775 42.340 118.435 ;
        RECT 42.535 117.775 42.800 118.435 ;
        RECT 43.015 117.775 43.260 118.435 ;
        RECT 41.235 117.605 41.405 117.775 ;
        RECT 43.430 117.605 43.600 118.605 ;
        RECT 43.945 118.565 45.540 118.735 ;
        RECT 45.775 118.615 46.055 119.415 ;
        RECT 43.945 118.275 44.270 118.565 ;
        RECT 45.370 118.445 45.540 118.565 ;
        RECT 44.465 118.225 45.180 118.395 ;
        RECT 45.370 118.275 46.095 118.445 ;
        RECT 46.265 118.275 46.540 119.245 ;
        RECT 40.735 117.080 41.065 117.590 ;
        RECT 41.235 117.435 43.600 117.605 ;
        RECT 43.945 117.535 44.300 118.105 ;
        RECT 44.470 117.775 45.180 118.225 ;
        RECT 45.925 118.105 46.095 118.275 ;
        RECT 45.350 117.775 45.755 118.105 ;
        RECT 45.925 117.775 46.200 118.105 ;
        RECT 45.925 117.605 46.095 117.775 ;
        RECT 44.485 117.435 46.095 117.605 ;
        RECT 46.370 117.540 46.540 118.275 ;
        RECT 46.710 118.235 46.880 119.415 ;
        RECT 47.740 118.785 48.025 119.245 ;
        RECT 48.195 118.955 48.465 119.415 ;
        RECT 47.740 118.565 48.695 118.785 ;
        RECT 47.625 117.835 48.315 118.395 ;
        RECT 41.235 116.865 41.565 117.265 ;
        RECT 42.615 117.095 42.945 117.435 ;
        RECT 43.115 116.865 43.445 117.265 ;
        RECT 43.950 116.865 44.285 117.365 ;
        RECT 44.485 117.085 44.655 117.435 ;
        RECT 44.855 116.865 45.185 117.265 ;
        RECT 45.355 117.085 45.525 117.435 ;
        RECT 45.695 116.865 46.075 117.265 ;
        RECT 46.265 117.195 46.540 117.540 ;
        RECT 46.710 116.865 46.880 117.780 ;
        RECT 48.485 117.665 48.695 118.565 ;
        RECT 47.740 117.495 48.695 117.665 ;
        RECT 48.865 118.395 49.265 119.245 ;
        RECT 49.455 118.785 49.735 119.245 ;
        RECT 50.255 118.955 50.580 119.415 ;
        RECT 49.455 118.565 50.580 118.785 ;
        RECT 48.865 117.835 49.960 118.395 ;
        RECT 50.130 118.105 50.580 118.565 ;
        RECT 50.750 118.275 51.135 119.245 ;
        RECT 51.965 118.745 52.245 119.415 ;
        RECT 52.415 118.525 52.715 119.075 ;
        RECT 52.915 118.695 53.245 119.415 ;
        RECT 53.435 118.695 53.895 119.245 ;
        RECT 47.740 117.035 48.025 117.495 ;
        RECT 48.195 116.865 48.465 117.325 ;
        RECT 48.865 117.035 49.265 117.835 ;
        RECT 50.130 117.775 50.685 118.105 ;
        RECT 50.130 117.665 50.580 117.775 ;
        RECT 49.455 117.495 50.580 117.665 ;
        RECT 50.855 117.605 51.135 118.275 ;
        RECT 51.780 118.105 52.045 118.465 ;
        RECT 52.415 118.355 53.355 118.525 ;
        RECT 53.185 118.105 53.355 118.355 ;
        RECT 51.780 117.855 52.455 118.105 ;
        RECT 52.675 117.855 53.015 118.105 ;
        RECT 53.185 117.775 53.475 118.105 ;
        RECT 53.185 117.685 53.355 117.775 ;
        RECT 49.455 117.035 49.735 117.495 ;
        RECT 50.255 116.865 50.580 117.325 ;
        RECT 50.750 117.035 51.135 117.605 ;
        RECT 51.965 117.495 53.355 117.685 ;
        RECT 51.965 117.135 52.295 117.495 ;
        RECT 53.645 117.325 53.895 118.695 ;
        RECT 54.070 118.275 54.390 119.415 ;
        RECT 54.570 118.105 54.765 119.155 ;
        RECT 54.945 118.565 55.275 119.245 ;
        RECT 55.475 118.615 55.730 119.415 ;
        RECT 55.905 118.980 61.250 119.415 ;
        RECT 54.945 118.285 55.295 118.565 ;
        RECT 54.130 118.055 54.390 118.105 ;
        RECT 54.125 117.885 54.390 118.055 ;
        RECT 54.130 117.775 54.390 117.885 ;
        RECT 54.570 117.775 54.955 118.105 ;
        RECT 55.125 117.905 55.295 118.285 ;
        RECT 55.485 118.075 55.730 118.435 ;
        RECT 55.125 117.735 55.645 117.905 ;
        RECT 52.915 116.865 53.165 117.325 ;
        RECT 53.335 117.035 53.895 117.325 ;
        RECT 54.070 117.395 55.285 117.565 ;
        RECT 54.070 117.045 54.360 117.395 ;
        RECT 54.555 116.865 54.885 117.225 ;
        RECT 55.055 117.090 55.285 117.395 ;
        RECT 55.475 117.375 55.645 117.735 ;
        RECT 57.490 117.410 57.830 118.240 ;
        RECT 59.310 117.730 59.660 118.980 ;
        RECT 61.425 118.250 61.715 119.415 ;
        RECT 61.885 118.325 63.555 119.415 ;
        RECT 63.725 118.860 64.330 119.415 ;
        RECT 64.505 118.905 64.985 119.245 ;
        RECT 65.155 118.870 65.410 119.415 ;
        RECT 63.725 118.760 64.340 118.860 ;
        RECT 64.155 118.735 64.340 118.760 ;
        RECT 61.885 117.635 62.635 118.155 ;
        RECT 62.805 117.805 63.555 118.325 ;
        RECT 63.725 118.140 63.985 118.590 ;
        RECT 64.155 118.490 64.485 118.735 ;
        RECT 64.655 118.415 65.410 118.665 ;
        RECT 65.580 118.545 65.855 119.245 ;
        RECT 64.640 118.380 65.410 118.415 ;
        RECT 64.625 118.370 65.410 118.380 ;
        RECT 64.620 118.355 65.515 118.370 ;
        RECT 64.600 118.340 65.515 118.355 ;
        RECT 64.580 118.330 65.515 118.340 ;
        RECT 64.555 118.320 65.515 118.330 ;
        RECT 64.485 118.290 65.515 118.320 ;
        RECT 64.465 118.260 65.515 118.290 ;
        RECT 64.445 118.230 65.515 118.260 ;
        RECT 64.415 118.205 65.515 118.230 ;
        RECT 64.380 118.170 65.515 118.205 ;
        RECT 64.350 118.165 65.515 118.170 ;
        RECT 64.350 118.160 64.740 118.165 ;
        RECT 64.350 118.150 64.715 118.160 ;
        RECT 64.350 118.145 64.700 118.150 ;
        RECT 64.350 118.140 64.685 118.145 ;
        RECT 63.725 118.135 64.685 118.140 ;
        RECT 63.725 118.125 64.675 118.135 ;
        RECT 63.725 118.120 64.665 118.125 ;
        RECT 63.725 118.110 64.655 118.120 ;
        RECT 63.725 118.100 64.650 118.110 ;
        RECT 63.725 118.095 64.645 118.100 ;
        RECT 63.725 118.080 64.635 118.095 ;
        RECT 63.725 118.065 64.630 118.080 ;
        RECT 63.725 118.040 64.620 118.065 ;
        RECT 63.725 117.970 64.615 118.040 ;
        RECT 55.475 117.205 55.675 117.375 ;
        RECT 55.475 117.170 55.645 117.205 ;
        RECT 55.905 116.865 61.250 117.410 ;
        RECT 61.425 116.865 61.715 117.590 ;
        RECT 61.885 116.865 63.555 117.635 ;
        RECT 63.725 117.415 64.275 117.800 ;
        RECT 64.445 117.245 64.615 117.970 ;
        RECT 63.725 117.075 64.615 117.245 ;
        RECT 64.785 117.570 65.115 117.995 ;
        RECT 65.285 117.770 65.515 118.165 ;
        RECT 64.785 117.085 65.005 117.570 ;
        RECT 65.685 117.515 65.855 118.545 ;
        RECT 65.175 116.865 65.425 117.405 ;
        RECT 65.595 117.035 65.855 117.515 ;
        RECT 66.025 118.275 66.410 119.245 ;
        RECT 66.580 118.955 66.905 119.415 ;
        RECT 67.425 118.785 67.705 119.245 ;
        RECT 66.580 118.565 67.705 118.785 ;
        RECT 66.025 117.605 66.305 118.275 ;
        RECT 66.580 118.105 67.030 118.565 ;
        RECT 67.895 118.395 68.295 119.245 ;
        RECT 68.695 118.955 68.965 119.415 ;
        RECT 69.135 118.785 69.420 119.245 ;
        RECT 66.475 117.775 67.030 118.105 ;
        RECT 67.200 117.835 68.295 118.395 ;
        RECT 66.580 117.665 67.030 117.775 ;
        RECT 66.025 117.035 66.410 117.605 ;
        RECT 66.580 117.495 67.705 117.665 ;
        RECT 66.580 116.865 66.905 117.325 ;
        RECT 67.425 117.035 67.705 117.495 ;
        RECT 67.895 117.035 68.295 117.835 ;
        RECT 68.465 118.565 69.420 118.785 ;
        RECT 68.465 117.665 68.675 118.565 ;
        RECT 69.725 118.525 69.985 119.235 ;
        RECT 70.155 118.705 70.485 119.415 ;
        RECT 70.655 118.525 70.885 119.235 ;
        RECT 68.845 117.835 69.535 118.395 ;
        RECT 69.725 118.285 70.885 118.525 ;
        RECT 71.065 118.505 71.335 119.235 ;
        RECT 71.515 118.685 71.855 119.415 ;
        RECT 71.065 118.285 71.835 118.505 ;
        RECT 69.715 117.775 70.015 118.105 ;
        RECT 70.195 117.795 70.720 118.105 ;
        RECT 70.900 117.795 71.365 118.105 ;
        RECT 68.465 117.495 69.420 117.665 ;
        RECT 68.695 116.865 68.965 117.325 ;
        RECT 69.135 117.035 69.420 117.495 ;
        RECT 69.725 116.865 70.015 117.595 ;
        RECT 70.195 117.155 70.425 117.795 ;
        RECT 71.545 117.615 71.835 118.285 ;
        RECT 70.605 117.415 71.835 117.615 ;
        RECT 70.605 117.045 70.915 117.415 ;
        RECT 71.095 116.865 71.765 117.235 ;
        RECT 72.025 117.045 72.285 119.235 ;
        RECT 72.465 118.545 72.740 119.245 ;
        RECT 72.910 118.870 73.165 119.415 ;
        RECT 73.335 118.905 73.815 119.245 ;
        RECT 73.990 118.860 74.595 119.415 ;
        RECT 73.980 118.760 74.595 118.860 ;
        RECT 73.980 118.735 74.165 118.760 ;
        RECT 72.465 117.515 72.635 118.545 ;
        RECT 72.910 118.415 73.665 118.665 ;
        RECT 73.835 118.490 74.165 118.735 ;
        RECT 75.775 118.745 75.945 119.245 ;
        RECT 76.115 118.915 76.445 119.415 ;
        RECT 72.910 118.380 73.680 118.415 ;
        RECT 72.910 118.370 73.695 118.380 ;
        RECT 72.805 118.355 73.700 118.370 ;
        RECT 72.805 118.340 73.720 118.355 ;
        RECT 72.805 118.330 73.740 118.340 ;
        RECT 72.805 118.320 73.765 118.330 ;
        RECT 72.805 118.290 73.835 118.320 ;
        RECT 72.805 118.260 73.855 118.290 ;
        RECT 72.805 118.230 73.875 118.260 ;
        RECT 72.805 118.205 73.905 118.230 ;
        RECT 72.805 118.170 73.940 118.205 ;
        RECT 72.805 118.165 73.970 118.170 ;
        RECT 72.805 117.770 73.035 118.165 ;
        RECT 73.580 118.160 73.970 118.165 ;
        RECT 73.605 118.150 73.970 118.160 ;
        RECT 73.620 118.145 73.970 118.150 ;
        RECT 73.635 118.140 73.970 118.145 ;
        RECT 74.335 118.140 74.595 118.590 ;
        RECT 75.775 118.575 76.440 118.745 ;
        RECT 73.635 118.135 74.595 118.140 ;
        RECT 73.645 118.125 74.595 118.135 ;
        RECT 73.655 118.120 74.595 118.125 ;
        RECT 73.665 118.110 74.595 118.120 ;
        RECT 73.670 118.100 74.595 118.110 ;
        RECT 73.675 118.095 74.595 118.100 ;
        RECT 73.685 118.080 74.595 118.095 ;
        RECT 73.690 118.065 74.595 118.080 ;
        RECT 73.700 118.040 74.595 118.065 ;
        RECT 73.205 117.570 73.535 117.995 ;
        RECT 72.465 117.035 72.725 117.515 ;
        RECT 72.895 116.865 73.145 117.405 ;
        RECT 73.315 117.085 73.535 117.570 ;
        RECT 73.705 117.970 74.595 118.040 ;
        RECT 73.705 117.245 73.875 117.970 ;
        RECT 74.045 117.415 74.595 117.800 ;
        RECT 75.690 117.755 76.040 118.405 ;
        RECT 76.210 117.585 76.440 118.575 ;
        RECT 75.775 117.415 76.440 117.585 ;
        RECT 73.705 117.075 74.595 117.245 ;
        RECT 75.775 117.125 75.945 117.415 ;
        RECT 76.115 116.865 76.445 117.245 ;
        RECT 76.615 117.125 76.800 119.245 ;
        RECT 77.040 118.955 77.305 119.415 ;
        RECT 77.475 118.820 77.725 119.245 ;
        RECT 77.935 118.970 79.040 119.140 ;
        RECT 77.420 118.690 77.725 118.820 ;
        RECT 76.970 117.495 77.250 118.445 ;
        RECT 77.420 117.585 77.590 118.690 ;
        RECT 77.760 117.905 78.000 118.500 ;
        RECT 78.170 118.435 78.700 118.800 ;
        RECT 78.170 117.735 78.340 118.435 ;
        RECT 78.870 118.355 79.040 118.970 ;
        RECT 79.210 118.615 79.380 119.415 ;
        RECT 79.550 118.915 79.800 119.245 ;
        RECT 80.025 118.945 80.910 119.115 ;
        RECT 78.870 118.265 79.380 118.355 ;
        RECT 77.420 117.455 77.645 117.585 ;
        RECT 77.815 117.515 78.340 117.735 ;
        RECT 78.510 118.095 79.380 118.265 ;
        RECT 77.055 116.865 77.305 117.325 ;
        RECT 77.475 117.315 77.645 117.455 ;
        RECT 78.510 117.315 78.680 118.095 ;
        RECT 79.210 118.025 79.380 118.095 ;
        RECT 78.890 117.845 79.090 117.875 ;
        RECT 79.550 117.845 79.720 118.915 ;
        RECT 79.890 118.025 80.080 118.745 ;
        RECT 78.890 117.545 79.720 117.845 ;
        RECT 80.250 117.815 80.570 118.775 ;
        RECT 77.475 117.145 77.810 117.315 ;
        RECT 78.005 117.145 78.680 117.315 ;
        RECT 79.000 116.865 79.370 117.365 ;
        RECT 79.550 117.315 79.720 117.545 ;
        RECT 80.105 117.485 80.570 117.815 ;
        RECT 80.740 118.105 80.910 118.945 ;
        RECT 81.090 118.915 81.405 119.415 ;
        RECT 81.635 118.685 81.975 119.245 ;
        RECT 81.080 118.310 81.975 118.685 ;
        RECT 82.145 118.405 82.315 119.415 ;
        RECT 81.785 118.105 81.975 118.310 ;
        RECT 82.485 118.355 82.815 119.200 ;
        RECT 83.045 118.545 83.320 119.245 ;
        RECT 83.490 118.870 83.745 119.415 ;
        RECT 83.915 118.905 84.395 119.245 ;
        RECT 84.570 118.860 85.175 119.415 ;
        RECT 84.560 118.760 85.175 118.860 ;
        RECT 84.560 118.735 84.745 118.760 ;
        RECT 82.485 118.275 82.875 118.355 ;
        RECT 82.660 118.225 82.875 118.275 ;
        RECT 80.740 117.775 81.615 118.105 ;
        RECT 81.785 117.775 82.535 118.105 ;
        RECT 80.740 117.315 80.910 117.775 ;
        RECT 81.785 117.605 81.985 117.775 ;
        RECT 82.705 117.645 82.875 118.225 ;
        RECT 82.650 117.605 82.875 117.645 ;
        RECT 79.550 117.145 79.955 117.315 ;
        RECT 80.125 117.145 80.910 117.315 ;
        RECT 81.185 116.865 81.395 117.395 ;
        RECT 81.655 117.080 81.985 117.605 ;
        RECT 82.495 117.520 82.875 117.605 ;
        RECT 82.155 116.865 82.325 117.475 ;
        RECT 82.495 117.085 82.825 117.520 ;
        RECT 83.045 117.515 83.215 118.545 ;
        RECT 83.490 118.415 84.245 118.665 ;
        RECT 84.415 118.490 84.745 118.735 ;
        RECT 83.490 118.380 84.260 118.415 ;
        RECT 83.490 118.370 84.275 118.380 ;
        RECT 83.385 118.355 84.280 118.370 ;
        RECT 83.385 118.340 84.300 118.355 ;
        RECT 83.385 118.330 84.320 118.340 ;
        RECT 83.385 118.320 84.345 118.330 ;
        RECT 83.385 118.290 84.415 118.320 ;
        RECT 83.385 118.260 84.435 118.290 ;
        RECT 83.385 118.230 84.455 118.260 ;
        RECT 83.385 118.205 84.485 118.230 ;
        RECT 83.385 118.170 84.520 118.205 ;
        RECT 83.385 118.165 84.550 118.170 ;
        RECT 83.385 117.770 83.615 118.165 ;
        RECT 84.160 118.160 84.550 118.165 ;
        RECT 84.185 118.150 84.550 118.160 ;
        RECT 84.200 118.145 84.550 118.150 ;
        RECT 84.215 118.140 84.550 118.145 ;
        RECT 84.915 118.140 85.175 118.590 ;
        RECT 85.355 118.445 85.685 119.230 ;
        RECT 85.355 118.275 86.035 118.445 ;
        RECT 86.215 118.275 86.545 119.415 ;
        RECT 84.215 118.135 85.175 118.140 ;
        RECT 84.225 118.125 85.175 118.135 ;
        RECT 84.235 118.120 85.175 118.125 ;
        RECT 84.245 118.110 85.175 118.120 ;
        RECT 84.250 118.100 85.175 118.110 ;
        RECT 84.255 118.095 85.175 118.100 ;
        RECT 84.265 118.080 85.175 118.095 ;
        RECT 84.270 118.065 85.175 118.080 ;
        RECT 84.280 118.040 85.175 118.065 ;
        RECT 83.785 117.570 84.115 117.995 ;
        RECT 83.865 117.545 84.115 117.570 ;
        RECT 83.045 117.035 83.305 117.515 ;
        RECT 83.475 116.865 83.725 117.405 ;
        RECT 83.895 117.085 84.115 117.545 ;
        RECT 84.285 117.970 85.175 118.040 ;
        RECT 84.285 117.245 84.455 117.970 ;
        RECT 85.345 117.855 85.695 118.105 ;
        RECT 84.625 117.415 85.175 117.800 ;
        RECT 85.865 117.675 86.035 118.275 ;
        RECT 87.185 118.250 87.475 119.415 ;
        RECT 87.735 118.745 87.905 119.245 ;
        RECT 88.075 118.915 88.405 119.415 ;
        RECT 87.735 118.575 88.400 118.745 ;
        RECT 86.205 117.855 86.555 118.105 ;
        RECT 87.650 117.755 88.000 118.405 ;
        RECT 84.285 117.075 85.175 117.245 ;
        RECT 85.365 116.865 85.605 117.675 ;
        RECT 85.775 117.035 86.105 117.675 ;
        RECT 86.275 116.865 86.545 117.675 ;
        RECT 87.185 116.865 87.475 117.590 ;
        RECT 88.170 117.585 88.400 118.575 ;
        RECT 87.735 117.415 88.400 117.585 ;
        RECT 87.735 117.125 87.905 117.415 ;
        RECT 88.075 116.865 88.405 117.245 ;
        RECT 88.575 117.125 88.760 119.245 ;
        RECT 89.000 118.955 89.265 119.415 ;
        RECT 89.435 118.820 89.685 119.245 ;
        RECT 89.895 118.970 91.000 119.140 ;
        RECT 89.380 118.690 89.685 118.820 ;
        RECT 88.930 117.495 89.210 118.445 ;
        RECT 89.380 117.585 89.550 118.690 ;
        RECT 89.720 117.905 89.960 118.500 ;
        RECT 90.130 118.435 90.660 118.800 ;
        RECT 90.130 117.735 90.300 118.435 ;
        RECT 90.830 118.355 91.000 118.970 ;
        RECT 91.170 118.615 91.340 119.415 ;
        RECT 91.510 118.915 91.760 119.245 ;
        RECT 91.985 118.945 92.870 119.115 ;
        RECT 90.830 118.265 91.340 118.355 ;
        RECT 89.380 117.455 89.605 117.585 ;
        RECT 89.775 117.515 90.300 117.735 ;
        RECT 90.470 118.095 91.340 118.265 ;
        RECT 89.015 116.865 89.265 117.325 ;
        RECT 89.435 117.315 89.605 117.455 ;
        RECT 90.470 117.315 90.640 118.095 ;
        RECT 91.170 118.025 91.340 118.095 ;
        RECT 90.850 117.845 91.050 117.875 ;
        RECT 91.510 117.845 91.680 118.915 ;
        RECT 91.850 118.025 92.040 118.745 ;
        RECT 90.850 117.545 91.680 117.845 ;
        RECT 92.210 117.815 92.530 118.775 ;
        RECT 89.435 117.145 89.770 117.315 ;
        RECT 89.965 117.145 90.640 117.315 ;
        RECT 90.960 116.865 91.330 117.365 ;
        RECT 91.510 117.315 91.680 117.545 ;
        RECT 92.065 117.485 92.530 117.815 ;
        RECT 92.700 118.105 92.870 118.945 ;
        RECT 93.050 118.915 93.365 119.415 ;
        RECT 93.595 118.685 93.935 119.245 ;
        RECT 93.040 118.310 93.935 118.685 ;
        RECT 94.105 118.405 94.275 119.415 ;
        RECT 93.745 118.105 93.935 118.310 ;
        RECT 94.445 118.355 94.775 119.200 ;
        RECT 96.015 118.745 96.185 119.245 ;
        RECT 96.355 118.915 96.685 119.415 ;
        RECT 96.015 118.575 96.680 118.745 ;
        RECT 94.445 118.275 94.835 118.355 ;
        RECT 94.620 118.225 94.835 118.275 ;
        RECT 92.700 117.775 93.575 118.105 ;
        RECT 93.745 117.775 94.495 118.105 ;
        RECT 92.700 117.315 92.870 117.775 ;
        RECT 93.745 117.605 93.945 117.775 ;
        RECT 94.665 117.645 94.835 118.225 ;
        RECT 95.930 117.755 96.280 118.405 ;
        RECT 94.610 117.605 94.835 117.645 ;
        RECT 91.510 117.145 91.915 117.315 ;
        RECT 92.085 117.145 92.870 117.315 ;
        RECT 93.145 116.865 93.355 117.395 ;
        RECT 93.615 117.080 93.945 117.605 ;
        RECT 94.455 117.520 94.835 117.605 ;
        RECT 96.450 117.585 96.680 118.575 ;
        RECT 94.115 116.865 94.285 117.475 ;
        RECT 94.455 117.085 94.785 117.520 ;
        RECT 96.015 117.415 96.680 117.585 ;
        RECT 96.015 117.125 96.185 117.415 ;
        RECT 96.355 116.865 96.685 117.245 ;
        RECT 96.855 117.125 97.040 119.245 ;
        RECT 97.280 118.955 97.545 119.415 ;
        RECT 97.715 118.820 97.965 119.245 ;
        RECT 98.175 118.970 99.280 119.140 ;
        RECT 97.660 118.690 97.965 118.820 ;
        RECT 97.210 117.495 97.490 118.445 ;
        RECT 97.660 117.585 97.830 118.690 ;
        RECT 98.000 117.905 98.240 118.500 ;
        RECT 98.410 118.435 98.940 118.800 ;
        RECT 98.410 117.735 98.580 118.435 ;
        RECT 99.110 118.355 99.280 118.970 ;
        RECT 99.450 118.615 99.620 119.415 ;
        RECT 99.790 118.915 100.040 119.245 ;
        RECT 100.265 118.945 101.150 119.115 ;
        RECT 99.110 118.265 99.620 118.355 ;
        RECT 97.660 117.455 97.885 117.585 ;
        RECT 98.055 117.515 98.580 117.735 ;
        RECT 98.750 118.095 99.620 118.265 ;
        RECT 97.295 116.865 97.545 117.325 ;
        RECT 97.715 117.315 97.885 117.455 ;
        RECT 98.750 117.315 98.920 118.095 ;
        RECT 99.450 118.025 99.620 118.095 ;
        RECT 99.130 117.845 99.330 117.875 ;
        RECT 99.790 117.845 99.960 118.915 ;
        RECT 100.130 118.025 100.320 118.745 ;
        RECT 99.130 117.545 99.960 117.845 ;
        RECT 100.490 117.815 100.810 118.775 ;
        RECT 97.715 117.145 98.050 117.315 ;
        RECT 98.245 117.145 98.920 117.315 ;
        RECT 99.240 116.865 99.610 117.365 ;
        RECT 99.790 117.315 99.960 117.545 ;
        RECT 100.345 117.485 100.810 117.815 ;
        RECT 100.980 118.105 101.150 118.945 ;
        RECT 101.330 118.915 101.645 119.415 ;
        RECT 101.875 118.685 102.215 119.245 ;
        RECT 101.320 118.310 102.215 118.685 ;
        RECT 102.385 118.405 102.555 119.415 ;
        RECT 102.025 118.105 102.215 118.310 ;
        RECT 102.725 118.355 103.055 119.200 ;
        RECT 102.725 118.275 103.115 118.355 ;
        RECT 103.285 118.325 106.795 119.415 ;
        RECT 102.900 118.225 103.115 118.275 ;
        RECT 100.980 117.775 101.855 118.105 ;
        RECT 102.025 117.775 102.775 118.105 ;
        RECT 100.980 117.315 101.150 117.775 ;
        RECT 102.025 117.605 102.225 117.775 ;
        RECT 102.945 117.645 103.115 118.225 ;
        RECT 102.890 117.605 103.115 117.645 ;
        RECT 99.790 117.145 100.195 117.315 ;
        RECT 100.365 117.145 101.150 117.315 ;
        RECT 101.425 116.865 101.635 117.395 ;
        RECT 101.895 117.080 102.225 117.605 ;
        RECT 102.735 117.520 103.115 117.605 ;
        RECT 103.285 117.635 104.935 118.155 ;
        RECT 105.105 117.805 106.795 118.325 ;
        RECT 106.965 118.305 107.225 119.245 ;
        RECT 107.395 119.015 107.725 119.415 ;
        RECT 108.870 119.150 109.125 119.245 ;
        RECT 107.985 118.980 109.125 119.150 ;
        RECT 109.295 119.035 109.625 119.205 ;
        RECT 107.985 118.755 108.155 118.980 ;
        RECT 107.395 118.585 108.155 118.755 ;
        RECT 108.870 118.845 109.125 118.980 ;
        RECT 102.395 116.865 102.565 117.475 ;
        RECT 102.735 117.085 103.065 117.520 ;
        RECT 103.285 116.865 106.795 117.635 ;
        RECT 106.965 117.590 107.140 118.305 ;
        RECT 107.395 118.105 107.565 118.585 ;
        RECT 108.420 118.495 108.590 118.685 ;
        RECT 108.870 118.675 109.280 118.845 ;
        RECT 107.310 117.775 107.565 118.105 ;
        RECT 107.790 117.775 108.120 118.395 ;
        RECT 108.420 118.325 108.940 118.495 ;
        RECT 108.290 117.775 108.580 118.155 ;
        RECT 108.770 117.605 108.940 118.325 ;
        RECT 106.965 117.035 107.225 117.590 ;
        RECT 108.060 117.435 108.940 117.605 ;
        RECT 109.110 117.650 109.280 118.675 ;
        RECT 109.455 118.785 109.625 119.035 ;
        RECT 109.795 118.955 110.045 119.415 ;
        RECT 110.215 118.785 110.395 119.245 ;
        RECT 109.455 118.615 110.395 118.785 ;
        RECT 109.480 118.135 109.960 118.435 ;
        RECT 109.110 117.480 109.460 117.650 ;
        RECT 109.700 117.545 109.960 118.135 ;
        RECT 110.160 117.545 110.420 118.435 ;
        RECT 111.625 118.275 111.835 119.415 ;
        RECT 112.005 118.265 112.335 119.245 ;
        RECT 112.505 118.275 112.735 119.415 ;
        RECT 107.395 116.865 107.825 117.310 ;
        RECT 108.060 117.035 108.230 117.435 ;
        RECT 108.400 116.865 109.120 117.265 ;
        RECT 109.290 117.035 109.460 117.480 ;
        RECT 110.035 116.865 110.435 117.375 ;
        RECT 111.625 116.865 111.835 117.685 ;
        RECT 112.005 117.665 112.255 118.265 ;
        RECT 112.945 118.250 113.235 119.415 ;
        RECT 113.495 118.745 113.665 119.245 ;
        RECT 113.835 118.915 114.165 119.415 ;
        RECT 113.495 118.575 114.160 118.745 ;
        RECT 112.425 117.855 112.755 118.105 ;
        RECT 113.410 117.755 113.760 118.405 ;
        RECT 112.005 117.035 112.335 117.665 ;
        RECT 112.505 116.865 112.735 117.685 ;
        RECT 112.945 116.865 113.235 117.590 ;
        RECT 113.930 117.585 114.160 118.575 ;
        RECT 113.495 117.415 114.160 117.585 ;
        RECT 113.495 117.125 113.665 117.415 ;
        RECT 113.835 116.865 114.165 117.245 ;
        RECT 114.335 117.125 114.520 119.245 ;
        RECT 114.760 118.955 115.025 119.415 ;
        RECT 115.195 118.820 115.445 119.245 ;
        RECT 115.655 118.970 116.760 119.140 ;
        RECT 115.140 118.690 115.445 118.820 ;
        RECT 114.690 117.495 114.970 118.445 ;
        RECT 115.140 117.585 115.310 118.690 ;
        RECT 115.480 117.905 115.720 118.500 ;
        RECT 115.890 118.435 116.420 118.800 ;
        RECT 115.890 117.735 116.060 118.435 ;
        RECT 116.590 118.355 116.760 118.970 ;
        RECT 116.930 118.615 117.100 119.415 ;
        RECT 117.270 118.915 117.520 119.245 ;
        RECT 117.745 118.945 118.630 119.115 ;
        RECT 116.590 118.265 117.100 118.355 ;
        RECT 115.140 117.455 115.365 117.585 ;
        RECT 115.535 117.515 116.060 117.735 ;
        RECT 116.230 118.095 117.100 118.265 ;
        RECT 114.775 116.865 115.025 117.325 ;
        RECT 115.195 117.315 115.365 117.455 ;
        RECT 116.230 117.315 116.400 118.095 ;
        RECT 116.930 118.025 117.100 118.095 ;
        RECT 116.610 117.845 116.810 117.875 ;
        RECT 117.270 117.845 117.440 118.915 ;
        RECT 117.610 118.025 117.800 118.745 ;
        RECT 116.610 117.545 117.440 117.845 ;
        RECT 117.970 117.815 118.290 118.775 ;
        RECT 115.195 117.145 115.530 117.315 ;
        RECT 115.725 117.145 116.400 117.315 ;
        RECT 116.720 116.865 117.090 117.365 ;
        RECT 117.270 117.315 117.440 117.545 ;
        RECT 117.825 117.485 118.290 117.815 ;
        RECT 118.460 118.105 118.630 118.945 ;
        RECT 118.810 118.915 119.125 119.415 ;
        RECT 119.355 118.685 119.695 119.245 ;
        RECT 118.800 118.310 119.695 118.685 ;
        RECT 119.865 118.405 120.035 119.415 ;
        RECT 119.505 118.105 119.695 118.310 ;
        RECT 120.205 118.355 120.535 119.200 ;
        RECT 120.205 118.275 120.595 118.355 ;
        RECT 120.775 118.275 121.105 119.415 ;
        RECT 121.635 118.445 121.965 119.230 ;
        RECT 121.285 118.275 121.965 118.445 ;
        RECT 122.145 118.325 123.355 119.415 ;
        RECT 123.615 118.745 123.785 119.245 ;
        RECT 123.955 118.915 124.285 119.415 ;
        RECT 123.615 118.575 124.280 118.745 ;
        RECT 120.380 118.225 120.595 118.275 ;
        RECT 118.460 117.775 119.335 118.105 ;
        RECT 119.505 117.775 120.255 118.105 ;
        RECT 118.460 117.315 118.630 117.775 ;
        RECT 119.505 117.605 119.705 117.775 ;
        RECT 120.425 117.645 120.595 118.225 ;
        RECT 120.765 117.855 121.115 118.105 ;
        RECT 121.285 117.675 121.455 118.275 ;
        RECT 121.625 117.855 121.975 118.105 ;
        RECT 120.370 117.605 120.595 117.645 ;
        RECT 117.270 117.145 117.675 117.315 ;
        RECT 117.845 117.145 118.630 117.315 ;
        RECT 118.905 116.865 119.115 117.395 ;
        RECT 119.375 117.080 119.705 117.605 ;
        RECT 120.215 117.520 120.595 117.605 ;
        RECT 119.875 116.865 120.045 117.475 ;
        RECT 120.215 117.085 120.545 117.520 ;
        RECT 120.775 116.865 121.045 117.675 ;
        RECT 121.215 117.035 121.545 117.675 ;
        RECT 121.715 116.865 121.955 117.675 ;
        RECT 122.145 117.615 122.665 118.155 ;
        RECT 122.835 117.785 123.355 118.325 ;
        RECT 123.530 117.755 123.880 118.405 ;
        RECT 122.145 116.865 123.355 117.615 ;
        RECT 124.050 117.585 124.280 118.575 ;
        RECT 123.615 117.415 124.280 117.585 ;
        RECT 123.615 117.125 123.785 117.415 ;
        RECT 123.955 116.865 124.285 117.245 ;
        RECT 124.455 117.125 124.640 119.245 ;
        RECT 124.880 118.955 125.145 119.415 ;
        RECT 125.315 118.820 125.565 119.245 ;
        RECT 125.775 118.970 126.880 119.140 ;
        RECT 125.260 118.690 125.565 118.820 ;
        RECT 124.810 117.495 125.090 118.445 ;
        RECT 125.260 117.585 125.430 118.690 ;
        RECT 125.600 117.905 125.840 118.500 ;
        RECT 126.010 118.435 126.540 118.800 ;
        RECT 126.010 117.735 126.180 118.435 ;
        RECT 126.710 118.355 126.880 118.970 ;
        RECT 127.050 118.615 127.220 119.415 ;
        RECT 127.390 118.915 127.640 119.245 ;
        RECT 127.865 118.945 128.750 119.115 ;
        RECT 126.710 118.265 127.220 118.355 ;
        RECT 125.260 117.455 125.485 117.585 ;
        RECT 125.655 117.515 126.180 117.735 ;
        RECT 126.350 118.095 127.220 118.265 ;
        RECT 124.895 116.865 125.145 117.325 ;
        RECT 125.315 117.315 125.485 117.455 ;
        RECT 126.350 117.315 126.520 118.095 ;
        RECT 127.050 118.025 127.220 118.095 ;
        RECT 126.730 117.845 126.930 117.875 ;
        RECT 127.390 117.845 127.560 118.915 ;
        RECT 127.730 118.025 127.920 118.745 ;
        RECT 126.730 117.545 127.560 117.845 ;
        RECT 128.090 117.815 128.410 118.775 ;
        RECT 125.315 117.145 125.650 117.315 ;
        RECT 125.845 117.145 126.520 117.315 ;
        RECT 126.840 116.865 127.210 117.365 ;
        RECT 127.390 117.315 127.560 117.545 ;
        RECT 127.945 117.485 128.410 117.815 ;
        RECT 128.580 118.105 128.750 118.945 ;
        RECT 128.930 118.915 129.245 119.415 ;
        RECT 129.475 118.685 129.815 119.245 ;
        RECT 128.920 118.310 129.815 118.685 ;
        RECT 129.985 118.405 130.155 119.415 ;
        RECT 129.625 118.105 129.815 118.310 ;
        RECT 130.325 118.355 130.655 119.200 ;
        RECT 130.325 118.275 130.715 118.355 ;
        RECT 130.500 118.225 130.715 118.275 ;
        RECT 128.580 117.775 129.455 118.105 ;
        RECT 129.625 117.775 130.375 118.105 ;
        RECT 128.580 117.315 128.750 117.775 ;
        RECT 129.625 117.605 129.825 117.775 ;
        RECT 130.545 117.645 130.715 118.225 ;
        RECT 130.490 117.605 130.715 117.645 ;
        RECT 127.390 117.145 127.795 117.315 ;
        RECT 127.965 117.145 128.750 117.315 ;
        RECT 129.025 116.865 129.235 117.395 ;
        RECT 129.495 117.080 129.825 117.605 ;
        RECT 130.335 117.520 130.715 117.605 ;
        RECT 129.995 116.865 130.165 117.475 ;
        RECT 130.335 117.085 130.665 117.520 ;
        RECT 130.895 117.035 131.155 119.245 ;
        RECT 131.325 118.615 132.135 119.415 ;
        RECT 132.305 118.445 132.635 119.245 ;
        RECT 132.820 118.615 133.560 119.415 ;
        RECT 133.730 118.445 133.980 119.245 ;
        RECT 131.495 118.275 133.980 118.445 ;
        RECT 131.495 118.105 131.665 118.275 ;
        RECT 134.150 118.105 134.335 119.195 ;
        RECT 134.530 118.615 134.855 119.415 ;
        RECT 131.325 117.775 131.665 118.105 ;
        RECT 132.065 117.855 132.545 118.105 ;
        RECT 131.495 117.685 131.665 117.775 ;
        RECT 131.495 117.515 132.165 117.685 ;
        RECT 131.335 116.865 131.645 117.345 ;
        RECT 131.825 117.035 132.165 117.515 ;
        RECT 132.335 117.170 132.545 117.855 ;
        RECT 132.725 117.170 132.995 118.105 ;
        RECT 133.245 117.775 133.505 118.105 ;
        RECT 133.850 117.855 134.335 118.105 ;
        RECT 134.505 117.855 134.835 118.440 ;
        RECT 135.025 118.275 135.410 119.245 ;
        RECT 135.580 118.955 135.905 119.415 ;
        RECT 136.425 118.785 136.705 119.245 ;
        RECT 135.580 118.565 136.705 118.785 ;
        RECT 133.245 117.170 133.490 117.775 ;
        RECT 133.670 117.485 134.855 117.655 ;
        RECT 133.670 117.035 133.960 117.485 ;
        RECT 134.130 116.865 134.420 117.315 ;
        RECT 134.590 117.035 134.855 117.485 ;
        RECT 135.025 117.605 135.305 118.275 ;
        RECT 135.580 118.105 136.030 118.565 ;
        RECT 136.895 118.395 137.295 119.245 ;
        RECT 137.695 118.955 137.965 119.415 ;
        RECT 138.135 118.785 138.420 119.245 ;
        RECT 135.475 117.775 136.030 118.105 ;
        RECT 136.200 117.835 137.295 118.395 ;
        RECT 135.580 117.665 136.030 117.775 ;
        RECT 135.025 117.035 135.410 117.605 ;
        RECT 135.580 117.495 136.705 117.665 ;
        RECT 135.580 116.865 135.905 117.325 ;
        RECT 136.425 117.035 136.705 117.495 ;
        RECT 136.895 117.035 137.295 117.835 ;
        RECT 137.465 118.565 138.420 118.785 ;
        RECT 137.465 117.665 137.675 118.565 ;
        RECT 137.845 117.835 138.535 118.395 ;
        RECT 138.705 118.250 138.995 119.415 ;
        RECT 139.225 118.355 139.555 119.200 ;
        RECT 139.725 118.405 139.895 119.415 ;
        RECT 140.065 118.685 140.405 119.245 ;
        RECT 140.635 118.915 140.950 119.415 ;
        RECT 141.130 118.945 142.015 119.115 ;
        RECT 139.165 118.275 139.555 118.355 ;
        RECT 140.065 118.310 140.960 118.685 ;
        RECT 139.165 118.225 139.380 118.275 ;
        RECT 137.465 117.495 138.420 117.665 ;
        RECT 139.165 117.645 139.335 118.225 ;
        RECT 140.065 118.105 140.255 118.310 ;
        RECT 141.130 118.105 141.300 118.945 ;
        RECT 142.240 118.915 142.490 119.245 ;
        RECT 139.505 117.775 140.255 118.105 ;
        RECT 140.425 117.775 141.300 118.105 ;
        RECT 139.165 117.605 139.390 117.645 ;
        RECT 140.055 117.605 140.255 117.775 ;
        RECT 137.695 116.865 137.965 117.325 ;
        RECT 138.135 117.035 138.420 117.495 ;
        RECT 138.705 116.865 138.995 117.590 ;
        RECT 139.165 117.520 139.545 117.605 ;
        RECT 139.215 117.085 139.545 117.520 ;
        RECT 139.715 116.865 139.885 117.475 ;
        RECT 140.055 117.080 140.385 117.605 ;
        RECT 140.645 116.865 140.855 117.395 ;
        RECT 141.130 117.315 141.300 117.775 ;
        RECT 141.470 117.815 141.790 118.775 ;
        RECT 141.960 118.025 142.150 118.745 ;
        RECT 142.320 117.845 142.490 118.915 ;
        RECT 142.660 118.615 142.830 119.415 ;
        RECT 143.000 118.970 144.105 119.140 ;
        RECT 143.000 118.355 143.170 118.970 ;
        RECT 144.315 118.820 144.565 119.245 ;
        RECT 144.735 118.955 145.000 119.415 ;
        RECT 143.340 118.435 143.870 118.800 ;
        RECT 144.315 118.690 144.620 118.820 ;
        RECT 142.660 118.265 143.170 118.355 ;
        RECT 142.660 118.095 143.530 118.265 ;
        RECT 142.660 118.025 142.830 118.095 ;
        RECT 142.950 117.845 143.150 117.875 ;
        RECT 141.470 117.485 141.935 117.815 ;
        RECT 142.320 117.545 143.150 117.845 ;
        RECT 142.320 117.315 142.490 117.545 ;
        RECT 141.130 117.145 141.915 117.315 ;
        RECT 142.085 117.145 142.490 117.315 ;
        RECT 142.670 116.865 143.040 117.365 ;
        RECT 143.360 117.315 143.530 118.095 ;
        RECT 143.700 117.735 143.870 118.435 ;
        RECT 144.040 117.905 144.280 118.500 ;
        RECT 143.700 117.515 144.225 117.735 ;
        RECT 144.450 117.585 144.620 118.690 ;
        RECT 144.395 117.455 144.620 117.585 ;
        RECT 144.790 117.495 145.070 118.445 ;
        RECT 144.395 117.315 144.565 117.455 ;
        RECT 143.360 117.145 144.035 117.315 ;
        RECT 144.230 117.145 144.565 117.315 ;
        RECT 144.735 116.865 144.985 117.325 ;
        RECT 145.240 117.125 145.425 119.245 ;
        RECT 145.595 118.915 145.925 119.415 ;
        RECT 146.095 118.745 146.265 119.245 ;
        RECT 145.600 118.575 146.265 118.745 ;
        RECT 145.600 117.585 145.830 118.575 ;
        RECT 146.000 117.755 146.350 118.405 ;
        RECT 146.525 118.325 148.195 119.415 ;
        RECT 148.455 118.745 148.625 119.245 ;
        RECT 148.795 118.915 149.125 119.415 ;
        RECT 148.455 118.575 149.120 118.745 ;
        RECT 146.525 117.635 147.275 118.155 ;
        RECT 147.445 117.805 148.195 118.325 ;
        RECT 148.370 117.755 148.720 118.405 ;
        RECT 145.600 117.415 146.265 117.585 ;
        RECT 145.595 116.865 145.925 117.245 ;
        RECT 146.095 117.125 146.265 117.415 ;
        RECT 146.525 116.865 148.195 117.635 ;
        RECT 148.890 117.585 149.120 118.575 ;
        RECT 148.455 117.415 149.120 117.585 ;
        RECT 148.455 117.125 148.625 117.415 ;
        RECT 148.795 116.865 149.125 117.245 ;
        RECT 149.295 117.125 149.480 119.245 ;
        RECT 149.720 118.955 149.985 119.415 ;
        RECT 150.155 118.820 150.405 119.245 ;
        RECT 150.615 118.970 151.720 119.140 ;
        RECT 150.100 118.690 150.405 118.820 ;
        RECT 149.650 117.495 149.930 118.445 ;
        RECT 150.100 117.585 150.270 118.690 ;
        RECT 150.440 117.905 150.680 118.500 ;
        RECT 150.850 118.435 151.380 118.800 ;
        RECT 150.850 117.735 151.020 118.435 ;
        RECT 151.550 118.355 151.720 118.970 ;
        RECT 151.890 118.615 152.060 119.415 ;
        RECT 152.230 118.915 152.480 119.245 ;
        RECT 152.705 118.945 153.590 119.115 ;
        RECT 151.550 118.265 152.060 118.355 ;
        RECT 150.100 117.455 150.325 117.585 ;
        RECT 150.495 117.515 151.020 117.735 ;
        RECT 151.190 118.095 152.060 118.265 ;
        RECT 149.735 116.865 149.985 117.325 ;
        RECT 150.155 117.315 150.325 117.455 ;
        RECT 151.190 117.315 151.360 118.095 ;
        RECT 151.890 118.025 152.060 118.095 ;
        RECT 151.570 117.845 151.770 117.875 ;
        RECT 152.230 117.845 152.400 118.915 ;
        RECT 152.570 118.025 152.760 118.745 ;
        RECT 151.570 117.545 152.400 117.845 ;
        RECT 152.930 117.815 153.250 118.775 ;
        RECT 150.155 117.145 150.490 117.315 ;
        RECT 150.685 117.145 151.360 117.315 ;
        RECT 151.680 116.865 152.050 117.365 ;
        RECT 152.230 117.315 152.400 117.545 ;
        RECT 152.785 117.485 153.250 117.815 ;
        RECT 153.420 118.105 153.590 118.945 ;
        RECT 153.770 118.915 154.085 119.415 ;
        RECT 154.315 118.685 154.655 119.245 ;
        RECT 153.760 118.310 154.655 118.685 ;
        RECT 154.825 118.405 154.995 119.415 ;
        RECT 154.465 118.105 154.655 118.310 ;
        RECT 155.165 118.355 155.495 119.200 ;
        RECT 155.165 118.275 155.555 118.355 ;
        RECT 155.340 118.225 155.555 118.275 ;
        RECT 153.420 117.775 154.295 118.105 ;
        RECT 154.465 117.775 155.215 118.105 ;
        RECT 153.420 117.315 153.590 117.775 ;
        RECT 154.465 117.605 154.665 117.775 ;
        RECT 155.385 117.645 155.555 118.225 ;
        RECT 155.725 118.325 156.935 119.415 ;
        RECT 155.725 117.785 156.245 118.325 ;
        RECT 155.330 117.605 155.555 117.645 ;
        RECT 156.415 117.615 156.935 118.155 ;
        RECT 152.230 117.145 152.635 117.315 ;
        RECT 152.805 117.145 153.590 117.315 ;
        RECT 153.865 116.865 154.075 117.395 ;
        RECT 154.335 117.080 154.665 117.605 ;
        RECT 155.175 117.520 155.555 117.605 ;
        RECT 154.835 116.865 155.005 117.475 ;
        RECT 155.175 117.085 155.505 117.520 ;
        RECT 155.725 116.865 156.935 117.615 ;
        RECT 22.700 116.695 157.020 116.865 ;
        RECT 22.785 115.945 23.995 116.695 ;
        RECT 24.255 116.145 24.425 116.435 ;
        RECT 24.595 116.315 24.925 116.695 ;
        RECT 24.255 115.975 24.920 116.145 ;
        RECT 22.785 115.405 23.305 115.945 ;
        RECT 23.475 115.235 23.995 115.775 ;
        RECT 22.785 114.145 23.995 115.235 ;
        RECT 24.170 115.155 24.520 115.805 ;
        RECT 24.690 114.985 24.920 115.975 ;
        RECT 24.255 114.815 24.920 114.985 ;
        RECT 24.255 114.315 24.425 114.815 ;
        RECT 24.595 114.145 24.925 114.645 ;
        RECT 25.095 114.315 25.280 116.435 ;
        RECT 25.535 116.235 25.785 116.695 ;
        RECT 25.955 116.245 26.290 116.415 ;
        RECT 26.485 116.245 27.160 116.415 ;
        RECT 25.955 116.105 26.125 116.245 ;
        RECT 25.450 115.115 25.730 116.065 ;
        RECT 25.900 115.975 26.125 116.105 ;
        RECT 25.900 114.870 26.070 115.975 ;
        RECT 26.295 115.825 26.820 116.045 ;
        RECT 26.240 115.060 26.480 115.655 ;
        RECT 26.650 115.125 26.820 115.825 ;
        RECT 26.990 115.465 27.160 116.245 ;
        RECT 27.480 116.195 27.850 116.695 ;
        RECT 28.030 116.245 28.435 116.415 ;
        RECT 28.605 116.245 29.390 116.415 ;
        RECT 28.030 116.015 28.200 116.245 ;
        RECT 27.370 115.715 28.200 116.015 ;
        RECT 28.585 115.745 29.050 116.075 ;
        RECT 27.370 115.685 27.570 115.715 ;
        RECT 27.690 115.465 27.860 115.535 ;
        RECT 26.990 115.295 27.860 115.465 ;
        RECT 27.350 115.205 27.860 115.295 ;
        RECT 25.900 114.740 26.205 114.870 ;
        RECT 26.650 114.760 27.180 115.125 ;
        RECT 25.520 114.145 25.785 114.605 ;
        RECT 25.955 114.315 26.205 114.740 ;
        RECT 27.350 114.590 27.520 115.205 ;
        RECT 26.415 114.420 27.520 114.590 ;
        RECT 27.690 114.145 27.860 114.945 ;
        RECT 28.030 114.645 28.200 115.715 ;
        RECT 28.370 114.815 28.560 115.535 ;
        RECT 28.730 114.785 29.050 115.745 ;
        RECT 29.220 115.785 29.390 116.245 ;
        RECT 29.665 116.165 29.875 116.695 ;
        RECT 30.135 115.955 30.465 116.480 ;
        RECT 30.635 116.085 30.805 116.695 ;
        RECT 30.975 116.040 31.305 116.475 ;
        RECT 31.615 116.145 31.785 116.435 ;
        RECT 31.955 116.315 32.285 116.695 ;
        RECT 30.975 115.955 31.355 116.040 ;
        RECT 31.615 115.975 32.280 116.145 ;
        RECT 30.265 115.785 30.465 115.955 ;
        RECT 31.130 115.915 31.355 115.955 ;
        RECT 29.220 115.455 30.095 115.785 ;
        RECT 30.265 115.455 31.015 115.785 ;
        RECT 28.030 114.315 28.280 114.645 ;
        RECT 29.220 114.615 29.390 115.455 ;
        RECT 30.265 115.250 30.455 115.455 ;
        RECT 31.185 115.335 31.355 115.915 ;
        RECT 31.140 115.285 31.355 115.335 ;
        RECT 29.560 114.875 30.455 115.250 ;
        RECT 30.965 115.205 31.355 115.285 ;
        RECT 28.505 114.445 29.390 114.615 ;
        RECT 29.570 114.145 29.885 114.645 ;
        RECT 30.115 114.315 30.455 114.875 ;
        RECT 30.625 114.145 30.795 115.155 ;
        RECT 30.965 114.360 31.295 115.205 ;
        RECT 31.530 115.155 31.880 115.805 ;
        RECT 32.050 114.985 32.280 115.975 ;
        RECT 31.615 114.815 32.280 114.985 ;
        RECT 31.615 114.315 31.785 114.815 ;
        RECT 31.955 114.145 32.285 114.645 ;
        RECT 32.455 114.315 32.640 116.435 ;
        RECT 32.895 116.235 33.145 116.695 ;
        RECT 33.315 116.245 33.650 116.415 ;
        RECT 33.845 116.245 34.520 116.415 ;
        RECT 33.315 116.105 33.485 116.245 ;
        RECT 32.810 115.115 33.090 116.065 ;
        RECT 33.260 115.975 33.485 116.105 ;
        RECT 33.260 114.870 33.430 115.975 ;
        RECT 33.655 115.825 34.180 116.045 ;
        RECT 33.600 115.060 33.840 115.655 ;
        RECT 34.010 115.125 34.180 115.825 ;
        RECT 34.350 115.465 34.520 116.245 ;
        RECT 34.840 116.195 35.210 116.695 ;
        RECT 35.390 116.245 35.795 116.415 ;
        RECT 35.965 116.245 36.750 116.415 ;
        RECT 35.390 116.015 35.560 116.245 ;
        RECT 34.730 115.715 35.560 116.015 ;
        RECT 35.945 115.745 36.410 116.075 ;
        RECT 34.730 115.685 34.930 115.715 ;
        RECT 35.050 115.465 35.220 115.535 ;
        RECT 34.350 115.295 35.220 115.465 ;
        RECT 34.710 115.205 35.220 115.295 ;
        RECT 33.260 114.740 33.565 114.870 ;
        RECT 34.010 114.760 34.540 115.125 ;
        RECT 32.880 114.145 33.145 114.605 ;
        RECT 33.315 114.315 33.565 114.740 ;
        RECT 34.710 114.590 34.880 115.205 ;
        RECT 33.775 114.420 34.880 114.590 ;
        RECT 35.050 114.145 35.220 114.945 ;
        RECT 35.390 114.645 35.560 115.715 ;
        RECT 35.730 114.815 35.920 115.535 ;
        RECT 36.090 114.785 36.410 115.745 ;
        RECT 36.580 115.785 36.750 116.245 ;
        RECT 37.025 116.165 37.235 116.695 ;
        RECT 37.495 115.955 37.825 116.480 ;
        RECT 37.995 116.085 38.165 116.695 ;
        RECT 38.335 116.040 38.665 116.475 ;
        RECT 38.335 115.955 38.715 116.040 ;
        RECT 37.625 115.785 37.825 115.955 ;
        RECT 38.490 115.915 38.715 115.955 ;
        RECT 36.580 115.455 37.455 115.785 ;
        RECT 37.625 115.455 38.375 115.785 ;
        RECT 35.390 114.315 35.640 114.645 ;
        RECT 36.580 114.615 36.750 115.455 ;
        RECT 37.625 115.250 37.815 115.455 ;
        RECT 38.545 115.335 38.715 115.915 ;
        RECT 38.885 115.945 40.095 116.695 ;
        RECT 40.265 115.955 40.625 116.330 ;
        RECT 40.890 115.955 41.060 116.695 ;
        RECT 41.340 116.125 41.510 116.330 ;
        RECT 41.340 115.955 41.880 116.125 ;
        RECT 38.885 115.405 39.405 115.945 ;
        RECT 38.500 115.285 38.715 115.335 ;
        RECT 36.920 114.875 37.815 115.250 ;
        RECT 38.325 115.205 38.715 115.285 ;
        RECT 39.575 115.235 40.095 115.775 ;
        RECT 35.865 114.445 36.750 114.615 ;
        RECT 36.930 114.145 37.245 114.645 ;
        RECT 37.475 114.315 37.815 114.875 ;
        RECT 37.985 114.145 38.155 115.155 ;
        RECT 38.325 114.360 38.655 115.205 ;
        RECT 38.885 114.145 40.095 115.235 ;
        RECT 40.265 115.300 40.520 115.955 ;
        RECT 40.690 115.455 41.040 115.785 ;
        RECT 41.210 115.455 41.540 115.785 ;
        RECT 40.265 114.315 40.605 115.300 ;
        RECT 40.775 114.915 41.040 115.455 ;
        RECT 41.710 115.255 41.880 115.955 ;
        RECT 41.255 115.085 41.880 115.255 ;
        RECT 42.050 115.325 42.220 116.525 ;
        RECT 42.450 116.045 42.780 116.525 ;
        RECT 42.950 116.225 43.120 116.695 ;
        RECT 43.290 116.045 43.620 116.510 ;
        RECT 42.450 115.875 43.620 116.045 ;
        RECT 44.405 115.955 44.790 116.525 ;
        RECT 44.960 116.235 45.285 116.695 ;
        RECT 45.805 116.065 46.085 116.525 ;
        RECT 42.390 115.495 42.960 115.705 ;
        RECT 43.130 115.495 43.775 115.705 ;
        RECT 42.050 114.915 42.755 115.325 ;
        RECT 44.405 115.285 44.685 115.955 ;
        RECT 44.960 115.895 46.085 116.065 ;
        RECT 44.960 115.785 45.410 115.895 ;
        RECT 44.855 115.455 45.410 115.785 ;
        RECT 46.275 115.725 46.675 116.525 ;
        RECT 47.075 116.235 47.345 116.695 ;
        RECT 47.515 116.065 47.800 116.525 ;
        RECT 40.775 114.745 42.755 114.915 ;
        RECT 40.775 114.145 41.185 114.575 ;
        RECT 41.930 114.145 42.260 114.565 ;
        RECT 42.430 114.315 42.755 114.745 ;
        RECT 43.230 114.145 43.560 115.245 ;
        RECT 44.405 114.315 44.790 115.285 ;
        RECT 44.960 114.995 45.410 115.455 ;
        RECT 45.580 115.165 46.675 115.725 ;
        RECT 44.960 114.775 46.085 114.995 ;
        RECT 44.960 114.145 45.285 114.605 ;
        RECT 45.805 114.315 46.085 114.775 ;
        RECT 46.275 114.315 46.675 115.165 ;
        RECT 46.845 115.895 47.800 116.065 ;
        RECT 48.545 115.970 48.835 116.695 ;
        RECT 49.095 116.145 49.265 116.435 ;
        RECT 49.435 116.315 49.765 116.695 ;
        RECT 49.095 115.975 49.760 116.145 ;
        RECT 46.845 114.995 47.055 115.895 ;
        RECT 47.225 115.165 47.915 115.725 ;
        RECT 46.845 114.775 47.800 114.995 ;
        RECT 47.075 114.145 47.345 114.605 ;
        RECT 47.515 114.315 47.800 114.775 ;
        RECT 48.545 114.145 48.835 115.310 ;
        RECT 49.010 115.155 49.360 115.805 ;
        RECT 49.530 114.985 49.760 115.975 ;
        RECT 49.095 114.815 49.760 114.985 ;
        RECT 49.095 114.315 49.265 114.815 ;
        RECT 49.435 114.145 49.765 114.645 ;
        RECT 49.935 114.315 50.120 116.435 ;
        RECT 50.375 116.235 50.625 116.695 ;
        RECT 50.795 116.245 51.130 116.415 ;
        RECT 51.325 116.245 52.000 116.415 ;
        RECT 50.795 116.105 50.965 116.245 ;
        RECT 50.290 115.115 50.570 116.065 ;
        RECT 50.740 115.975 50.965 116.105 ;
        RECT 50.740 114.870 50.910 115.975 ;
        RECT 51.135 115.825 51.660 116.045 ;
        RECT 51.080 115.060 51.320 115.655 ;
        RECT 51.490 115.125 51.660 115.825 ;
        RECT 51.830 115.465 52.000 116.245 ;
        RECT 52.320 116.195 52.690 116.695 ;
        RECT 52.870 116.245 53.275 116.415 ;
        RECT 53.445 116.245 54.230 116.415 ;
        RECT 52.870 116.015 53.040 116.245 ;
        RECT 52.210 115.715 53.040 116.015 ;
        RECT 53.425 115.745 53.890 116.075 ;
        RECT 52.210 115.685 52.410 115.715 ;
        RECT 52.530 115.465 52.700 115.535 ;
        RECT 51.830 115.295 52.700 115.465 ;
        RECT 52.190 115.205 52.700 115.295 ;
        RECT 50.740 114.740 51.045 114.870 ;
        RECT 51.490 114.760 52.020 115.125 ;
        RECT 50.360 114.145 50.625 114.605 ;
        RECT 50.795 114.315 51.045 114.740 ;
        RECT 52.190 114.590 52.360 115.205 ;
        RECT 51.255 114.420 52.360 114.590 ;
        RECT 52.530 114.145 52.700 114.945 ;
        RECT 52.870 114.645 53.040 115.715 ;
        RECT 53.210 114.815 53.400 115.535 ;
        RECT 53.570 114.785 53.890 115.745 ;
        RECT 54.060 115.785 54.230 116.245 ;
        RECT 54.505 116.165 54.715 116.695 ;
        RECT 54.975 115.955 55.305 116.480 ;
        RECT 55.475 116.085 55.645 116.695 ;
        RECT 55.815 116.040 56.145 116.475 ;
        RECT 55.815 115.955 56.195 116.040 ;
        RECT 55.105 115.785 55.305 115.955 ;
        RECT 55.970 115.915 56.195 115.955 ;
        RECT 54.060 115.455 54.935 115.785 ;
        RECT 55.105 115.455 55.855 115.785 ;
        RECT 52.870 114.315 53.120 114.645 ;
        RECT 54.060 114.615 54.230 115.455 ;
        RECT 55.105 115.250 55.295 115.455 ;
        RECT 56.025 115.335 56.195 115.915 ;
        RECT 55.980 115.285 56.195 115.335 ;
        RECT 54.400 114.875 55.295 115.250 ;
        RECT 55.805 115.205 56.195 115.285 ;
        RECT 56.365 115.955 56.750 116.525 ;
        RECT 56.920 116.235 57.245 116.695 ;
        RECT 57.765 116.065 58.045 116.525 ;
        RECT 56.365 115.285 56.645 115.955 ;
        RECT 56.920 115.895 58.045 116.065 ;
        RECT 56.920 115.785 57.370 115.895 ;
        RECT 56.815 115.455 57.370 115.785 ;
        RECT 58.235 115.725 58.635 116.525 ;
        RECT 59.035 116.235 59.305 116.695 ;
        RECT 59.475 116.065 59.760 116.525 ;
        RECT 60.215 116.180 60.385 116.695 ;
        RECT 53.345 114.445 54.230 114.615 ;
        RECT 54.410 114.145 54.725 114.645 ;
        RECT 54.955 114.315 55.295 114.875 ;
        RECT 55.465 114.145 55.635 115.155 ;
        RECT 55.805 114.360 56.135 115.205 ;
        RECT 56.365 114.315 56.750 115.285 ;
        RECT 56.920 114.995 57.370 115.455 ;
        RECT 57.540 115.165 58.635 115.725 ;
        RECT 56.920 114.775 58.045 114.995 ;
        RECT 56.920 114.145 57.245 114.605 ;
        RECT 57.765 114.315 58.045 114.775 ;
        RECT 58.235 114.315 58.635 115.165 ;
        RECT 58.805 115.895 59.760 116.065 ;
        RECT 60.555 116.040 60.885 116.475 ;
        RECT 61.055 116.085 61.225 116.695 ;
        RECT 60.505 115.955 60.885 116.040 ;
        RECT 61.395 115.955 61.725 116.480 ;
        RECT 61.985 116.165 62.195 116.695 ;
        RECT 62.470 116.245 63.255 116.415 ;
        RECT 63.425 116.245 63.830 116.415 ;
        RECT 60.505 115.915 60.730 115.955 ;
        RECT 58.805 114.995 59.015 115.895 ;
        RECT 59.185 115.165 59.875 115.725 ;
        RECT 60.505 115.335 60.675 115.915 ;
        RECT 61.395 115.785 61.595 115.955 ;
        RECT 62.470 115.785 62.640 116.245 ;
        RECT 60.845 115.455 61.595 115.785 ;
        RECT 61.765 115.455 62.640 115.785 ;
        RECT 60.505 115.285 60.720 115.335 ;
        RECT 60.505 115.205 60.895 115.285 ;
        RECT 58.805 114.775 59.760 114.995 ;
        RECT 59.035 114.145 59.305 114.605 ;
        RECT 59.475 114.315 59.760 114.775 ;
        RECT 60.225 114.145 60.395 115.060 ;
        RECT 60.565 114.360 60.895 115.205 ;
        RECT 61.405 115.250 61.595 115.455 ;
        RECT 61.065 114.145 61.235 115.155 ;
        RECT 61.405 114.875 62.300 115.250 ;
        RECT 61.405 114.315 61.745 114.875 ;
        RECT 61.975 114.145 62.290 114.645 ;
        RECT 62.470 114.615 62.640 115.455 ;
        RECT 62.810 115.745 63.275 116.075 ;
        RECT 63.660 116.015 63.830 116.245 ;
        RECT 64.010 116.195 64.380 116.695 ;
        RECT 64.700 116.245 65.375 116.415 ;
        RECT 65.570 116.245 65.905 116.415 ;
        RECT 62.810 114.785 63.130 115.745 ;
        RECT 63.660 115.715 64.490 116.015 ;
        RECT 63.300 114.815 63.490 115.535 ;
        RECT 63.660 114.645 63.830 115.715 ;
        RECT 64.290 115.685 64.490 115.715 ;
        RECT 64.000 115.465 64.170 115.535 ;
        RECT 64.700 115.465 64.870 116.245 ;
        RECT 65.735 116.105 65.905 116.245 ;
        RECT 66.075 116.235 66.325 116.695 ;
        RECT 64.000 115.295 64.870 115.465 ;
        RECT 65.040 115.825 65.565 116.045 ;
        RECT 65.735 115.975 65.960 116.105 ;
        RECT 64.000 115.205 64.510 115.295 ;
        RECT 62.470 114.445 63.355 114.615 ;
        RECT 63.580 114.315 63.830 114.645 ;
        RECT 64.000 114.145 64.170 114.945 ;
        RECT 64.340 114.590 64.510 115.205 ;
        RECT 65.040 115.125 65.210 115.825 ;
        RECT 64.680 114.760 65.210 115.125 ;
        RECT 65.380 115.060 65.620 115.655 ;
        RECT 65.790 114.870 65.960 115.975 ;
        RECT 66.130 115.115 66.410 116.065 ;
        RECT 65.655 114.740 65.960 114.870 ;
        RECT 64.340 114.420 65.445 114.590 ;
        RECT 65.655 114.315 65.905 114.740 ;
        RECT 66.075 114.145 66.340 114.605 ;
        RECT 66.580 114.315 66.765 116.435 ;
        RECT 66.935 116.315 67.265 116.695 ;
        RECT 67.435 116.145 67.605 116.435 ;
        RECT 67.865 116.315 68.755 116.485 ;
        RECT 66.940 115.975 67.605 116.145 ;
        RECT 66.940 114.985 67.170 115.975 ;
        RECT 67.340 115.155 67.690 115.805 ;
        RECT 67.865 115.760 68.415 116.145 ;
        RECT 68.585 115.590 68.755 116.315 ;
        RECT 67.865 115.520 68.755 115.590 ;
        RECT 68.925 115.990 69.145 116.475 ;
        RECT 69.315 116.155 69.565 116.695 ;
        RECT 69.735 116.045 69.995 116.525 ;
        RECT 68.925 115.565 69.255 115.990 ;
        RECT 67.865 115.495 68.760 115.520 ;
        RECT 67.865 115.480 68.770 115.495 ;
        RECT 67.865 115.465 68.775 115.480 ;
        RECT 67.865 115.460 68.785 115.465 ;
        RECT 67.865 115.450 68.790 115.460 ;
        RECT 67.865 115.440 68.795 115.450 ;
        RECT 67.865 115.435 68.805 115.440 ;
        RECT 67.865 115.425 68.815 115.435 ;
        RECT 67.865 115.420 68.825 115.425 ;
        RECT 66.940 114.815 67.605 114.985 ;
        RECT 67.865 114.970 68.125 115.420 ;
        RECT 68.490 115.415 68.825 115.420 ;
        RECT 68.490 115.410 68.840 115.415 ;
        RECT 68.490 115.400 68.855 115.410 ;
        RECT 68.490 115.395 68.880 115.400 ;
        RECT 69.425 115.395 69.655 115.790 ;
        RECT 68.490 115.390 69.655 115.395 ;
        RECT 68.520 115.355 69.655 115.390 ;
        RECT 68.555 115.330 69.655 115.355 ;
        RECT 68.585 115.300 69.655 115.330 ;
        RECT 68.605 115.270 69.655 115.300 ;
        RECT 68.625 115.240 69.655 115.270 ;
        RECT 68.695 115.230 69.655 115.240 ;
        RECT 68.720 115.220 69.655 115.230 ;
        RECT 68.740 115.205 69.655 115.220 ;
        RECT 68.760 115.190 69.655 115.205 ;
        RECT 68.765 115.180 69.550 115.190 ;
        RECT 68.780 115.145 69.550 115.180 ;
        RECT 66.935 114.145 67.265 114.645 ;
        RECT 67.435 114.315 67.605 114.815 ;
        RECT 68.295 114.825 68.625 115.070 ;
        RECT 68.795 114.895 69.550 115.145 ;
        RECT 69.825 115.015 69.995 116.045 ;
        RECT 68.295 114.800 68.480 114.825 ;
        RECT 67.865 114.700 68.480 114.800 ;
        RECT 67.865 114.145 68.470 114.700 ;
        RECT 68.645 114.315 69.125 114.655 ;
        RECT 69.295 114.145 69.550 114.690 ;
        RECT 69.720 114.315 69.995 115.015 ;
        RECT 70.165 115.955 70.550 116.525 ;
        RECT 70.720 116.235 71.045 116.695 ;
        RECT 71.565 116.065 71.845 116.525 ;
        RECT 70.165 115.285 70.445 115.955 ;
        RECT 70.720 115.895 71.845 116.065 ;
        RECT 70.720 115.785 71.170 115.895 ;
        RECT 70.615 115.455 71.170 115.785 ;
        RECT 72.035 115.725 72.435 116.525 ;
        RECT 72.835 116.235 73.105 116.695 ;
        RECT 73.275 116.065 73.560 116.525 ;
        RECT 70.165 114.315 70.550 115.285 ;
        RECT 70.720 114.995 71.170 115.455 ;
        RECT 71.340 115.165 72.435 115.725 ;
        RECT 70.720 114.775 71.845 114.995 ;
        RECT 70.720 114.145 71.045 114.605 ;
        RECT 71.565 114.315 71.845 114.775 ;
        RECT 72.035 114.315 72.435 115.165 ;
        RECT 72.605 115.895 73.560 116.065 ;
        RECT 74.305 115.970 74.595 116.695 ;
        RECT 72.605 114.995 72.815 115.895 ;
        RECT 72.985 115.165 73.675 115.725 ;
        RECT 72.605 114.775 73.560 114.995 ;
        RECT 72.835 114.145 73.105 114.605 ;
        RECT 73.275 114.315 73.560 114.775 ;
        RECT 74.305 114.145 74.595 115.310 ;
        RECT 74.775 114.325 75.035 116.515 ;
        RECT 75.295 116.325 75.965 116.695 ;
        RECT 76.145 116.145 76.455 116.515 ;
        RECT 75.225 115.945 76.455 116.145 ;
        RECT 75.225 115.275 75.515 115.945 ;
        RECT 76.635 115.765 76.865 116.405 ;
        RECT 77.045 115.965 77.335 116.695 ;
        RECT 75.695 115.455 76.160 115.765 ;
        RECT 76.340 115.455 76.865 115.765 ;
        RECT 77.045 115.455 77.345 115.785 ;
        RECT 75.225 115.055 75.995 115.275 ;
        RECT 75.205 114.145 75.545 114.875 ;
        RECT 75.725 114.325 75.995 115.055 ;
        RECT 76.175 115.035 77.335 115.275 ;
        RECT 76.175 114.325 76.405 115.035 ;
        RECT 76.575 114.145 76.905 114.855 ;
        RECT 77.075 114.325 77.335 115.035 ;
        RECT 77.535 114.325 77.795 116.515 ;
        RECT 78.055 116.325 78.725 116.695 ;
        RECT 78.905 116.145 79.215 116.515 ;
        RECT 77.985 115.945 79.215 116.145 ;
        RECT 77.985 115.275 78.275 115.945 ;
        RECT 79.395 115.765 79.625 116.405 ;
        RECT 79.805 115.965 80.095 116.695 ;
        RECT 80.375 116.145 80.545 116.435 ;
        RECT 80.715 116.315 81.045 116.695 ;
        RECT 80.375 115.975 81.040 116.145 ;
        RECT 78.455 115.455 78.920 115.765 ;
        RECT 79.100 115.455 79.625 115.765 ;
        RECT 79.805 115.455 80.105 115.785 ;
        RECT 77.985 115.055 78.755 115.275 ;
        RECT 77.965 114.145 78.305 114.875 ;
        RECT 78.485 114.325 78.755 115.055 ;
        RECT 78.935 115.035 80.095 115.275 ;
        RECT 80.290 115.155 80.640 115.805 ;
        RECT 78.935 114.325 79.165 115.035 ;
        RECT 79.335 114.145 79.665 114.855 ;
        RECT 79.835 114.325 80.095 115.035 ;
        RECT 80.810 114.985 81.040 115.975 ;
        RECT 80.375 114.815 81.040 114.985 ;
        RECT 80.375 114.315 80.545 114.815 ;
        RECT 80.715 114.145 81.045 114.645 ;
        RECT 81.215 114.315 81.400 116.435 ;
        RECT 81.655 116.235 81.905 116.695 ;
        RECT 82.075 116.245 82.410 116.415 ;
        RECT 82.605 116.245 83.280 116.415 ;
        RECT 82.075 116.105 82.245 116.245 ;
        RECT 81.570 115.115 81.850 116.065 ;
        RECT 82.020 115.975 82.245 116.105 ;
        RECT 82.020 114.870 82.190 115.975 ;
        RECT 82.415 115.825 82.940 116.045 ;
        RECT 82.360 115.060 82.600 115.655 ;
        RECT 82.770 115.125 82.940 115.825 ;
        RECT 83.110 115.465 83.280 116.245 ;
        RECT 83.600 116.195 83.970 116.695 ;
        RECT 84.150 116.245 84.555 116.415 ;
        RECT 84.725 116.245 85.510 116.415 ;
        RECT 84.150 116.015 84.320 116.245 ;
        RECT 83.490 115.715 84.320 116.015 ;
        RECT 84.705 115.745 85.170 116.075 ;
        RECT 83.490 115.685 83.690 115.715 ;
        RECT 83.810 115.465 83.980 115.535 ;
        RECT 83.110 115.295 83.980 115.465 ;
        RECT 83.470 115.205 83.980 115.295 ;
        RECT 82.020 114.740 82.325 114.870 ;
        RECT 82.770 114.760 83.300 115.125 ;
        RECT 81.640 114.145 81.905 114.605 ;
        RECT 82.075 114.315 82.325 114.740 ;
        RECT 83.470 114.590 83.640 115.205 ;
        RECT 82.535 114.420 83.640 114.590 ;
        RECT 83.810 114.145 83.980 114.945 ;
        RECT 84.150 114.645 84.320 115.715 ;
        RECT 84.490 114.815 84.680 115.535 ;
        RECT 84.850 114.785 85.170 115.745 ;
        RECT 85.340 115.785 85.510 116.245 ;
        RECT 85.785 116.165 85.995 116.695 ;
        RECT 86.255 115.955 86.585 116.480 ;
        RECT 86.755 116.085 86.925 116.695 ;
        RECT 87.095 116.040 87.425 116.475 ;
        RECT 87.595 116.180 87.765 116.695 ;
        RECT 87.095 115.955 87.475 116.040 ;
        RECT 86.385 115.785 86.585 115.955 ;
        RECT 87.250 115.915 87.475 115.955 ;
        RECT 85.340 115.455 86.215 115.785 ;
        RECT 86.385 115.455 87.135 115.785 ;
        RECT 84.150 114.315 84.400 114.645 ;
        RECT 85.340 114.615 85.510 115.455 ;
        RECT 86.385 115.250 86.575 115.455 ;
        RECT 87.305 115.335 87.475 115.915 ;
        RECT 87.260 115.285 87.475 115.335 ;
        RECT 85.680 114.875 86.575 115.250 ;
        RECT 87.085 115.205 87.475 115.285 ;
        RECT 84.625 114.445 85.510 114.615 ;
        RECT 85.690 114.145 86.005 114.645 ;
        RECT 86.235 114.315 86.575 114.875 ;
        RECT 86.745 114.145 86.915 115.155 ;
        RECT 87.085 114.360 87.415 115.205 ;
        RECT 87.585 114.145 87.755 115.060 ;
        RECT 89.035 114.325 89.295 116.515 ;
        RECT 89.555 116.325 90.225 116.695 ;
        RECT 90.405 116.145 90.715 116.515 ;
        RECT 89.485 115.945 90.715 116.145 ;
        RECT 89.485 115.275 89.775 115.945 ;
        RECT 90.895 115.765 91.125 116.405 ;
        RECT 91.305 115.965 91.595 116.695 ;
        RECT 91.785 115.945 92.995 116.695 ;
        RECT 93.170 116.295 93.505 116.695 ;
        RECT 93.675 116.125 93.880 116.525 ;
        RECT 94.090 116.215 94.365 116.695 ;
        RECT 94.575 116.195 94.835 116.525 ;
        RECT 93.195 115.955 93.880 116.125 ;
        RECT 89.955 115.455 90.420 115.765 ;
        RECT 90.600 115.455 91.125 115.765 ;
        RECT 91.305 115.455 91.605 115.785 ;
        RECT 91.785 115.405 92.305 115.945 ;
        RECT 89.485 115.055 90.255 115.275 ;
        RECT 89.465 114.145 89.805 114.875 ;
        RECT 89.985 114.325 90.255 115.055 ;
        RECT 90.435 115.035 91.595 115.275 ;
        RECT 92.475 115.235 92.995 115.775 ;
        RECT 90.435 114.325 90.665 115.035 ;
        RECT 90.835 114.145 91.165 114.855 ;
        RECT 91.335 114.325 91.595 115.035 ;
        RECT 91.785 114.145 92.995 115.235 ;
        RECT 93.195 114.925 93.535 115.955 ;
        RECT 93.705 115.285 93.955 115.785 ;
        RECT 94.135 115.455 94.495 116.035 ;
        RECT 94.665 115.285 94.835 116.195 ;
        RECT 95.005 115.925 97.595 116.695 ;
        RECT 98.315 116.355 98.485 116.390 ;
        RECT 98.285 116.185 98.485 116.355 ;
        RECT 95.005 115.405 96.215 115.925 ;
        RECT 98.315 115.825 98.485 116.185 ;
        RECT 98.675 116.165 98.905 116.470 ;
        RECT 99.075 116.335 99.405 116.695 ;
        RECT 99.600 116.165 99.890 116.515 ;
        RECT 98.675 115.995 99.890 116.165 ;
        RECT 100.065 115.970 100.355 116.695 ;
        RECT 100.525 116.150 105.870 116.695 ;
        RECT 93.705 115.115 94.835 115.285 ;
        RECT 96.385 115.235 97.595 115.755 ;
        RECT 98.315 115.655 98.835 115.825 ;
        RECT 93.195 114.750 93.860 114.925 ;
        RECT 93.170 114.145 93.505 114.570 ;
        RECT 93.675 114.345 93.860 114.750 ;
        RECT 94.065 114.145 94.395 114.925 ;
        RECT 94.565 114.345 94.835 115.115 ;
        RECT 95.005 114.145 97.595 115.235 ;
        RECT 98.230 115.125 98.475 115.485 ;
        RECT 98.665 115.275 98.835 115.655 ;
        RECT 99.005 115.455 99.390 115.785 ;
        RECT 99.570 115.675 99.830 115.785 ;
        RECT 99.570 115.505 99.835 115.675 ;
        RECT 99.570 115.455 99.830 115.505 ;
        RECT 98.665 114.995 99.015 115.275 ;
        RECT 98.230 114.145 98.485 114.945 ;
        RECT 98.685 114.315 99.015 114.995 ;
        RECT 99.195 114.405 99.390 115.455 ;
        RECT 102.110 115.320 102.450 116.150 ;
        RECT 106.045 115.925 109.555 116.695 ;
        RECT 110.300 116.065 110.585 116.525 ;
        RECT 110.755 116.235 111.025 116.695 ;
        RECT 99.570 114.145 99.890 115.285 ;
        RECT 100.065 114.145 100.355 115.310 ;
        RECT 103.930 114.580 104.280 115.830 ;
        RECT 106.045 115.405 107.695 115.925 ;
        RECT 110.300 115.895 111.255 116.065 ;
        RECT 107.865 115.235 109.555 115.755 ;
        RECT 100.525 114.145 105.870 114.580 ;
        RECT 106.045 114.145 109.555 115.235 ;
        RECT 110.185 115.165 110.875 115.725 ;
        RECT 111.045 114.995 111.255 115.895 ;
        RECT 110.300 114.775 111.255 114.995 ;
        RECT 111.425 115.725 111.825 116.525 ;
        RECT 112.015 116.065 112.295 116.525 ;
        RECT 112.815 116.235 113.140 116.695 ;
        RECT 112.015 115.895 113.140 116.065 ;
        RECT 113.310 115.955 113.695 116.525 ;
        RECT 113.885 115.965 114.175 116.695 ;
        RECT 112.690 115.785 113.140 115.895 ;
        RECT 111.425 115.165 112.520 115.725 ;
        RECT 112.690 115.455 113.245 115.785 ;
        RECT 110.300 114.315 110.585 114.775 ;
        RECT 110.755 114.145 111.025 114.605 ;
        RECT 111.425 114.315 111.825 115.165 ;
        RECT 112.690 114.995 113.140 115.455 ;
        RECT 113.415 115.285 113.695 115.955 ;
        RECT 113.875 115.455 114.175 115.785 ;
        RECT 114.355 115.765 114.585 116.405 ;
        RECT 114.765 116.145 115.075 116.515 ;
        RECT 115.255 116.325 115.925 116.695 ;
        RECT 114.765 115.945 115.995 116.145 ;
        RECT 114.355 115.455 114.880 115.765 ;
        RECT 115.060 115.455 115.525 115.765 ;
        RECT 112.015 114.775 113.140 114.995 ;
        RECT 112.015 114.315 112.295 114.775 ;
        RECT 112.815 114.145 113.140 114.605 ;
        RECT 113.310 114.315 113.695 115.285 ;
        RECT 115.705 115.275 115.995 115.945 ;
        RECT 113.885 115.035 115.045 115.275 ;
        RECT 113.885 114.325 114.145 115.035 ;
        RECT 114.315 114.145 114.645 114.855 ;
        RECT 114.815 114.325 115.045 115.035 ;
        RECT 115.225 115.055 115.995 115.275 ;
        RECT 115.225 114.325 115.495 115.055 ;
        RECT 115.675 114.145 116.015 114.875 ;
        RECT 116.185 114.325 116.445 116.515 ;
        RECT 116.625 115.925 118.295 116.695 ;
        RECT 118.465 115.955 118.850 116.525 ;
        RECT 119.020 116.235 119.345 116.695 ;
        RECT 119.865 116.065 120.145 116.525 ;
        RECT 116.625 115.405 117.375 115.925 ;
        RECT 117.545 115.235 118.295 115.755 ;
        RECT 116.625 114.145 118.295 115.235 ;
        RECT 118.465 115.285 118.745 115.955 ;
        RECT 119.020 115.895 120.145 116.065 ;
        RECT 119.020 115.785 119.470 115.895 ;
        RECT 118.915 115.455 119.470 115.785 ;
        RECT 120.335 115.725 120.735 116.525 ;
        RECT 121.135 116.235 121.405 116.695 ;
        RECT 121.575 116.065 121.860 116.525 ;
        RECT 118.465 114.315 118.850 115.285 ;
        RECT 119.020 114.995 119.470 115.455 ;
        RECT 119.640 115.165 120.735 115.725 ;
        RECT 119.020 114.775 120.145 114.995 ;
        RECT 119.020 114.145 119.345 114.605 ;
        RECT 119.865 114.315 120.145 114.775 ;
        RECT 120.335 114.315 120.735 115.165 ;
        RECT 120.905 115.895 121.860 116.065 ;
        RECT 122.145 115.925 125.655 116.695 ;
        RECT 125.825 115.970 126.115 116.695 ;
        RECT 127.210 116.020 127.485 116.365 ;
        RECT 127.675 116.295 128.055 116.695 ;
        RECT 128.225 116.125 128.395 116.475 ;
        RECT 128.565 116.295 128.895 116.695 ;
        RECT 129.065 116.125 129.320 116.475 ;
        RECT 120.905 114.995 121.115 115.895 ;
        RECT 121.285 115.165 121.975 115.725 ;
        RECT 122.145 115.405 123.795 115.925 ;
        RECT 123.965 115.235 125.655 115.755 ;
        RECT 120.905 114.775 121.860 114.995 ;
        RECT 121.135 114.145 121.405 114.605 ;
        RECT 121.575 114.315 121.860 114.775 ;
        RECT 122.145 114.145 125.655 115.235 ;
        RECT 125.825 114.145 126.115 115.310 ;
        RECT 127.210 115.285 127.380 116.020 ;
        RECT 127.655 115.955 129.320 116.125 ;
        RECT 127.655 115.785 127.825 115.955 ;
        RECT 129.505 115.875 129.765 116.695 ;
        RECT 129.935 115.875 130.265 116.295 ;
        RECT 130.445 116.125 130.705 116.525 ;
        RECT 130.875 116.295 131.205 116.695 ;
        RECT 131.375 116.125 131.545 116.475 ;
        RECT 131.715 116.295 132.090 116.695 ;
        RECT 130.445 115.955 132.110 116.125 ;
        RECT 132.280 116.020 132.555 116.365 ;
        RECT 130.015 115.785 130.265 115.875 ;
        RECT 131.940 115.785 132.110 115.955 ;
        RECT 127.550 115.455 127.825 115.785 ;
        RECT 127.995 115.455 128.820 115.785 ;
        RECT 128.990 115.455 129.335 115.785 ;
        RECT 129.510 115.455 129.845 115.705 ;
        RECT 130.015 115.455 130.730 115.785 ;
        RECT 130.945 115.455 131.770 115.785 ;
        RECT 131.940 115.455 132.215 115.785 ;
        RECT 127.655 115.285 127.825 115.455 ;
        RECT 127.210 114.315 127.485 115.285 ;
        RECT 127.655 115.115 128.315 115.285 ;
        RECT 128.625 115.165 128.820 115.455 ;
        RECT 128.145 114.995 128.315 115.115 ;
        RECT 128.990 114.995 129.315 115.285 ;
        RECT 127.695 114.145 127.975 114.945 ;
        RECT 128.145 114.825 129.315 114.995 ;
        RECT 128.145 114.365 129.335 114.655 ;
        RECT 129.505 114.145 129.765 115.285 ;
        RECT 130.015 114.895 130.185 115.455 ;
        RECT 130.445 114.995 130.775 115.285 ;
        RECT 130.945 115.165 131.190 115.455 ;
        RECT 131.940 115.285 132.110 115.455 ;
        RECT 132.385 115.285 132.555 116.020 ;
        RECT 131.450 115.115 132.110 115.285 ;
        RECT 131.450 114.995 131.620 115.115 ;
        RECT 130.445 114.825 131.620 114.995 ;
        RECT 130.005 114.325 131.620 114.655 ;
        RECT 131.790 114.145 132.070 114.945 ;
        RECT 132.280 114.315 132.555 115.285 ;
        RECT 132.760 115.955 133.375 116.525 ;
        RECT 133.545 116.185 133.760 116.695 ;
        RECT 133.990 116.185 134.270 116.515 ;
        RECT 134.450 116.185 134.690 116.695 ;
        RECT 135.190 116.185 135.430 116.695 ;
        RECT 135.610 116.185 135.890 116.515 ;
        RECT 136.120 116.185 136.335 116.695 ;
        RECT 132.760 114.935 133.075 115.955 ;
        RECT 133.245 115.285 133.415 115.785 ;
        RECT 133.665 115.455 133.930 116.015 ;
        RECT 134.100 115.285 134.270 116.185 ;
        RECT 134.440 115.455 134.795 116.015 ;
        RECT 135.085 115.455 135.440 116.015 ;
        RECT 135.610 115.285 135.780 116.185 ;
        RECT 135.950 115.455 136.215 116.015 ;
        RECT 136.505 115.955 137.120 116.525 ;
        RECT 136.465 115.285 136.635 115.785 ;
        RECT 133.245 115.115 134.670 115.285 ;
        RECT 132.760 114.315 133.295 114.935 ;
        RECT 133.465 114.145 133.795 114.945 ;
        RECT 134.280 114.940 134.670 115.115 ;
        RECT 135.210 115.115 136.635 115.285 ;
        RECT 135.210 114.940 135.600 115.115 ;
        RECT 136.085 114.145 136.415 114.945 ;
        RECT 136.805 114.935 137.120 115.955 ;
        RECT 136.585 114.315 137.120 114.935 ;
        RECT 137.325 116.195 137.585 116.525 ;
        RECT 137.795 116.215 138.070 116.695 ;
        RECT 137.325 115.285 137.495 116.195 ;
        RECT 138.280 116.125 138.485 116.525 ;
        RECT 138.655 116.295 138.990 116.695 ;
        RECT 137.665 115.455 138.025 116.035 ;
        RECT 138.280 115.955 138.965 116.125 ;
        RECT 138.205 115.285 138.455 115.785 ;
        RECT 137.325 115.115 138.455 115.285 ;
        RECT 137.325 114.345 137.595 115.115 ;
        RECT 138.625 114.925 138.965 115.955 ;
        RECT 137.765 114.145 138.095 114.925 ;
        RECT 138.300 114.750 138.965 114.925 ;
        RECT 139.200 115.955 139.815 116.525 ;
        RECT 139.985 116.185 140.200 116.695 ;
        RECT 140.430 116.185 140.710 116.515 ;
        RECT 140.890 116.185 141.130 116.695 ;
        RECT 139.200 114.935 139.515 115.955 ;
        RECT 139.685 115.285 139.855 115.785 ;
        RECT 140.105 115.455 140.370 116.015 ;
        RECT 140.540 115.285 140.710 116.185 ;
        RECT 140.880 115.455 141.235 116.015 ;
        RECT 141.465 115.945 142.675 116.695 ;
        RECT 142.960 116.065 143.245 116.525 ;
        RECT 143.415 116.235 143.685 116.695 ;
        RECT 141.465 115.405 141.985 115.945 ;
        RECT 142.960 115.895 143.915 116.065 ;
        RECT 139.685 115.115 141.110 115.285 ;
        RECT 142.155 115.235 142.675 115.775 ;
        RECT 138.300 114.345 138.485 114.750 ;
        RECT 138.655 114.145 138.990 114.570 ;
        RECT 139.200 114.315 139.735 114.935 ;
        RECT 139.905 114.145 140.235 114.945 ;
        RECT 140.720 114.940 141.110 115.115 ;
        RECT 141.465 114.145 142.675 115.235 ;
        RECT 142.845 115.165 143.535 115.725 ;
        RECT 143.705 114.995 143.915 115.895 ;
        RECT 142.960 114.775 143.915 114.995 ;
        RECT 144.085 115.725 144.485 116.525 ;
        RECT 144.675 116.065 144.955 116.525 ;
        RECT 145.475 116.235 145.800 116.695 ;
        RECT 144.675 115.895 145.800 116.065 ;
        RECT 145.970 115.955 146.355 116.525 ;
        RECT 145.350 115.785 145.800 115.895 ;
        RECT 144.085 115.165 145.180 115.725 ;
        RECT 145.350 115.455 145.905 115.785 ;
        RECT 142.960 114.315 143.245 114.775 ;
        RECT 143.415 114.145 143.685 114.605 ;
        RECT 144.085 114.315 144.485 115.165 ;
        RECT 145.350 114.995 145.800 115.455 ;
        RECT 146.075 115.285 146.355 115.955 ;
        RECT 144.675 114.775 145.800 114.995 ;
        RECT 144.675 114.315 144.955 114.775 ;
        RECT 145.475 114.145 145.800 114.605 ;
        RECT 145.970 114.315 146.355 115.285 ;
        RECT 146.525 115.895 146.865 116.525 ;
        RECT 147.035 115.895 147.285 116.695 ;
        RECT 147.475 116.045 147.805 116.525 ;
        RECT 147.975 116.235 148.200 116.695 ;
        RECT 148.370 116.045 148.700 116.525 ;
        RECT 146.525 115.335 146.700 115.895 ;
        RECT 147.475 115.875 148.700 116.045 ;
        RECT 149.330 115.915 149.830 116.525 ;
        RECT 150.205 115.945 151.415 116.695 ;
        RECT 151.585 115.970 151.875 116.695 ;
        RECT 146.870 115.535 147.565 115.705 ;
        RECT 146.525 115.285 146.755 115.335 ;
        RECT 147.395 115.285 147.565 115.535 ;
        RECT 147.740 115.505 148.160 115.705 ;
        RECT 148.330 115.505 148.660 115.705 ;
        RECT 148.830 115.505 149.160 115.705 ;
        RECT 149.330 115.285 149.500 115.915 ;
        RECT 149.685 115.455 150.035 115.705 ;
        RECT 150.205 115.405 150.725 115.945 ;
        RECT 152.045 115.895 152.385 116.525 ;
        RECT 152.555 115.895 152.805 116.695 ;
        RECT 152.995 116.045 153.325 116.525 ;
        RECT 153.495 116.235 153.720 116.695 ;
        RECT 153.890 116.045 154.220 116.525 ;
        RECT 146.525 114.315 146.865 115.285 ;
        RECT 147.035 114.145 147.205 115.285 ;
        RECT 147.395 115.115 149.830 115.285 ;
        RECT 150.895 115.235 151.415 115.775 ;
        RECT 147.475 114.145 147.725 114.945 ;
        RECT 148.370 114.315 148.700 115.115 ;
        RECT 149.000 114.145 149.330 114.945 ;
        RECT 149.500 114.315 149.830 115.115 ;
        RECT 150.205 114.145 151.415 115.235 ;
        RECT 151.585 114.145 151.875 115.310 ;
        RECT 152.045 115.285 152.220 115.895 ;
        RECT 152.995 115.875 154.220 116.045 ;
        RECT 154.850 115.915 155.350 116.525 ;
        RECT 155.725 115.945 156.935 116.695 ;
        RECT 152.390 115.535 153.085 115.705 ;
        RECT 152.915 115.285 153.085 115.535 ;
        RECT 153.260 115.505 153.680 115.705 ;
        RECT 153.850 115.505 154.180 115.705 ;
        RECT 154.350 115.505 154.680 115.705 ;
        RECT 154.850 115.285 155.020 115.915 ;
        RECT 155.205 115.455 155.555 115.705 ;
        RECT 152.045 114.315 152.385 115.285 ;
        RECT 152.555 114.145 152.725 115.285 ;
        RECT 152.915 115.115 155.350 115.285 ;
        RECT 152.995 114.145 153.245 114.945 ;
        RECT 153.890 114.315 154.220 115.115 ;
        RECT 154.520 114.145 154.850 114.945 ;
        RECT 155.020 114.315 155.350 115.115 ;
        RECT 155.725 115.235 156.245 115.775 ;
        RECT 156.415 115.405 156.935 115.945 ;
        RECT 155.725 114.145 156.935 115.235 ;
        RECT 22.700 113.975 157.020 114.145 ;
        RECT 22.785 112.885 23.995 113.975 ;
        RECT 24.165 112.885 25.835 113.975 ;
        RECT 22.785 112.175 23.305 112.715 ;
        RECT 23.475 112.345 23.995 112.885 ;
        RECT 24.165 112.195 24.915 112.715 ;
        RECT 25.085 112.365 25.835 112.885 ;
        RECT 26.465 112.835 26.850 113.805 ;
        RECT 27.020 113.515 27.345 113.975 ;
        RECT 27.865 113.345 28.145 113.805 ;
        RECT 27.020 113.125 28.145 113.345 ;
        RECT 22.785 111.425 23.995 112.175 ;
        RECT 24.165 111.425 25.835 112.195 ;
        RECT 26.465 112.165 26.745 112.835 ;
        RECT 27.020 112.665 27.470 113.125 ;
        RECT 28.335 112.955 28.735 113.805 ;
        RECT 29.135 113.515 29.405 113.975 ;
        RECT 29.575 113.345 29.860 113.805 ;
        RECT 26.915 112.335 27.470 112.665 ;
        RECT 27.640 112.395 28.735 112.955 ;
        RECT 27.020 112.225 27.470 112.335 ;
        RECT 26.465 111.595 26.850 112.165 ;
        RECT 27.020 112.055 28.145 112.225 ;
        RECT 27.020 111.425 27.345 111.885 ;
        RECT 27.865 111.595 28.145 112.055 ;
        RECT 28.335 111.595 28.735 112.395 ;
        RECT 28.905 113.125 29.860 113.345 ;
        RECT 28.905 112.225 29.115 113.125 ;
        RECT 29.285 112.395 29.975 112.955 ;
        RECT 30.145 112.835 30.530 113.805 ;
        RECT 30.700 113.515 31.025 113.975 ;
        RECT 31.545 113.345 31.825 113.805 ;
        RECT 30.700 113.125 31.825 113.345 ;
        RECT 28.905 112.055 29.860 112.225 ;
        RECT 29.135 111.425 29.405 111.885 ;
        RECT 29.575 111.595 29.860 112.055 ;
        RECT 30.145 112.165 30.425 112.835 ;
        RECT 30.700 112.665 31.150 113.125 ;
        RECT 32.015 112.955 32.415 113.805 ;
        RECT 32.815 113.515 33.085 113.975 ;
        RECT 33.255 113.345 33.540 113.805 ;
        RECT 30.595 112.335 31.150 112.665 ;
        RECT 31.320 112.395 32.415 112.955 ;
        RECT 30.700 112.225 31.150 112.335 ;
        RECT 30.145 111.595 30.530 112.165 ;
        RECT 30.700 112.055 31.825 112.225 ;
        RECT 30.700 111.425 31.025 111.885 ;
        RECT 31.545 111.595 31.825 112.055 ;
        RECT 32.015 111.595 32.415 112.395 ;
        RECT 32.585 113.125 33.540 113.345 ;
        RECT 32.585 112.225 32.795 113.125 ;
        RECT 32.965 112.395 33.655 112.955 ;
        RECT 33.825 112.885 35.495 113.975 ;
        RECT 32.585 112.055 33.540 112.225 ;
        RECT 32.815 111.425 33.085 111.885 ;
        RECT 33.255 111.595 33.540 112.055 ;
        RECT 33.825 112.195 34.575 112.715 ;
        RECT 34.745 112.365 35.495 112.885 ;
        RECT 35.665 112.810 35.955 113.975 ;
        RECT 36.125 113.105 36.400 113.805 ;
        RECT 36.570 113.430 36.825 113.975 ;
        RECT 36.995 113.465 37.475 113.805 ;
        RECT 37.650 113.420 38.255 113.975 ;
        RECT 37.640 113.320 38.255 113.420 ;
        RECT 37.640 113.295 37.825 113.320 ;
        RECT 33.825 111.425 35.495 112.195 ;
        RECT 35.665 111.425 35.955 112.150 ;
        RECT 36.125 112.075 36.295 113.105 ;
        RECT 36.570 112.975 37.325 113.225 ;
        RECT 37.495 113.050 37.825 113.295 ;
        RECT 38.515 113.305 38.685 113.805 ;
        RECT 38.855 113.475 39.185 113.975 ;
        RECT 36.570 112.940 37.340 112.975 ;
        RECT 36.570 112.930 37.355 112.940 ;
        RECT 36.465 112.915 37.360 112.930 ;
        RECT 36.465 112.900 37.380 112.915 ;
        RECT 36.465 112.890 37.400 112.900 ;
        RECT 36.465 112.880 37.425 112.890 ;
        RECT 36.465 112.850 37.495 112.880 ;
        RECT 36.465 112.820 37.515 112.850 ;
        RECT 36.465 112.790 37.535 112.820 ;
        RECT 36.465 112.765 37.565 112.790 ;
        RECT 36.465 112.730 37.600 112.765 ;
        RECT 36.465 112.725 37.630 112.730 ;
        RECT 36.465 112.330 36.695 112.725 ;
        RECT 37.240 112.720 37.630 112.725 ;
        RECT 37.265 112.710 37.630 112.720 ;
        RECT 37.280 112.705 37.630 112.710 ;
        RECT 37.295 112.700 37.630 112.705 ;
        RECT 37.995 112.700 38.255 113.150 ;
        RECT 38.515 113.135 39.180 113.305 ;
        RECT 37.295 112.695 38.255 112.700 ;
        RECT 37.305 112.685 38.255 112.695 ;
        RECT 37.315 112.680 38.255 112.685 ;
        RECT 37.325 112.670 38.255 112.680 ;
        RECT 37.330 112.660 38.255 112.670 ;
        RECT 37.335 112.655 38.255 112.660 ;
        RECT 37.345 112.640 38.255 112.655 ;
        RECT 37.350 112.625 38.255 112.640 ;
        RECT 37.360 112.600 38.255 112.625 ;
        RECT 36.865 112.130 37.195 112.555 ;
        RECT 36.125 111.595 36.385 112.075 ;
        RECT 36.555 111.425 36.805 111.965 ;
        RECT 36.975 111.645 37.195 112.130 ;
        RECT 37.365 112.530 38.255 112.600 ;
        RECT 37.365 111.805 37.535 112.530 ;
        RECT 37.705 111.975 38.255 112.360 ;
        RECT 38.430 112.315 38.780 112.965 ;
        RECT 38.950 112.145 39.180 113.135 ;
        RECT 38.515 111.975 39.180 112.145 ;
        RECT 37.365 111.635 38.255 111.805 ;
        RECT 38.515 111.685 38.685 111.975 ;
        RECT 38.855 111.425 39.185 111.805 ;
        RECT 39.355 111.685 39.540 113.805 ;
        RECT 39.780 113.515 40.045 113.975 ;
        RECT 40.215 113.380 40.465 113.805 ;
        RECT 40.675 113.530 41.780 113.700 ;
        RECT 40.160 113.250 40.465 113.380 ;
        RECT 39.710 112.055 39.990 113.005 ;
        RECT 40.160 112.145 40.330 113.250 ;
        RECT 40.500 112.465 40.740 113.060 ;
        RECT 40.910 112.995 41.440 113.360 ;
        RECT 40.910 112.295 41.080 112.995 ;
        RECT 41.610 112.915 41.780 113.530 ;
        RECT 41.950 113.175 42.120 113.975 ;
        RECT 42.290 113.475 42.540 113.805 ;
        RECT 42.765 113.505 43.650 113.675 ;
        RECT 41.610 112.825 42.120 112.915 ;
        RECT 40.160 112.015 40.385 112.145 ;
        RECT 40.555 112.075 41.080 112.295 ;
        RECT 41.250 112.655 42.120 112.825 ;
        RECT 39.795 111.425 40.045 111.885 ;
        RECT 40.215 111.875 40.385 112.015 ;
        RECT 41.250 111.875 41.420 112.655 ;
        RECT 41.950 112.585 42.120 112.655 ;
        RECT 41.630 112.405 41.830 112.435 ;
        RECT 42.290 112.405 42.460 113.475 ;
        RECT 42.630 112.585 42.820 113.305 ;
        RECT 41.630 112.105 42.460 112.405 ;
        RECT 42.990 112.375 43.310 113.335 ;
        RECT 40.215 111.705 40.550 111.875 ;
        RECT 40.745 111.705 41.420 111.875 ;
        RECT 41.740 111.425 42.110 111.925 ;
        RECT 42.290 111.875 42.460 112.105 ;
        RECT 42.845 112.045 43.310 112.375 ;
        RECT 43.480 112.665 43.650 113.505 ;
        RECT 43.830 113.475 44.145 113.975 ;
        RECT 44.375 113.245 44.715 113.805 ;
        RECT 43.820 112.870 44.715 113.245 ;
        RECT 44.885 112.965 45.055 113.975 ;
        RECT 44.525 112.665 44.715 112.870 ;
        RECT 45.225 112.915 45.555 113.760 ;
        RECT 45.225 112.835 45.615 112.915 ;
        RECT 45.785 112.885 46.995 113.975 ;
        RECT 45.400 112.785 45.615 112.835 ;
        RECT 43.480 112.335 44.355 112.665 ;
        RECT 44.525 112.335 45.275 112.665 ;
        RECT 43.480 111.875 43.650 112.335 ;
        RECT 44.525 112.165 44.725 112.335 ;
        RECT 45.445 112.205 45.615 112.785 ;
        RECT 45.390 112.165 45.615 112.205 ;
        RECT 42.290 111.705 42.695 111.875 ;
        RECT 42.865 111.705 43.650 111.875 ;
        RECT 43.925 111.425 44.135 111.955 ;
        RECT 44.395 111.640 44.725 112.165 ;
        RECT 45.235 112.080 45.615 112.165 ;
        RECT 45.785 112.175 46.305 112.715 ;
        RECT 46.475 112.345 46.995 112.885 ;
        RECT 47.175 112.835 47.505 113.975 ;
        RECT 48.035 113.005 48.365 113.790 ;
        RECT 47.685 112.835 48.365 113.005 ;
        RECT 48.545 112.885 51.135 113.975 ;
        RECT 47.165 112.415 47.515 112.665 ;
        RECT 47.685 112.235 47.855 112.835 ;
        RECT 48.025 112.415 48.375 112.665 ;
        RECT 44.895 111.425 45.065 112.035 ;
        RECT 45.235 111.645 45.565 112.080 ;
        RECT 45.785 111.425 46.995 112.175 ;
        RECT 47.175 111.425 47.445 112.235 ;
        RECT 47.615 111.595 47.945 112.235 ;
        RECT 48.115 111.425 48.355 112.235 ;
        RECT 48.545 112.195 49.755 112.715 ;
        RECT 49.925 112.365 51.135 112.885 ;
        RECT 51.305 112.835 51.690 113.805 ;
        RECT 51.860 113.515 52.185 113.975 ;
        RECT 52.705 113.345 52.985 113.805 ;
        RECT 51.860 113.125 52.985 113.345 ;
        RECT 48.545 111.425 51.135 112.195 ;
        RECT 51.305 112.165 51.585 112.835 ;
        RECT 51.860 112.665 52.310 113.125 ;
        RECT 53.175 112.955 53.575 113.805 ;
        RECT 53.975 113.515 54.245 113.975 ;
        RECT 54.415 113.345 54.700 113.805 ;
        RECT 51.755 112.335 52.310 112.665 ;
        RECT 52.480 112.395 53.575 112.955 ;
        RECT 51.860 112.225 52.310 112.335 ;
        RECT 51.305 111.595 51.690 112.165 ;
        RECT 51.860 112.055 52.985 112.225 ;
        RECT 51.860 111.425 52.185 111.885 ;
        RECT 52.705 111.595 52.985 112.055 ;
        RECT 53.175 111.595 53.575 112.395 ;
        RECT 53.745 113.125 54.700 113.345 ;
        RECT 53.745 112.225 53.955 113.125 ;
        RECT 54.985 113.105 55.260 113.805 ;
        RECT 55.430 113.430 55.685 113.975 ;
        RECT 55.855 113.465 56.335 113.805 ;
        RECT 56.510 113.420 57.115 113.975 ;
        RECT 56.500 113.320 57.115 113.420 ;
        RECT 56.500 113.295 56.685 113.320 ;
        RECT 54.125 112.395 54.815 112.955 ;
        RECT 53.745 112.055 54.700 112.225 ;
        RECT 53.975 111.425 54.245 111.885 ;
        RECT 54.415 111.595 54.700 112.055 ;
        RECT 54.985 112.075 55.155 113.105 ;
        RECT 55.430 112.975 56.185 113.225 ;
        RECT 56.355 113.050 56.685 113.295 ;
        RECT 55.430 112.940 56.200 112.975 ;
        RECT 55.430 112.930 56.215 112.940 ;
        RECT 55.325 112.915 56.220 112.930 ;
        RECT 55.325 112.900 56.240 112.915 ;
        RECT 55.325 112.890 56.260 112.900 ;
        RECT 55.325 112.880 56.285 112.890 ;
        RECT 55.325 112.850 56.355 112.880 ;
        RECT 55.325 112.820 56.375 112.850 ;
        RECT 55.325 112.790 56.395 112.820 ;
        RECT 55.325 112.765 56.425 112.790 ;
        RECT 55.325 112.730 56.460 112.765 ;
        RECT 55.325 112.725 56.490 112.730 ;
        RECT 55.325 112.330 55.555 112.725 ;
        RECT 56.100 112.720 56.490 112.725 ;
        RECT 56.125 112.710 56.490 112.720 ;
        RECT 56.140 112.705 56.490 112.710 ;
        RECT 56.155 112.700 56.490 112.705 ;
        RECT 56.855 112.700 57.115 113.150 ;
        RECT 57.295 113.005 57.625 113.805 ;
        RECT 57.795 113.175 58.025 113.975 ;
        RECT 58.195 113.005 58.525 113.805 ;
        RECT 57.295 112.835 58.525 113.005 ;
        RECT 58.695 112.835 58.950 113.975 ;
        RECT 59.125 112.885 60.795 113.975 ;
        RECT 56.155 112.695 57.115 112.700 ;
        RECT 56.165 112.685 57.115 112.695 ;
        RECT 56.175 112.680 57.115 112.685 ;
        RECT 56.185 112.670 57.115 112.680 ;
        RECT 56.190 112.660 57.115 112.670 ;
        RECT 56.195 112.655 57.115 112.660 ;
        RECT 56.205 112.640 57.115 112.655 ;
        RECT 56.210 112.625 57.115 112.640 ;
        RECT 56.220 112.600 57.115 112.625 ;
        RECT 55.725 112.130 56.055 112.555 ;
        RECT 55.805 112.105 56.055 112.130 ;
        RECT 54.985 111.595 55.245 112.075 ;
        RECT 55.415 111.425 55.665 111.965 ;
        RECT 55.835 111.645 56.055 112.105 ;
        RECT 56.225 112.530 57.115 112.600 ;
        RECT 56.225 111.805 56.395 112.530 ;
        RECT 56.565 111.975 57.115 112.360 ;
        RECT 57.285 112.335 57.595 112.665 ;
        RECT 57.295 111.935 57.625 112.165 ;
        RECT 57.800 112.105 58.175 112.665 ;
        RECT 58.345 111.935 58.525 112.835 ;
        RECT 58.710 112.085 58.930 112.665 ;
        RECT 59.125 112.195 59.875 112.715 ;
        RECT 60.045 112.365 60.795 112.885 ;
        RECT 61.425 112.810 61.715 113.975 ;
        RECT 61.885 113.305 62.200 113.805 ;
        RECT 62.370 113.475 62.620 113.975 ;
        RECT 62.790 113.305 63.040 113.805 ;
        RECT 63.210 113.475 63.460 113.975 ;
        RECT 63.630 113.305 63.880 113.805 ;
        RECT 64.190 113.465 64.440 113.805 ;
        RECT 64.610 113.475 64.860 113.975 ;
        RECT 65.030 113.635 66.155 113.805 ;
        RECT 65.030 113.465 65.355 113.635 ;
        RECT 65.905 113.475 66.155 113.635 ;
        RECT 66.425 113.475 66.675 113.975 ;
        RECT 61.885 113.295 63.880 113.305 ;
        RECT 65.525 113.305 65.735 113.465 ;
        RECT 66.845 113.305 67.095 113.465 ;
        RECT 61.885 113.125 65.280 113.295 ;
        RECT 65.525 113.135 67.095 113.305 ;
        RECT 67.265 113.135 67.695 113.975 ;
        RECT 61.885 112.235 62.115 113.125 ;
        RECT 65.110 112.965 65.280 113.125 ;
        RECT 66.845 112.965 67.095 113.135 ;
        RECT 62.590 112.785 64.900 112.955 ;
        RECT 65.110 112.795 66.605 112.965 ;
        RECT 62.590 112.625 62.760 112.785 ;
        RECT 62.285 112.415 62.760 112.625 ;
        RECT 64.730 112.625 64.900 112.785 ;
        RECT 63.055 112.415 64.505 112.615 ;
        RECT 64.730 112.415 65.755 112.625 ;
        RECT 66.435 112.585 66.605 112.795 ;
        RECT 66.845 112.755 67.695 112.965 ;
        RECT 67.925 112.915 68.255 113.760 ;
        RECT 68.425 112.965 68.595 113.975 ;
        RECT 68.765 113.245 69.105 113.805 ;
        RECT 69.335 113.475 69.650 113.975 ;
        RECT 69.830 113.505 70.715 113.675 ;
        RECT 66.435 112.415 67.095 112.585 ;
        RECT 56.225 111.635 57.115 111.805 ;
        RECT 57.295 111.595 58.525 111.935 ;
        RECT 58.695 111.425 58.950 111.915 ;
        RECT 59.125 111.425 60.795 112.195 ;
        RECT 61.425 111.425 61.715 112.150 ;
        RECT 61.885 111.985 62.660 112.235 ;
        RECT 62.830 112.065 63.920 112.245 ;
        RECT 62.830 111.815 63.080 112.065 ;
        RECT 61.905 111.595 63.080 111.815 ;
        RECT 63.250 111.425 63.420 111.895 ;
        RECT 63.590 111.595 63.920 112.065 ;
        RECT 64.230 111.425 64.400 112.245 ;
        RECT 64.570 112.065 67.135 112.245 ;
        RECT 64.570 111.595 64.900 112.065 ;
        RECT 65.070 111.425 65.240 111.895 ;
        RECT 65.410 111.595 65.775 112.065 ;
        RECT 66.805 111.985 67.135 112.065 ;
        RECT 65.945 111.425 66.115 111.895 ;
        RECT 67.305 111.815 67.695 112.755 ;
        RECT 67.865 112.835 68.255 112.915 ;
        RECT 68.765 112.870 69.660 113.245 ;
        RECT 67.865 112.785 68.080 112.835 ;
        RECT 67.865 112.205 68.035 112.785 ;
        RECT 68.765 112.665 68.955 112.870 ;
        RECT 69.830 112.665 70.000 113.505 ;
        RECT 70.940 113.475 71.190 113.805 ;
        RECT 68.205 112.335 68.955 112.665 ;
        RECT 69.125 112.335 70.000 112.665 ;
        RECT 67.865 112.165 68.090 112.205 ;
        RECT 68.755 112.165 68.955 112.335 ;
        RECT 67.865 112.080 68.245 112.165 ;
        RECT 66.385 111.645 67.695 111.815 ;
        RECT 67.915 111.645 68.245 112.080 ;
        RECT 68.415 111.425 68.585 112.035 ;
        RECT 68.755 111.640 69.085 112.165 ;
        RECT 69.345 111.425 69.555 111.955 ;
        RECT 69.830 111.875 70.000 112.335 ;
        RECT 70.170 112.375 70.490 113.335 ;
        RECT 70.660 112.585 70.850 113.305 ;
        RECT 71.020 112.405 71.190 113.475 ;
        RECT 71.360 113.175 71.530 113.975 ;
        RECT 71.700 113.530 72.805 113.700 ;
        RECT 71.700 112.915 71.870 113.530 ;
        RECT 73.015 113.380 73.265 113.805 ;
        RECT 73.435 113.515 73.700 113.975 ;
        RECT 72.040 112.995 72.570 113.360 ;
        RECT 73.015 113.250 73.320 113.380 ;
        RECT 71.360 112.825 71.870 112.915 ;
        RECT 71.360 112.655 72.230 112.825 ;
        RECT 71.360 112.585 71.530 112.655 ;
        RECT 71.650 112.405 71.850 112.435 ;
        RECT 70.170 112.045 70.635 112.375 ;
        RECT 71.020 112.105 71.850 112.405 ;
        RECT 71.020 111.875 71.190 112.105 ;
        RECT 69.830 111.705 70.615 111.875 ;
        RECT 70.785 111.705 71.190 111.875 ;
        RECT 71.370 111.425 71.740 111.925 ;
        RECT 72.060 111.875 72.230 112.655 ;
        RECT 72.400 112.295 72.570 112.995 ;
        RECT 72.740 112.465 72.980 113.060 ;
        RECT 72.400 112.075 72.925 112.295 ;
        RECT 73.150 112.145 73.320 113.250 ;
        RECT 73.095 112.015 73.320 112.145 ;
        RECT 73.490 112.055 73.770 113.005 ;
        RECT 73.095 111.875 73.265 112.015 ;
        RECT 72.060 111.705 72.735 111.875 ;
        RECT 72.930 111.705 73.265 111.875 ;
        RECT 73.435 111.425 73.685 111.885 ;
        RECT 73.940 111.685 74.125 113.805 ;
        RECT 74.295 113.475 74.625 113.975 ;
        RECT 74.795 113.305 74.965 113.805 ;
        RECT 75.225 113.540 80.570 113.975 ;
        RECT 74.300 113.135 74.965 113.305 ;
        RECT 74.300 112.145 74.530 113.135 ;
        RECT 74.700 112.315 75.050 112.965 ;
        RECT 74.300 111.975 74.965 112.145 ;
        RECT 74.295 111.425 74.625 111.805 ;
        RECT 74.795 111.685 74.965 111.975 ;
        RECT 76.810 111.970 77.150 112.800 ;
        RECT 78.630 112.290 78.980 113.540 ;
        RECT 75.225 111.425 80.570 111.970 ;
        RECT 80.755 111.605 81.015 113.795 ;
        RECT 81.185 113.245 81.525 113.975 ;
        RECT 81.705 113.065 81.975 113.795 ;
        RECT 81.205 112.845 81.975 113.065 ;
        RECT 82.155 113.085 82.385 113.795 ;
        RECT 82.555 113.265 82.885 113.975 ;
        RECT 83.055 113.085 83.315 113.795 ;
        RECT 82.155 112.845 83.315 113.085 ;
        RECT 83.505 113.105 83.780 113.805 ;
        RECT 83.950 113.430 84.205 113.975 ;
        RECT 84.375 113.465 84.855 113.805 ;
        RECT 85.030 113.420 85.635 113.975 ;
        RECT 85.020 113.320 85.635 113.420 ;
        RECT 85.020 113.295 85.205 113.320 ;
        RECT 81.205 112.175 81.495 112.845 ;
        RECT 81.675 112.355 82.140 112.665 ;
        RECT 82.320 112.355 82.845 112.665 ;
        RECT 81.205 111.975 82.435 112.175 ;
        RECT 81.275 111.425 81.945 111.795 ;
        RECT 82.125 111.605 82.435 111.975 ;
        RECT 82.615 111.715 82.845 112.355 ;
        RECT 83.025 112.335 83.325 112.665 ;
        RECT 83.025 111.425 83.315 112.155 ;
        RECT 83.505 112.075 83.675 113.105 ;
        RECT 83.950 112.975 84.705 113.225 ;
        RECT 84.875 113.050 85.205 113.295 ;
        RECT 83.950 112.940 84.720 112.975 ;
        RECT 83.950 112.930 84.735 112.940 ;
        RECT 83.845 112.915 84.740 112.930 ;
        RECT 83.845 112.900 84.760 112.915 ;
        RECT 83.845 112.890 84.780 112.900 ;
        RECT 83.845 112.880 84.805 112.890 ;
        RECT 83.845 112.850 84.875 112.880 ;
        RECT 83.845 112.820 84.895 112.850 ;
        RECT 83.845 112.790 84.915 112.820 ;
        RECT 83.845 112.765 84.945 112.790 ;
        RECT 83.845 112.730 84.980 112.765 ;
        RECT 83.845 112.725 85.010 112.730 ;
        RECT 83.845 112.330 84.075 112.725 ;
        RECT 84.620 112.720 85.010 112.725 ;
        RECT 84.645 112.710 85.010 112.720 ;
        RECT 84.660 112.705 85.010 112.710 ;
        RECT 84.675 112.700 85.010 112.705 ;
        RECT 85.375 112.700 85.635 113.150 ;
        RECT 85.805 112.885 87.015 113.975 ;
        RECT 84.675 112.695 85.635 112.700 ;
        RECT 84.685 112.685 85.635 112.695 ;
        RECT 84.695 112.680 85.635 112.685 ;
        RECT 84.705 112.670 85.635 112.680 ;
        RECT 84.710 112.660 85.635 112.670 ;
        RECT 84.715 112.655 85.635 112.660 ;
        RECT 84.725 112.640 85.635 112.655 ;
        RECT 84.730 112.625 85.635 112.640 ;
        RECT 84.740 112.600 85.635 112.625 ;
        RECT 84.245 112.130 84.575 112.555 ;
        RECT 83.505 111.595 83.765 112.075 ;
        RECT 83.935 111.425 84.185 111.965 ;
        RECT 84.355 111.645 84.575 112.130 ;
        RECT 84.745 112.530 85.635 112.600 ;
        RECT 84.745 111.805 84.915 112.530 ;
        RECT 85.085 111.975 85.635 112.360 ;
        RECT 85.805 112.175 86.325 112.715 ;
        RECT 86.495 112.345 87.015 112.885 ;
        RECT 87.185 112.810 87.475 113.975 ;
        RECT 87.645 112.885 91.155 113.975 ;
        RECT 91.325 113.420 91.930 113.975 ;
        RECT 92.105 113.465 92.585 113.805 ;
        RECT 92.755 113.430 93.010 113.975 ;
        RECT 91.325 113.320 91.940 113.420 ;
        RECT 91.755 113.295 91.940 113.320 ;
        RECT 87.645 112.195 89.295 112.715 ;
        RECT 89.465 112.365 91.155 112.885 ;
        RECT 91.325 112.700 91.585 113.150 ;
        RECT 91.755 113.050 92.085 113.295 ;
        RECT 92.255 112.975 93.010 113.225 ;
        RECT 93.180 113.105 93.455 113.805 ;
        RECT 93.715 113.305 93.885 113.805 ;
        RECT 94.055 113.475 94.385 113.975 ;
        RECT 93.715 113.135 94.380 113.305 ;
        RECT 92.240 112.940 93.010 112.975 ;
        RECT 92.225 112.930 93.010 112.940 ;
        RECT 92.220 112.915 93.115 112.930 ;
        RECT 92.200 112.900 93.115 112.915 ;
        RECT 92.180 112.890 93.115 112.900 ;
        RECT 92.155 112.880 93.115 112.890 ;
        RECT 92.085 112.850 93.115 112.880 ;
        RECT 92.065 112.820 93.115 112.850 ;
        RECT 92.045 112.790 93.115 112.820 ;
        RECT 92.015 112.765 93.115 112.790 ;
        RECT 91.980 112.730 93.115 112.765 ;
        RECT 91.950 112.725 93.115 112.730 ;
        RECT 91.950 112.720 92.340 112.725 ;
        RECT 91.950 112.710 92.315 112.720 ;
        RECT 91.950 112.705 92.300 112.710 ;
        RECT 91.950 112.700 92.285 112.705 ;
        RECT 91.325 112.695 92.285 112.700 ;
        RECT 91.325 112.685 92.275 112.695 ;
        RECT 91.325 112.680 92.265 112.685 ;
        RECT 91.325 112.670 92.255 112.680 ;
        RECT 91.325 112.660 92.250 112.670 ;
        RECT 91.325 112.655 92.245 112.660 ;
        RECT 91.325 112.640 92.235 112.655 ;
        RECT 91.325 112.625 92.230 112.640 ;
        RECT 91.325 112.600 92.220 112.625 ;
        RECT 91.325 112.530 92.215 112.600 ;
        RECT 84.745 111.635 85.635 111.805 ;
        RECT 85.805 111.425 87.015 112.175 ;
        RECT 87.185 111.425 87.475 112.150 ;
        RECT 87.645 111.425 91.155 112.195 ;
        RECT 91.325 111.975 91.875 112.360 ;
        RECT 92.045 111.805 92.215 112.530 ;
        RECT 91.325 111.635 92.215 111.805 ;
        RECT 92.385 112.130 92.715 112.555 ;
        RECT 92.885 112.330 93.115 112.725 ;
        RECT 92.385 111.645 92.605 112.130 ;
        RECT 93.285 112.075 93.455 113.105 ;
        RECT 93.630 112.315 93.980 112.965 ;
        RECT 94.150 112.145 94.380 113.135 ;
        RECT 92.775 111.425 93.025 111.965 ;
        RECT 93.195 111.595 93.455 112.075 ;
        RECT 93.715 111.975 94.380 112.145 ;
        RECT 93.715 111.685 93.885 111.975 ;
        RECT 94.055 111.425 94.385 111.805 ;
        RECT 94.555 111.685 94.740 113.805 ;
        RECT 94.980 113.515 95.245 113.975 ;
        RECT 95.415 113.380 95.665 113.805 ;
        RECT 95.875 113.530 96.980 113.700 ;
        RECT 95.360 113.250 95.665 113.380 ;
        RECT 94.910 112.055 95.190 113.005 ;
        RECT 95.360 112.145 95.530 113.250 ;
        RECT 95.700 112.465 95.940 113.060 ;
        RECT 96.110 112.995 96.640 113.360 ;
        RECT 96.110 112.295 96.280 112.995 ;
        RECT 96.810 112.915 96.980 113.530 ;
        RECT 97.150 113.175 97.320 113.975 ;
        RECT 97.490 113.475 97.740 113.805 ;
        RECT 97.965 113.505 98.850 113.675 ;
        RECT 96.810 112.825 97.320 112.915 ;
        RECT 95.360 112.015 95.585 112.145 ;
        RECT 95.755 112.075 96.280 112.295 ;
        RECT 96.450 112.655 97.320 112.825 ;
        RECT 94.995 111.425 95.245 111.885 ;
        RECT 95.415 111.875 95.585 112.015 ;
        RECT 96.450 111.875 96.620 112.655 ;
        RECT 97.150 112.585 97.320 112.655 ;
        RECT 96.830 112.405 97.030 112.435 ;
        RECT 97.490 112.405 97.660 113.475 ;
        RECT 97.830 112.585 98.020 113.305 ;
        RECT 96.830 112.105 97.660 112.405 ;
        RECT 98.190 112.375 98.510 113.335 ;
        RECT 95.415 111.705 95.750 111.875 ;
        RECT 95.945 111.705 96.620 111.875 ;
        RECT 96.940 111.425 97.310 111.925 ;
        RECT 97.490 111.875 97.660 112.105 ;
        RECT 98.045 112.045 98.510 112.375 ;
        RECT 98.680 112.665 98.850 113.505 ;
        RECT 99.030 113.475 99.345 113.975 ;
        RECT 99.575 113.245 99.915 113.805 ;
        RECT 99.020 112.870 99.915 113.245 ;
        RECT 100.085 112.965 100.255 113.975 ;
        RECT 99.725 112.665 99.915 112.870 ;
        RECT 100.425 112.915 100.755 113.760 ;
        RECT 100.925 113.060 101.095 113.975 ;
        RECT 102.455 113.305 102.625 113.805 ;
        RECT 102.795 113.475 103.125 113.975 ;
        RECT 102.455 113.135 103.120 113.305 ;
        RECT 100.425 112.835 100.815 112.915 ;
        RECT 100.600 112.785 100.815 112.835 ;
        RECT 98.680 112.335 99.555 112.665 ;
        RECT 99.725 112.335 100.475 112.665 ;
        RECT 98.680 111.875 98.850 112.335 ;
        RECT 99.725 112.165 99.925 112.335 ;
        RECT 100.645 112.205 100.815 112.785 ;
        RECT 102.370 112.315 102.720 112.965 ;
        RECT 100.590 112.165 100.815 112.205 ;
        RECT 97.490 111.705 97.895 111.875 ;
        RECT 98.065 111.705 98.850 111.875 ;
        RECT 99.125 111.425 99.335 111.955 ;
        RECT 99.595 111.640 99.925 112.165 ;
        RECT 100.435 112.080 100.815 112.165 ;
        RECT 102.890 112.145 103.120 113.135 ;
        RECT 100.095 111.425 100.265 112.035 ;
        RECT 100.435 111.645 100.765 112.080 ;
        RECT 102.455 111.975 103.120 112.145 ;
        RECT 100.935 111.425 101.105 111.940 ;
        RECT 102.455 111.685 102.625 111.975 ;
        RECT 102.795 111.425 103.125 111.805 ;
        RECT 103.295 111.685 103.480 113.805 ;
        RECT 103.720 113.515 103.985 113.975 ;
        RECT 104.155 113.380 104.405 113.805 ;
        RECT 104.615 113.530 105.720 113.700 ;
        RECT 104.100 113.250 104.405 113.380 ;
        RECT 103.650 112.055 103.930 113.005 ;
        RECT 104.100 112.145 104.270 113.250 ;
        RECT 104.440 112.465 104.680 113.060 ;
        RECT 104.850 112.995 105.380 113.360 ;
        RECT 104.850 112.295 105.020 112.995 ;
        RECT 105.550 112.915 105.720 113.530 ;
        RECT 105.890 113.175 106.060 113.975 ;
        RECT 106.230 113.475 106.480 113.805 ;
        RECT 106.705 113.505 107.590 113.675 ;
        RECT 105.550 112.825 106.060 112.915 ;
        RECT 104.100 112.015 104.325 112.145 ;
        RECT 104.495 112.075 105.020 112.295 ;
        RECT 105.190 112.655 106.060 112.825 ;
        RECT 103.735 111.425 103.985 111.885 ;
        RECT 104.155 111.875 104.325 112.015 ;
        RECT 105.190 111.875 105.360 112.655 ;
        RECT 105.890 112.585 106.060 112.655 ;
        RECT 105.570 112.405 105.770 112.435 ;
        RECT 106.230 112.405 106.400 113.475 ;
        RECT 106.570 112.585 106.760 113.305 ;
        RECT 105.570 112.105 106.400 112.405 ;
        RECT 106.930 112.375 107.250 113.335 ;
        RECT 104.155 111.705 104.490 111.875 ;
        RECT 104.685 111.705 105.360 111.875 ;
        RECT 105.680 111.425 106.050 111.925 ;
        RECT 106.230 111.875 106.400 112.105 ;
        RECT 106.785 112.045 107.250 112.375 ;
        RECT 107.420 112.665 107.590 113.505 ;
        RECT 107.770 113.475 108.085 113.975 ;
        RECT 108.315 113.245 108.655 113.805 ;
        RECT 107.760 112.870 108.655 113.245 ;
        RECT 108.825 112.965 108.995 113.975 ;
        RECT 108.465 112.665 108.655 112.870 ;
        RECT 109.165 112.915 109.495 113.760 ;
        RECT 109.725 113.105 110.000 113.805 ;
        RECT 110.170 113.430 110.425 113.975 ;
        RECT 110.595 113.465 111.075 113.805 ;
        RECT 111.250 113.420 111.855 113.975 ;
        RECT 111.240 113.320 111.855 113.420 ;
        RECT 111.240 113.295 111.425 113.320 ;
        RECT 109.165 112.835 109.555 112.915 ;
        RECT 109.340 112.785 109.555 112.835 ;
        RECT 107.420 112.335 108.295 112.665 ;
        RECT 108.465 112.335 109.215 112.665 ;
        RECT 107.420 111.875 107.590 112.335 ;
        RECT 108.465 112.165 108.665 112.335 ;
        RECT 109.385 112.205 109.555 112.785 ;
        RECT 109.330 112.165 109.555 112.205 ;
        RECT 106.230 111.705 106.635 111.875 ;
        RECT 106.805 111.705 107.590 111.875 ;
        RECT 107.865 111.425 108.075 111.955 ;
        RECT 108.335 111.640 108.665 112.165 ;
        RECT 109.175 112.080 109.555 112.165 ;
        RECT 108.835 111.425 109.005 112.035 ;
        RECT 109.175 111.645 109.505 112.080 ;
        RECT 109.725 112.075 109.895 113.105 ;
        RECT 110.170 112.975 110.925 113.225 ;
        RECT 111.095 113.050 111.425 113.295 ;
        RECT 110.170 112.940 110.940 112.975 ;
        RECT 110.170 112.930 110.955 112.940 ;
        RECT 110.065 112.915 110.960 112.930 ;
        RECT 110.065 112.900 110.980 112.915 ;
        RECT 110.065 112.890 111.000 112.900 ;
        RECT 110.065 112.880 111.025 112.890 ;
        RECT 110.065 112.850 111.095 112.880 ;
        RECT 110.065 112.820 111.115 112.850 ;
        RECT 110.065 112.790 111.135 112.820 ;
        RECT 110.065 112.765 111.165 112.790 ;
        RECT 110.065 112.730 111.200 112.765 ;
        RECT 110.065 112.725 111.230 112.730 ;
        RECT 110.065 112.330 110.295 112.725 ;
        RECT 110.840 112.720 111.230 112.725 ;
        RECT 110.865 112.710 111.230 112.720 ;
        RECT 110.880 112.705 111.230 112.710 ;
        RECT 110.895 112.700 111.230 112.705 ;
        RECT 111.595 112.700 111.855 113.150 ;
        RECT 112.945 112.810 113.235 113.975 ;
        RECT 113.405 112.885 114.615 113.975 ;
        RECT 110.895 112.695 111.855 112.700 ;
        RECT 110.905 112.685 111.855 112.695 ;
        RECT 110.915 112.680 111.855 112.685 ;
        RECT 110.925 112.670 111.855 112.680 ;
        RECT 110.930 112.660 111.855 112.670 ;
        RECT 110.935 112.655 111.855 112.660 ;
        RECT 110.945 112.640 111.855 112.655 ;
        RECT 110.950 112.625 111.855 112.640 ;
        RECT 110.960 112.600 111.855 112.625 ;
        RECT 110.465 112.130 110.795 112.555 ;
        RECT 109.725 111.595 109.985 112.075 ;
        RECT 110.155 111.425 110.405 111.965 ;
        RECT 110.575 111.645 110.795 112.130 ;
        RECT 110.965 112.530 111.855 112.600 ;
        RECT 110.965 111.805 111.135 112.530 ;
        RECT 111.305 111.975 111.855 112.360 ;
        RECT 113.405 112.175 113.925 112.715 ;
        RECT 114.095 112.345 114.615 112.885 ;
        RECT 114.785 113.105 115.060 113.805 ;
        RECT 115.230 113.430 115.485 113.975 ;
        RECT 115.655 113.465 116.135 113.805 ;
        RECT 116.310 113.420 116.915 113.975 ;
        RECT 116.300 113.320 116.915 113.420 ;
        RECT 116.300 113.295 116.485 113.320 ;
        RECT 110.965 111.635 111.855 111.805 ;
        RECT 112.945 111.425 113.235 112.150 ;
        RECT 113.405 111.425 114.615 112.175 ;
        RECT 114.785 112.075 114.955 113.105 ;
        RECT 115.230 112.975 115.985 113.225 ;
        RECT 116.155 113.050 116.485 113.295 ;
        RECT 115.230 112.940 116.000 112.975 ;
        RECT 115.230 112.930 116.015 112.940 ;
        RECT 115.125 112.915 116.020 112.930 ;
        RECT 115.125 112.900 116.040 112.915 ;
        RECT 115.125 112.890 116.060 112.900 ;
        RECT 115.125 112.880 116.085 112.890 ;
        RECT 115.125 112.850 116.155 112.880 ;
        RECT 115.125 112.820 116.175 112.850 ;
        RECT 115.125 112.790 116.195 112.820 ;
        RECT 115.125 112.765 116.225 112.790 ;
        RECT 115.125 112.730 116.260 112.765 ;
        RECT 115.125 112.725 116.290 112.730 ;
        RECT 115.125 112.330 115.355 112.725 ;
        RECT 115.900 112.720 116.290 112.725 ;
        RECT 115.925 112.710 116.290 112.720 ;
        RECT 115.940 112.705 116.290 112.710 ;
        RECT 115.955 112.700 116.290 112.705 ;
        RECT 116.655 112.700 116.915 113.150 ;
        RECT 117.605 112.835 117.815 113.975 ;
        RECT 115.955 112.695 116.915 112.700 ;
        RECT 115.965 112.685 116.915 112.695 ;
        RECT 115.975 112.680 116.915 112.685 ;
        RECT 115.985 112.670 116.915 112.680 ;
        RECT 115.990 112.660 116.915 112.670 ;
        RECT 115.995 112.655 116.915 112.660 ;
        RECT 116.005 112.640 116.915 112.655 ;
        RECT 116.010 112.625 116.915 112.640 ;
        RECT 116.020 112.600 116.915 112.625 ;
        RECT 115.525 112.130 115.855 112.555 ;
        RECT 114.785 111.595 115.045 112.075 ;
        RECT 115.215 111.425 115.465 111.965 ;
        RECT 115.635 111.645 115.855 112.130 ;
        RECT 116.025 112.530 116.915 112.600 ;
        RECT 117.985 112.825 118.315 113.805 ;
        RECT 118.485 112.835 118.715 113.975 ;
        RECT 119.960 113.345 120.245 113.805 ;
        RECT 120.415 113.515 120.685 113.975 ;
        RECT 119.960 113.125 120.915 113.345 ;
        RECT 116.025 111.805 116.195 112.530 ;
        RECT 116.365 111.975 116.915 112.360 ;
        RECT 116.025 111.635 116.915 111.805 ;
        RECT 117.605 111.425 117.815 112.245 ;
        RECT 117.985 112.225 118.235 112.825 ;
        RECT 118.405 112.415 118.735 112.665 ;
        RECT 119.845 112.395 120.535 112.955 ;
        RECT 117.985 111.595 118.315 112.225 ;
        RECT 118.485 111.425 118.715 112.245 ;
        RECT 120.705 112.225 120.915 113.125 ;
        RECT 119.960 112.055 120.915 112.225 ;
        RECT 121.085 112.955 121.485 113.805 ;
        RECT 121.675 113.345 121.955 113.805 ;
        RECT 122.475 113.515 122.800 113.975 ;
        RECT 121.675 113.125 122.800 113.345 ;
        RECT 121.085 112.395 122.180 112.955 ;
        RECT 122.350 112.665 122.800 113.125 ;
        RECT 122.970 112.835 123.355 113.805 ;
        RECT 123.530 113.175 123.785 113.975 ;
        RECT 123.985 113.125 124.315 113.805 ;
        RECT 119.960 111.595 120.245 112.055 ;
        RECT 120.415 111.425 120.685 111.885 ;
        RECT 121.085 111.595 121.485 112.395 ;
        RECT 122.350 112.335 122.905 112.665 ;
        RECT 122.350 112.225 122.800 112.335 ;
        RECT 121.675 112.055 122.800 112.225 ;
        RECT 123.075 112.165 123.355 112.835 ;
        RECT 123.530 112.635 123.775 112.995 ;
        RECT 123.965 112.845 124.315 113.125 ;
        RECT 123.965 112.465 124.135 112.845 ;
        RECT 124.495 112.665 124.690 113.715 ;
        RECT 124.870 112.835 125.190 113.975 ;
        RECT 125.365 112.885 127.035 113.975 ;
        RECT 121.675 111.595 121.955 112.055 ;
        RECT 122.475 111.425 122.800 111.885 ;
        RECT 122.970 111.595 123.355 112.165 ;
        RECT 123.615 112.295 124.135 112.465 ;
        RECT 124.305 112.335 124.690 112.665 ;
        RECT 124.870 112.615 125.130 112.665 ;
        RECT 124.870 112.445 125.135 112.615 ;
        RECT 124.870 112.335 125.130 112.445 ;
        RECT 123.615 111.935 123.785 112.295 ;
        RECT 125.365 112.195 126.115 112.715 ;
        RECT 126.285 112.365 127.035 112.885 ;
        RECT 127.670 112.835 127.925 113.975 ;
        RECT 128.095 113.005 128.425 113.805 ;
        RECT 128.595 113.175 128.825 113.975 ;
        RECT 128.995 113.005 129.325 113.805 ;
        RECT 128.095 112.835 129.325 113.005 ;
        RECT 129.690 113.005 130.080 113.180 ;
        RECT 130.565 113.175 130.895 113.975 ;
        RECT 131.065 113.185 131.600 113.805 ;
        RECT 129.690 112.835 131.115 113.005 ;
        RECT 123.585 111.765 123.785 111.935 ;
        RECT 123.615 111.730 123.785 111.765 ;
        RECT 123.975 111.955 125.190 112.125 ;
        RECT 123.975 111.650 124.205 111.955 ;
        RECT 124.375 111.425 124.705 111.785 ;
        RECT 124.900 111.605 125.190 111.955 ;
        RECT 125.365 111.425 127.035 112.195 ;
        RECT 127.690 112.085 127.910 112.665 ;
        RECT 128.095 111.935 128.275 112.835 ;
        RECT 128.445 112.105 128.820 112.665 ;
        RECT 129.025 112.335 129.335 112.665 ;
        RECT 128.995 111.935 129.325 112.165 ;
        RECT 129.565 112.105 129.920 112.665 ;
        RECT 130.090 111.935 130.260 112.835 ;
        RECT 130.430 112.105 130.695 112.665 ;
        RECT 130.945 112.335 131.115 112.835 ;
        RECT 131.285 112.165 131.600 113.185 ;
        RECT 132.010 113.005 132.340 113.805 ;
        RECT 132.510 113.175 132.840 113.975 ;
        RECT 133.140 113.005 133.470 113.805 ;
        RECT 134.115 113.175 134.365 113.975 ;
        RECT 132.010 112.835 134.445 113.005 ;
        RECT 134.635 112.835 134.805 113.975 ;
        RECT 134.975 112.835 135.315 113.805 ;
        RECT 136.130 113.005 136.520 113.180 ;
        RECT 137.005 113.175 137.335 113.975 ;
        RECT 137.505 113.185 138.040 113.805 ;
        RECT 136.130 112.835 137.555 113.005 ;
        RECT 131.805 112.415 132.155 112.665 ;
        RECT 132.340 112.205 132.510 112.835 ;
        RECT 132.680 112.415 133.010 112.615 ;
        RECT 133.180 112.415 133.510 112.615 ;
        RECT 133.680 112.415 134.100 112.615 ;
        RECT 134.275 112.585 134.445 112.835 ;
        RECT 134.275 112.415 134.970 112.585 ;
        RECT 127.670 111.425 127.925 111.915 ;
        RECT 128.095 111.595 129.325 111.935 ;
        RECT 129.670 111.425 129.910 111.935 ;
        RECT 130.090 111.605 130.370 111.935 ;
        RECT 130.600 111.425 130.815 111.935 ;
        RECT 130.985 111.595 131.600 112.165 ;
        RECT 132.010 111.595 132.510 112.205 ;
        RECT 133.140 112.075 134.365 112.245 ;
        RECT 135.140 112.225 135.315 112.835 ;
        RECT 133.140 111.595 133.470 112.075 ;
        RECT 133.640 111.425 133.865 111.885 ;
        RECT 134.035 111.595 134.365 112.075 ;
        RECT 134.555 111.425 134.805 112.225 ;
        RECT 134.975 111.595 135.315 112.225 ;
        RECT 136.005 112.105 136.360 112.665 ;
        RECT 136.530 111.935 136.700 112.835 ;
        RECT 136.870 112.105 137.135 112.665 ;
        RECT 137.385 112.335 137.555 112.835 ;
        RECT 137.725 112.165 138.040 113.185 ;
        RECT 138.705 112.810 138.995 113.975 ;
        RECT 139.165 112.835 139.550 113.805 ;
        RECT 139.720 113.515 140.045 113.975 ;
        RECT 140.565 113.345 140.845 113.805 ;
        RECT 139.720 113.125 140.845 113.345 ;
        RECT 136.110 111.425 136.350 111.935 ;
        RECT 136.530 111.605 136.810 111.935 ;
        RECT 137.040 111.425 137.255 111.935 ;
        RECT 137.425 111.595 138.040 112.165 ;
        RECT 139.165 112.165 139.445 112.835 ;
        RECT 139.720 112.665 140.170 113.125 ;
        RECT 141.035 112.955 141.435 113.805 ;
        RECT 141.835 113.515 142.105 113.975 ;
        RECT 142.275 113.345 142.560 113.805 ;
        RECT 139.615 112.335 140.170 112.665 ;
        RECT 140.340 112.395 141.435 112.955 ;
        RECT 139.720 112.225 140.170 112.335 ;
        RECT 138.705 111.425 138.995 112.150 ;
        RECT 139.165 111.595 139.550 112.165 ;
        RECT 139.720 112.055 140.845 112.225 ;
        RECT 139.720 111.425 140.045 111.885 ;
        RECT 140.565 111.595 140.845 112.055 ;
        RECT 141.035 111.595 141.435 112.395 ;
        RECT 141.605 113.125 142.560 113.345 ;
        RECT 141.605 112.225 141.815 113.125 ;
        RECT 141.985 112.395 142.675 112.955 ;
        RECT 142.850 112.825 143.110 113.975 ;
        RECT 143.285 112.900 143.540 113.805 ;
        RECT 143.710 113.215 144.040 113.975 ;
        RECT 144.255 113.045 144.425 113.805 ;
        RECT 141.605 112.055 142.560 112.225 ;
        RECT 141.835 111.425 142.105 111.885 ;
        RECT 142.275 111.595 142.560 112.055 ;
        RECT 142.850 111.425 143.110 112.265 ;
        RECT 143.285 112.170 143.455 112.900 ;
        RECT 143.710 112.875 144.425 113.045 ;
        RECT 144.890 113.005 145.220 113.805 ;
        RECT 145.390 113.175 145.720 113.975 ;
        RECT 146.020 113.005 146.350 113.805 ;
        RECT 146.995 113.175 147.245 113.975 ;
        RECT 143.710 112.665 143.880 112.875 ;
        RECT 144.890 112.835 147.325 113.005 ;
        RECT 147.515 112.835 147.685 113.975 ;
        RECT 147.855 112.835 148.195 113.805 ;
        RECT 148.455 113.305 148.625 113.805 ;
        RECT 148.795 113.475 149.125 113.975 ;
        RECT 148.455 113.135 149.120 113.305 ;
        RECT 143.625 112.335 143.880 112.665 ;
        RECT 143.285 111.595 143.540 112.170 ;
        RECT 143.710 112.145 143.880 112.335 ;
        RECT 144.160 112.325 144.515 112.695 ;
        RECT 144.685 112.415 145.035 112.665 ;
        RECT 145.220 112.205 145.390 112.835 ;
        RECT 145.560 112.415 145.890 112.615 ;
        RECT 146.060 112.415 146.390 112.615 ;
        RECT 146.560 112.415 146.980 112.615 ;
        RECT 147.155 112.585 147.325 112.835 ;
        RECT 147.155 112.415 147.850 112.585 ;
        RECT 148.020 112.275 148.195 112.835 ;
        RECT 148.370 112.315 148.720 112.965 ;
        RECT 143.710 111.975 144.425 112.145 ;
        RECT 143.710 111.425 144.040 111.805 ;
        RECT 144.255 111.595 144.425 111.975 ;
        RECT 144.890 111.595 145.390 112.205 ;
        RECT 146.020 112.075 147.245 112.245 ;
        RECT 147.965 112.225 148.195 112.275 ;
        RECT 146.020 111.595 146.350 112.075 ;
        RECT 146.520 111.425 146.745 111.885 ;
        RECT 146.915 111.595 147.245 112.075 ;
        RECT 147.435 111.425 147.685 112.225 ;
        RECT 147.855 111.595 148.195 112.225 ;
        RECT 148.890 112.145 149.120 113.135 ;
        RECT 148.455 111.975 149.120 112.145 ;
        RECT 148.455 111.685 148.625 111.975 ;
        RECT 148.795 111.425 149.125 111.805 ;
        RECT 149.295 111.685 149.480 113.805 ;
        RECT 149.720 113.515 149.985 113.975 ;
        RECT 150.155 113.380 150.405 113.805 ;
        RECT 150.615 113.530 151.720 113.700 ;
        RECT 150.100 113.250 150.405 113.380 ;
        RECT 149.650 112.055 149.930 113.005 ;
        RECT 150.100 112.145 150.270 113.250 ;
        RECT 150.440 112.465 150.680 113.060 ;
        RECT 150.850 112.995 151.380 113.360 ;
        RECT 150.850 112.295 151.020 112.995 ;
        RECT 151.550 112.915 151.720 113.530 ;
        RECT 151.890 113.175 152.060 113.975 ;
        RECT 152.230 113.475 152.480 113.805 ;
        RECT 152.705 113.505 153.590 113.675 ;
        RECT 151.550 112.825 152.060 112.915 ;
        RECT 150.100 112.015 150.325 112.145 ;
        RECT 150.495 112.075 151.020 112.295 ;
        RECT 151.190 112.655 152.060 112.825 ;
        RECT 149.735 111.425 149.985 111.885 ;
        RECT 150.155 111.875 150.325 112.015 ;
        RECT 151.190 111.875 151.360 112.655 ;
        RECT 151.890 112.585 152.060 112.655 ;
        RECT 151.570 112.405 151.770 112.435 ;
        RECT 152.230 112.405 152.400 113.475 ;
        RECT 152.570 112.585 152.760 113.305 ;
        RECT 151.570 112.105 152.400 112.405 ;
        RECT 152.930 112.375 153.250 113.335 ;
        RECT 150.155 111.705 150.490 111.875 ;
        RECT 150.685 111.705 151.360 111.875 ;
        RECT 151.680 111.425 152.050 111.925 ;
        RECT 152.230 111.875 152.400 112.105 ;
        RECT 152.785 112.045 153.250 112.375 ;
        RECT 153.420 112.665 153.590 113.505 ;
        RECT 153.770 113.475 154.085 113.975 ;
        RECT 154.315 113.245 154.655 113.805 ;
        RECT 153.760 112.870 154.655 113.245 ;
        RECT 154.825 112.965 154.995 113.975 ;
        RECT 154.465 112.665 154.655 112.870 ;
        RECT 155.165 112.915 155.495 113.760 ;
        RECT 155.165 112.835 155.555 112.915 ;
        RECT 155.340 112.785 155.555 112.835 ;
        RECT 153.420 112.335 154.295 112.665 ;
        RECT 154.465 112.335 155.215 112.665 ;
        RECT 153.420 111.875 153.590 112.335 ;
        RECT 154.465 112.165 154.665 112.335 ;
        RECT 155.385 112.205 155.555 112.785 ;
        RECT 155.725 112.885 156.935 113.975 ;
        RECT 155.725 112.345 156.245 112.885 ;
        RECT 155.330 112.165 155.555 112.205 ;
        RECT 156.415 112.175 156.935 112.715 ;
        RECT 152.230 111.705 152.635 111.875 ;
        RECT 152.805 111.705 153.590 111.875 ;
        RECT 153.865 111.425 154.075 111.955 ;
        RECT 154.335 111.640 154.665 112.165 ;
        RECT 155.175 112.080 155.555 112.165 ;
        RECT 154.835 111.425 155.005 112.035 ;
        RECT 155.175 111.645 155.505 112.080 ;
        RECT 155.725 111.425 156.935 112.175 ;
        RECT 22.700 111.255 157.020 111.425 ;
        RECT 22.785 110.505 23.995 111.255 ;
        RECT 22.785 109.965 23.305 110.505 ;
        RECT 24.165 110.485 26.755 111.255 ;
        RECT 23.475 109.795 23.995 110.335 ;
        RECT 24.165 109.965 25.375 110.485 ;
        RECT 25.545 109.795 26.755 110.315 ;
        RECT 22.785 108.705 23.995 109.795 ;
        RECT 24.165 108.705 26.755 109.795 ;
        RECT 26.925 110.310 27.265 111.085 ;
        RECT 27.435 110.795 27.605 111.255 ;
        RECT 27.845 110.820 28.205 111.085 ;
        RECT 27.845 110.815 28.200 110.820 ;
        RECT 27.845 110.805 28.195 110.815 ;
        RECT 27.845 110.800 28.190 110.805 ;
        RECT 27.845 110.790 28.185 110.800 ;
        RECT 28.835 110.795 29.005 111.255 ;
        RECT 27.845 110.785 28.180 110.790 ;
        RECT 27.845 110.775 28.170 110.785 ;
        RECT 27.845 110.765 28.160 110.775 ;
        RECT 27.845 110.625 28.145 110.765 ;
        RECT 27.435 110.435 28.145 110.625 ;
        RECT 28.335 110.625 28.665 110.705 ;
        RECT 29.175 110.625 29.515 111.085 ;
        RECT 28.335 110.435 29.515 110.625 ;
        RECT 29.685 110.485 31.355 111.255 ;
        RECT 31.985 110.605 32.245 111.085 ;
        RECT 32.415 110.795 32.745 111.255 ;
        RECT 32.935 110.615 33.135 111.035 ;
        RECT 26.925 108.875 27.205 110.310 ;
        RECT 27.435 109.865 27.720 110.435 ;
        RECT 27.905 110.035 28.375 110.265 ;
        RECT 28.545 110.245 28.875 110.265 ;
        RECT 28.545 110.065 28.995 110.245 ;
        RECT 29.185 110.065 29.515 110.265 ;
        RECT 27.435 109.650 28.585 109.865 ;
        RECT 27.375 108.705 28.085 109.480 ;
        RECT 28.255 108.875 28.585 109.650 ;
        RECT 28.780 108.950 28.995 110.065 ;
        RECT 29.285 109.725 29.515 110.065 ;
        RECT 29.685 109.965 30.435 110.485 ;
        RECT 30.605 109.795 31.355 110.315 ;
        RECT 29.175 108.705 29.505 109.425 ;
        RECT 29.685 108.705 31.355 109.795 ;
        RECT 31.985 109.575 32.155 110.605 ;
        RECT 32.325 109.915 32.555 110.345 ;
        RECT 32.725 110.095 33.135 110.615 ;
        RECT 33.305 110.770 34.095 111.035 ;
        RECT 33.305 109.915 33.560 110.770 ;
        RECT 34.275 110.435 34.605 110.855 ;
        RECT 34.775 110.435 35.035 111.255 ;
        RECT 35.205 110.710 40.550 111.255 ;
        RECT 40.725 110.710 46.070 111.255 ;
        RECT 34.275 110.345 34.525 110.435 ;
        RECT 33.730 110.095 34.525 110.345 ;
        RECT 32.325 109.745 34.115 109.915 ;
        RECT 31.985 108.875 32.260 109.575 ;
        RECT 32.430 109.450 33.145 109.745 ;
        RECT 33.365 109.385 33.695 109.575 ;
        RECT 32.470 108.705 32.685 109.250 ;
        RECT 32.855 108.875 33.330 109.215 ;
        RECT 33.500 109.210 33.695 109.385 ;
        RECT 33.865 109.380 34.115 109.745 ;
        RECT 33.500 108.705 34.115 109.210 ;
        RECT 34.355 108.875 34.525 110.095 ;
        RECT 34.695 109.385 35.035 110.265 ;
        RECT 36.790 109.880 37.130 110.710 ;
        RECT 34.775 108.705 35.035 109.215 ;
        RECT 38.610 109.140 38.960 110.390 ;
        RECT 42.310 109.880 42.650 110.710 ;
        RECT 46.245 110.485 47.915 111.255 ;
        RECT 48.545 110.530 48.835 111.255 ;
        RECT 49.005 110.485 50.675 111.255 ;
        RECT 50.880 110.515 51.495 111.085 ;
        RECT 51.665 110.745 51.880 111.255 ;
        RECT 52.110 110.745 52.390 111.075 ;
        RECT 52.570 110.745 52.810 111.255 ;
        RECT 53.695 110.915 53.865 110.950 ;
        RECT 53.665 110.745 53.865 110.915 ;
        RECT 44.130 109.140 44.480 110.390 ;
        RECT 46.245 109.965 46.995 110.485 ;
        RECT 47.165 109.795 47.915 110.315 ;
        RECT 49.005 109.965 49.755 110.485 ;
        RECT 35.205 108.705 40.550 109.140 ;
        RECT 40.725 108.705 46.070 109.140 ;
        RECT 46.245 108.705 47.915 109.795 ;
        RECT 48.545 108.705 48.835 109.870 ;
        RECT 49.925 109.795 50.675 110.315 ;
        RECT 49.005 108.705 50.675 109.795 ;
        RECT 50.880 109.495 51.195 110.515 ;
        RECT 51.365 109.845 51.535 110.345 ;
        RECT 51.785 110.015 52.050 110.575 ;
        RECT 52.220 109.845 52.390 110.745 ;
        RECT 52.560 110.015 52.915 110.575 ;
        RECT 53.695 110.385 53.865 110.745 ;
        RECT 54.055 110.725 54.285 111.030 ;
        RECT 54.455 110.895 54.785 111.255 ;
        RECT 54.980 110.725 55.270 111.075 ;
        RECT 54.055 110.555 55.270 110.725 ;
        RECT 55.445 110.515 55.910 111.060 ;
        RECT 53.695 110.215 54.215 110.385 ;
        RECT 51.365 109.675 52.790 109.845 ;
        RECT 53.610 109.685 53.855 110.045 ;
        RECT 54.045 109.835 54.215 110.215 ;
        RECT 54.385 110.015 54.770 110.345 ;
        RECT 54.950 110.235 55.210 110.345 ;
        RECT 54.950 110.065 55.215 110.235 ;
        RECT 54.950 110.015 55.210 110.065 ;
        RECT 50.880 108.875 51.415 109.495 ;
        RECT 51.585 108.705 51.915 109.505 ;
        RECT 52.400 109.500 52.790 109.675 ;
        RECT 54.045 109.555 54.395 109.835 ;
        RECT 53.610 108.705 53.865 109.505 ;
        RECT 54.065 108.875 54.395 109.555 ;
        RECT 54.575 108.965 54.770 110.015 ;
        RECT 54.950 108.705 55.270 109.845 ;
        RECT 55.445 109.555 55.615 110.515 ;
        RECT 56.415 110.435 56.585 111.255 ;
        RECT 56.755 110.605 57.085 111.085 ;
        RECT 57.255 110.865 57.605 111.255 ;
        RECT 57.775 110.685 58.005 111.085 ;
        RECT 57.495 110.605 58.005 110.685 ;
        RECT 56.755 110.515 58.005 110.605 ;
        RECT 58.175 110.515 58.495 110.995 ;
        RECT 58.665 110.710 64.010 111.255 ;
        RECT 65.105 110.875 65.995 111.045 ;
        RECT 56.755 110.435 57.665 110.515 ;
        RECT 55.785 109.895 56.030 110.345 ;
        RECT 56.290 110.065 56.985 110.265 ;
        RECT 57.155 110.095 57.755 110.265 ;
        RECT 57.155 109.895 57.325 110.095 ;
        RECT 57.985 109.925 58.155 110.345 ;
        RECT 55.785 109.725 57.325 109.895 ;
        RECT 57.495 109.755 58.155 109.925 ;
        RECT 57.495 109.555 57.665 109.755 ;
        RECT 58.325 109.585 58.495 110.515 ;
        RECT 60.250 109.880 60.590 110.710 ;
        RECT 55.445 109.385 57.665 109.555 ;
        RECT 57.835 109.385 58.495 109.585 ;
        RECT 55.445 108.705 55.745 109.215 ;
        RECT 55.915 108.875 56.245 109.385 ;
        RECT 57.835 109.215 58.005 109.385 ;
        RECT 56.415 108.705 57.045 109.215 ;
        RECT 57.625 109.045 58.005 109.215 ;
        RECT 58.175 108.705 58.475 109.215 ;
        RECT 62.070 109.140 62.420 110.390 ;
        RECT 65.105 110.320 65.655 110.705 ;
        RECT 65.825 110.150 65.995 110.875 ;
        RECT 65.105 110.080 65.995 110.150 ;
        RECT 66.165 110.550 66.385 111.035 ;
        RECT 66.555 110.715 66.805 111.255 ;
        RECT 66.975 110.605 67.235 111.085 ;
        RECT 66.165 110.125 66.495 110.550 ;
        RECT 65.105 110.055 66.000 110.080 ;
        RECT 65.105 110.040 66.010 110.055 ;
        RECT 65.105 110.025 66.015 110.040 ;
        RECT 65.105 110.020 66.025 110.025 ;
        RECT 65.105 110.010 66.030 110.020 ;
        RECT 65.105 110.000 66.035 110.010 ;
        RECT 65.105 109.995 66.045 110.000 ;
        RECT 65.105 109.985 66.055 109.995 ;
        RECT 65.105 109.980 66.065 109.985 ;
        RECT 65.105 109.530 65.365 109.980 ;
        RECT 65.730 109.975 66.065 109.980 ;
        RECT 65.730 109.970 66.080 109.975 ;
        RECT 65.730 109.960 66.095 109.970 ;
        RECT 65.730 109.955 66.120 109.960 ;
        RECT 66.665 109.955 66.895 110.350 ;
        RECT 65.730 109.950 66.895 109.955 ;
        RECT 65.760 109.915 66.895 109.950 ;
        RECT 65.795 109.890 66.895 109.915 ;
        RECT 65.825 109.860 66.895 109.890 ;
        RECT 65.845 109.830 66.895 109.860 ;
        RECT 65.865 109.800 66.895 109.830 ;
        RECT 65.935 109.790 66.895 109.800 ;
        RECT 65.960 109.780 66.895 109.790 ;
        RECT 65.980 109.765 66.895 109.780 ;
        RECT 66.000 109.750 66.895 109.765 ;
        RECT 66.005 109.740 66.790 109.750 ;
        RECT 66.020 109.705 66.790 109.740 ;
        RECT 65.535 109.385 65.865 109.630 ;
        RECT 66.035 109.455 66.790 109.705 ;
        RECT 67.065 109.575 67.235 110.605 ;
        RECT 67.415 110.445 67.685 111.255 ;
        RECT 67.855 110.445 68.185 111.085 ;
        RECT 68.355 110.445 68.595 111.255 ;
        RECT 69.725 110.525 70.015 111.255 ;
        RECT 67.405 110.015 67.755 110.265 ;
        RECT 67.925 109.845 68.095 110.445 ;
        RECT 68.265 110.015 68.615 110.265 ;
        RECT 69.715 110.015 70.015 110.345 ;
        RECT 70.195 110.325 70.425 110.965 ;
        RECT 70.605 110.705 70.915 111.075 ;
        RECT 71.095 110.885 71.765 111.255 ;
        RECT 70.605 110.505 71.835 110.705 ;
        RECT 70.195 110.015 70.720 110.325 ;
        RECT 70.900 110.015 71.365 110.325 ;
        RECT 65.535 109.360 65.720 109.385 ;
        RECT 65.105 109.260 65.720 109.360 ;
        RECT 58.665 108.705 64.010 109.140 ;
        RECT 65.105 108.705 65.710 109.260 ;
        RECT 65.885 108.875 66.365 109.215 ;
        RECT 66.535 108.705 66.790 109.250 ;
        RECT 66.960 108.875 67.235 109.575 ;
        RECT 67.415 108.705 67.745 109.845 ;
        RECT 67.925 109.675 68.605 109.845 ;
        RECT 71.545 109.835 71.835 110.505 ;
        RECT 68.275 108.890 68.605 109.675 ;
        RECT 69.725 109.595 70.885 109.835 ;
        RECT 69.725 108.885 69.985 109.595 ;
        RECT 70.155 108.705 70.485 109.415 ;
        RECT 70.655 108.885 70.885 109.595 ;
        RECT 71.065 109.615 71.835 109.835 ;
        RECT 71.065 108.885 71.335 109.615 ;
        RECT 71.515 108.705 71.855 109.435 ;
        RECT 72.025 108.885 72.285 111.075 ;
        RECT 72.465 110.485 74.135 111.255 ;
        RECT 74.305 110.530 74.595 111.255 ;
        RECT 75.315 110.705 75.485 110.995 ;
        RECT 75.655 110.875 75.985 111.255 ;
        RECT 75.315 110.535 75.980 110.705 ;
        RECT 72.465 109.965 73.215 110.485 ;
        RECT 73.385 109.795 74.135 110.315 ;
        RECT 72.465 108.705 74.135 109.795 ;
        RECT 74.305 108.705 74.595 109.870 ;
        RECT 75.230 109.715 75.580 110.365 ;
        RECT 75.750 109.545 75.980 110.535 ;
        RECT 75.315 109.375 75.980 109.545 ;
        RECT 75.315 108.875 75.485 109.375 ;
        RECT 75.655 108.705 75.985 109.205 ;
        RECT 76.155 108.875 76.340 110.995 ;
        RECT 76.595 110.795 76.845 111.255 ;
        RECT 77.015 110.805 77.350 110.975 ;
        RECT 77.545 110.805 78.220 110.975 ;
        RECT 77.015 110.665 77.185 110.805 ;
        RECT 76.510 109.675 76.790 110.625 ;
        RECT 76.960 110.535 77.185 110.665 ;
        RECT 76.960 109.430 77.130 110.535 ;
        RECT 77.355 110.385 77.880 110.605 ;
        RECT 77.300 109.620 77.540 110.215 ;
        RECT 77.710 109.685 77.880 110.385 ;
        RECT 78.050 110.025 78.220 110.805 ;
        RECT 78.540 110.755 78.910 111.255 ;
        RECT 79.090 110.805 79.495 110.975 ;
        RECT 79.665 110.805 80.450 110.975 ;
        RECT 79.090 110.575 79.260 110.805 ;
        RECT 78.430 110.275 79.260 110.575 ;
        RECT 79.645 110.305 80.110 110.635 ;
        RECT 78.430 110.245 78.630 110.275 ;
        RECT 78.750 110.025 78.920 110.095 ;
        RECT 78.050 109.855 78.920 110.025 ;
        RECT 78.410 109.765 78.920 109.855 ;
        RECT 76.960 109.300 77.265 109.430 ;
        RECT 77.710 109.320 78.240 109.685 ;
        RECT 76.580 108.705 76.845 109.165 ;
        RECT 77.015 108.875 77.265 109.300 ;
        RECT 78.410 109.150 78.580 109.765 ;
        RECT 77.475 108.980 78.580 109.150 ;
        RECT 78.750 108.705 78.920 109.505 ;
        RECT 79.090 109.205 79.260 110.275 ;
        RECT 79.430 109.375 79.620 110.095 ;
        RECT 79.790 109.345 80.110 110.305 ;
        RECT 80.280 110.345 80.450 110.805 ;
        RECT 80.725 110.725 80.935 111.255 ;
        RECT 81.195 110.515 81.525 111.040 ;
        RECT 81.695 110.645 81.865 111.255 ;
        RECT 82.035 110.600 82.365 111.035 ;
        RECT 82.035 110.515 82.415 110.600 ;
        RECT 81.325 110.345 81.525 110.515 ;
        RECT 82.190 110.475 82.415 110.515 ;
        RECT 80.280 110.015 81.155 110.345 ;
        RECT 81.325 110.015 82.075 110.345 ;
        RECT 79.090 108.875 79.340 109.205 ;
        RECT 80.280 109.175 80.450 110.015 ;
        RECT 81.325 109.810 81.515 110.015 ;
        RECT 82.245 109.895 82.415 110.475 ;
        RECT 82.585 110.485 85.175 111.255 ;
        RECT 85.895 110.705 86.065 110.995 ;
        RECT 86.235 110.875 86.565 111.255 ;
        RECT 85.895 110.535 86.560 110.705 ;
        RECT 82.585 109.965 83.795 110.485 ;
        RECT 82.200 109.845 82.415 109.895 ;
        RECT 80.620 109.435 81.515 109.810 ;
        RECT 82.025 109.765 82.415 109.845 ;
        RECT 83.965 109.795 85.175 110.315 ;
        RECT 79.565 109.005 80.450 109.175 ;
        RECT 80.630 108.705 80.945 109.205 ;
        RECT 81.175 108.875 81.515 109.435 ;
        RECT 81.685 108.705 81.855 109.715 ;
        RECT 82.025 108.920 82.355 109.765 ;
        RECT 82.585 108.705 85.175 109.795 ;
        RECT 85.810 109.715 86.160 110.365 ;
        RECT 86.330 109.545 86.560 110.535 ;
        RECT 85.895 109.375 86.560 109.545 ;
        RECT 85.895 108.875 86.065 109.375 ;
        RECT 86.235 108.705 86.565 109.205 ;
        RECT 86.735 108.875 86.920 110.995 ;
        RECT 87.175 110.795 87.425 111.255 ;
        RECT 87.595 110.805 87.930 110.975 ;
        RECT 88.125 110.805 88.800 110.975 ;
        RECT 87.595 110.665 87.765 110.805 ;
        RECT 87.090 109.675 87.370 110.625 ;
        RECT 87.540 110.535 87.765 110.665 ;
        RECT 87.540 109.430 87.710 110.535 ;
        RECT 87.935 110.385 88.460 110.605 ;
        RECT 87.880 109.620 88.120 110.215 ;
        RECT 88.290 109.685 88.460 110.385 ;
        RECT 88.630 110.025 88.800 110.805 ;
        RECT 89.120 110.755 89.490 111.255 ;
        RECT 89.670 110.805 90.075 110.975 ;
        RECT 90.245 110.805 91.030 110.975 ;
        RECT 89.670 110.575 89.840 110.805 ;
        RECT 89.010 110.275 89.840 110.575 ;
        RECT 90.225 110.305 90.690 110.635 ;
        RECT 89.010 110.245 89.210 110.275 ;
        RECT 89.330 110.025 89.500 110.095 ;
        RECT 88.630 109.855 89.500 110.025 ;
        RECT 88.990 109.765 89.500 109.855 ;
        RECT 87.540 109.300 87.845 109.430 ;
        RECT 88.290 109.320 88.820 109.685 ;
        RECT 87.160 108.705 87.425 109.165 ;
        RECT 87.595 108.875 87.845 109.300 ;
        RECT 88.990 109.150 89.160 109.765 ;
        RECT 88.055 108.980 89.160 109.150 ;
        RECT 89.330 108.705 89.500 109.505 ;
        RECT 89.670 109.205 89.840 110.275 ;
        RECT 90.010 109.375 90.200 110.095 ;
        RECT 90.370 109.345 90.690 110.305 ;
        RECT 90.860 110.345 91.030 110.805 ;
        RECT 91.305 110.725 91.515 111.255 ;
        RECT 91.775 110.515 92.105 111.040 ;
        RECT 92.275 110.645 92.445 111.255 ;
        RECT 92.615 110.600 92.945 111.035 ;
        RECT 92.615 110.515 92.995 110.600 ;
        RECT 91.905 110.345 92.105 110.515 ;
        RECT 92.770 110.475 92.995 110.515 ;
        RECT 90.860 110.015 91.735 110.345 ;
        RECT 91.905 110.015 92.655 110.345 ;
        RECT 89.670 108.875 89.920 109.205 ;
        RECT 90.860 109.175 91.030 110.015 ;
        RECT 91.905 109.810 92.095 110.015 ;
        RECT 92.825 109.895 92.995 110.475 ;
        RECT 92.780 109.845 92.995 109.895 ;
        RECT 91.200 109.435 92.095 109.810 ;
        RECT 92.605 109.765 92.995 109.845 ;
        RECT 93.165 110.515 93.550 111.085 ;
        RECT 93.720 110.795 94.045 111.255 ;
        RECT 94.565 110.625 94.845 111.085 ;
        RECT 93.165 109.845 93.445 110.515 ;
        RECT 93.720 110.455 94.845 110.625 ;
        RECT 93.720 110.345 94.170 110.455 ;
        RECT 93.615 110.015 94.170 110.345 ;
        RECT 95.035 110.285 95.435 111.085 ;
        RECT 95.835 110.795 96.105 111.255 ;
        RECT 96.275 110.625 96.560 111.085 ;
        RECT 90.145 109.005 91.030 109.175 ;
        RECT 91.210 108.705 91.525 109.205 ;
        RECT 91.755 108.875 92.095 109.435 ;
        RECT 92.265 108.705 92.435 109.715 ;
        RECT 92.605 108.920 92.935 109.765 ;
        RECT 93.165 108.875 93.550 109.845 ;
        RECT 93.720 109.555 94.170 110.015 ;
        RECT 94.340 109.725 95.435 110.285 ;
        RECT 93.720 109.335 94.845 109.555 ;
        RECT 93.720 108.705 94.045 109.165 ;
        RECT 94.565 108.875 94.845 109.335 ;
        RECT 95.035 108.875 95.435 109.725 ;
        RECT 95.605 110.455 96.560 110.625 ;
        RECT 95.605 109.555 95.815 110.455 ;
        RECT 95.985 109.725 96.675 110.285 ;
        RECT 95.605 109.335 96.560 109.555 ;
        RECT 95.835 108.705 96.105 109.165 ;
        RECT 96.275 108.875 96.560 109.335 ;
        RECT 96.855 108.885 97.115 111.075 ;
        RECT 97.375 110.885 98.045 111.255 ;
        RECT 98.225 110.705 98.535 111.075 ;
        RECT 97.305 110.505 98.535 110.705 ;
        RECT 97.305 109.835 97.595 110.505 ;
        RECT 98.715 110.325 98.945 110.965 ;
        RECT 99.125 110.525 99.415 111.255 ;
        RECT 100.065 110.530 100.355 111.255 ;
        RECT 100.545 110.445 100.785 111.255 ;
        RECT 100.955 110.445 101.285 111.085 ;
        RECT 101.455 110.445 101.725 111.255 ;
        RECT 101.905 110.485 104.495 111.255 ;
        RECT 97.775 110.015 98.240 110.325 ;
        RECT 98.420 110.015 98.945 110.325 ;
        RECT 99.125 110.015 99.425 110.345 ;
        RECT 100.525 110.015 100.875 110.265 ;
        RECT 97.305 109.615 98.075 109.835 ;
        RECT 97.285 108.705 97.625 109.435 ;
        RECT 97.805 108.885 98.075 109.615 ;
        RECT 98.255 109.595 99.415 109.835 ;
        RECT 98.255 108.885 98.485 109.595 ;
        RECT 98.655 108.705 98.985 109.415 ;
        RECT 99.155 108.885 99.415 109.595 ;
        RECT 100.065 108.705 100.355 109.870 ;
        RECT 101.045 109.845 101.215 110.445 ;
        RECT 101.385 110.015 101.735 110.265 ;
        RECT 101.905 109.965 103.115 110.485 ;
        RECT 100.535 109.675 101.215 109.845 ;
        RECT 100.535 108.890 100.865 109.675 ;
        RECT 101.395 108.705 101.725 109.845 ;
        RECT 103.285 109.795 104.495 110.315 ;
        RECT 101.905 108.705 104.495 109.795 ;
        RECT 104.675 108.885 104.935 111.075 ;
        RECT 105.195 110.885 105.865 111.255 ;
        RECT 106.045 110.705 106.355 111.075 ;
        RECT 105.125 110.505 106.355 110.705 ;
        RECT 105.125 109.835 105.415 110.505 ;
        RECT 106.535 110.325 106.765 110.965 ;
        RECT 106.945 110.525 107.235 111.255 ;
        RECT 107.485 110.435 107.695 111.255 ;
        RECT 107.865 110.455 108.195 111.085 ;
        RECT 105.595 110.015 106.060 110.325 ;
        RECT 106.240 110.015 106.765 110.325 ;
        RECT 106.945 110.015 107.245 110.345 ;
        RECT 107.865 109.855 108.115 110.455 ;
        RECT 108.365 110.435 108.595 111.255 ;
        RECT 108.805 110.710 114.150 111.255 ;
        RECT 108.285 110.015 108.615 110.265 ;
        RECT 110.390 109.880 110.730 110.710 ;
        RECT 114.425 110.410 114.595 111.255 ;
        RECT 114.765 110.530 115.020 111.085 ;
        RECT 115.190 110.810 115.620 111.255 ;
        RECT 115.855 110.685 116.025 111.085 ;
        RECT 116.195 110.855 116.930 111.255 ;
        RECT 105.125 109.615 105.895 109.835 ;
        RECT 105.105 108.705 105.445 109.435 ;
        RECT 105.625 108.885 105.895 109.615 ;
        RECT 106.075 109.595 107.235 109.835 ;
        RECT 106.075 108.885 106.305 109.595 ;
        RECT 106.475 108.705 106.805 109.415 ;
        RECT 106.975 108.885 107.235 109.595 ;
        RECT 107.485 108.705 107.695 109.845 ;
        RECT 107.865 108.875 108.195 109.855 ;
        RECT 108.365 108.705 108.595 109.845 ;
        RECT 112.210 109.140 112.560 110.390 ;
        RECT 108.805 108.705 114.150 109.140 ;
        RECT 114.425 108.705 114.595 109.895 ;
        RECT 114.765 109.815 114.935 110.530 ;
        RECT 115.855 110.515 116.750 110.685 ;
        RECT 117.100 110.640 117.270 111.085 ;
        RECT 117.845 110.745 118.245 111.255 ;
        RECT 115.105 110.015 115.360 110.345 ;
        RECT 114.765 108.875 115.020 109.815 ;
        RECT 115.190 109.535 115.360 110.015 ;
        RECT 115.585 109.725 115.915 110.345 ;
        RECT 116.085 110.235 116.375 110.345 ;
        RECT 116.085 110.065 116.395 110.235 ;
        RECT 116.085 109.965 116.375 110.065 ;
        RECT 116.580 109.795 116.750 110.515 ;
        RECT 116.215 109.625 116.750 109.795 ;
        RECT 116.920 110.470 117.270 110.640 ;
        RECT 118.515 110.600 118.845 111.035 ;
        RECT 119.015 110.645 119.185 111.255 ;
        RECT 115.190 109.365 115.950 109.535 ;
        RECT 116.215 109.435 116.385 109.625 ;
        RECT 116.920 109.445 117.090 110.470 ;
        RECT 117.510 109.985 117.770 110.575 ;
        RECT 117.290 109.895 117.770 109.985 ;
        RECT 117.970 110.405 118.235 110.575 ;
        RECT 118.465 110.515 118.845 110.600 ;
        RECT 119.355 110.515 119.685 111.040 ;
        RECT 119.945 110.725 120.155 111.255 ;
        RECT 120.430 110.805 121.215 110.975 ;
        RECT 121.385 110.805 121.790 110.975 ;
        RECT 118.465 110.475 118.690 110.515 ;
        RECT 117.290 109.725 117.775 109.895 ;
        RECT 117.290 109.685 117.770 109.725 ;
        RECT 117.970 109.685 118.230 110.405 ;
        RECT 118.465 109.895 118.635 110.475 ;
        RECT 119.355 110.345 119.555 110.515 ;
        RECT 120.430 110.345 120.600 110.805 ;
        RECT 118.805 110.015 119.555 110.345 ;
        RECT 119.725 110.015 120.600 110.345 ;
        RECT 118.465 109.845 118.680 109.895 ;
        RECT 118.465 109.765 118.855 109.845 ;
        RECT 115.780 109.140 115.950 109.365 ;
        RECT 116.680 109.275 117.090 109.445 ;
        RECT 117.275 109.335 118.205 109.505 ;
        RECT 116.680 109.140 116.910 109.275 ;
        RECT 115.190 108.705 115.520 109.105 ;
        RECT 115.780 108.970 116.910 109.140 ;
        RECT 117.275 109.085 117.445 109.335 ;
        RECT 116.740 108.875 116.910 108.970 ;
        RECT 117.115 108.915 117.445 109.085 ;
        RECT 117.615 108.705 117.865 109.165 ;
        RECT 118.035 108.875 118.205 109.335 ;
        RECT 118.525 108.920 118.855 109.765 ;
        RECT 119.365 109.810 119.555 110.015 ;
        RECT 119.025 108.705 119.195 109.715 ;
        RECT 119.365 109.435 120.260 109.810 ;
        RECT 119.365 108.875 119.705 109.435 ;
        RECT 119.935 108.705 120.250 109.205 ;
        RECT 120.430 109.175 120.600 110.015 ;
        RECT 120.770 110.305 121.235 110.635 ;
        RECT 121.620 110.575 121.790 110.805 ;
        RECT 121.970 110.755 122.340 111.255 ;
        RECT 122.660 110.805 123.335 110.975 ;
        RECT 123.530 110.805 123.865 110.975 ;
        RECT 120.770 109.345 121.090 110.305 ;
        RECT 121.620 110.275 122.450 110.575 ;
        RECT 121.260 109.375 121.450 110.095 ;
        RECT 121.620 109.205 121.790 110.275 ;
        RECT 122.250 110.245 122.450 110.275 ;
        RECT 121.960 110.025 122.130 110.095 ;
        RECT 122.660 110.025 122.830 110.805 ;
        RECT 123.695 110.665 123.865 110.805 ;
        RECT 124.035 110.795 124.285 111.255 ;
        RECT 121.960 109.855 122.830 110.025 ;
        RECT 123.000 110.385 123.525 110.605 ;
        RECT 123.695 110.535 123.920 110.665 ;
        RECT 121.960 109.765 122.470 109.855 ;
        RECT 120.430 109.005 121.315 109.175 ;
        RECT 121.540 108.875 121.790 109.205 ;
        RECT 121.960 108.705 122.130 109.505 ;
        RECT 122.300 109.150 122.470 109.765 ;
        RECT 123.000 109.685 123.170 110.385 ;
        RECT 122.640 109.320 123.170 109.685 ;
        RECT 123.340 109.620 123.580 110.215 ;
        RECT 123.750 109.430 123.920 110.535 ;
        RECT 124.090 109.675 124.370 110.625 ;
        RECT 123.615 109.300 123.920 109.430 ;
        RECT 122.300 108.980 123.405 109.150 ;
        RECT 123.615 108.875 123.865 109.300 ;
        RECT 124.035 108.705 124.300 109.165 ;
        RECT 124.540 108.875 124.725 110.995 ;
        RECT 124.895 110.875 125.225 111.255 ;
        RECT 125.395 110.705 125.565 110.995 ;
        RECT 124.900 110.535 125.565 110.705 ;
        RECT 124.900 109.545 125.130 110.535 ;
        RECT 125.825 110.530 126.115 111.255 ;
        RECT 126.285 110.485 128.875 111.255 ;
        RECT 129.160 110.625 129.445 111.085 ;
        RECT 129.615 110.795 129.885 111.255 ;
        RECT 125.300 109.715 125.650 110.365 ;
        RECT 126.285 109.965 127.495 110.485 ;
        RECT 129.160 110.455 130.115 110.625 ;
        RECT 124.900 109.375 125.565 109.545 ;
        RECT 124.895 108.705 125.225 109.205 ;
        RECT 125.395 108.875 125.565 109.375 ;
        RECT 125.825 108.705 126.115 109.870 ;
        RECT 127.665 109.795 128.875 110.315 ;
        RECT 126.285 108.705 128.875 109.795 ;
        RECT 129.045 109.725 129.735 110.285 ;
        RECT 129.905 109.555 130.115 110.455 ;
        RECT 129.160 109.335 130.115 109.555 ;
        RECT 130.285 110.285 130.685 111.085 ;
        RECT 130.875 110.625 131.155 111.085 ;
        RECT 131.675 110.795 132.000 111.255 ;
        RECT 130.875 110.455 132.000 110.625 ;
        RECT 132.170 110.515 132.555 111.085 ;
        RECT 132.815 110.705 132.985 110.995 ;
        RECT 133.155 110.875 133.485 111.255 ;
        RECT 132.815 110.535 133.480 110.705 ;
        RECT 131.550 110.345 132.000 110.455 ;
        RECT 130.285 109.725 131.380 110.285 ;
        RECT 131.550 110.015 132.105 110.345 ;
        RECT 129.160 108.875 129.445 109.335 ;
        RECT 129.615 108.705 129.885 109.165 ;
        RECT 130.285 108.875 130.685 109.725 ;
        RECT 131.550 109.555 132.000 110.015 ;
        RECT 132.275 109.845 132.555 110.515 ;
        RECT 130.875 109.335 132.000 109.555 ;
        RECT 130.875 108.875 131.155 109.335 ;
        RECT 131.675 108.705 132.000 109.165 ;
        RECT 132.170 108.875 132.555 109.845 ;
        RECT 132.730 109.715 133.080 110.365 ;
        RECT 133.250 109.545 133.480 110.535 ;
        RECT 132.815 109.375 133.480 109.545 ;
        RECT 132.815 108.875 132.985 109.375 ;
        RECT 133.155 108.705 133.485 109.205 ;
        RECT 133.655 108.875 133.840 110.995 ;
        RECT 134.095 110.795 134.345 111.255 ;
        RECT 134.515 110.805 134.850 110.975 ;
        RECT 135.045 110.805 135.720 110.975 ;
        RECT 134.515 110.665 134.685 110.805 ;
        RECT 134.010 109.675 134.290 110.625 ;
        RECT 134.460 110.535 134.685 110.665 ;
        RECT 134.460 109.430 134.630 110.535 ;
        RECT 134.855 110.385 135.380 110.605 ;
        RECT 134.800 109.620 135.040 110.215 ;
        RECT 135.210 109.685 135.380 110.385 ;
        RECT 135.550 110.025 135.720 110.805 ;
        RECT 136.040 110.755 136.410 111.255 ;
        RECT 136.590 110.805 136.995 110.975 ;
        RECT 137.165 110.805 137.950 110.975 ;
        RECT 136.590 110.575 136.760 110.805 ;
        RECT 135.930 110.275 136.760 110.575 ;
        RECT 137.145 110.305 137.610 110.635 ;
        RECT 135.930 110.245 136.130 110.275 ;
        RECT 136.250 110.025 136.420 110.095 ;
        RECT 135.550 109.855 136.420 110.025 ;
        RECT 135.910 109.765 136.420 109.855 ;
        RECT 134.460 109.300 134.765 109.430 ;
        RECT 135.210 109.320 135.740 109.685 ;
        RECT 134.080 108.705 134.345 109.165 ;
        RECT 134.515 108.875 134.765 109.300 ;
        RECT 135.910 109.150 136.080 109.765 ;
        RECT 134.975 108.980 136.080 109.150 ;
        RECT 136.250 108.705 136.420 109.505 ;
        RECT 136.590 109.205 136.760 110.275 ;
        RECT 136.930 109.375 137.120 110.095 ;
        RECT 137.290 109.345 137.610 110.305 ;
        RECT 137.780 110.345 137.950 110.805 ;
        RECT 138.225 110.725 138.435 111.255 ;
        RECT 138.695 110.515 139.025 111.040 ;
        RECT 139.195 110.645 139.365 111.255 ;
        RECT 139.535 110.600 139.865 111.035 ;
        RECT 140.135 110.600 140.465 111.035 ;
        RECT 140.635 110.645 140.805 111.255 ;
        RECT 139.535 110.515 139.915 110.600 ;
        RECT 138.825 110.345 139.025 110.515 ;
        RECT 139.690 110.475 139.915 110.515 ;
        RECT 137.780 110.015 138.655 110.345 ;
        RECT 138.825 110.015 139.575 110.345 ;
        RECT 136.590 108.875 136.840 109.205 ;
        RECT 137.780 109.175 137.950 110.015 ;
        RECT 138.825 109.810 139.015 110.015 ;
        RECT 139.745 109.895 139.915 110.475 ;
        RECT 139.700 109.845 139.915 109.895 ;
        RECT 138.120 109.435 139.015 109.810 ;
        RECT 139.525 109.765 139.915 109.845 ;
        RECT 140.085 110.515 140.465 110.600 ;
        RECT 140.975 110.515 141.305 111.040 ;
        RECT 141.565 110.725 141.775 111.255 ;
        RECT 142.050 110.805 142.835 110.975 ;
        RECT 143.005 110.805 143.410 110.975 ;
        RECT 140.085 110.475 140.310 110.515 ;
        RECT 140.085 109.895 140.255 110.475 ;
        RECT 140.975 110.345 141.175 110.515 ;
        RECT 142.050 110.345 142.220 110.805 ;
        RECT 140.425 110.015 141.175 110.345 ;
        RECT 141.345 110.015 142.220 110.345 ;
        RECT 140.085 109.845 140.300 109.895 ;
        RECT 140.085 109.765 140.475 109.845 ;
        RECT 137.065 109.005 137.950 109.175 ;
        RECT 138.130 108.705 138.445 109.205 ;
        RECT 138.675 108.875 139.015 109.435 ;
        RECT 139.185 108.705 139.355 109.715 ;
        RECT 139.525 108.920 139.855 109.765 ;
        RECT 140.145 108.920 140.475 109.765 ;
        RECT 140.985 109.810 141.175 110.015 ;
        RECT 140.645 108.705 140.815 109.715 ;
        RECT 140.985 109.435 141.880 109.810 ;
        RECT 140.985 108.875 141.325 109.435 ;
        RECT 141.555 108.705 141.870 109.205 ;
        RECT 142.050 109.175 142.220 110.015 ;
        RECT 142.390 110.305 142.855 110.635 ;
        RECT 143.240 110.575 143.410 110.805 ;
        RECT 143.590 110.755 143.960 111.255 ;
        RECT 144.280 110.805 144.955 110.975 ;
        RECT 145.150 110.805 145.485 110.975 ;
        RECT 142.390 109.345 142.710 110.305 ;
        RECT 143.240 110.275 144.070 110.575 ;
        RECT 142.880 109.375 143.070 110.095 ;
        RECT 143.240 109.205 143.410 110.275 ;
        RECT 143.870 110.245 144.070 110.275 ;
        RECT 143.580 110.025 143.750 110.095 ;
        RECT 144.280 110.025 144.450 110.805 ;
        RECT 145.315 110.665 145.485 110.805 ;
        RECT 145.655 110.795 145.905 111.255 ;
        RECT 143.580 109.855 144.450 110.025 ;
        RECT 144.620 110.385 145.145 110.605 ;
        RECT 145.315 110.535 145.540 110.665 ;
        RECT 143.580 109.765 144.090 109.855 ;
        RECT 142.050 109.005 142.935 109.175 ;
        RECT 143.160 108.875 143.410 109.205 ;
        RECT 143.580 108.705 143.750 109.505 ;
        RECT 143.920 109.150 144.090 109.765 ;
        RECT 144.620 109.685 144.790 110.385 ;
        RECT 144.260 109.320 144.790 109.685 ;
        RECT 144.960 109.620 145.200 110.215 ;
        RECT 145.370 109.430 145.540 110.535 ;
        RECT 145.710 109.675 145.990 110.625 ;
        RECT 145.235 109.300 145.540 109.430 ;
        RECT 143.920 108.980 145.025 109.150 ;
        RECT 145.235 108.875 145.485 109.300 ;
        RECT 145.655 108.705 145.920 109.165 ;
        RECT 146.160 108.875 146.345 110.995 ;
        RECT 146.515 110.875 146.845 111.255 ;
        RECT 147.015 110.705 147.185 110.995 ;
        RECT 146.520 110.535 147.185 110.705 ;
        RECT 146.520 109.545 146.750 110.535 ;
        RECT 147.445 110.515 147.830 111.085 ;
        RECT 148.000 110.795 148.325 111.255 ;
        RECT 148.845 110.625 149.125 111.085 ;
        RECT 146.920 109.715 147.270 110.365 ;
        RECT 147.445 109.845 147.725 110.515 ;
        RECT 148.000 110.455 149.125 110.625 ;
        RECT 148.000 110.345 148.450 110.455 ;
        RECT 147.895 110.015 148.450 110.345 ;
        RECT 149.315 110.285 149.715 111.085 ;
        RECT 150.115 110.795 150.385 111.255 ;
        RECT 150.555 110.625 150.840 111.085 ;
        RECT 146.520 109.375 147.185 109.545 ;
        RECT 146.515 108.705 146.845 109.205 ;
        RECT 147.015 108.875 147.185 109.375 ;
        RECT 147.445 108.875 147.830 109.845 ;
        RECT 148.000 109.555 148.450 110.015 ;
        RECT 148.620 109.725 149.715 110.285 ;
        RECT 148.000 109.335 149.125 109.555 ;
        RECT 148.000 108.705 148.325 109.165 ;
        RECT 148.845 108.875 149.125 109.335 ;
        RECT 149.315 108.875 149.715 109.725 ;
        RECT 149.885 110.455 150.840 110.625 ;
        RECT 151.585 110.530 151.875 111.255 ;
        RECT 152.045 110.515 152.430 111.085 ;
        RECT 152.600 110.795 152.925 111.255 ;
        RECT 153.445 110.625 153.725 111.085 ;
        RECT 149.885 109.555 150.095 110.455 ;
        RECT 150.265 109.725 150.955 110.285 ;
        RECT 149.885 109.335 150.840 109.555 ;
        RECT 150.115 108.705 150.385 109.165 ;
        RECT 150.555 108.875 150.840 109.335 ;
        RECT 151.585 108.705 151.875 109.870 ;
        RECT 152.045 109.845 152.325 110.515 ;
        RECT 152.600 110.455 153.725 110.625 ;
        RECT 152.600 110.345 153.050 110.455 ;
        RECT 152.495 110.015 153.050 110.345 ;
        RECT 153.915 110.285 154.315 111.085 ;
        RECT 154.715 110.795 154.985 111.255 ;
        RECT 155.155 110.625 155.440 111.085 ;
        RECT 152.045 108.875 152.430 109.845 ;
        RECT 152.600 109.555 153.050 110.015 ;
        RECT 153.220 109.725 154.315 110.285 ;
        RECT 152.600 109.335 153.725 109.555 ;
        RECT 152.600 108.705 152.925 109.165 ;
        RECT 153.445 108.875 153.725 109.335 ;
        RECT 153.915 108.875 154.315 109.725 ;
        RECT 154.485 110.455 155.440 110.625 ;
        RECT 155.725 110.505 156.935 111.255 ;
        RECT 154.485 109.555 154.695 110.455 ;
        RECT 154.865 109.725 155.555 110.285 ;
        RECT 155.725 109.795 156.245 110.335 ;
        RECT 156.415 109.965 156.935 110.505 ;
        RECT 154.485 109.335 155.440 109.555 ;
        RECT 154.715 108.705 154.985 109.165 ;
        RECT 155.155 108.875 155.440 109.335 ;
        RECT 155.725 108.705 156.935 109.795 ;
        RECT 22.700 108.535 157.020 108.705 ;
        RECT 22.785 107.445 23.995 108.535 ;
        RECT 24.165 108.100 29.510 108.535 ;
        RECT 22.785 106.735 23.305 107.275 ;
        RECT 23.475 106.905 23.995 107.445 ;
        RECT 22.785 105.985 23.995 106.735 ;
        RECT 25.750 106.530 26.090 107.360 ;
        RECT 27.570 106.850 27.920 108.100 ;
        RECT 29.685 107.445 32.275 108.535 ;
        RECT 29.685 106.755 30.895 107.275 ;
        RECT 31.065 106.925 32.275 107.445 ;
        RECT 32.465 107.645 32.725 108.355 ;
        RECT 32.895 107.825 33.225 108.535 ;
        RECT 33.395 107.645 33.625 108.355 ;
        RECT 32.465 107.405 33.625 107.645 ;
        RECT 33.805 107.625 34.075 108.355 ;
        RECT 34.255 107.805 34.595 108.535 ;
        RECT 33.805 107.405 34.575 107.625 ;
        RECT 32.455 106.895 32.755 107.225 ;
        RECT 32.935 106.915 33.460 107.225 ;
        RECT 33.640 106.915 34.105 107.225 ;
        RECT 24.165 105.985 29.510 106.530 ;
        RECT 29.685 105.985 32.275 106.755 ;
        RECT 32.465 105.985 32.755 106.715 ;
        RECT 32.935 106.275 33.165 106.915 ;
        RECT 34.285 106.735 34.575 107.405 ;
        RECT 33.345 106.535 34.575 106.735 ;
        RECT 33.345 106.165 33.655 106.535 ;
        RECT 33.835 105.985 34.505 106.355 ;
        RECT 34.765 106.165 35.025 108.355 ;
        RECT 35.665 107.370 35.955 108.535 ;
        RECT 36.135 107.925 36.465 108.355 ;
        RECT 36.645 108.095 36.840 108.535 ;
        RECT 37.010 107.925 37.340 108.355 ;
        RECT 36.135 107.755 37.340 107.925 ;
        RECT 36.135 107.425 37.030 107.755 ;
        RECT 37.510 107.585 37.785 108.355 ;
        RECT 37.200 107.395 37.785 107.585 ;
        RECT 37.965 107.445 39.635 108.535 ;
        RECT 36.140 106.895 36.435 107.225 ;
        RECT 36.615 106.895 37.030 107.225 ;
        RECT 35.665 105.985 35.955 106.710 ;
        RECT 36.135 105.985 36.435 106.715 ;
        RECT 36.615 106.275 36.845 106.895 ;
        RECT 37.200 106.725 37.375 107.395 ;
        RECT 37.045 106.545 37.375 106.725 ;
        RECT 37.545 106.575 37.785 107.225 ;
        RECT 37.965 106.755 38.715 107.275 ;
        RECT 38.885 106.925 39.635 107.445 ;
        RECT 39.805 107.395 40.065 108.535 ;
        RECT 40.235 107.385 40.565 108.365 ;
        RECT 40.735 107.395 41.015 108.535 ;
        RECT 41.185 107.395 41.570 108.365 ;
        RECT 41.740 108.075 42.065 108.535 ;
        RECT 42.585 107.905 42.865 108.365 ;
        RECT 41.740 107.685 42.865 107.905 ;
        RECT 39.825 106.975 40.160 107.225 ;
        RECT 40.330 106.785 40.500 107.385 ;
        RECT 40.670 106.955 41.005 107.225 ;
        RECT 37.045 106.165 37.270 106.545 ;
        RECT 37.440 105.985 37.770 106.375 ;
        RECT 37.965 105.985 39.635 106.755 ;
        RECT 39.805 106.155 40.500 106.785 ;
        RECT 40.705 105.985 41.015 106.785 ;
        RECT 41.185 106.725 41.465 107.395 ;
        RECT 41.740 107.225 42.190 107.685 ;
        RECT 43.055 107.515 43.455 108.365 ;
        RECT 43.855 108.075 44.125 108.535 ;
        RECT 44.295 107.905 44.580 108.365 ;
        RECT 41.635 106.895 42.190 107.225 ;
        RECT 42.360 106.955 43.455 107.515 ;
        RECT 41.740 106.785 42.190 106.895 ;
        RECT 41.185 106.155 41.570 106.725 ;
        RECT 41.740 106.615 42.865 106.785 ;
        RECT 41.740 105.985 42.065 106.445 ;
        RECT 42.585 106.155 42.865 106.615 ;
        RECT 43.055 106.155 43.455 106.955 ;
        RECT 43.625 107.685 44.580 107.905 ;
        RECT 43.625 106.785 43.835 107.685 ;
        RECT 45.785 107.665 46.060 108.365 ;
        RECT 46.230 107.990 46.485 108.535 ;
        RECT 46.655 108.025 47.135 108.365 ;
        RECT 47.310 107.980 47.915 108.535 ;
        RECT 47.300 107.880 47.915 107.980 ;
        RECT 47.300 107.855 47.485 107.880 ;
        RECT 44.005 106.955 44.695 107.515 ;
        RECT 43.625 106.615 44.580 106.785 ;
        RECT 43.855 105.985 44.125 106.445 ;
        RECT 44.295 106.155 44.580 106.615 ;
        RECT 45.785 106.635 45.955 107.665 ;
        RECT 46.230 107.535 46.985 107.785 ;
        RECT 47.155 107.610 47.485 107.855 ;
        RECT 46.230 107.500 47.000 107.535 ;
        RECT 46.230 107.490 47.015 107.500 ;
        RECT 46.125 107.475 47.020 107.490 ;
        RECT 46.125 107.460 47.040 107.475 ;
        RECT 46.125 107.450 47.060 107.460 ;
        RECT 46.125 107.440 47.085 107.450 ;
        RECT 46.125 107.410 47.155 107.440 ;
        RECT 46.125 107.380 47.175 107.410 ;
        RECT 46.125 107.350 47.195 107.380 ;
        RECT 46.125 107.325 47.225 107.350 ;
        RECT 46.125 107.290 47.260 107.325 ;
        RECT 46.125 107.285 47.290 107.290 ;
        RECT 46.125 106.890 46.355 107.285 ;
        RECT 46.900 107.280 47.290 107.285 ;
        RECT 46.925 107.270 47.290 107.280 ;
        RECT 46.940 107.265 47.290 107.270 ;
        RECT 46.955 107.260 47.290 107.265 ;
        RECT 47.655 107.260 47.915 107.710 ;
        RECT 46.955 107.255 47.915 107.260 ;
        RECT 46.965 107.245 47.915 107.255 ;
        RECT 46.975 107.240 47.915 107.245 ;
        RECT 46.985 107.230 47.915 107.240 ;
        RECT 46.990 107.220 47.915 107.230 ;
        RECT 46.995 107.215 47.915 107.220 ;
        RECT 47.005 107.200 47.915 107.215 ;
        RECT 47.010 107.185 47.915 107.200 ;
        RECT 47.020 107.160 47.915 107.185 ;
        RECT 46.525 106.690 46.855 107.115 ;
        RECT 45.785 106.155 46.045 106.635 ;
        RECT 46.215 105.985 46.465 106.525 ;
        RECT 46.635 106.205 46.855 106.690 ;
        RECT 47.025 107.090 47.915 107.160 ;
        RECT 47.025 106.365 47.195 107.090 ;
        RECT 48.085 106.930 48.365 108.365 ;
        RECT 48.535 107.760 49.245 108.535 ;
        RECT 49.415 107.590 49.745 108.365 ;
        RECT 48.595 107.375 49.745 107.590 ;
        RECT 47.365 106.535 47.915 106.920 ;
        RECT 47.025 106.195 47.915 106.365 ;
        RECT 48.085 106.155 48.425 106.930 ;
        RECT 48.595 106.805 48.880 107.375 ;
        RECT 49.065 106.975 49.535 107.205 ;
        RECT 49.940 107.175 50.155 108.290 ;
        RECT 50.335 107.815 50.665 108.535 ;
        RECT 50.855 107.945 51.115 108.335 ;
        RECT 51.285 108.125 51.615 108.535 ;
        RECT 50.855 107.745 51.615 107.945 ;
        RECT 50.445 107.175 50.675 107.515 ;
        RECT 49.705 106.995 50.155 107.175 ;
        RECT 49.705 106.975 50.035 106.995 ;
        RECT 50.345 106.975 50.675 107.175 ;
        RECT 50.865 106.875 51.095 107.565 ;
        RECT 51.275 107.065 51.615 107.745 ;
        RECT 51.805 107.245 52.135 108.355 ;
        RECT 52.305 107.625 52.495 108.355 ;
        RECT 52.665 107.805 52.995 108.535 ;
        RECT 53.175 107.625 53.345 108.355 ;
        RECT 54.525 108.025 54.825 108.535 ;
        RECT 54.995 107.855 55.325 108.365 ;
        RECT 55.495 108.025 56.125 108.535 ;
        RECT 56.705 108.025 57.085 108.195 ;
        RECT 57.255 108.025 57.555 108.535 ;
        RECT 56.915 107.855 57.085 108.025 ;
        RECT 52.305 107.425 53.345 107.625 ;
        RECT 54.525 107.685 56.745 107.855 ;
        RECT 48.595 106.615 49.305 106.805 ;
        RECT 49.005 106.475 49.305 106.615 ;
        RECT 49.495 106.615 50.675 106.805 ;
        RECT 51.275 106.615 51.505 107.065 ;
        RECT 51.805 106.945 52.340 107.245 ;
        RECT 49.495 106.535 49.825 106.615 ;
        RECT 49.005 106.465 49.320 106.475 ;
        RECT 49.005 106.455 49.330 106.465 ;
        RECT 49.005 106.450 49.340 106.455 ;
        RECT 48.595 105.985 48.765 106.445 ;
        RECT 49.005 106.440 49.345 106.450 ;
        RECT 49.005 106.435 49.350 106.440 ;
        RECT 49.005 106.425 49.355 106.435 ;
        RECT 49.005 106.420 49.360 106.425 ;
        RECT 49.005 106.155 49.365 106.420 ;
        RECT 49.995 105.985 50.165 106.445 ;
        RECT 50.335 106.155 50.675 106.615 ;
        RECT 51.125 106.165 51.505 106.615 ;
        RECT 51.685 105.985 51.915 106.765 ;
        RECT 52.095 106.695 52.340 106.945 ;
        RECT 52.520 106.895 52.915 107.245 ;
        RECT 53.110 106.895 53.400 107.245 ;
        RECT 52.095 106.165 52.525 106.695 ;
        RECT 52.705 106.275 52.915 106.895 ;
        RECT 54.525 106.725 54.695 107.685 ;
        RECT 54.865 107.345 56.405 107.515 ;
        RECT 54.865 106.895 55.110 107.345 ;
        RECT 55.370 106.975 56.065 107.175 ;
        RECT 56.235 107.145 56.405 107.345 ;
        RECT 56.575 107.485 56.745 107.685 ;
        RECT 56.915 107.655 57.575 107.855 ;
        RECT 56.575 107.315 57.235 107.485 ;
        RECT 56.235 106.975 56.835 107.145 ;
        RECT 57.065 106.895 57.235 107.315 ;
        RECT 53.085 105.985 53.415 106.715 ;
        RECT 54.525 106.180 54.990 106.725 ;
        RECT 55.495 105.985 55.665 106.805 ;
        RECT 55.835 106.725 56.745 106.805 ;
        RECT 57.405 106.725 57.575 107.655 ;
        RECT 57.745 107.445 61.255 108.535 ;
        RECT 55.835 106.635 57.085 106.725 ;
        RECT 55.835 106.155 56.165 106.635 ;
        RECT 56.575 106.555 57.085 106.635 ;
        RECT 56.335 105.985 56.685 106.375 ;
        RECT 56.855 106.155 57.085 106.555 ;
        RECT 57.255 106.245 57.575 106.725 ;
        RECT 57.745 106.755 59.395 107.275 ;
        RECT 59.565 106.925 61.255 107.445 ;
        RECT 61.425 107.370 61.715 108.535 ;
        RECT 61.885 107.445 63.095 108.535 ;
        RECT 57.745 105.985 61.255 106.755 ;
        RECT 61.885 106.735 62.405 107.275 ;
        RECT 62.575 106.905 63.095 107.445 ;
        RECT 63.270 107.390 63.565 108.535 ;
        RECT 61.425 105.985 61.715 106.710 ;
        RECT 61.885 105.985 63.095 106.735 ;
        RECT 63.270 105.985 63.565 106.805 ;
        RECT 63.735 106.535 63.965 108.235 ;
        RECT 64.180 107.730 64.435 108.535 ;
        RECT 64.635 107.920 64.965 108.365 ;
        RECT 65.135 108.090 65.410 108.535 ;
        RECT 65.645 107.920 65.975 108.365 ;
        RECT 64.635 107.740 65.975 107.920 ;
        RECT 66.435 107.560 66.765 108.225 ;
        RECT 64.180 107.390 66.765 107.560 ;
        RECT 66.955 107.565 67.285 108.350 ;
        RECT 66.955 107.395 67.635 107.565 ;
        RECT 67.815 107.395 68.145 108.535 ;
        RECT 68.325 107.445 69.995 108.535 ;
        RECT 64.180 106.775 64.490 107.390 ;
        RECT 64.660 106.945 64.990 107.175 ;
        RECT 65.160 106.945 65.630 107.175 ;
        RECT 65.800 107.005 66.255 107.175 ;
        RECT 65.800 106.945 66.250 107.005 ;
        RECT 66.440 106.945 66.775 107.175 ;
        RECT 66.945 106.975 67.295 107.225 ;
        RECT 67.465 106.795 67.635 107.395 ;
        RECT 67.805 106.975 68.155 107.225 ;
        RECT 64.180 106.595 66.765 106.775 ;
        RECT 63.735 106.155 63.955 106.535 ;
        RECT 64.125 105.985 64.975 106.345 ;
        RECT 65.455 106.175 65.785 106.595 ;
        RECT 65.990 105.985 66.265 106.425 ;
        RECT 66.435 106.175 66.765 106.595 ;
        RECT 66.965 105.985 67.205 106.795 ;
        RECT 67.375 106.155 67.705 106.795 ;
        RECT 67.875 105.985 68.145 106.795 ;
        RECT 68.325 106.755 69.075 107.275 ;
        RECT 69.245 106.925 69.995 107.445 ;
        RECT 68.325 105.985 69.995 106.755 ;
        RECT 70.635 106.165 70.895 108.355 ;
        RECT 71.065 107.805 71.405 108.535 ;
        RECT 71.585 107.625 71.855 108.355 ;
        RECT 71.085 107.405 71.855 107.625 ;
        RECT 72.035 107.645 72.265 108.355 ;
        RECT 72.435 107.825 72.765 108.535 ;
        RECT 72.935 107.645 73.195 108.355 ;
        RECT 74.420 107.905 74.705 108.365 ;
        RECT 74.875 108.075 75.145 108.535 ;
        RECT 74.420 107.685 75.375 107.905 ;
        RECT 72.035 107.405 73.195 107.645 ;
        RECT 71.085 106.735 71.375 107.405 ;
        RECT 71.555 106.915 72.020 107.225 ;
        RECT 72.200 106.915 72.725 107.225 ;
        RECT 71.085 106.535 72.315 106.735 ;
        RECT 71.155 105.985 71.825 106.355 ;
        RECT 72.005 106.165 72.315 106.535 ;
        RECT 72.495 106.275 72.725 106.915 ;
        RECT 72.905 106.895 73.205 107.225 ;
        RECT 74.305 106.955 74.995 107.515 ;
        RECT 75.165 106.785 75.375 107.685 ;
        RECT 72.905 105.985 73.195 106.715 ;
        RECT 74.420 106.615 75.375 106.785 ;
        RECT 75.545 107.515 75.945 108.365 ;
        RECT 76.135 107.905 76.415 108.365 ;
        RECT 76.935 108.075 77.260 108.535 ;
        RECT 76.135 107.685 77.260 107.905 ;
        RECT 75.545 106.955 76.640 107.515 ;
        RECT 76.810 107.225 77.260 107.685 ;
        RECT 77.430 107.395 77.815 108.365 ;
        RECT 74.420 106.155 74.705 106.615 ;
        RECT 74.875 105.985 75.145 106.445 ;
        RECT 75.545 106.155 75.945 106.955 ;
        RECT 76.810 106.895 77.365 107.225 ;
        RECT 76.810 106.785 77.260 106.895 ;
        RECT 76.135 106.615 77.260 106.785 ;
        RECT 77.535 106.725 77.815 107.395 ;
        RECT 77.990 107.390 78.285 108.535 ;
        RECT 76.135 106.155 76.415 106.615 ;
        RECT 76.935 105.985 77.260 106.445 ;
        RECT 77.430 106.155 77.815 106.725 ;
        RECT 77.990 105.985 78.285 106.805 ;
        RECT 78.455 106.535 78.685 108.235 ;
        RECT 78.900 107.730 79.155 108.535 ;
        RECT 79.355 107.920 79.685 108.365 ;
        RECT 79.855 108.090 80.130 108.535 ;
        RECT 80.365 107.920 80.695 108.365 ;
        RECT 79.355 107.740 80.695 107.920 ;
        RECT 81.155 107.560 81.485 108.225 ;
        RECT 78.900 107.390 81.485 107.560 ;
        RECT 81.665 107.395 82.050 108.365 ;
        RECT 82.220 108.075 82.545 108.535 ;
        RECT 83.065 107.905 83.345 108.365 ;
        RECT 82.220 107.685 83.345 107.905 ;
        RECT 78.900 106.775 79.210 107.390 ;
        RECT 79.380 106.945 79.710 107.175 ;
        RECT 79.880 106.945 80.350 107.175 ;
        RECT 80.520 107.005 80.975 107.175 ;
        RECT 80.520 106.945 80.970 107.005 ;
        RECT 81.160 106.945 81.495 107.175 ;
        RECT 78.900 106.595 81.485 106.775 ;
        RECT 78.455 106.155 78.675 106.535 ;
        RECT 78.845 105.985 79.695 106.345 ;
        RECT 80.175 106.175 80.505 106.595 ;
        RECT 80.710 105.985 80.985 106.425 ;
        RECT 81.155 106.175 81.485 106.595 ;
        RECT 81.665 106.725 81.945 107.395 ;
        RECT 82.220 107.225 82.670 107.685 ;
        RECT 83.535 107.515 83.935 108.365 ;
        RECT 84.335 108.075 84.605 108.535 ;
        RECT 84.775 107.905 85.060 108.365 ;
        RECT 82.115 106.895 82.670 107.225 ;
        RECT 82.840 106.955 83.935 107.515 ;
        RECT 82.220 106.785 82.670 106.895 ;
        RECT 81.665 106.155 82.050 106.725 ;
        RECT 82.220 106.615 83.345 106.785 ;
        RECT 82.220 105.985 82.545 106.445 ;
        RECT 83.065 106.155 83.345 106.615 ;
        RECT 83.535 106.155 83.935 106.955 ;
        RECT 84.105 107.685 85.060 107.905 ;
        RECT 84.105 106.785 84.315 107.685 ;
        RECT 85.355 107.565 85.685 108.350 ;
        RECT 84.485 106.955 85.175 107.515 ;
        RECT 85.355 107.395 86.035 107.565 ;
        RECT 86.215 107.395 86.545 108.535 ;
        RECT 85.345 106.975 85.695 107.225 ;
        RECT 85.865 106.795 86.035 107.395 ;
        RECT 87.185 107.370 87.475 108.535 ;
        RECT 86.205 106.975 86.555 107.225 ;
        RECT 84.105 106.615 85.060 106.785 ;
        RECT 84.335 105.985 84.605 106.445 ;
        RECT 84.775 106.155 85.060 106.615 ;
        RECT 85.365 105.985 85.605 106.795 ;
        RECT 85.775 106.155 86.105 106.795 ;
        RECT 86.275 105.985 86.545 106.795 ;
        RECT 87.185 105.985 87.475 106.710 ;
        RECT 88.115 106.165 88.375 108.355 ;
        RECT 88.545 107.805 88.885 108.535 ;
        RECT 89.065 107.625 89.335 108.355 ;
        RECT 88.565 107.405 89.335 107.625 ;
        RECT 89.515 107.645 89.745 108.355 ;
        RECT 89.915 107.825 90.245 108.535 ;
        RECT 90.415 107.645 90.675 108.355 ;
        RECT 89.515 107.405 90.675 107.645 ;
        RECT 90.865 107.665 91.140 108.365 ;
        RECT 91.310 107.990 91.565 108.535 ;
        RECT 91.735 108.025 92.215 108.365 ;
        RECT 92.390 107.980 92.995 108.535 ;
        RECT 92.380 107.880 92.995 107.980 ;
        RECT 92.380 107.855 92.565 107.880 ;
        RECT 88.565 106.735 88.855 107.405 ;
        RECT 89.035 106.915 89.500 107.225 ;
        RECT 89.680 106.915 90.205 107.225 ;
        RECT 88.565 106.535 89.795 106.735 ;
        RECT 88.635 105.985 89.305 106.355 ;
        RECT 89.485 106.165 89.795 106.535 ;
        RECT 89.975 106.275 90.205 106.915 ;
        RECT 90.385 106.895 90.685 107.225 ;
        RECT 90.385 105.985 90.675 106.715 ;
        RECT 90.865 106.635 91.035 107.665 ;
        RECT 91.310 107.535 92.065 107.785 ;
        RECT 92.235 107.610 92.565 107.855 ;
        RECT 91.310 107.500 92.080 107.535 ;
        RECT 91.310 107.490 92.095 107.500 ;
        RECT 91.205 107.475 92.100 107.490 ;
        RECT 91.205 107.460 92.120 107.475 ;
        RECT 91.205 107.450 92.140 107.460 ;
        RECT 91.205 107.440 92.165 107.450 ;
        RECT 91.205 107.410 92.235 107.440 ;
        RECT 91.205 107.380 92.255 107.410 ;
        RECT 91.205 107.350 92.275 107.380 ;
        RECT 91.205 107.325 92.305 107.350 ;
        RECT 91.205 107.290 92.340 107.325 ;
        RECT 91.205 107.285 92.370 107.290 ;
        RECT 91.205 106.890 91.435 107.285 ;
        RECT 91.980 107.280 92.370 107.285 ;
        RECT 92.005 107.270 92.370 107.280 ;
        RECT 92.020 107.265 92.370 107.270 ;
        RECT 92.035 107.260 92.370 107.265 ;
        RECT 92.735 107.260 92.995 107.710 ;
        RECT 93.165 107.445 95.755 108.535 ;
        RECT 92.035 107.255 92.995 107.260 ;
        RECT 92.045 107.245 92.995 107.255 ;
        RECT 92.055 107.240 92.995 107.245 ;
        RECT 92.065 107.230 92.995 107.240 ;
        RECT 92.070 107.220 92.995 107.230 ;
        RECT 92.075 107.215 92.995 107.220 ;
        RECT 92.085 107.200 92.995 107.215 ;
        RECT 92.090 107.185 92.995 107.200 ;
        RECT 92.100 107.160 92.995 107.185 ;
        RECT 91.605 106.690 91.935 107.115 ;
        RECT 90.865 106.155 91.125 106.635 ;
        RECT 91.295 105.985 91.545 106.525 ;
        RECT 91.715 106.205 91.935 106.690 ;
        RECT 92.105 107.090 92.995 107.160 ;
        RECT 92.105 106.365 92.275 107.090 ;
        RECT 92.445 106.535 92.995 106.920 ;
        RECT 93.165 106.755 94.375 107.275 ;
        RECT 94.545 106.925 95.755 107.445 ;
        RECT 96.390 107.390 96.685 108.535 ;
        RECT 92.105 106.195 92.995 106.365 ;
        RECT 93.165 105.985 95.755 106.755 ;
        RECT 96.390 105.985 96.685 106.805 ;
        RECT 96.855 106.535 97.085 108.235 ;
        RECT 97.300 107.730 97.555 108.535 ;
        RECT 97.755 107.920 98.085 108.365 ;
        RECT 98.255 108.090 98.530 108.535 ;
        RECT 98.765 107.920 99.095 108.365 ;
        RECT 97.755 107.740 99.095 107.920 ;
        RECT 99.555 107.560 99.885 108.225 ;
        RECT 100.065 107.980 100.670 108.535 ;
        RECT 100.845 108.025 101.325 108.365 ;
        RECT 101.495 107.990 101.750 108.535 ;
        RECT 100.065 107.880 100.680 107.980 ;
        RECT 100.495 107.855 100.680 107.880 ;
        RECT 97.300 107.390 99.885 107.560 ;
        RECT 97.300 106.775 97.610 107.390 ;
        RECT 100.065 107.260 100.325 107.710 ;
        RECT 100.495 107.610 100.825 107.855 ;
        RECT 100.995 107.535 101.750 107.785 ;
        RECT 101.920 107.665 102.195 108.365 ;
        RECT 100.980 107.500 101.750 107.535 ;
        RECT 100.965 107.490 101.750 107.500 ;
        RECT 100.960 107.475 101.855 107.490 ;
        RECT 100.940 107.460 101.855 107.475 ;
        RECT 100.920 107.450 101.855 107.460 ;
        RECT 100.895 107.440 101.855 107.450 ;
        RECT 100.825 107.410 101.855 107.440 ;
        RECT 100.805 107.380 101.855 107.410 ;
        RECT 100.785 107.350 101.855 107.380 ;
        RECT 100.755 107.325 101.855 107.350 ;
        RECT 100.720 107.290 101.855 107.325 ;
        RECT 100.690 107.285 101.855 107.290 ;
        RECT 100.690 107.280 101.080 107.285 ;
        RECT 100.690 107.270 101.055 107.280 ;
        RECT 100.690 107.265 101.040 107.270 ;
        RECT 100.690 107.260 101.025 107.265 ;
        RECT 100.065 107.255 101.025 107.260 ;
        RECT 100.065 107.245 101.015 107.255 ;
        RECT 100.065 107.240 101.005 107.245 ;
        RECT 100.065 107.230 100.995 107.240 ;
        RECT 100.065 107.220 100.990 107.230 ;
        RECT 100.065 107.215 100.985 107.220 ;
        RECT 100.065 107.200 100.975 107.215 ;
        RECT 100.065 107.185 100.970 107.200 ;
        RECT 97.780 106.945 98.110 107.175 ;
        RECT 98.280 106.945 98.750 107.175 ;
        RECT 98.920 107.005 99.375 107.175 ;
        RECT 98.920 106.945 99.370 107.005 ;
        RECT 99.560 106.945 99.895 107.175 ;
        RECT 100.065 107.160 100.960 107.185 ;
        RECT 100.065 107.090 100.955 107.160 ;
        RECT 97.300 106.595 99.885 106.775 ;
        RECT 96.855 106.155 97.075 106.535 ;
        RECT 97.245 105.985 98.095 106.345 ;
        RECT 98.575 106.175 98.905 106.595 ;
        RECT 99.110 105.985 99.385 106.425 ;
        RECT 99.555 106.175 99.885 106.595 ;
        RECT 100.065 106.535 100.615 106.920 ;
        RECT 100.785 106.365 100.955 107.090 ;
        RECT 100.065 106.195 100.955 106.365 ;
        RECT 101.125 106.690 101.455 107.115 ;
        RECT 101.625 106.890 101.855 107.285 ;
        RECT 101.125 106.205 101.345 106.690 ;
        RECT 102.025 106.635 102.195 107.665 ;
        RECT 101.515 105.985 101.765 106.525 ;
        RECT 101.935 106.155 102.195 106.635 ;
        RECT 102.365 107.395 102.750 108.365 ;
        RECT 102.920 108.075 103.245 108.535 ;
        RECT 103.765 107.905 104.045 108.365 ;
        RECT 102.920 107.685 104.045 107.905 ;
        RECT 102.365 106.725 102.645 107.395 ;
        RECT 102.920 107.225 103.370 107.685 ;
        RECT 104.235 107.515 104.635 108.365 ;
        RECT 105.035 108.075 105.305 108.535 ;
        RECT 105.475 107.905 105.760 108.365 ;
        RECT 102.815 106.895 103.370 107.225 ;
        RECT 103.540 106.955 104.635 107.515 ;
        RECT 102.920 106.785 103.370 106.895 ;
        RECT 102.365 106.155 102.750 106.725 ;
        RECT 102.920 106.615 104.045 106.785 ;
        RECT 102.920 105.985 103.245 106.445 ;
        RECT 103.765 106.155 104.045 106.615 ;
        RECT 104.235 106.155 104.635 106.955 ;
        RECT 104.805 107.685 105.760 107.905 ;
        RECT 104.805 106.785 105.015 107.685 ;
        RECT 105.185 106.955 105.875 107.515 ;
        RECT 106.045 107.425 106.305 108.365 ;
        RECT 106.475 108.135 106.805 108.535 ;
        RECT 107.950 108.270 108.205 108.365 ;
        RECT 107.065 108.100 108.205 108.270 ;
        RECT 108.375 108.155 108.705 108.325 ;
        RECT 107.065 107.875 107.235 108.100 ;
        RECT 106.475 107.705 107.235 107.875 ;
        RECT 107.950 107.965 108.205 108.100 ;
        RECT 104.805 106.615 105.760 106.785 ;
        RECT 105.035 105.985 105.305 106.445 ;
        RECT 105.475 106.155 105.760 106.615 ;
        RECT 106.045 106.710 106.220 107.425 ;
        RECT 106.475 107.225 106.645 107.705 ;
        RECT 107.500 107.615 107.670 107.805 ;
        RECT 107.950 107.795 108.360 107.965 ;
        RECT 106.390 106.895 106.645 107.225 ;
        RECT 106.870 106.895 107.200 107.515 ;
        RECT 107.500 107.445 108.020 107.615 ;
        RECT 107.370 106.895 107.660 107.275 ;
        RECT 107.850 106.725 108.020 107.445 ;
        RECT 106.045 106.155 106.305 106.710 ;
        RECT 107.140 106.555 108.020 106.725 ;
        RECT 108.190 106.770 108.360 107.795 ;
        RECT 108.535 107.905 108.705 108.155 ;
        RECT 108.875 108.075 109.125 108.535 ;
        RECT 109.295 107.905 109.475 108.365 ;
        RECT 108.535 107.735 109.475 107.905 ;
        RECT 108.560 107.255 109.040 107.555 ;
        RECT 108.190 106.600 108.540 106.770 ;
        RECT 108.780 106.665 109.040 107.255 ;
        RECT 109.240 106.665 109.500 107.555 ;
        RECT 106.475 105.985 106.905 106.430 ;
        RECT 107.140 106.155 107.310 106.555 ;
        RECT 107.480 105.985 108.200 106.385 ;
        RECT 108.370 106.155 108.540 106.600 ;
        RECT 109.115 105.985 109.515 106.495 ;
        RECT 109.735 106.165 109.995 108.355 ;
        RECT 110.165 107.805 110.505 108.535 ;
        RECT 110.685 107.625 110.955 108.355 ;
        RECT 110.185 107.405 110.955 107.625 ;
        RECT 111.135 107.645 111.365 108.355 ;
        RECT 111.535 107.825 111.865 108.535 ;
        RECT 112.035 107.645 112.295 108.355 ;
        RECT 111.135 107.405 112.295 107.645 ;
        RECT 110.185 106.735 110.475 107.405 ;
        RECT 112.945 107.370 113.235 108.535 ;
        RECT 113.495 107.865 113.665 108.365 ;
        RECT 113.835 108.035 114.165 108.535 ;
        RECT 113.495 107.695 114.160 107.865 ;
        RECT 110.655 106.915 111.120 107.225 ;
        RECT 111.300 106.915 111.825 107.225 ;
        RECT 110.185 106.535 111.415 106.735 ;
        RECT 110.255 105.985 110.925 106.355 ;
        RECT 111.105 106.165 111.415 106.535 ;
        RECT 111.595 106.275 111.825 106.915 ;
        RECT 112.005 106.895 112.305 107.225 ;
        RECT 113.410 106.875 113.760 107.525 ;
        RECT 112.005 105.985 112.295 106.715 ;
        RECT 112.945 105.985 113.235 106.710 ;
        RECT 113.930 106.705 114.160 107.695 ;
        RECT 113.495 106.535 114.160 106.705 ;
        RECT 113.495 106.245 113.665 106.535 ;
        RECT 113.835 105.985 114.165 106.365 ;
        RECT 114.335 106.245 114.520 108.365 ;
        RECT 114.760 108.075 115.025 108.535 ;
        RECT 115.195 107.940 115.445 108.365 ;
        RECT 115.655 108.090 116.760 108.260 ;
        RECT 115.140 107.810 115.445 107.940 ;
        RECT 114.690 106.615 114.970 107.565 ;
        RECT 115.140 106.705 115.310 107.810 ;
        RECT 115.480 107.025 115.720 107.620 ;
        RECT 115.890 107.555 116.420 107.920 ;
        RECT 115.890 106.855 116.060 107.555 ;
        RECT 116.590 107.475 116.760 108.090 ;
        RECT 116.930 107.735 117.100 108.535 ;
        RECT 117.270 108.035 117.520 108.365 ;
        RECT 117.745 108.065 118.630 108.235 ;
        RECT 116.590 107.385 117.100 107.475 ;
        RECT 115.140 106.575 115.365 106.705 ;
        RECT 115.535 106.635 116.060 106.855 ;
        RECT 116.230 107.215 117.100 107.385 ;
        RECT 114.775 105.985 115.025 106.445 ;
        RECT 115.195 106.435 115.365 106.575 ;
        RECT 116.230 106.435 116.400 107.215 ;
        RECT 116.930 107.145 117.100 107.215 ;
        RECT 116.610 106.965 116.810 106.995 ;
        RECT 117.270 106.965 117.440 108.035 ;
        RECT 117.610 107.145 117.800 107.865 ;
        RECT 116.610 106.665 117.440 106.965 ;
        RECT 117.970 106.935 118.290 107.895 ;
        RECT 115.195 106.265 115.530 106.435 ;
        RECT 115.725 106.265 116.400 106.435 ;
        RECT 116.720 105.985 117.090 106.485 ;
        RECT 117.270 106.435 117.440 106.665 ;
        RECT 117.825 106.605 118.290 106.935 ;
        RECT 118.460 107.225 118.630 108.065 ;
        RECT 118.810 108.035 119.125 108.535 ;
        RECT 119.355 107.805 119.695 108.365 ;
        RECT 118.800 107.430 119.695 107.805 ;
        RECT 119.865 107.525 120.035 108.535 ;
        RECT 119.505 107.225 119.695 107.430 ;
        RECT 120.205 107.475 120.535 108.320 ;
        RECT 120.775 107.585 121.050 108.355 ;
        RECT 121.220 107.925 121.550 108.355 ;
        RECT 121.720 108.095 121.915 108.535 ;
        RECT 122.095 107.925 122.425 108.355 ;
        RECT 121.220 107.755 122.425 107.925 ;
        RECT 120.205 107.395 120.595 107.475 ;
        RECT 120.775 107.395 121.360 107.585 ;
        RECT 121.530 107.425 122.425 107.755 ;
        RECT 123.125 107.475 123.455 108.320 ;
        RECT 123.625 107.525 123.795 108.535 ;
        RECT 123.965 107.805 124.305 108.365 ;
        RECT 124.535 108.035 124.850 108.535 ;
        RECT 125.030 108.065 125.915 108.235 ;
        RECT 120.380 107.345 120.595 107.395 ;
        RECT 118.460 106.895 119.335 107.225 ;
        RECT 119.505 106.895 120.255 107.225 ;
        RECT 118.460 106.435 118.630 106.895 ;
        RECT 119.505 106.725 119.705 106.895 ;
        RECT 120.425 106.765 120.595 107.345 ;
        RECT 120.370 106.725 120.595 106.765 ;
        RECT 117.270 106.265 117.675 106.435 ;
        RECT 117.845 106.265 118.630 106.435 ;
        RECT 118.905 105.985 119.115 106.515 ;
        RECT 119.375 106.200 119.705 106.725 ;
        RECT 120.215 106.640 120.595 106.725 ;
        RECT 119.875 105.985 120.045 106.595 ;
        RECT 120.215 106.205 120.545 106.640 ;
        RECT 120.775 106.575 121.015 107.225 ;
        RECT 121.185 106.725 121.360 107.395 ;
        RECT 123.065 107.395 123.455 107.475 ;
        RECT 123.965 107.430 124.860 107.805 ;
        RECT 123.065 107.345 123.280 107.395 ;
        RECT 121.530 106.895 121.945 107.225 ;
        RECT 122.125 106.895 122.420 107.225 ;
        RECT 121.185 106.545 121.515 106.725 ;
        RECT 120.790 105.985 121.120 106.375 ;
        RECT 121.290 106.165 121.515 106.545 ;
        RECT 121.715 106.275 121.945 106.895 ;
        RECT 123.065 106.765 123.235 107.345 ;
        RECT 123.965 107.225 124.155 107.430 ;
        RECT 125.030 107.225 125.200 108.065 ;
        RECT 126.140 108.035 126.390 108.365 ;
        RECT 123.405 106.895 124.155 107.225 ;
        RECT 124.325 106.895 125.200 107.225 ;
        RECT 123.065 106.725 123.290 106.765 ;
        RECT 123.955 106.725 124.155 106.895 ;
        RECT 122.125 105.985 122.425 106.715 ;
        RECT 123.065 106.640 123.445 106.725 ;
        RECT 123.115 106.205 123.445 106.640 ;
        RECT 123.615 105.985 123.785 106.595 ;
        RECT 123.955 106.200 124.285 106.725 ;
        RECT 124.545 105.985 124.755 106.515 ;
        RECT 125.030 106.435 125.200 106.895 ;
        RECT 125.370 106.935 125.690 107.895 ;
        RECT 125.860 107.145 126.050 107.865 ;
        RECT 126.220 106.965 126.390 108.035 ;
        RECT 126.560 107.735 126.730 108.535 ;
        RECT 126.900 108.090 128.005 108.260 ;
        RECT 126.900 107.475 127.070 108.090 ;
        RECT 128.215 107.940 128.465 108.365 ;
        RECT 128.635 108.075 128.900 108.535 ;
        RECT 127.240 107.555 127.770 107.920 ;
        RECT 128.215 107.810 128.520 107.940 ;
        RECT 126.560 107.385 127.070 107.475 ;
        RECT 126.560 107.215 127.430 107.385 ;
        RECT 126.560 107.145 126.730 107.215 ;
        RECT 126.850 106.965 127.050 106.995 ;
        RECT 125.370 106.605 125.835 106.935 ;
        RECT 126.220 106.665 127.050 106.965 ;
        RECT 126.220 106.435 126.390 106.665 ;
        RECT 125.030 106.265 125.815 106.435 ;
        RECT 125.985 106.265 126.390 106.435 ;
        RECT 126.570 105.985 126.940 106.485 ;
        RECT 127.260 106.435 127.430 107.215 ;
        RECT 127.600 106.855 127.770 107.555 ;
        RECT 127.940 107.025 128.180 107.620 ;
        RECT 127.600 106.635 128.125 106.855 ;
        RECT 128.350 106.705 128.520 107.810 ;
        RECT 128.295 106.575 128.520 106.705 ;
        RECT 128.690 106.615 128.970 107.565 ;
        RECT 128.295 106.435 128.465 106.575 ;
        RECT 127.260 106.265 127.935 106.435 ;
        RECT 128.130 106.265 128.465 106.435 ;
        RECT 128.635 105.985 128.885 106.445 ;
        RECT 129.140 106.245 129.325 108.365 ;
        RECT 129.495 108.035 129.825 108.535 ;
        RECT 129.995 107.865 130.165 108.365 ;
        RECT 129.500 107.695 130.165 107.865 ;
        RECT 130.540 107.905 130.825 108.365 ;
        RECT 130.995 108.075 131.265 108.535 ;
        RECT 129.500 106.705 129.730 107.695 ;
        RECT 130.540 107.685 131.495 107.905 ;
        RECT 129.900 106.875 130.250 107.525 ;
        RECT 130.425 106.955 131.115 107.515 ;
        RECT 131.285 106.785 131.495 107.685 ;
        RECT 129.500 106.535 130.165 106.705 ;
        RECT 129.495 105.985 129.825 106.365 ;
        RECT 129.995 106.245 130.165 106.535 ;
        RECT 130.540 106.615 131.495 106.785 ;
        RECT 131.665 107.515 132.065 108.365 ;
        RECT 132.255 107.905 132.535 108.365 ;
        RECT 133.055 108.075 133.380 108.535 ;
        RECT 132.255 107.685 133.380 107.905 ;
        RECT 131.665 106.955 132.760 107.515 ;
        RECT 132.930 107.225 133.380 107.685 ;
        RECT 133.550 107.395 133.935 108.365 ;
        RECT 130.540 106.155 130.825 106.615 ;
        RECT 130.995 105.985 131.265 106.445 ;
        RECT 131.665 106.155 132.065 106.955 ;
        RECT 132.930 106.895 133.485 107.225 ;
        RECT 132.930 106.785 133.380 106.895 ;
        RECT 132.255 106.615 133.380 106.785 ;
        RECT 133.655 106.725 133.935 107.395 ;
        RECT 132.255 106.155 132.535 106.615 ;
        RECT 133.055 105.985 133.380 106.445 ;
        RECT 133.550 106.155 133.935 106.725 ;
        RECT 134.105 107.395 134.445 108.365 ;
        RECT 134.615 107.395 134.785 108.535 ;
        RECT 135.055 107.735 135.305 108.535 ;
        RECT 135.950 107.565 136.280 108.365 ;
        RECT 136.580 107.735 136.910 108.535 ;
        RECT 137.080 107.565 137.410 108.365 ;
        RECT 134.975 107.395 137.410 107.565 ;
        RECT 134.105 106.835 134.280 107.395 ;
        RECT 134.975 107.145 135.145 107.395 ;
        RECT 134.450 106.975 135.145 107.145 ;
        RECT 135.320 106.975 135.740 107.175 ;
        RECT 135.910 106.975 136.240 107.175 ;
        RECT 136.410 106.975 136.740 107.175 ;
        RECT 134.105 106.785 134.335 106.835 ;
        RECT 134.105 106.155 134.445 106.785 ;
        RECT 134.615 105.985 134.865 106.785 ;
        RECT 135.055 106.635 136.280 106.805 ;
        RECT 135.055 106.155 135.385 106.635 ;
        RECT 135.555 105.985 135.780 106.445 ;
        RECT 135.950 106.155 136.280 106.635 ;
        RECT 136.910 106.765 137.080 107.395 ;
        RECT 138.705 107.370 138.995 108.535 ;
        RECT 139.165 107.445 140.835 108.535 ;
        RECT 141.120 107.905 141.405 108.365 ;
        RECT 141.575 108.075 141.845 108.535 ;
        RECT 141.120 107.685 142.075 107.905 ;
        RECT 137.265 106.975 137.615 107.225 ;
        RECT 136.910 106.155 137.410 106.765 ;
        RECT 139.165 106.755 139.915 107.275 ;
        RECT 140.085 106.925 140.835 107.445 ;
        RECT 141.005 106.955 141.695 107.515 ;
        RECT 141.865 106.785 142.075 107.685 ;
        RECT 138.705 105.985 138.995 106.710 ;
        RECT 139.165 105.985 140.835 106.755 ;
        RECT 141.120 106.615 142.075 106.785 ;
        RECT 142.245 107.515 142.645 108.365 ;
        RECT 142.835 107.905 143.115 108.365 ;
        RECT 143.635 108.075 143.960 108.535 ;
        RECT 142.835 107.685 143.960 107.905 ;
        RECT 142.245 106.955 143.340 107.515 ;
        RECT 143.510 107.225 143.960 107.685 ;
        RECT 144.130 107.395 144.515 108.365 ;
        RECT 141.120 106.155 141.405 106.615 ;
        RECT 141.575 105.985 141.845 106.445 ;
        RECT 142.245 106.155 142.645 106.955 ;
        RECT 143.510 106.895 144.065 107.225 ;
        RECT 143.510 106.785 143.960 106.895 ;
        RECT 142.835 106.615 143.960 106.785 ;
        RECT 144.235 106.725 144.515 107.395 ;
        RECT 142.835 106.155 143.115 106.615 ;
        RECT 143.635 105.985 143.960 106.445 ;
        RECT 144.130 106.155 144.515 106.725 ;
        RECT 144.685 107.395 144.955 108.365 ;
        RECT 145.165 107.735 145.445 108.535 ;
        RECT 145.615 108.025 147.270 108.315 ;
        RECT 147.535 107.865 147.705 108.365 ;
        RECT 147.875 108.035 148.205 108.535 ;
        RECT 145.680 107.685 147.270 107.855 ;
        RECT 147.535 107.695 148.200 107.865 ;
        RECT 145.680 107.565 145.850 107.685 ;
        RECT 145.125 107.395 145.850 107.565 ;
        RECT 144.685 106.660 144.855 107.395 ;
        RECT 145.125 107.225 145.295 107.395 ;
        RECT 145.025 106.895 145.295 107.225 ;
        RECT 145.465 106.895 145.870 107.225 ;
        RECT 146.040 106.895 146.750 107.515 ;
        RECT 146.950 107.395 147.270 107.685 ;
        RECT 145.125 106.725 145.295 106.895 ;
        RECT 144.685 106.315 144.955 106.660 ;
        RECT 145.125 106.555 146.735 106.725 ;
        RECT 146.920 106.655 147.270 107.225 ;
        RECT 147.450 106.875 147.800 107.525 ;
        RECT 147.970 106.705 148.200 107.695 ;
        RECT 145.145 105.985 145.525 106.385 ;
        RECT 145.695 106.205 145.865 106.555 ;
        RECT 146.035 105.985 146.365 106.385 ;
        RECT 146.565 106.205 146.735 106.555 ;
        RECT 147.535 106.535 148.200 106.705 ;
        RECT 146.935 105.985 147.265 106.485 ;
        RECT 147.535 106.245 147.705 106.535 ;
        RECT 147.875 105.985 148.205 106.365 ;
        RECT 148.375 106.245 148.560 108.365 ;
        RECT 148.800 108.075 149.065 108.535 ;
        RECT 149.235 107.940 149.485 108.365 ;
        RECT 149.695 108.090 150.800 108.260 ;
        RECT 149.180 107.810 149.485 107.940 ;
        RECT 148.730 106.615 149.010 107.565 ;
        RECT 149.180 106.705 149.350 107.810 ;
        RECT 149.520 107.025 149.760 107.620 ;
        RECT 149.930 107.555 150.460 107.920 ;
        RECT 149.930 106.855 150.100 107.555 ;
        RECT 150.630 107.475 150.800 108.090 ;
        RECT 150.970 107.735 151.140 108.535 ;
        RECT 151.310 108.035 151.560 108.365 ;
        RECT 151.785 108.065 152.670 108.235 ;
        RECT 150.630 107.385 151.140 107.475 ;
        RECT 149.180 106.575 149.405 106.705 ;
        RECT 149.575 106.635 150.100 106.855 ;
        RECT 150.270 107.215 151.140 107.385 ;
        RECT 148.815 105.985 149.065 106.445 ;
        RECT 149.235 106.435 149.405 106.575 ;
        RECT 150.270 106.435 150.440 107.215 ;
        RECT 150.970 107.145 151.140 107.215 ;
        RECT 150.650 106.965 150.850 106.995 ;
        RECT 151.310 106.965 151.480 108.035 ;
        RECT 151.650 107.145 151.840 107.865 ;
        RECT 150.650 106.665 151.480 106.965 ;
        RECT 152.010 106.935 152.330 107.895 ;
        RECT 149.235 106.265 149.570 106.435 ;
        RECT 149.765 106.265 150.440 106.435 ;
        RECT 150.760 105.985 151.130 106.485 ;
        RECT 151.310 106.435 151.480 106.665 ;
        RECT 151.865 106.605 152.330 106.935 ;
        RECT 152.500 107.225 152.670 108.065 ;
        RECT 152.850 108.035 153.165 108.535 ;
        RECT 153.395 107.805 153.735 108.365 ;
        RECT 152.840 107.430 153.735 107.805 ;
        RECT 153.905 107.525 154.075 108.535 ;
        RECT 153.545 107.225 153.735 107.430 ;
        RECT 154.245 107.475 154.575 108.320 ;
        RECT 154.245 107.395 154.635 107.475 ;
        RECT 154.420 107.345 154.635 107.395 ;
        RECT 152.500 106.895 153.375 107.225 ;
        RECT 153.545 106.895 154.295 107.225 ;
        RECT 152.500 106.435 152.670 106.895 ;
        RECT 153.545 106.725 153.745 106.895 ;
        RECT 154.465 106.765 154.635 107.345 ;
        RECT 155.725 107.445 156.935 108.535 ;
        RECT 155.725 106.905 156.245 107.445 ;
        RECT 154.410 106.725 154.635 106.765 ;
        RECT 156.415 106.735 156.935 107.275 ;
        RECT 151.310 106.265 151.715 106.435 ;
        RECT 151.885 106.265 152.670 106.435 ;
        RECT 152.945 105.985 153.155 106.515 ;
        RECT 153.415 106.200 153.745 106.725 ;
        RECT 154.255 106.640 154.635 106.725 ;
        RECT 153.915 105.985 154.085 106.595 ;
        RECT 154.255 106.205 154.585 106.640 ;
        RECT 155.725 105.985 156.935 106.735 ;
        RECT 22.700 105.815 157.020 105.985 ;
        RECT 22.785 105.065 23.995 105.815 ;
        RECT 24.165 105.270 29.510 105.815 ;
        RECT 30.935 105.415 31.265 105.815 ;
        RECT 22.785 104.525 23.305 105.065 ;
        RECT 23.475 104.355 23.995 104.895 ;
        RECT 25.750 104.440 26.090 105.270 ;
        RECT 31.435 105.245 31.765 105.585 ;
        RECT 32.815 105.415 33.145 105.815 ;
        RECT 30.780 105.075 33.145 105.245 ;
        RECT 33.315 105.090 33.645 105.600 ;
        RECT 33.915 105.265 34.085 105.555 ;
        RECT 34.255 105.435 34.585 105.815 ;
        RECT 33.915 105.095 34.580 105.265 ;
        RECT 22.785 103.265 23.995 104.355 ;
        RECT 27.570 103.700 27.920 104.950 ;
        RECT 30.780 104.075 30.950 105.075 ;
        RECT 32.975 104.905 33.145 105.075 ;
        RECT 31.120 104.245 31.365 104.905 ;
        RECT 31.580 104.245 31.845 104.905 ;
        RECT 32.040 104.245 32.325 104.905 ;
        RECT 32.500 104.575 32.805 104.905 ;
        RECT 32.975 104.575 33.285 104.905 ;
        RECT 32.500 104.245 32.715 104.575 ;
        RECT 30.780 103.905 31.235 104.075 ;
        RECT 24.165 103.265 29.510 103.700 ;
        RECT 30.905 103.475 31.235 103.905 ;
        RECT 31.415 103.905 32.705 104.075 ;
        RECT 31.415 103.485 31.665 103.905 ;
        RECT 31.895 103.265 32.225 103.735 ;
        RECT 32.455 103.485 32.705 103.905 ;
        RECT 32.895 103.265 33.145 104.405 ;
        RECT 33.455 104.325 33.645 105.090 ;
        RECT 33.315 103.475 33.645 104.325 ;
        RECT 33.830 104.275 34.180 104.925 ;
        RECT 34.350 104.105 34.580 105.095 ;
        RECT 33.915 103.935 34.580 104.105 ;
        RECT 33.915 103.435 34.085 103.935 ;
        RECT 34.255 103.265 34.585 103.765 ;
        RECT 34.755 103.435 34.940 105.555 ;
        RECT 35.195 105.355 35.445 105.815 ;
        RECT 35.615 105.365 35.950 105.535 ;
        RECT 36.145 105.365 36.820 105.535 ;
        RECT 35.615 105.225 35.785 105.365 ;
        RECT 35.110 104.235 35.390 105.185 ;
        RECT 35.560 105.095 35.785 105.225 ;
        RECT 35.560 103.990 35.730 105.095 ;
        RECT 35.955 104.945 36.480 105.165 ;
        RECT 35.900 104.180 36.140 104.775 ;
        RECT 36.310 104.245 36.480 104.945 ;
        RECT 36.650 104.585 36.820 105.365 ;
        RECT 37.140 105.315 37.510 105.815 ;
        RECT 37.690 105.365 38.095 105.535 ;
        RECT 38.265 105.365 39.050 105.535 ;
        RECT 37.690 105.135 37.860 105.365 ;
        RECT 37.030 104.835 37.860 105.135 ;
        RECT 38.245 104.865 38.710 105.195 ;
        RECT 37.030 104.805 37.230 104.835 ;
        RECT 37.350 104.585 37.520 104.655 ;
        RECT 36.650 104.415 37.520 104.585 ;
        RECT 37.010 104.325 37.520 104.415 ;
        RECT 35.560 103.860 35.865 103.990 ;
        RECT 36.310 103.880 36.840 104.245 ;
        RECT 35.180 103.265 35.445 103.725 ;
        RECT 35.615 103.435 35.865 103.860 ;
        RECT 37.010 103.710 37.180 104.325 ;
        RECT 36.075 103.540 37.180 103.710 ;
        RECT 37.350 103.265 37.520 104.065 ;
        RECT 37.690 103.765 37.860 104.835 ;
        RECT 38.030 103.935 38.220 104.655 ;
        RECT 38.390 103.905 38.710 104.865 ;
        RECT 38.880 104.905 39.050 105.365 ;
        RECT 39.325 105.285 39.535 105.815 ;
        RECT 39.795 105.075 40.125 105.600 ;
        RECT 40.295 105.205 40.465 105.815 ;
        RECT 40.635 105.160 40.965 105.595 ;
        RECT 41.275 105.265 41.445 105.555 ;
        RECT 41.615 105.435 41.945 105.815 ;
        RECT 40.635 105.075 41.015 105.160 ;
        RECT 41.275 105.095 41.940 105.265 ;
        RECT 39.925 104.905 40.125 105.075 ;
        RECT 40.790 105.035 41.015 105.075 ;
        RECT 38.880 104.575 39.755 104.905 ;
        RECT 39.925 104.575 40.675 104.905 ;
        RECT 37.690 103.435 37.940 103.765 ;
        RECT 38.880 103.735 39.050 104.575 ;
        RECT 39.925 104.370 40.115 104.575 ;
        RECT 40.845 104.455 41.015 105.035 ;
        RECT 40.800 104.405 41.015 104.455 ;
        RECT 39.220 103.995 40.115 104.370 ;
        RECT 40.625 104.325 41.015 104.405 ;
        RECT 38.165 103.565 39.050 103.735 ;
        RECT 39.230 103.265 39.545 103.765 ;
        RECT 39.775 103.435 40.115 103.995 ;
        RECT 40.285 103.265 40.455 104.275 ;
        RECT 40.625 103.480 40.955 104.325 ;
        RECT 41.190 104.275 41.540 104.925 ;
        RECT 41.710 104.105 41.940 105.095 ;
        RECT 41.275 103.935 41.940 104.105 ;
        RECT 41.275 103.435 41.445 103.935 ;
        RECT 41.615 103.265 41.945 103.765 ;
        RECT 42.115 103.435 42.300 105.555 ;
        RECT 42.555 105.355 42.805 105.815 ;
        RECT 42.975 105.365 43.310 105.535 ;
        RECT 43.505 105.365 44.180 105.535 ;
        RECT 42.975 105.225 43.145 105.365 ;
        RECT 42.470 104.235 42.750 105.185 ;
        RECT 42.920 105.095 43.145 105.225 ;
        RECT 42.920 103.990 43.090 105.095 ;
        RECT 43.315 104.945 43.840 105.165 ;
        RECT 43.260 104.180 43.500 104.775 ;
        RECT 43.670 104.245 43.840 104.945 ;
        RECT 44.010 104.585 44.180 105.365 ;
        RECT 44.500 105.315 44.870 105.815 ;
        RECT 45.050 105.365 45.455 105.535 ;
        RECT 45.625 105.365 46.410 105.535 ;
        RECT 45.050 105.135 45.220 105.365 ;
        RECT 44.390 104.835 45.220 105.135 ;
        RECT 45.605 104.865 46.070 105.195 ;
        RECT 44.390 104.805 44.590 104.835 ;
        RECT 44.710 104.585 44.880 104.655 ;
        RECT 44.010 104.415 44.880 104.585 ;
        RECT 44.370 104.325 44.880 104.415 ;
        RECT 42.920 103.860 43.225 103.990 ;
        RECT 43.670 103.880 44.200 104.245 ;
        RECT 42.540 103.265 42.805 103.725 ;
        RECT 42.975 103.435 43.225 103.860 ;
        RECT 44.370 103.710 44.540 104.325 ;
        RECT 43.435 103.540 44.540 103.710 ;
        RECT 44.710 103.265 44.880 104.065 ;
        RECT 45.050 103.765 45.220 104.835 ;
        RECT 45.390 103.935 45.580 104.655 ;
        RECT 45.750 103.905 46.070 104.865 ;
        RECT 46.240 104.905 46.410 105.365 ;
        RECT 46.685 105.285 46.895 105.815 ;
        RECT 47.155 105.075 47.485 105.600 ;
        RECT 47.655 105.205 47.825 105.815 ;
        RECT 47.995 105.160 48.325 105.595 ;
        RECT 47.995 105.075 48.375 105.160 ;
        RECT 48.545 105.090 48.835 105.815 ;
        RECT 47.285 104.905 47.485 105.075 ;
        RECT 48.150 105.035 48.375 105.075 ;
        RECT 46.240 104.575 47.115 104.905 ;
        RECT 47.285 104.575 48.035 104.905 ;
        RECT 45.050 103.435 45.300 103.765 ;
        RECT 46.240 103.735 46.410 104.575 ;
        RECT 47.285 104.370 47.475 104.575 ;
        RECT 48.205 104.455 48.375 105.035 ;
        RECT 49.005 105.045 50.675 105.815 ;
        RECT 50.960 105.185 51.245 105.645 ;
        RECT 51.415 105.355 51.685 105.815 ;
        RECT 49.005 104.525 49.755 105.045 ;
        RECT 50.960 105.015 51.915 105.185 ;
        RECT 48.160 104.405 48.375 104.455 ;
        RECT 46.580 103.995 47.475 104.370 ;
        RECT 47.985 104.325 48.375 104.405 ;
        RECT 45.525 103.565 46.410 103.735 ;
        RECT 46.590 103.265 46.905 103.765 ;
        RECT 47.135 103.435 47.475 103.995 ;
        RECT 47.645 103.265 47.815 104.275 ;
        RECT 47.985 103.480 48.315 104.325 ;
        RECT 48.545 103.265 48.835 104.430 ;
        RECT 49.925 104.355 50.675 104.875 ;
        RECT 49.005 103.265 50.675 104.355 ;
        RECT 50.845 104.285 51.535 104.845 ;
        RECT 51.705 104.115 51.915 105.015 ;
        RECT 50.960 103.895 51.915 104.115 ;
        RECT 52.085 104.845 52.485 105.645 ;
        RECT 52.675 105.185 52.955 105.645 ;
        RECT 53.475 105.355 53.800 105.815 ;
        RECT 52.675 105.015 53.800 105.185 ;
        RECT 53.970 105.075 54.355 105.645 ;
        RECT 53.350 104.905 53.800 105.015 ;
        RECT 52.085 104.285 53.180 104.845 ;
        RECT 53.350 104.575 53.905 104.905 ;
        RECT 50.960 103.435 51.245 103.895 ;
        RECT 51.415 103.265 51.685 103.725 ;
        RECT 52.085 103.435 52.485 104.285 ;
        RECT 53.350 104.115 53.800 104.575 ;
        RECT 54.075 104.405 54.355 105.075 ;
        RECT 54.525 105.015 54.835 105.815 ;
        RECT 55.040 105.015 55.735 105.645 ;
        RECT 54.535 104.575 54.870 104.845 ;
        RECT 55.040 104.415 55.210 105.015 ;
        RECT 55.965 104.995 56.175 105.815 ;
        RECT 56.345 105.015 56.675 105.645 ;
        RECT 55.380 104.575 55.715 104.825 ;
        RECT 56.345 104.415 56.595 105.015 ;
        RECT 56.845 104.995 57.075 105.815 ;
        RECT 57.285 105.075 57.670 105.645 ;
        RECT 57.840 105.355 58.165 105.815 ;
        RECT 58.685 105.185 58.965 105.645 ;
        RECT 56.765 104.575 57.095 104.825 ;
        RECT 52.675 103.895 53.800 104.115 ;
        RECT 52.675 103.435 52.955 103.895 ;
        RECT 53.475 103.265 53.800 103.725 ;
        RECT 53.970 103.435 54.355 104.405 ;
        RECT 54.525 103.265 54.805 104.405 ;
        RECT 54.975 103.435 55.305 104.415 ;
        RECT 55.475 103.265 55.735 104.405 ;
        RECT 55.965 103.265 56.175 104.405 ;
        RECT 56.345 103.435 56.675 104.415 ;
        RECT 57.285 104.405 57.565 105.075 ;
        RECT 57.840 105.015 58.965 105.185 ;
        RECT 57.840 104.905 58.290 105.015 ;
        RECT 57.735 104.575 58.290 104.905 ;
        RECT 59.155 104.845 59.555 105.645 ;
        RECT 59.955 105.355 60.225 105.815 ;
        RECT 60.395 105.185 60.680 105.645 ;
        RECT 56.845 103.265 57.075 104.405 ;
        RECT 57.285 103.435 57.670 104.405 ;
        RECT 57.840 104.115 58.290 104.575 ;
        RECT 58.460 104.285 59.555 104.845 ;
        RECT 57.840 103.895 58.965 104.115 ;
        RECT 57.840 103.265 58.165 103.725 ;
        RECT 58.685 103.435 58.965 103.895 ;
        RECT 59.155 103.435 59.555 104.285 ;
        RECT 59.725 105.015 60.680 105.185 ;
        RECT 59.725 104.115 59.935 105.015 ;
        RECT 60.105 104.285 60.795 104.845 ;
        RECT 61.890 104.215 62.225 105.635 ;
        RECT 62.405 105.445 63.150 105.815 ;
        RECT 63.715 105.275 63.970 105.635 ;
        RECT 64.150 105.445 64.480 105.815 ;
        RECT 64.660 105.275 64.885 105.635 ;
        RECT 62.400 105.085 64.885 105.275 ;
        RECT 62.400 104.395 62.625 105.085 ;
        RECT 65.575 105.005 65.845 105.815 ;
        RECT 66.015 105.005 66.345 105.645 ;
        RECT 66.515 105.005 66.755 105.815 ;
        RECT 67.035 105.265 67.205 105.555 ;
        RECT 67.375 105.435 67.705 105.815 ;
        RECT 67.035 105.095 67.700 105.265 ;
        RECT 62.825 104.575 63.105 104.905 ;
        RECT 63.285 104.575 63.860 104.905 ;
        RECT 64.040 104.575 64.475 104.905 ;
        RECT 64.655 104.575 64.925 104.905 ;
        RECT 65.565 104.575 65.915 104.825 ;
        RECT 66.085 104.405 66.255 105.005 ;
        RECT 66.425 104.575 66.775 104.825 ;
        RECT 62.400 104.215 64.895 104.395 ;
        RECT 59.725 103.895 60.680 104.115 ;
        RECT 59.955 103.265 60.225 103.725 ;
        RECT 60.395 103.435 60.680 103.895 ;
        RECT 61.890 103.445 62.155 104.215 ;
        RECT 62.325 103.265 62.655 103.985 ;
        RECT 62.845 103.805 64.035 104.035 ;
        RECT 62.845 103.445 63.105 103.805 ;
        RECT 63.275 103.265 63.605 103.635 ;
        RECT 63.775 103.445 64.035 103.805 ;
        RECT 64.605 103.445 64.895 104.215 ;
        RECT 65.575 103.265 65.905 104.405 ;
        RECT 66.085 104.235 66.765 104.405 ;
        RECT 66.950 104.275 67.300 104.925 ;
        RECT 66.435 103.450 66.765 104.235 ;
        RECT 67.470 104.105 67.700 105.095 ;
        RECT 67.035 103.935 67.700 104.105 ;
        RECT 67.035 103.435 67.205 103.935 ;
        RECT 67.375 103.265 67.705 103.765 ;
        RECT 67.875 103.435 68.060 105.555 ;
        RECT 68.315 105.355 68.565 105.815 ;
        RECT 68.735 105.365 69.070 105.535 ;
        RECT 69.265 105.365 69.940 105.535 ;
        RECT 68.735 105.225 68.905 105.365 ;
        RECT 68.230 104.235 68.510 105.185 ;
        RECT 68.680 105.095 68.905 105.225 ;
        RECT 68.680 103.990 68.850 105.095 ;
        RECT 69.075 104.945 69.600 105.165 ;
        RECT 69.020 104.180 69.260 104.775 ;
        RECT 69.430 104.245 69.600 104.945 ;
        RECT 69.770 104.585 69.940 105.365 ;
        RECT 70.260 105.315 70.630 105.815 ;
        RECT 70.810 105.365 71.215 105.535 ;
        RECT 71.385 105.365 72.170 105.535 ;
        RECT 70.810 105.135 70.980 105.365 ;
        RECT 70.150 104.835 70.980 105.135 ;
        RECT 71.365 104.865 71.830 105.195 ;
        RECT 70.150 104.805 70.350 104.835 ;
        RECT 70.470 104.585 70.640 104.655 ;
        RECT 69.770 104.415 70.640 104.585 ;
        RECT 70.130 104.325 70.640 104.415 ;
        RECT 68.680 103.860 68.985 103.990 ;
        RECT 69.430 103.880 69.960 104.245 ;
        RECT 68.300 103.265 68.565 103.725 ;
        RECT 68.735 103.435 68.985 103.860 ;
        RECT 70.130 103.710 70.300 104.325 ;
        RECT 69.195 103.540 70.300 103.710 ;
        RECT 70.470 103.265 70.640 104.065 ;
        RECT 70.810 103.765 70.980 104.835 ;
        RECT 71.150 103.935 71.340 104.655 ;
        RECT 71.510 103.905 71.830 104.865 ;
        RECT 72.000 104.905 72.170 105.365 ;
        RECT 72.445 105.285 72.655 105.815 ;
        RECT 72.915 105.075 73.245 105.600 ;
        RECT 73.415 105.205 73.585 105.815 ;
        RECT 73.755 105.160 74.085 105.595 ;
        RECT 73.755 105.075 74.135 105.160 ;
        RECT 74.305 105.090 74.595 105.815 ;
        RECT 74.765 105.165 75.025 105.645 ;
        RECT 75.195 105.275 75.445 105.815 ;
        RECT 73.045 104.905 73.245 105.075 ;
        RECT 73.910 105.035 74.135 105.075 ;
        RECT 72.000 104.575 72.875 104.905 ;
        RECT 73.045 104.575 73.795 104.905 ;
        RECT 70.810 103.435 71.060 103.765 ;
        RECT 72.000 103.735 72.170 104.575 ;
        RECT 73.045 104.370 73.235 104.575 ;
        RECT 73.965 104.455 74.135 105.035 ;
        RECT 73.920 104.405 74.135 104.455 ;
        RECT 72.340 103.995 73.235 104.370 ;
        RECT 73.745 104.325 74.135 104.405 ;
        RECT 71.285 103.565 72.170 103.735 ;
        RECT 72.350 103.265 72.665 103.765 ;
        RECT 72.895 103.435 73.235 103.995 ;
        RECT 73.405 103.265 73.575 104.275 ;
        RECT 73.745 103.480 74.075 104.325 ;
        RECT 74.305 103.265 74.595 104.430 ;
        RECT 74.765 104.135 74.935 105.165 ;
        RECT 75.615 105.135 75.835 105.595 ;
        RECT 75.585 105.110 75.835 105.135 ;
        RECT 75.105 104.515 75.335 104.910 ;
        RECT 75.505 104.685 75.835 105.110 ;
        RECT 76.005 105.435 76.895 105.605 ;
        RECT 76.005 104.710 76.175 105.435 ;
        RECT 76.345 104.880 76.895 105.265 ;
        RECT 76.005 104.640 76.895 104.710 ;
        RECT 76.000 104.615 76.895 104.640 ;
        RECT 75.990 104.600 76.895 104.615 ;
        RECT 75.985 104.585 76.895 104.600 ;
        RECT 75.975 104.580 76.895 104.585 ;
        RECT 75.970 104.570 76.895 104.580 ;
        RECT 75.965 104.560 76.895 104.570 ;
        RECT 75.955 104.555 76.895 104.560 ;
        RECT 75.945 104.545 76.895 104.555 ;
        RECT 75.935 104.540 76.895 104.545 ;
        RECT 75.935 104.535 76.270 104.540 ;
        RECT 75.920 104.530 76.270 104.535 ;
        RECT 75.905 104.520 76.270 104.530 ;
        RECT 75.880 104.515 76.270 104.520 ;
        RECT 75.105 104.510 76.270 104.515 ;
        RECT 75.105 104.475 76.240 104.510 ;
        RECT 75.105 104.450 76.205 104.475 ;
        RECT 75.105 104.420 76.175 104.450 ;
        RECT 75.105 104.390 76.155 104.420 ;
        RECT 75.105 104.360 76.135 104.390 ;
        RECT 75.105 104.350 76.065 104.360 ;
        RECT 75.105 104.340 76.040 104.350 ;
        RECT 75.105 104.325 76.020 104.340 ;
        RECT 75.105 104.310 76.000 104.325 ;
        RECT 75.210 104.300 75.995 104.310 ;
        RECT 75.210 104.265 75.980 104.300 ;
        RECT 74.765 103.435 75.040 104.135 ;
        RECT 75.210 104.015 75.965 104.265 ;
        RECT 76.135 103.945 76.465 104.190 ;
        RECT 76.635 104.090 76.895 104.540 ;
        RECT 76.280 103.920 76.465 103.945 ;
        RECT 76.280 103.820 76.895 103.920 ;
        RECT 75.210 103.265 75.465 103.810 ;
        RECT 75.635 103.435 76.115 103.775 ;
        RECT 76.290 103.265 76.895 103.820 ;
        RECT 77.535 103.445 77.795 105.635 ;
        RECT 78.055 105.445 78.725 105.815 ;
        RECT 78.905 105.265 79.215 105.635 ;
        RECT 77.985 105.065 79.215 105.265 ;
        RECT 77.985 104.395 78.275 105.065 ;
        RECT 79.395 104.885 79.625 105.525 ;
        RECT 79.805 105.085 80.095 105.815 ;
        RECT 80.285 105.165 80.545 105.645 ;
        RECT 80.715 105.275 80.965 105.815 ;
        RECT 78.455 104.575 78.920 104.885 ;
        RECT 79.100 104.575 79.625 104.885 ;
        RECT 79.805 104.575 80.105 104.905 ;
        RECT 77.985 104.175 78.755 104.395 ;
        RECT 77.965 103.265 78.305 103.995 ;
        RECT 78.485 103.445 78.755 104.175 ;
        RECT 78.935 104.155 80.095 104.395 ;
        RECT 78.935 103.445 79.165 104.155 ;
        RECT 79.335 103.265 79.665 103.975 ;
        RECT 79.835 103.445 80.095 104.155 ;
        RECT 80.285 104.135 80.455 105.165 ;
        RECT 81.135 105.110 81.355 105.595 ;
        RECT 80.625 104.515 80.855 104.910 ;
        RECT 81.025 104.685 81.355 105.110 ;
        RECT 81.525 105.435 82.415 105.605 ;
        RECT 81.525 104.710 81.695 105.435 ;
        RECT 81.865 104.880 82.415 105.265 ;
        RECT 82.585 105.045 84.255 105.815 ;
        RECT 81.525 104.640 82.415 104.710 ;
        RECT 81.520 104.615 82.415 104.640 ;
        RECT 81.510 104.600 82.415 104.615 ;
        RECT 81.505 104.585 82.415 104.600 ;
        RECT 81.495 104.580 82.415 104.585 ;
        RECT 81.490 104.570 82.415 104.580 ;
        RECT 81.485 104.560 82.415 104.570 ;
        RECT 81.475 104.555 82.415 104.560 ;
        RECT 81.465 104.545 82.415 104.555 ;
        RECT 81.455 104.540 82.415 104.545 ;
        RECT 81.455 104.535 81.790 104.540 ;
        RECT 81.440 104.530 81.790 104.535 ;
        RECT 81.425 104.520 81.790 104.530 ;
        RECT 81.400 104.515 81.790 104.520 ;
        RECT 80.625 104.510 81.790 104.515 ;
        RECT 80.625 104.475 81.760 104.510 ;
        RECT 80.625 104.450 81.725 104.475 ;
        RECT 80.625 104.420 81.695 104.450 ;
        RECT 80.625 104.390 81.675 104.420 ;
        RECT 80.625 104.360 81.655 104.390 ;
        RECT 80.625 104.350 81.585 104.360 ;
        RECT 80.625 104.340 81.560 104.350 ;
        RECT 80.625 104.325 81.540 104.340 ;
        RECT 80.625 104.310 81.520 104.325 ;
        RECT 80.730 104.300 81.515 104.310 ;
        RECT 80.730 104.265 81.500 104.300 ;
        RECT 80.285 103.435 80.560 104.135 ;
        RECT 80.730 104.015 81.485 104.265 ;
        RECT 81.655 103.945 81.985 104.190 ;
        RECT 82.155 104.090 82.415 104.540 ;
        RECT 82.585 104.525 83.335 105.045 ;
        RECT 84.905 105.005 85.145 105.815 ;
        RECT 85.315 105.005 85.645 105.645 ;
        RECT 85.815 105.005 86.085 105.815 ;
        RECT 86.265 105.270 91.610 105.815 ;
        RECT 83.505 104.355 84.255 104.875 ;
        RECT 84.885 104.575 85.235 104.825 ;
        RECT 85.405 104.405 85.575 105.005 ;
        RECT 85.745 104.575 86.095 104.825 ;
        RECT 87.850 104.440 88.190 105.270 ;
        RECT 81.800 103.920 81.985 103.945 ;
        RECT 81.800 103.820 82.415 103.920 ;
        RECT 80.730 103.265 80.985 103.810 ;
        RECT 81.155 103.435 81.635 103.775 ;
        RECT 81.810 103.265 82.415 103.820 ;
        RECT 82.585 103.265 84.255 104.355 ;
        RECT 84.895 104.235 85.575 104.405 ;
        RECT 84.895 103.450 85.225 104.235 ;
        RECT 85.755 103.265 86.085 104.405 ;
        RECT 89.670 103.700 90.020 104.950 ;
        RECT 92.250 104.215 92.585 105.635 ;
        RECT 92.765 105.445 93.510 105.815 ;
        RECT 94.075 105.275 94.330 105.635 ;
        RECT 94.510 105.445 94.840 105.815 ;
        RECT 95.020 105.275 95.245 105.635 ;
        RECT 92.760 105.085 95.245 105.275 ;
        RECT 92.760 104.395 92.985 105.085 ;
        RECT 95.465 105.075 95.850 105.645 ;
        RECT 96.020 105.355 96.345 105.815 ;
        RECT 96.865 105.185 97.145 105.645 ;
        RECT 93.185 104.575 93.465 104.905 ;
        RECT 93.645 104.575 94.220 104.905 ;
        RECT 94.400 104.575 94.835 104.905 ;
        RECT 95.015 104.575 95.285 104.905 ;
        RECT 95.465 104.405 95.745 105.075 ;
        RECT 96.020 105.015 97.145 105.185 ;
        RECT 96.020 104.905 96.470 105.015 ;
        RECT 95.915 104.575 96.470 104.905 ;
        RECT 97.335 104.845 97.735 105.645 ;
        RECT 98.135 105.355 98.405 105.815 ;
        RECT 98.575 105.185 98.860 105.645 ;
        RECT 92.760 104.215 95.255 104.395 ;
        RECT 86.265 103.265 91.610 103.700 ;
        RECT 92.250 103.445 92.515 104.215 ;
        RECT 92.685 103.265 93.015 103.985 ;
        RECT 93.205 103.805 94.395 104.035 ;
        RECT 93.205 103.445 93.465 103.805 ;
        RECT 93.635 103.265 93.965 103.635 ;
        RECT 94.135 103.445 94.395 103.805 ;
        RECT 94.965 103.445 95.255 104.215 ;
        RECT 95.465 103.435 95.850 104.405 ;
        RECT 96.020 104.115 96.470 104.575 ;
        RECT 96.640 104.285 97.735 104.845 ;
        RECT 96.020 103.895 97.145 104.115 ;
        RECT 96.020 103.265 96.345 103.725 ;
        RECT 96.865 103.435 97.145 103.895 ;
        RECT 97.335 103.435 97.735 104.285 ;
        RECT 97.905 105.015 98.860 105.185 ;
        RECT 100.065 105.090 100.355 105.815 ;
        RECT 97.905 104.115 98.115 105.015 ;
        RECT 100.545 105.005 100.785 105.815 ;
        RECT 100.955 105.005 101.285 105.645 ;
        RECT 101.455 105.005 101.725 105.815 ;
        RECT 101.955 105.160 102.285 105.595 ;
        RECT 102.455 105.205 102.625 105.815 ;
        RECT 101.905 105.075 102.285 105.160 ;
        RECT 102.795 105.075 103.125 105.600 ;
        RECT 103.385 105.285 103.595 105.815 ;
        RECT 103.870 105.365 104.655 105.535 ;
        RECT 104.825 105.365 105.230 105.535 ;
        RECT 101.905 105.035 102.130 105.075 ;
        RECT 98.285 104.285 98.975 104.845 ;
        RECT 100.525 104.575 100.875 104.825 ;
        RECT 97.905 103.895 98.860 104.115 ;
        RECT 98.135 103.265 98.405 103.725 ;
        RECT 98.575 103.435 98.860 103.895 ;
        RECT 100.065 103.265 100.355 104.430 ;
        RECT 101.045 104.405 101.215 105.005 ;
        RECT 101.385 104.575 101.735 104.825 ;
        RECT 101.905 104.455 102.075 105.035 ;
        RECT 102.795 104.905 102.995 105.075 ;
        RECT 103.870 104.905 104.040 105.365 ;
        RECT 102.245 104.575 102.995 104.905 ;
        RECT 103.165 104.575 104.040 104.905 ;
        RECT 101.905 104.405 102.120 104.455 ;
        RECT 100.535 104.235 101.215 104.405 ;
        RECT 100.535 103.450 100.865 104.235 ;
        RECT 101.395 103.265 101.725 104.405 ;
        RECT 101.905 104.325 102.295 104.405 ;
        RECT 101.965 103.480 102.295 104.325 ;
        RECT 102.805 104.370 102.995 104.575 ;
        RECT 102.465 103.265 102.635 104.275 ;
        RECT 102.805 103.995 103.700 104.370 ;
        RECT 102.805 103.435 103.145 103.995 ;
        RECT 103.375 103.265 103.690 103.765 ;
        RECT 103.870 103.735 104.040 104.575 ;
        RECT 104.210 104.865 104.675 105.195 ;
        RECT 105.060 105.135 105.230 105.365 ;
        RECT 105.410 105.315 105.780 105.815 ;
        RECT 106.100 105.365 106.775 105.535 ;
        RECT 106.970 105.365 107.305 105.535 ;
        RECT 104.210 103.905 104.530 104.865 ;
        RECT 105.060 104.835 105.890 105.135 ;
        RECT 104.700 103.935 104.890 104.655 ;
        RECT 105.060 103.765 105.230 104.835 ;
        RECT 105.690 104.805 105.890 104.835 ;
        RECT 105.400 104.585 105.570 104.655 ;
        RECT 106.100 104.585 106.270 105.365 ;
        RECT 107.135 105.225 107.305 105.365 ;
        RECT 107.475 105.355 107.725 105.815 ;
        RECT 105.400 104.415 106.270 104.585 ;
        RECT 106.440 104.945 106.965 105.165 ;
        RECT 107.135 105.095 107.360 105.225 ;
        RECT 105.400 104.325 105.910 104.415 ;
        RECT 103.870 103.565 104.755 103.735 ;
        RECT 104.980 103.435 105.230 103.765 ;
        RECT 105.400 103.265 105.570 104.065 ;
        RECT 105.740 103.710 105.910 104.325 ;
        RECT 106.440 104.245 106.610 104.945 ;
        RECT 106.080 103.880 106.610 104.245 ;
        RECT 106.780 104.180 107.020 104.775 ;
        RECT 107.190 103.990 107.360 105.095 ;
        RECT 107.530 104.235 107.810 105.185 ;
        RECT 107.055 103.860 107.360 103.990 ;
        RECT 105.740 103.540 106.845 103.710 ;
        RECT 107.055 103.435 107.305 103.860 ;
        RECT 107.475 103.265 107.740 103.725 ;
        RECT 107.980 103.435 108.165 105.555 ;
        RECT 108.335 105.435 108.665 105.815 ;
        RECT 108.835 105.265 109.005 105.555 ;
        RECT 108.340 105.095 109.005 105.265 ;
        RECT 108.340 104.105 108.570 105.095 ;
        RECT 110.205 105.085 110.495 105.815 ;
        RECT 108.740 104.275 109.090 104.925 ;
        RECT 110.195 104.575 110.495 104.905 ;
        RECT 110.675 104.885 110.905 105.525 ;
        RECT 111.085 105.265 111.395 105.635 ;
        RECT 111.575 105.445 112.245 105.815 ;
        RECT 111.085 105.065 112.315 105.265 ;
        RECT 110.675 104.575 111.200 104.885 ;
        RECT 111.380 104.575 111.845 104.885 ;
        RECT 112.025 104.395 112.315 105.065 ;
        RECT 110.205 104.155 111.365 104.395 ;
        RECT 108.340 103.935 109.005 104.105 ;
        RECT 108.335 103.265 108.665 103.765 ;
        RECT 108.835 103.435 109.005 103.935 ;
        RECT 110.205 103.445 110.465 104.155 ;
        RECT 110.635 103.265 110.965 103.975 ;
        RECT 111.135 103.445 111.365 104.155 ;
        RECT 111.545 104.175 112.315 104.395 ;
        RECT 111.545 103.445 111.815 104.175 ;
        RECT 111.995 103.265 112.335 103.995 ;
        RECT 112.505 103.445 112.765 105.635 ;
        RECT 112.945 105.165 113.205 105.645 ;
        RECT 113.375 105.275 113.625 105.815 ;
        RECT 112.945 104.135 113.115 105.165 ;
        RECT 113.795 105.110 114.015 105.595 ;
        RECT 113.285 104.515 113.515 104.910 ;
        RECT 113.685 104.685 114.015 105.110 ;
        RECT 114.185 105.435 115.075 105.605 ;
        RECT 114.185 104.710 114.355 105.435 ;
        RECT 114.525 104.880 115.075 105.265 ;
        RECT 115.245 105.045 116.915 105.815 ;
        RECT 117.085 105.075 117.470 105.645 ;
        RECT 117.640 105.355 117.965 105.815 ;
        RECT 118.485 105.185 118.765 105.645 ;
        RECT 114.185 104.640 115.075 104.710 ;
        RECT 114.180 104.615 115.075 104.640 ;
        RECT 114.170 104.600 115.075 104.615 ;
        RECT 114.165 104.585 115.075 104.600 ;
        RECT 114.155 104.580 115.075 104.585 ;
        RECT 114.150 104.570 115.075 104.580 ;
        RECT 114.145 104.560 115.075 104.570 ;
        RECT 114.135 104.555 115.075 104.560 ;
        RECT 114.125 104.545 115.075 104.555 ;
        RECT 114.115 104.540 115.075 104.545 ;
        RECT 114.115 104.535 114.450 104.540 ;
        RECT 114.100 104.530 114.450 104.535 ;
        RECT 114.085 104.520 114.450 104.530 ;
        RECT 114.060 104.515 114.450 104.520 ;
        RECT 113.285 104.510 114.450 104.515 ;
        RECT 113.285 104.475 114.420 104.510 ;
        RECT 113.285 104.450 114.385 104.475 ;
        RECT 113.285 104.420 114.355 104.450 ;
        RECT 113.285 104.390 114.335 104.420 ;
        RECT 113.285 104.360 114.315 104.390 ;
        RECT 113.285 104.350 114.245 104.360 ;
        RECT 113.285 104.340 114.220 104.350 ;
        RECT 113.285 104.325 114.200 104.340 ;
        RECT 113.285 104.310 114.180 104.325 ;
        RECT 113.390 104.300 114.175 104.310 ;
        RECT 113.390 104.265 114.160 104.300 ;
        RECT 112.945 103.435 113.220 104.135 ;
        RECT 113.390 104.015 114.145 104.265 ;
        RECT 114.315 103.945 114.645 104.190 ;
        RECT 114.815 104.090 115.075 104.540 ;
        RECT 115.245 104.525 115.995 105.045 ;
        RECT 116.165 104.355 116.915 104.875 ;
        RECT 114.460 103.920 114.645 103.945 ;
        RECT 114.460 103.820 115.075 103.920 ;
        RECT 113.390 103.265 113.645 103.810 ;
        RECT 113.815 103.435 114.295 103.775 ;
        RECT 114.470 103.265 115.075 103.820 ;
        RECT 115.245 103.265 116.915 104.355 ;
        RECT 117.085 104.405 117.365 105.075 ;
        RECT 117.640 105.015 118.765 105.185 ;
        RECT 117.640 104.905 118.090 105.015 ;
        RECT 117.535 104.575 118.090 104.905 ;
        RECT 118.955 104.845 119.355 105.645 ;
        RECT 119.755 105.355 120.025 105.815 ;
        RECT 120.195 105.185 120.480 105.645 ;
        RECT 117.085 103.435 117.470 104.405 ;
        RECT 117.640 104.115 118.090 104.575 ;
        RECT 118.260 104.285 119.355 104.845 ;
        RECT 117.640 103.895 118.765 104.115 ;
        RECT 117.640 103.265 117.965 103.725 ;
        RECT 118.485 103.435 118.765 103.895 ;
        RECT 118.955 103.435 119.355 104.285 ;
        RECT 119.525 105.015 120.480 105.185 ;
        RECT 120.765 105.045 124.275 105.815 ;
        RECT 124.445 105.065 125.655 105.815 ;
        RECT 125.825 105.090 126.115 105.815 ;
        RECT 119.525 104.115 119.735 105.015 ;
        RECT 119.905 104.285 120.595 104.845 ;
        RECT 120.765 104.525 122.415 105.045 ;
        RECT 122.585 104.355 124.275 104.875 ;
        RECT 124.445 104.525 124.965 105.065 ;
        RECT 126.285 105.045 127.955 105.815 ;
        RECT 128.290 105.305 128.530 105.815 ;
        RECT 128.710 105.305 128.990 105.635 ;
        RECT 129.220 105.305 129.435 105.815 ;
        RECT 125.135 104.355 125.655 104.895 ;
        RECT 126.285 104.525 127.035 105.045 ;
        RECT 119.525 103.895 120.480 104.115 ;
        RECT 119.755 103.265 120.025 103.725 ;
        RECT 120.195 103.435 120.480 103.895 ;
        RECT 120.765 103.265 124.275 104.355 ;
        RECT 124.445 103.265 125.655 104.355 ;
        RECT 125.825 103.265 126.115 104.430 ;
        RECT 127.205 104.355 127.955 104.875 ;
        RECT 128.185 104.575 128.540 105.135 ;
        RECT 128.710 104.405 128.880 105.305 ;
        RECT 129.050 104.575 129.315 105.135 ;
        RECT 129.605 105.075 130.220 105.645 ;
        RECT 129.565 104.405 129.735 104.905 ;
        RECT 126.285 103.265 127.955 104.355 ;
        RECT 128.310 104.235 129.735 104.405 ;
        RECT 128.310 104.060 128.700 104.235 ;
        RECT 129.185 103.265 129.515 104.065 ;
        RECT 129.905 104.055 130.220 105.075 ;
        RECT 129.685 103.435 130.220 104.055 ;
        RECT 130.425 105.015 130.765 105.645 ;
        RECT 130.935 105.015 131.185 105.815 ;
        RECT 131.375 105.165 131.705 105.645 ;
        RECT 131.875 105.355 132.100 105.815 ;
        RECT 132.270 105.165 132.600 105.645 ;
        RECT 130.425 104.405 130.600 105.015 ;
        RECT 131.375 104.995 132.600 105.165 ;
        RECT 133.230 105.035 133.730 105.645 ;
        RECT 134.310 105.035 134.810 105.645 ;
        RECT 130.770 104.655 131.465 104.825 ;
        RECT 131.295 104.405 131.465 104.655 ;
        RECT 131.640 104.625 132.060 104.825 ;
        RECT 132.230 104.625 132.560 104.825 ;
        RECT 132.730 104.625 133.060 104.825 ;
        RECT 133.230 104.405 133.400 105.035 ;
        RECT 133.585 104.575 133.935 104.825 ;
        RECT 134.105 104.575 134.455 104.825 ;
        RECT 134.640 104.405 134.810 105.035 ;
        RECT 135.440 105.165 135.770 105.645 ;
        RECT 135.940 105.355 136.165 105.815 ;
        RECT 136.335 105.165 136.665 105.645 ;
        RECT 135.440 104.995 136.665 105.165 ;
        RECT 136.855 105.015 137.105 105.815 ;
        RECT 137.275 105.015 137.615 105.645 ;
        RECT 137.900 105.185 138.185 105.645 ;
        RECT 138.355 105.355 138.625 105.815 ;
        RECT 137.900 105.015 138.855 105.185 ;
        RECT 134.980 104.625 135.310 104.825 ;
        RECT 135.480 104.625 135.810 104.825 ;
        RECT 135.980 104.625 136.400 104.825 ;
        RECT 136.575 104.655 137.270 104.825 ;
        RECT 136.575 104.405 136.745 104.655 ;
        RECT 137.440 104.455 137.615 105.015 ;
        RECT 137.385 104.405 137.615 104.455 ;
        RECT 130.425 103.435 130.765 104.405 ;
        RECT 130.935 103.265 131.105 104.405 ;
        RECT 131.295 104.235 133.730 104.405 ;
        RECT 131.375 103.265 131.625 104.065 ;
        RECT 132.270 103.435 132.600 104.235 ;
        RECT 132.900 103.265 133.230 104.065 ;
        RECT 133.400 103.435 133.730 104.235 ;
        RECT 134.310 104.235 136.745 104.405 ;
        RECT 134.310 103.435 134.640 104.235 ;
        RECT 134.810 103.265 135.140 104.065 ;
        RECT 135.440 103.435 135.770 104.235 ;
        RECT 136.415 103.265 136.665 104.065 ;
        RECT 136.935 103.265 137.105 104.405 ;
        RECT 137.275 103.435 137.615 104.405 ;
        RECT 137.785 104.285 138.475 104.845 ;
        RECT 138.645 104.115 138.855 105.015 ;
        RECT 137.900 103.895 138.855 104.115 ;
        RECT 139.025 104.845 139.425 105.645 ;
        RECT 139.615 105.185 139.895 105.645 ;
        RECT 140.415 105.355 140.740 105.815 ;
        RECT 139.615 105.015 140.740 105.185 ;
        RECT 140.910 105.075 141.295 105.645 ;
        RECT 140.290 104.905 140.740 105.015 ;
        RECT 139.025 104.285 140.120 104.845 ;
        RECT 140.290 104.575 140.845 104.905 ;
        RECT 137.900 103.435 138.185 103.895 ;
        RECT 138.355 103.265 138.625 103.725 ;
        RECT 139.025 103.435 139.425 104.285 ;
        RECT 140.290 104.115 140.740 104.575 ;
        RECT 141.015 104.405 141.295 105.075 ;
        RECT 141.670 105.035 142.170 105.645 ;
        RECT 141.465 104.575 141.815 104.825 ;
        RECT 142.000 104.405 142.170 105.035 ;
        RECT 142.800 105.165 143.130 105.645 ;
        RECT 143.300 105.355 143.525 105.815 ;
        RECT 143.695 105.165 144.025 105.645 ;
        RECT 142.800 104.995 144.025 105.165 ;
        RECT 144.215 105.015 144.465 105.815 ;
        RECT 144.635 105.015 144.975 105.645 ;
        RECT 142.340 104.625 142.670 104.825 ;
        RECT 142.840 104.625 143.170 104.825 ;
        RECT 143.340 104.625 143.760 104.825 ;
        RECT 143.935 104.655 144.630 104.825 ;
        RECT 143.935 104.405 144.105 104.655 ;
        RECT 144.800 104.405 144.975 105.015 ;
        RECT 139.615 103.895 140.740 104.115 ;
        RECT 139.615 103.435 139.895 103.895 ;
        RECT 140.415 103.265 140.740 103.725 ;
        RECT 140.910 103.435 141.295 104.405 ;
        RECT 141.670 104.235 144.105 104.405 ;
        RECT 141.670 103.435 142.000 104.235 ;
        RECT 142.170 103.265 142.500 104.065 ;
        RECT 142.800 103.435 143.130 104.235 ;
        RECT 143.775 103.265 144.025 104.065 ;
        RECT 144.295 103.265 144.465 104.405 ;
        RECT 144.635 103.435 144.975 104.405 ;
        RECT 145.145 105.075 145.530 105.645 ;
        RECT 145.700 105.355 146.025 105.815 ;
        RECT 146.545 105.185 146.825 105.645 ;
        RECT 145.145 104.405 145.425 105.075 ;
        RECT 145.700 105.015 146.825 105.185 ;
        RECT 145.700 104.905 146.150 105.015 ;
        RECT 145.595 104.575 146.150 104.905 ;
        RECT 147.015 104.845 147.415 105.645 ;
        RECT 147.815 105.355 148.085 105.815 ;
        RECT 148.255 105.185 148.540 105.645 ;
        RECT 145.145 103.435 145.530 104.405 ;
        RECT 145.700 104.115 146.150 104.575 ;
        RECT 146.320 104.285 147.415 104.845 ;
        RECT 145.700 103.895 146.825 104.115 ;
        RECT 145.700 103.265 146.025 103.725 ;
        RECT 146.545 103.435 146.825 103.895 ;
        RECT 147.015 103.435 147.415 104.285 ;
        RECT 147.585 105.015 148.540 105.185 ;
        RECT 148.860 105.075 149.475 105.645 ;
        RECT 149.645 105.305 149.860 105.815 ;
        RECT 150.090 105.305 150.370 105.635 ;
        RECT 150.550 105.305 150.790 105.815 ;
        RECT 147.585 104.115 147.795 105.015 ;
        RECT 147.965 104.285 148.655 104.845 ;
        RECT 147.585 103.895 148.540 104.115 ;
        RECT 147.815 103.265 148.085 103.725 ;
        RECT 148.255 103.435 148.540 103.895 ;
        RECT 148.860 104.055 149.175 105.075 ;
        RECT 149.345 104.405 149.515 104.905 ;
        RECT 149.765 104.575 150.030 105.135 ;
        RECT 150.200 104.405 150.370 105.305 ;
        RECT 150.540 104.575 150.895 105.135 ;
        RECT 151.585 105.090 151.875 105.815 ;
        RECT 152.045 105.075 152.430 105.645 ;
        RECT 152.600 105.355 152.925 105.815 ;
        RECT 153.445 105.185 153.725 105.645 ;
        RECT 149.345 104.235 150.770 104.405 ;
        RECT 148.860 103.435 149.395 104.055 ;
        RECT 149.565 103.265 149.895 104.065 ;
        RECT 150.380 104.060 150.770 104.235 ;
        RECT 151.585 103.265 151.875 104.430 ;
        RECT 152.045 104.405 152.325 105.075 ;
        RECT 152.600 105.015 153.725 105.185 ;
        RECT 152.600 104.905 153.050 105.015 ;
        RECT 152.495 104.575 153.050 104.905 ;
        RECT 153.915 104.845 154.315 105.645 ;
        RECT 154.715 105.355 154.985 105.815 ;
        RECT 155.155 105.185 155.440 105.645 ;
        RECT 152.045 103.435 152.430 104.405 ;
        RECT 152.600 104.115 153.050 104.575 ;
        RECT 153.220 104.285 154.315 104.845 ;
        RECT 152.600 103.895 153.725 104.115 ;
        RECT 152.600 103.265 152.925 103.725 ;
        RECT 153.445 103.435 153.725 103.895 ;
        RECT 153.915 103.435 154.315 104.285 ;
        RECT 154.485 105.015 155.440 105.185 ;
        RECT 155.725 105.065 156.935 105.815 ;
        RECT 154.485 104.115 154.695 105.015 ;
        RECT 154.865 104.285 155.555 104.845 ;
        RECT 155.725 104.355 156.245 104.895 ;
        RECT 156.415 104.525 156.935 105.065 ;
        RECT 154.485 103.895 155.440 104.115 ;
        RECT 154.715 103.265 154.985 103.725 ;
        RECT 155.155 103.435 155.440 103.895 ;
        RECT 155.725 103.265 156.935 104.355 ;
        RECT 22.700 103.095 157.020 103.265 ;
        RECT 22.785 102.005 23.995 103.095 ;
        RECT 24.165 102.660 29.510 103.095 ;
        RECT 22.785 101.295 23.305 101.835 ;
        RECT 23.475 101.465 23.995 102.005 ;
        RECT 22.785 100.545 23.995 101.295 ;
        RECT 25.750 101.090 26.090 101.920 ;
        RECT 27.570 101.410 27.920 102.660 ;
        RECT 29.870 102.125 30.260 102.300 ;
        RECT 30.745 102.295 31.075 103.095 ;
        RECT 31.245 102.305 31.780 102.925 ;
        RECT 29.870 101.955 31.295 102.125 ;
        RECT 29.745 101.225 30.100 101.785 ;
        RECT 24.165 100.545 29.510 101.090 ;
        RECT 30.270 101.055 30.440 101.955 ;
        RECT 30.610 101.225 30.875 101.785 ;
        RECT 31.125 101.455 31.295 101.955 ;
        RECT 31.465 101.285 31.780 102.305 ;
        RECT 32.995 102.475 33.165 102.905 ;
        RECT 33.335 102.645 33.665 103.095 ;
        RECT 32.995 102.245 33.670 102.475 ;
        RECT 29.850 100.545 30.090 101.055 ;
        RECT 30.270 100.725 30.550 101.055 ;
        RECT 30.780 100.545 30.995 101.055 ;
        RECT 31.165 100.715 31.780 101.285 ;
        RECT 32.965 101.225 33.265 102.075 ;
        RECT 33.435 101.595 33.670 102.245 ;
        RECT 33.840 101.935 34.125 102.880 ;
        RECT 34.305 102.625 34.990 103.095 ;
        RECT 34.300 102.105 34.995 102.415 ;
        RECT 35.170 102.040 35.475 102.825 ;
        RECT 33.840 101.785 34.700 101.935 ;
        RECT 35.265 101.905 35.475 102.040 ;
        RECT 35.665 101.930 35.955 103.095 ;
        RECT 36.125 102.020 36.395 102.925 ;
        RECT 36.565 102.335 36.895 103.095 ;
        RECT 37.075 102.165 37.245 102.925 ;
        RECT 33.840 101.765 35.125 101.785 ;
        RECT 33.435 101.265 33.970 101.595 ;
        RECT 34.140 101.405 35.125 101.765 ;
        RECT 33.435 101.115 33.655 101.265 ;
        RECT 32.910 100.545 33.245 101.050 ;
        RECT 33.415 100.740 33.655 101.115 ;
        RECT 34.140 101.070 34.310 101.405 ;
        RECT 35.300 101.235 35.475 101.905 ;
        RECT 33.935 100.875 34.310 101.070 ;
        RECT 33.935 100.730 34.105 100.875 ;
        RECT 34.670 100.545 35.065 101.040 ;
        RECT 35.235 100.715 35.475 101.235 ;
        RECT 35.665 100.545 35.955 101.270 ;
        RECT 36.125 101.220 36.295 102.020 ;
        RECT 36.580 101.995 37.245 102.165 ;
        RECT 37.505 102.005 39.175 103.095 ;
        RECT 36.580 101.850 36.750 101.995 ;
        RECT 36.465 101.520 36.750 101.850 ;
        RECT 36.580 101.265 36.750 101.520 ;
        RECT 36.985 101.445 37.315 101.815 ;
        RECT 37.505 101.315 38.255 101.835 ;
        RECT 38.425 101.485 39.175 102.005 ;
        RECT 39.805 101.955 40.065 103.095 ;
        RECT 40.235 101.945 40.565 102.925 ;
        RECT 40.735 101.955 41.015 103.095 ;
        RECT 41.220 102.305 41.755 102.925 ;
        RECT 39.825 101.535 40.160 101.785 ;
        RECT 40.330 101.395 40.500 101.945 ;
        RECT 40.670 101.515 41.005 101.785 ;
        RECT 40.325 101.345 40.500 101.395 ;
        RECT 36.125 100.715 36.385 101.220 ;
        RECT 36.580 101.095 37.245 101.265 ;
        RECT 36.565 100.545 36.895 100.925 ;
        RECT 37.075 100.715 37.245 101.095 ;
        RECT 37.505 100.545 39.175 101.315 ;
        RECT 39.805 100.715 40.500 101.345 ;
        RECT 40.705 100.545 41.015 101.345 ;
        RECT 41.220 101.285 41.535 102.305 ;
        RECT 41.925 102.295 42.255 103.095 ;
        RECT 42.740 102.125 43.130 102.300 ;
        RECT 41.705 101.955 43.130 102.125 ;
        RECT 44.405 102.020 44.675 102.925 ;
        RECT 44.845 102.335 45.175 103.095 ;
        RECT 45.355 102.165 45.525 102.925 ;
        RECT 41.705 101.455 41.875 101.955 ;
        RECT 41.220 100.715 41.835 101.285 ;
        RECT 42.125 101.225 42.390 101.785 ;
        RECT 42.560 101.055 42.730 101.955 ;
        RECT 42.900 101.225 43.255 101.785 ;
        RECT 44.405 101.220 44.575 102.020 ;
        RECT 44.860 101.995 45.525 102.165 ;
        RECT 45.785 102.005 49.295 103.095 ;
        RECT 49.525 102.035 49.855 102.880 ;
        RECT 50.025 102.085 50.195 103.095 ;
        RECT 50.365 102.365 50.705 102.925 ;
        RECT 50.935 102.595 51.250 103.095 ;
        RECT 51.430 102.625 52.315 102.795 ;
        RECT 44.860 101.850 45.030 101.995 ;
        RECT 44.745 101.520 45.030 101.850 ;
        RECT 44.860 101.265 45.030 101.520 ;
        RECT 45.265 101.445 45.595 101.815 ;
        RECT 45.785 101.315 47.435 101.835 ;
        RECT 47.605 101.485 49.295 102.005 ;
        RECT 49.465 101.955 49.855 102.035 ;
        RECT 50.365 101.990 51.260 102.365 ;
        RECT 49.465 101.905 49.680 101.955 ;
        RECT 49.465 101.325 49.635 101.905 ;
        RECT 50.365 101.785 50.555 101.990 ;
        RECT 51.430 101.785 51.600 102.625 ;
        RECT 52.540 102.595 52.790 102.925 ;
        RECT 49.805 101.455 50.555 101.785 ;
        RECT 50.725 101.455 51.600 101.785 ;
        RECT 42.005 100.545 42.220 101.055 ;
        RECT 42.450 100.725 42.730 101.055 ;
        RECT 42.910 100.545 43.150 101.055 ;
        RECT 44.405 100.715 44.665 101.220 ;
        RECT 44.860 101.095 45.525 101.265 ;
        RECT 44.845 100.545 45.175 100.925 ;
        RECT 45.355 100.715 45.525 101.095 ;
        RECT 45.785 100.545 49.295 101.315 ;
        RECT 49.465 101.285 49.690 101.325 ;
        RECT 50.355 101.285 50.555 101.455 ;
        RECT 49.465 101.200 49.845 101.285 ;
        RECT 49.515 100.765 49.845 101.200 ;
        RECT 50.015 100.545 50.185 101.155 ;
        RECT 50.355 100.760 50.685 101.285 ;
        RECT 50.945 100.545 51.155 101.075 ;
        RECT 51.430 100.995 51.600 101.455 ;
        RECT 51.770 101.495 52.090 102.455 ;
        RECT 52.260 101.705 52.450 102.425 ;
        RECT 52.620 101.525 52.790 102.595 ;
        RECT 52.960 102.295 53.130 103.095 ;
        RECT 53.300 102.650 54.405 102.820 ;
        RECT 53.300 102.035 53.470 102.650 ;
        RECT 54.615 102.500 54.865 102.925 ;
        RECT 55.035 102.635 55.300 103.095 ;
        RECT 53.640 102.115 54.170 102.480 ;
        RECT 54.615 102.370 54.920 102.500 ;
        RECT 52.960 101.945 53.470 102.035 ;
        RECT 52.960 101.775 53.830 101.945 ;
        RECT 52.960 101.705 53.130 101.775 ;
        RECT 53.250 101.525 53.450 101.555 ;
        RECT 51.770 101.165 52.235 101.495 ;
        RECT 52.620 101.225 53.450 101.525 ;
        RECT 52.620 100.995 52.790 101.225 ;
        RECT 51.430 100.825 52.215 100.995 ;
        RECT 52.385 100.825 52.790 100.995 ;
        RECT 52.970 100.545 53.340 101.045 ;
        RECT 53.660 100.995 53.830 101.775 ;
        RECT 54.000 101.415 54.170 102.115 ;
        RECT 54.340 101.585 54.580 102.180 ;
        RECT 54.000 101.195 54.525 101.415 ;
        RECT 54.750 101.265 54.920 102.370 ;
        RECT 54.695 101.135 54.920 101.265 ;
        RECT 55.090 101.175 55.370 102.125 ;
        RECT 54.695 100.995 54.865 101.135 ;
        RECT 53.660 100.825 54.335 100.995 ;
        RECT 54.530 100.825 54.865 100.995 ;
        RECT 55.035 100.545 55.285 101.005 ;
        RECT 55.540 100.805 55.725 102.925 ;
        RECT 55.895 102.595 56.225 103.095 ;
        RECT 56.395 102.425 56.565 102.925 ;
        RECT 55.900 102.255 56.565 102.425 ;
        RECT 55.900 101.265 56.130 102.255 ;
        RECT 56.300 101.435 56.650 102.085 ;
        RECT 56.825 102.005 58.035 103.095 ;
        RECT 56.825 101.295 57.345 101.835 ;
        RECT 57.515 101.465 58.035 102.005 ;
        RECT 58.210 102.145 58.475 102.915 ;
        RECT 58.645 102.375 58.975 103.095 ;
        RECT 59.165 102.555 59.425 102.915 ;
        RECT 59.595 102.725 59.925 103.095 ;
        RECT 60.095 102.555 60.355 102.915 ;
        RECT 59.165 102.325 60.355 102.555 ;
        RECT 60.925 102.145 61.215 102.915 ;
        RECT 55.900 101.095 56.565 101.265 ;
        RECT 55.895 100.545 56.225 100.925 ;
        RECT 56.395 100.805 56.565 101.095 ;
        RECT 56.825 100.545 58.035 101.295 ;
        RECT 58.210 100.725 58.545 102.145 ;
        RECT 58.720 101.965 61.215 102.145 ;
        RECT 58.720 101.275 58.945 101.965 ;
        RECT 61.425 101.930 61.715 103.095 ;
        RECT 61.885 102.005 63.555 103.095 ;
        RECT 63.785 102.745 65.855 102.915 ;
        RECT 63.785 102.245 64.045 102.745 ;
        RECT 64.715 102.715 65.855 102.745 ;
        RECT 64.215 102.245 64.545 102.565 ;
        RECT 64.715 102.245 64.905 102.715 ;
        RECT 59.145 101.455 59.425 101.785 ;
        RECT 59.605 101.455 60.180 101.785 ;
        RECT 60.360 101.455 60.795 101.785 ;
        RECT 60.975 101.455 61.245 101.785 ;
        RECT 61.885 101.315 62.635 101.835 ;
        RECT 62.805 101.485 63.555 102.005 ;
        RECT 63.740 101.455 64.045 102.075 ;
        RECT 64.215 101.315 64.495 102.245 ;
        RECT 65.075 102.115 65.405 102.535 ;
        RECT 65.575 102.295 65.855 102.715 ;
        RECT 66.075 102.295 66.305 103.095 ;
        RECT 66.485 102.115 66.755 102.925 ;
        RECT 66.935 102.295 67.165 103.095 ;
        RECT 67.345 102.115 67.615 102.925 ;
        RECT 67.795 102.295 68.025 103.095 ;
        RECT 64.675 101.745 64.895 102.075 ;
        RECT 65.075 101.915 67.615 102.115 ;
        RECT 67.815 101.745 68.140 102.115 ;
        RECT 68.335 101.955 68.665 103.095 ;
        RECT 69.195 102.125 69.525 102.910 ;
        RECT 69.705 102.660 75.050 103.095 ;
        RECT 68.845 101.955 69.525 102.125 ;
        RECT 64.675 101.495 65.425 101.745 ;
        RECT 66.010 101.495 66.720 101.745 ;
        RECT 67.380 101.495 68.140 101.745 ;
        RECT 68.325 101.535 68.675 101.785 ;
        RECT 68.845 101.355 69.015 101.955 ;
        RECT 69.185 101.535 69.535 101.785 ;
        RECT 58.720 101.085 61.205 101.275 ;
        RECT 58.725 100.545 59.470 100.915 ;
        RECT 60.035 100.725 60.290 101.085 ;
        RECT 60.470 100.545 60.800 100.915 ;
        RECT 60.980 100.725 61.205 101.085 ;
        RECT 61.425 100.545 61.715 101.270 ;
        RECT 61.885 100.545 63.555 101.315 ;
        RECT 63.785 100.545 64.035 101.275 ;
        RECT 64.215 101.115 66.785 101.315 ;
        RECT 64.215 100.715 64.475 101.115 ;
        RECT 64.645 100.545 64.975 100.935 ;
        RECT 65.145 100.745 65.335 101.115 ;
        RECT 66.965 101.095 68.075 101.315 ;
        RECT 66.965 100.935 67.135 101.095 ;
        RECT 65.505 100.545 65.835 100.935 ;
        RECT 66.025 100.725 67.135 100.935 ;
        RECT 67.315 100.545 67.645 100.915 ;
        RECT 67.825 100.725 68.075 101.095 ;
        RECT 68.335 100.545 68.605 101.355 ;
        RECT 68.775 100.715 69.105 101.355 ;
        RECT 69.275 100.545 69.515 101.355 ;
        RECT 71.290 101.090 71.630 101.920 ;
        RECT 73.110 101.410 73.460 102.660 ;
        RECT 75.225 102.005 76.435 103.095 ;
        RECT 75.225 101.295 75.745 101.835 ;
        RECT 75.915 101.465 76.435 102.005 ;
        RECT 69.705 100.545 75.050 101.090 ;
        RECT 75.225 100.545 76.435 101.295 ;
        RECT 76.615 100.725 76.875 102.915 ;
        RECT 77.045 102.365 77.385 103.095 ;
        RECT 77.565 102.185 77.835 102.915 ;
        RECT 77.065 101.965 77.835 102.185 ;
        RECT 78.015 102.205 78.245 102.915 ;
        RECT 78.415 102.385 78.745 103.095 ;
        RECT 78.915 102.205 79.175 102.915 ;
        RECT 78.015 101.965 79.175 102.205 ;
        RECT 79.830 102.145 80.095 102.915 ;
        RECT 80.265 102.375 80.595 103.095 ;
        RECT 80.785 102.555 81.045 102.915 ;
        RECT 81.215 102.725 81.545 103.095 ;
        RECT 81.715 102.555 81.975 102.915 ;
        RECT 80.785 102.325 81.975 102.555 ;
        RECT 82.545 102.145 82.835 102.915 ;
        RECT 77.065 101.295 77.355 101.965 ;
        RECT 77.535 101.475 78.000 101.785 ;
        RECT 78.180 101.475 78.705 101.785 ;
        RECT 77.065 101.095 78.295 101.295 ;
        RECT 77.135 100.545 77.805 100.915 ;
        RECT 77.985 100.725 78.295 101.095 ;
        RECT 78.475 100.835 78.705 101.475 ;
        RECT 78.885 101.455 79.185 101.785 ;
        RECT 78.885 100.545 79.175 101.275 ;
        RECT 79.830 100.725 80.165 102.145 ;
        RECT 80.340 101.965 82.835 102.145 ;
        RECT 80.340 101.275 80.565 101.965 ;
        RECT 83.050 101.950 83.345 103.095 ;
        RECT 80.765 101.455 81.045 101.785 ;
        RECT 81.225 101.455 81.800 101.785 ;
        RECT 81.980 101.455 82.415 101.785 ;
        RECT 82.595 101.455 82.865 101.785 ;
        RECT 80.340 101.085 82.825 101.275 ;
        RECT 80.345 100.545 81.090 100.915 ;
        RECT 81.655 100.725 81.910 101.085 ;
        RECT 82.090 100.545 82.420 100.915 ;
        RECT 82.600 100.725 82.825 101.085 ;
        RECT 83.050 100.545 83.345 101.365 ;
        RECT 83.515 101.095 83.745 102.795 ;
        RECT 83.960 102.290 84.215 103.095 ;
        RECT 84.415 102.480 84.745 102.925 ;
        RECT 84.915 102.650 85.190 103.095 ;
        RECT 85.425 102.480 85.755 102.925 ;
        RECT 84.415 102.300 85.755 102.480 ;
        RECT 86.215 102.120 86.545 102.785 ;
        RECT 83.960 101.950 86.545 102.120 ;
        RECT 83.960 101.335 84.270 101.950 ;
        RECT 87.185 101.930 87.475 103.095 ;
        RECT 87.735 102.425 87.905 102.925 ;
        RECT 88.075 102.595 88.405 103.095 ;
        RECT 87.735 102.255 88.400 102.425 ;
        RECT 84.440 101.505 84.770 101.735 ;
        RECT 84.940 101.505 85.410 101.735 ;
        RECT 85.580 101.565 86.035 101.735 ;
        RECT 85.580 101.505 86.030 101.565 ;
        RECT 86.220 101.505 86.555 101.735 ;
        RECT 87.650 101.435 88.000 102.085 ;
        RECT 83.960 101.155 86.545 101.335 ;
        RECT 83.515 100.715 83.735 101.095 ;
        RECT 83.905 100.545 84.755 100.905 ;
        RECT 85.235 100.735 85.565 101.155 ;
        RECT 85.770 100.545 86.045 100.985 ;
        RECT 86.215 100.735 86.545 101.155 ;
        RECT 87.185 100.545 87.475 101.270 ;
        RECT 88.170 101.265 88.400 102.255 ;
        RECT 87.735 101.095 88.400 101.265 ;
        RECT 87.735 100.805 87.905 101.095 ;
        RECT 88.075 100.545 88.405 100.925 ;
        RECT 88.575 100.805 88.760 102.925 ;
        RECT 89.000 102.635 89.265 103.095 ;
        RECT 89.435 102.500 89.685 102.925 ;
        RECT 89.895 102.650 91.000 102.820 ;
        RECT 89.380 102.370 89.685 102.500 ;
        RECT 88.930 101.175 89.210 102.125 ;
        RECT 89.380 101.265 89.550 102.370 ;
        RECT 89.720 101.585 89.960 102.180 ;
        RECT 90.130 102.115 90.660 102.480 ;
        RECT 90.130 101.415 90.300 102.115 ;
        RECT 90.830 102.035 91.000 102.650 ;
        RECT 91.170 102.295 91.340 103.095 ;
        RECT 91.510 102.595 91.760 102.925 ;
        RECT 91.985 102.625 92.870 102.795 ;
        RECT 90.830 101.945 91.340 102.035 ;
        RECT 89.380 101.135 89.605 101.265 ;
        RECT 89.775 101.195 90.300 101.415 ;
        RECT 90.470 101.775 91.340 101.945 ;
        RECT 89.015 100.545 89.265 101.005 ;
        RECT 89.435 100.995 89.605 101.135 ;
        RECT 90.470 100.995 90.640 101.775 ;
        RECT 91.170 101.705 91.340 101.775 ;
        RECT 90.850 101.525 91.050 101.555 ;
        RECT 91.510 101.525 91.680 102.595 ;
        RECT 91.850 101.705 92.040 102.425 ;
        RECT 90.850 101.225 91.680 101.525 ;
        RECT 92.210 101.495 92.530 102.455 ;
        RECT 89.435 100.825 89.770 100.995 ;
        RECT 89.965 100.825 90.640 100.995 ;
        RECT 90.960 100.545 91.330 101.045 ;
        RECT 91.510 100.995 91.680 101.225 ;
        RECT 92.065 101.165 92.530 101.495 ;
        RECT 92.700 101.785 92.870 102.625 ;
        RECT 93.050 102.595 93.365 103.095 ;
        RECT 93.595 102.365 93.935 102.925 ;
        RECT 93.040 101.990 93.935 102.365 ;
        RECT 94.105 102.085 94.275 103.095 ;
        RECT 93.745 101.785 93.935 101.990 ;
        RECT 94.445 102.035 94.775 102.880 ;
        RECT 95.005 102.225 95.280 102.925 ;
        RECT 95.450 102.550 95.705 103.095 ;
        RECT 95.875 102.585 96.355 102.925 ;
        RECT 96.530 102.540 97.135 103.095 ;
        RECT 96.520 102.440 97.135 102.540 ;
        RECT 96.520 102.415 96.705 102.440 ;
        RECT 94.445 101.955 94.835 102.035 ;
        RECT 94.620 101.905 94.835 101.955 ;
        RECT 92.700 101.455 93.575 101.785 ;
        RECT 93.745 101.455 94.495 101.785 ;
        RECT 92.700 100.995 92.870 101.455 ;
        RECT 93.745 101.285 93.945 101.455 ;
        RECT 94.665 101.325 94.835 101.905 ;
        RECT 94.610 101.285 94.835 101.325 ;
        RECT 91.510 100.825 91.915 100.995 ;
        RECT 92.085 100.825 92.870 100.995 ;
        RECT 93.145 100.545 93.355 101.075 ;
        RECT 93.615 100.760 93.945 101.285 ;
        RECT 94.455 101.200 94.835 101.285 ;
        RECT 94.115 100.545 94.285 101.155 ;
        RECT 94.455 100.765 94.785 101.200 ;
        RECT 95.005 101.195 95.175 102.225 ;
        RECT 95.450 102.095 96.205 102.345 ;
        RECT 96.375 102.170 96.705 102.415 ;
        RECT 95.450 102.060 96.220 102.095 ;
        RECT 95.450 102.050 96.235 102.060 ;
        RECT 95.345 102.035 96.240 102.050 ;
        RECT 95.345 102.020 96.260 102.035 ;
        RECT 95.345 102.010 96.280 102.020 ;
        RECT 95.345 102.000 96.305 102.010 ;
        RECT 95.345 101.970 96.375 102.000 ;
        RECT 95.345 101.940 96.395 101.970 ;
        RECT 95.345 101.910 96.415 101.940 ;
        RECT 95.345 101.885 96.445 101.910 ;
        RECT 95.345 101.850 96.480 101.885 ;
        RECT 95.345 101.845 96.510 101.850 ;
        RECT 95.345 101.450 95.575 101.845 ;
        RECT 96.120 101.840 96.510 101.845 ;
        RECT 96.145 101.830 96.510 101.840 ;
        RECT 96.160 101.825 96.510 101.830 ;
        RECT 96.175 101.820 96.510 101.825 ;
        RECT 96.875 101.820 97.135 102.270 ;
        RECT 97.310 101.950 97.605 103.095 ;
        RECT 96.175 101.815 97.135 101.820 ;
        RECT 96.185 101.805 97.135 101.815 ;
        RECT 96.195 101.800 97.135 101.805 ;
        RECT 96.205 101.790 97.135 101.800 ;
        RECT 96.210 101.780 97.135 101.790 ;
        RECT 96.215 101.775 97.135 101.780 ;
        RECT 96.225 101.760 97.135 101.775 ;
        RECT 96.230 101.745 97.135 101.760 ;
        RECT 96.240 101.720 97.135 101.745 ;
        RECT 95.745 101.250 96.075 101.675 ;
        RECT 95.825 101.225 96.075 101.250 ;
        RECT 95.005 100.715 95.265 101.195 ;
        RECT 95.435 100.545 95.685 101.085 ;
        RECT 95.855 100.765 96.075 101.225 ;
        RECT 96.245 101.650 97.135 101.720 ;
        RECT 96.245 100.925 96.415 101.650 ;
        RECT 96.585 101.095 97.135 101.480 ;
        RECT 96.245 100.755 97.135 100.925 ;
        RECT 97.310 100.545 97.605 101.365 ;
        RECT 97.775 101.095 98.005 102.795 ;
        RECT 98.220 102.290 98.475 103.095 ;
        RECT 98.675 102.480 99.005 102.925 ;
        RECT 99.175 102.650 99.450 103.095 ;
        RECT 99.685 102.480 100.015 102.925 ;
        RECT 98.675 102.300 100.015 102.480 ;
        RECT 100.475 102.120 100.805 102.785 ;
        RECT 98.220 101.950 100.805 102.120 ;
        RECT 100.995 101.955 101.325 103.095 ;
        RECT 101.855 102.125 102.185 102.910 ;
        RECT 101.505 101.955 102.185 102.125 ;
        RECT 102.375 102.125 102.705 102.910 ;
        RECT 102.375 101.955 103.055 102.125 ;
        RECT 103.235 101.955 103.565 103.095 ;
        RECT 103.745 102.660 109.090 103.095 ;
        RECT 98.220 101.335 98.530 101.950 ;
        RECT 98.700 101.505 99.030 101.735 ;
        RECT 99.200 101.505 99.670 101.735 ;
        RECT 99.840 101.565 100.295 101.735 ;
        RECT 99.840 101.505 100.290 101.565 ;
        RECT 100.480 101.505 100.815 101.735 ;
        RECT 100.985 101.535 101.335 101.785 ;
        RECT 101.505 101.355 101.675 101.955 ;
        RECT 101.845 101.535 102.195 101.785 ;
        RECT 102.365 101.535 102.715 101.785 ;
        RECT 102.885 101.355 103.055 101.955 ;
        RECT 103.225 101.535 103.575 101.785 ;
        RECT 98.220 101.155 100.805 101.335 ;
        RECT 97.775 100.715 97.995 101.095 ;
        RECT 98.165 100.545 99.015 100.905 ;
        RECT 99.495 100.735 99.825 101.155 ;
        RECT 100.030 100.545 100.305 100.985 ;
        RECT 100.475 100.735 100.805 101.155 ;
        RECT 100.995 100.545 101.265 101.355 ;
        RECT 101.435 100.715 101.765 101.355 ;
        RECT 101.935 100.545 102.175 101.355 ;
        RECT 102.385 100.545 102.625 101.355 ;
        RECT 102.795 100.715 103.125 101.355 ;
        RECT 103.295 100.545 103.565 101.355 ;
        RECT 105.330 101.090 105.670 101.920 ;
        RECT 107.150 101.410 107.500 102.660 ;
        RECT 109.265 102.005 112.775 103.095 ;
        RECT 109.265 101.315 110.915 101.835 ;
        RECT 111.085 101.485 112.775 102.005 ;
        RECT 112.945 101.930 113.235 103.095 ;
        RECT 113.405 101.955 113.665 103.095 ;
        RECT 113.835 101.945 114.165 102.925 ;
        RECT 114.335 101.955 114.615 103.095 ;
        RECT 115.765 102.035 116.095 102.880 ;
        RECT 116.265 102.085 116.435 103.095 ;
        RECT 116.605 102.365 116.945 102.925 ;
        RECT 117.175 102.595 117.490 103.095 ;
        RECT 117.670 102.625 118.555 102.795 ;
        RECT 115.705 101.955 116.095 102.035 ;
        RECT 116.605 101.990 117.500 102.365 ;
        RECT 113.425 101.535 113.760 101.785 ;
        RECT 113.930 101.345 114.100 101.945 ;
        RECT 115.705 101.905 115.920 101.955 ;
        RECT 114.270 101.515 114.605 101.785 ;
        RECT 103.745 100.545 109.090 101.090 ;
        RECT 109.265 100.545 112.775 101.315 ;
        RECT 112.945 100.545 113.235 101.270 ;
        RECT 113.405 100.715 114.100 101.345 ;
        RECT 114.305 100.545 114.615 101.345 ;
        RECT 115.705 101.325 115.875 101.905 ;
        RECT 116.605 101.785 116.795 101.990 ;
        RECT 117.670 101.785 117.840 102.625 ;
        RECT 118.780 102.595 119.030 102.925 ;
        RECT 116.045 101.455 116.795 101.785 ;
        RECT 116.965 101.455 117.840 101.785 ;
        RECT 115.705 101.285 115.930 101.325 ;
        RECT 116.595 101.285 116.795 101.455 ;
        RECT 115.705 101.200 116.085 101.285 ;
        RECT 115.755 100.765 116.085 101.200 ;
        RECT 116.255 100.545 116.425 101.155 ;
        RECT 116.595 100.760 116.925 101.285 ;
        RECT 117.185 100.545 117.395 101.075 ;
        RECT 117.670 100.995 117.840 101.455 ;
        RECT 118.010 101.495 118.330 102.455 ;
        RECT 118.500 101.705 118.690 102.425 ;
        RECT 118.860 101.525 119.030 102.595 ;
        RECT 119.200 102.295 119.370 103.095 ;
        RECT 119.540 102.650 120.645 102.820 ;
        RECT 119.540 102.035 119.710 102.650 ;
        RECT 120.855 102.500 121.105 102.925 ;
        RECT 121.275 102.635 121.540 103.095 ;
        RECT 119.880 102.115 120.410 102.480 ;
        RECT 120.855 102.370 121.160 102.500 ;
        RECT 119.200 101.945 119.710 102.035 ;
        RECT 119.200 101.775 120.070 101.945 ;
        RECT 119.200 101.705 119.370 101.775 ;
        RECT 119.490 101.525 119.690 101.555 ;
        RECT 118.010 101.165 118.475 101.495 ;
        RECT 118.860 101.225 119.690 101.525 ;
        RECT 118.860 100.995 119.030 101.225 ;
        RECT 117.670 100.825 118.455 100.995 ;
        RECT 118.625 100.825 119.030 100.995 ;
        RECT 119.210 100.545 119.580 101.045 ;
        RECT 119.900 100.995 120.070 101.775 ;
        RECT 120.240 101.415 120.410 102.115 ;
        RECT 120.580 101.585 120.820 102.180 ;
        RECT 120.240 101.195 120.765 101.415 ;
        RECT 120.990 101.265 121.160 102.370 ;
        RECT 120.935 101.135 121.160 101.265 ;
        RECT 121.330 101.175 121.610 102.125 ;
        RECT 120.935 100.995 121.105 101.135 ;
        RECT 119.900 100.825 120.575 100.995 ;
        RECT 120.770 100.825 121.105 100.995 ;
        RECT 121.275 100.545 121.525 101.005 ;
        RECT 121.780 100.805 121.965 102.925 ;
        RECT 122.135 102.595 122.465 103.095 ;
        RECT 122.635 102.425 122.805 102.925 ;
        RECT 122.140 102.255 122.805 102.425 ;
        RECT 122.140 101.265 122.370 102.255 ;
        RECT 122.540 101.435 122.890 102.085 ;
        RECT 123.065 102.005 124.735 103.095 ;
        RECT 124.995 102.425 125.165 102.925 ;
        RECT 125.335 102.595 125.665 103.095 ;
        RECT 124.995 102.255 125.660 102.425 ;
        RECT 123.065 101.315 123.815 101.835 ;
        RECT 123.985 101.485 124.735 102.005 ;
        RECT 124.910 101.435 125.260 102.085 ;
        RECT 122.140 101.095 122.805 101.265 ;
        RECT 122.135 100.545 122.465 100.925 ;
        RECT 122.635 100.805 122.805 101.095 ;
        RECT 123.065 100.545 124.735 101.315 ;
        RECT 125.430 101.265 125.660 102.255 ;
        RECT 124.995 101.095 125.660 101.265 ;
        RECT 124.995 100.805 125.165 101.095 ;
        RECT 125.335 100.545 125.665 100.925 ;
        RECT 125.835 100.805 126.020 102.925 ;
        RECT 126.260 102.635 126.525 103.095 ;
        RECT 126.695 102.500 126.945 102.925 ;
        RECT 127.155 102.650 128.260 102.820 ;
        RECT 126.640 102.370 126.945 102.500 ;
        RECT 126.190 101.175 126.470 102.125 ;
        RECT 126.640 101.265 126.810 102.370 ;
        RECT 126.980 101.585 127.220 102.180 ;
        RECT 127.390 102.115 127.920 102.480 ;
        RECT 127.390 101.415 127.560 102.115 ;
        RECT 128.090 102.035 128.260 102.650 ;
        RECT 128.430 102.295 128.600 103.095 ;
        RECT 128.770 102.595 129.020 102.925 ;
        RECT 129.245 102.625 130.130 102.795 ;
        RECT 128.090 101.945 128.600 102.035 ;
        RECT 126.640 101.135 126.865 101.265 ;
        RECT 127.035 101.195 127.560 101.415 ;
        RECT 127.730 101.775 128.600 101.945 ;
        RECT 126.275 100.545 126.525 101.005 ;
        RECT 126.695 100.995 126.865 101.135 ;
        RECT 127.730 100.995 127.900 101.775 ;
        RECT 128.430 101.705 128.600 101.775 ;
        RECT 128.110 101.525 128.310 101.555 ;
        RECT 128.770 101.525 128.940 102.595 ;
        RECT 129.110 101.705 129.300 102.425 ;
        RECT 128.110 101.225 128.940 101.525 ;
        RECT 129.470 101.495 129.790 102.455 ;
        RECT 126.695 100.825 127.030 100.995 ;
        RECT 127.225 100.825 127.900 100.995 ;
        RECT 128.220 100.545 128.590 101.045 ;
        RECT 128.770 100.995 128.940 101.225 ;
        RECT 129.325 101.165 129.790 101.495 ;
        RECT 129.960 101.785 130.130 102.625 ;
        RECT 130.310 102.595 130.625 103.095 ;
        RECT 130.855 102.365 131.195 102.925 ;
        RECT 130.300 101.990 131.195 102.365 ;
        RECT 131.365 102.085 131.535 103.095 ;
        RECT 131.005 101.785 131.195 101.990 ;
        RECT 131.705 102.035 132.035 102.880 ;
        RECT 131.705 101.955 132.095 102.035 ;
        RECT 131.880 101.905 132.095 101.955 ;
        RECT 129.960 101.455 130.835 101.785 ;
        RECT 131.005 101.455 131.755 101.785 ;
        RECT 129.960 100.995 130.130 101.455 ;
        RECT 131.005 101.285 131.205 101.455 ;
        RECT 131.925 101.325 132.095 101.905 ;
        RECT 131.870 101.285 132.095 101.325 ;
        RECT 128.770 100.825 129.175 100.995 ;
        RECT 129.345 100.825 130.130 100.995 ;
        RECT 130.405 100.545 130.615 101.075 ;
        RECT 130.875 100.760 131.205 101.285 ;
        RECT 131.715 101.200 132.095 101.285 ;
        RECT 132.265 101.955 132.650 102.925 ;
        RECT 132.820 102.635 133.145 103.095 ;
        RECT 133.665 102.465 133.945 102.925 ;
        RECT 132.820 102.245 133.945 102.465 ;
        RECT 132.265 101.285 132.545 101.955 ;
        RECT 132.820 101.785 133.270 102.245 ;
        RECT 134.135 102.075 134.535 102.925 ;
        RECT 134.935 102.635 135.205 103.095 ;
        RECT 135.375 102.465 135.660 102.925 ;
        RECT 132.715 101.455 133.270 101.785 ;
        RECT 133.440 101.515 134.535 102.075 ;
        RECT 132.820 101.345 133.270 101.455 ;
        RECT 131.375 100.545 131.545 101.155 ;
        RECT 131.715 100.765 132.045 101.200 ;
        RECT 132.265 100.715 132.650 101.285 ;
        RECT 132.820 101.175 133.945 101.345 ;
        RECT 132.820 100.545 133.145 101.005 ;
        RECT 133.665 100.715 133.945 101.175 ;
        RECT 134.135 100.715 134.535 101.515 ;
        RECT 134.705 102.245 135.660 102.465 ;
        RECT 134.705 101.345 134.915 102.245 ;
        RECT 135.085 101.515 135.775 102.075 ;
        RECT 135.945 101.955 136.215 102.925 ;
        RECT 136.425 102.295 136.705 103.095 ;
        RECT 136.875 102.585 138.530 102.875 ;
        RECT 136.940 102.245 138.530 102.415 ;
        RECT 136.940 102.125 137.110 102.245 ;
        RECT 136.385 101.955 137.110 102.125 ;
        RECT 134.705 101.175 135.660 101.345 ;
        RECT 134.935 100.545 135.205 101.005 ;
        RECT 135.375 100.715 135.660 101.175 ;
        RECT 135.945 101.220 136.115 101.955 ;
        RECT 136.385 101.785 136.555 101.955 ;
        RECT 137.300 101.905 138.015 102.075 ;
        RECT 138.210 101.955 138.530 102.245 ;
        RECT 138.705 101.930 138.995 103.095 ;
        RECT 139.175 101.985 139.470 103.095 ;
        RECT 136.285 101.455 136.555 101.785 ;
        RECT 136.725 101.455 137.130 101.785 ;
        RECT 137.300 101.455 138.010 101.905 ;
        RECT 139.650 101.785 139.900 102.920 ;
        RECT 140.070 101.985 140.330 103.095 ;
        RECT 140.500 102.195 140.760 102.920 ;
        RECT 140.930 102.365 141.190 103.095 ;
        RECT 141.360 102.195 141.620 102.920 ;
        RECT 141.790 102.365 142.050 103.095 ;
        RECT 142.220 102.195 142.480 102.920 ;
        RECT 142.650 102.365 142.910 103.095 ;
        RECT 143.080 102.195 143.340 102.920 ;
        RECT 143.510 102.365 143.805 103.095 ;
        RECT 140.500 101.955 143.810 102.195 ;
        RECT 144.430 102.125 144.760 102.925 ;
        RECT 144.930 102.295 145.260 103.095 ;
        RECT 145.560 102.125 145.890 102.925 ;
        RECT 146.535 102.295 146.785 103.095 ;
        RECT 144.430 101.955 146.865 102.125 ;
        RECT 147.055 101.955 147.225 103.095 ;
        RECT 147.395 101.955 147.735 102.925 ;
        RECT 148.455 102.425 148.625 102.925 ;
        RECT 148.795 102.595 149.125 103.095 ;
        RECT 148.455 102.255 149.120 102.425 ;
        RECT 136.385 101.285 136.555 101.455 ;
        RECT 135.945 100.875 136.215 101.220 ;
        RECT 136.385 101.115 137.995 101.285 ;
        RECT 138.180 101.215 138.530 101.785 ;
        RECT 136.405 100.545 136.785 100.945 ;
        RECT 136.955 100.765 137.125 101.115 ;
        RECT 137.295 100.545 137.625 100.945 ;
        RECT 137.825 100.765 137.995 101.115 ;
        RECT 138.195 100.545 138.525 101.045 ;
        RECT 138.705 100.545 138.995 101.270 ;
        RECT 139.165 101.175 139.480 101.785 ;
        RECT 139.650 101.535 142.670 101.785 ;
        RECT 139.225 100.545 139.470 101.005 ;
        RECT 139.650 100.725 139.900 101.535 ;
        RECT 142.840 101.365 143.810 101.955 ;
        RECT 144.225 101.535 144.575 101.785 ;
        RECT 140.500 101.195 143.810 101.365 ;
        RECT 144.760 101.325 144.930 101.955 ;
        RECT 145.100 101.535 145.430 101.735 ;
        RECT 145.600 101.535 145.930 101.735 ;
        RECT 146.100 101.535 146.520 101.735 ;
        RECT 146.695 101.705 146.865 101.955 ;
        RECT 146.695 101.535 147.390 101.705 ;
        RECT 140.070 100.545 140.330 101.070 ;
        RECT 140.500 100.740 140.760 101.195 ;
        RECT 140.930 100.545 141.190 101.025 ;
        RECT 141.360 100.740 141.620 101.195 ;
        RECT 141.790 100.545 142.050 101.025 ;
        RECT 142.220 100.740 142.480 101.195 ;
        RECT 142.650 100.545 142.910 101.025 ;
        RECT 143.080 100.740 143.340 101.195 ;
        RECT 143.510 100.545 143.810 101.025 ;
        RECT 144.430 100.715 144.930 101.325 ;
        RECT 145.560 101.195 146.785 101.365 ;
        RECT 147.560 101.345 147.735 101.955 ;
        RECT 148.370 101.435 148.720 102.085 ;
        RECT 145.560 100.715 145.890 101.195 ;
        RECT 146.060 100.545 146.285 101.005 ;
        RECT 146.455 100.715 146.785 101.195 ;
        RECT 146.975 100.545 147.225 101.345 ;
        RECT 147.395 100.715 147.735 101.345 ;
        RECT 148.890 101.265 149.120 102.255 ;
        RECT 148.455 101.095 149.120 101.265 ;
        RECT 148.455 100.805 148.625 101.095 ;
        RECT 148.795 100.545 149.125 100.925 ;
        RECT 149.295 100.805 149.480 102.925 ;
        RECT 149.720 102.635 149.985 103.095 ;
        RECT 150.155 102.500 150.405 102.925 ;
        RECT 150.615 102.650 151.720 102.820 ;
        RECT 150.100 102.370 150.405 102.500 ;
        RECT 149.650 101.175 149.930 102.125 ;
        RECT 150.100 101.265 150.270 102.370 ;
        RECT 150.440 101.585 150.680 102.180 ;
        RECT 150.850 102.115 151.380 102.480 ;
        RECT 150.850 101.415 151.020 102.115 ;
        RECT 151.550 102.035 151.720 102.650 ;
        RECT 151.890 102.295 152.060 103.095 ;
        RECT 152.230 102.595 152.480 102.925 ;
        RECT 152.705 102.625 153.590 102.795 ;
        RECT 151.550 101.945 152.060 102.035 ;
        RECT 150.100 101.135 150.325 101.265 ;
        RECT 150.495 101.195 151.020 101.415 ;
        RECT 151.190 101.775 152.060 101.945 ;
        RECT 149.735 100.545 149.985 101.005 ;
        RECT 150.155 100.995 150.325 101.135 ;
        RECT 151.190 100.995 151.360 101.775 ;
        RECT 151.890 101.705 152.060 101.775 ;
        RECT 151.570 101.525 151.770 101.555 ;
        RECT 152.230 101.525 152.400 102.595 ;
        RECT 152.570 101.705 152.760 102.425 ;
        RECT 151.570 101.225 152.400 101.525 ;
        RECT 152.930 101.495 153.250 102.455 ;
        RECT 150.155 100.825 150.490 100.995 ;
        RECT 150.685 100.825 151.360 100.995 ;
        RECT 151.680 100.545 152.050 101.045 ;
        RECT 152.230 100.995 152.400 101.225 ;
        RECT 152.785 101.165 153.250 101.495 ;
        RECT 153.420 101.785 153.590 102.625 ;
        RECT 153.770 102.595 154.085 103.095 ;
        RECT 154.315 102.365 154.655 102.925 ;
        RECT 153.760 101.990 154.655 102.365 ;
        RECT 154.825 102.085 154.995 103.095 ;
        RECT 154.465 101.785 154.655 101.990 ;
        RECT 155.165 102.035 155.495 102.880 ;
        RECT 155.165 101.955 155.555 102.035 ;
        RECT 155.340 101.905 155.555 101.955 ;
        RECT 153.420 101.455 154.295 101.785 ;
        RECT 154.465 101.455 155.215 101.785 ;
        RECT 153.420 100.995 153.590 101.455 ;
        RECT 154.465 101.285 154.665 101.455 ;
        RECT 155.385 101.325 155.555 101.905 ;
        RECT 155.725 102.005 156.935 103.095 ;
        RECT 155.725 101.465 156.245 102.005 ;
        RECT 155.330 101.285 155.555 101.325 ;
        RECT 156.415 101.295 156.935 101.835 ;
        RECT 152.230 100.825 152.635 100.995 ;
        RECT 152.805 100.825 153.590 100.995 ;
        RECT 153.865 100.545 154.075 101.075 ;
        RECT 154.335 100.760 154.665 101.285 ;
        RECT 155.175 101.200 155.555 101.285 ;
        RECT 154.835 100.545 155.005 101.155 ;
        RECT 155.175 100.765 155.505 101.200 ;
        RECT 155.725 100.545 156.935 101.295 ;
        RECT 22.700 100.375 157.020 100.545 ;
        RECT 22.785 99.625 23.995 100.375 ;
        RECT 24.255 99.825 24.425 100.115 ;
        RECT 24.595 99.995 24.925 100.375 ;
        RECT 24.255 99.655 24.920 99.825 ;
        RECT 22.785 99.085 23.305 99.625 ;
        RECT 23.475 98.915 23.995 99.455 ;
        RECT 22.785 97.825 23.995 98.915 ;
        RECT 24.170 98.835 24.520 99.485 ;
        RECT 24.690 98.665 24.920 99.655 ;
        RECT 24.255 98.495 24.920 98.665 ;
        RECT 24.255 97.995 24.425 98.495 ;
        RECT 24.595 97.825 24.925 98.325 ;
        RECT 25.095 97.995 25.280 100.115 ;
        RECT 25.535 99.915 25.785 100.375 ;
        RECT 25.955 99.925 26.290 100.095 ;
        RECT 26.485 99.925 27.160 100.095 ;
        RECT 25.955 99.785 26.125 99.925 ;
        RECT 25.450 98.795 25.730 99.745 ;
        RECT 25.900 99.655 26.125 99.785 ;
        RECT 25.900 98.550 26.070 99.655 ;
        RECT 26.295 99.505 26.820 99.725 ;
        RECT 26.240 98.740 26.480 99.335 ;
        RECT 26.650 98.805 26.820 99.505 ;
        RECT 26.990 99.145 27.160 99.925 ;
        RECT 27.480 99.875 27.850 100.375 ;
        RECT 28.030 99.925 28.435 100.095 ;
        RECT 28.605 99.925 29.390 100.095 ;
        RECT 28.030 99.695 28.200 99.925 ;
        RECT 27.370 99.395 28.200 99.695 ;
        RECT 28.585 99.425 29.050 99.755 ;
        RECT 27.370 99.365 27.570 99.395 ;
        RECT 27.690 99.145 27.860 99.215 ;
        RECT 26.990 98.975 27.860 99.145 ;
        RECT 27.350 98.885 27.860 98.975 ;
        RECT 25.900 98.420 26.205 98.550 ;
        RECT 26.650 98.440 27.180 98.805 ;
        RECT 25.520 97.825 25.785 98.285 ;
        RECT 25.955 97.995 26.205 98.420 ;
        RECT 27.350 98.270 27.520 98.885 ;
        RECT 26.415 98.100 27.520 98.270 ;
        RECT 27.690 97.825 27.860 98.625 ;
        RECT 28.030 98.325 28.200 99.395 ;
        RECT 28.370 98.495 28.560 99.215 ;
        RECT 28.730 98.465 29.050 99.425 ;
        RECT 29.220 99.465 29.390 99.925 ;
        RECT 29.665 99.845 29.875 100.375 ;
        RECT 30.135 99.635 30.465 100.160 ;
        RECT 30.635 99.765 30.805 100.375 ;
        RECT 30.975 99.720 31.305 100.155 ;
        RECT 32.445 99.725 32.705 100.205 ;
        RECT 32.875 99.835 33.125 100.375 ;
        RECT 30.975 99.635 31.355 99.720 ;
        RECT 30.265 99.465 30.465 99.635 ;
        RECT 31.130 99.595 31.355 99.635 ;
        RECT 29.220 99.135 30.095 99.465 ;
        RECT 30.265 99.135 31.015 99.465 ;
        RECT 28.030 97.995 28.280 98.325 ;
        RECT 29.220 98.295 29.390 99.135 ;
        RECT 30.265 98.930 30.455 99.135 ;
        RECT 31.185 99.015 31.355 99.595 ;
        RECT 31.140 98.965 31.355 99.015 ;
        RECT 29.560 98.555 30.455 98.930 ;
        RECT 30.965 98.885 31.355 98.965 ;
        RECT 28.505 98.125 29.390 98.295 ;
        RECT 29.570 97.825 29.885 98.325 ;
        RECT 30.115 97.995 30.455 98.555 ;
        RECT 30.625 97.825 30.795 98.835 ;
        RECT 30.965 98.040 31.295 98.885 ;
        RECT 32.445 98.695 32.615 99.725 ;
        RECT 33.295 99.670 33.515 100.155 ;
        RECT 32.785 99.075 33.015 99.470 ;
        RECT 33.185 99.245 33.515 99.670 ;
        RECT 33.685 99.995 34.575 100.165 ;
        RECT 33.685 99.270 33.855 99.995 ;
        RECT 34.025 99.440 34.575 99.825 ;
        RECT 34.945 99.745 35.275 100.105 ;
        RECT 35.895 99.915 36.145 100.375 ;
        RECT 36.315 99.915 36.875 100.205 ;
        RECT 34.945 99.555 36.335 99.745 ;
        RECT 36.165 99.465 36.335 99.555 ;
        RECT 33.685 99.200 34.575 99.270 ;
        RECT 33.680 99.175 34.575 99.200 ;
        RECT 33.670 99.160 34.575 99.175 ;
        RECT 33.665 99.145 34.575 99.160 ;
        RECT 33.655 99.140 34.575 99.145 ;
        RECT 33.650 99.130 34.575 99.140 ;
        RECT 33.645 99.120 34.575 99.130 ;
        RECT 33.635 99.115 34.575 99.120 ;
        RECT 33.625 99.105 34.575 99.115 ;
        RECT 33.615 99.100 34.575 99.105 ;
        RECT 33.615 99.095 33.950 99.100 ;
        RECT 33.600 99.090 33.950 99.095 ;
        RECT 33.585 99.080 33.950 99.090 ;
        RECT 33.560 99.075 33.950 99.080 ;
        RECT 32.785 99.070 33.950 99.075 ;
        RECT 32.785 99.035 33.920 99.070 ;
        RECT 32.785 99.010 33.885 99.035 ;
        RECT 32.785 98.980 33.855 99.010 ;
        RECT 32.785 98.950 33.835 98.980 ;
        RECT 32.785 98.920 33.815 98.950 ;
        RECT 32.785 98.910 33.745 98.920 ;
        RECT 32.785 98.900 33.720 98.910 ;
        RECT 32.785 98.885 33.700 98.900 ;
        RECT 32.785 98.870 33.680 98.885 ;
        RECT 32.890 98.860 33.675 98.870 ;
        RECT 32.890 98.825 33.660 98.860 ;
        RECT 32.445 97.995 32.720 98.695 ;
        RECT 32.890 98.575 33.645 98.825 ;
        RECT 33.815 98.505 34.145 98.750 ;
        RECT 34.315 98.650 34.575 99.100 ;
        RECT 34.760 99.135 35.435 99.385 ;
        RECT 35.655 99.135 35.995 99.385 ;
        RECT 36.165 99.135 36.455 99.465 ;
        RECT 34.760 98.775 35.025 99.135 ;
        RECT 36.165 98.885 36.335 99.135 ;
        RECT 35.395 98.715 36.335 98.885 ;
        RECT 33.960 98.480 34.145 98.505 ;
        RECT 33.960 98.380 34.575 98.480 ;
        RECT 32.890 97.825 33.145 98.370 ;
        RECT 33.315 97.995 33.795 98.335 ;
        RECT 33.970 97.825 34.575 98.380 ;
        RECT 34.945 97.825 35.225 98.495 ;
        RECT 35.395 98.165 35.695 98.715 ;
        RECT 36.625 98.545 36.875 99.915 ;
        RECT 37.045 99.575 37.740 100.205 ;
        RECT 37.945 99.575 38.255 100.375 ;
        RECT 38.425 99.830 43.770 100.375 ;
        RECT 37.565 99.525 37.740 99.575 ;
        RECT 37.065 99.135 37.400 99.385 ;
        RECT 37.570 98.975 37.740 99.525 ;
        RECT 37.910 99.135 38.245 99.405 ;
        RECT 40.010 99.000 40.350 99.830 ;
        RECT 43.945 99.605 47.455 100.375 ;
        RECT 48.545 99.650 48.835 100.375 ;
        RECT 49.005 99.830 54.350 100.375 ;
        RECT 35.895 97.825 36.225 98.545 ;
        RECT 36.415 97.995 36.875 98.545 ;
        RECT 37.045 97.825 37.305 98.965 ;
        RECT 37.475 97.995 37.805 98.975 ;
        RECT 37.975 97.825 38.255 98.965 ;
        RECT 41.830 98.260 42.180 99.510 ;
        RECT 43.945 99.085 45.595 99.605 ;
        RECT 45.765 98.915 47.455 99.435 ;
        RECT 50.590 99.000 50.930 99.830 ;
        RECT 55.445 99.635 55.910 100.180 ;
        RECT 38.425 97.825 43.770 98.260 ;
        RECT 43.945 97.825 47.455 98.915 ;
        RECT 48.545 97.825 48.835 98.990 ;
        RECT 52.410 98.260 52.760 99.510 ;
        RECT 55.445 98.675 55.615 99.635 ;
        RECT 56.415 99.555 56.585 100.375 ;
        RECT 56.755 99.725 57.085 100.205 ;
        RECT 57.255 99.985 57.605 100.375 ;
        RECT 57.775 99.805 58.005 100.205 ;
        RECT 57.495 99.725 58.005 99.805 ;
        RECT 56.755 99.635 58.005 99.725 ;
        RECT 58.175 99.635 58.495 100.115 ;
        RECT 56.755 99.555 57.665 99.635 ;
        RECT 55.785 99.015 56.030 99.465 ;
        RECT 56.290 99.185 56.985 99.385 ;
        RECT 57.155 99.215 57.755 99.385 ;
        RECT 57.155 99.015 57.325 99.215 ;
        RECT 57.985 99.045 58.155 99.465 ;
        RECT 55.785 98.845 57.325 99.015 ;
        RECT 57.495 98.875 58.155 99.045 ;
        RECT 57.495 98.675 57.665 98.875 ;
        RECT 58.325 98.705 58.495 99.635 ;
        RECT 58.665 99.605 62.175 100.375 ;
        RECT 58.665 99.085 60.315 99.605 ;
        RECT 62.350 99.555 62.645 100.375 ;
        RECT 62.815 99.825 63.035 100.205 ;
        RECT 63.205 100.015 64.055 100.375 ;
        RECT 60.485 98.915 62.175 99.435 ;
        RECT 55.445 98.505 57.665 98.675 ;
        RECT 57.835 98.505 58.495 98.705 ;
        RECT 49.005 97.825 54.350 98.260 ;
        RECT 55.445 97.825 55.745 98.335 ;
        RECT 55.915 97.995 56.245 98.505 ;
        RECT 57.835 98.335 58.005 98.505 ;
        RECT 56.415 97.825 57.045 98.335 ;
        RECT 57.625 98.165 58.005 98.335 ;
        RECT 58.175 97.825 58.475 98.335 ;
        RECT 58.665 97.825 62.175 98.915 ;
        RECT 62.350 97.825 62.645 98.970 ;
        RECT 62.815 98.125 63.045 99.825 ;
        RECT 64.535 99.765 64.865 100.185 ;
        RECT 65.070 99.935 65.345 100.375 ;
        RECT 65.515 99.765 65.845 100.185 ;
        RECT 63.260 99.585 65.845 99.765 ;
        RECT 66.025 99.605 69.535 100.375 ;
        RECT 69.705 99.625 70.915 100.375 ;
        RECT 63.260 98.970 63.570 99.585 ;
        RECT 63.740 99.185 64.070 99.415 ;
        RECT 64.240 99.185 64.710 99.415 ;
        RECT 64.880 99.355 65.330 99.415 ;
        RECT 64.880 99.185 65.335 99.355 ;
        RECT 65.520 99.185 65.855 99.415 ;
        RECT 66.025 99.085 67.675 99.605 ;
        RECT 63.260 98.800 65.845 98.970 ;
        RECT 67.845 98.915 69.535 99.435 ;
        RECT 69.705 99.085 70.225 99.625 ;
        RECT 71.085 99.575 71.780 100.205 ;
        RECT 71.985 99.575 72.295 100.375 ;
        RECT 72.465 99.605 74.135 100.375 ;
        RECT 74.305 99.650 74.595 100.375 ;
        RECT 74.855 99.825 75.025 100.115 ;
        RECT 75.195 99.995 75.525 100.375 ;
        RECT 74.855 99.655 75.520 99.825 ;
        RECT 70.395 98.915 70.915 99.455 ;
        RECT 71.105 99.135 71.440 99.385 ;
        RECT 71.610 98.975 71.780 99.575 ;
        RECT 71.950 99.135 72.285 99.405 ;
        RECT 72.465 99.085 73.215 99.605 ;
        RECT 63.260 97.825 63.515 98.630 ;
        RECT 63.715 98.440 65.055 98.620 ;
        RECT 63.715 97.995 64.045 98.440 ;
        RECT 64.215 97.825 64.490 98.270 ;
        RECT 64.725 97.995 65.055 98.440 ;
        RECT 65.515 98.135 65.845 98.800 ;
        RECT 66.025 97.825 69.535 98.915 ;
        RECT 69.705 97.825 70.915 98.915 ;
        RECT 71.085 97.825 71.345 98.965 ;
        RECT 71.515 97.995 71.845 98.975 ;
        RECT 72.015 97.825 72.295 98.965 ;
        RECT 73.385 98.915 74.135 99.435 ;
        RECT 72.465 97.825 74.135 98.915 ;
        RECT 74.305 97.825 74.595 98.990 ;
        RECT 74.770 98.835 75.120 99.485 ;
        RECT 75.290 98.665 75.520 99.655 ;
        RECT 74.855 98.495 75.520 98.665 ;
        RECT 74.855 97.995 75.025 98.495 ;
        RECT 75.195 97.825 75.525 98.325 ;
        RECT 75.695 97.995 75.880 100.115 ;
        RECT 76.135 99.915 76.385 100.375 ;
        RECT 76.555 99.925 76.890 100.095 ;
        RECT 77.085 99.925 77.760 100.095 ;
        RECT 76.555 99.785 76.725 99.925 ;
        RECT 76.050 98.795 76.330 99.745 ;
        RECT 76.500 99.655 76.725 99.785 ;
        RECT 76.500 98.550 76.670 99.655 ;
        RECT 76.895 99.505 77.420 99.725 ;
        RECT 76.840 98.740 77.080 99.335 ;
        RECT 77.250 98.805 77.420 99.505 ;
        RECT 77.590 99.145 77.760 99.925 ;
        RECT 78.080 99.875 78.450 100.375 ;
        RECT 78.630 99.925 79.035 100.095 ;
        RECT 79.205 99.925 79.990 100.095 ;
        RECT 78.630 99.695 78.800 99.925 ;
        RECT 77.970 99.395 78.800 99.695 ;
        RECT 79.185 99.425 79.650 99.755 ;
        RECT 77.970 99.365 78.170 99.395 ;
        RECT 78.290 99.145 78.460 99.215 ;
        RECT 77.590 98.975 78.460 99.145 ;
        RECT 77.950 98.885 78.460 98.975 ;
        RECT 76.500 98.420 76.805 98.550 ;
        RECT 77.250 98.440 77.780 98.805 ;
        RECT 76.120 97.825 76.385 98.285 ;
        RECT 76.555 97.995 76.805 98.420 ;
        RECT 77.950 98.270 78.120 98.885 ;
        RECT 77.015 98.100 78.120 98.270 ;
        RECT 78.290 97.825 78.460 98.625 ;
        RECT 78.630 98.325 78.800 99.395 ;
        RECT 78.970 98.495 79.160 99.215 ;
        RECT 79.330 98.465 79.650 99.425 ;
        RECT 79.820 99.465 79.990 99.925 ;
        RECT 80.265 99.845 80.475 100.375 ;
        RECT 80.735 99.635 81.065 100.160 ;
        RECT 81.235 99.765 81.405 100.375 ;
        RECT 81.575 99.720 81.905 100.155 ;
        RECT 81.575 99.635 81.955 99.720 ;
        RECT 80.865 99.465 81.065 99.635 ;
        RECT 81.730 99.595 81.955 99.635 ;
        RECT 79.820 99.135 80.695 99.465 ;
        RECT 80.865 99.135 81.615 99.465 ;
        RECT 78.630 97.995 78.880 98.325 ;
        RECT 79.820 98.295 79.990 99.135 ;
        RECT 80.865 98.930 81.055 99.135 ;
        RECT 81.785 99.015 81.955 99.595 ;
        RECT 82.130 99.555 82.425 100.375 ;
        RECT 82.595 99.825 82.815 100.205 ;
        RECT 82.985 100.015 83.835 100.375 ;
        RECT 81.740 98.965 81.955 99.015 ;
        RECT 80.160 98.555 81.055 98.930 ;
        RECT 81.565 98.885 81.955 98.965 ;
        RECT 79.105 98.125 79.990 98.295 ;
        RECT 80.170 97.825 80.485 98.325 ;
        RECT 80.715 97.995 81.055 98.555 ;
        RECT 81.225 97.825 81.395 98.835 ;
        RECT 81.565 98.040 81.895 98.885 ;
        RECT 82.130 97.825 82.425 98.970 ;
        RECT 82.595 98.125 82.825 99.825 ;
        RECT 84.315 99.765 84.645 100.185 ;
        RECT 84.850 99.935 85.125 100.375 ;
        RECT 85.295 99.765 85.625 100.185 ;
        RECT 83.040 99.585 85.625 99.765 ;
        RECT 85.805 99.605 89.315 100.375 ;
        RECT 83.040 98.970 83.350 99.585 ;
        RECT 83.520 99.185 83.850 99.415 ;
        RECT 84.020 99.185 84.490 99.415 ;
        RECT 84.660 99.355 85.110 99.415 ;
        RECT 84.660 99.185 85.115 99.355 ;
        RECT 85.300 99.185 85.635 99.415 ;
        RECT 85.805 99.085 87.455 99.605 ;
        RECT 83.040 98.800 85.625 98.970 ;
        RECT 87.625 98.915 89.315 99.435 ;
        RECT 83.040 97.825 83.295 98.630 ;
        RECT 83.495 98.440 84.835 98.620 ;
        RECT 83.495 97.995 83.825 98.440 ;
        RECT 83.995 97.825 84.270 98.270 ;
        RECT 84.505 97.995 84.835 98.440 ;
        RECT 85.295 98.135 85.625 98.800 ;
        RECT 85.805 97.825 89.315 98.915 ;
        RECT 89.495 98.005 89.755 100.195 ;
        RECT 90.015 100.005 90.685 100.375 ;
        RECT 90.865 99.825 91.175 100.195 ;
        RECT 89.945 99.625 91.175 99.825 ;
        RECT 89.945 98.955 90.235 99.625 ;
        RECT 91.355 99.445 91.585 100.085 ;
        RECT 91.765 99.645 92.055 100.375 ;
        RECT 92.245 99.605 95.755 100.375 ;
        RECT 90.415 99.135 90.880 99.445 ;
        RECT 91.060 99.135 91.585 99.445 ;
        RECT 91.765 99.135 92.065 99.465 ;
        RECT 92.245 99.085 93.895 99.605 ;
        RECT 96.390 99.555 96.685 100.375 ;
        RECT 96.855 99.825 97.075 100.205 ;
        RECT 97.245 100.015 98.095 100.375 ;
        RECT 89.945 98.735 90.715 98.955 ;
        RECT 89.925 97.825 90.265 98.555 ;
        RECT 90.445 98.005 90.715 98.735 ;
        RECT 90.895 98.715 92.055 98.955 ;
        RECT 94.065 98.915 95.755 99.435 ;
        RECT 90.895 98.005 91.125 98.715 ;
        RECT 91.295 97.825 91.625 98.535 ;
        RECT 91.795 98.005 92.055 98.715 ;
        RECT 92.245 97.825 95.755 98.915 ;
        RECT 96.390 97.825 96.685 98.970 ;
        RECT 96.855 98.125 97.085 99.825 ;
        RECT 98.575 99.765 98.905 100.185 ;
        RECT 99.110 99.935 99.385 100.375 ;
        RECT 99.555 99.765 99.885 100.185 ;
        RECT 97.300 99.585 99.885 99.765 ;
        RECT 100.065 99.650 100.355 100.375 ;
        RECT 100.525 99.605 104.035 100.375 ;
        RECT 105.215 99.825 105.385 100.115 ;
        RECT 105.555 99.995 105.885 100.375 ;
        RECT 105.215 99.655 105.880 99.825 ;
        RECT 97.300 98.970 97.610 99.585 ;
        RECT 97.780 99.185 98.110 99.415 ;
        RECT 98.280 99.185 98.750 99.415 ;
        RECT 98.920 99.355 99.370 99.415 ;
        RECT 98.920 99.185 99.375 99.355 ;
        RECT 99.560 99.185 99.895 99.415 ;
        RECT 100.525 99.085 102.175 99.605 ;
        RECT 97.300 98.800 99.885 98.970 ;
        RECT 97.300 97.825 97.555 98.630 ;
        RECT 97.755 98.440 99.095 98.620 ;
        RECT 97.755 97.995 98.085 98.440 ;
        RECT 98.255 97.825 98.530 98.270 ;
        RECT 98.765 97.995 99.095 98.440 ;
        RECT 99.555 98.135 99.885 98.800 ;
        RECT 100.065 97.825 100.355 98.990 ;
        RECT 102.345 98.915 104.035 99.435 ;
        RECT 100.525 97.825 104.035 98.915 ;
        RECT 105.130 98.835 105.480 99.485 ;
        RECT 105.650 98.665 105.880 99.655 ;
        RECT 105.215 98.495 105.880 98.665 ;
        RECT 105.215 97.995 105.385 98.495 ;
        RECT 105.555 97.825 105.885 98.325 ;
        RECT 106.055 97.995 106.240 100.115 ;
        RECT 106.495 99.915 106.745 100.375 ;
        RECT 106.915 99.925 107.250 100.095 ;
        RECT 107.445 99.925 108.120 100.095 ;
        RECT 106.915 99.785 107.085 99.925 ;
        RECT 106.410 98.795 106.690 99.745 ;
        RECT 106.860 99.655 107.085 99.785 ;
        RECT 106.860 98.550 107.030 99.655 ;
        RECT 107.255 99.505 107.780 99.725 ;
        RECT 107.200 98.740 107.440 99.335 ;
        RECT 107.610 98.805 107.780 99.505 ;
        RECT 107.950 99.145 108.120 99.925 ;
        RECT 108.440 99.875 108.810 100.375 ;
        RECT 108.990 99.925 109.395 100.095 ;
        RECT 109.565 99.925 110.350 100.095 ;
        RECT 108.990 99.695 109.160 99.925 ;
        RECT 108.330 99.395 109.160 99.695 ;
        RECT 109.545 99.425 110.010 99.755 ;
        RECT 108.330 99.365 108.530 99.395 ;
        RECT 108.650 99.145 108.820 99.215 ;
        RECT 107.950 98.975 108.820 99.145 ;
        RECT 108.310 98.885 108.820 98.975 ;
        RECT 106.860 98.420 107.165 98.550 ;
        RECT 107.610 98.440 108.140 98.805 ;
        RECT 106.480 97.825 106.745 98.285 ;
        RECT 106.915 97.995 107.165 98.420 ;
        RECT 108.310 98.270 108.480 98.885 ;
        RECT 107.375 98.100 108.480 98.270 ;
        RECT 108.650 97.825 108.820 98.625 ;
        RECT 108.990 98.325 109.160 99.395 ;
        RECT 109.330 98.495 109.520 99.215 ;
        RECT 109.690 98.465 110.010 99.425 ;
        RECT 110.180 99.465 110.350 99.925 ;
        RECT 110.625 99.845 110.835 100.375 ;
        RECT 111.095 99.635 111.425 100.160 ;
        RECT 111.595 99.765 111.765 100.375 ;
        RECT 111.935 99.720 112.265 100.155 ;
        RECT 111.935 99.635 112.315 99.720 ;
        RECT 111.225 99.465 111.425 99.635 ;
        RECT 112.090 99.595 112.315 99.635 ;
        RECT 110.180 99.135 111.055 99.465 ;
        RECT 111.225 99.135 111.975 99.465 ;
        RECT 108.990 97.995 109.240 98.325 ;
        RECT 110.180 98.295 110.350 99.135 ;
        RECT 111.225 98.930 111.415 99.135 ;
        RECT 112.145 99.015 112.315 99.595 ;
        RECT 112.100 98.965 112.315 99.015 ;
        RECT 110.520 98.555 111.415 98.930 ;
        RECT 111.925 98.885 112.315 98.965 ;
        RECT 112.945 99.635 113.330 100.205 ;
        RECT 113.500 99.915 113.825 100.375 ;
        RECT 114.345 99.745 114.625 100.205 ;
        RECT 112.945 98.965 113.225 99.635 ;
        RECT 113.500 99.575 114.625 99.745 ;
        RECT 113.500 99.465 113.950 99.575 ;
        RECT 113.395 99.135 113.950 99.465 ;
        RECT 114.815 99.405 115.215 100.205 ;
        RECT 115.615 99.915 115.885 100.375 ;
        RECT 116.055 99.745 116.340 100.205 ;
        RECT 109.465 98.125 110.350 98.295 ;
        RECT 110.530 97.825 110.845 98.325 ;
        RECT 111.075 97.995 111.415 98.555 ;
        RECT 111.585 97.825 111.755 98.835 ;
        RECT 111.925 98.040 112.255 98.885 ;
        RECT 112.945 97.995 113.330 98.965 ;
        RECT 113.500 98.675 113.950 99.135 ;
        RECT 114.120 98.845 115.215 99.405 ;
        RECT 113.500 98.455 114.625 98.675 ;
        RECT 113.500 97.825 113.825 98.285 ;
        RECT 114.345 97.995 114.625 98.455 ;
        RECT 114.815 97.995 115.215 98.845 ;
        RECT 115.385 99.575 116.340 99.745 ;
        RECT 116.640 99.595 116.935 100.375 ;
        RECT 117.495 99.845 117.840 100.205 ;
        RECT 118.300 100.015 118.630 100.375 ;
        RECT 118.835 99.845 119.155 100.205 ;
        RECT 117.495 99.675 119.155 99.845 ;
        RECT 115.385 98.675 115.595 99.575 ;
        RECT 115.765 98.845 116.455 99.405 ;
        RECT 116.685 98.965 117.185 99.425 ;
        RECT 117.355 99.135 117.965 99.465 ;
        RECT 118.145 99.215 118.475 99.385 ;
        RECT 118.145 98.965 118.470 99.215 ;
        RECT 116.685 98.785 118.470 98.965 ;
        RECT 115.385 98.455 116.340 98.675 ;
        RECT 115.615 97.825 115.885 98.285 ;
        RECT 116.055 97.995 116.340 98.455 ;
        RECT 116.650 98.435 118.685 98.605 ;
        RECT 116.650 98.355 117.760 98.435 ;
        RECT 116.650 97.995 116.910 98.355 ;
        RECT 117.080 97.825 117.410 98.185 ;
        RECT 117.590 97.995 117.760 98.355 ;
        RECT 118.015 97.825 118.185 98.265 ;
        RECT 118.355 98.175 118.685 98.435 ;
        RECT 118.855 98.345 119.155 99.675 ;
        RECT 119.335 99.635 119.665 100.375 ;
        RECT 119.845 99.635 120.285 100.195 ;
        RECT 120.455 99.635 120.905 100.375 ;
        RECT 121.075 99.805 121.245 100.205 ;
        RECT 121.415 99.975 121.835 100.375 ;
        RECT 122.005 99.805 122.235 100.205 ;
        RECT 121.075 99.635 122.235 99.805 ;
        RECT 122.405 99.635 122.895 100.205 ;
        RECT 119.340 98.835 119.615 99.465 ;
        RECT 119.325 98.175 119.630 98.665 ;
        RECT 118.355 97.995 119.630 98.175 ;
        RECT 119.845 98.625 120.155 99.635 ;
        RECT 120.325 99.015 120.495 99.465 ;
        RECT 120.665 99.185 121.055 99.465 ;
        RECT 121.240 99.135 121.485 99.465 ;
        RECT 120.325 98.845 121.115 99.015 ;
        RECT 119.845 97.995 120.285 98.625 ;
        RECT 120.460 97.825 120.775 98.675 ;
        RECT 120.945 98.165 121.115 98.845 ;
        RECT 121.285 98.335 121.485 99.135 ;
        RECT 121.685 98.335 121.935 99.465 ;
        RECT 122.150 99.135 122.555 99.465 ;
        RECT 122.725 98.965 122.895 99.635 ;
        RECT 122.125 98.795 122.895 98.965 ;
        RECT 123.065 99.915 123.625 100.205 ;
        RECT 123.795 99.915 124.045 100.375 ;
        RECT 122.125 98.165 122.375 98.795 ;
        RECT 120.945 97.995 122.375 98.165 ;
        RECT 122.555 97.825 122.885 98.625 ;
        RECT 123.065 98.545 123.315 99.915 ;
        RECT 124.665 99.745 124.995 100.105 ;
        RECT 123.605 99.555 124.995 99.745 ;
        RECT 125.825 99.650 126.115 100.375 ;
        RECT 126.285 99.605 127.955 100.375 ;
        RECT 128.675 99.825 128.845 100.205 ;
        RECT 129.060 99.995 129.390 100.375 ;
        RECT 128.675 99.655 129.390 99.825 ;
        RECT 123.605 99.465 123.775 99.555 ;
        RECT 123.485 99.135 123.775 99.465 ;
        RECT 123.945 99.135 124.285 99.385 ;
        RECT 124.505 99.135 125.180 99.385 ;
        RECT 123.605 98.885 123.775 99.135 ;
        RECT 123.605 98.715 124.545 98.885 ;
        RECT 124.915 98.775 125.180 99.135 ;
        RECT 126.285 99.085 127.035 99.605 ;
        RECT 123.065 97.995 123.525 98.545 ;
        RECT 123.715 97.825 124.045 98.545 ;
        RECT 124.245 98.165 124.545 98.715 ;
        RECT 124.715 97.825 124.995 98.495 ;
        RECT 125.825 97.825 126.115 98.990 ;
        RECT 127.205 98.915 127.955 99.435 ;
        RECT 128.585 99.105 128.940 99.475 ;
        RECT 129.220 99.465 129.390 99.655 ;
        RECT 129.560 99.630 129.815 100.205 ;
        RECT 129.220 99.135 129.475 99.465 ;
        RECT 129.220 98.925 129.390 99.135 ;
        RECT 126.285 97.825 127.955 98.915 ;
        RECT 128.675 98.755 129.390 98.925 ;
        RECT 129.645 98.900 129.815 99.630 ;
        RECT 129.990 99.535 130.250 100.375 ;
        RECT 130.425 99.605 133.015 100.375 ;
        RECT 133.235 99.720 133.565 100.155 ;
        RECT 133.735 99.765 133.905 100.375 ;
        RECT 133.185 99.635 133.565 99.720 ;
        RECT 134.075 99.635 134.405 100.160 ;
        RECT 134.665 99.845 134.875 100.375 ;
        RECT 135.150 99.925 135.935 100.095 ;
        RECT 136.105 99.925 136.510 100.095 ;
        RECT 130.425 99.085 131.635 99.605 ;
        RECT 133.185 99.595 133.410 99.635 ;
        RECT 128.675 97.995 128.845 98.755 ;
        RECT 129.060 97.825 129.390 98.585 ;
        RECT 129.560 97.995 129.815 98.900 ;
        RECT 129.990 97.825 130.250 98.975 ;
        RECT 131.805 98.915 133.015 99.435 ;
        RECT 130.425 97.825 133.015 98.915 ;
        RECT 133.185 99.015 133.355 99.595 ;
        RECT 134.075 99.465 134.275 99.635 ;
        RECT 135.150 99.465 135.320 99.925 ;
        RECT 133.525 99.135 134.275 99.465 ;
        RECT 134.445 99.135 135.320 99.465 ;
        RECT 133.185 98.965 133.400 99.015 ;
        RECT 133.185 98.885 133.575 98.965 ;
        RECT 133.245 98.040 133.575 98.885 ;
        RECT 134.085 98.930 134.275 99.135 ;
        RECT 133.745 97.825 133.915 98.835 ;
        RECT 134.085 98.555 134.980 98.930 ;
        RECT 134.085 97.995 134.425 98.555 ;
        RECT 134.655 97.825 134.970 98.325 ;
        RECT 135.150 98.295 135.320 99.135 ;
        RECT 135.490 99.425 135.955 99.755 ;
        RECT 136.340 99.695 136.510 99.925 ;
        RECT 136.690 99.875 137.060 100.375 ;
        RECT 137.380 99.925 138.055 100.095 ;
        RECT 138.250 99.925 138.585 100.095 ;
        RECT 135.490 98.465 135.810 99.425 ;
        RECT 136.340 99.395 137.170 99.695 ;
        RECT 135.980 98.495 136.170 99.215 ;
        RECT 136.340 98.325 136.510 99.395 ;
        RECT 136.970 99.365 137.170 99.395 ;
        RECT 136.680 99.145 136.850 99.215 ;
        RECT 137.380 99.145 137.550 99.925 ;
        RECT 138.415 99.785 138.585 99.925 ;
        RECT 138.755 99.915 139.005 100.375 ;
        RECT 136.680 98.975 137.550 99.145 ;
        RECT 137.720 99.505 138.245 99.725 ;
        RECT 138.415 99.655 138.640 99.785 ;
        RECT 136.680 98.885 137.190 98.975 ;
        RECT 135.150 98.125 136.035 98.295 ;
        RECT 136.260 97.995 136.510 98.325 ;
        RECT 136.680 97.825 136.850 98.625 ;
        RECT 137.020 98.270 137.190 98.885 ;
        RECT 137.720 98.805 137.890 99.505 ;
        RECT 137.360 98.440 137.890 98.805 ;
        RECT 138.060 98.740 138.300 99.335 ;
        RECT 138.470 98.550 138.640 99.655 ;
        RECT 138.810 98.795 139.090 99.745 ;
        RECT 138.335 98.420 138.640 98.550 ;
        RECT 137.020 98.100 138.125 98.270 ;
        RECT 138.335 97.995 138.585 98.420 ;
        RECT 138.755 97.825 139.020 98.285 ;
        RECT 139.260 97.995 139.445 100.115 ;
        RECT 139.615 99.995 139.945 100.375 ;
        RECT 140.115 99.825 140.285 100.115 ;
        RECT 139.620 99.655 140.285 99.825 ;
        RECT 139.620 98.665 139.850 99.655 ;
        RECT 140.750 99.595 141.250 100.205 ;
        RECT 140.020 98.835 140.370 99.485 ;
        RECT 140.545 99.135 140.895 99.385 ;
        RECT 141.080 98.965 141.250 99.595 ;
        RECT 141.880 99.725 142.210 100.205 ;
        RECT 142.380 99.915 142.605 100.375 ;
        RECT 142.775 99.725 143.105 100.205 ;
        RECT 141.880 99.555 143.105 99.725 ;
        RECT 143.295 99.575 143.545 100.375 ;
        RECT 143.715 99.575 144.055 100.205 ;
        RECT 144.340 99.745 144.625 100.205 ;
        RECT 144.795 99.915 145.065 100.375 ;
        RECT 144.340 99.575 145.295 99.745 ;
        RECT 141.420 99.185 141.750 99.385 ;
        RECT 141.920 99.185 142.250 99.385 ;
        RECT 142.420 99.185 142.840 99.385 ;
        RECT 143.015 99.215 143.710 99.385 ;
        RECT 143.015 98.965 143.185 99.215 ;
        RECT 143.880 99.015 144.055 99.575 ;
        RECT 143.825 98.965 144.055 99.015 ;
        RECT 140.750 98.795 143.185 98.965 ;
        RECT 139.620 98.495 140.285 98.665 ;
        RECT 139.615 97.825 139.945 98.325 ;
        RECT 140.115 97.995 140.285 98.495 ;
        RECT 140.750 97.995 141.080 98.795 ;
        RECT 141.250 97.825 141.580 98.625 ;
        RECT 141.880 97.995 142.210 98.795 ;
        RECT 142.855 97.825 143.105 98.625 ;
        RECT 143.375 97.825 143.545 98.965 ;
        RECT 143.715 97.995 144.055 98.965 ;
        RECT 144.225 98.845 144.915 99.405 ;
        RECT 145.085 98.675 145.295 99.575 ;
        RECT 144.340 98.455 145.295 98.675 ;
        RECT 145.465 99.405 145.865 100.205 ;
        RECT 146.055 99.745 146.335 100.205 ;
        RECT 146.855 99.915 147.180 100.375 ;
        RECT 146.055 99.575 147.180 99.745 ;
        RECT 147.350 99.635 147.735 100.205 ;
        RECT 146.730 99.465 147.180 99.575 ;
        RECT 145.465 98.845 146.560 99.405 ;
        RECT 146.730 99.135 147.285 99.465 ;
        RECT 144.340 97.995 144.625 98.455 ;
        RECT 144.795 97.825 145.065 98.285 ;
        RECT 145.465 97.995 145.865 98.845 ;
        RECT 146.730 98.675 147.180 99.135 ;
        RECT 147.455 98.965 147.735 99.635 ;
        RECT 146.055 98.455 147.180 98.675 ;
        RECT 146.055 97.995 146.335 98.455 ;
        RECT 146.855 97.825 147.180 98.285 ;
        RECT 147.350 97.995 147.735 98.965 ;
        RECT 147.905 99.575 148.245 100.205 ;
        RECT 148.415 99.575 148.665 100.375 ;
        RECT 148.855 99.725 149.185 100.205 ;
        RECT 149.355 99.915 149.580 100.375 ;
        RECT 149.750 99.725 150.080 100.205 ;
        RECT 147.905 98.965 148.080 99.575 ;
        RECT 148.855 99.555 150.080 99.725 ;
        RECT 150.710 99.595 151.210 100.205 ;
        RECT 151.585 99.650 151.875 100.375 ;
        RECT 152.045 99.635 152.430 100.205 ;
        RECT 152.600 99.915 152.925 100.375 ;
        RECT 153.445 99.745 153.725 100.205 ;
        RECT 148.250 99.215 148.945 99.385 ;
        RECT 148.775 98.965 148.945 99.215 ;
        RECT 149.120 99.185 149.540 99.385 ;
        RECT 149.710 99.185 150.040 99.385 ;
        RECT 150.210 99.185 150.540 99.385 ;
        RECT 150.710 98.965 150.880 99.595 ;
        RECT 151.065 99.135 151.415 99.385 ;
        RECT 147.905 97.995 148.245 98.965 ;
        RECT 148.415 97.825 148.585 98.965 ;
        RECT 148.775 98.795 151.210 98.965 ;
        RECT 148.855 97.825 149.105 98.625 ;
        RECT 149.750 97.995 150.080 98.795 ;
        RECT 150.380 97.825 150.710 98.625 ;
        RECT 150.880 97.995 151.210 98.795 ;
        RECT 151.585 97.825 151.875 98.990 ;
        RECT 152.045 98.965 152.325 99.635 ;
        RECT 152.600 99.575 153.725 99.745 ;
        RECT 152.600 99.465 153.050 99.575 ;
        RECT 152.495 99.135 153.050 99.465 ;
        RECT 153.915 99.405 154.315 100.205 ;
        RECT 154.715 99.915 154.985 100.375 ;
        RECT 155.155 99.745 155.440 100.205 ;
        RECT 152.045 97.995 152.430 98.965 ;
        RECT 152.600 98.675 153.050 99.135 ;
        RECT 153.220 98.845 154.315 99.405 ;
        RECT 152.600 98.455 153.725 98.675 ;
        RECT 152.600 97.825 152.925 98.285 ;
        RECT 153.445 97.995 153.725 98.455 ;
        RECT 153.915 97.995 154.315 98.845 ;
        RECT 154.485 99.575 155.440 99.745 ;
        RECT 155.725 99.625 156.935 100.375 ;
        RECT 154.485 98.675 154.695 99.575 ;
        RECT 154.865 98.845 155.555 99.405 ;
        RECT 155.725 98.915 156.245 99.455 ;
        RECT 156.415 99.085 156.935 99.625 ;
        RECT 154.485 98.455 155.440 98.675 ;
        RECT 154.715 97.825 154.985 98.285 ;
        RECT 155.155 97.995 155.440 98.455 ;
        RECT 155.725 97.825 156.935 98.915 ;
        RECT 22.700 97.655 157.020 97.825 ;
        RECT 22.785 96.565 23.995 97.655 ;
        RECT 24.165 96.565 25.375 97.655 ;
        RECT 22.785 95.855 23.305 96.395 ;
        RECT 23.475 96.025 23.995 96.565 ;
        RECT 24.165 95.855 24.685 96.395 ;
        RECT 24.855 96.025 25.375 96.565 ;
        RECT 25.545 96.580 25.815 97.485 ;
        RECT 25.985 96.895 26.315 97.655 ;
        RECT 26.495 96.725 26.665 97.485 ;
        RECT 22.785 95.105 23.995 95.855 ;
        RECT 24.165 95.105 25.375 95.855 ;
        RECT 25.545 95.780 25.715 96.580 ;
        RECT 26.000 96.555 26.665 96.725 ;
        RECT 26.925 96.565 29.515 97.655 ;
        RECT 26.000 96.410 26.170 96.555 ;
        RECT 25.885 96.080 26.170 96.410 ;
        RECT 26.000 95.825 26.170 96.080 ;
        RECT 26.405 96.005 26.735 96.375 ;
        RECT 26.925 95.875 28.135 96.395 ;
        RECT 28.305 96.045 29.515 96.565 ;
        RECT 29.715 96.555 30.090 97.655 ;
        RECT 30.565 96.645 30.890 97.485 ;
        RECT 31.060 96.895 31.390 97.655 ;
        RECT 31.560 96.725 31.835 97.230 ;
        RECT 30.565 96.475 31.175 96.645 ;
        RECT 29.685 96.095 30.165 96.305 ;
        RECT 30.335 96.095 30.835 96.305 ;
        RECT 25.545 95.275 25.805 95.780 ;
        RECT 26.000 95.655 26.665 95.825 ;
        RECT 25.985 95.105 26.315 95.485 ;
        RECT 26.495 95.275 26.665 95.655 ;
        RECT 26.925 95.105 29.515 95.875 ;
        RECT 29.695 95.755 30.790 95.925 ;
        RECT 29.695 95.290 30.025 95.755 ;
        RECT 30.195 95.105 30.365 95.575 ;
        RECT 30.620 95.505 30.790 95.755 ;
        RECT 31.005 95.845 31.175 96.475 ;
        RECT 31.345 96.555 31.835 96.725 ;
        RECT 31.345 96.015 31.640 96.555 ;
        RECT 32.005 96.365 32.275 97.465 ;
        RECT 31.825 96.015 32.275 96.365 ;
        RECT 32.445 96.515 32.720 97.485 ;
        RECT 32.930 96.855 33.210 97.655 ;
        RECT 33.380 97.145 34.995 97.475 ;
        RECT 33.380 96.805 34.555 96.975 ;
        RECT 33.380 96.685 33.550 96.805 ;
        RECT 32.890 96.515 33.550 96.685 ;
        RECT 31.470 95.845 31.640 96.015 ;
        RECT 31.005 95.665 31.245 95.845 ;
        RECT 31.470 95.675 31.780 95.845 ;
        RECT 30.540 95.275 30.870 95.505 ;
        RECT 31.075 95.275 31.245 95.665 ;
        RECT 31.590 95.515 31.780 95.675 ;
        RECT 32.000 95.105 32.275 95.845 ;
        RECT 32.445 95.780 32.615 96.515 ;
        RECT 32.890 96.345 33.060 96.515 ;
        RECT 33.810 96.345 34.055 96.635 ;
        RECT 34.225 96.515 34.555 96.805 ;
        RECT 34.815 96.345 34.985 96.905 ;
        RECT 35.235 96.515 35.495 97.655 ;
        RECT 35.665 96.490 35.955 97.655 ;
        RECT 37.135 96.985 37.305 97.485 ;
        RECT 37.475 97.155 37.805 97.655 ;
        RECT 37.135 96.815 37.800 96.985 ;
        RECT 32.785 96.015 33.060 96.345 ;
        RECT 33.230 96.015 34.055 96.345 ;
        RECT 34.270 96.015 34.985 96.345 ;
        RECT 35.155 96.095 35.490 96.345 ;
        RECT 32.890 95.845 33.060 96.015 ;
        RECT 34.735 95.925 34.985 96.015 ;
        RECT 37.050 95.995 37.400 96.645 ;
        RECT 32.445 95.435 32.720 95.780 ;
        RECT 32.890 95.675 34.555 95.845 ;
        RECT 32.910 95.105 33.285 95.505 ;
        RECT 33.455 95.325 33.625 95.675 ;
        RECT 33.795 95.105 34.125 95.505 ;
        RECT 34.295 95.275 34.555 95.675 ;
        RECT 34.735 95.505 35.065 95.925 ;
        RECT 35.235 95.105 35.495 95.925 ;
        RECT 35.665 95.105 35.955 95.830 ;
        RECT 37.570 95.825 37.800 96.815 ;
        RECT 37.135 95.655 37.800 95.825 ;
        RECT 37.135 95.365 37.305 95.655 ;
        RECT 37.475 95.105 37.805 95.485 ;
        RECT 37.975 95.365 38.160 97.485 ;
        RECT 38.400 97.195 38.665 97.655 ;
        RECT 38.835 97.060 39.085 97.485 ;
        RECT 39.295 97.210 40.400 97.380 ;
        RECT 38.780 96.930 39.085 97.060 ;
        RECT 38.330 95.735 38.610 96.685 ;
        RECT 38.780 95.825 38.950 96.930 ;
        RECT 39.120 96.145 39.360 96.740 ;
        RECT 39.530 96.675 40.060 97.040 ;
        RECT 39.530 95.975 39.700 96.675 ;
        RECT 40.230 96.595 40.400 97.210 ;
        RECT 40.570 96.855 40.740 97.655 ;
        RECT 40.910 97.155 41.160 97.485 ;
        RECT 41.385 97.185 42.270 97.355 ;
        RECT 40.230 96.505 40.740 96.595 ;
        RECT 38.780 95.695 39.005 95.825 ;
        RECT 39.175 95.755 39.700 95.975 ;
        RECT 39.870 96.335 40.740 96.505 ;
        RECT 38.415 95.105 38.665 95.565 ;
        RECT 38.835 95.555 39.005 95.695 ;
        RECT 39.870 95.555 40.040 96.335 ;
        RECT 40.570 96.265 40.740 96.335 ;
        RECT 40.250 96.085 40.450 96.115 ;
        RECT 40.910 96.085 41.080 97.155 ;
        RECT 41.250 96.265 41.440 96.985 ;
        RECT 40.250 95.785 41.080 96.085 ;
        RECT 41.610 96.055 41.930 97.015 ;
        RECT 38.835 95.385 39.170 95.555 ;
        RECT 39.365 95.385 40.040 95.555 ;
        RECT 40.360 95.105 40.730 95.605 ;
        RECT 40.910 95.555 41.080 95.785 ;
        RECT 41.465 95.725 41.930 96.055 ;
        RECT 42.100 96.345 42.270 97.185 ;
        RECT 42.450 97.155 42.765 97.655 ;
        RECT 42.995 96.925 43.335 97.485 ;
        RECT 42.440 96.550 43.335 96.925 ;
        RECT 43.505 96.645 43.675 97.655 ;
        RECT 43.145 96.345 43.335 96.550 ;
        RECT 43.845 96.595 44.175 97.440 ;
        RECT 44.495 96.985 44.665 97.485 ;
        RECT 44.835 97.155 45.165 97.655 ;
        RECT 44.495 96.815 45.160 96.985 ;
        RECT 43.845 96.515 44.235 96.595 ;
        RECT 44.020 96.465 44.235 96.515 ;
        RECT 42.100 96.015 42.975 96.345 ;
        RECT 43.145 96.015 43.895 96.345 ;
        RECT 42.100 95.555 42.270 96.015 ;
        RECT 43.145 95.845 43.345 96.015 ;
        RECT 44.065 95.885 44.235 96.465 ;
        RECT 44.410 95.995 44.760 96.645 ;
        RECT 44.010 95.845 44.235 95.885 ;
        RECT 40.910 95.385 41.315 95.555 ;
        RECT 41.485 95.385 42.270 95.555 ;
        RECT 42.545 95.105 42.755 95.635 ;
        RECT 43.015 95.320 43.345 95.845 ;
        RECT 43.855 95.760 44.235 95.845 ;
        RECT 44.930 95.825 45.160 96.815 ;
        RECT 43.515 95.105 43.685 95.715 ;
        RECT 43.855 95.325 44.185 95.760 ;
        RECT 44.495 95.655 45.160 95.825 ;
        RECT 44.495 95.365 44.665 95.655 ;
        RECT 44.835 95.105 45.165 95.485 ;
        RECT 45.335 95.365 45.520 97.485 ;
        RECT 45.760 97.195 46.025 97.655 ;
        RECT 46.195 97.060 46.445 97.485 ;
        RECT 46.655 97.210 47.760 97.380 ;
        RECT 46.140 96.930 46.445 97.060 ;
        RECT 45.690 95.735 45.970 96.685 ;
        RECT 46.140 95.825 46.310 96.930 ;
        RECT 46.480 96.145 46.720 96.740 ;
        RECT 46.890 96.675 47.420 97.040 ;
        RECT 46.890 95.975 47.060 96.675 ;
        RECT 47.590 96.595 47.760 97.210 ;
        RECT 47.930 96.855 48.100 97.655 ;
        RECT 48.270 97.155 48.520 97.485 ;
        RECT 48.745 97.185 49.630 97.355 ;
        RECT 47.590 96.505 48.100 96.595 ;
        RECT 46.140 95.695 46.365 95.825 ;
        RECT 46.535 95.755 47.060 95.975 ;
        RECT 47.230 96.335 48.100 96.505 ;
        RECT 45.775 95.105 46.025 95.565 ;
        RECT 46.195 95.555 46.365 95.695 ;
        RECT 47.230 95.555 47.400 96.335 ;
        RECT 47.930 96.265 48.100 96.335 ;
        RECT 47.610 96.085 47.810 96.115 ;
        RECT 48.270 96.085 48.440 97.155 ;
        RECT 48.610 96.265 48.800 96.985 ;
        RECT 47.610 95.785 48.440 96.085 ;
        RECT 48.970 96.055 49.290 97.015 ;
        RECT 46.195 95.385 46.530 95.555 ;
        RECT 46.725 95.385 47.400 95.555 ;
        RECT 47.720 95.105 48.090 95.605 ;
        RECT 48.270 95.555 48.440 95.785 ;
        RECT 48.825 95.725 49.290 96.055 ;
        RECT 49.460 96.345 49.630 97.185 ;
        RECT 49.810 97.155 50.125 97.655 ;
        RECT 50.355 96.925 50.695 97.485 ;
        RECT 49.800 96.550 50.695 96.925 ;
        RECT 50.865 96.645 51.035 97.655 ;
        RECT 50.505 96.345 50.695 96.550 ;
        RECT 51.205 96.595 51.535 97.440 ;
        RECT 51.205 96.515 51.595 96.595 ;
        RECT 51.765 96.565 55.275 97.655 ;
        RECT 51.380 96.465 51.595 96.515 ;
        RECT 49.460 96.015 50.335 96.345 ;
        RECT 50.505 96.015 51.255 96.345 ;
        RECT 49.460 95.555 49.630 96.015 ;
        RECT 50.505 95.845 50.705 96.015 ;
        RECT 51.425 95.885 51.595 96.465 ;
        RECT 51.370 95.845 51.595 95.885 ;
        RECT 48.270 95.385 48.675 95.555 ;
        RECT 48.845 95.385 49.630 95.555 ;
        RECT 49.905 95.105 50.115 95.635 ;
        RECT 50.375 95.320 50.705 95.845 ;
        RECT 51.215 95.760 51.595 95.845 ;
        RECT 51.765 95.875 53.415 96.395 ;
        RECT 53.585 96.045 55.275 96.565 ;
        RECT 55.535 96.725 55.705 97.485 ;
        RECT 55.885 96.895 56.215 97.655 ;
        RECT 55.535 96.555 56.200 96.725 ;
        RECT 56.385 96.580 56.655 97.485 ;
        RECT 56.030 96.410 56.200 96.555 ;
        RECT 55.465 96.005 55.795 96.375 ;
        RECT 56.030 96.080 56.315 96.410 ;
        RECT 50.875 95.105 51.045 95.715 ;
        RECT 51.215 95.325 51.545 95.760 ;
        RECT 51.765 95.105 55.275 95.875 ;
        RECT 56.030 95.825 56.200 96.080 ;
        RECT 55.535 95.655 56.200 95.825 ;
        RECT 56.485 95.780 56.655 96.580 ;
        RECT 56.825 96.565 60.335 97.655 ;
        RECT 55.535 95.275 55.705 95.655 ;
        RECT 55.885 95.105 56.215 95.485 ;
        RECT 56.395 95.275 56.655 95.780 ;
        RECT 56.825 95.875 58.475 96.395 ;
        RECT 58.645 96.045 60.335 96.565 ;
        RECT 61.425 96.490 61.715 97.655 ;
        RECT 61.885 96.565 65.395 97.655 ;
        RECT 65.610 97.305 66.885 97.485 ;
        RECT 65.610 96.815 65.915 97.305 ;
        RECT 61.885 95.875 63.535 96.395 ;
        RECT 63.705 96.045 65.395 96.565 ;
        RECT 65.625 96.015 65.900 96.645 ;
        RECT 56.825 95.105 60.335 95.875 ;
        RECT 61.425 95.105 61.715 95.830 ;
        RECT 61.885 95.105 65.395 95.875 ;
        RECT 65.575 95.105 65.905 95.845 ;
        RECT 66.085 95.805 66.385 97.135 ;
        RECT 66.555 97.045 66.885 97.305 ;
        RECT 67.055 97.215 67.225 97.655 ;
        RECT 67.480 97.125 67.650 97.485 ;
        RECT 67.830 97.295 68.160 97.655 ;
        RECT 68.330 97.125 68.590 97.485 ;
        RECT 67.480 97.045 68.590 97.125 ;
        RECT 66.555 96.875 68.590 97.045 ;
        RECT 68.900 97.025 69.185 97.485 ;
        RECT 69.355 97.195 69.625 97.655 ;
        RECT 68.900 96.805 69.855 97.025 ;
        RECT 66.770 96.515 68.555 96.695 ;
        RECT 66.770 96.265 67.095 96.515 ;
        RECT 66.765 96.095 67.095 96.265 ;
        RECT 67.275 96.015 67.885 96.345 ;
        RECT 68.055 96.055 68.555 96.515 ;
        RECT 68.785 96.075 69.475 96.635 ;
        RECT 69.645 95.905 69.855 96.805 ;
        RECT 66.085 95.635 67.745 95.805 ;
        RECT 66.085 95.275 66.405 95.635 ;
        RECT 66.610 95.105 66.940 95.465 ;
        RECT 67.400 95.275 67.745 95.635 ;
        RECT 68.305 95.105 68.600 95.885 ;
        RECT 68.900 95.735 69.855 95.905 ;
        RECT 70.025 96.635 70.425 97.485 ;
        RECT 70.615 97.025 70.895 97.485 ;
        RECT 71.415 97.195 71.740 97.655 ;
        RECT 70.615 96.805 71.740 97.025 ;
        RECT 70.025 96.075 71.120 96.635 ;
        RECT 71.290 96.345 71.740 96.805 ;
        RECT 71.910 96.515 72.295 97.485 ;
        RECT 72.475 96.545 72.770 97.655 ;
        RECT 68.900 95.275 69.185 95.735 ;
        RECT 69.355 95.105 69.625 95.565 ;
        RECT 70.025 95.275 70.425 96.075 ;
        RECT 71.290 96.015 71.845 96.345 ;
        RECT 71.290 95.905 71.740 96.015 ;
        RECT 70.615 95.735 71.740 95.905 ;
        RECT 72.015 95.845 72.295 96.515 ;
        RECT 72.950 96.345 73.200 97.480 ;
        RECT 73.370 96.545 73.630 97.655 ;
        RECT 73.800 96.755 74.060 97.480 ;
        RECT 74.230 96.925 74.490 97.655 ;
        RECT 74.660 96.755 74.920 97.480 ;
        RECT 75.090 96.925 75.350 97.655 ;
        RECT 75.520 96.755 75.780 97.480 ;
        RECT 75.950 96.925 76.210 97.655 ;
        RECT 76.380 96.755 76.640 97.480 ;
        RECT 76.810 96.925 77.105 97.655 ;
        RECT 78.445 96.785 78.720 97.485 ;
        RECT 78.890 97.110 79.145 97.655 ;
        RECT 79.315 97.145 79.795 97.485 ;
        RECT 79.970 97.100 80.575 97.655 ;
        RECT 79.960 97.000 80.575 97.100 ;
        RECT 79.960 96.975 80.145 97.000 ;
        RECT 73.800 96.515 77.110 96.755 ;
        RECT 70.615 95.275 70.895 95.735 ;
        RECT 71.415 95.105 71.740 95.565 ;
        RECT 71.910 95.275 72.295 95.845 ;
        RECT 72.465 95.735 72.780 96.345 ;
        RECT 72.950 96.095 75.970 96.345 ;
        RECT 72.525 95.105 72.770 95.565 ;
        RECT 72.950 95.285 73.200 96.095 ;
        RECT 76.140 95.925 77.110 96.515 ;
        RECT 73.800 95.755 77.110 95.925 ;
        RECT 78.445 95.755 78.615 96.785 ;
        RECT 78.890 96.655 79.645 96.905 ;
        RECT 79.815 96.730 80.145 96.975 ;
        RECT 78.890 96.620 79.660 96.655 ;
        RECT 78.890 96.610 79.675 96.620 ;
        RECT 78.785 96.595 79.680 96.610 ;
        RECT 78.785 96.580 79.700 96.595 ;
        RECT 78.785 96.570 79.720 96.580 ;
        RECT 78.785 96.560 79.745 96.570 ;
        RECT 78.785 96.530 79.815 96.560 ;
        RECT 78.785 96.500 79.835 96.530 ;
        RECT 78.785 96.470 79.855 96.500 ;
        RECT 78.785 96.445 79.885 96.470 ;
        RECT 78.785 96.410 79.920 96.445 ;
        RECT 78.785 96.405 79.950 96.410 ;
        RECT 78.785 96.010 79.015 96.405 ;
        RECT 79.560 96.400 79.950 96.405 ;
        RECT 79.585 96.390 79.950 96.400 ;
        RECT 79.600 96.385 79.950 96.390 ;
        RECT 79.615 96.380 79.950 96.385 ;
        RECT 80.315 96.380 80.575 96.830 ;
        RECT 79.615 96.375 80.575 96.380 ;
        RECT 79.625 96.365 80.575 96.375 ;
        RECT 79.635 96.360 80.575 96.365 ;
        RECT 79.645 96.350 80.575 96.360 ;
        RECT 79.650 96.340 80.575 96.350 ;
        RECT 79.655 96.335 80.575 96.340 ;
        RECT 79.665 96.320 80.575 96.335 ;
        RECT 79.670 96.305 80.575 96.320 ;
        RECT 79.680 96.280 80.575 96.305 ;
        RECT 79.185 95.810 79.515 96.235 ;
        RECT 73.370 95.105 73.630 95.630 ;
        RECT 73.800 95.300 74.060 95.755 ;
        RECT 74.230 95.105 74.490 95.585 ;
        RECT 74.660 95.300 74.920 95.755 ;
        RECT 75.090 95.105 75.350 95.585 ;
        RECT 75.520 95.300 75.780 95.755 ;
        RECT 75.950 95.105 76.210 95.585 ;
        RECT 76.380 95.300 76.640 95.755 ;
        RECT 76.810 95.105 77.110 95.585 ;
        RECT 78.445 95.275 78.705 95.755 ;
        RECT 78.875 95.105 79.125 95.645 ;
        RECT 79.295 95.325 79.515 95.810 ;
        RECT 79.685 96.210 80.575 96.280 ;
        RECT 80.745 96.515 81.130 97.485 ;
        RECT 81.300 97.195 81.625 97.655 ;
        RECT 82.145 97.025 82.425 97.485 ;
        RECT 81.300 96.805 82.425 97.025 ;
        RECT 79.685 95.485 79.855 96.210 ;
        RECT 80.025 95.655 80.575 96.040 ;
        RECT 80.745 95.845 81.025 96.515 ;
        RECT 81.300 96.345 81.750 96.805 ;
        RECT 82.615 96.635 83.015 97.485 ;
        RECT 83.415 97.195 83.685 97.655 ;
        RECT 83.855 97.025 84.140 97.485 ;
        RECT 81.195 96.015 81.750 96.345 ;
        RECT 81.920 96.075 83.015 96.635 ;
        RECT 81.300 95.905 81.750 96.015 ;
        RECT 79.685 95.315 80.575 95.485 ;
        RECT 80.745 95.275 81.130 95.845 ;
        RECT 81.300 95.735 82.425 95.905 ;
        RECT 81.300 95.105 81.625 95.565 ;
        RECT 82.145 95.275 82.425 95.735 ;
        RECT 82.615 95.275 83.015 96.075 ;
        RECT 83.185 96.805 84.140 97.025 ;
        RECT 83.185 95.905 83.395 96.805 ;
        RECT 84.435 96.685 84.765 97.470 ;
        RECT 83.565 96.075 84.255 96.635 ;
        RECT 84.435 96.515 85.115 96.685 ;
        RECT 85.295 96.515 85.625 97.655 ;
        RECT 85.805 96.565 87.015 97.655 ;
        RECT 84.425 96.095 84.775 96.345 ;
        RECT 84.945 95.915 85.115 96.515 ;
        RECT 85.285 96.095 85.635 96.345 ;
        RECT 83.185 95.735 84.140 95.905 ;
        RECT 83.415 95.105 83.685 95.565 ;
        RECT 83.855 95.275 84.140 95.735 ;
        RECT 84.445 95.105 84.685 95.915 ;
        RECT 84.855 95.275 85.185 95.915 ;
        RECT 85.355 95.105 85.625 95.915 ;
        RECT 85.805 95.855 86.325 96.395 ;
        RECT 86.495 96.025 87.015 96.565 ;
        RECT 87.185 96.490 87.475 97.655 ;
        RECT 87.645 96.565 89.315 97.655 ;
        RECT 89.945 97.100 90.550 97.655 ;
        RECT 90.725 97.145 91.205 97.485 ;
        RECT 91.375 97.110 91.630 97.655 ;
        RECT 89.945 97.000 90.560 97.100 ;
        RECT 90.375 96.975 90.560 97.000 ;
        RECT 87.645 95.875 88.395 96.395 ;
        RECT 88.565 96.045 89.315 96.565 ;
        RECT 89.945 96.380 90.205 96.830 ;
        RECT 90.375 96.730 90.705 96.975 ;
        RECT 90.875 96.655 91.630 96.905 ;
        RECT 91.800 96.785 92.075 97.485 ;
        RECT 90.860 96.620 91.630 96.655 ;
        RECT 90.845 96.610 91.630 96.620 ;
        RECT 90.840 96.595 91.735 96.610 ;
        RECT 90.820 96.580 91.735 96.595 ;
        RECT 90.800 96.570 91.735 96.580 ;
        RECT 90.775 96.560 91.735 96.570 ;
        RECT 90.705 96.530 91.735 96.560 ;
        RECT 90.685 96.500 91.735 96.530 ;
        RECT 90.665 96.470 91.735 96.500 ;
        RECT 90.635 96.445 91.735 96.470 ;
        RECT 90.600 96.410 91.735 96.445 ;
        RECT 90.570 96.405 91.735 96.410 ;
        RECT 90.570 96.400 90.960 96.405 ;
        RECT 90.570 96.390 90.935 96.400 ;
        RECT 90.570 96.385 90.920 96.390 ;
        RECT 90.570 96.380 90.905 96.385 ;
        RECT 89.945 96.375 90.905 96.380 ;
        RECT 89.945 96.365 90.895 96.375 ;
        RECT 89.945 96.360 90.885 96.365 ;
        RECT 89.945 96.350 90.875 96.360 ;
        RECT 89.945 96.340 90.870 96.350 ;
        RECT 89.945 96.335 90.865 96.340 ;
        RECT 89.945 96.320 90.855 96.335 ;
        RECT 89.945 96.305 90.850 96.320 ;
        RECT 89.945 96.280 90.840 96.305 ;
        RECT 89.945 96.210 90.835 96.280 ;
        RECT 85.805 95.105 87.015 95.855 ;
        RECT 87.185 95.105 87.475 95.830 ;
        RECT 87.645 95.105 89.315 95.875 ;
        RECT 89.945 95.655 90.495 96.040 ;
        RECT 90.665 95.485 90.835 96.210 ;
        RECT 89.945 95.315 90.835 95.485 ;
        RECT 91.005 95.810 91.335 96.235 ;
        RECT 91.505 96.010 91.735 96.405 ;
        RECT 91.005 95.785 91.255 95.810 ;
        RECT 91.005 95.325 91.225 95.785 ;
        RECT 91.905 95.755 92.075 96.785 ;
        RECT 92.245 96.565 93.915 97.655 ;
        RECT 91.395 95.105 91.645 95.645 ;
        RECT 91.815 95.275 92.075 95.755 ;
        RECT 92.245 95.875 92.995 96.395 ;
        RECT 93.165 96.045 93.915 96.565 ;
        RECT 94.730 96.685 95.120 96.860 ;
        RECT 95.605 96.855 95.935 97.655 ;
        RECT 96.105 96.865 96.640 97.485 ;
        RECT 94.730 96.515 96.155 96.685 ;
        RECT 92.245 95.105 93.915 95.875 ;
        RECT 94.605 95.785 94.960 96.345 ;
        RECT 95.130 95.615 95.300 96.515 ;
        RECT 95.470 95.785 95.735 96.345 ;
        RECT 95.985 96.015 96.155 96.515 ;
        RECT 96.325 95.845 96.640 96.865 ;
        RECT 96.845 96.515 97.105 97.655 ;
        RECT 97.275 96.505 97.605 97.485 ;
        RECT 97.775 96.515 98.055 97.655 ;
        RECT 98.225 96.565 100.815 97.655 ;
        RECT 96.865 96.095 97.200 96.345 ;
        RECT 97.370 95.905 97.540 96.505 ;
        RECT 97.710 96.075 98.045 96.345 ;
        RECT 94.710 95.105 94.950 95.615 ;
        RECT 95.130 95.285 95.410 95.615 ;
        RECT 95.640 95.105 95.855 95.615 ;
        RECT 96.025 95.275 96.640 95.845 ;
        RECT 96.845 95.275 97.540 95.905 ;
        RECT 97.745 95.105 98.055 95.905 ;
        RECT 98.225 95.875 99.435 96.395 ;
        RECT 99.605 96.045 100.815 96.565 ;
        RECT 101.445 96.580 101.715 97.485 ;
        RECT 101.885 96.895 102.215 97.655 ;
        RECT 102.395 96.725 102.565 97.485 ;
        RECT 98.225 95.105 100.815 95.875 ;
        RECT 101.445 95.780 101.615 96.580 ;
        RECT 101.900 96.555 102.565 96.725 ;
        RECT 102.825 96.565 106.335 97.655 ;
        RECT 101.900 96.410 102.070 96.555 ;
        RECT 101.785 96.080 102.070 96.410 ;
        RECT 101.900 95.825 102.070 96.080 ;
        RECT 102.305 96.005 102.635 96.375 ;
        RECT 102.825 95.875 104.475 96.395 ;
        RECT 104.645 96.045 106.335 96.565 ;
        RECT 107.425 96.580 107.695 97.485 ;
        RECT 107.865 96.895 108.195 97.655 ;
        RECT 108.375 96.725 108.545 97.485 ;
        RECT 101.445 95.275 101.705 95.780 ;
        RECT 101.900 95.655 102.565 95.825 ;
        RECT 101.885 95.105 102.215 95.485 ;
        RECT 102.395 95.275 102.565 95.655 ;
        RECT 102.825 95.105 106.335 95.875 ;
        RECT 107.425 95.780 107.595 96.580 ;
        RECT 107.880 96.555 108.545 96.725 ;
        RECT 109.285 96.600 109.590 97.385 ;
        RECT 109.770 97.185 110.455 97.655 ;
        RECT 109.765 96.665 110.460 96.975 ;
        RECT 107.880 96.410 108.050 96.555 ;
        RECT 107.765 96.080 108.050 96.410 ;
        RECT 109.285 96.465 109.495 96.600 ;
        RECT 110.635 96.495 110.920 97.440 ;
        RECT 111.095 97.205 111.425 97.655 ;
        RECT 111.595 97.035 111.765 97.465 ;
        RECT 107.880 95.825 108.050 96.080 ;
        RECT 108.285 96.005 108.615 96.375 ;
        RECT 107.425 95.275 107.685 95.780 ;
        RECT 107.880 95.655 108.545 95.825 ;
        RECT 107.865 95.105 108.195 95.485 ;
        RECT 108.375 95.275 108.545 95.655 ;
        RECT 109.285 95.795 109.460 96.465 ;
        RECT 110.060 96.345 110.920 96.495 ;
        RECT 109.635 96.325 110.920 96.345 ;
        RECT 111.090 96.805 111.765 97.035 ;
        RECT 109.635 95.965 110.620 96.325 ;
        RECT 111.090 96.155 111.325 96.805 ;
        RECT 109.285 95.275 109.525 95.795 ;
        RECT 110.450 95.630 110.620 95.965 ;
        RECT 110.790 95.825 111.325 96.155 ;
        RECT 111.105 95.675 111.325 95.825 ;
        RECT 111.495 95.785 111.795 96.635 ;
        RECT 112.945 96.490 113.235 97.655 ;
        RECT 113.405 96.515 113.665 97.655 ;
        RECT 113.835 96.505 114.165 97.485 ;
        RECT 114.335 96.515 114.615 97.655 ;
        RECT 115.890 96.685 116.280 96.860 ;
        RECT 116.765 96.855 117.095 97.655 ;
        RECT 117.265 96.865 117.800 97.485 ;
        RECT 115.890 96.515 117.315 96.685 ;
        RECT 113.425 96.095 113.760 96.345 ;
        RECT 113.930 95.905 114.100 96.505 ;
        RECT 114.270 96.075 114.605 96.345 ;
        RECT 109.695 95.105 110.090 95.600 ;
        RECT 110.450 95.435 110.825 95.630 ;
        RECT 110.655 95.290 110.825 95.435 ;
        RECT 111.105 95.300 111.345 95.675 ;
        RECT 111.515 95.105 111.850 95.610 ;
        RECT 112.945 95.105 113.235 95.830 ;
        RECT 113.405 95.275 114.100 95.905 ;
        RECT 114.305 95.105 114.615 95.905 ;
        RECT 115.765 95.785 116.120 96.345 ;
        RECT 116.290 95.615 116.460 96.515 ;
        RECT 116.630 95.785 116.895 96.345 ;
        RECT 117.145 96.015 117.315 96.515 ;
        RECT 117.485 95.845 117.800 96.865 ;
        RECT 118.015 96.685 118.345 97.470 ;
        RECT 118.015 96.515 118.695 96.685 ;
        RECT 118.875 96.515 119.205 97.655 ;
        RECT 120.490 96.685 120.880 96.860 ;
        RECT 121.365 96.855 121.695 97.655 ;
        RECT 121.865 96.865 122.400 97.485 ;
        RECT 120.490 96.515 121.915 96.685 ;
        RECT 118.005 96.095 118.355 96.345 ;
        RECT 118.525 95.915 118.695 96.515 ;
        RECT 118.865 96.095 119.215 96.345 ;
        RECT 115.870 95.105 116.110 95.615 ;
        RECT 116.290 95.285 116.570 95.615 ;
        RECT 116.800 95.105 117.015 95.615 ;
        RECT 117.185 95.275 117.800 95.845 ;
        RECT 118.025 95.105 118.265 95.915 ;
        RECT 118.435 95.275 118.765 95.915 ;
        RECT 118.935 95.105 119.205 95.915 ;
        RECT 120.365 95.785 120.720 96.345 ;
        RECT 120.890 95.615 121.060 96.515 ;
        RECT 121.230 95.785 121.495 96.345 ;
        RECT 121.745 96.015 121.915 96.515 ;
        RECT 122.085 95.845 122.400 96.865 ;
        RECT 122.615 96.705 122.890 97.475 ;
        RECT 123.060 97.045 123.390 97.475 ;
        RECT 123.560 97.215 123.755 97.655 ;
        RECT 123.935 97.045 124.265 97.475 ;
        RECT 123.060 96.875 124.265 97.045 ;
        RECT 122.615 96.515 123.200 96.705 ;
        RECT 123.370 96.545 124.265 96.875 ;
        RECT 124.445 96.565 126.115 97.655 ;
        RECT 120.470 95.105 120.710 95.615 ;
        RECT 120.890 95.285 121.170 95.615 ;
        RECT 121.400 95.105 121.615 95.615 ;
        RECT 121.785 95.275 122.400 95.845 ;
        RECT 122.615 95.695 122.855 96.345 ;
        RECT 123.025 95.845 123.200 96.515 ;
        RECT 123.370 96.015 123.785 96.345 ;
        RECT 123.965 96.015 124.260 96.345 ;
        RECT 123.025 95.665 123.355 95.845 ;
        RECT 122.630 95.105 122.960 95.495 ;
        RECT 123.130 95.285 123.355 95.665 ;
        RECT 123.555 95.395 123.785 96.015 ;
        RECT 124.445 95.875 125.195 96.395 ;
        RECT 125.365 96.045 126.115 96.565 ;
        RECT 126.345 96.515 126.555 97.655 ;
        RECT 126.725 96.505 127.055 97.485 ;
        RECT 127.225 96.515 127.455 97.655 ;
        RECT 127.675 96.515 128.005 97.655 ;
        RECT 128.535 96.685 128.865 97.470 ;
        RECT 129.045 97.220 134.390 97.655 ;
        RECT 128.185 96.515 128.865 96.685 ;
        RECT 123.965 95.105 124.265 95.835 ;
        RECT 124.445 95.105 126.115 95.875 ;
        RECT 126.345 95.105 126.555 95.925 ;
        RECT 126.725 95.905 126.975 96.505 ;
        RECT 127.145 96.095 127.475 96.345 ;
        RECT 127.665 96.095 128.015 96.345 ;
        RECT 126.725 95.275 127.055 95.905 ;
        RECT 127.225 95.105 127.455 95.925 ;
        RECT 128.185 95.915 128.355 96.515 ;
        RECT 128.525 96.095 128.875 96.345 ;
        RECT 127.675 95.105 127.945 95.915 ;
        RECT 128.115 95.275 128.445 95.915 ;
        RECT 128.615 95.105 128.855 95.915 ;
        RECT 130.630 95.650 130.970 96.480 ;
        RECT 132.450 95.970 132.800 97.220 ;
        RECT 134.565 96.565 135.775 97.655 ;
        RECT 134.565 95.855 135.085 96.395 ;
        RECT 135.255 96.025 135.775 96.565 ;
        RECT 135.980 96.865 136.515 97.485 ;
        RECT 129.045 95.105 134.390 95.650 ;
        RECT 134.565 95.105 135.775 95.855 ;
        RECT 135.980 95.845 136.295 96.865 ;
        RECT 136.685 96.855 137.015 97.655 ;
        RECT 137.500 96.685 137.890 96.860 ;
        RECT 136.465 96.515 137.890 96.685 ;
        RECT 136.465 96.015 136.635 96.515 ;
        RECT 135.980 95.275 136.595 95.845 ;
        RECT 136.885 95.785 137.150 96.345 ;
        RECT 137.320 95.615 137.490 96.515 ;
        RECT 138.705 96.490 138.995 97.655 ;
        RECT 139.225 96.595 139.555 97.440 ;
        RECT 139.725 96.645 139.895 97.655 ;
        RECT 140.065 96.925 140.405 97.485 ;
        RECT 140.635 97.155 140.950 97.655 ;
        RECT 141.130 97.185 142.015 97.355 ;
        RECT 139.165 96.515 139.555 96.595 ;
        RECT 140.065 96.550 140.960 96.925 ;
        RECT 139.165 96.465 139.380 96.515 ;
        RECT 137.660 95.785 138.015 96.345 ;
        RECT 139.165 95.885 139.335 96.465 ;
        RECT 140.065 96.345 140.255 96.550 ;
        RECT 141.130 96.345 141.300 97.185 ;
        RECT 142.240 97.155 142.490 97.485 ;
        RECT 139.505 96.015 140.255 96.345 ;
        RECT 140.425 96.015 141.300 96.345 ;
        RECT 139.165 95.845 139.390 95.885 ;
        RECT 140.055 95.845 140.255 96.015 ;
        RECT 136.765 95.105 136.980 95.615 ;
        RECT 137.210 95.285 137.490 95.615 ;
        RECT 137.670 95.105 137.910 95.615 ;
        RECT 138.705 95.105 138.995 95.830 ;
        RECT 139.165 95.760 139.545 95.845 ;
        RECT 139.215 95.325 139.545 95.760 ;
        RECT 139.715 95.105 139.885 95.715 ;
        RECT 140.055 95.320 140.385 95.845 ;
        RECT 140.645 95.105 140.855 95.635 ;
        RECT 141.130 95.555 141.300 96.015 ;
        RECT 141.470 96.055 141.790 97.015 ;
        RECT 141.960 96.265 142.150 96.985 ;
        RECT 142.320 96.085 142.490 97.155 ;
        RECT 142.660 96.855 142.830 97.655 ;
        RECT 143.000 97.210 144.105 97.380 ;
        RECT 143.000 96.595 143.170 97.210 ;
        RECT 144.315 97.060 144.565 97.485 ;
        RECT 144.735 97.195 145.000 97.655 ;
        RECT 143.340 96.675 143.870 97.040 ;
        RECT 144.315 96.930 144.620 97.060 ;
        RECT 142.660 96.505 143.170 96.595 ;
        RECT 142.660 96.335 143.530 96.505 ;
        RECT 142.660 96.265 142.830 96.335 ;
        RECT 142.950 96.085 143.150 96.115 ;
        RECT 141.470 95.725 141.935 96.055 ;
        RECT 142.320 95.785 143.150 96.085 ;
        RECT 142.320 95.555 142.490 95.785 ;
        RECT 141.130 95.385 141.915 95.555 ;
        RECT 142.085 95.385 142.490 95.555 ;
        RECT 142.670 95.105 143.040 95.605 ;
        RECT 143.360 95.555 143.530 96.335 ;
        RECT 143.700 95.975 143.870 96.675 ;
        RECT 144.040 96.145 144.280 96.740 ;
        RECT 143.700 95.755 144.225 95.975 ;
        RECT 144.450 95.825 144.620 96.930 ;
        RECT 144.395 95.695 144.620 95.825 ;
        RECT 144.790 95.735 145.070 96.685 ;
        RECT 144.395 95.555 144.565 95.695 ;
        RECT 143.360 95.385 144.035 95.555 ;
        RECT 144.230 95.385 144.565 95.555 ;
        RECT 144.735 95.105 144.985 95.565 ;
        RECT 145.240 95.365 145.425 97.485 ;
        RECT 145.595 97.155 145.925 97.655 ;
        RECT 146.095 96.985 146.265 97.485 ;
        RECT 145.600 96.815 146.265 96.985 ;
        RECT 145.600 95.825 145.830 96.815 ;
        RECT 146.000 95.995 146.350 96.645 ;
        RECT 146.525 96.565 147.735 97.655 ;
        RECT 147.995 96.985 148.165 97.485 ;
        RECT 148.335 97.155 148.665 97.655 ;
        RECT 147.995 96.815 148.660 96.985 ;
        RECT 146.525 95.855 147.045 96.395 ;
        RECT 147.215 96.025 147.735 96.565 ;
        RECT 147.910 95.995 148.260 96.645 ;
        RECT 145.600 95.655 146.265 95.825 ;
        RECT 145.595 95.105 145.925 95.485 ;
        RECT 146.095 95.365 146.265 95.655 ;
        RECT 146.525 95.105 147.735 95.855 ;
        RECT 148.430 95.825 148.660 96.815 ;
        RECT 147.995 95.655 148.660 95.825 ;
        RECT 147.995 95.365 148.165 95.655 ;
        RECT 148.335 95.105 148.665 95.485 ;
        RECT 148.835 95.365 149.020 97.485 ;
        RECT 149.260 97.195 149.525 97.655 ;
        RECT 149.695 97.060 149.945 97.485 ;
        RECT 150.155 97.210 151.260 97.380 ;
        RECT 149.640 96.930 149.945 97.060 ;
        RECT 149.190 95.735 149.470 96.685 ;
        RECT 149.640 95.825 149.810 96.930 ;
        RECT 149.980 96.145 150.220 96.740 ;
        RECT 150.390 96.675 150.920 97.040 ;
        RECT 150.390 95.975 150.560 96.675 ;
        RECT 151.090 96.595 151.260 97.210 ;
        RECT 151.430 96.855 151.600 97.655 ;
        RECT 151.770 97.155 152.020 97.485 ;
        RECT 152.245 97.185 153.130 97.355 ;
        RECT 151.090 96.505 151.600 96.595 ;
        RECT 149.640 95.695 149.865 95.825 ;
        RECT 150.035 95.755 150.560 95.975 ;
        RECT 150.730 96.335 151.600 96.505 ;
        RECT 149.275 95.105 149.525 95.565 ;
        RECT 149.695 95.555 149.865 95.695 ;
        RECT 150.730 95.555 150.900 96.335 ;
        RECT 151.430 96.265 151.600 96.335 ;
        RECT 151.110 96.085 151.310 96.115 ;
        RECT 151.770 96.085 151.940 97.155 ;
        RECT 152.110 96.265 152.300 96.985 ;
        RECT 151.110 95.785 151.940 96.085 ;
        RECT 152.470 96.055 152.790 97.015 ;
        RECT 149.695 95.385 150.030 95.555 ;
        RECT 150.225 95.385 150.900 95.555 ;
        RECT 151.220 95.105 151.590 95.605 ;
        RECT 151.770 95.555 151.940 95.785 ;
        RECT 152.325 95.725 152.790 96.055 ;
        RECT 152.960 96.345 153.130 97.185 ;
        RECT 153.310 97.155 153.625 97.655 ;
        RECT 153.855 96.925 154.195 97.485 ;
        RECT 153.300 96.550 154.195 96.925 ;
        RECT 154.365 96.645 154.535 97.655 ;
        RECT 154.005 96.345 154.195 96.550 ;
        RECT 154.705 96.595 155.035 97.440 ;
        RECT 154.705 96.515 155.095 96.595 ;
        RECT 154.880 96.465 155.095 96.515 ;
        RECT 152.960 96.015 153.835 96.345 ;
        RECT 154.005 96.015 154.755 96.345 ;
        RECT 152.960 95.555 153.130 96.015 ;
        RECT 154.005 95.845 154.205 96.015 ;
        RECT 154.925 95.885 155.095 96.465 ;
        RECT 155.725 96.565 156.935 97.655 ;
        RECT 155.725 96.025 156.245 96.565 ;
        RECT 154.870 95.845 155.095 95.885 ;
        RECT 156.415 95.855 156.935 96.395 ;
        RECT 151.770 95.385 152.175 95.555 ;
        RECT 152.345 95.385 153.130 95.555 ;
        RECT 153.405 95.105 153.615 95.635 ;
        RECT 153.875 95.320 154.205 95.845 ;
        RECT 154.715 95.760 155.095 95.845 ;
        RECT 154.375 95.105 154.545 95.715 ;
        RECT 154.715 95.325 155.045 95.760 ;
        RECT 155.725 95.105 156.935 95.855 ;
        RECT 22.700 94.935 157.020 95.105 ;
        RECT 22.785 94.185 23.995 94.935 ;
        RECT 24.165 94.390 29.510 94.935 ;
        RECT 22.785 93.645 23.305 94.185 ;
        RECT 23.475 93.475 23.995 94.015 ;
        RECT 25.750 93.560 26.090 94.390 ;
        RECT 29.685 94.165 32.275 94.935 ;
        RECT 22.785 92.385 23.995 93.475 ;
        RECT 27.570 92.820 27.920 94.070 ;
        RECT 29.685 93.645 30.895 94.165 ;
        RECT 32.465 94.125 32.705 94.935 ;
        RECT 32.875 94.125 33.205 94.765 ;
        RECT 33.375 94.125 33.645 94.935 ;
        RECT 33.825 94.165 35.495 94.935 ;
        RECT 36.370 94.455 36.670 94.935 ;
        RECT 36.840 94.285 37.100 94.740 ;
        RECT 37.270 94.455 37.530 94.935 ;
        RECT 37.700 94.285 37.960 94.740 ;
        RECT 38.130 94.455 38.390 94.935 ;
        RECT 38.560 94.285 38.820 94.740 ;
        RECT 38.990 94.455 39.250 94.935 ;
        RECT 39.420 94.285 39.680 94.740 ;
        RECT 39.850 94.410 40.110 94.935 ;
        RECT 31.065 93.475 32.275 93.995 ;
        RECT 32.445 93.695 32.795 93.945 ;
        RECT 32.965 93.525 33.135 94.125 ;
        RECT 33.305 93.695 33.655 93.945 ;
        RECT 33.825 93.645 34.575 94.165 ;
        RECT 36.370 94.115 39.680 94.285 ;
        RECT 24.165 92.385 29.510 92.820 ;
        RECT 29.685 92.385 32.275 93.475 ;
        RECT 32.455 93.355 33.135 93.525 ;
        RECT 32.455 92.570 32.785 93.355 ;
        RECT 33.315 92.385 33.645 93.525 ;
        RECT 34.745 93.475 35.495 93.995 ;
        RECT 33.825 92.385 35.495 93.475 ;
        RECT 36.370 93.525 37.340 94.115 ;
        RECT 40.280 93.945 40.530 94.755 ;
        RECT 40.710 94.475 40.955 94.935 ;
        RECT 37.510 93.695 40.530 93.945 ;
        RECT 40.700 93.695 41.015 94.305 ;
        RECT 41.185 94.260 41.445 94.765 ;
        RECT 41.625 94.555 41.955 94.935 ;
        RECT 42.135 94.385 42.305 94.765 ;
        RECT 42.565 94.390 47.910 94.935 ;
        RECT 36.370 93.285 39.680 93.525 ;
        RECT 36.375 92.385 36.670 93.115 ;
        RECT 36.840 92.560 37.100 93.285 ;
        RECT 37.270 92.385 37.530 93.115 ;
        RECT 37.700 92.560 37.960 93.285 ;
        RECT 38.130 92.385 38.390 93.115 ;
        RECT 38.560 92.560 38.820 93.285 ;
        RECT 38.990 92.385 39.250 93.115 ;
        RECT 39.420 92.560 39.680 93.285 ;
        RECT 39.850 92.385 40.110 93.495 ;
        RECT 40.280 92.560 40.530 93.695 ;
        RECT 40.710 92.385 41.005 93.495 ;
        RECT 41.185 93.460 41.355 94.260 ;
        RECT 41.640 94.215 42.305 94.385 ;
        RECT 41.640 93.960 41.810 94.215 ;
        RECT 41.525 93.630 41.810 93.960 ;
        RECT 42.045 93.665 42.375 94.035 ;
        RECT 41.640 93.485 41.810 93.630 ;
        RECT 44.150 93.560 44.490 94.390 ;
        RECT 48.545 94.210 48.835 94.935 ;
        RECT 49.005 94.260 49.265 94.765 ;
        RECT 49.445 94.555 49.775 94.935 ;
        RECT 49.955 94.385 50.125 94.765 ;
        RECT 41.185 92.555 41.455 93.460 ;
        RECT 41.640 93.315 42.305 93.485 ;
        RECT 41.625 92.385 41.955 93.145 ;
        RECT 42.135 92.555 42.305 93.315 ;
        RECT 45.970 92.820 46.320 94.070 ;
        RECT 42.565 92.385 47.910 92.820 ;
        RECT 48.545 92.385 48.835 93.550 ;
        RECT 49.005 93.460 49.175 94.260 ;
        RECT 49.460 94.215 50.125 94.385 ;
        RECT 49.460 93.960 49.630 94.215 ;
        RECT 51.305 94.115 51.565 94.935 ;
        RECT 51.735 94.115 52.065 94.535 ;
        RECT 52.245 94.450 53.035 94.715 ;
        RECT 49.345 93.630 49.630 93.960 ;
        RECT 49.865 93.665 50.195 94.035 ;
        RECT 51.815 94.025 52.065 94.115 ;
        RECT 49.460 93.485 49.630 93.630 ;
        RECT 49.005 92.555 49.275 93.460 ;
        RECT 49.460 93.315 50.125 93.485 ;
        RECT 49.445 92.385 49.775 93.145 ;
        RECT 49.955 92.555 50.125 93.315 ;
        RECT 51.305 93.065 51.645 93.945 ;
        RECT 51.815 93.775 52.610 94.025 ;
        RECT 51.305 92.385 51.565 92.895 ;
        RECT 51.815 92.555 51.985 93.775 ;
        RECT 52.780 93.595 53.035 94.450 ;
        RECT 53.205 94.295 53.405 94.715 ;
        RECT 53.595 94.475 53.925 94.935 ;
        RECT 53.205 93.775 53.615 94.295 ;
        RECT 54.095 94.285 54.355 94.765 ;
        RECT 53.785 93.595 54.015 94.025 ;
        RECT 52.225 93.425 54.015 93.595 ;
        RECT 52.225 93.060 52.475 93.425 ;
        RECT 52.645 93.065 52.975 93.255 ;
        RECT 53.195 93.130 53.910 93.425 ;
        RECT 54.185 93.255 54.355 94.285 ;
        RECT 54.615 94.385 54.785 94.675 ;
        RECT 54.955 94.555 55.285 94.935 ;
        RECT 54.615 94.215 55.280 94.385 ;
        RECT 54.530 93.395 54.880 94.045 ;
        RECT 52.645 92.890 52.840 93.065 ;
        RECT 52.225 92.385 52.840 92.890 ;
        RECT 53.010 92.555 53.485 92.895 ;
        RECT 53.655 92.385 53.870 92.930 ;
        RECT 54.080 92.555 54.355 93.255 ;
        RECT 55.050 93.225 55.280 94.215 ;
        RECT 54.615 93.055 55.280 93.225 ;
        RECT 54.615 92.555 54.785 93.055 ;
        RECT 54.955 92.385 55.285 92.885 ;
        RECT 55.455 92.555 55.640 94.675 ;
        RECT 55.895 94.475 56.145 94.935 ;
        RECT 56.315 94.485 56.650 94.655 ;
        RECT 56.845 94.485 57.520 94.655 ;
        RECT 56.315 94.345 56.485 94.485 ;
        RECT 55.810 93.355 56.090 94.305 ;
        RECT 56.260 94.215 56.485 94.345 ;
        RECT 56.260 93.110 56.430 94.215 ;
        RECT 56.655 94.065 57.180 94.285 ;
        RECT 56.600 93.300 56.840 93.895 ;
        RECT 57.010 93.365 57.180 94.065 ;
        RECT 57.350 93.705 57.520 94.485 ;
        RECT 57.840 94.435 58.210 94.935 ;
        RECT 58.390 94.485 58.795 94.655 ;
        RECT 58.965 94.485 59.750 94.655 ;
        RECT 58.390 94.255 58.560 94.485 ;
        RECT 57.730 93.955 58.560 94.255 ;
        RECT 58.945 93.985 59.410 94.315 ;
        RECT 57.730 93.925 57.930 93.955 ;
        RECT 58.050 93.705 58.220 93.775 ;
        RECT 57.350 93.535 58.220 93.705 ;
        RECT 57.710 93.445 58.220 93.535 ;
        RECT 56.260 92.980 56.565 93.110 ;
        RECT 57.010 93.000 57.540 93.365 ;
        RECT 55.880 92.385 56.145 92.845 ;
        RECT 56.315 92.555 56.565 92.980 ;
        RECT 57.710 92.830 57.880 93.445 ;
        RECT 56.775 92.660 57.880 92.830 ;
        RECT 58.050 92.385 58.220 93.185 ;
        RECT 58.390 92.885 58.560 93.955 ;
        RECT 58.730 93.055 58.920 93.775 ;
        RECT 59.090 93.025 59.410 93.985 ;
        RECT 59.580 94.025 59.750 94.485 ;
        RECT 60.025 94.405 60.235 94.935 ;
        RECT 60.495 94.195 60.825 94.720 ;
        RECT 60.995 94.325 61.165 94.935 ;
        RECT 61.335 94.280 61.665 94.715 ;
        RECT 61.975 94.385 62.145 94.765 ;
        RECT 62.325 94.555 62.655 94.935 ;
        RECT 61.335 94.195 61.715 94.280 ;
        RECT 61.975 94.215 62.640 94.385 ;
        RECT 62.835 94.260 63.095 94.765 ;
        RECT 60.625 94.025 60.825 94.195 ;
        RECT 61.490 94.155 61.715 94.195 ;
        RECT 59.580 93.695 60.455 94.025 ;
        RECT 60.625 93.695 61.375 94.025 ;
        RECT 58.390 92.555 58.640 92.885 ;
        RECT 59.580 92.855 59.750 93.695 ;
        RECT 60.625 93.490 60.815 93.695 ;
        RECT 61.545 93.575 61.715 94.155 ;
        RECT 61.905 93.665 62.235 94.035 ;
        RECT 62.470 93.960 62.640 94.215 ;
        RECT 61.500 93.525 61.715 93.575 ;
        RECT 59.920 93.115 60.815 93.490 ;
        RECT 61.325 93.445 61.715 93.525 ;
        RECT 62.470 93.630 62.755 93.960 ;
        RECT 62.470 93.485 62.640 93.630 ;
        RECT 58.865 92.685 59.750 92.855 ;
        RECT 59.930 92.385 60.245 92.885 ;
        RECT 60.475 92.555 60.815 93.115 ;
        RECT 60.985 92.385 61.155 93.395 ;
        RECT 61.325 92.600 61.655 93.445 ;
        RECT 61.975 93.315 62.640 93.485 ;
        RECT 62.925 93.460 63.095 94.260 ;
        RECT 61.975 92.555 62.145 93.315 ;
        RECT 62.325 92.385 62.655 93.145 ;
        RECT 62.825 92.555 63.095 93.460 ;
        RECT 63.285 94.245 63.525 94.765 ;
        RECT 63.695 94.440 64.090 94.935 ;
        RECT 64.655 94.605 64.825 94.750 ;
        RECT 64.450 94.410 64.825 94.605 ;
        RECT 63.285 93.575 63.460 94.245 ;
        RECT 64.450 94.075 64.620 94.410 ;
        RECT 65.105 94.365 65.345 94.740 ;
        RECT 65.515 94.430 65.850 94.935 ;
        RECT 66.115 94.385 66.285 94.675 ;
        RECT 66.455 94.555 66.785 94.935 ;
        RECT 65.105 94.215 65.325 94.365 ;
        RECT 63.635 93.715 64.620 94.075 ;
        RECT 64.790 93.885 65.325 94.215 ;
        RECT 63.635 93.695 64.920 93.715 ;
        RECT 63.285 93.440 63.495 93.575 ;
        RECT 64.060 93.545 64.920 93.695 ;
        RECT 63.285 92.655 63.590 93.440 ;
        RECT 63.765 93.065 64.460 93.375 ;
        RECT 63.770 92.385 64.455 92.855 ;
        RECT 64.635 92.600 64.920 93.545 ;
        RECT 65.090 93.235 65.325 93.885 ;
        RECT 65.495 93.405 65.795 94.255 ;
        RECT 66.115 94.215 66.780 94.385 ;
        RECT 66.030 93.395 66.380 94.045 ;
        RECT 65.090 93.005 65.765 93.235 ;
        RECT 66.550 93.225 66.780 94.215 ;
        RECT 65.095 92.385 65.425 92.835 ;
        RECT 65.595 92.575 65.765 93.005 ;
        RECT 66.115 93.055 66.780 93.225 ;
        RECT 66.115 92.555 66.285 93.055 ;
        RECT 66.455 92.385 66.785 92.885 ;
        RECT 66.955 92.555 67.140 94.675 ;
        RECT 67.395 94.475 67.645 94.935 ;
        RECT 67.815 94.485 68.150 94.655 ;
        RECT 68.345 94.485 69.020 94.655 ;
        RECT 67.815 94.345 67.985 94.485 ;
        RECT 67.310 93.355 67.590 94.305 ;
        RECT 67.760 94.215 67.985 94.345 ;
        RECT 67.760 93.110 67.930 94.215 ;
        RECT 68.155 94.065 68.680 94.285 ;
        RECT 68.100 93.300 68.340 93.895 ;
        RECT 68.510 93.365 68.680 94.065 ;
        RECT 68.850 93.705 69.020 94.485 ;
        RECT 69.340 94.435 69.710 94.935 ;
        RECT 69.890 94.485 70.295 94.655 ;
        RECT 70.465 94.485 71.250 94.655 ;
        RECT 69.890 94.255 70.060 94.485 ;
        RECT 69.230 93.955 70.060 94.255 ;
        RECT 70.445 93.985 70.910 94.315 ;
        RECT 69.230 93.925 69.430 93.955 ;
        RECT 69.550 93.705 69.720 93.775 ;
        RECT 68.850 93.535 69.720 93.705 ;
        RECT 69.210 93.445 69.720 93.535 ;
        RECT 67.760 92.980 68.065 93.110 ;
        RECT 68.510 93.000 69.040 93.365 ;
        RECT 67.380 92.385 67.645 92.845 ;
        RECT 67.815 92.555 68.065 92.980 ;
        RECT 69.210 92.830 69.380 93.445 ;
        RECT 68.275 92.660 69.380 92.830 ;
        RECT 69.550 92.385 69.720 93.185 ;
        RECT 69.890 92.885 70.060 93.955 ;
        RECT 70.230 93.055 70.420 93.775 ;
        RECT 70.590 93.025 70.910 93.985 ;
        RECT 71.080 94.025 71.250 94.485 ;
        RECT 71.525 94.405 71.735 94.935 ;
        RECT 71.995 94.195 72.325 94.720 ;
        RECT 72.495 94.325 72.665 94.935 ;
        RECT 72.835 94.280 73.165 94.715 ;
        RECT 72.835 94.195 73.215 94.280 ;
        RECT 74.305 94.210 74.595 94.935 ;
        RECT 74.930 94.425 75.170 94.935 ;
        RECT 75.350 94.425 75.630 94.755 ;
        RECT 75.860 94.425 76.075 94.935 ;
        RECT 72.125 94.025 72.325 94.195 ;
        RECT 72.990 94.155 73.215 94.195 ;
        RECT 71.080 93.695 71.955 94.025 ;
        RECT 72.125 93.695 72.875 94.025 ;
        RECT 69.890 92.555 70.140 92.885 ;
        RECT 71.080 92.855 71.250 93.695 ;
        RECT 72.125 93.490 72.315 93.695 ;
        RECT 73.045 93.575 73.215 94.155 ;
        RECT 74.825 93.695 75.180 94.255 ;
        RECT 73.000 93.525 73.215 93.575 ;
        RECT 71.420 93.115 72.315 93.490 ;
        RECT 72.825 93.445 73.215 93.525 ;
        RECT 70.365 92.685 71.250 92.855 ;
        RECT 71.430 92.385 71.745 92.885 ;
        RECT 71.975 92.555 72.315 93.115 ;
        RECT 72.485 92.385 72.655 93.395 ;
        RECT 72.825 92.600 73.155 93.445 ;
        RECT 74.305 92.385 74.595 93.550 ;
        RECT 75.350 93.525 75.520 94.425 ;
        RECT 75.690 93.695 75.955 94.255 ;
        RECT 76.245 94.195 76.860 94.765 ;
        RECT 76.205 93.525 76.375 94.025 ;
        RECT 74.950 93.355 76.375 93.525 ;
        RECT 74.950 93.180 75.340 93.355 ;
        RECT 75.825 92.385 76.155 93.185 ;
        RECT 76.545 93.175 76.860 94.195 ;
        RECT 77.065 94.165 79.655 94.935 ;
        RECT 79.825 94.475 80.385 94.765 ;
        RECT 80.555 94.475 80.805 94.935 ;
        RECT 77.065 93.645 78.275 94.165 ;
        RECT 78.445 93.475 79.655 93.995 ;
        RECT 76.325 92.555 76.860 93.175 ;
        RECT 77.065 92.385 79.655 93.475 ;
        RECT 79.825 93.105 80.075 94.475 ;
        RECT 81.425 94.305 81.755 94.665 ;
        RECT 80.365 94.115 81.755 94.305 ;
        RECT 80.365 94.025 80.535 94.115 ;
        RECT 80.245 93.695 80.535 94.025 ;
        RECT 80.705 93.695 81.045 93.945 ;
        RECT 81.265 93.695 81.940 93.945 ;
        RECT 80.365 93.445 80.535 93.695 ;
        RECT 80.365 93.275 81.305 93.445 ;
        RECT 81.675 93.335 81.940 93.695 ;
        RECT 79.825 92.555 80.285 93.105 ;
        RECT 80.475 92.385 80.805 93.105 ;
        RECT 81.005 92.725 81.305 93.275 ;
        RECT 81.475 92.385 81.755 93.055 ;
        RECT 82.135 92.565 82.395 94.755 ;
        RECT 82.655 94.565 83.325 94.935 ;
        RECT 83.505 94.385 83.815 94.755 ;
        RECT 82.585 94.185 83.815 94.385 ;
        RECT 82.585 93.515 82.875 94.185 ;
        RECT 83.995 94.005 84.225 94.645 ;
        RECT 84.405 94.205 84.695 94.935 ;
        RECT 85.215 94.535 85.545 94.935 ;
        RECT 85.715 94.365 86.045 94.705 ;
        RECT 87.095 94.535 87.425 94.935 ;
        RECT 85.060 94.195 87.425 94.365 ;
        RECT 87.595 94.210 87.925 94.720 ;
        RECT 88.195 94.385 88.365 94.675 ;
        RECT 88.535 94.555 88.865 94.935 ;
        RECT 88.195 94.215 88.860 94.385 ;
        RECT 83.055 93.695 83.520 94.005 ;
        RECT 83.700 93.695 84.225 94.005 ;
        RECT 84.405 93.695 84.705 94.025 ;
        RECT 82.585 93.295 83.355 93.515 ;
        RECT 82.565 92.385 82.905 93.115 ;
        RECT 83.085 92.565 83.355 93.295 ;
        RECT 83.535 93.275 84.695 93.515 ;
        RECT 83.535 92.565 83.765 93.275 ;
        RECT 83.935 92.385 84.265 93.095 ;
        RECT 84.435 92.565 84.695 93.275 ;
        RECT 85.060 93.195 85.230 94.195 ;
        RECT 87.255 94.025 87.425 94.195 ;
        RECT 85.400 93.365 85.645 94.025 ;
        RECT 85.860 93.365 86.125 94.025 ;
        RECT 86.320 93.365 86.605 94.025 ;
        RECT 86.780 93.695 87.085 94.025 ;
        RECT 87.255 93.695 87.565 94.025 ;
        RECT 86.780 93.365 86.995 93.695 ;
        RECT 85.060 93.025 85.515 93.195 ;
        RECT 85.185 92.595 85.515 93.025 ;
        RECT 85.695 93.025 86.985 93.195 ;
        RECT 85.695 92.605 85.945 93.025 ;
        RECT 86.175 92.385 86.505 92.855 ;
        RECT 86.735 92.605 86.985 93.025 ;
        RECT 87.175 92.385 87.425 93.525 ;
        RECT 87.735 93.445 87.925 94.210 ;
        RECT 87.595 92.595 87.925 93.445 ;
        RECT 88.110 93.395 88.460 94.045 ;
        RECT 88.630 93.225 88.860 94.215 ;
        RECT 88.195 93.055 88.860 93.225 ;
        RECT 88.195 92.555 88.365 93.055 ;
        RECT 88.535 92.385 88.865 92.885 ;
        RECT 89.035 92.555 89.220 94.675 ;
        RECT 89.475 94.475 89.725 94.935 ;
        RECT 89.895 94.485 90.230 94.655 ;
        RECT 90.425 94.485 91.100 94.655 ;
        RECT 89.895 94.345 90.065 94.485 ;
        RECT 89.390 93.355 89.670 94.305 ;
        RECT 89.840 94.215 90.065 94.345 ;
        RECT 89.840 93.110 90.010 94.215 ;
        RECT 90.235 94.065 90.760 94.285 ;
        RECT 90.180 93.300 90.420 93.895 ;
        RECT 90.590 93.365 90.760 94.065 ;
        RECT 90.930 93.705 91.100 94.485 ;
        RECT 91.420 94.435 91.790 94.935 ;
        RECT 91.970 94.485 92.375 94.655 ;
        RECT 92.545 94.485 93.330 94.655 ;
        RECT 91.970 94.255 92.140 94.485 ;
        RECT 91.310 93.955 92.140 94.255 ;
        RECT 92.525 93.985 92.990 94.315 ;
        RECT 91.310 93.925 91.510 93.955 ;
        RECT 91.630 93.705 91.800 93.775 ;
        RECT 90.930 93.535 91.800 93.705 ;
        RECT 91.290 93.445 91.800 93.535 ;
        RECT 89.840 92.980 90.145 93.110 ;
        RECT 90.590 93.000 91.120 93.365 ;
        RECT 89.460 92.385 89.725 92.845 ;
        RECT 89.895 92.555 90.145 92.980 ;
        RECT 91.290 92.830 91.460 93.445 ;
        RECT 90.355 92.660 91.460 92.830 ;
        RECT 91.630 92.385 91.800 93.185 ;
        RECT 91.970 92.885 92.140 93.955 ;
        RECT 92.310 93.055 92.500 93.775 ;
        RECT 92.670 93.025 92.990 93.985 ;
        RECT 93.160 94.025 93.330 94.485 ;
        RECT 93.605 94.405 93.815 94.935 ;
        RECT 94.075 94.195 94.405 94.720 ;
        RECT 94.575 94.325 94.745 94.935 ;
        RECT 94.915 94.280 95.245 94.715 ;
        RECT 95.475 94.575 97.545 94.765 ;
        RECT 97.775 94.575 98.105 94.935 ;
        RECT 98.635 94.575 98.965 94.935 ;
        RECT 99.495 94.575 99.825 94.935 ;
        RECT 96.425 94.555 97.545 94.575 ;
        RECT 94.915 94.195 95.295 94.280 ;
        RECT 94.205 94.025 94.405 94.195 ;
        RECT 95.070 94.155 95.295 94.195 ;
        RECT 93.160 93.695 94.035 94.025 ;
        RECT 94.205 93.695 94.955 94.025 ;
        RECT 91.970 92.555 92.220 92.885 ;
        RECT 93.160 92.855 93.330 93.695 ;
        RECT 94.205 93.490 94.395 93.695 ;
        RECT 95.125 93.575 95.295 94.155 ;
        RECT 95.080 93.525 95.295 93.575 ;
        RECT 93.500 93.115 94.395 93.490 ;
        RECT 94.905 93.445 95.295 93.525 ;
        RECT 92.445 92.685 93.330 92.855 ;
        RECT 93.510 92.385 93.825 92.885 ;
        RECT 94.055 92.555 94.395 93.115 ;
        RECT 94.565 92.385 94.735 93.395 ;
        RECT 94.905 92.600 95.235 93.445 ;
        RECT 95.465 93.050 95.755 94.025 ;
        RECT 95.925 93.480 96.255 94.350 ;
        RECT 96.425 94.130 96.615 94.555 ;
        RECT 99.135 94.385 99.325 94.505 ;
        RECT 96.785 94.175 99.325 94.385 ;
        RECT 99.495 93.945 99.835 94.255 ;
        RECT 100.065 94.210 100.355 94.935 ;
        RECT 100.615 94.385 100.785 94.675 ;
        RECT 100.955 94.555 101.285 94.935 ;
        RECT 100.615 94.215 101.280 94.385 ;
        RECT 96.425 93.655 97.285 93.945 ;
        RECT 97.745 93.665 98.715 93.945 ;
        RECT 98.885 93.775 99.835 93.945 ;
        RECT 98.940 93.725 99.835 93.775 ;
        RECT 95.925 93.310 98.535 93.480 ;
        RECT 95.495 92.385 95.755 92.845 ;
        RECT 95.925 92.555 96.185 93.310 ;
        RECT 96.355 92.385 96.685 93.105 ;
        RECT 96.855 92.555 97.045 93.310 ;
        RECT 97.215 92.385 97.545 93.105 ;
        RECT 97.775 92.725 98.035 92.920 ;
        RECT 98.205 92.895 98.535 93.310 ;
        RECT 98.705 93.325 99.825 93.495 ;
        RECT 98.705 92.725 98.895 93.325 ;
        RECT 97.775 92.555 98.895 92.725 ;
        RECT 99.065 92.385 99.395 93.155 ;
        RECT 99.565 92.555 99.825 93.325 ;
        RECT 100.065 92.385 100.355 93.550 ;
        RECT 100.530 93.395 100.880 94.045 ;
        RECT 101.050 93.225 101.280 94.215 ;
        RECT 100.615 93.055 101.280 93.225 ;
        RECT 100.615 92.555 100.785 93.055 ;
        RECT 100.955 92.385 101.285 92.885 ;
        RECT 101.455 92.555 101.640 94.675 ;
        RECT 101.895 94.475 102.145 94.935 ;
        RECT 102.315 94.485 102.650 94.655 ;
        RECT 102.845 94.485 103.520 94.655 ;
        RECT 102.315 94.345 102.485 94.485 ;
        RECT 101.810 93.355 102.090 94.305 ;
        RECT 102.260 94.215 102.485 94.345 ;
        RECT 102.260 93.110 102.430 94.215 ;
        RECT 102.655 94.065 103.180 94.285 ;
        RECT 102.600 93.300 102.840 93.895 ;
        RECT 103.010 93.365 103.180 94.065 ;
        RECT 103.350 93.705 103.520 94.485 ;
        RECT 103.840 94.435 104.210 94.935 ;
        RECT 104.390 94.485 104.795 94.655 ;
        RECT 104.965 94.485 105.750 94.655 ;
        RECT 104.390 94.255 104.560 94.485 ;
        RECT 103.730 93.955 104.560 94.255 ;
        RECT 104.945 93.985 105.410 94.315 ;
        RECT 103.730 93.925 103.930 93.955 ;
        RECT 104.050 93.705 104.220 93.775 ;
        RECT 103.350 93.535 104.220 93.705 ;
        RECT 103.710 93.445 104.220 93.535 ;
        RECT 102.260 92.980 102.565 93.110 ;
        RECT 103.010 93.000 103.540 93.365 ;
        RECT 101.880 92.385 102.145 92.845 ;
        RECT 102.315 92.555 102.565 92.980 ;
        RECT 103.710 92.830 103.880 93.445 ;
        RECT 102.775 92.660 103.880 92.830 ;
        RECT 104.050 92.385 104.220 93.185 ;
        RECT 104.390 92.885 104.560 93.955 ;
        RECT 104.730 93.055 104.920 93.775 ;
        RECT 105.090 93.025 105.410 93.985 ;
        RECT 105.580 94.025 105.750 94.485 ;
        RECT 106.025 94.405 106.235 94.935 ;
        RECT 106.495 94.195 106.825 94.720 ;
        RECT 106.995 94.325 107.165 94.935 ;
        RECT 107.335 94.280 107.665 94.715 ;
        RECT 108.130 94.455 108.430 94.935 ;
        RECT 108.600 94.285 108.860 94.740 ;
        RECT 109.030 94.455 109.290 94.935 ;
        RECT 109.460 94.285 109.720 94.740 ;
        RECT 109.890 94.455 110.150 94.935 ;
        RECT 110.320 94.285 110.580 94.740 ;
        RECT 110.750 94.455 111.010 94.935 ;
        RECT 111.180 94.285 111.440 94.740 ;
        RECT 111.610 94.410 111.870 94.935 ;
        RECT 107.335 94.195 107.715 94.280 ;
        RECT 106.625 94.025 106.825 94.195 ;
        RECT 107.490 94.155 107.715 94.195 ;
        RECT 105.580 93.695 106.455 94.025 ;
        RECT 106.625 93.695 107.375 94.025 ;
        RECT 104.390 92.555 104.640 92.885 ;
        RECT 105.580 92.855 105.750 93.695 ;
        RECT 106.625 93.490 106.815 93.695 ;
        RECT 107.545 93.575 107.715 94.155 ;
        RECT 107.500 93.525 107.715 93.575 ;
        RECT 105.920 93.115 106.815 93.490 ;
        RECT 107.325 93.445 107.715 93.525 ;
        RECT 108.130 94.115 111.440 94.285 ;
        RECT 108.130 93.525 109.100 94.115 ;
        RECT 112.040 93.945 112.290 94.755 ;
        RECT 112.470 94.475 112.715 94.935 ;
        RECT 109.270 93.695 112.290 93.945 ;
        RECT 112.460 93.695 112.775 94.305 ;
        RECT 112.955 94.210 113.285 94.720 ;
        RECT 113.455 94.535 113.785 94.935 ;
        RECT 114.835 94.365 115.165 94.705 ;
        RECT 115.335 94.535 115.665 94.935 ;
        RECT 104.865 92.685 105.750 92.855 ;
        RECT 105.930 92.385 106.245 92.885 ;
        RECT 106.475 92.555 106.815 93.115 ;
        RECT 106.985 92.385 107.155 93.395 ;
        RECT 107.325 92.600 107.655 93.445 ;
        RECT 108.130 93.285 111.440 93.525 ;
        RECT 108.135 92.385 108.430 93.115 ;
        RECT 108.600 92.560 108.860 93.285 ;
        RECT 109.030 92.385 109.290 93.115 ;
        RECT 109.460 92.560 109.720 93.285 ;
        RECT 109.890 92.385 110.150 93.115 ;
        RECT 110.320 92.560 110.580 93.285 ;
        RECT 110.750 92.385 111.010 93.115 ;
        RECT 111.180 92.560 111.440 93.285 ;
        RECT 111.610 92.385 111.870 93.495 ;
        RECT 112.040 92.560 112.290 93.695 ;
        RECT 112.470 92.385 112.765 93.495 ;
        RECT 112.955 93.445 113.145 94.210 ;
        RECT 113.455 94.195 115.820 94.365 ;
        RECT 113.455 94.025 113.625 94.195 ;
        RECT 113.315 93.695 113.625 94.025 ;
        RECT 113.795 93.695 114.100 94.025 ;
        RECT 112.955 92.595 113.285 93.445 ;
        RECT 113.455 92.385 113.705 93.525 ;
        RECT 113.885 93.365 114.100 93.695 ;
        RECT 114.275 93.365 114.560 94.025 ;
        RECT 114.755 93.365 115.020 94.025 ;
        RECT 115.235 93.365 115.480 94.025 ;
        RECT 115.650 93.195 115.820 94.195 ;
        RECT 113.895 93.025 115.185 93.195 ;
        RECT 113.895 92.605 114.145 93.025 ;
        RECT 114.375 92.385 114.705 92.855 ;
        RECT 114.935 92.605 115.185 93.025 ;
        RECT 115.365 93.025 115.820 93.195 ;
        RECT 116.630 93.335 116.965 94.755 ;
        RECT 117.145 94.565 117.890 94.935 ;
        RECT 118.455 94.395 118.710 94.755 ;
        RECT 118.890 94.565 119.220 94.935 ;
        RECT 119.400 94.395 119.625 94.755 ;
        RECT 117.140 94.205 119.625 94.395 ;
        RECT 117.140 93.515 117.365 94.205 ;
        RECT 120.765 94.195 121.125 94.570 ;
        RECT 121.390 94.195 121.560 94.935 ;
        RECT 121.840 94.365 122.010 94.570 ;
        RECT 121.840 94.195 122.380 94.365 ;
        RECT 117.565 93.695 117.845 94.025 ;
        RECT 118.025 93.695 118.600 94.025 ;
        RECT 118.780 93.695 119.215 94.025 ;
        RECT 119.395 93.695 119.665 94.025 ;
        RECT 120.765 93.540 121.020 94.195 ;
        RECT 121.190 93.695 121.540 94.025 ;
        RECT 121.710 93.695 122.040 94.025 ;
        RECT 117.140 93.335 119.635 93.515 ;
        RECT 115.365 92.595 115.695 93.025 ;
        RECT 116.630 92.565 116.895 93.335 ;
        RECT 117.065 92.385 117.395 93.105 ;
        RECT 117.585 92.925 118.775 93.155 ;
        RECT 117.585 92.565 117.845 92.925 ;
        RECT 118.015 92.385 118.345 92.755 ;
        RECT 118.515 92.565 118.775 92.925 ;
        RECT 119.345 92.565 119.635 93.335 ;
        RECT 120.765 92.555 121.105 93.540 ;
        RECT 121.275 93.155 121.540 93.695 ;
        RECT 122.210 93.495 122.380 94.195 ;
        RECT 121.755 93.325 122.380 93.495 ;
        RECT 122.550 93.565 122.720 94.765 ;
        RECT 122.950 94.285 123.280 94.765 ;
        RECT 123.450 94.465 123.620 94.935 ;
        RECT 123.790 94.285 124.120 94.750 ;
        RECT 122.950 94.115 124.120 94.285 ;
        RECT 124.465 94.125 124.705 94.935 ;
        RECT 124.875 94.125 125.205 94.765 ;
        RECT 125.375 94.125 125.645 94.935 ;
        RECT 125.825 94.210 126.115 94.935 ;
        RECT 126.375 94.385 126.545 94.675 ;
        RECT 126.715 94.555 127.045 94.935 ;
        RECT 126.375 94.215 127.040 94.385 ;
        RECT 122.890 93.735 123.460 93.945 ;
        RECT 123.630 93.735 124.275 93.945 ;
        RECT 124.445 93.695 124.795 93.945 ;
        RECT 122.550 93.155 123.255 93.565 ;
        RECT 124.965 93.525 125.135 94.125 ;
        RECT 125.305 93.695 125.655 93.945 ;
        RECT 121.275 92.985 123.255 93.155 ;
        RECT 121.275 92.385 121.685 92.815 ;
        RECT 122.430 92.385 122.760 92.805 ;
        RECT 122.930 92.555 123.255 92.985 ;
        RECT 123.730 92.385 124.060 93.485 ;
        RECT 124.455 93.355 125.135 93.525 ;
        RECT 124.455 92.570 124.785 93.355 ;
        RECT 125.315 92.385 125.645 93.525 ;
        RECT 125.825 92.385 126.115 93.550 ;
        RECT 126.290 93.395 126.640 94.045 ;
        RECT 126.810 93.225 127.040 94.215 ;
        RECT 126.375 93.055 127.040 93.225 ;
        RECT 126.375 92.555 126.545 93.055 ;
        RECT 126.715 92.385 127.045 92.885 ;
        RECT 127.215 92.555 127.400 94.675 ;
        RECT 127.655 94.475 127.905 94.935 ;
        RECT 128.075 94.485 128.410 94.655 ;
        RECT 128.605 94.485 129.280 94.655 ;
        RECT 128.075 94.345 128.245 94.485 ;
        RECT 127.570 93.355 127.850 94.305 ;
        RECT 128.020 94.215 128.245 94.345 ;
        RECT 128.020 93.110 128.190 94.215 ;
        RECT 128.415 94.065 128.940 94.285 ;
        RECT 128.360 93.300 128.600 93.895 ;
        RECT 128.770 93.365 128.940 94.065 ;
        RECT 129.110 93.705 129.280 94.485 ;
        RECT 129.600 94.435 129.970 94.935 ;
        RECT 130.150 94.485 130.555 94.655 ;
        RECT 130.725 94.485 131.510 94.655 ;
        RECT 130.150 94.255 130.320 94.485 ;
        RECT 129.490 93.955 130.320 94.255 ;
        RECT 130.705 93.985 131.170 94.315 ;
        RECT 129.490 93.925 129.690 93.955 ;
        RECT 129.810 93.705 129.980 93.775 ;
        RECT 129.110 93.535 129.980 93.705 ;
        RECT 129.470 93.445 129.980 93.535 ;
        RECT 128.020 92.980 128.325 93.110 ;
        RECT 128.770 93.000 129.300 93.365 ;
        RECT 127.640 92.385 127.905 92.845 ;
        RECT 128.075 92.555 128.325 92.980 ;
        RECT 129.470 92.830 129.640 93.445 ;
        RECT 128.535 92.660 129.640 92.830 ;
        RECT 129.810 92.385 129.980 93.185 ;
        RECT 130.150 92.885 130.320 93.955 ;
        RECT 130.490 93.055 130.680 93.775 ;
        RECT 130.850 93.025 131.170 93.985 ;
        RECT 131.340 94.025 131.510 94.485 ;
        RECT 131.785 94.405 131.995 94.935 ;
        RECT 132.255 94.195 132.585 94.720 ;
        RECT 132.755 94.325 132.925 94.935 ;
        RECT 133.095 94.280 133.425 94.715 ;
        RECT 133.810 94.425 134.050 94.935 ;
        RECT 134.230 94.425 134.510 94.755 ;
        RECT 134.740 94.425 134.955 94.935 ;
        RECT 133.095 94.195 133.475 94.280 ;
        RECT 132.385 94.025 132.585 94.195 ;
        RECT 133.250 94.155 133.475 94.195 ;
        RECT 131.340 93.695 132.215 94.025 ;
        RECT 132.385 93.695 133.135 94.025 ;
        RECT 130.150 92.555 130.400 92.885 ;
        RECT 131.340 92.855 131.510 93.695 ;
        RECT 132.385 93.490 132.575 93.695 ;
        RECT 133.305 93.575 133.475 94.155 ;
        RECT 133.705 93.695 134.060 94.255 ;
        RECT 133.260 93.525 133.475 93.575 ;
        RECT 134.230 93.525 134.400 94.425 ;
        RECT 134.570 93.695 134.835 94.255 ;
        RECT 135.125 94.195 135.740 94.765 ;
        RECT 135.085 93.525 135.255 94.025 ;
        RECT 131.680 93.115 132.575 93.490 ;
        RECT 133.085 93.445 133.475 93.525 ;
        RECT 130.625 92.685 131.510 92.855 ;
        RECT 131.690 92.385 132.005 92.885 ;
        RECT 132.235 92.555 132.575 93.115 ;
        RECT 132.745 92.385 132.915 93.395 ;
        RECT 133.085 92.600 133.415 93.445 ;
        RECT 133.830 93.355 135.255 93.525 ;
        RECT 133.830 93.180 134.220 93.355 ;
        RECT 134.705 92.385 135.035 93.185 ;
        RECT 135.425 93.175 135.740 94.195 ;
        RECT 135.205 92.555 135.740 93.175 ;
        RECT 136.440 94.195 137.055 94.765 ;
        RECT 137.225 94.425 137.440 94.935 ;
        RECT 137.670 94.425 137.950 94.755 ;
        RECT 138.130 94.425 138.370 94.935 ;
        RECT 136.440 93.175 136.755 94.195 ;
        RECT 136.925 93.525 137.095 94.025 ;
        RECT 137.345 93.695 137.610 94.255 ;
        RECT 137.780 93.525 137.950 94.425 ;
        RECT 138.120 93.695 138.475 94.255 ;
        RECT 138.705 94.135 139.400 94.765 ;
        RECT 139.605 94.135 139.915 94.935 ;
        RECT 140.085 94.135 140.780 94.765 ;
        RECT 140.985 94.135 141.295 94.935 ;
        RECT 142.090 94.425 142.330 94.935 ;
        RECT 142.510 94.425 142.790 94.755 ;
        RECT 143.020 94.425 143.235 94.935 ;
        RECT 138.725 93.695 139.060 93.945 ;
        RECT 139.230 93.535 139.400 94.135 ;
        RECT 139.570 93.695 139.905 93.965 ;
        RECT 140.105 93.695 140.440 93.945 ;
        RECT 140.610 93.535 140.780 94.135 ;
        RECT 140.950 93.695 141.285 93.965 ;
        RECT 141.985 93.695 142.340 94.255 ;
        RECT 136.925 93.355 138.350 93.525 ;
        RECT 136.440 92.555 136.975 93.175 ;
        RECT 137.145 92.385 137.475 93.185 ;
        RECT 137.960 93.180 138.350 93.355 ;
        RECT 138.705 92.385 138.965 93.525 ;
        RECT 139.135 92.555 139.465 93.535 ;
        RECT 139.635 92.385 139.915 93.525 ;
        RECT 140.085 92.385 140.345 93.525 ;
        RECT 140.515 92.555 140.845 93.535 ;
        RECT 142.510 93.525 142.680 94.425 ;
        RECT 142.850 93.695 143.115 94.255 ;
        RECT 143.405 94.195 144.020 94.765 ;
        RECT 143.365 93.525 143.535 94.025 ;
        RECT 141.015 92.385 141.295 93.525 ;
        RECT 142.110 93.355 143.535 93.525 ;
        RECT 142.110 93.180 142.500 93.355 ;
        RECT 142.985 92.385 143.315 93.185 ;
        RECT 143.705 93.175 144.020 94.195 ;
        RECT 143.485 92.555 144.020 93.175 ;
        RECT 144.225 94.195 144.610 94.765 ;
        RECT 144.780 94.475 145.105 94.935 ;
        RECT 145.625 94.305 145.905 94.765 ;
        RECT 144.225 93.525 144.505 94.195 ;
        RECT 144.780 94.135 145.905 94.305 ;
        RECT 144.780 94.025 145.230 94.135 ;
        RECT 144.675 93.695 145.230 94.025 ;
        RECT 146.095 93.965 146.495 94.765 ;
        RECT 146.895 94.475 147.165 94.935 ;
        RECT 147.335 94.305 147.620 94.765 ;
        RECT 144.225 92.555 144.610 93.525 ;
        RECT 144.780 93.235 145.230 93.695 ;
        RECT 145.400 93.405 146.495 93.965 ;
        RECT 144.780 93.015 145.905 93.235 ;
        RECT 144.780 92.385 145.105 92.845 ;
        RECT 145.625 92.555 145.905 93.015 ;
        RECT 146.095 92.555 146.495 93.405 ;
        RECT 146.665 94.135 147.620 94.305 ;
        RECT 147.905 94.135 148.245 94.765 ;
        RECT 148.415 94.135 148.665 94.935 ;
        RECT 148.855 94.285 149.185 94.765 ;
        RECT 149.355 94.475 149.580 94.935 ;
        RECT 149.750 94.285 150.080 94.765 ;
        RECT 146.665 93.235 146.875 94.135 ;
        RECT 147.045 93.405 147.735 93.965 ;
        RECT 147.905 93.525 148.080 94.135 ;
        RECT 148.855 94.115 150.080 94.285 ;
        RECT 150.710 94.155 151.210 94.765 ;
        RECT 151.585 94.210 151.875 94.935 ;
        RECT 152.045 94.195 152.430 94.765 ;
        RECT 152.600 94.475 152.925 94.935 ;
        RECT 153.445 94.305 153.725 94.765 ;
        RECT 148.250 93.775 148.945 93.945 ;
        RECT 148.775 93.525 148.945 93.775 ;
        RECT 149.120 93.745 149.540 93.945 ;
        RECT 149.710 93.745 150.040 93.945 ;
        RECT 150.210 93.745 150.540 93.945 ;
        RECT 150.710 93.525 150.880 94.155 ;
        RECT 151.065 93.695 151.415 93.945 ;
        RECT 146.665 93.015 147.620 93.235 ;
        RECT 146.895 92.385 147.165 92.845 ;
        RECT 147.335 92.555 147.620 93.015 ;
        RECT 147.905 92.555 148.245 93.525 ;
        RECT 148.415 92.385 148.585 93.525 ;
        RECT 148.775 93.355 151.210 93.525 ;
        RECT 148.855 92.385 149.105 93.185 ;
        RECT 149.750 92.555 150.080 93.355 ;
        RECT 150.380 92.385 150.710 93.185 ;
        RECT 150.880 92.555 151.210 93.355 ;
        RECT 151.585 92.385 151.875 93.550 ;
        RECT 152.045 93.525 152.325 94.195 ;
        RECT 152.600 94.135 153.725 94.305 ;
        RECT 152.600 94.025 153.050 94.135 ;
        RECT 152.495 93.695 153.050 94.025 ;
        RECT 153.915 93.965 154.315 94.765 ;
        RECT 154.715 94.475 154.985 94.935 ;
        RECT 155.155 94.305 155.440 94.765 ;
        RECT 152.045 92.555 152.430 93.525 ;
        RECT 152.600 93.235 153.050 93.695 ;
        RECT 153.220 93.405 154.315 93.965 ;
        RECT 152.600 93.015 153.725 93.235 ;
        RECT 152.600 92.385 152.925 92.845 ;
        RECT 153.445 92.555 153.725 93.015 ;
        RECT 153.915 92.555 154.315 93.405 ;
        RECT 154.485 94.135 155.440 94.305 ;
        RECT 155.725 94.185 156.935 94.935 ;
        RECT 154.485 93.235 154.695 94.135 ;
        RECT 154.865 93.405 155.555 93.965 ;
        RECT 155.725 93.475 156.245 94.015 ;
        RECT 156.415 93.645 156.935 94.185 ;
        RECT 154.485 93.015 155.440 93.235 ;
        RECT 154.715 92.385 154.985 92.845 ;
        RECT 155.155 92.555 155.440 93.015 ;
        RECT 155.725 92.385 156.935 93.475 ;
        RECT 22.700 92.215 157.020 92.385 ;
        RECT 22.785 91.125 23.995 92.215 ;
        RECT 24.255 91.545 24.425 92.045 ;
        RECT 24.595 91.715 24.925 92.215 ;
        RECT 24.255 91.375 24.920 91.545 ;
        RECT 22.785 90.415 23.305 90.955 ;
        RECT 23.475 90.585 23.995 91.125 ;
        RECT 24.170 90.555 24.520 91.205 ;
        RECT 22.785 89.665 23.995 90.415 ;
        RECT 24.690 90.385 24.920 91.375 ;
        RECT 24.255 90.215 24.920 90.385 ;
        RECT 24.255 89.925 24.425 90.215 ;
        RECT 24.595 89.665 24.925 90.045 ;
        RECT 25.095 89.925 25.280 92.045 ;
        RECT 25.520 91.755 25.785 92.215 ;
        RECT 25.955 91.620 26.205 92.045 ;
        RECT 26.415 91.770 27.520 91.940 ;
        RECT 25.900 91.490 26.205 91.620 ;
        RECT 25.450 90.295 25.730 91.245 ;
        RECT 25.900 90.385 26.070 91.490 ;
        RECT 26.240 90.705 26.480 91.300 ;
        RECT 26.650 91.235 27.180 91.600 ;
        RECT 26.650 90.535 26.820 91.235 ;
        RECT 27.350 91.155 27.520 91.770 ;
        RECT 27.690 91.415 27.860 92.215 ;
        RECT 28.030 91.715 28.280 92.045 ;
        RECT 28.505 91.745 29.390 91.915 ;
        RECT 27.350 91.065 27.860 91.155 ;
        RECT 25.900 90.255 26.125 90.385 ;
        RECT 26.295 90.315 26.820 90.535 ;
        RECT 26.990 90.895 27.860 91.065 ;
        RECT 25.535 89.665 25.785 90.125 ;
        RECT 25.955 90.115 26.125 90.255 ;
        RECT 26.990 90.115 27.160 90.895 ;
        RECT 27.690 90.825 27.860 90.895 ;
        RECT 27.370 90.645 27.570 90.675 ;
        RECT 28.030 90.645 28.200 91.715 ;
        RECT 28.370 90.825 28.560 91.545 ;
        RECT 27.370 90.345 28.200 90.645 ;
        RECT 28.730 90.615 29.050 91.575 ;
        RECT 25.955 89.945 26.290 90.115 ;
        RECT 26.485 89.945 27.160 90.115 ;
        RECT 27.480 89.665 27.850 90.165 ;
        RECT 28.030 90.115 28.200 90.345 ;
        RECT 28.585 90.285 29.050 90.615 ;
        RECT 29.220 90.905 29.390 91.745 ;
        RECT 29.570 91.715 29.885 92.215 ;
        RECT 30.115 91.485 30.455 92.045 ;
        RECT 29.560 91.110 30.455 91.485 ;
        RECT 30.625 91.205 30.795 92.215 ;
        RECT 30.265 90.905 30.455 91.110 ;
        RECT 30.965 91.155 31.295 92.000 ;
        RECT 30.965 91.075 31.355 91.155 ;
        RECT 32.450 91.075 32.705 92.215 ;
        RECT 32.900 91.665 34.095 91.995 ;
        RECT 31.140 91.025 31.355 91.075 ;
        RECT 29.220 90.575 30.095 90.905 ;
        RECT 30.265 90.575 31.015 90.905 ;
        RECT 29.220 90.115 29.390 90.575 ;
        RECT 30.265 90.405 30.465 90.575 ;
        RECT 31.185 90.445 31.355 91.025 ;
        RECT 32.955 90.905 33.125 91.465 ;
        RECT 33.350 91.245 33.770 91.495 ;
        RECT 34.275 91.415 34.555 92.215 ;
        RECT 33.350 91.075 34.595 91.245 ;
        RECT 34.765 91.075 35.035 92.045 ;
        RECT 34.425 90.905 34.595 91.075 ;
        RECT 34.805 91.025 35.035 91.075 ;
        RECT 35.665 91.050 35.955 92.215 ;
        RECT 36.135 91.155 36.465 92.005 ;
        RECT 32.450 90.655 32.785 90.905 ;
        RECT 32.955 90.575 33.695 90.905 ;
        RECT 34.425 90.575 34.655 90.905 ;
        RECT 32.955 90.485 33.205 90.575 ;
        RECT 31.130 90.405 31.355 90.445 ;
        RECT 28.030 89.945 28.435 90.115 ;
        RECT 28.605 89.945 29.390 90.115 ;
        RECT 29.665 89.665 29.875 90.195 ;
        RECT 30.135 89.880 30.465 90.405 ;
        RECT 30.975 90.320 31.355 90.405 ;
        RECT 30.635 89.665 30.805 90.275 ;
        RECT 30.975 89.885 31.305 90.320 ;
        RECT 32.470 90.315 33.205 90.485 ;
        RECT 34.425 90.405 34.595 90.575 ;
        RECT 32.470 89.845 32.780 90.315 ;
        RECT 33.855 90.235 34.595 90.405 ;
        RECT 34.865 90.340 35.035 91.025 ;
        RECT 36.135 90.390 36.325 91.155 ;
        RECT 36.635 91.075 36.885 92.215 ;
        RECT 37.075 91.575 37.325 91.995 ;
        RECT 37.555 91.745 37.885 92.215 ;
        RECT 38.115 91.575 38.365 91.995 ;
        RECT 37.075 91.405 38.365 91.575 ;
        RECT 38.545 91.575 38.875 92.005 ;
        RECT 40.265 91.660 40.870 92.215 ;
        RECT 41.045 91.705 41.525 92.045 ;
        RECT 41.695 91.670 41.950 92.215 ;
        RECT 38.545 91.405 39.000 91.575 ;
        RECT 40.265 91.560 40.880 91.660 ;
        RECT 37.065 90.905 37.280 91.235 ;
        RECT 36.495 90.575 36.805 90.905 ;
        RECT 36.975 90.575 37.280 90.905 ;
        RECT 37.455 90.575 37.740 91.235 ;
        RECT 37.935 90.575 38.200 91.235 ;
        RECT 38.415 90.575 38.660 91.235 ;
        RECT 36.635 90.405 36.805 90.575 ;
        RECT 38.830 90.405 39.000 91.405 ;
        RECT 40.695 91.535 40.880 91.560 ;
        RECT 40.265 90.940 40.525 91.390 ;
        RECT 40.695 91.290 41.025 91.535 ;
        RECT 41.195 91.215 41.950 91.465 ;
        RECT 42.120 91.345 42.395 92.045 ;
        RECT 41.180 91.180 41.950 91.215 ;
        RECT 41.165 91.170 41.950 91.180 ;
        RECT 41.160 91.155 42.055 91.170 ;
        RECT 41.140 91.140 42.055 91.155 ;
        RECT 41.120 91.130 42.055 91.140 ;
        RECT 41.095 91.120 42.055 91.130 ;
        RECT 41.025 91.090 42.055 91.120 ;
        RECT 41.005 91.060 42.055 91.090 ;
        RECT 40.985 91.030 42.055 91.060 ;
        RECT 40.955 91.005 42.055 91.030 ;
        RECT 40.920 90.970 42.055 91.005 ;
        RECT 40.890 90.965 42.055 90.970 ;
        RECT 40.890 90.960 41.280 90.965 ;
        RECT 40.890 90.950 41.255 90.960 ;
        RECT 40.890 90.945 41.240 90.950 ;
        RECT 40.890 90.940 41.225 90.945 ;
        RECT 40.265 90.935 41.225 90.940 ;
        RECT 40.265 90.925 41.215 90.935 ;
        RECT 40.265 90.920 41.205 90.925 ;
        RECT 40.265 90.910 41.195 90.920 ;
        RECT 40.265 90.900 41.190 90.910 ;
        RECT 40.265 90.895 41.185 90.900 ;
        RECT 40.265 90.880 41.175 90.895 ;
        RECT 40.265 90.865 41.170 90.880 ;
        RECT 40.265 90.840 41.160 90.865 ;
        RECT 40.265 90.770 41.155 90.840 ;
        RECT 32.950 89.665 33.685 90.145 ;
        RECT 33.855 89.885 34.025 90.235 ;
        RECT 34.195 89.665 34.575 90.065 ;
        RECT 34.765 89.995 35.035 90.340 ;
        RECT 35.665 89.665 35.955 90.390 ;
        RECT 36.135 89.880 36.465 90.390 ;
        RECT 36.635 90.235 39.000 90.405 ;
        RECT 36.635 89.665 36.965 90.065 ;
        RECT 38.015 89.895 38.345 90.235 ;
        RECT 40.265 90.215 40.815 90.600 ;
        RECT 38.515 89.665 38.845 90.065 ;
        RECT 40.985 90.045 41.155 90.770 ;
        RECT 40.265 89.875 41.155 90.045 ;
        RECT 41.325 90.370 41.655 90.795 ;
        RECT 41.825 90.570 42.055 90.965 ;
        RECT 41.325 89.885 41.545 90.370 ;
        RECT 42.225 90.315 42.395 91.345 ;
        RECT 41.715 89.665 41.965 90.205 ;
        RECT 42.135 89.835 42.395 90.315 ;
        RECT 42.570 91.265 42.835 92.035 ;
        RECT 43.005 91.495 43.335 92.215 ;
        RECT 43.525 91.675 43.785 92.035 ;
        RECT 43.955 91.845 44.285 92.215 ;
        RECT 44.455 91.675 44.715 92.035 ;
        RECT 43.525 91.445 44.715 91.675 ;
        RECT 45.285 91.265 45.575 92.035 ;
        RECT 42.570 89.845 42.905 91.265 ;
        RECT 43.080 91.085 45.575 91.265 ;
        RECT 43.080 90.395 43.305 91.085 ;
        RECT 46.305 91.075 46.515 92.215 ;
        RECT 46.685 91.065 47.015 92.045 ;
        RECT 47.185 91.075 47.415 92.215 ;
        RECT 47.625 91.705 47.885 92.215 ;
        RECT 43.505 90.575 43.785 90.905 ;
        RECT 43.965 90.575 44.540 90.905 ;
        RECT 44.720 90.575 45.155 90.905 ;
        RECT 45.335 90.575 45.605 90.905 ;
        RECT 43.080 90.205 45.565 90.395 ;
        RECT 43.085 89.665 43.830 90.035 ;
        RECT 44.395 89.845 44.650 90.205 ;
        RECT 44.830 89.665 45.160 90.035 ;
        RECT 45.340 89.845 45.565 90.205 ;
        RECT 46.305 89.665 46.515 90.485 ;
        RECT 46.685 90.465 46.935 91.065 ;
        RECT 47.105 90.655 47.435 90.905 ;
        RECT 47.625 90.655 47.965 91.535 ;
        RECT 48.135 90.825 48.305 92.045 ;
        RECT 48.545 91.710 49.160 92.215 ;
        RECT 48.545 91.175 48.795 91.540 ;
        RECT 48.965 91.535 49.160 91.710 ;
        RECT 49.330 91.705 49.805 92.045 ;
        RECT 49.975 91.670 50.190 92.215 ;
        RECT 48.965 91.345 49.295 91.535 ;
        RECT 49.515 91.175 50.230 91.470 ;
        RECT 50.400 91.345 50.675 92.045 ;
        RECT 48.545 91.005 50.335 91.175 ;
        RECT 48.135 90.575 48.930 90.825 ;
        RECT 48.135 90.485 48.385 90.575 ;
        RECT 46.685 89.835 47.015 90.465 ;
        RECT 47.185 89.665 47.415 90.485 ;
        RECT 47.625 89.665 47.885 90.485 ;
        RECT 48.055 90.065 48.385 90.485 ;
        RECT 49.100 90.150 49.355 91.005 ;
        RECT 48.565 89.885 49.355 90.150 ;
        RECT 49.525 90.305 49.935 90.825 ;
        RECT 50.105 90.575 50.335 91.005 ;
        RECT 50.505 90.315 50.675 91.345 ;
        RECT 49.525 89.885 49.725 90.305 ;
        RECT 49.915 89.665 50.245 90.125 ;
        RECT 50.415 89.835 50.675 90.315 ;
        RECT 50.845 91.075 51.185 92.045 ;
        RECT 51.355 91.075 51.525 92.215 ;
        RECT 51.795 91.415 52.045 92.215 ;
        RECT 52.690 91.245 53.020 92.045 ;
        RECT 53.320 91.415 53.650 92.215 ;
        RECT 53.820 91.245 54.150 92.045 ;
        RECT 51.715 91.075 54.150 91.245 ;
        RECT 55.045 91.075 55.255 92.215 ;
        RECT 50.845 91.025 51.075 91.075 ;
        RECT 50.845 90.465 51.020 91.025 ;
        RECT 51.715 90.825 51.885 91.075 ;
        RECT 51.190 90.655 51.885 90.825 ;
        RECT 52.060 90.655 52.480 90.855 ;
        RECT 52.650 90.655 52.980 90.855 ;
        RECT 53.150 90.655 53.480 90.855 ;
        RECT 50.845 89.835 51.185 90.465 ;
        RECT 51.355 89.665 51.605 90.465 ;
        RECT 51.795 90.315 53.020 90.485 ;
        RECT 51.795 89.835 52.125 90.315 ;
        RECT 52.295 89.665 52.520 90.125 ;
        RECT 52.690 89.835 53.020 90.315 ;
        RECT 53.650 90.445 53.820 91.075 ;
        RECT 55.425 91.065 55.755 92.045 ;
        RECT 55.925 91.075 56.155 92.215 ;
        RECT 54.005 90.655 54.355 90.905 ;
        RECT 53.650 89.835 54.150 90.445 ;
        RECT 55.045 89.665 55.255 90.485 ;
        RECT 55.425 90.465 55.675 91.065 ;
        RECT 55.845 90.655 56.175 90.905 ;
        RECT 55.425 89.835 55.755 90.465 ;
        RECT 55.925 89.665 56.155 90.485 ;
        RECT 56.380 89.845 56.660 92.035 ;
        RECT 56.850 91.075 57.135 92.215 ;
        RECT 57.400 91.565 57.570 92.035 ;
        RECT 57.745 91.735 58.075 92.215 ;
        RECT 58.245 91.565 58.425 92.035 ;
        RECT 57.400 91.365 58.425 91.565 ;
        RECT 56.860 90.395 57.120 90.905 ;
        RECT 57.330 90.575 57.590 91.195 ;
        RECT 57.785 90.575 58.210 91.195 ;
        RECT 58.595 90.925 58.925 92.035 ;
        RECT 59.095 91.805 59.445 92.215 ;
        RECT 59.615 91.625 59.855 92.015 ;
        RECT 58.380 90.625 58.925 90.925 ;
        RECT 59.105 91.425 59.855 91.625 ;
        RECT 59.105 90.745 59.445 91.425 ;
        RECT 58.380 90.395 58.600 90.625 ;
        RECT 56.860 90.205 58.600 90.395 ;
        RECT 56.860 89.665 57.590 90.035 ;
        RECT 58.170 89.845 58.600 90.205 ;
        RECT 58.770 89.665 59.015 90.445 ;
        RECT 59.215 89.845 59.445 90.745 ;
        RECT 59.625 89.905 59.855 91.245 ;
        RECT 60.045 91.075 60.305 92.215 ;
        RECT 60.475 91.065 60.805 92.045 ;
        RECT 60.975 91.075 61.255 92.215 ;
        RECT 60.565 91.025 60.740 91.065 ;
        RECT 61.425 91.050 61.715 92.215 ;
        RECT 62.070 91.245 62.460 91.420 ;
        RECT 62.945 91.415 63.275 92.215 ;
        RECT 63.445 91.425 63.980 92.045 ;
        RECT 62.070 91.075 63.495 91.245 ;
        RECT 60.065 90.655 60.400 90.905 ;
        RECT 60.570 90.465 60.740 91.025 ;
        RECT 60.910 90.635 61.245 90.905 ;
        RECT 60.045 89.835 60.740 90.465 ;
        RECT 60.945 89.665 61.255 90.465 ;
        RECT 61.425 89.665 61.715 90.390 ;
        RECT 61.945 90.345 62.300 90.905 ;
        RECT 62.470 90.175 62.640 91.075 ;
        RECT 62.810 90.345 63.075 90.905 ;
        RECT 63.325 90.575 63.495 91.075 ;
        RECT 63.665 90.405 63.980 91.425 ;
        RECT 64.185 91.125 65.855 92.215 ;
        RECT 62.050 89.665 62.290 90.175 ;
        RECT 62.470 89.845 62.750 90.175 ;
        RECT 62.980 89.665 63.195 90.175 ;
        RECT 63.365 89.835 63.980 90.405 ;
        RECT 64.185 90.435 64.935 90.955 ;
        RECT 65.105 90.605 65.855 91.125 ;
        RECT 66.495 91.155 66.825 92.005 ;
        RECT 64.185 89.665 65.855 90.435 ;
        RECT 66.495 90.390 66.685 91.155 ;
        RECT 66.995 91.075 67.245 92.215 ;
        RECT 67.435 91.575 67.685 91.995 ;
        RECT 67.915 91.745 68.245 92.215 ;
        RECT 68.475 91.575 68.725 91.995 ;
        RECT 67.435 91.405 68.725 91.575 ;
        RECT 68.905 91.575 69.235 92.005 ;
        RECT 68.905 91.405 69.360 91.575 ;
        RECT 67.425 90.905 67.640 91.235 ;
        RECT 66.855 90.575 67.165 90.905 ;
        RECT 67.335 90.575 67.640 90.905 ;
        RECT 67.815 90.575 68.100 91.235 ;
        RECT 68.295 90.575 68.560 91.235 ;
        RECT 68.775 90.575 69.020 91.235 ;
        RECT 66.995 90.405 67.165 90.575 ;
        RECT 69.190 90.405 69.360 91.405 ;
        RECT 66.495 89.880 66.825 90.390 ;
        RECT 66.995 90.235 69.360 90.405 ;
        RECT 66.995 89.665 67.325 90.065 ;
        RECT 68.375 89.895 68.705 90.235 ;
        RECT 68.875 89.665 69.205 90.065 ;
        RECT 69.715 89.845 69.975 92.035 ;
        RECT 70.145 91.485 70.485 92.215 ;
        RECT 70.665 91.305 70.935 92.035 ;
        RECT 70.165 91.085 70.935 91.305 ;
        RECT 71.115 91.325 71.345 92.035 ;
        RECT 71.515 91.505 71.845 92.215 ;
        RECT 72.015 91.325 72.275 92.035 ;
        RECT 71.115 91.085 72.275 91.325 ;
        RECT 70.165 90.415 70.455 91.085 ;
        RECT 72.465 91.075 72.725 92.215 ;
        RECT 72.895 91.065 73.225 92.045 ;
        RECT 73.395 91.075 73.675 92.215 ;
        RECT 73.845 91.125 77.355 92.215 ;
        RECT 70.635 90.595 71.100 90.905 ;
        RECT 71.280 90.595 71.805 90.905 ;
        RECT 70.165 90.215 71.395 90.415 ;
        RECT 70.235 89.665 70.905 90.035 ;
        RECT 71.085 89.845 71.395 90.215 ;
        RECT 71.575 89.955 71.805 90.595 ;
        RECT 71.985 90.575 72.285 90.905 ;
        RECT 72.485 90.655 72.820 90.905 ;
        RECT 72.990 90.515 73.160 91.065 ;
        RECT 73.330 90.635 73.665 90.905 ;
        RECT 72.985 90.465 73.160 90.515 ;
        RECT 71.985 89.665 72.275 90.395 ;
        RECT 72.465 89.835 73.160 90.465 ;
        RECT 73.365 89.665 73.675 90.465 ;
        RECT 73.845 90.435 75.495 90.955 ;
        RECT 75.665 90.605 77.355 91.125 ;
        RECT 77.985 91.060 78.325 92.045 ;
        RECT 78.495 91.785 78.905 92.215 ;
        RECT 79.650 91.795 79.980 92.215 ;
        RECT 80.150 91.615 80.475 92.045 ;
        RECT 78.495 91.445 80.475 91.615 ;
        RECT 73.845 89.665 77.355 90.435 ;
        RECT 77.985 90.405 78.240 91.060 ;
        RECT 78.495 90.905 78.760 91.445 ;
        RECT 78.975 91.105 79.600 91.275 ;
        RECT 78.410 90.575 78.760 90.905 ;
        RECT 78.930 90.575 79.260 90.905 ;
        RECT 79.430 90.405 79.600 91.105 ;
        RECT 77.985 90.030 78.345 90.405 ;
        RECT 78.045 90.005 78.215 90.030 ;
        RECT 78.610 89.665 78.780 90.405 ;
        RECT 79.060 90.235 79.600 90.405 ;
        RECT 79.770 91.035 80.475 91.445 ;
        RECT 80.950 91.115 81.280 92.215 ;
        RECT 81.675 91.155 82.005 92.005 ;
        RECT 79.060 90.030 79.230 90.235 ;
        RECT 79.770 89.835 79.940 91.035 ;
        RECT 81.675 91.025 81.895 91.155 ;
        RECT 82.175 91.075 82.425 92.215 ;
        RECT 82.615 91.575 82.865 91.995 ;
        RECT 83.095 91.745 83.425 92.215 ;
        RECT 83.655 91.575 83.905 91.995 ;
        RECT 82.615 91.405 83.905 91.575 ;
        RECT 84.085 91.575 84.415 92.005 ;
        RECT 84.085 91.405 84.540 91.575 ;
        RECT 80.110 90.655 80.680 90.865 ;
        RECT 80.850 90.655 81.495 90.865 ;
        RECT 80.170 90.315 81.340 90.485 ;
        RECT 80.170 89.835 80.500 90.315 ;
        RECT 80.670 89.665 80.840 90.135 ;
        RECT 81.010 89.850 81.340 90.315 ;
        RECT 81.675 90.390 81.865 91.025 ;
        RECT 82.605 90.905 82.820 91.235 ;
        RECT 82.035 90.575 82.345 90.905 ;
        RECT 82.515 90.575 82.820 90.905 ;
        RECT 82.995 90.575 83.280 91.235 ;
        RECT 83.475 90.575 83.740 91.235 ;
        RECT 83.955 90.575 84.200 91.235 ;
        RECT 82.175 90.405 82.345 90.575 ;
        RECT 84.370 90.405 84.540 91.405 ;
        RECT 84.885 91.125 86.555 92.215 ;
        RECT 81.675 89.880 82.005 90.390 ;
        RECT 82.175 90.235 84.540 90.405 ;
        RECT 84.885 90.435 85.635 90.955 ;
        RECT 85.805 90.605 86.555 91.125 ;
        RECT 87.185 91.050 87.475 92.215 ;
        RECT 87.665 91.160 87.970 91.945 ;
        RECT 88.150 91.745 88.835 92.215 ;
        RECT 88.145 91.225 88.840 91.535 ;
        RECT 82.175 89.665 82.505 90.065 ;
        RECT 83.555 89.895 83.885 90.235 ;
        RECT 84.055 89.665 84.385 90.065 ;
        RECT 84.885 89.665 86.555 90.435 ;
        RECT 87.185 89.665 87.475 90.390 ;
        RECT 87.665 90.355 87.840 91.160 ;
        RECT 89.015 91.055 89.300 92.000 ;
        RECT 89.475 91.765 89.805 92.215 ;
        RECT 89.975 91.595 90.145 92.025 ;
        RECT 88.440 90.905 89.300 91.055 ;
        RECT 88.015 90.885 89.300 90.905 ;
        RECT 89.470 91.365 90.145 91.595 ;
        RECT 88.015 90.525 89.000 90.885 ;
        RECT 89.470 90.715 89.705 91.365 ;
        RECT 87.665 89.835 87.905 90.355 ;
        RECT 88.830 90.190 89.000 90.525 ;
        RECT 89.170 90.385 89.705 90.715 ;
        RECT 89.485 90.235 89.705 90.385 ;
        RECT 89.875 90.345 90.175 91.195 ;
        RECT 90.405 91.140 90.675 92.045 ;
        RECT 90.845 91.455 91.175 92.215 ;
        RECT 91.355 91.285 91.525 92.045 ;
        RECT 90.405 90.340 90.575 91.140 ;
        RECT 90.860 91.115 91.525 91.285 ;
        RECT 91.785 91.125 93.455 92.215 ;
        RECT 90.860 90.970 91.030 91.115 ;
        RECT 90.745 90.640 91.030 90.970 ;
        RECT 90.860 90.385 91.030 90.640 ;
        RECT 91.265 90.565 91.595 90.935 ;
        RECT 91.785 90.435 92.535 90.955 ;
        RECT 92.705 90.605 93.455 91.125 ;
        RECT 94.090 91.265 94.355 92.035 ;
        RECT 94.525 91.495 94.855 92.215 ;
        RECT 95.045 91.675 95.305 92.035 ;
        RECT 95.475 91.845 95.805 92.215 ;
        RECT 95.975 91.675 96.235 92.035 ;
        RECT 95.045 91.445 96.235 91.675 ;
        RECT 96.805 91.265 97.095 92.035 ;
        RECT 88.075 89.665 88.470 90.160 ;
        RECT 88.830 89.995 89.205 90.190 ;
        RECT 89.035 89.850 89.205 89.995 ;
        RECT 89.485 89.860 89.725 90.235 ;
        RECT 89.895 89.665 90.230 90.170 ;
        RECT 90.405 89.835 90.665 90.340 ;
        RECT 90.860 90.215 91.525 90.385 ;
        RECT 90.845 89.665 91.175 90.045 ;
        RECT 91.355 89.835 91.525 90.215 ;
        RECT 91.785 89.665 93.455 90.435 ;
        RECT 94.090 89.845 94.425 91.265 ;
        RECT 94.600 91.085 97.095 91.265 ;
        RECT 94.600 90.395 94.825 91.085 ;
        RECT 97.825 91.075 98.035 92.215 ;
        RECT 98.205 91.065 98.535 92.045 ;
        RECT 98.705 91.075 98.935 92.215 ;
        RECT 99.145 91.705 99.405 92.215 ;
        RECT 95.025 90.575 95.305 90.905 ;
        RECT 95.485 90.575 96.060 90.905 ;
        RECT 96.240 90.575 96.675 90.905 ;
        RECT 96.855 90.575 97.125 90.905 ;
        RECT 94.600 90.205 97.085 90.395 ;
        RECT 94.605 89.665 95.350 90.035 ;
        RECT 95.915 89.845 96.170 90.205 ;
        RECT 96.350 89.665 96.680 90.035 ;
        RECT 96.860 89.845 97.085 90.205 ;
        RECT 97.825 89.665 98.035 90.485 ;
        RECT 98.205 90.465 98.455 91.065 ;
        RECT 98.625 90.655 98.955 90.905 ;
        RECT 99.145 90.655 99.485 91.535 ;
        RECT 99.655 90.825 99.825 92.045 ;
        RECT 100.065 91.710 100.680 92.215 ;
        RECT 100.065 91.175 100.315 91.540 ;
        RECT 100.485 91.535 100.680 91.710 ;
        RECT 100.850 91.705 101.325 92.045 ;
        RECT 101.495 91.670 101.710 92.215 ;
        RECT 100.485 91.345 100.815 91.535 ;
        RECT 101.035 91.175 101.750 91.470 ;
        RECT 101.920 91.345 102.195 92.045 ;
        RECT 100.065 91.005 101.855 91.175 ;
        RECT 99.655 90.575 100.450 90.825 ;
        RECT 99.655 90.485 99.905 90.575 ;
        RECT 98.205 89.835 98.535 90.465 ;
        RECT 98.705 89.665 98.935 90.485 ;
        RECT 99.145 89.665 99.405 90.485 ;
        RECT 99.575 90.065 99.905 90.485 ;
        RECT 100.620 90.150 100.875 91.005 ;
        RECT 100.085 89.885 100.875 90.150 ;
        RECT 101.045 90.305 101.455 90.825 ;
        RECT 101.625 90.575 101.855 91.005 ;
        RECT 102.025 90.315 102.195 91.345 ;
        RECT 101.045 89.885 101.245 90.305 ;
        RECT 101.435 89.665 101.765 90.125 ;
        RECT 101.935 89.835 102.195 90.315 ;
        RECT 103.285 91.075 103.625 92.045 ;
        RECT 103.795 91.075 103.965 92.215 ;
        RECT 104.235 91.415 104.485 92.215 ;
        RECT 105.130 91.245 105.460 92.045 ;
        RECT 105.760 91.415 106.090 92.215 ;
        RECT 106.260 91.245 106.590 92.045 ;
        RECT 104.155 91.075 106.590 91.245 ;
        RECT 106.965 91.125 108.175 92.215 ;
        RECT 103.285 90.465 103.460 91.075 ;
        RECT 104.155 90.825 104.325 91.075 ;
        RECT 103.630 90.655 104.325 90.825 ;
        RECT 104.500 90.655 104.920 90.855 ;
        RECT 105.090 90.655 105.420 90.855 ;
        RECT 105.590 90.655 105.920 90.855 ;
        RECT 103.285 89.835 103.625 90.465 ;
        RECT 103.795 89.665 104.045 90.465 ;
        RECT 104.235 90.315 105.460 90.485 ;
        RECT 104.235 89.835 104.565 90.315 ;
        RECT 104.735 89.665 104.960 90.125 ;
        RECT 105.130 89.835 105.460 90.315 ;
        RECT 106.090 90.445 106.260 91.075 ;
        RECT 106.445 90.655 106.795 90.905 ;
        RECT 106.090 89.835 106.590 90.445 ;
        RECT 106.965 90.415 107.485 90.955 ;
        RECT 107.655 90.585 108.175 91.125 ;
        RECT 106.965 89.665 108.175 90.415 ;
        RECT 108.355 89.845 108.615 92.035 ;
        RECT 108.785 91.485 109.125 92.215 ;
        RECT 109.305 91.305 109.575 92.035 ;
        RECT 108.805 91.085 109.575 91.305 ;
        RECT 109.755 91.325 109.985 92.035 ;
        RECT 110.155 91.505 110.485 92.215 ;
        RECT 110.655 91.325 110.915 92.035 ;
        RECT 109.755 91.085 110.915 91.325 ;
        RECT 108.805 90.415 109.095 91.085 ;
        RECT 111.105 91.075 111.365 92.215 ;
        RECT 111.535 91.065 111.865 92.045 ;
        RECT 112.035 91.075 112.315 92.215 ;
        RECT 109.275 90.595 109.740 90.905 ;
        RECT 109.920 90.595 110.445 90.905 ;
        RECT 108.805 90.215 110.035 90.415 ;
        RECT 108.875 89.665 109.545 90.035 ;
        RECT 109.725 89.845 110.035 90.215 ;
        RECT 110.215 89.955 110.445 90.595 ;
        RECT 110.625 90.575 110.925 90.905 ;
        RECT 111.125 90.655 111.460 90.905 ;
        RECT 111.630 90.465 111.800 91.065 ;
        RECT 112.945 91.050 113.235 92.215 ;
        RECT 113.405 91.345 113.680 92.045 ;
        RECT 113.850 91.670 114.105 92.215 ;
        RECT 114.275 91.705 114.755 92.045 ;
        RECT 114.930 91.660 115.535 92.215 ;
        RECT 114.920 91.560 115.535 91.660 ;
        RECT 114.920 91.535 115.105 91.560 ;
        RECT 111.970 90.635 112.305 90.905 ;
        RECT 110.625 89.665 110.915 90.395 ;
        RECT 111.105 89.835 111.800 90.465 ;
        RECT 112.005 89.665 112.315 90.465 ;
        RECT 112.945 89.665 113.235 90.390 ;
        RECT 113.405 90.315 113.575 91.345 ;
        RECT 113.850 91.215 114.605 91.465 ;
        RECT 114.775 91.290 115.105 91.535 ;
        RECT 113.850 91.180 114.620 91.215 ;
        RECT 113.850 91.170 114.635 91.180 ;
        RECT 113.745 91.155 114.640 91.170 ;
        RECT 113.745 91.140 114.660 91.155 ;
        RECT 113.745 91.130 114.680 91.140 ;
        RECT 113.745 91.120 114.705 91.130 ;
        RECT 113.745 91.090 114.775 91.120 ;
        RECT 113.745 91.060 114.795 91.090 ;
        RECT 113.745 91.030 114.815 91.060 ;
        RECT 113.745 91.005 114.845 91.030 ;
        RECT 113.745 90.970 114.880 91.005 ;
        RECT 113.745 90.965 114.910 90.970 ;
        RECT 113.745 90.570 113.975 90.965 ;
        RECT 114.520 90.960 114.910 90.965 ;
        RECT 114.545 90.950 114.910 90.960 ;
        RECT 114.560 90.945 114.910 90.950 ;
        RECT 114.575 90.940 114.910 90.945 ;
        RECT 115.275 90.940 115.535 91.390 ;
        RECT 115.705 91.125 116.915 92.215 ;
        RECT 117.115 91.755 117.375 92.215 ;
        RECT 114.575 90.935 115.535 90.940 ;
        RECT 114.585 90.925 115.535 90.935 ;
        RECT 114.595 90.920 115.535 90.925 ;
        RECT 114.605 90.910 115.535 90.920 ;
        RECT 114.610 90.900 115.535 90.910 ;
        RECT 114.615 90.895 115.535 90.900 ;
        RECT 114.625 90.880 115.535 90.895 ;
        RECT 114.630 90.865 115.535 90.880 ;
        RECT 114.640 90.840 115.535 90.865 ;
        RECT 114.145 90.370 114.475 90.795 ;
        RECT 113.405 89.835 113.665 90.315 ;
        RECT 113.835 89.665 114.085 90.205 ;
        RECT 114.255 89.885 114.475 90.370 ;
        RECT 114.645 90.770 115.535 90.840 ;
        RECT 114.645 90.045 114.815 90.770 ;
        RECT 114.985 90.215 115.535 90.600 ;
        RECT 115.705 90.415 116.225 90.955 ;
        RECT 116.395 90.585 116.915 91.125 ;
        RECT 117.085 90.575 117.375 91.550 ;
        RECT 117.545 91.290 117.805 92.045 ;
        RECT 117.975 91.495 118.305 92.215 ;
        RECT 118.475 91.290 118.665 92.045 ;
        RECT 118.835 91.495 119.165 92.215 ;
        RECT 119.395 91.875 120.515 92.045 ;
        RECT 119.395 91.680 119.655 91.875 ;
        RECT 119.825 91.290 120.155 91.705 ;
        RECT 117.545 91.120 120.155 91.290 ;
        RECT 120.325 91.275 120.515 91.875 ;
        RECT 120.685 91.445 121.015 92.215 ;
        RECT 121.185 91.275 121.445 92.045 ;
        RECT 114.645 89.875 115.535 90.045 ;
        RECT 115.705 89.665 116.915 90.415 ;
        RECT 117.545 90.250 117.875 91.120 ;
        RECT 120.325 91.105 121.445 91.275 ;
        RECT 121.685 91.125 125.195 92.215 ;
        RECT 125.365 91.125 126.575 92.215 ;
        RECT 118.045 90.655 118.905 90.945 ;
        RECT 119.365 90.655 120.335 90.935 ;
        RECT 120.560 90.825 121.455 90.875 ;
        RECT 120.505 90.655 121.455 90.825 ;
        RECT 118.045 90.045 118.235 90.470 ;
        RECT 118.405 90.215 120.945 90.425 ;
        RECT 121.115 90.345 121.455 90.655 ;
        RECT 121.685 90.435 123.335 90.955 ;
        RECT 123.505 90.605 125.195 91.125 ;
        RECT 120.755 90.095 120.945 90.215 ;
        RECT 118.045 90.025 119.165 90.045 ;
        RECT 117.095 89.835 119.165 90.025 ;
        RECT 119.395 89.665 119.725 90.025 ;
        RECT 120.255 89.665 120.585 90.025 ;
        RECT 121.115 89.665 121.445 90.025 ;
        RECT 121.685 89.665 125.195 90.435 ;
        RECT 125.365 90.415 125.885 90.955 ;
        RECT 126.055 90.585 126.575 91.125 ;
        RECT 126.755 91.605 127.085 92.035 ;
        RECT 127.265 91.775 127.460 92.215 ;
        RECT 127.630 91.605 127.960 92.035 ;
        RECT 126.755 91.435 127.960 91.605 ;
        RECT 126.755 91.105 127.650 91.435 ;
        RECT 128.130 91.265 128.405 92.035 ;
        RECT 127.820 91.075 128.405 91.265 ;
        RECT 128.595 91.155 128.925 92.005 ;
        RECT 126.760 90.575 127.055 90.905 ;
        RECT 127.235 90.575 127.650 90.905 ;
        RECT 125.365 89.665 126.575 90.415 ;
        RECT 126.755 89.665 127.055 90.395 ;
        RECT 127.235 89.955 127.465 90.575 ;
        RECT 127.820 90.405 127.995 91.075 ;
        RECT 127.665 90.225 127.995 90.405 ;
        RECT 128.165 90.255 128.405 90.905 ;
        RECT 128.595 90.390 128.785 91.155 ;
        RECT 129.095 91.075 129.345 92.215 ;
        RECT 129.535 91.575 129.785 91.995 ;
        RECT 130.015 91.745 130.345 92.215 ;
        RECT 130.575 91.575 130.825 91.995 ;
        RECT 129.535 91.405 130.825 91.575 ;
        RECT 131.005 91.575 131.335 92.005 ;
        RECT 131.005 91.405 131.460 91.575 ;
        RECT 129.525 90.905 129.740 91.235 ;
        RECT 128.955 90.575 129.265 90.905 ;
        RECT 129.435 90.575 129.740 90.905 ;
        RECT 129.915 90.575 130.200 91.235 ;
        RECT 130.395 90.575 130.660 91.235 ;
        RECT 130.875 90.575 131.120 91.235 ;
        RECT 129.095 90.405 129.265 90.575 ;
        RECT 131.290 90.405 131.460 91.405 ;
        RECT 131.805 91.125 134.395 92.215 ;
        RECT 127.665 89.845 127.890 90.225 ;
        RECT 128.060 89.665 128.390 90.055 ;
        RECT 128.595 89.880 128.925 90.390 ;
        RECT 129.095 90.235 131.460 90.405 ;
        RECT 131.805 90.435 133.015 90.955 ;
        RECT 133.185 90.605 134.395 91.125 ;
        RECT 135.030 91.265 135.295 92.035 ;
        RECT 135.465 91.495 135.795 92.215 ;
        RECT 135.985 91.675 136.245 92.035 ;
        RECT 136.415 91.845 136.745 92.215 ;
        RECT 136.915 91.675 137.175 92.035 ;
        RECT 135.985 91.445 137.175 91.675 ;
        RECT 137.745 91.265 138.035 92.035 ;
        RECT 129.095 89.665 129.425 90.065 ;
        RECT 130.475 89.895 130.805 90.235 ;
        RECT 130.975 89.665 131.305 90.065 ;
        RECT 131.805 89.665 134.395 90.435 ;
        RECT 135.030 89.845 135.365 91.265 ;
        RECT 135.540 91.085 138.035 91.265 ;
        RECT 135.540 90.395 135.765 91.085 ;
        RECT 138.705 91.050 138.995 92.215 ;
        RECT 139.165 91.125 141.755 92.215 ;
        RECT 135.965 90.575 136.245 90.905 ;
        RECT 136.425 90.575 137.000 90.905 ;
        RECT 137.180 90.575 137.615 90.905 ;
        RECT 137.795 90.575 138.065 90.905 ;
        RECT 139.165 90.435 140.375 90.955 ;
        RECT 140.545 90.605 141.755 91.125 ;
        RECT 142.015 91.285 142.185 92.045 ;
        RECT 142.365 91.455 142.695 92.215 ;
        RECT 142.015 91.115 142.680 91.285 ;
        RECT 142.865 91.140 143.135 92.045 ;
        RECT 143.395 91.545 143.565 92.045 ;
        RECT 143.735 91.715 144.065 92.215 ;
        RECT 143.395 91.375 144.060 91.545 ;
        RECT 142.510 90.970 142.680 91.115 ;
        RECT 141.945 90.565 142.275 90.935 ;
        RECT 142.510 90.640 142.795 90.970 ;
        RECT 135.540 90.205 138.025 90.395 ;
        RECT 135.545 89.665 136.290 90.035 ;
        RECT 136.855 89.845 137.110 90.205 ;
        RECT 137.290 89.665 137.620 90.035 ;
        RECT 137.800 89.845 138.025 90.205 ;
        RECT 138.705 89.665 138.995 90.390 ;
        RECT 139.165 89.665 141.755 90.435 ;
        RECT 142.510 90.385 142.680 90.640 ;
        RECT 142.015 90.215 142.680 90.385 ;
        RECT 142.965 90.340 143.135 91.140 ;
        RECT 143.310 90.555 143.660 91.205 ;
        RECT 143.830 90.385 144.060 91.375 ;
        RECT 142.015 89.835 142.185 90.215 ;
        RECT 142.365 89.665 142.695 90.045 ;
        RECT 142.875 89.835 143.135 90.340 ;
        RECT 143.395 90.215 144.060 90.385 ;
        RECT 143.395 89.925 143.565 90.215 ;
        RECT 143.735 89.665 144.065 90.045 ;
        RECT 144.235 89.925 144.420 92.045 ;
        RECT 144.660 91.755 144.925 92.215 ;
        RECT 145.095 91.620 145.345 92.045 ;
        RECT 145.555 91.770 146.660 91.940 ;
        RECT 145.040 91.490 145.345 91.620 ;
        RECT 144.590 90.295 144.870 91.245 ;
        RECT 145.040 90.385 145.210 91.490 ;
        RECT 145.380 90.705 145.620 91.300 ;
        RECT 145.790 91.235 146.320 91.600 ;
        RECT 145.790 90.535 145.960 91.235 ;
        RECT 146.490 91.155 146.660 91.770 ;
        RECT 146.830 91.415 147.000 92.215 ;
        RECT 147.170 91.715 147.420 92.045 ;
        RECT 147.645 91.745 148.530 91.915 ;
        RECT 146.490 91.065 147.000 91.155 ;
        RECT 145.040 90.255 145.265 90.385 ;
        RECT 145.435 90.315 145.960 90.535 ;
        RECT 146.130 90.895 147.000 91.065 ;
        RECT 144.675 89.665 144.925 90.125 ;
        RECT 145.095 90.115 145.265 90.255 ;
        RECT 146.130 90.115 146.300 90.895 ;
        RECT 146.830 90.825 147.000 90.895 ;
        RECT 146.510 90.645 146.710 90.675 ;
        RECT 147.170 90.645 147.340 91.715 ;
        RECT 147.510 90.825 147.700 91.545 ;
        RECT 146.510 90.345 147.340 90.645 ;
        RECT 147.870 90.615 148.190 91.575 ;
        RECT 145.095 89.945 145.430 90.115 ;
        RECT 145.625 89.945 146.300 90.115 ;
        RECT 146.620 89.665 146.990 90.165 ;
        RECT 147.170 90.115 147.340 90.345 ;
        RECT 147.725 90.285 148.190 90.615 ;
        RECT 148.360 90.905 148.530 91.745 ;
        RECT 148.710 91.715 149.025 92.215 ;
        RECT 149.255 91.485 149.595 92.045 ;
        RECT 148.700 91.110 149.595 91.485 ;
        RECT 149.765 91.205 149.935 92.215 ;
        RECT 149.405 90.905 149.595 91.110 ;
        RECT 150.105 91.155 150.435 92.000 ;
        RECT 150.105 91.075 150.495 91.155 ;
        RECT 150.280 91.025 150.495 91.075 ;
        RECT 148.360 90.575 149.235 90.905 ;
        RECT 149.405 90.575 150.155 90.905 ;
        RECT 148.360 90.115 148.530 90.575 ;
        RECT 149.405 90.405 149.605 90.575 ;
        RECT 150.325 90.445 150.495 91.025 ;
        RECT 150.270 90.405 150.495 90.445 ;
        RECT 147.170 89.945 147.575 90.115 ;
        RECT 147.745 89.945 148.530 90.115 ;
        RECT 148.805 89.665 149.015 90.195 ;
        RECT 149.275 89.880 149.605 90.405 ;
        RECT 150.115 90.320 150.495 90.405 ;
        RECT 151.585 91.075 151.970 92.045 ;
        RECT 152.140 91.755 152.465 92.215 ;
        RECT 152.985 91.585 153.265 92.045 ;
        RECT 152.140 91.365 153.265 91.585 ;
        RECT 151.585 90.405 151.865 91.075 ;
        RECT 152.140 90.905 152.590 91.365 ;
        RECT 153.455 91.195 153.855 92.045 ;
        RECT 154.255 91.755 154.525 92.215 ;
        RECT 154.695 91.585 154.980 92.045 ;
        RECT 152.035 90.575 152.590 90.905 ;
        RECT 152.760 90.635 153.855 91.195 ;
        RECT 152.140 90.465 152.590 90.575 ;
        RECT 149.775 89.665 149.945 90.275 ;
        RECT 150.115 89.885 150.445 90.320 ;
        RECT 151.585 89.835 151.970 90.405 ;
        RECT 152.140 90.295 153.265 90.465 ;
        RECT 152.140 89.665 152.465 90.125 ;
        RECT 152.985 89.835 153.265 90.295 ;
        RECT 153.455 89.835 153.855 90.635 ;
        RECT 154.025 91.365 154.980 91.585 ;
        RECT 154.025 90.465 154.235 91.365 ;
        RECT 154.405 90.635 155.095 91.195 ;
        RECT 155.725 91.125 156.935 92.215 ;
        RECT 155.725 90.585 156.245 91.125 ;
        RECT 154.025 90.295 154.980 90.465 ;
        RECT 156.415 90.415 156.935 90.955 ;
        RECT 154.255 89.665 154.525 90.125 ;
        RECT 154.695 89.835 154.980 90.295 ;
        RECT 155.725 89.665 156.935 90.415 ;
        RECT 22.700 89.495 157.020 89.665 ;
        RECT 22.785 88.745 23.995 89.495 ;
        RECT 24.165 88.950 29.510 89.495 ;
        RECT 22.785 88.205 23.305 88.745 ;
        RECT 23.475 88.035 23.995 88.575 ;
        RECT 25.750 88.120 26.090 88.950 ;
        RECT 30.155 88.685 30.425 89.495 ;
        RECT 30.595 88.685 30.925 89.325 ;
        RECT 31.095 88.685 31.335 89.495 ;
        RECT 31.525 88.695 31.835 89.495 ;
        RECT 32.040 88.695 32.735 89.325 ;
        RECT 32.905 88.695 33.245 89.325 ;
        RECT 33.415 88.695 33.665 89.495 ;
        RECT 33.855 88.845 34.185 89.325 ;
        RECT 34.355 89.035 34.580 89.495 ;
        RECT 34.750 88.845 35.080 89.325 ;
        RECT 22.785 86.945 23.995 88.035 ;
        RECT 27.570 87.380 27.920 88.630 ;
        RECT 30.145 88.255 30.495 88.505 ;
        RECT 30.665 88.085 30.835 88.685 ;
        RECT 32.040 88.645 32.215 88.695 ;
        RECT 31.005 88.255 31.355 88.505 ;
        RECT 31.535 88.255 31.870 88.525 ;
        RECT 32.040 88.095 32.210 88.645 ;
        RECT 32.380 88.255 32.715 88.505 ;
        RECT 32.905 88.135 33.080 88.695 ;
        RECT 33.855 88.675 35.080 88.845 ;
        RECT 35.710 88.715 36.210 89.325 ;
        RECT 36.610 89.105 36.940 89.495 ;
        RECT 37.110 88.935 37.335 89.315 ;
        RECT 33.250 88.335 33.945 88.505 ;
        RECT 24.165 86.945 29.510 87.380 ;
        RECT 30.155 86.945 30.485 88.085 ;
        RECT 30.665 87.915 31.345 88.085 ;
        RECT 31.015 87.130 31.345 87.915 ;
        RECT 31.525 86.945 31.805 88.085 ;
        RECT 31.975 87.115 32.305 88.095 ;
        RECT 32.905 88.085 33.135 88.135 ;
        RECT 33.775 88.085 33.945 88.335 ;
        RECT 34.120 88.305 34.540 88.505 ;
        RECT 34.710 88.305 35.040 88.505 ;
        RECT 35.210 88.305 35.540 88.505 ;
        RECT 35.710 88.085 35.880 88.715 ;
        RECT 36.065 88.255 36.415 88.505 ;
        RECT 36.595 88.255 36.835 88.905 ;
        RECT 37.005 88.755 37.335 88.935 ;
        RECT 37.005 88.085 37.180 88.755 ;
        RECT 37.535 88.585 37.765 89.205 ;
        RECT 37.945 88.765 38.245 89.495 ;
        RECT 38.425 88.725 40.095 89.495 ;
        RECT 40.265 89.035 40.825 89.325 ;
        RECT 40.995 89.035 41.245 89.495 ;
        RECT 37.350 88.255 37.765 88.585 ;
        RECT 37.945 88.255 38.240 88.585 ;
        RECT 38.425 88.205 39.175 88.725 ;
        RECT 32.475 86.945 32.735 88.085 ;
        RECT 32.905 87.115 33.245 88.085 ;
        RECT 33.415 86.945 33.585 88.085 ;
        RECT 33.775 87.915 36.210 88.085 ;
        RECT 33.855 86.945 34.105 87.745 ;
        RECT 34.750 87.115 35.080 87.915 ;
        RECT 35.380 86.945 35.710 87.745 ;
        RECT 35.880 87.115 36.210 87.915 ;
        RECT 36.595 87.895 37.180 88.085 ;
        RECT 36.595 87.125 36.870 87.895 ;
        RECT 37.350 87.725 38.245 88.055 ;
        RECT 39.345 88.035 40.095 88.555 ;
        RECT 37.040 87.555 38.245 87.725 ;
        RECT 37.040 87.125 37.370 87.555 ;
        RECT 37.540 86.945 37.735 87.385 ;
        RECT 37.915 87.125 38.245 87.555 ;
        RECT 38.425 86.945 40.095 88.035 ;
        RECT 40.265 87.665 40.515 89.035 ;
        RECT 41.865 88.865 42.195 89.225 ;
        RECT 40.805 88.675 42.195 88.865 ;
        RECT 42.565 88.735 43.275 89.325 ;
        RECT 43.785 88.965 44.115 89.325 ;
        RECT 44.315 89.135 44.645 89.495 ;
        RECT 44.815 88.965 45.145 89.325 ;
        RECT 45.490 88.985 45.730 89.495 ;
        RECT 45.910 88.985 46.190 89.315 ;
        RECT 46.420 88.985 46.635 89.495 ;
        RECT 43.785 88.755 45.145 88.965 ;
        RECT 40.805 88.585 40.975 88.675 ;
        RECT 40.685 88.255 40.975 88.585 ;
        RECT 42.565 88.645 42.795 88.735 ;
        RECT 41.145 88.255 41.485 88.505 ;
        RECT 41.705 88.255 42.380 88.505 ;
        RECT 40.805 88.005 40.975 88.255 ;
        RECT 40.805 87.835 41.745 88.005 ;
        RECT 42.115 87.895 42.380 88.255 ;
        RECT 40.265 87.115 40.725 87.665 ;
        RECT 40.915 86.945 41.245 87.665 ;
        RECT 41.445 87.285 41.745 87.835 ;
        RECT 42.565 87.765 42.770 88.645 ;
        RECT 42.940 87.965 43.270 88.505 ;
        RECT 43.445 88.255 43.940 88.585 ;
        RECT 44.260 88.255 44.635 88.585 ;
        RECT 44.845 88.255 45.155 88.585 ;
        RECT 45.385 88.255 45.740 88.815 ;
        RECT 43.445 87.965 43.770 88.255 ;
        RECT 43.965 87.765 44.295 87.985 ;
        RECT 41.915 86.945 42.195 87.615 ;
        RECT 42.565 87.535 44.295 87.765 ;
        RECT 42.565 87.115 43.265 87.535 ;
        RECT 43.465 86.945 43.795 87.305 ;
        RECT 43.965 87.135 44.295 87.535 ;
        RECT 44.465 87.330 44.635 88.255 ;
        RECT 45.910 88.085 46.080 88.985 ;
        RECT 46.250 88.255 46.515 88.815 ;
        RECT 46.805 88.755 47.420 89.325 ;
        RECT 48.545 88.770 48.835 89.495 ;
        RECT 46.765 88.085 46.935 88.585 ;
        RECT 44.815 86.945 45.145 88.005 ;
        RECT 45.510 87.915 46.935 88.085 ;
        RECT 45.510 87.740 45.900 87.915 ;
        RECT 46.385 86.945 46.715 87.745 ;
        RECT 47.105 87.735 47.420 88.755 ;
        RECT 46.885 87.115 47.420 87.735 ;
        RECT 48.545 86.945 48.835 88.110 ;
        RECT 49.930 87.895 50.265 89.315 ;
        RECT 50.445 89.125 51.190 89.495 ;
        RECT 51.755 88.955 52.010 89.315 ;
        RECT 52.190 89.125 52.520 89.495 ;
        RECT 52.700 88.955 52.925 89.315 ;
        RECT 53.310 88.985 53.550 89.495 ;
        RECT 53.730 88.985 54.010 89.315 ;
        RECT 54.240 88.985 54.455 89.495 ;
        RECT 50.440 88.765 52.925 88.955 ;
        RECT 50.440 88.075 50.665 88.765 ;
        RECT 50.865 88.255 51.145 88.585 ;
        RECT 51.325 88.255 51.900 88.585 ;
        RECT 52.080 88.255 52.515 88.585 ;
        RECT 52.695 88.255 52.965 88.585 ;
        RECT 53.205 88.255 53.560 88.815 ;
        RECT 53.730 88.085 53.900 88.985 ;
        RECT 54.070 88.255 54.335 88.815 ;
        RECT 54.625 88.755 55.240 89.325 ;
        RECT 54.585 88.085 54.755 88.585 ;
        RECT 50.440 87.895 52.935 88.075 ;
        RECT 49.930 87.125 50.195 87.895 ;
        RECT 50.365 86.945 50.695 87.665 ;
        RECT 50.885 87.485 52.075 87.715 ;
        RECT 50.885 87.125 51.145 87.485 ;
        RECT 51.315 86.945 51.645 87.315 ;
        RECT 51.815 87.125 52.075 87.485 ;
        RECT 52.645 87.125 52.935 87.895 ;
        RECT 53.330 87.915 54.755 88.085 ;
        RECT 53.330 87.740 53.720 87.915 ;
        RECT 54.205 86.945 54.535 87.745 ;
        RECT 54.925 87.735 55.240 88.755 ;
        RECT 55.445 88.725 57.115 89.495 ;
        RECT 57.285 88.845 57.545 89.325 ;
        RECT 57.715 89.035 58.045 89.495 ;
        RECT 58.235 88.855 58.435 89.275 ;
        RECT 55.445 88.205 56.195 88.725 ;
        RECT 56.365 88.035 57.115 88.555 ;
        RECT 54.705 87.115 55.240 87.735 ;
        RECT 55.445 86.945 57.115 88.035 ;
        RECT 57.285 87.815 57.455 88.845 ;
        RECT 57.625 88.155 57.855 88.585 ;
        RECT 58.025 88.335 58.435 88.855 ;
        RECT 58.605 89.010 59.395 89.275 ;
        RECT 58.605 88.155 58.860 89.010 ;
        RECT 59.575 88.675 59.905 89.095 ;
        RECT 60.075 88.675 60.335 89.495 ;
        RECT 60.505 88.950 65.850 89.495 ;
        RECT 66.025 88.950 71.370 89.495 ;
        RECT 59.575 88.585 59.825 88.675 ;
        RECT 59.030 88.335 59.825 88.585 ;
        RECT 57.625 87.985 59.415 88.155 ;
        RECT 57.285 87.115 57.560 87.815 ;
        RECT 57.730 87.690 58.445 87.985 ;
        RECT 58.665 87.625 58.995 87.815 ;
        RECT 57.770 86.945 57.985 87.490 ;
        RECT 58.155 87.115 58.630 87.455 ;
        RECT 58.800 87.450 58.995 87.625 ;
        RECT 59.165 87.620 59.415 87.985 ;
        RECT 58.800 86.945 59.415 87.450 ;
        RECT 59.655 87.115 59.825 88.335 ;
        RECT 59.995 87.625 60.335 88.505 ;
        RECT 62.090 88.120 62.430 88.950 ;
        RECT 60.075 86.945 60.335 87.455 ;
        RECT 63.910 87.380 64.260 88.630 ;
        RECT 67.610 88.120 67.950 88.950 ;
        RECT 71.545 88.725 74.135 89.495 ;
        RECT 74.305 88.770 74.595 89.495 ;
        RECT 74.855 88.945 75.025 89.235 ;
        RECT 75.195 89.115 75.525 89.495 ;
        RECT 74.855 88.775 75.520 88.945 ;
        RECT 69.430 87.380 69.780 88.630 ;
        RECT 71.545 88.205 72.755 88.725 ;
        RECT 72.925 88.035 74.135 88.555 ;
        RECT 60.505 86.945 65.850 87.380 ;
        RECT 66.025 86.945 71.370 87.380 ;
        RECT 71.545 86.945 74.135 88.035 ;
        RECT 74.305 86.945 74.595 88.110 ;
        RECT 74.770 87.955 75.120 88.605 ;
        RECT 75.290 87.785 75.520 88.775 ;
        RECT 74.855 87.615 75.520 87.785 ;
        RECT 74.855 87.115 75.025 87.615 ;
        RECT 75.195 86.945 75.525 87.445 ;
        RECT 75.695 87.115 75.880 89.235 ;
        RECT 76.135 89.035 76.385 89.495 ;
        RECT 76.555 89.045 76.890 89.215 ;
        RECT 77.085 89.045 77.760 89.215 ;
        RECT 76.555 88.905 76.725 89.045 ;
        RECT 76.050 87.915 76.330 88.865 ;
        RECT 76.500 88.775 76.725 88.905 ;
        RECT 76.500 87.670 76.670 88.775 ;
        RECT 76.895 88.625 77.420 88.845 ;
        RECT 76.840 87.860 77.080 88.455 ;
        RECT 77.250 87.925 77.420 88.625 ;
        RECT 77.590 88.265 77.760 89.045 ;
        RECT 78.080 88.995 78.450 89.495 ;
        RECT 78.630 89.045 79.035 89.215 ;
        RECT 79.205 89.045 79.990 89.215 ;
        RECT 78.630 88.815 78.800 89.045 ;
        RECT 77.970 88.515 78.800 88.815 ;
        RECT 79.185 88.545 79.650 88.875 ;
        RECT 77.970 88.485 78.170 88.515 ;
        RECT 78.290 88.265 78.460 88.335 ;
        RECT 77.590 88.095 78.460 88.265 ;
        RECT 77.950 88.005 78.460 88.095 ;
        RECT 76.500 87.540 76.805 87.670 ;
        RECT 77.250 87.560 77.780 87.925 ;
        RECT 76.120 86.945 76.385 87.405 ;
        RECT 76.555 87.115 76.805 87.540 ;
        RECT 77.950 87.390 78.120 88.005 ;
        RECT 77.015 87.220 78.120 87.390 ;
        RECT 78.290 86.945 78.460 87.745 ;
        RECT 78.630 87.445 78.800 88.515 ;
        RECT 78.970 87.615 79.160 88.335 ;
        RECT 79.330 87.585 79.650 88.545 ;
        RECT 79.820 88.585 79.990 89.045 ;
        RECT 80.265 88.965 80.475 89.495 ;
        RECT 80.735 88.755 81.065 89.280 ;
        RECT 81.235 88.885 81.405 89.495 ;
        RECT 81.575 88.840 81.905 89.275 ;
        RECT 82.290 88.985 82.530 89.495 ;
        RECT 82.710 88.985 82.990 89.315 ;
        RECT 83.220 88.985 83.435 89.495 ;
        RECT 81.575 88.755 81.955 88.840 ;
        RECT 80.865 88.585 81.065 88.755 ;
        RECT 81.730 88.715 81.955 88.755 ;
        RECT 79.820 88.255 80.695 88.585 ;
        RECT 80.865 88.255 81.615 88.585 ;
        RECT 78.630 87.115 78.880 87.445 ;
        RECT 79.820 87.415 79.990 88.255 ;
        RECT 80.865 88.050 81.055 88.255 ;
        RECT 81.785 88.135 81.955 88.715 ;
        RECT 82.185 88.255 82.540 88.815 ;
        RECT 81.740 88.085 81.955 88.135 ;
        RECT 82.710 88.085 82.880 88.985 ;
        RECT 83.050 88.255 83.315 88.815 ;
        RECT 83.605 88.755 84.220 89.325 ;
        RECT 85.435 88.945 85.605 89.325 ;
        RECT 85.785 89.115 86.115 89.495 ;
        RECT 85.435 88.775 86.100 88.945 ;
        RECT 86.295 88.820 86.555 89.325 ;
        RECT 83.565 88.085 83.735 88.585 ;
        RECT 80.160 87.675 81.055 88.050 ;
        RECT 81.565 88.005 81.955 88.085 ;
        RECT 79.105 87.245 79.990 87.415 ;
        RECT 80.170 86.945 80.485 87.445 ;
        RECT 80.715 87.115 81.055 87.675 ;
        RECT 81.225 86.945 81.395 87.955 ;
        RECT 81.565 87.160 81.895 88.005 ;
        RECT 82.310 87.915 83.735 88.085 ;
        RECT 82.310 87.740 82.700 87.915 ;
        RECT 83.185 86.945 83.515 87.745 ;
        RECT 83.905 87.735 84.220 88.755 ;
        RECT 85.365 88.225 85.695 88.595 ;
        RECT 85.930 88.520 86.100 88.775 ;
        RECT 85.930 88.190 86.215 88.520 ;
        RECT 85.930 88.045 86.100 88.190 ;
        RECT 83.685 87.115 84.220 87.735 ;
        RECT 85.435 87.875 86.100 88.045 ;
        RECT 86.385 88.020 86.555 88.820 ;
        RECT 87.645 88.695 87.955 89.495 ;
        RECT 88.160 88.695 88.855 89.325 ;
        RECT 89.025 88.950 94.370 89.495 ;
        RECT 94.545 88.950 99.890 89.495 ;
        RECT 87.655 88.255 87.990 88.525 ;
        RECT 88.160 88.095 88.330 88.695 ;
        RECT 88.500 88.255 88.835 88.505 ;
        RECT 90.610 88.120 90.950 88.950 ;
        RECT 85.435 87.115 85.605 87.875 ;
        RECT 85.785 86.945 86.115 87.705 ;
        RECT 86.285 87.115 86.555 88.020 ;
        RECT 87.645 86.945 87.925 88.085 ;
        RECT 88.095 87.115 88.425 88.095 ;
        RECT 88.595 86.945 88.855 88.085 ;
        RECT 92.430 87.380 92.780 88.630 ;
        RECT 96.130 88.120 96.470 88.950 ;
        RECT 100.065 88.770 100.355 89.495 ;
        RECT 100.525 88.725 102.195 89.495 ;
        RECT 97.950 87.380 98.300 88.630 ;
        RECT 100.525 88.205 101.275 88.725 ;
        RECT 89.025 86.945 94.370 87.380 ;
        RECT 94.545 86.945 99.890 87.380 ;
        RECT 100.065 86.945 100.355 88.110 ;
        RECT 101.445 88.035 102.195 88.555 ;
        RECT 100.525 86.945 102.195 88.035 ;
        RECT 102.370 87.895 102.705 89.315 ;
        RECT 102.885 89.125 103.630 89.495 ;
        RECT 104.195 88.955 104.450 89.315 ;
        RECT 104.630 89.125 104.960 89.495 ;
        RECT 105.140 88.955 105.365 89.315 ;
        RECT 102.880 88.765 105.365 88.955 ;
        RECT 102.880 88.075 103.105 88.765 ;
        RECT 105.645 88.675 105.855 89.495 ;
        RECT 106.025 88.695 106.355 89.325 ;
        RECT 103.305 88.255 103.585 88.585 ;
        RECT 103.765 88.255 104.340 88.585 ;
        RECT 104.520 88.255 104.955 88.585 ;
        RECT 105.135 88.255 105.405 88.585 ;
        RECT 106.025 88.095 106.275 88.695 ;
        RECT 106.525 88.675 106.755 89.495 ;
        RECT 107.000 88.755 107.615 89.325 ;
        RECT 107.785 88.985 108.000 89.495 ;
        RECT 108.230 88.985 108.510 89.315 ;
        RECT 108.690 88.985 108.930 89.495 ;
        RECT 106.445 88.255 106.775 88.505 ;
        RECT 102.880 87.895 105.375 88.075 ;
        RECT 102.370 87.125 102.635 87.895 ;
        RECT 102.805 86.945 103.135 87.665 ;
        RECT 103.325 87.485 104.515 87.715 ;
        RECT 103.325 87.125 103.585 87.485 ;
        RECT 103.755 86.945 104.085 87.315 ;
        RECT 104.255 87.125 104.515 87.485 ;
        RECT 105.085 87.125 105.375 87.895 ;
        RECT 105.645 86.945 105.855 88.085 ;
        RECT 106.025 87.115 106.355 88.095 ;
        RECT 106.525 86.945 106.755 88.085 ;
        RECT 107.000 87.735 107.315 88.755 ;
        RECT 107.485 88.085 107.655 88.585 ;
        RECT 107.905 88.255 108.170 88.815 ;
        RECT 108.340 88.085 108.510 88.985 ;
        RECT 109.355 88.945 109.525 89.325 ;
        RECT 109.705 89.115 110.035 89.495 ;
        RECT 108.680 88.255 109.035 88.815 ;
        RECT 109.355 88.775 110.020 88.945 ;
        RECT 110.215 88.820 110.475 89.325 ;
        RECT 109.285 88.225 109.615 88.595 ;
        RECT 109.850 88.520 110.020 88.775 ;
        RECT 109.850 88.190 110.135 88.520 ;
        RECT 107.485 87.915 108.910 88.085 ;
        RECT 109.850 88.045 110.020 88.190 ;
        RECT 107.000 87.115 107.535 87.735 ;
        RECT 107.705 86.945 108.035 87.745 ;
        RECT 108.520 87.740 108.910 87.915 ;
        RECT 109.355 87.875 110.020 88.045 ;
        RECT 110.305 88.020 110.475 88.820 ;
        RECT 110.735 88.945 110.905 89.235 ;
        RECT 111.075 89.115 111.405 89.495 ;
        RECT 110.735 88.775 111.400 88.945 ;
        RECT 109.355 87.115 109.525 87.875 ;
        RECT 109.705 86.945 110.035 87.705 ;
        RECT 110.205 87.115 110.475 88.020 ;
        RECT 110.650 87.955 111.000 88.605 ;
        RECT 111.170 87.785 111.400 88.775 ;
        RECT 110.735 87.615 111.400 87.785 ;
        RECT 110.735 87.115 110.905 87.615 ;
        RECT 111.075 86.945 111.405 87.445 ;
        RECT 111.575 87.115 111.760 89.235 ;
        RECT 112.015 89.035 112.265 89.495 ;
        RECT 112.435 89.045 112.770 89.215 ;
        RECT 112.965 89.045 113.640 89.215 ;
        RECT 112.435 88.905 112.605 89.045 ;
        RECT 111.930 87.915 112.210 88.865 ;
        RECT 112.380 88.775 112.605 88.905 ;
        RECT 112.380 87.670 112.550 88.775 ;
        RECT 112.775 88.625 113.300 88.845 ;
        RECT 112.720 87.860 112.960 88.455 ;
        RECT 113.130 87.925 113.300 88.625 ;
        RECT 113.470 88.265 113.640 89.045 ;
        RECT 113.960 88.995 114.330 89.495 ;
        RECT 114.510 89.045 114.915 89.215 ;
        RECT 115.085 89.045 115.870 89.215 ;
        RECT 114.510 88.815 114.680 89.045 ;
        RECT 113.850 88.515 114.680 88.815 ;
        RECT 115.065 88.545 115.530 88.875 ;
        RECT 113.850 88.485 114.050 88.515 ;
        RECT 114.170 88.265 114.340 88.335 ;
        RECT 113.470 88.095 114.340 88.265 ;
        RECT 113.830 88.005 114.340 88.095 ;
        RECT 112.380 87.540 112.685 87.670 ;
        RECT 113.130 87.560 113.660 87.925 ;
        RECT 112.000 86.945 112.265 87.405 ;
        RECT 112.435 87.115 112.685 87.540 ;
        RECT 113.830 87.390 114.000 88.005 ;
        RECT 112.895 87.220 114.000 87.390 ;
        RECT 114.170 86.945 114.340 87.745 ;
        RECT 114.510 87.445 114.680 88.515 ;
        RECT 114.850 87.615 115.040 88.335 ;
        RECT 115.210 87.585 115.530 88.545 ;
        RECT 115.700 88.585 115.870 89.045 ;
        RECT 116.145 88.965 116.355 89.495 ;
        RECT 116.615 88.755 116.945 89.280 ;
        RECT 117.115 88.885 117.285 89.495 ;
        RECT 117.455 88.840 117.785 89.275 ;
        RECT 117.455 88.755 117.835 88.840 ;
        RECT 116.745 88.585 116.945 88.755 ;
        RECT 117.610 88.715 117.835 88.755 ;
        RECT 115.700 88.255 116.575 88.585 ;
        RECT 116.745 88.255 117.495 88.585 ;
        RECT 114.510 87.115 114.760 87.445 ;
        RECT 115.700 87.415 115.870 88.255 ;
        RECT 116.745 88.050 116.935 88.255 ;
        RECT 117.665 88.135 117.835 88.715 ;
        RECT 117.620 88.085 117.835 88.135 ;
        RECT 116.040 87.675 116.935 88.050 ;
        RECT 117.445 88.005 117.835 88.085 ;
        RECT 118.040 88.755 118.655 89.325 ;
        RECT 118.825 88.985 119.040 89.495 ;
        RECT 119.270 88.985 119.550 89.315 ;
        RECT 119.730 88.985 119.970 89.495 ;
        RECT 114.985 87.245 115.870 87.415 ;
        RECT 116.050 86.945 116.365 87.445 ;
        RECT 116.595 87.115 116.935 87.675 ;
        RECT 117.105 86.945 117.275 87.955 ;
        RECT 117.445 87.160 117.775 88.005 ;
        RECT 118.040 87.735 118.355 88.755 ;
        RECT 118.525 88.085 118.695 88.585 ;
        RECT 118.945 88.255 119.210 88.815 ;
        RECT 119.380 88.085 119.550 88.985 ;
        RECT 119.720 88.255 120.075 88.815 ;
        RECT 120.305 88.695 120.615 89.495 ;
        RECT 120.820 88.695 121.515 89.325 ;
        RECT 121.685 88.725 125.195 89.495 ;
        RECT 125.825 88.770 126.115 89.495 ;
        RECT 126.745 89.115 127.635 89.285 ;
        RECT 120.315 88.255 120.650 88.525 ;
        RECT 120.820 88.095 120.990 88.695 ;
        RECT 121.160 88.255 121.495 88.505 ;
        RECT 121.685 88.205 123.335 88.725 ;
        RECT 126.745 88.560 127.295 88.945 ;
        RECT 118.525 87.915 119.950 88.085 ;
        RECT 118.040 87.115 118.575 87.735 ;
        RECT 118.745 86.945 119.075 87.745 ;
        RECT 119.560 87.740 119.950 87.915 ;
        RECT 120.305 86.945 120.585 88.085 ;
        RECT 120.755 87.115 121.085 88.095 ;
        RECT 121.255 86.945 121.515 88.085 ;
        RECT 123.505 88.035 125.195 88.555 ;
        RECT 127.465 88.390 127.635 89.115 ;
        RECT 126.745 88.320 127.635 88.390 ;
        RECT 127.805 88.815 128.025 89.275 ;
        RECT 128.195 88.955 128.445 89.495 ;
        RECT 128.615 88.845 128.875 89.325 ;
        RECT 129.045 88.950 134.390 89.495 ;
        RECT 135.035 89.135 137.105 89.325 ;
        RECT 137.335 89.135 137.665 89.495 ;
        RECT 138.195 89.135 138.525 89.495 ;
        RECT 139.055 89.135 139.385 89.495 ;
        RECT 135.985 89.115 137.105 89.135 ;
        RECT 127.805 88.790 128.055 88.815 ;
        RECT 127.805 88.365 128.135 88.790 ;
        RECT 126.745 88.295 127.640 88.320 ;
        RECT 126.745 88.280 127.650 88.295 ;
        RECT 126.745 88.265 127.655 88.280 ;
        RECT 126.745 88.260 127.665 88.265 ;
        RECT 126.745 88.250 127.670 88.260 ;
        RECT 126.745 88.240 127.675 88.250 ;
        RECT 126.745 88.235 127.685 88.240 ;
        RECT 126.745 88.225 127.695 88.235 ;
        RECT 126.745 88.220 127.705 88.225 ;
        RECT 121.685 86.945 125.195 88.035 ;
        RECT 125.825 86.945 126.115 88.110 ;
        RECT 126.745 87.770 127.005 88.220 ;
        RECT 127.370 88.215 127.705 88.220 ;
        RECT 127.370 88.210 127.720 88.215 ;
        RECT 127.370 88.200 127.735 88.210 ;
        RECT 127.370 88.195 127.760 88.200 ;
        RECT 128.305 88.195 128.535 88.590 ;
        RECT 127.370 88.190 128.535 88.195 ;
        RECT 127.400 88.155 128.535 88.190 ;
        RECT 127.435 88.130 128.535 88.155 ;
        RECT 127.465 88.100 128.535 88.130 ;
        RECT 127.485 88.070 128.535 88.100 ;
        RECT 127.505 88.040 128.535 88.070 ;
        RECT 127.575 88.030 128.535 88.040 ;
        RECT 127.600 88.020 128.535 88.030 ;
        RECT 127.620 88.005 128.535 88.020 ;
        RECT 127.640 87.990 128.535 88.005 ;
        RECT 127.645 87.980 128.430 87.990 ;
        RECT 127.660 87.945 128.430 87.980 ;
        RECT 127.175 87.625 127.505 87.870 ;
        RECT 127.675 87.695 128.430 87.945 ;
        RECT 128.705 87.815 128.875 88.845 ;
        RECT 130.630 88.120 130.970 88.950 ;
        RECT 127.175 87.600 127.360 87.625 ;
        RECT 126.745 87.500 127.360 87.600 ;
        RECT 126.745 86.945 127.350 87.500 ;
        RECT 127.525 87.115 128.005 87.455 ;
        RECT 128.175 86.945 128.430 87.490 ;
        RECT 128.600 87.115 128.875 87.815 ;
        RECT 132.450 87.380 132.800 88.630 ;
        RECT 135.025 87.610 135.315 88.585 ;
        RECT 135.485 88.040 135.815 88.910 ;
        RECT 135.985 88.690 136.175 89.115 ;
        RECT 138.695 88.945 138.885 89.065 ;
        RECT 136.345 88.735 138.885 88.945 ;
        RECT 139.055 88.505 139.395 88.815 ;
        RECT 140.145 88.675 140.355 89.495 ;
        RECT 140.525 88.695 140.855 89.325 ;
        RECT 135.985 88.215 136.845 88.505 ;
        RECT 137.305 88.225 138.275 88.505 ;
        RECT 138.445 88.335 139.395 88.505 ;
        RECT 138.500 88.285 139.395 88.335 ;
        RECT 140.525 88.095 140.775 88.695 ;
        RECT 141.025 88.675 141.255 89.495 ;
        RECT 141.925 88.695 142.265 89.325 ;
        RECT 142.435 88.695 142.685 89.495 ;
        RECT 142.875 88.845 143.205 89.325 ;
        RECT 143.375 89.035 143.600 89.495 ;
        RECT 143.770 88.845 144.100 89.325 ;
        RECT 140.945 88.255 141.275 88.505 ;
        RECT 141.925 88.135 142.100 88.695 ;
        RECT 142.875 88.675 144.100 88.845 ;
        RECT 144.730 88.715 145.230 89.325 ;
        RECT 145.655 88.955 145.880 89.315 ;
        RECT 146.060 89.125 146.390 89.495 ;
        RECT 146.570 88.955 146.825 89.315 ;
        RECT 147.390 89.125 148.135 89.495 ;
        RECT 145.655 88.765 148.140 88.955 ;
        RECT 142.270 88.335 142.965 88.505 ;
        RECT 135.485 87.870 138.095 88.040 ;
        RECT 129.045 86.945 134.390 87.380 ;
        RECT 135.055 86.945 135.315 87.405 ;
        RECT 135.485 87.115 135.745 87.870 ;
        RECT 135.915 86.945 136.245 87.665 ;
        RECT 136.415 87.115 136.605 87.870 ;
        RECT 136.775 86.945 137.105 87.665 ;
        RECT 137.335 87.285 137.595 87.480 ;
        RECT 137.765 87.455 138.095 87.870 ;
        RECT 138.265 87.885 139.385 88.055 ;
        RECT 138.265 87.285 138.455 87.885 ;
        RECT 137.335 87.115 138.455 87.285 ;
        RECT 138.625 86.945 138.955 87.715 ;
        RECT 139.125 87.115 139.385 87.885 ;
        RECT 140.145 86.945 140.355 88.085 ;
        RECT 140.525 87.115 140.855 88.095 ;
        RECT 141.925 88.085 142.155 88.135 ;
        RECT 142.795 88.085 142.965 88.335 ;
        RECT 143.140 88.305 143.560 88.505 ;
        RECT 143.730 88.305 144.060 88.505 ;
        RECT 144.230 88.305 144.560 88.505 ;
        RECT 144.730 88.085 144.900 88.715 ;
        RECT 145.085 88.255 145.435 88.505 ;
        RECT 145.615 88.255 145.885 88.585 ;
        RECT 146.065 88.255 146.500 88.585 ;
        RECT 146.680 88.255 147.255 88.585 ;
        RECT 147.435 88.255 147.715 88.585 ;
        RECT 141.025 86.945 141.255 88.085 ;
        RECT 141.925 87.115 142.265 88.085 ;
        RECT 142.435 86.945 142.605 88.085 ;
        RECT 142.795 87.915 145.230 88.085 ;
        RECT 147.915 88.075 148.140 88.765 ;
        RECT 142.875 86.945 143.125 87.745 ;
        RECT 143.770 87.115 144.100 87.915 ;
        RECT 144.400 86.945 144.730 87.745 ;
        RECT 144.900 87.115 145.230 87.915 ;
        RECT 145.645 87.895 148.140 88.075 ;
        RECT 148.315 87.895 148.650 89.315 ;
        RECT 148.990 88.985 149.230 89.495 ;
        RECT 149.410 88.985 149.690 89.315 ;
        RECT 149.920 88.985 150.135 89.495 ;
        RECT 148.885 88.255 149.240 88.815 ;
        RECT 149.410 88.085 149.580 88.985 ;
        RECT 149.750 88.255 150.015 88.815 ;
        RECT 150.305 88.755 150.920 89.325 ;
        RECT 151.585 88.770 151.875 89.495 ;
        RECT 152.210 88.985 152.450 89.495 ;
        RECT 152.630 88.985 152.910 89.315 ;
        RECT 153.140 88.985 153.355 89.495 ;
        RECT 150.265 88.085 150.435 88.585 ;
        RECT 145.645 87.125 145.935 87.895 ;
        RECT 146.505 87.485 147.695 87.715 ;
        RECT 146.505 87.125 146.765 87.485 ;
        RECT 146.935 86.945 147.265 87.315 ;
        RECT 147.435 87.125 147.695 87.485 ;
        RECT 147.885 86.945 148.215 87.665 ;
        RECT 148.385 87.125 148.650 87.895 ;
        RECT 149.010 87.915 150.435 88.085 ;
        RECT 149.010 87.740 149.400 87.915 ;
        RECT 149.885 86.945 150.215 87.745 ;
        RECT 150.605 87.735 150.920 88.755 ;
        RECT 152.105 88.255 152.460 88.815 ;
        RECT 150.385 87.115 150.920 87.735 ;
        RECT 151.585 86.945 151.875 88.110 ;
        RECT 152.630 88.085 152.800 88.985 ;
        RECT 152.970 88.255 153.235 88.815 ;
        RECT 153.525 88.755 154.140 89.325 ;
        RECT 153.485 88.085 153.655 88.585 ;
        RECT 152.230 87.915 153.655 88.085 ;
        RECT 152.230 87.740 152.620 87.915 ;
        RECT 153.105 86.945 153.435 87.745 ;
        RECT 153.825 87.735 154.140 88.755 ;
        RECT 154.345 88.745 155.555 89.495 ;
        RECT 155.725 88.745 156.935 89.495 ;
        RECT 154.345 88.205 154.865 88.745 ;
        RECT 155.035 88.035 155.555 88.575 ;
        RECT 153.605 87.115 154.140 87.735 ;
        RECT 154.345 86.945 155.555 88.035 ;
        RECT 155.725 88.035 156.245 88.575 ;
        RECT 156.415 88.205 156.935 88.745 ;
        RECT 155.725 86.945 156.935 88.035 ;
        RECT 22.700 86.775 157.020 86.945 ;
        RECT 22.785 85.685 23.995 86.775 ;
        RECT 24.165 86.340 29.510 86.775 ;
        RECT 22.785 84.975 23.305 85.515 ;
        RECT 23.475 85.145 23.995 85.685 ;
        RECT 22.785 84.225 23.995 84.975 ;
        RECT 25.750 84.770 26.090 85.600 ;
        RECT 27.570 85.090 27.920 86.340 ;
        RECT 29.685 85.685 33.195 86.775 ;
        RECT 29.685 84.995 31.335 85.515 ;
        RECT 31.505 85.165 33.195 85.685 ;
        RECT 34.285 85.635 34.545 86.775 ;
        RECT 34.715 85.625 35.045 86.605 ;
        RECT 35.215 85.635 35.495 86.775 ;
        RECT 34.305 85.215 34.640 85.465 ;
        RECT 34.810 85.025 34.980 85.625 ;
        RECT 35.665 85.610 35.955 86.775 ;
        RECT 36.310 85.805 36.700 85.980 ;
        RECT 37.185 85.975 37.515 86.775 ;
        RECT 37.685 85.985 38.220 86.605 ;
        RECT 36.310 85.635 37.735 85.805 ;
        RECT 35.150 85.195 35.485 85.465 ;
        RECT 24.165 84.225 29.510 84.770 ;
        RECT 29.685 84.225 33.195 84.995 ;
        RECT 34.285 84.395 34.980 85.025 ;
        RECT 35.185 84.225 35.495 85.025 ;
        RECT 35.665 84.225 35.955 84.950 ;
        RECT 36.185 84.905 36.540 85.465 ;
        RECT 36.710 84.735 36.880 85.635 ;
        RECT 37.050 84.905 37.315 85.465 ;
        RECT 37.565 85.135 37.735 85.635 ;
        RECT 37.905 84.965 38.220 85.985 ;
        RECT 36.290 84.225 36.530 84.735 ;
        RECT 36.710 84.405 36.990 84.735 ;
        RECT 37.220 84.225 37.435 84.735 ;
        RECT 37.605 84.395 38.220 84.965 ;
        RECT 38.425 85.905 38.700 86.605 ;
        RECT 38.870 86.230 39.125 86.775 ;
        RECT 39.295 86.265 39.775 86.605 ;
        RECT 39.950 86.220 40.555 86.775 ;
        RECT 39.940 86.120 40.555 86.220 ;
        RECT 39.940 86.095 40.125 86.120 ;
        RECT 38.425 84.875 38.595 85.905 ;
        RECT 38.870 85.775 39.625 86.025 ;
        RECT 39.795 85.850 40.125 86.095 ;
        RECT 40.915 86.050 41.245 86.775 ;
        RECT 38.870 85.740 39.640 85.775 ;
        RECT 38.870 85.730 39.655 85.740 ;
        RECT 38.765 85.715 39.660 85.730 ;
        RECT 38.765 85.700 39.680 85.715 ;
        RECT 38.765 85.690 39.700 85.700 ;
        RECT 38.765 85.680 39.725 85.690 ;
        RECT 38.765 85.650 39.795 85.680 ;
        RECT 38.765 85.620 39.815 85.650 ;
        RECT 38.765 85.590 39.835 85.620 ;
        RECT 38.765 85.565 39.865 85.590 ;
        RECT 38.765 85.530 39.900 85.565 ;
        RECT 38.765 85.525 39.930 85.530 ;
        RECT 38.765 85.130 38.995 85.525 ;
        RECT 39.540 85.520 39.930 85.525 ;
        RECT 39.565 85.510 39.930 85.520 ;
        RECT 39.580 85.505 39.930 85.510 ;
        RECT 39.595 85.500 39.930 85.505 ;
        RECT 40.295 85.500 40.555 85.950 ;
        RECT 39.595 85.495 40.555 85.500 ;
        RECT 39.605 85.485 40.555 85.495 ;
        RECT 39.615 85.480 40.555 85.485 ;
        RECT 39.625 85.470 40.555 85.480 ;
        RECT 39.630 85.460 40.555 85.470 ;
        RECT 39.635 85.455 40.555 85.460 ;
        RECT 39.645 85.440 40.555 85.455 ;
        RECT 39.650 85.425 40.555 85.440 ;
        RECT 39.660 85.400 40.555 85.425 ;
        RECT 39.165 84.930 39.495 85.355 ;
        RECT 39.245 84.905 39.495 84.930 ;
        RECT 38.425 84.395 38.685 84.875 ;
        RECT 38.855 84.225 39.105 84.765 ;
        RECT 39.275 84.445 39.495 84.905 ;
        RECT 39.665 85.330 40.555 85.400 ;
        RECT 39.665 84.605 39.835 85.330 ;
        RECT 40.005 84.775 40.555 85.160 ;
        RECT 39.665 84.435 40.555 84.605 ;
        RECT 40.725 84.395 41.245 85.880 ;
        RECT 41.415 85.055 41.935 86.605 ;
        RECT 43.025 85.635 43.285 86.775 ;
        RECT 43.455 85.625 43.785 86.605 ;
        RECT 43.955 85.635 44.235 86.775 ;
        RECT 43.045 85.215 43.380 85.465 ;
        RECT 43.550 85.025 43.720 85.625 ;
        RECT 43.890 85.195 44.225 85.465 ;
        RECT 44.405 85.055 44.925 86.605 ;
        RECT 45.095 86.050 45.425 86.775 ;
        RECT 41.415 84.225 41.755 84.885 ;
        RECT 43.025 84.395 43.720 85.025 ;
        RECT 43.925 84.225 44.235 85.025 ;
        RECT 44.585 84.225 44.925 84.885 ;
        RECT 45.095 84.395 45.615 85.880 ;
        RECT 45.785 85.685 49.295 86.775 ;
        RECT 45.785 84.995 47.435 85.515 ;
        RECT 47.605 85.165 49.295 85.685 ;
        RECT 49.465 85.635 49.725 86.775 ;
        RECT 49.895 85.625 50.225 86.605 ;
        RECT 50.395 85.635 50.675 86.775 ;
        RECT 49.485 85.215 49.820 85.465 ;
        RECT 49.990 85.025 50.160 85.625 ;
        RECT 50.330 85.195 50.665 85.465 ;
        RECT 51.765 85.055 52.285 86.605 ;
        RECT 52.455 86.050 52.785 86.775 ;
        RECT 45.785 84.225 49.295 84.995 ;
        RECT 49.465 84.395 50.160 85.025 ;
        RECT 50.365 84.225 50.675 85.025 ;
        RECT 51.945 84.225 52.285 84.885 ;
        RECT 52.455 84.395 52.975 85.880 ;
        RECT 53.145 85.685 54.815 86.775 ;
        RECT 53.145 84.995 53.895 85.515 ;
        RECT 54.065 85.165 54.815 85.685 ;
        RECT 55.630 85.805 56.020 85.980 ;
        RECT 56.505 85.975 56.835 86.775 ;
        RECT 57.005 85.985 57.540 86.605 ;
        RECT 57.745 86.220 58.350 86.775 ;
        RECT 58.525 86.265 59.005 86.605 ;
        RECT 59.175 86.230 59.430 86.775 ;
        RECT 57.745 86.120 58.360 86.220 ;
        RECT 55.630 85.635 57.055 85.805 ;
        RECT 53.145 84.225 54.815 84.995 ;
        RECT 55.505 84.905 55.860 85.465 ;
        RECT 56.030 84.735 56.200 85.635 ;
        RECT 56.370 84.905 56.635 85.465 ;
        RECT 56.885 85.135 57.055 85.635 ;
        RECT 57.225 84.965 57.540 85.985 ;
        RECT 58.175 86.095 58.360 86.120 ;
        RECT 57.745 85.500 58.005 85.950 ;
        RECT 58.175 85.850 58.505 86.095 ;
        RECT 58.675 85.775 59.430 86.025 ;
        RECT 59.600 85.905 59.875 86.605 ;
        RECT 58.660 85.740 59.430 85.775 ;
        RECT 58.645 85.730 59.430 85.740 ;
        RECT 58.640 85.715 59.535 85.730 ;
        RECT 58.620 85.700 59.535 85.715 ;
        RECT 58.600 85.690 59.535 85.700 ;
        RECT 58.575 85.680 59.535 85.690 ;
        RECT 58.505 85.650 59.535 85.680 ;
        RECT 58.485 85.620 59.535 85.650 ;
        RECT 58.465 85.590 59.535 85.620 ;
        RECT 58.435 85.565 59.535 85.590 ;
        RECT 58.400 85.530 59.535 85.565 ;
        RECT 58.370 85.525 59.535 85.530 ;
        RECT 58.370 85.520 58.760 85.525 ;
        RECT 58.370 85.510 58.735 85.520 ;
        RECT 58.370 85.505 58.720 85.510 ;
        RECT 58.370 85.500 58.705 85.505 ;
        RECT 57.745 85.495 58.705 85.500 ;
        RECT 57.745 85.485 58.695 85.495 ;
        RECT 57.745 85.480 58.685 85.485 ;
        RECT 57.745 85.470 58.675 85.480 ;
        RECT 57.745 85.460 58.670 85.470 ;
        RECT 57.745 85.455 58.665 85.460 ;
        RECT 57.745 85.440 58.655 85.455 ;
        RECT 57.745 85.425 58.650 85.440 ;
        RECT 57.745 85.400 58.640 85.425 ;
        RECT 57.745 85.330 58.635 85.400 ;
        RECT 55.610 84.225 55.850 84.735 ;
        RECT 56.030 84.405 56.310 84.735 ;
        RECT 56.540 84.225 56.755 84.735 ;
        RECT 56.925 84.395 57.540 84.965 ;
        RECT 57.745 84.775 58.295 85.160 ;
        RECT 58.465 84.605 58.635 85.330 ;
        RECT 57.745 84.435 58.635 84.605 ;
        RECT 58.805 84.930 59.135 85.355 ;
        RECT 59.305 85.130 59.535 85.525 ;
        RECT 58.805 84.445 59.025 84.930 ;
        RECT 59.705 84.875 59.875 85.905 ;
        RECT 60.045 85.685 61.255 86.775 ;
        RECT 59.195 84.225 59.445 84.765 ;
        RECT 59.615 84.395 59.875 84.875 ;
        RECT 60.045 84.975 60.565 85.515 ;
        RECT 60.735 85.145 61.255 85.685 ;
        RECT 61.425 85.610 61.715 86.775 ;
        RECT 61.885 85.685 64.475 86.775 ;
        RECT 64.645 86.220 65.250 86.775 ;
        RECT 65.425 86.265 65.905 86.605 ;
        RECT 66.075 86.230 66.330 86.775 ;
        RECT 64.645 86.120 65.260 86.220 ;
        RECT 65.075 86.095 65.260 86.120 ;
        RECT 61.885 84.995 63.095 85.515 ;
        RECT 63.265 85.165 64.475 85.685 ;
        RECT 64.645 85.500 64.905 85.950 ;
        RECT 65.075 85.850 65.405 86.095 ;
        RECT 65.575 85.775 66.330 86.025 ;
        RECT 66.500 85.905 66.775 86.605 ;
        RECT 65.560 85.740 66.330 85.775 ;
        RECT 65.545 85.730 66.330 85.740 ;
        RECT 65.540 85.715 66.435 85.730 ;
        RECT 65.520 85.700 66.435 85.715 ;
        RECT 65.500 85.690 66.435 85.700 ;
        RECT 65.475 85.680 66.435 85.690 ;
        RECT 65.405 85.650 66.435 85.680 ;
        RECT 65.385 85.620 66.435 85.650 ;
        RECT 65.365 85.590 66.435 85.620 ;
        RECT 65.335 85.565 66.435 85.590 ;
        RECT 65.300 85.530 66.435 85.565 ;
        RECT 65.270 85.525 66.435 85.530 ;
        RECT 65.270 85.520 65.660 85.525 ;
        RECT 65.270 85.510 65.635 85.520 ;
        RECT 65.270 85.505 65.620 85.510 ;
        RECT 65.270 85.500 65.605 85.505 ;
        RECT 64.645 85.495 65.605 85.500 ;
        RECT 64.645 85.485 65.595 85.495 ;
        RECT 64.645 85.480 65.585 85.485 ;
        RECT 64.645 85.470 65.575 85.480 ;
        RECT 64.645 85.460 65.570 85.470 ;
        RECT 64.645 85.455 65.565 85.460 ;
        RECT 64.645 85.440 65.555 85.455 ;
        RECT 64.645 85.425 65.550 85.440 ;
        RECT 64.645 85.400 65.540 85.425 ;
        RECT 64.645 85.330 65.535 85.400 ;
        RECT 60.045 84.225 61.255 84.975 ;
        RECT 61.425 84.225 61.715 84.950 ;
        RECT 61.885 84.225 64.475 84.995 ;
        RECT 64.645 84.775 65.195 85.160 ;
        RECT 65.365 84.605 65.535 85.330 ;
        RECT 64.645 84.435 65.535 84.605 ;
        RECT 65.705 84.930 66.035 85.355 ;
        RECT 66.205 85.130 66.435 85.525 ;
        RECT 65.705 84.905 65.955 84.930 ;
        RECT 65.705 84.445 65.925 84.905 ;
        RECT 66.605 84.875 66.775 85.905 ;
        RECT 66.095 84.225 66.345 84.765 ;
        RECT 66.515 84.395 66.775 84.875 ;
        RECT 66.950 85.825 67.215 86.595 ;
        RECT 67.385 86.055 67.715 86.775 ;
        RECT 67.905 86.235 68.165 86.595 ;
        RECT 68.335 86.405 68.665 86.775 ;
        RECT 68.835 86.235 69.095 86.595 ;
        RECT 67.905 86.005 69.095 86.235 ;
        RECT 69.665 85.825 69.955 86.595 ;
        RECT 70.195 86.315 70.455 86.775 ;
        RECT 66.950 84.405 67.285 85.825 ;
        RECT 67.460 85.645 69.955 85.825 ;
        RECT 67.460 84.955 67.685 85.645 ;
        RECT 67.885 85.135 68.165 85.465 ;
        RECT 68.345 85.135 68.920 85.465 ;
        RECT 69.100 85.135 69.535 85.465 ;
        RECT 69.715 85.135 69.985 85.465 ;
        RECT 70.165 85.135 70.455 86.110 ;
        RECT 70.625 85.850 70.885 86.605 ;
        RECT 71.055 86.055 71.385 86.775 ;
        RECT 71.555 85.850 71.745 86.605 ;
        RECT 71.915 86.055 72.245 86.775 ;
        RECT 72.475 86.435 73.595 86.605 ;
        RECT 72.475 86.240 72.735 86.435 ;
        RECT 72.905 85.850 73.235 86.265 ;
        RECT 70.625 85.680 73.235 85.850 ;
        RECT 73.405 85.835 73.595 86.435 ;
        RECT 73.765 86.005 74.095 86.775 ;
        RECT 74.265 85.835 74.525 86.605 ;
        RECT 67.460 84.765 69.945 84.955 ;
        RECT 70.625 84.810 70.955 85.680 ;
        RECT 73.405 85.665 74.525 85.835 ;
        RECT 74.765 85.685 77.355 86.775 ;
        RECT 71.125 85.215 71.985 85.505 ;
        RECT 72.445 85.215 73.415 85.495 ;
        RECT 73.640 85.385 74.535 85.435 ;
        RECT 73.585 85.215 74.535 85.385 ;
        RECT 67.465 84.225 68.210 84.595 ;
        RECT 68.775 84.405 69.030 84.765 ;
        RECT 69.210 84.225 69.540 84.595 ;
        RECT 69.720 84.405 69.945 84.765 ;
        RECT 71.125 84.605 71.315 85.030 ;
        RECT 71.485 84.775 74.025 84.985 ;
        RECT 74.195 84.905 74.535 85.215 ;
        RECT 74.765 84.995 75.975 85.515 ;
        RECT 76.145 85.165 77.355 85.685 ;
        RECT 77.525 86.055 77.985 86.605 ;
        RECT 78.175 86.055 78.505 86.775 ;
        RECT 73.835 84.655 74.025 84.775 ;
        RECT 71.125 84.585 72.245 84.605 ;
        RECT 70.175 84.395 72.245 84.585 ;
        RECT 72.475 84.225 72.805 84.585 ;
        RECT 73.335 84.225 73.665 84.585 ;
        RECT 74.195 84.225 74.525 84.585 ;
        RECT 74.765 84.225 77.355 84.995 ;
        RECT 77.525 84.685 77.775 86.055 ;
        RECT 78.705 85.885 79.005 86.435 ;
        RECT 79.175 86.105 79.455 86.775 ;
        RECT 78.065 85.715 79.005 85.885 ;
        RECT 79.835 85.825 80.110 86.595 ;
        RECT 80.280 86.165 80.610 86.595 ;
        RECT 80.780 86.335 80.975 86.775 ;
        RECT 81.155 86.165 81.485 86.595 ;
        RECT 80.280 85.995 81.485 86.165 ;
        RECT 78.065 85.465 78.235 85.715 ;
        RECT 79.375 85.465 79.640 85.825 ;
        RECT 79.835 85.635 80.420 85.825 ;
        RECT 80.590 85.665 81.485 85.995 ;
        RECT 81.675 85.635 82.005 86.775 ;
        RECT 82.535 85.805 82.865 86.590 ;
        RECT 82.185 85.635 82.865 85.805 ;
        RECT 83.045 85.685 85.635 86.775 ;
        RECT 77.945 85.135 78.235 85.465 ;
        RECT 78.405 85.215 78.745 85.465 ;
        RECT 78.965 85.215 79.640 85.465 ;
        RECT 78.065 85.045 78.235 85.135 ;
        RECT 78.065 84.855 79.455 85.045 ;
        RECT 77.525 84.395 78.085 84.685 ;
        RECT 78.255 84.225 78.505 84.685 ;
        RECT 79.125 84.495 79.455 84.855 ;
        RECT 79.835 84.815 80.075 85.465 ;
        RECT 80.245 84.965 80.420 85.635 ;
        RECT 80.590 85.135 81.005 85.465 ;
        RECT 81.185 85.135 81.480 85.465 ;
        RECT 81.665 85.215 82.015 85.465 ;
        RECT 80.245 84.785 80.575 84.965 ;
        RECT 79.850 84.225 80.180 84.615 ;
        RECT 80.350 84.405 80.575 84.785 ;
        RECT 80.775 84.515 81.005 85.135 ;
        RECT 82.185 85.035 82.355 85.635 ;
        RECT 82.525 85.215 82.875 85.465 ;
        RECT 81.185 84.225 81.485 84.955 ;
        RECT 81.675 84.225 81.945 85.035 ;
        RECT 82.115 84.395 82.445 85.035 ;
        RECT 82.615 84.225 82.855 85.035 ;
        RECT 83.045 84.995 84.255 85.515 ;
        RECT 84.425 85.165 85.635 85.685 ;
        RECT 85.805 85.635 86.065 86.775 ;
        RECT 86.235 85.625 86.565 86.605 ;
        RECT 86.735 85.635 87.015 86.775 ;
        RECT 85.825 85.215 86.160 85.465 ;
        RECT 86.330 85.025 86.500 85.625 ;
        RECT 87.185 85.610 87.475 86.775 ;
        RECT 87.705 85.715 88.035 86.560 ;
        RECT 88.205 85.765 88.375 86.775 ;
        RECT 88.545 86.045 88.885 86.605 ;
        RECT 89.115 86.275 89.430 86.775 ;
        RECT 89.610 86.305 90.495 86.475 ;
        RECT 87.645 85.635 88.035 85.715 ;
        RECT 88.545 85.670 89.440 86.045 ;
        RECT 87.645 85.585 87.860 85.635 ;
        RECT 86.670 85.195 87.005 85.465 ;
        RECT 83.045 84.225 85.635 84.995 ;
        RECT 85.805 84.395 86.500 85.025 ;
        RECT 86.705 84.225 87.015 85.025 ;
        RECT 87.645 85.005 87.815 85.585 ;
        RECT 88.545 85.465 88.735 85.670 ;
        RECT 89.610 85.465 89.780 86.305 ;
        RECT 90.720 86.275 90.970 86.605 ;
        RECT 87.985 85.135 88.735 85.465 ;
        RECT 88.905 85.135 89.780 85.465 ;
        RECT 87.645 84.965 87.870 85.005 ;
        RECT 88.535 84.965 88.735 85.135 ;
        RECT 87.185 84.225 87.475 84.950 ;
        RECT 87.645 84.880 88.025 84.965 ;
        RECT 87.695 84.445 88.025 84.880 ;
        RECT 88.195 84.225 88.365 84.835 ;
        RECT 88.535 84.440 88.865 84.965 ;
        RECT 89.125 84.225 89.335 84.755 ;
        RECT 89.610 84.675 89.780 85.135 ;
        RECT 89.950 85.175 90.270 86.135 ;
        RECT 90.440 85.385 90.630 86.105 ;
        RECT 90.800 85.205 90.970 86.275 ;
        RECT 91.140 85.975 91.310 86.775 ;
        RECT 91.480 86.330 92.585 86.500 ;
        RECT 91.480 85.715 91.650 86.330 ;
        RECT 92.795 86.180 93.045 86.605 ;
        RECT 93.215 86.315 93.480 86.775 ;
        RECT 91.820 85.795 92.350 86.160 ;
        RECT 92.795 86.050 93.100 86.180 ;
        RECT 91.140 85.625 91.650 85.715 ;
        RECT 91.140 85.455 92.010 85.625 ;
        RECT 91.140 85.385 91.310 85.455 ;
        RECT 91.430 85.205 91.630 85.235 ;
        RECT 89.950 84.845 90.415 85.175 ;
        RECT 90.800 84.905 91.630 85.205 ;
        RECT 90.800 84.675 90.970 84.905 ;
        RECT 89.610 84.505 90.395 84.675 ;
        RECT 90.565 84.505 90.970 84.675 ;
        RECT 91.150 84.225 91.520 84.725 ;
        RECT 91.840 84.675 92.010 85.455 ;
        RECT 92.180 85.095 92.350 85.795 ;
        RECT 92.520 85.265 92.760 85.860 ;
        RECT 92.180 84.875 92.705 85.095 ;
        RECT 92.930 84.945 93.100 86.050 ;
        RECT 92.875 84.815 93.100 84.945 ;
        RECT 93.270 84.855 93.550 85.805 ;
        RECT 92.875 84.675 93.045 84.815 ;
        RECT 91.840 84.505 92.515 84.675 ;
        RECT 92.710 84.505 93.045 84.675 ;
        RECT 93.215 84.225 93.465 84.685 ;
        RECT 93.720 84.485 93.905 86.605 ;
        RECT 94.075 86.275 94.405 86.775 ;
        RECT 94.575 86.105 94.745 86.605 ;
        RECT 94.080 85.935 94.745 86.105 ;
        RECT 95.500 85.985 96.035 86.605 ;
        RECT 94.080 84.945 94.310 85.935 ;
        RECT 94.480 85.115 94.830 85.765 ;
        RECT 95.500 84.965 95.815 85.985 ;
        RECT 96.205 85.975 96.535 86.775 ;
        RECT 97.020 85.805 97.410 85.980 ;
        RECT 95.985 85.635 97.410 85.805 ;
        RECT 97.765 85.635 98.025 86.775 ;
        RECT 95.985 85.135 96.155 85.635 ;
        RECT 94.080 84.775 94.745 84.945 ;
        RECT 94.075 84.225 94.405 84.605 ;
        RECT 94.575 84.485 94.745 84.775 ;
        RECT 95.500 84.395 96.115 84.965 ;
        RECT 96.405 84.905 96.670 85.465 ;
        RECT 96.840 84.735 97.010 85.635 ;
        RECT 98.195 85.625 98.525 86.605 ;
        RECT 98.695 85.635 98.975 86.775 ;
        RECT 100.065 85.905 100.340 86.605 ;
        RECT 100.550 86.230 100.765 86.775 ;
        RECT 100.935 86.265 101.410 86.605 ;
        RECT 101.580 86.270 102.195 86.775 ;
        RECT 101.580 86.095 101.775 86.270 ;
        RECT 97.180 84.905 97.535 85.465 ;
        RECT 97.785 85.215 98.120 85.465 ;
        RECT 98.290 85.025 98.460 85.625 ;
        RECT 98.630 85.195 98.965 85.465 ;
        RECT 96.285 84.225 96.500 84.735 ;
        RECT 96.730 84.405 97.010 84.735 ;
        RECT 97.190 84.225 97.430 84.735 ;
        RECT 97.765 84.395 98.460 85.025 ;
        RECT 98.665 84.225 98.975 85.025 ;
        RECT 100.065 84.875 100.235 85.905 ;
        RECT 100.510 85.735 101.225 86.030 ;
        RECT 101.445 85.905 101.775 86.095 ;
        RECT 101.945 85.735 102.195 86.100 ;
        RECT 100.405 85.565 102.195 85.735 ;
        RECT 100.405 85.135 100.635 85.565 ;
        RECT 100.065 84.395 100.325 84.875 ;
        RECT 100.805 84.865 101.215 85.385 ;
        RECT 100.495 84.225 100.825 84.685 ;
        RECT 101.015 84.445 101.215 84.865 ;
        RECT 101.385 84.710 101.640 85.565 ;
        RECT 102.435 85.385 102.605 86.605 ;
        RECT 102.855 86.265 103.115 86.775 ;
        RECT 101.810 85.135 102.605 85.385 ;
        RECT 102.775 85.215 103.115 86.095 ;
        RECT 103.285 85.685 105.875 86.775 ;
        RECT 102.355 85.045 102.605 85.135 ;
        RECT 101.385 84.445 102.175 84.710 ;
        RECT 102.355 84.625 102.685 85.045 ;
        RECT 102.855 84.225 103.115 85.045 ;
        RECT 103.285 84.995 104.495 85.515 ;
        RECT 104.665 85.165 105.875 85.685 ;
        RECT 106.045 85.635 106.305 86.775 ;
        RECT 106.475 85.625 106.805 86.605 ;
        RECT 106.975 85.635 107.255 86.775 ;
        RECT 107.425 86.340 112.770 86.775 ;
        RECT 106.065 85.215 106.400 85.465 ;
        RECT 106.570 85.025 106.740 85.625 ;
        RECT 106.910 85.195 107.245 85.465 ;
        RECT 103.285 84.225 105.875 84.995 ;
        RECT 106.045 84.395 106.740 85.025 ;
        RECT 106.945 84.225 107.255 85.025 ;
        RECT 109.010 84.770 109.350 85.600 ;
        RECT 110.830 85.090 111.180 86.340 ;
        RECT 112.945 85.610 113.235 86.775 ;
        RECT 113.405 86.340 118.750 86.775 ;
        RECT 118.925 86.340 124.270 86.775 ;
        RECT 107.425 84.225 112.770 84.770 ;
        RECT 112.945 84.225 113.235 84.950 ;
        RECT 114.990 84.770 115.330 85.600 ;
        RECT 116.810 85.090 117.160 86.340 ;
        RECT 120.510 84.770 120.850 85.600 ;
        RECT 122.330 85.090 122.680 86.340 ;
        RECT 124.445 85.685 127.035 86.775 ;
        RECT 124.445 84.995 125.655 85.515 ;
        RECT 125.825 85.165 127.035 85.685 ;
        RECT 127.295 85.845 127.465 86.605 ;
        RECT 127.645 86.015 127.975 86.775 ;
        RECT 127.295 85.675 127.960 85.845 ;
        RECT 128.145 85.700 128.415 86.605 ;
        RECT 128.675 86.105 128.845 86.605 ;
        RECT 129.015 86.275 129.345 86.775 ;
        RECT 128.675 85.935 129.340 86.105 ;
        RECT 127.790 85.530 127.960 85.675 ;
        RECT 127.225 85.125 127.555 85.495 ;
        RECT 127.790 85.200 128.075 85.530 ;
        RECT 113.405 84.225 118.750 84.770 ;
        RECT 118.925 84.225 124.270 84.770 ;
        RECT 124.445 84.225 127.035 84.995 ;
        RECT 127.790 84.945 127.960 85.200 ;
        RECT 127.295 84.775 127.960 84.945 ;
        RECT 128.245 84.900 128.415 85.700 ;
        RECT 128.590 85.115 128.940 85.765 ;
        RECT 129.110 84.945 129.340 85.935 ;
        RECT 127.295 84.395 127.465 84.775 ;
        RECT 127.645 84.225 127.975 84.605 ;
        RECT 128.155 84.395 128.415 84.900 ;
        RECT 128.675 84.775 129.340 84.945 ;
        RECT 128.675 84.485 128.845 84.775 ;
        RECT 129.015 84.225 129.345 84.605 ;
        RECT 129.515 84.485 129.700 86.605 ;
        RECT 129.940 86.315 130.205 86.775 ;
        RECT 130.375 86.180 130.625 86.605 ;
        RECT 130.835 86.330 131.940 86.500 ;
        RECT 130.320 86.050 130.625 86.180 ;
        RECT 129.870 84.855 130.150 85.805 ;
        RECT 130.320 84.945 130.490 86.050 ;
        RECT 130.660 85.265 130.900 85.860 ;
        RECT 131.070 85.795 131.600 86.160 ;
        RECT 131.070 85.095 131.240 85.795 ;
        RECT 131.770 85.715 131.940 86.330 ;
        RECT 132.110 85.975 132.280 86.775 ;
        RECT 132.450 86.275 132.700 86.605 ;
        RECT 132.925 86.305 133.810 86.475 ;
        RECT 131.770 85.625 132.280 85.715 ;
        RECT 130.320 84.815 130.545 84.945 ;
        RECT 130.715 84.875 131.240 85.095 ;
        RECT 131.410 85.455 132.280 85.625 ;
        RECT 129.955 84.225 130.205 84.685 ;
        RECT 130.375 84.675 130.545 84.815 ;
        RECT 131.410 84.675 131.580 85.455 ;
        RECT 132.110 85.385 132.280 85.455 ;
        RECT 131.790 85.205 131.990 85.235 ;
        RECT 132.450 85.205 132.620 86.275 ;
        RECT 132.790 85.385 132.980 86.105 ;
        RECT 131.790 84.905 132.620 85.205 ;
        RECT 133.150 85.175 133.470 86.135 ;
        RECT 130.375 84.505 130.710 84.675 ;
        RECT 130.905 84.505 131.580 84.675 ;
        RECT 131.900 84.225 132.270 84.725 ;
        RECT 132.450 84.675 132.620 84.905 ;
        RECT 133.005 84.845 133.470 85.175 ;
        RECT 133.640 85.465 133.810 86.305 ;
        RECT 133.990 86.275 134.305 86.775 ;
        RECT 134.535 86.045 134.875 86.605 ;
        RECT 133.980 85.670 134.875 86.045 ;
        RECT 135.045 85.765 135.215 86.775 ;
        RECT 134.685 85.465 134.875 85.670 ;
        RECT 135.385 85.715 135.715 86.560 ;
        RECT 136.130 85.805 136.520 85.980 ;
        RECT 137.005 85.975 137.335 86.775 ;
        RECT 137.505 85.985 138.040 86.605 ;
        RECT 135.385 85.635 135.775 85.715 ;
        RECT 136.130 85.635 137.555 85.805 ;
        RECT 135.560 85.585 135.775 85.635 ;
        RECT 133.640 85.135 134.515 85.465 ;
        RECT 134.685 85.135 135.435 85.465 ;
        RECT 133.640 84.675 133.810 85.135 ;
        RECT 134.685 84.965 134.885 85.135 ;
        RECT 135.605 85.005 135.775 85.585 ;
        RECT 135.550 84.965 135.775 85.005 ;
        RECT 132.450 84.505 132.855 84.675 ;
        RECT 133.025 84.505 133.810 84.675 ;
        RECT 134.085 84.225 134.295 84.755 ;
        RECT 134.555 84.440 134.885 84.965 ;
        RECT 135.395 84.880 135.775 84.965 ;
        RECT 136.005 84.905 136.360 85.465 ;
        RECT 135.055 84.225 135.225 84.835 ;
        RECT 135.395 84.445 135.725 84.880 ;
        RECT 136.530 84.735 136.700 85.635 ;
        RECT 136.870 84.905 137.135 85.465 ;
        RECT 137.385 85.135 137.555 85.635 ;
        RECT 137.725 84.965 138.040 85.985 ;
        RECT 138.705 85.610 138.995 86.775 ;
        RECT 140.085 86.265 140.345 86.775 ;
        RECT 140.085 85.215 140.425 86.095 ;
        RECT 140.595 85.385 140.765 86.605 ;
        RECT 141.005 86.270 141.620 86.775 ;
        RECT 141.005 85.735 141.255 86.100 ;
        RECT 141.425 86.095 141.620 86.270 ;
        RECT 141.790 86.265 142.265 86.605 ;
        RECT 142.435 86.230 142.650 86.775 ;
        RECT 141.425 85.905 141.755 86.095 ;
        RECT 141.975 85.735 142.690 86.030 ;
        RECT 142.860 85.905 143.135 86.605 ;
        RECT 141.005 85.565 142.795 85.735 ;
        RECT 140.595 85.135 141.390 85.385 ;
        RECT 140.595 85.045 140.845 85.135 ;
        RECT 136.110 84.225 136.350 84.735 ;
        RECT 136.530 84.405 136.810 84.735 ;
        RECT 137.040 84.225 137.255 84.735 ;
        RECT 137.425 84.395 138.040 84.965 ;
        RECT 138.705 84.225 138.995 84.950 ;
        RECT 140.085 84.225 140.345 85.045 ;
        RECT 140.515 84.625 140.845 85.045 ;
        RECT 141.560 84.710 141.815 85.565 ;
        RECT 141.025 84.445 141.815 84.710 ;
        RECT 141.985 84.865 142.395 85.385 ;
        RECT 142.565 85.135 142.795 85.565 ;
        RECT 142.965 84.875 143.135 85.905 ;
        RECT 143.305 85.685 145.895 86.775 ;
        RECT 141.985 84.445 142.185 84.865 ;
        RECT 142.375 84.225 142.705 84.685 ;
        RECT 142.875 84.395 143.135 84.875 ;
        RECT 143.305 84.995 144.515 85.515 ;
        RECT 144.685 85.165 145.895 85.685 ;
        RECT 146.065 85.635 146.325 86.775 ;
        RECT 146.495 85.625 146.825 86.605 ;
        RECT 146.995 85.635 147.275 86.775 ;
        RECT 147.445 85.685 148.655 86.775 ;
        RECT 146.085 85.215 146.420 85.465 ;
        RECT 146.590 85.025 146.760 85.625 ;
        RECT 146.930 85.195 147.265 85.465 ;
        RECT 143.305 84.225 145.895 84.995 ;
        RECT 146.065 84.395 146.760 85.025 ;
        RECT 146.965 84.225 147.275 85.025 ;
        RECT 147.445 84.975 147.965 85.515 ;
        RECT 148.135 85.145 148.655 85.685 ;
        RECT 148.860 85.985 149.395 86.605 ;
        RECT 147.445 84.225 148.655 84.975 ;
        RECT 148.860 84.965 149.175 85.985 ;
        RECT 149.565 85.975 149.895 86.775 ;
        RECT 150.380 85.805 150.770 85.980 ;
        RECT 149.345 85.635 150.770 85.805 ;
        RECT 151.125 85.685 154.635 86.775 ;
        RECT 149.345 85.135 149.515 85.635 ;
        RECT 148.860 84.395 149.475 84.965 ;
        RECT 149.765 84.905 150.030 85.465 ;
        RECT 150.200 84.735 150.370 85.635 ;
        RECT 150.540 84.905 150.895 85.465 ;
        RECT 151.125 84.995 152.775 85.515 ;
        RECT 152.945 85.165 154.635 85.685 ;
        RECT 155.725 85.685 156.935 86.775 ;
        RECT 155.725 85.145 156.245 85.685 ;
        RECT 149.645 84.225 149.860 84.735 ;
        RECT 150.090 84.405 150.370 84.735 ;
        RECT 150.550 84.225 150.790 84.735 ;
        RECT 151.125 84.225 154.635 84.995 ;
        RECT 156.415 84.975 156.935 85.515 ;
        RECT 155.725 84.225 156.935 84.975 ;
        RECT 22.700 84.055 157.020 84.225 ;
        RECT 22.785 83.305 23.995 84.055 ;
        RECT 22.785 82.765 23.305 83.305 ;
        RECT 24.165 83.285 25.835 84.055 ;
        RECT 26.185 83.395 26.525 84.055 ;
        RECT 23.475 82.595 23.995 83.135 ;
        RECT 24.165 82.765 24.915 83.285 ;
        RECT 25.085 82.595 25.835 83.115 ;
        RECT 22.785 81.505 23.995 82.595 ;
        RECT 24.165 81.505 25.835 82.595 ;
        RECT 26.005 81.675 26.525 83.225 ;
        RECT 26.695 82.400 27.215 83.885 ;
        RECT 27.385 83.285 30.895 84.055 ;
        RECT 31.985 83.380 32.245 83.885 ;
        RECT 32.425 83.675 32.755 84.055 ;
        RECT 32.935 83.505 33.105 83.885 ;
        RECT 27.385 82.765 29.035 83.285 ;
        RECT 29.205 82.595 30.895 83.115 ;
        RECT 26.695 81.505 27.025 82.230 ;
        RECT 27.385 81.505 30.895 82.595 ;
        RECT 31.985 82.580 32.155 83.380 ;
        RECT 32.440 83.335 33.105 83.505 ;
        RECT 32.440 83.080 32.610 83.335 ;
        RECT 33.365 83.285 35.035 84.055 ;
        RECT 32.325 82.750 32.610 83.080 ;
        RECT 32.845 82.785 33.175 83.155 ;
        RECT 33.365 82.765 34.115 83.285 ;
        RECT 35.205 83.255 35.515 84.055 ;
        RECT 35.720 83.255 36.415 83.885 ;
        RECT 37.505 83.395 37.765 83.725 ;
        RECT 37.960 83.425 38.185 84.055 ;
        RECT 38.400 83.420 38.645 83.880 ;
        RECT 38.895 83.595 39.165 84.055 ;
        RECT 39.335 83.605 40.175 83.775 ;
        RECT 40.735 83.695 41.065 84.055 ;
        RECT 32.440 82.605 32.610 82.750 ;
        RECT 31.985 81.675 32.255 82.580 ;
        RECT 32.440 82.435 33.105 82.605 ;
        RECT 34.285 82.595 35.035 83.115 ;
        RECT 35.215 82.815 35.550 83.085 ;
        RECT 35.720 82.655 35.890 83.255 ;
        RECT 36.060 82.815 36.395 83.065 ;
        RECT 32.425 81.505 32.755 82.265 ;
        RECT 32.935 81.675 33.105 82.435 ;
        RECT 33.365 81.505 35.035 82.595 ;
        RECT 35.205 81.505 35.485 82.645 ;
        RECT 35.655 81.675 35.985 82.655 ;
        RECT 36.155 81.505 36.415 82.645 ;
        RECT 37.505 82.470 37.675 83.395 ;
        RECT 38.400 83.145 38.570 83.420 ;
        RECT 39.335 83.145 39.505 83.605 ;
        RECT 41.235 83.525 41.430 83.795 ;
        RECT 37.845 82.815 38.570 83.145 ;
        RECT 38.740 82.815 39.505 83.145 ;
        RECT 38.400 82.605 38.570 82.815 ;
        RECT 39.295 82.690 39.505 82.815 ;
        RECT 39.675 83.100 40.380 83.405 ;
        RECT 40.825 83.375 41.430 83.525 ;
        RECT 40.620 83.355 41.430 83.375 ;
        RECT 37.505 81.685 37.765 82.470 ;
        RECT 37.935 81.505 38.220 82.570 ;
        RECT 38.400 82.275 39.125 82.605 ;
        RECT 38.400 81.705 38.645 82.275 ;
        RECT 39.295 82.130 39.485 82.690 ;
        RECT 39.675 82.580 39.990 83.100 ;
        RECT 40.620 82.905 40.995 83.355 ;
        RECT 39.655 82.230 39.990 82.580 ;
        RECT 40.160 82.135 40.495 82.785 ;
        RECT 40.825 82.645 40.995 82.905 ;
        RECT 41.175 82.815 41.505 83.185 ;
        RECT 40.825 82.475 41.510 82.645 ;
        RECT 39.295 82.105 39.510 82.130 ;
        RECT 39.295 82.095 39.535 82.105 ;
        RECT 39.295 82.075 39.550 82.095 ;
        RECT 39.310 82.055 39.550 82.075 ;
        RECT 39.320 82.050 39.550 82.055 ;
        RECT 39.320 82.035 39.645 82.050 ;
        RECT 38.845 81.505 39.165 81.965 ;
        RECT 39.335 81.885 39.645 82.035 ;
        RECT 39.335 81.715 40.195 81.885 ;
        RECT 40.695 81.505 40.985 82.305 ;
        RECT 41.155 81.725 41.510 82.475 ;
        RECT 41.755 82.455 41.925 83.795 ;
        RECT 42.095 83.675 42.425 84.055 ;
        RECT 42.595 83.505 42.765 83.795 ;
        RECT 42.160 83.335 42.765 83.505 ;
        RECT 43.115 83.505 43.285 83.795 ;
        RECT 43.455 83.675 43.785 84.055 ;
        RECT 43.115 83.335 43.720 83.505 ;
        RECT 42.160 83.070 42.330 83.335 ;
        RECT 42.100 82.740 42.330 83.070 ;
        RECT 41.700 81.675 41.925 82.455 ;
        RECT 42.160 82.345 42.330 82.740 ;
        RECT 42.610 82.515 42.855 83.155 ;
        RECT 43.025 82.515 43.270 83.155 ;
        RECT 43.550 83.070 43.720 83.335 ;
        RECT 43.550 82.740 43.780 83.070 ;
        RECT 43.550 82.345 43.720 82.740 ;
        RECT 42.160 82.175 42.765 82.345 ;
        RECT 42.095 81.505 42.425 82.005 ;
        RECT 42.595 81.675 42.765 82.175 ;
        RECT 43.115 82.175 43.720 82.345 ;
        RECT 43.955 82.455 44.125 83.795 ;
        RECT 44.450 83.525 44.645 83.795 ;
        RECT 44.815 83.695 45.145 84.055 ;
        RECT 45.705 83.605 46.545 83.775 ;
        RECT 44.450 83.375 45.055 83.525 ;
        RECT 44.450 83.355 45.260 83.375 ;
        RECT 44.375 82.815 44.705 83.185 ;
        RECT 44.885 82.905 45.260 83.355 ;
        RECT 45.500 83.100 46.205 83.405 ;
        RECT 44.885 82.645 45.055 82.905 ;
        RECT 44.370 82.475 45.055 82.645 ;
        RECT 43.115 81.675 43.285 82.175 ;
        RECT 43.455 81.505 43.785 82.005 ;
        RECT 43.955 81.675 44.180 82.455 ;
        RECT 44.370 81.725 44.725 82.475 ;
        RECT 44.895 81.505 45.185 82.305 ;
        RECT 45.385 82.135 45.720 82.785 ;
        RECT 45.890 82.580 46.205 83.100 ;
        RECT 46.375 83.145 46.545 83.605 ;
        RECT 46.715 83.595 46.985 84.055 ;
        RECT 47.235 83.420 47.480 83.880 ;
        RECT 47.695 83.425 47.920 84.055 ;
        RECT 47.310 83.145 47.480 83.420 ;
        RECT 48.115 83.395 48.375 83.725 ;
        RECT 46.375 82.815 47.140 83.145 ;
        RECT 47.310 82.815 48.035 83.145 ;
        RECT 46.375 82.690 46.585 82.815 ;
        RECT 45.890 82.230 46.225 82.580 ;
        RECT 46.395 82.130 46.585 82.690 ;
        RECT 47.310 82.605 47.480 82.815 ;
        RECT 46.755 82.275 47.480 82.605 ;
        RECT 46.370 82.105 46.585 82.130 ;
        RECT 46.345 82.095 46.585 82.105 ;
        RECT 46.330 82.075 46.585 82.095 ;
        RECT 46.330 82.055 46.570 82.075 ;
        RECT 46.330 82.050 46.560 82.055 ;
        RECT 46.235 82.035 46.560 82.050 ;
        RECT 46.235 81.885 46.545 82.035 ;
        RECT 45.685 81.715 46.545 81.885 ;
        RECT 46.715 81.505 47.035 81.965 ;
        RECT 47.235 81.705 47.480 82.275 ;
        RECT 47.660 81.505 47.945 82.570 ;
        RECT 48.205 82.470 48.375 83.395 ;
        RECT 48.545 83.330 48.835 84.055 ;
        RECT 50.015 83.505 50.185 83.795 ;
        RECT 50.355 83.675 50.685 84.055 ;
        RECT 50.015 83.335 50.620 83.505 ;
        RECT 48.115 81.685 48.375 82.470 ;
        RECT 48.545 81.505 48.835 82.670 ;
        RECT 49.925 82.515 50.170 83.155 ;
        RECT 50.450 83.070 50.620 83.335 ;
        RECT 50.450 82.740 50.680 83.070 ;
        RECT 50.450 82.345 50.620 82.740 ;
        RECT 50.015 82.175 50.620 82.345 ;
        RECT 50.855 82.455 51.025 83.795 ;
        RECT 51.350 83.525 51.545 83.795 ;
        RECT 51.715 83.695 52.045 84.055 ;
        RECT 52.605 83.605 53.445 83.775 ;
        RECT 51.350 83.375 51.955 83.525 ;
        RECT 51.350 83.355 52.160 83.375 ;
        RECT 51.275 82.815 51.605 83.185 ;
        RECT 51.785 82.905 52.160 83.355 ;
        RECT 52.400 83.100 53.105 83.405 ;
        RECT 51.785 82.645 51.955 82.905 ;
        RECT 51.270 82.475 51.955 82.645 ;
        RECT 50.015 81.675 50.185 82.175 ;
        RECT 50.355 81.505 50.685 82.005 ;
        RECT 50.855 81.675 51.080 82.455 ;
        RECT 51.270 81.725 51.625 82.475 ;
        RECT 51.795 81.505 52.085 82.305 ;
        RECT 52.285 82.135 52.620 82.785 ;
        RECT 52.790 82.580 53.105 83.100 ;
        RECT 53.275 83.145 53.445 83.605 ;
        RECT 53.615 83.595 53.885 84.055 ;
        RECT 54.135 83.420 54.380 83.880 ;
        RECT 54.595 83.425 54.820 84.055 ;
        RECT 54.210 83.145 54.380 83.420 ;
        RECT 55.015 83.395 55.275 83.725 ;
        RECT 55.495 83.400 55.825 83.835 ;
        RECT 55.995 83.445 56.165 84.055 ;
        RECT 53.275 82.815 54.040 83.145 ;
        RECT 54.210 82.815 54.935 83.145 ;
        RECT 53.275 82.690 53.485 82.815 ;
        RECT 52.790 82.230 53.125 82.580 ;
        RECT 53.295 82.130 53.485 82.690 ;
        RECT 54.210 82.605 54.380 82.815 ;
        RECT 53.655 82.275 54.380 82.605 ;
        RECT 53.270 82.105 53.485 82.130 ;
        RECT 53.245 82.095 53.485 82.105 ;
        RECT 53.230 82.075 53.485 82.095 ;
        RECT 53.230 82.055 53.470 82.075 ;
        RECT 53.230 82.050 53.460 82.055 ;
        RECT 53.135 82.035 53.460 82.050 ;
        RECT 53.135 81.885 53.445 82.035 ;
        RECT 52.585 81.715 53.445 81.885 ;
        RECT 53.615 81.505 53.935 81.965 ;
        RECT 54.135 81.705 54.380 82.275 ;
        RECT 54.560 81.505 54.845 82.570 ;
        RECT 55.105 82.470 55.275 83.395 ;
        RECT 55.445 83.315 55.825 83.400 ;
        RECT 56.335 83.315 56.665 83.840 ;
        RECT 56.925 83.525 57.135 84.055 ;
        RECT 57.410 83.605 58.195 83.775 ;
        RECT 58.365 83.605 58.770 83.775 ;
        RECT 55.445 83.275 55.670 83.315 ;
        RECT 55.445 82.695 55.615 83.275 ;
        RECT 56.335 83.145 56.535 83.315 ;
        RECT 57.410 83.145 57.580 83.605 ;
        RECT 55.785 82.815 56.535 83.145 ;
        RECT 56.705 82.815 57.580 83.145 ;
        RECT 55.445 82.645 55.660 82.695 ;
        RECT 55.445 82.565 55.835 82.645 ;
        RECT 55.015 81.685 55.275 82.470 ;
        RECT 55.505 81.720 55.835 82.565 ;
        RECT 56.345 82.610 56.535 82.815 ;
        RECT 56.005 81.505 56.175 82.515 ;
        RECT 56.345 82.235 57.240 82.610 ;
        RECT 56.345 81.675 56.685 82.235 ;
        RECT 56.915 81.505 57.230 82.005 ;
        RECT 57.410 81.975 57.580 82.815 ;
        RECT 57.750 83.105 58.215 83.435 ;
        RECT 58.600 83.375 58.770 83.605 ;
        RECT 58.950 83.555 59.320 84.055 ;
        RECT 59.640 83.605 60.315 83.775 ;
        RECT 60.510 83.605 60.845 83.775 ;
        RECT 57.750 82.145 58.070 83.105 ;
        RECT 58.600 83.075 59.430 83.375 ;
        RECT 58.240 82.175 58.430 82.895 ;
        RECT 58.600 82.005 58.770 83.075 ;
        RECT 59.230 83.045 59.430 83.075 ;
        RECT 58.940 82.825 59.110 82.895 ;
        RECT 59.640 82.825 59.810 83.605 ;
        RECT 60.675 83.465 60.845 83.605 ;
        RECT 61.015 83.595 61.265 84.055 ;
        RECT 58.940 82.655 59.810 82.825 ;
        RECT 59.980 83.185 60.505 83.405 ;
        RECT 60.675 83.335 60.900 83.465 ;
        RECT 58.940 82.565 59.450 82.655 ;
        RECT 57.410 81.805 58.295 81.975 ;
        RECT 58.520 81.675 58.770 82.005 ;
        RECT 58.940 81.505 59.110 82.305 ;
        RECT 59.280 81.950 59.450 82.565 ;
        RECT 59.980 82.485 60.150 83.185 ;
        RECT 59.620 82.120 60.150 82.485 ;
        RECT 60.320 82.420 60.560 83.015 ;
        RECT 60.730 82.230 60.900 83.335 ;
        RECT 61.070 82.475 61.350 83.425 ;
        RECT 60.595 82.100 60.900 82.230 ;
        RECT 59.280 81.780 60.385 81.950 ;
        RECT 60.595 81.675 60.845 82.100 ;
        RECT 61.015 81.505 61.280 81.965 ;
        RECT 61.520 81.675 61.705 83.795 ;
        RECT 61.875 83.675 62.205 84.055 ;
        RECT 62.375 83.505 62.545 83.795 ;
        RECT 61.880 83.335 62.545 83.505 ;
        RECT 62.895 83.505 63.065 83.795 ;
        RECT 63.235 83.675 63.565 84.055 ;
        RECT 62.895 83.335 63.560 83.505 ;
        RECT 61.880 82.345 62.110 83.335 ;
        RECT 62.280 82.515 62.630 83.165 ;
        RECT 62.810 82.515 63.160 83.165 ;
        RECT 63.330 82.345 63.560 83.335 ;
        RECT 61.880 82.175 62.545 82.345 ;
        RECT 61.875 81.505 62.205 82.005 ;
        RECT 62.375 81.675 62.545 82.175 ;
        RECT 62.895 82.175 63.560 82.345 ;
        RECT 62.895 81.675 63.065 82.175 ;
        RECT 63.235 81.505 63.565 82.005 ;
        RECT 63.735 81.675 63.920 83.795 ;
        RECT 64.175 83.595 64.425 84.055 ;
        RECT 64.595 83.605 64.930 83.775 ;
        RECT 65.125 83.605 65.800 83.775 ;
        RECT 64.595 83.465 64.765 83.605 ;
        RECT 64.090 82.475 64.370 83.425 ;
        RECT 64.540 83.335 64.765 83.465 ;
        RECT 64.540 82.230 64.710 83.335 ;
        RECT 64.935 83.185 65.460 83.405 ;
        RECT 64.880 82.420 65.120 83.015 ;
        RECT 65.290 82.485 65.460 83.185 ;
        RECT 65.630 82.825 65.800 83.605 ;
        RECT 66.120 83.555 66.490 84.055 ;
        RECT 66.670 83.605 67.075 83.775 ;
        RECT 67.245 83.605 68.030 83.775 ;
        RECT 66.670 83.375 66.840 83.605 ;
        RECT 66.010 83.075 66.840 83.375 ;
        RECT 67.225 83.105 67.690 83.435 ;
        RECT 66.010 83.045 66.210 83.075 ;
        RECT 66.330 82.825 66.500 82.895 ;
        RECT 65.630 82.655 66.500 82.825 ;
        RECT 65.990 82.565 66.500 82.655 ;
        RECT 64.540 82.100 64.845 82.230 ;
        RECT 65.290 82.120 65.820 82.485 ;
        RECT 64.160 81.505 64.425 81.965 ;
        RECT 64.595 81.675 64.845 82.100 ;
        RECT 65.990 81.950 66.160 82.565 ;
        RECT 65.055 81.780 66.160 81.950 ;
        RECT 66.330 81.505 66.500 82.305 ;
        RECT 66.670 82.005 66.840 83.075 ;
        RECT 67.010 82.175 67.200 82.895 ;
        RECT 67.370 82.145 67.690 83.105 ;
        RECT 67.860 83.145 68.030 83.605 ;
        RECT 68.305 83.525 68.515 84.055 ;
        RECT 68.775 83.315 69.105 83.840 ;
        RECT 69.275 83.445 69.445 84.055 ;
        RECT 69.615 83.400 69.945 83.835 ;
        RECT 69.615 83.315 69.995 83.400 ;
        RECT 68.905 83.145 69.105 83.315 ;
        RECT 69.770 83.275 69.995 83.315 ;
        RECT 67.860 82.815 68.735 83.145 ;
        RECT 68.905 82.815 69.655 83.145 ;
        RECT 66.670 81.675 66.920 82.005 ;
        RECT 67.860 81.975 68.030 82.815 ;
        RECT 68.905 82.610 69.095 82.815 ;
        RECT 69.825 82.695 69.995 83.275 ;
        RECT 69.780 82.645 69.995 82.695 ;
        RECT 68.200 82.235 69.095 82.610 ;
        RECT 69.605 82.565 69.995 82.645 ;
        RECT 70.200 83.315 70.815 83.885 ;
        RECT 70.985 83.545 71.200 84.055 ;
        RECT 71.430 83.545 71.710 83.875 ;
        RECT 71.890 83.545 72.130 84.055 ;
        RECT 67.145 81.805 68.030 81.975 ;
        RECT 68.210 81.505 68.525 82.005 ;
        RECT 68.755 81.675 69.095 82.235 ;
        RECT 69.265 81.505 69.435 82.515 ;
        RECT 69.605 81.720 69.935 82.565 ;
        RECT 70.200 82.295 70.515 83.315 ;
        RECT 70.685 82.645 70.855 83.145 ;
        RECT 71.105 82.815 71.370 83.375 ;
        RECT 71.540 82.645 71.710 83.545 ;
        RECT 71.880 82.815 72.235 83.375 ;
        RECT 72.465 83.255 73.160 83.885 ;
        RECT 73.365 83.255 73.675 84.055 ;
        RECT 74.305 83.330 74.595 84.055 ;
        RECT 74.765 83.510 80.110 84.055 ;
        RECT 72.485 82.815 72.820 83.065 ;
        RECT 72.990 82.655 73.160 83.255 ;
        RECT 73.330 82.815 73.665 83.085 ;
        RECT 76.350 82.680 76.690 83.510 ;
        RECT 80.285 83.285 81.955 84.055 ;
        RECT 82.305 83.395 82.645 84.055 ;
        RECT 70.685 82.475 72.110 82.645 ;
        RECT 70.200 81.675 70.735 82.295 ;
        RECT 70.905 81.505 71.235 82.305 ;
        RECT 71.720 82.300 72.110 82.475 ;
        RECT 72.465 81.505 72.725 82.645 ;
        RECT 72.895 81.675 73.225 82.655 ;
        RECT 73.395 81.505 73.675 82.645 ;
        RECT 74.305 81.505 74.595 82.670 ;
        RECT 78.170 81.940 78.520 83.190 ;
        RECT 80.285 82.765 81.035 83.285 ;
        RECT 81.205 82.595 81.955 83.115 ;
        RECT 74.765 81.505 80.110 81.940 ;
        RECT 80.285 81.505 81.955 82.595 ;
        RECT 82.125 81.675 82.645 83.225 ;
        RECT 82.815 82.400 83.335 83.885 ;
        RECT 83.505 83.510 88.850 84.055 ;
        RECT 89.190 83.545 89.430 84.055 ;
        RECT 89.610 83.545 89.890 83.875 ;
        RECT 90.120 83.545 90.335 84.055 ;
        RECT 85.090 82.680 85.430 83.510 ;
        RECT 82.815 81.505 83.145 82.230 ;
        RECT 86.910 81.940 87.260 83.190 ;
        RECT 89.085 82.815 89.440 83.375 ;
        RECT 89.610 82.645 89.780 83.545 ;
        RECT 89.950 82.815 90.215 83.375 ;
        RECT 90.505 83.315 91.120 83.885 ;
        RECT 91.835 83.400 92.165 83.835 ;
        RECT 92.335 83.445 92.505 84.055 ;
        RECT 90.465 82.645 90.635 83.145 ;
        RECT 89.210 82.475 90.635 82.645 ;
        RECT 89.210 82.300 89.600 82.475 ;
        RECT 83.505 81.505 88.850 81.940 ;
        RECT 90.085 81.505 90.415 82.305 ;
        RECT 90.805 82.295 91.120 83.315 ;
        RECT 91.785 83.315 92.165 83.400 ;
        RECT 92.675 83.315 93.005 83.840 ;
        RECT 93.265 83.525 93.475 84.055 ;
        RECT 93.750 83.605 94.535 83.775 ;
        RECT 94.705 83.605 95.110 83.775 ;
        RECT 91.785 83.275 92.010 83.315 ;
        RECT 91.785 82.695 91.955 83.275 ;
        RECT 92.675 83.145 92.875 83.315 ;
        RECT 93.750 83.145 93.920 83.605 ;
        RECT 92.125 82.815 92.875 83.145 ;
        RECT 93.045 82.815 93.920 83.145 ;
        RECT 91.785 82.645 92.000 82.695 ;
        RECT 91.785 82.565 92.175 82.645 ;
        RECT 90.585 81.675 91.120 82.295 ;
        RECT 91.845 81.720 92.175 82.565 ;
        RECT 92.685 82.610 92.875 82.815 ;
        RECT 92.345 81.505 92.515 82.515 ;
        RECT 92.685 82.235 93.580 82.610 ;
        RECT 92.685 81.675 93.025 82.235 ;
        RECT 93.255 81.505 93.570 82.005 ;
        RECT 93.750 81.975 93.920 82.815 ;
        RECT 94.090 83.105 94.555 83.435 ;
        RECT 94.940 83.375 95.110 83.605 ;
        RECT 95.290 83.555 95.660 84.055 ;
        RECT 95.980 83.605 96.655 83.775 ;
        RECT 96.850 83.605 97.185 83.775 ;
        RECT 94.090 82.145 94.410 83.105 ;
        RECT 94.940 83.075 95.770 83.375 ;
        RECT 94.580 82.175 94.770 82.895 ;
        RECT 94.940 82.005 95.110 83.075 ;
        RECT 95.570 83.045 95.770 83.075 ;
        RECT 95.280 82.825 95.450 82.895 ;
        RECT 95.980 82.825 96.150 83.605 ;
        RECT 97.015 83.465 97.185 83.605 ;
        RECT 97.355 83.595 97.605 84.055 ;
        RECT 95.280 82.655 96.150 82.825 ;
        RECT 96.320 83.185 96.845 83.405 ;
        RECT 97.015 83.335 97.240 83.465 ;
        RECT 95.280 82.565 95.790 82.655 ;
        RECT 93.750 81.805 94.635 81.975 ;
        RECT 94.860 81.675 95.110 82.005 ;
        RECT 95.280 81.505 95.450 82.305 ;
        RECT 95.620 81.950 95.790 82.565 ;
        RECT 96.320 82.485 96.490 83.185 ;
        RECT 95.960 82.120 96.490 82.485 ;
        RECT 96.660 82.420 96.900 83.015 ;
        RECT 97.070 82.230 97.240 83.335 ;
        RECT 97.410 82.475 97.690 83.425 ;
        RECT 96.935 82.100 97.240 82.230 ;
        RECT 95.620 81.780 96.725 81.950 ;
        RECT 96.935 81.675 97.185 82.100 ;
        RECT 97.355 81.505 97.620 81.965 ;
        RECT 97.860 81.675 98.045 83.795 ;
        RECT 98.215 83.675 98.545 84.055 ;
        RECT 98.715 83.505 98.885 83.795 ;
        RECT 98.220 83.335 98.885 83.505 ;
        RECT 98.220 82.345 98.450 83.335 ;
        RECT 100.065 83.330 100.355 84.055 ;
        RECT 101.075 83.505 101.245 83.885 ;
        RECT 101.425 83.675 101.755 84.055 ;
        RECT 101.075 83.335 101.740 83.505 ;
        RECT 101.935 83.380 102.195 83.885 ;
        RECT 98.620 82.515 98.970 83.165 ;
        RECT 101.005 82.785 101.335 83.155 ;
        RECT 101.570 83.080 101.740 83.335 ;
        RECT 101.570 82.750 101.855 83.080 ;
        RECT 98.220 82.175 98.885 82.345 ;
        RECT 98.215 81.505 98.545 82.005 ;
        RECT 98.715 81.675 98.885 82.175 ;
        RECT 100.065 81.505 100.355 82.670 ;
        RECT 101.570 82.605 101.740 82.750 ;
        RECT 101.075 82.435 101.740 82.605 ;
        RECT 102.025 82.580 102.195 83.380 ;
        RECT 101.075 81.675 101.245 82.435 ;
        RECT 101.425 81.505 101.755 82.265 ;
        RECT 101.925 81.675 102.195 82.580 ;
        RECT 102.380 81.685 102.660 83.875 ;
        RECT 102.860 83.685 103.590 84.055 ;
        RECT 104.170 83.515 104.600 83.875 ;
        RECT 102.860 83.325 104.600 83.515 ;
        RECT 102.860 82.815 103.120 83.325 ;
        RECT 102.850 81.505 103.135 82.645 ;
        RECT 103.330 82.525 103.590 83.145 ;
        RECT 103.785 82.525 104.210 83.145 ;
        RECT 104.380 83.095 104.600 83.325 ;
        RECT 104.770 83.275 105.015 84.055 ;
        RECT 104.380 82.795 104.925 83.095 ;
        RECT 105.215 82.975 105.445 83.875 ;
        RECT 103.400 82.155 104.425 82.355 ;
        RECT 103.400 81.685 103.570 82.155 ;
        RECT 103.745 81.505 104.075 81.985 ;
        RECT 104.245 81.685 104.425 82.155 ;
        RECT 104.595 81.685 104.925 82.795 ;
        RECT 105.105 82.295 105.445 82.975 ;
        RECT 105.625 82.475 105.855 83.815 ;
        RECT 106.045 83.405 106.305 83.885 ;
        RECT 106.475 83.595 106.805 84.055 ;
        RECT 106.995 83.415 107.195 83.835 ;
        RECT 106.045 82.375 106.215 83.405 ;
        RECT 106.385 82.715 106.615 83.145 ;
        RECT 106.785 82.895 107.195 83.415 ;
        RECT 107.365 83.570 108.155 83.835 ;
        RECT 107.365 82.715 107.620 83.570 ;
        RECT 108.335 83.235 108.665 83.655 ;
        RECT 108.835 83.235 109.095 84.055 ;
        RECT 109.430 83.545 109.670 84.055 ;
        RECT 109.850 83.545 110.130 83.875 ;
        RECT 110.360 83.545 110.575 84.055 ;
        RECT 108.335 83.145 108.585 83.235 ;
        RECT 107.790 82.895 108.585 83.145 ;
        RECT 106.385 82.545 108.175 82.715 ;
        RECT 105.105 82.095 105.855 82.295 ;
        RECT 105.095 81.505 105.445 81.915 ;
        RECT 105.615 81.705 105.855 82.095 ;
        RECT 106.045 81.675 106.320 82.375 ;
        RECT 106.490 82.250 107.205 82.545 ;
        RECT 107.425 82.185 107.755 82.375 ;
        RECT 106.530 81.505 106.745 82.050 ;
        RECT 106.915 81.675 107.390 82.015 ;
        RECT 107.560 82.010 107.755 82.185 ;
        RECT 107.925 82.180 108.175 82.545 ;
        RECT 107.560 81.505 108.175 82.010 ;
        RECT 108.415 81.675 108.585 82.895 ;
        RECT 108.755 82.185 109.095 83.065 ;
        RECT 109.325 82.815 109.680 83.375 ;
        RECT 109.850 82.645 110.020 83.545 ;
        RECT 110.190 82.815 110.455 83.375 ;
        RECT 110.745 83.315 111.360 83.885 ;
        RECT 111.745 83.395 112.085 84.055 ;
        RECT 110.705 82.645 110.875 83.145 ;
        RECT 109.450 82.475 110.875 82.645 ;
        RECT 109.450 82.300 109.840 82.475 ;
        RECT 108.835 81.505 109.095 82.015 ;
        RECT 110.325 81.505 110.655 82.305 ;
        RECT 111.045 82.295 111.360 83.315 ;
        RECT 110.825 81.675 111.360 82.295 ;
        RECT 111.565 81.675 112.085 83.225 ;
        RECT 112.255 82.400 112.775 83.885 ;
        RECT 112.945 83.285 114.615 84.055 ;
        RECT 114.965 83.395 115.305 84.055 ;
        RECT 112.945 82.765 113.695 83.285 ;
        RECT 113.865 82.595 114.615 83.115 ;
        RECT 112.255 81.505 112.585 82.230 ;
        RECT 112.945 81.505 114.615 82.595 ;
        RECT 114.785 81.675 115.305 83.225 ;
        RECT 115.475 82.400 115.995 83.885 ;
        RECT 116.805 83.395 117.145 84.055 ;
        RECT 115.475 81.505 115.805 82.230 ;
        RECT 116.625 81.675 117.145 83.225 ;
        RECT 117.315 82.400 117.835 83.885 ;
        RECT 118.555 83.505 118.725 83.795 ;
        RECT 118.895 83.675 119.225 84.055 ;
        RECT 118.555 83.335 119.160 83.505 ;
        RECT 118.465 82.515 118.710 83.155 ;
        RECT 118.990 83.070 119.160 83.335 ;
        RECT 118.990 82.740 119.220 83.070 ;
        RECT 118.990 82.345 119.160 82.740 ;
        RECT 117.315 81.505 117.645 82.230 ;
        RECT 118.555 82.175 119.160 82.345 ;
        RECT 119.395 82.455 119.565 83.795 ;
        RECT 119.890 83.525 120.085 83.795 ;
        RECT 120.255 83.695 120.585 84.055 ;
        RECT 121.145 83.605 121.985 83.775 ;
        RECT 119.890 83.375 120.495 83.525 ;
        RECT 119.890 83.355 120.700 83.375 ;
        RECT 119.815 82.815 120.145 83.185 ;
        RECT 120.325 82.905 120.700 83.355 ;
        RECT 120.940 83.100 121.645 83.405 ;
        RECT 120.325 82.645 120.495 82.905 ;
        RECT 119.810 82.475 120.495 82.645 ;
        RECT 118.555 81.675 118.725 82.175 ;
        RECT 118.895 81.505 119.225 82.005 ;
        RECT 119.395 81.675 119.620 82.455 ;
        RECT 119.810 81.725 120.165 82.475 ;
        RECT 120.335 81.505 120.625 82.305 ;
        RECT 120.825 82.135 121.160 82.785 ;
        RECT 121.330 82.580 121.645 83.100 ;
        RECT 121.815 83.145 121.985 83.605 ;
        RECT 122.155 83.595 122.425 84.055 ;
        RECT 122.675 83.420 122.920 83.880 ;
        RECT 123.135 83.425 123.360 84.055 ;
        RECT 122.750 83.145 122.920 83.420 ;
        RECT 123.555 83.395 123.815 83.725 ;
        RECT 121.815 82.815 122.580 83.145 ;
        RECT 122.750 82.815 123.475 83.145 ;
        RECT 121.815 82.690 122.025 82.815 ;
        RECT 121.330 82.230 121.665 82.580 ;
        RECT 121.835 82.130 122.025 82.690 ;
        RECT 122.750 82.605 122.920 82.815 ;
        RECT 122.195 82.275 122.920 82.605 ;
        RECT 121.810 82.105 122.025 82.130 ;
        RECT 121.785 82.095 122.025 82.105 ;
        RECT 121.770 82.075 122.025 82.095 ;
        RECT 121.770 82.055 122.010 82.075 ;
        RECT 121.770 82.050 122.000 82.055 ;
        RECT 121.675 82.035 122.000 82.050 ;
        RECT 121.675 81.885 121.985 82.035 ;
        RECT 121.125 81.715 121.985 81.885 ;
        RECT 122.155 81.505 122.475 81.965 ;
        RECT 122.675 81.705 122.920 82.275 ;
        RECT 123.100 81.505 123.385 82.570 ;
        RECT 123.645 82.470 123.815 83.395 ;
        RECT 123.555 81.685 123.815 82.470 ;
        RECT 124.445 83.380 124.705 83.885 ;
        RECT 124.885 83.675 125.215 84.055 ;
        RECT 125.395 83.505 125.565 83.885 ;
        RECT 124.445 82.580 124.615 83.380 ;
        RECT 124.900 83.335 125.565 83.505 ;
        RECT 124.900 83.080 125.070 83.335 ;
        RECT 125.825 83.330 126.115 84.055 ;
        RECT 126.285 83.405 126.545 83.885 ;
        RECT 126.715 83.515 126.965 84.055 ;
        RECT 124.785 82.750 125.070 83.080 ;
        RECT 125.305 82.785 125.635 83.155 ;
        RECT 124.900 82.605 125.070 82.750 ;
        RECT 124.445 81.675 124.715 82.580 ;
        RECT 124.900 82.435 125.565 82.605 ;
        RECT 124.885 81.505 125.215 82.265 ;
        RECT 125.395 81.675 125.565 82.435 ;
        RECT 125.825 81.505 126.115 82.670 ;
        RECT 126.285 82.375 126.455 83.405 ;
        RECT 127.135 83.350 127.355 83.835 ;
        RECT 126.625 82.755 126.855 83.150 ;
        RECT 127.025 82.925 127.355 83.350 ;
        RECT 127.525 83.675 128.415 83.845 ;
        RECT 127.525 82.950 127.695 83.675 ;
        RECT 128.750 83.545 128.990 84.055 ;
        RECT 129.170 83.545 129.450 83.875 ;
        RECT 129.680 83.545 129.895 84.055 ;
        RECT 127.865 83.120 128.415 83.505 ;
        RECT 127.525 82.880 128.415 82.950 ;
        RECT 127.520 82.855 128.415 82.880 ;
        RECT 127.510 82.840 128.415 82.855 ;
        RECT 127.505 82.825 128.415 82.840 ;
        RECT 127.495 82.820 128.415 82.825 ;
        RECT 127.490 82.810 128.415 82.820 ;
        RECT 128.645 82.815 129.000 83.375 ;
        RECT 127.485 82.800 128.415 82.810 ;
        RECT 127.475 82.795 128.415 82.800 ;
        RECT 127.465 82.785 128.415 82.795 ;
        RECT 127.455 82.780 128.415 82.785 ;
        RECT 127.455 82.775 127.790 82.780 ;
        RECT 127.440 82.770 127.790 82.775 ;
        RECT 127.425 82.760 127.790 82.770 ;
        RECT 127.400 82.755 127.790 82.760 ;
        RECT 126.625 82.750 127.790 82.755 ;
        RECT 126.625 82.715 127.760 82.750 ;
        RECT 126.625 82.690 127.725 82.715 ;
        RECT 126.625 82.660 127.695 82.690 ;
        RECT 126.625 82.630 127.675 82.660 ;
        RECT 126.625 82.600 127.655 82.630 ;
        RECT 126.625 82.590 127.585 82.600 ;
        RECT 126.625 82.580 127.560 82.590 ;
        RECT 126.625 82.565 127.540 82.580 ;
        RECT 126.625 82.550 127.520 82.565 ;
        RECT 126.730 82.540 127.515 82.550 ;
        RECT 126.730 82.505 127.500 82.540 ;
        RECT 126.285 81.675 126.560 82.375 ;
        RECT 126.730 82.255 127.485 82.505 ;
        RECT 127.655 82.185 127.985 82.430 ;
        RECT 128.155 82.330 128.415 82.780 ;
        RECT 129.170 82.645 129.340 83.545 ;
        RECT 129.510 82.815 129.775 83.375 ;
        RECT 130.065 83.315 130.680 83.885 ;
        RECT 130.025 82.645 130.195 83.145 ;
        RECT 128.770 82.475 130.195 82.645 ;
        RECT 128.770 82.300 129.160 82.475 ;
        RECT 127.800 82.160 127.985 82.185 ;
        RECT 127.800 82.060 128.415 82.160 ;
        RECT 126.730 81.505 126.985 82.050 ;
        RECT 127.155 81.675 127.635 82.015 ;
        RECT 127.810 81.505 128.415 82.060 ;
        RECT 129.645 81.505 129.975 82.305 ;
        RECT 130.365 82.295 130.680 83.315 ;
        RECT 130.885 83.285 132.555 84.055 ;
        RECT 132.905 83.395 133.245 84.055 ;
        RECT 130.885 82.765 131.635 83.285 ;
        RECT 131.805 82.595 132.555 83.115 ;
        RECT 130.145 81.675 130.680 82.295 ;
        RECT 130.885 81.505 132.555 82.595 ;
        RECT 132.725 81.675 133.245 83.225 ;
        RECT 133.415 82.400 133.935 83.885 ;
        RECT 134.565 83.255 135.260 83.885 ;
        RECT 135.465 83.255 135.775 84.055 ;
        RECT 135.945 83.510 141.290 84.055 ;
        RECT 134.585 82.815 134.920 83.065 ;
        RECT 135.090 82.655 135.260 83.255 ;
        RECT 135.430 82.815 135.765 83.085 ;
        RECT 137.530 82.680 137.870 83.510 ;
        RECT 141.465 83.235 141.725 84.055 ;
        RECT 141.895 83.235 142.225 83.655 ;
        RECT 142.405 83.570 143.195 83.835 ;
        RECT 133.415 81.505 133.745 82.230 ;
        RECT 134.565 81.505 134.825 82.645 ;
        RECT 134.995 81.675 135.325 82.655 ;
        RECT 135.495 81.505 135.775 82.645 ;
        RECT 139.350 81.940 139.700 83.190 ;
        RECT 141.975 83.145 142.225 83.235 ;
        RECT 141.465 82.185 141.805 83.065 ;
        RECT 141.975 82.895 142.770 83.145 ;
        RECT 135.945 81.505 141.290 81.940 ;
        RECT 141.465 81.505 141.725 82.015 ;
        RECT 141.975 81.675 142.145 82.895 ;
        RECT 142.940 82.715 143.195 83.570 ;
        RECT 143.365 83.415 143.565 83.835 ;
        RECT 143.755 83.595 144.085 84.055 ;
        RECT 143.365 82.895 143.775 83.415 ;
        RECT 144.255 83.405 144.515 83.885 ;
        RECT 143.945 82.715 144.175 83.145 ;
        RECT 142.385 82.545 144.175 82.715 ;
        RECT 142.385 82.180 142.635 82.545 ;
        RECT 142.805 82.185 143.135 82.375 ;
        RECT 143.355 82.250 144.070 82.545 ;
        RECT 144.345 82.375 144.515 83.405 ;
        RECT 144.745 83.235 144.955 84.055 ;
        RECT 145.125 83.255 145.455 83.885 ;
        RECT 145.125 82.655 145.375 83.255 ;
        RECT 145.625 83.235 145.855 84.055 ;
        RECT 146.155 83.505 146.325 83.885 ;
        RECT 146.505 83.675 146.835 84.055 ;
        RECT 146.155 83.335 146.820 83.505 ;
        RECT 147.015 83.380 147.275 83.885 ;
        RECT 145.545 82.815 145.875 83.065 ;
        RECT 146.085 82.785 146.415 83.155 ;
        RECT 146.650 83.080 146.820 83.335 ;
        RECT 146.650 82.750 146.935 83.080 ;
        RECT 142.805 82.010 143.000 82.185 ;
        RECT 142.385 81.505 143.000 82.010 ;
        RECT 143.170 81.675 143.645 82.015 ;
        RECT 143.815 81.505 144.030 82.050 ;
        RECT 144.240 81.675 144.515 82.375 ;
        RECT 144.745 81.505 144.955 82.645 ;
        RECT 145.125 81.675 145.455 82.655 ;
        RECT 145.625 81.505 145.855 82.645 ;
        RECT 146.650 82.605 146.820 82.750 ;
        RECT 146.155 82.435 146.820 82.605 ;
        RECT 147.105 82.580 147.275 83.380 ;
        RECT 147.445 83.255 148.140 83.885 ;
        RECT 148.345 83.255 148.655 84.055 ;
        RECT 148.825 83.285 151.415 84.055 ;
        RECT 151.585 83.330 151.875 84.055 ;
        RECT 152.045 83.285 155.555 84.055 ;
        RECT 155.725 83.305 156.935 84.055 ;
        RECT 147.465 82.815 147.800 83.065 ;
        RECT 147.970 82.695 148.140 83.255 ;
        RECT 148.310 82.815 148.645 83.085 ;
        RECT 148.825 82.765 150.035 83.285 ;
        RECT 147.965 82.655 148.140 82.695 ;
        RECT 146.155 81.675 146.325 82.435 ;
        RECT 146.505 81.505 146.835 82.265 ;
        RECT 147.005 81.675 147.275 82.580 ;
        RECT 147.445 81.505 147.705 82.645 ;
        RECT 147.875 81.675 148.205 82.655 ;
        RECT 148.375 81.505 148.655 82.645 ;
        RECT 150.205 82.595 151.415 83.115 ;
        RECT 152.045 82.765 153.695 83.285 ;
        RECT 148.825 81.505 151.415 82.595 ;
        RECT 151.585 81.505 151.875 82.670 ;
        RECT 153.865 82.595 155.555 83.115 ;
        RECT 152.045 81.505 155.555 82.595 ;
        RECT 155.725 82.595 156.245 83.135 ;
        RECT 156.415 82.765 156.935 83.305 ;
        RECT 155.725 81.505 156.935 82.595 ;
        RECT 22.700 81.335 157.020 81.505 ;
        RECT 22.785 80.245 23.995 81.335 ;
        RECT 24.165 80.245 26.755 81.335 ;
        RECT 22.785 79.535 23.305 80.075 ;
        RECT 23.475 79.705 23.995 80.245 ;
        RECT 24.165 79.555 25.375 80.075 ;
        RECT 25.545 79.725 26.755 80.245 ;
        RECT 26.925 80.260 27.195 81.165 ;
        RECT 27.365 80.575 27.695 81.335 ;
        RECT 27.875 80.405 28.045 81.165 ;
        RECT 28.395 80.665 28.565 81.165 ;
        RECT 28.735 80.835 29.065 81.335 ;
        RECT 28.395 80.495 29.060 80.665 ;
        RECT 22.785 78.785 23.995 79.535 ;
        RECT 24.165 78.785 26.755 79.555 ;
        RECT 26.925 79.460 27.095 80.260 ;
        RECT 27.380 80.235 28.045 80.405 ;
        RECT 27.380 80.090 27.550 80.235 ;
        RECT 27.265 79.760 27.550 80.090 ;
        RECT 27.380 79.505 27.550 79.760 ;
        RECT 27.785 79.685 28.115 80.055 ;
        RECT 28.310 79.675 28.660 80.325 ;
        RECT 28.830 79.505 29.060 80.495 ;
        RECT 26.925 78.955 27.185 79.460 ;
        RECT 27.380 79.335 28.045 79.505 ;
        RECT 27.365 78.785 27.695 79.165 ;
        RECT 27.875 78.955 28.045 79.335 ;
        RECT 28.395 79.335 29.060 79.505 ;
        RECT 28.395 79.045 28.565 79.335 ;
        RECT 28.735 78.785 29.065 79.165 ;
        RECT 29.235 79.045 29.420 81.165 ;
        RECT 29.660 80.875 29.925 81.335 ;
        RECT 30.095 80.740 30.345 81.165 ;
        RECT 30.555 80.890 31.660 81.060 ;
        RECT 30.040 80.610 30.345 80.740 ;
        RECT 29.590 79.415 29.870 80.365 ;
        RECT 30.040 79.505 30.210 80.610 ;
        RECT 30.380 79.825 30.620 80.420 ;
        RECT 30.790 80.355 31.320 80.720 ;
        RECT 30.790 79.655 30.960 80.355 ;
        RECT 31.490 80.275 31.660 80.890 ;
        RECT 31.830 80.535 32.000 81.335 ;
        RECT 32.170 80.835 32.420 81.165 ;
        RECT 32.645 80.865 33.530 81.035 ;
        RECT 31.490 80.185 32.000 80.275 ;
        RECT 30.040 79.375 30.265 79.505 ;
        RECT 30.435 79.435 30.960 79.655 ;
        RECT 31.130 80.015 32.000 80.185 ;
        RECT 29.675 78.785 29.925 79.245 ;
        RECT 30.095 79.235 30.265 79.375 ;
        RECT 31.130 79.235 31.300 80.015 ;
        RECT 31.830 79.945 32.000 80.015 ;
        RECT 31.510 79.765 31.710 79.795 ;
        RECT 32.170 79.765 32.340 80.835 ;
        RECT 32.510 79.945 32.700 80.665 ;
        RECT 31.510 79.465 32.340 79.765 ;
        RECT 32.870 79.735 33.190 80.695 ;
        RECT 30.095 79.065 30.430 79.235 ;
        RECT 30.625 79.065 31.300 79.235 ;
        RECT 31.620 78.785 31.990 79.285 ;
        RECT 32.170 79.235 32.340 79.465 ;
        RECT 32.725 79.405 33.190 79.735 ;
        RECT 33.360 80.025 33.530 80.865 ;
        RECT 33.710 80.835 34.025 81.335 ;
        RECT 34.255 80.605 34.595 81.165 ;
        RECT 33.700 80.230 34.595 80.605 ;
        RECT 34.765 80.325 34.935 81.335 ;
        RECT 34.405 80.025 34.595 80.230 ;
        RECT 35.105 80.275 35.435 81.120 ;
        RECT 35.105 80.195 35.495 80.275 ;
        RECT 35.280 80.145 35.495 80.195 ;
        RECT 35.665 80.170 35.955 81.335 ;
        RECT 36.310 80.365 36.700 80.540 ;
        RECT 37.185 80.535 37.515 81.335 ;
        RECT 37.685 80.545 38.220 81.165 ;
        RECT 39.535 80.610 39.865 81.335 ;
        RECT 36.310 80.195 37.735 80.365 ;
        RECT 33.360 79.695 34.235 80.025 ;
        RECT 34.405 79.695 35.155 80.025 ;
        RECT 33.360 79.235 33.530 79.695 ;
        RECT 34.405 79.525 34.605 79.695 ;
        RECT 35.325 79.565 35.495 80.145 ;
        RECT 35.270 79.525 35.495 79.565 ;
        RECT 32.170 79.065 32.575 79.235 ;
        RECT 32.745 79.065 33.530 79.235 ;
        RECT 33.805 78.785 34.015 79.315 ;
        RECT 34.275 79.000 34.605 79.525 ;
        RECT 35.115 79.440 35.495 79.525 ;
        RECT 34.775 78.785 34.945 79.395 ;
        RECT 35.115 79.005 35.445 79.440 ;
        RECT 35.665 78.785 35.955 79.510 ;
        RECT 36.185 79.465 36.540 80.025 ;
        RECT 36.710 79.295 36.880 80.195 ;
        RECT 37.050 79.465 37.315 80.025 ;
        RECT 37.565 79.695 37.735 80.195 ;
        RECT 37.905 79.525 38.220 80.545 ;
        RECT 36.290 78.785 36.530 79.295 ;
        RECT 36.710 78.965 36.990 79.295 ;
        RECT 37.220 78.785 37.435 79.295 ;
        RECT 37.605 78.955 38.220 79.525 ;
        RECT 39.345 78.955 39.865 80.440 ;
        RECT 40.035 79.615 40.555 81.165 ;
        RECT 40.815 80.665 40.985 81.165 ;
        RECT 41.155 80.835 41.485 81.335 ;
        RECT 40.815 80.495 41.420 80.665 ;
        RECT 40.725 79.685 40.970 80.325 ;
        RECT 41.250 80.100 41.420 80.495 ;
        RECT 41.655 80.385 41.880 81.165 ;
        RECT 41.250 79.770 41.480 80.100 ;
        RECT 41.250 79.505 41.420 79.770 ;
        RECT 40.035 78.785 40.375 79.445 ;
        RECT 40.815 79.335 41.420 79.505 ;
        RECT 40.815 79.045 40.985 79.335 ;
        RECT 41.155 78.785 41.485 79.165 ;
        RECT 41.655 79.045 41.825 80.385 ;
        RECT 42.070 80.365 42.425 81.115 ;
        RECT 42.595 80.535 42.885 81.335 ;
        RECT 43.385 80.955 44.245 81.125 ;
        RECT 43.935 80.805 44.245 80.955 ;
        RECT 44.415 80.875 44.735 81.335 ;
        RECT 43.935 80.790 44.260 80.805 ;
        RECT 44.030 80.785 44.260 80.790 ;
        RECT 44.030 80.765 44.270 80.785 ;
        RECT 44.030 80.745 44.285 80.765 ;
        RECT 44.045 80.735 44.285 80.745 ;
        RECT 44.070 80.710 44.285 80.735 ;
        RECT 42.070 80.195 42.755 80.365 ;
        RECT 42.075 79.655 42.405 80.025 ;
        RECT 42.585 79.935 42.755 80.195 ;
        RECT 43.085 80.055 43.420 80.705 ;
        RECT 43.590 80.260 43.925 80.610 ;
        RECT 42.585 79.485 42.960 79.935 ;
        RECT 43.590 79.740 43.905 80.260 ;
        RECT 44.095 80.150 44.285 80.710 ;
        RECT 44.935 80.565 45.180 81.135 ;
        RECT 44.455 80.235 45.180 80.565 ;
        RECT 45.360 80.270 45.645 81.335 ;
        RECT 45.815 80.370 46.075 81.155 ;
        RECT 42.150 79.465 42.960 79.485 ;
        RECT 42.150 79.315 42.755 79.465 ;
        RECT 43.200 79.435 43.905 79.740 ;
        RECT 44.075 80.025 44.285 80.150 ;
        RECT 45.010 80.025 45.180 80.235 ;
        RECT 44.075 79.695 44.840 80.025 ;
        RECT 45.010 79.695 45.735 80.025 ;
        RECT 42.150 79.045 42.345 79.315 ;
        RECT 44.075 79.235 44.245 79.695 ;
        RECT 45.010 79.420 45.180 79.695 ;
        RECT 45.905 79.445 46.075 80.370 ;
        RECT 46.255 80.195 46.585 81.335 ;
        RECT 47.115 80.365 47.445 81.150 ;
        RECT 46.765 80.195 47.445 80.365 ;
        RECT 47.625 80.245 49.295 81.335 ;
        RECT 46.245 79.775 46.595 80.025 ;
        RECT 46.765 79.595 46.935 80.195 ;
        RECT 47.105 79.775 47.455 80.025 ;
        RECT 42.515 78.785 42.845 79.145 ;
        RECT 43.405 79.065 44.245 79.235 ;
        RECT 44.415 78.785 44.685 79.245 ;
        RECT 44.935 78.960 45.180 79.420 ;
        RECT 45.395 78.785 45.620 79.415 ;
        RECT 45.815 79.115 46.075 79.445 ;
        RECT 46.255 78.785 46.525 79.595 ;
        RECT 46.695 78.955 47.025 79.595 ;
        RECT 47.195 78.785 47.435 79.595 ;
        RECT 47.625 79.555 48.375 80.075 ;
        RECT 48.545 79.725 49.295 80.245 ;
        RECT 49.925 80.195 50.185 81.335 ;
        RECT 50.355 80.185 50.685 81.165 ;
        RECT 50.855 80.195 51.135 81.335 ;
        RECT 51.315 80.275 51.645 81.125 ;
        RECT 50.445 80.145 50.620 80.185 ;
        RECT 49.945 79.775 50.280 80.025 ;
        RECT 50.450 79.585 50.620 80.145 ;
        RECT 50.790 79.755 51.125 80.025 ;
        RECT 47.625 78.785 49.295 79.555 ;
        RECT 49.925 78.955 50.620 79.585 ;
        RECT 50.825 78.785 51.135 79.585 ;
        RECT 51.315 79.510 51.505 80.275 ;
        RECT 51.815 80.195 52.065 81.335 ;
        RECT 52.255 80.695 52.505 81.115 ;
        RECT 52.735 80.865 53.065 81.335 ;
        RECT 53.295 80.695 53.545 81.115 ;
        RECT 52.255 80.525 53.545 80.695 ;
        RECT 53.725 80.695 54.055 81.125 ;
        RECT 53.725 80.525 54.180 80.695 ;
        RECT 52.245 80.025 52.460 80.355 ;
        RECT 51.675 79.695 51.985 80.025 ;
        RECT 52.155 79.695 52.460 80.025 ;
        RECT 52.635 79.695 52.920 80.355 ;
        RECT 53.115 79.695 53.380 80.355 ;
        RECT 53.595 79.695 53.840 80.355 ;
        RECT 51.815 79.525 51.985 79.695 ;
        RECT 54.010 79.525 54.180 80.525 ;
        RECT 54.535 80.365 54.865 81.150 ;
        RECT 54.535 80.195 55.215 80.365 ;
        RECT 55.395 80.195 55.725 81.335 ;
        RECT 55.905 80.245 57.115 81.335 ;
        RECT 54.525 79.775 54.875 80.025 ;
        RECT 55.045 79.595 55.215 80.195 ;
        RECT 55.385 79.775 55.735 80.025 ;
        RECT 51.315 79.000 51.645 79.510 ;
        RECT 51.815 79.355 54.180 79.525 ;
        RECT 51.815 78.785 52.145 79.185 ;
        RECT 53.195 79.015 53.525 79.355 ;
        RECT 53.695 78.785 54.025 79.185 ;
        RECT 54.545 78.785 54.785 79.595 ;
        RECT 54.955 78.955 55.285 79.595 ;
        RECT 55.455 78.785 55.725 79.595 ;
        RECT 55.905 79.535 56.425 80.075 ;
        RECT 56.595 79.705 57.115 80.245 ;
        RECT 57.285 80.195 57.565 81.335 ;
        RECT 57.735 80.185 58.065 81.165 ;
        RECT 58.235 80.195 58.495 81.335 ;
        RECT 59.215 80.405 59.385 81.165 ;
        RECT 59.565 80.575 59.895 81.335 ;
        RECT 59.215 80.235 59.880 80.405 ;
        RECT 60.065 80.260 60.335 81.165 ;
        RECT 57.295 79.755 57.630 80.025 ;
        RECT 57.800 79.585 57.970 80.185 ;
        RECT 59.710 80.090 59.880 80.235 ;
        RECT 58.140 79.775 58.475 80.025 ;
        RECT 59.145 79.685 59.475 80.055 ;
        RECT 59.710 79.760 59.995 80.090 ;
        RECT 55.905 78.785 57.115 79.535 ;
        RECT 57.285 78.785 57.595 79.585 ;
        RECT 57.800 78.955 58.495 79.585 ;
        RECT 59.710 79.505 59.880 79.760 ;
        RECT 59.215 79.335 59.880 79.505 ;
        RECT 60.165 79.460 60.335 80.260 ;
        RECT 61.425 80.170 61.715 81.335 ;
        RECT 61.885 80.245 64.475 81.335 ;
        RECT 61.885 79.555 63.095 80.075 ;
        RECT 63.265 79.725 64.475 80.245 ;
        RECT 65.105 80.260 65.375 81.165 ;
        RECT 65.545 80.575 65.875 81.335 ;
        RECT 66.055 80.405 66.225 81.165 ;
        RECT 59.215 78.955 59.385 79.335 ;
        RECT 59.565 78.785 59.895 79.165 ;
        RECT 60.075 78.955 60.335 79.460 ;
        RECT 61.425 78.785 61.715 79.510 ;
        RECT 61.885 78.785 64.475 79.555 ;
        RECT 65.105 79.460 65.275 80.260 ;
        RECT 65.560 80.235 66.225 80.405 ;
        RECT 66.485 80.245 69.995 81.335 ;
        RECT 70.165 80.245 71.375 81.335 ;
        RECT 71.735 80.610 72.065 81.335 ;
        RECT 65.560 80.090 65.730 80.235 ;
        RECT 65.445 79.760 65.730 80.090 ;
        RECT 65.560 79.505 65.730 79.760 ;
        RECT 65.965 79.685 66.295 80.055 ;
        RECT 66.485 79.555 68.135 80.075 ;
        RECT 68.305 79.725 69.995 80.245 ;
        RECT 65.105 78.955 65.365 79.460 ;
        RECT 65.560 79.335 66.225 79.505 ;
        RECT 65.545 78.785 65.875 79.165 ;
        RECT 66.055 78.955 66.225 79.335 ;
        RECT 66.485 78.785 69.995 79.555 ;
        RECT 70.165 79.535 70.685 80.075 ;
        RECT 70.855 79.705 71.375 80.245 ;
        RECT 70.165 78.785 71.375 79.535 ;
        RECT 71.545 78.955 72.065 80.440 ;
        RECT 72.235 79.615 72.755 81.165 ;
        RECT 73.015 80.665 73.185 81.165 ;
        RECT 73.355 80.835 73.685 81.335 ;
        RECT 73.015 80.495 73.620 80.665 ;
        RECT 72.925 79.685 73.170 80.325 ;
        RECT 73.450 80.100 73.620 80.495 ;
        RECT 73.855 80.385 74.080 81.165 ;
        RECT 73.450 79.770 73.680 80.100 ;
        RECT 73.450 79.505 73.620 79.770 ;
        RECT 72.235 78.785 72.575 79.445 ;
        RECT 73.015 79.335 73.620 79.505 ;
        RECT 73.015 79.045 73.185 79.335 ;
        RECT 73.355 78.785 73.685 79.165 ;
        RECT 73.855 79.045 74.025 80.385 ;
        RECT 74.270 80.365 74.625 81.115 ;
        RECT 74.795 80.535 75.085 81.335 ;
        RECT 75.585 80.955 76.445 81.125 ;
        RECT 76.135 80.805 76.445 80.955 ;
        RECT 76.615 80.875 76.935 81.335 ;
        RECT 76.135 80.790 76.460 80.805 ;
        RECT 76.230 80.785 76.460 80.790 ;
        RECT 76.230 80.765 76.470 80.785 ;
        RECT 76.230 80.745 76.485 80.765 ;
        RECT 76.245 80.735 76.485 80.745 ;
        RECT 76.270 80.710 76.485 80.735 ;
        RECT 74.270 80.195 74.955 80.365 ;
        RECT 74.275 79.655 74.605 80.025 ;
        RECT 74.785 79.935 74.955 80.195 ;
        RECT 75.285 80.055 75.620 80.705 ;
        RECT 75.790 80.260 76.125 80.610 ;
        RECT 74.785 79.485 75.160 79.935 ;
        RECT 75.790 79.740 76.105 80.260 ;
        RECT 76.295 80.150 76.485 80.710 ;
        RECT 77.135 80.565 77.380 81.135 ;
        RECT 76.655 80.235 77.380 80.565 ;
        RECT 77.560 80.270 77.845 81.335 ;
        RECT 78.015 80.370 78.275 81.155 ;
        RECT 74.350 79.465 75.160 79.485 ;
        RECT 74.350 79.315 74.955 79.465 ;
        RECT 75.400 79.435 76.105 79.740 ;
        RECT 76.275 80.025 76.485 80.150 ;
        RECT 77.210 80.025 77.380 80.235 ;
        RECT 76.275 79.695 77.040 80.025 ;
        RECT 77.210 79.695 77.935 80.025 ;
        RECT 74.350 79.045 74.545 79.315 ;
        RECT 76.275 79.235 76.445 79.695 ;
        RECT 77.210 79.420 77.380 79.695 ;
        RECT 78.105 79.445 78.275 80.370 ;
        RECT 79.550 80.365 79.940 80.540 ;
        RECT 80.425 80.535 80.755 81.335 ;
        RECT 80.925 80.545 81.460 81.165 ;
        RECT 79.550 80.195 80.975 80.365 ;
        RECT 79.425 79.465 79.780 80.025 ;
        RECT 74.715 78.785 75.045 79.145 ;
        RECT 75.605 79.065 76.445 79.235 ;
        RECT 76.615 78.785 76.885 79.245 ;
        RECT 77.135 78.960 77.380 79.420 ;
        RECT 77.595 78.785 77.820 79.415 ;
        RECT 78.015 79.115 78.275 79.445 ;
        RECT 79.950 79.295 80.120 80.195 ;
        RECT 80.290 79.465 80.555 80.025 ;
        RECT 80.805 79.695 80.975 80.195 ;
        RECT 81.145 79.525 81.460 80.545 ;
        RECT 81.755 80.665 81.925 81.165 ;
        RECT 82.095 80.835 82.425 81.335 ;
        RECT 81.755 80.495 82.360 80.665 ;
        RECT 81.665 79.685 81.910 80.325 ;
        RECT 82.190 80.100 82.360 80.495 ;
        RECT 82.595 80.385 82.820 81.165 ;
        RECT 82.190 79.770 82.420 80.100 ;
        RECT 79.530 78.785 79.770 79.295 ;
        RECT 79.950 78.965 80.230 79.295 ;
        RECT 80.460 78.785 80.675 79.295 ;
        RECT 80.845 78.955 81.460 79.525 ;
        RECT 82.190 79.505 82.360 79.770 ;
        RECT 81.755 79.335 82.360 79.505 ;
        RECT 81.755 79.045 81.925 79.335 ;
        RECT 82.095 78.785 82.425 79.165 ;
        RECT 82.595 79.045 82.765 80.385 ;
        RECT 83.010 80.365 83.365 81.115 ;
        RECT 83.535 80.535 83.825 81.335 ;
        RECT 84.325 80.955 85.185 81.125 ;
        RECT 84.875 80.805 85.185 80.955 ;
        RECT 85.355 80.875 85.675 81.335 ;
        RECT 84.875 80.790 85.200 80.805 ;
        RECT 84.970 80.785 85.200 80.790 ;
        RECT 84.970 80.765 85.210 80.785 ;
        RECT 84.970 80.745 85.225 80.765 ;
        RECT 84.985 80.735 85.225 80.745 ;
        RECT 85.010 80.710 85.225 80.735 ;
        RECT 83.010 80.195 83.695 80.365 ;
        RECT 83.015 79.655 83.345 80.025 ;
        RECT 83.525 79.935 83.695 80.195 ;
        RECT 84.025 80.055 84.360 80.705 ;
        RECT 84.530 80.260 84.865 80.610 ;
        RECT 83.525 79.485 83.900 79.935 ;
        RECT 84.530 79.740 84.845 80.260 ;
        RECT 85.035 80.150 85.225 80.710 ;
        RECT 85.875 80.565 86.120 81.135 ;
        RECT 85.395 80.235 86.120 80.565 ;
        RECT 86.300 80.270 86.585 81.335 ;
        RECT 86.755 80.370 87.015 81.155 ;
        RECT 83.090 79.465 83.900 79.485 ;
        RECT 83.090 79.315 83.695 79.465 ;
        RECT 84.140 79.435 84.845 79.740 ;
        RECT 85.015 80.025 85.225 80.150 ;
        RECT 85.950 80.025 86.120 80.235 ;
        RECT 85.015 79.695 85.780 80.025 ;
        RECT 85.950 79.695 86.675 80.025 ;
        RECT 83.090 79.045 83.285 79.315 ;
        RECT 85.015 79.235 85.185 79.695 ;
        RECT 85.950 79.420 86.120 79.695 ;
        RECT 86.845 79.445 87.015 80.370 ;
        RECT 87.185 80.170 87.475 81.335 ;
        RECT 87.735 80.665 87.905 81.165 ;
        RECT 88.075 80.835 88.405 81.335 ;
        RECT 87.735 80.495 88.340 80.665 ;
        RECT 87.645 79.685 87.890 80.325 ;
        RECT 88.170 80.100 88.340 80.495 ;
        RECT 88.575 80.385 88.800 81.165 ;
        RECT 88.170 79.770 88.400 80.100 ;
        RECT 83.455 78.785 83.785 79.145 ;
        RECT 84.345 79.065 85.185 79.235 ;
        RECT 85.355 78.785 85.625 79.245 ;
        RECT 85.875 78.960 86.120 79.420 ;
        RECT 86.335 78.785 86.560 79.415 ;
        RECT 86.755 79.115 87.015 79.445 ;
        RECT 87.185 78.785 87.475 79.510 ;
        RECT 88.170 79.505 88.340 79.770 ;
        RECT 87.735 79.335 88.340 79.505 ;
        RECT 87.735 79.045 87.905 79.335 ;
        RECT 88.075 78.785 88.405 79.165 ;
        RECT 88.575 79.045 88.745 80.385 ;
        RECT 88.990 80.365 89.345 81.115 ;
        RECT 89.515 80.535 89.805 81.335 ;
        RECT 90.305 80.955 91.165 81.125 ;
        RECT 90.855 80.805 91.165 80.955 ;
        RECT 91.335 80.875 91.655 81.335 ;
        RECT 90.855 80.790 91.180 80.805 ;
        RECT 90.950 80.785 91.180 80.790 ;
        RECT 90.950 80.765 91.190 80.785 ;
        RECT 90.950 80.745 91.205 80.765 ;
        RECT 90.965 80.735 91.205 80.745 ;
        RECT 90.990 80.710 91.205 80.735 ;
        RECT 88.990 80.195 89.675 80.365 ;
        RECT 88.995 79.655 89.325 80.025 ;
        RECT 89.505 79.935 89.675 80.195 ;
        RECT 90.005 80.055 90.340 80.705 ;
        RECT 90.510 80.260 90.845 80.610 ;
        RECT 89.505 79.485 89.880 79.935 ;
        RECT 90.510 79.740 90.825 80.260 ;
        RECT 91.015 80.150 91.205 80.710 ;
        RECT 91.855 80.565 92.100 81.135 ;
        RECT 91.375 80.235 92.100 80.565 ;
        RECT 92.280 80.270 92.565 81.335 ;
        RECT 92.735 80.370 92.995 81.155 ;
        RECT 89.070 79.465 89.880 79.485 ;
        RECT 89.070 79.315 89.675 79.465 ;
        RECT 90.120 79.435 90.825 79.740 ;
        RECT 90.995 80.025 91.205 80.150 ;
        RECT 91.930 80.025 92.100 80.235 ;
        RECT 90.995 79.695 91.760 80.025 ;
        RECT 91.930 79.695 92.655 80.025 ;
        RECT 89.070 79.045 89.265 79.315 ;
        RECT 90.995 79.235 91.165 79.695 ;
        RECT 91.930 79.420 92.100 79.695 ;
        RECT 92.825 79.445 92.995 80.370 ;
        RECT 93.165 80.245 94.835 81.335 ;
        RECT 95.465 80.780 96.070 81.335 ;
        RECT 96.245 80.825 96.725 81.165 ;
        RECT 96.895 80.790 97.150 81.335 ;
        RECT 95.465 80.680 96.080 80.780 ;
        RECT 95.895 80.655 96.080 80.680 ;
        RECT 89.435 78.785 89.765 79.145 ;
        RECT 90.325 79.065 91.165 79.235 ;
        RECT 91.335 78.785 91.605 79.245 ;
        RECT 91.855 78.960 92.100 79.420 ;
        RECT 92.315 78.785 92.540 79.415 ;
        RECT 92.735 79.115 92.995 79.445 ;
        RECT 93.165 79.555 93.915 80.075 ;
        RECT 94.085 79.725 94.835 80.245 ;
        RECT 95.465 80.060 95.725 80.510 ;
        RECT 95.895 80.410 96.225 80.655 ;
        RECT 96.395 80.335 97.150 80.585 ;
        RECT 97.320 80.465 97.595 81.165 ;
        RECT 96.380 80.300 97.150 80.335 ;
        RECT 96.365 80.290 97.150 80.300 ;
        RECT 96.360 80.275 97.255 80.290 ;
        RECT 96.340 80.260 97.255 80.275 ;
        RECT 96.320 80.250 97.255 80.260 ;
        RECT 96.295 80.240 97.255 80.250 ;
        RECT 96.225 80.210 97.255 80.240 ;
        RECT 96.205 80.180 97.255 80.210 ;
        RECT 96.185 80.150 97.255 80.180 ;
        RECT 96.155 80.125 97.255 80.150 ;
        RECT 96.120 80.090 97.255 80.125 ;
        RECT 96.090 80.085 97.255 80.090 ;
        RECT 96.090 80.080 96.480 80.085 ;
        RECT 96.090 80.070 96.455 80.080 ;
        RECT 96.090 80.065 96.440 80.070 ;
        RECT 96.090 80.060 96.425 80.065 ;
        RECT 95.465 80.055 96.425 80.060 ;
        RECT 95.465 80.045 96.415 80.055 ;
        RECT 95.465 80.040 96.405 80.045 ;
        RECT 95.465 80.030 96.395 80.040 ;
        RECT 95.465 80.020 96.390 80.030 ;
        RECT 95.465 80.015 96.385 80.020 ;
        RECT 95.465 80.000 96.375 80.015 ;
        RECT 95.465 79.985 96.370 80.000 ;
        RECT 95.465 79.960 96.360 79.985 ;
        RECT 95.465 79.890 96.355 79.960 ;
        RECT 93.165 78.785 94.835 79.555 ;
        RECT 95.465 79.335 96.015 79.720 ;
        RECT 96.185 79.165 96.355 79.890 ;
        RECT 95.465 78.995 96.355 79.165 ;
        RECT 96.525 79.490 96.855 79.915 ;
        RECT 97.025 79.690 97.255 80.085 ;
        RECT 96.525 79.465 96.775 79.490 ;
        RECT 96.525 79.005 96.745 79.465 ;
        RECT 97.425 79.435 97.595 80.465 ;
        RECT 96.915 78.785 97.165 79.325 ;
        RECT 97.335 78.955 97.595 79.435 ;
        RECT 97.765 80.260 98.035 81.165 ;
        RECT 98.205 80.575 98.535 81.335 ;
        RECT 98.715 80.405 98.885 81.165 ;
        RECT 97.765 79.460 97.935 80.260 ;
        RECT 98.220 80.235 98.885 80.405 ;
        RECT 99.145 80.245 100.815 81.335 ;
        RECT 101.075 80.665 101.245 81.165 ;
        RECT 101.415 80.835 101.745 81.335 ;
        RECT 101.075 80.495 101.740 80.665 ;
        RECT 98.220 80.090 98.390 80.235 ;
        RECT 98.105 79.760 98.390 80.090 ;
        RECT 98.220 79.505 98.390 79.760 ;
        RECT 98.625 79.685 98.955 80.055 ;
        RECT 99.145 79.555 99.895 80.075 ;
        RECT 100.065 79.725 100.815 80.245 ;
        RECT 100.990 79.675 101.340 80.325 ;
        RECT 97.765 78.955 98.025 79.460 ;
        RECT 98.220 79.335 98.885 79.505 ;
        RECT 98.205 78.785 98.535 79.165 ;
        RECT 98.715 78.955 98.885 79.335 ;
        RECT 99.145 78.785 100.815 79.555 ;
        RECT 101.510 79.505 101.740 80.495 ;
        RECT 101.075 79.335 101.740 79.505 ;
        RECT 101.075 79.045 101.245 79.335 ;
        RECT 101.415 78.785 101.745 79.165 ;
        RECT 101.915 79.045 102.100 81.165 ;
        RECT 102.340 80.875 102.605 81.335 ;
        RECT 102.775 80.740 103.025 81.165 ;
        RECT 103.235 80.890 104.340 81.060 ;
        RECT 102.720 80.610 103.025 80.740 ;
        RECT 102.270 79.415 102.550 80.365 ;
        RECT 102.720 79.505 102.890 80.610 ;
        RECT 103.060 79.825 103.300 80.420 ;
        RECT 103.470 80.355 104.000 80.720 ;
        RECT 103.470 79.655 103.640 80.355 ;
        RECT 104.170 80.275 104.340 80.890 ;
        RECT 104.510 80.535 104.680 81.335 ;
        RECT 104.850 80.835 105.100 81.165 ;
        RECT 105.325 80.865 106.210 81.035 ;
        RECT 104.170 80.185 104.680 80.275 ;
        RECT 102.720 79.375 102.945 79.505 ;
        RECT 103.115 79.435 103.640 79.655 ;
        RECT 103.810 80.015 104.680 80.185 ;
        RECT 102.355 78.785 102.605 79.245 ;
        RECT 102.775 79.235 102.945 79.375 ;
        RECT 103.810 79.235 103.980 80.015 ;
        RECT 104.510 79.945 104.680 80.015 ;
        RECT 104.190 79.765 104.390 79.795 ;
        RECT 104.850 79.765 105.020 80.835 ;
        RECT 105.190 79.945 105.380 80.665 ;
        RECT 104.190 79.465 105.020 79.765 ;
        RECT 105.550 79.735 105.870 80.695 ;
        RECT 102.775 79.065 103.110 79.235 ;
        RECT 103.305 79.065 103.980 79.235 ;
        RECT 104.300 78.785 104.670 79.285 ;
        RECT 104.850 79.235 105.020 79.465 ;
        RECT 105.405 79.405 105.870 79.735 ;
        RECT 106.040 80.025 106.210 80.865 ;
        RECT 106.390 80.835 106.705 81.335 ;
        RECT 106.935 80.605 107.275 81.165 ;
        RECT 106.380 80.230 107.275 80.605 ;
        RECT 107.445 80.325 107.615 81.335 ;
        RECT 107.085 80.025 107.275 80.230 ;
        RECT 107.785 80.275 108.115 81.120 ;
        RECT 107.785 80.195 108.175 80.275 ;
        RECT 108.345 80.245 109.555 81.335 ;
        RECT 107.960 80.145 108.175 80.195 ;
        RECT 106.040 79.695 106.915 80.025 ;
        RECT 107.085 79.695 107.835 80.025 ;
        RECT 106.040 79.235 106.210 79.695 ;
        RECT 107.085 79.525 107.285 79.695 ;
        RECT 108.005 79.565 108.175 80.145 ;
        RECT 107.950 79.525 108.175 79.565 ;
        RECT 104.850 79.065 105.255 79.235 ;
        RECT 105.425 79.065 106.210 79.235 ;
        RECT 106.485 78.785 106.695 79.315 ;
        RECT 106.955 79.000 107.285 79.525 ;
        RECT 107.795 79.440 108.175 79.525 ;
        RECT 108.345 79.535 108.865 80.075 ;
        RECT 109.035 79.705 109.555 80.245 ;
        RECT 109.735 80.365 110.065 81.150 ;
        RECT 109.735 80.195 110.415 80.365 ;
        RECT 110.595 80.195 110.925 81.335 ;
        RECT 111.105 80.245 112.775 81.335 ;
        RECT 109.725 79.775 110.075 80.025 ;
        RECT 110.245 79.595 110.415 80.195 ;
        RECT 110.585 79.775 110.935 80.025 ;
        RECT 107.455 78.785 107.625 79.395 ;
        RECT 107.795 79.005 108.125 79.440 ;
        RECT 108.345 78.785 109.555 79.535 ;
        RECT 109.745 78.785 109.985 79.595 ;
        RECT 110.155 78.955 110.485 79.595 ;
        RECT 110.655 78.785 110.925 79.595 ;
        RECT 111.105 79.555 111.855 80.075 ;
        RECT 112.025 79.725 112.775 80.245 ;
        RECT 112.945 80.170 113.235 81.335 ;
        RECT 114.415 80.665 114.585 81.165 ;
        RECT 114.755 80.835 115.085 81.335 ;
        RECT 114.415 80.495 115.020 80.665 ;
        RECT 114.325 79.685 114.570 80.325 ;
        RECT 114.850 80.100 115.020 80.495 ;
        RECT 115.255 80.385 115.480 81.165 ;
        RECT 114.850 79.770 115.080 80.100 ;
        RECT 111.105 78.785 112.775 79.555 ;
        RECT 112.945 78.785 113.235 79.510 ;
        RECT 114.850 79.505 115.020 79.770 ;
        RECT 114.415 79.335 115.020 79.505 ;
        RECT 114.415 79.045 114.585 79.335 ;
        RECT 114.755 78.785 115.085 79.165 ;
        RECT 115.255 79.045 115.425 80.385 ;
        RECT 115.670 80.365 116.025 81.115 ;
        RECT 116.195 80.535 116.485 81.335 ;
        RECT 116.985 80.955 117.845 81.125 ;
        RECT 117.535 80.805 117.845 80.955 ;
        RECT 118.015 80.875 118.335 81.335 ;
        RECT 117.535 80.790 117.860 80.805 ;
        RECT 117.630 80.785 117.860 80.790 ;
        RECT 117.630 80.765 117.870 80.785 ;
        RECT 117.630 80.745 117.885 80.765 ;
        RECT 117.645 80.735 117.885 80.745 ;
        RECT 117.670 80.710 117.885 80.735 ;
        RECT 115.670 80.195 116.355 80.365 ;
        RECT 115.675 79.655 116.005 80.025 ;
        RECT 116.185 79.935 116.355 80.195 ;
        RECT 116.685 80.055 117.020 80.705 ;
        RECT 117.190 80.260 117.525 80.610 ;
        RECT 116.185 79.485 116.560 79.935 ;
        RECT 117.190 79.740 117.505 80.260 ;
        RECT 117.695 80.150 117.885 80.710 ;
        RECT 118.535 80.565 118.780 81.135 ;
        RECT 118.055 80.235 118.780 80.565 ;
        RECT 118.960 80.270 119.245 81.335 ;
        RECT 119.415 80.370 119.675 81.155 ;
        RECT 115.750 79.465 116.560 79.485 ;
        RECT 115.750 79.315 116.355 79.465 ;
        RECT 116.800 79.435 117.505 79.740 ;
        RECT 117.675 80.025 117.885 80.150 ;
        RECT 118.610 80.025 118.780 80.235 ;
        RECT 117.675 79.695 118.440 80.025 ;
        RECT 118.610 79.695 119.335 80.025 ;
        RECT 115.750 79.045 115.945 79.315 ;
        RECT 117.675 79.235 117.845 79.695 ;
        RECT 118.610 79.420 118.780 79.695 ;
        RECT 119.505 79.445 119.675 80.370 ;
        RECT 119.845 79.615 120.365 81.165 ;
        RECT 120.535 80.610 120.865 81.335 ;
        RECT 121.315 80.665 121.485 81.165 ;
        RECT 121.655 80.835 121.985 81.335 ;
        RECT 121.315 80.495 121.980 80.665 ;
        RECT 116.115 78.785 116.445 79.145 ;
        RECT 117.005 79.065 117.845 79.235 ;
        RECT 118.015 78.785 118.285 79.245 ;
        RECT 118.535 78.960 118.780 79.420 ;
        RECT 118.995 78.785 119.220 79.415 ;
        RECT 119.415 79.115 119.675 79.445 ;
        RECT 120.025 78.785 120.365 79.445 ;
        RECT 120.535 78.955 121.055 80.440 ;
        RECT 121.230 79.675 121.580 80.325 ;
        RECT 121.750 79.505 121.980 80.495 ;
        RECT 121.315 79.335 121.980 79.505 ;
        RECT 121.315 79.045 121.485 79.335 ;
        RECT 121.655 78.785 121.985 79.165 ;
        RECT 122.155 79.045 122.340 81.165 ;
        RECT 122.580 80.875 122.845 81.335 ;
        RECT 123.015 80.740 123.265 81.165 ;
        RECT 123.475 80.890 124.580 81.060 ;
        RECT 122.960 80.610 123.265 80.740 ;
        RECT 122.510 79.415 122.790 80.365 ;
        RECT 122.960 79.505 123.130 80.610 ;
        RECT 123.300 79.825 123.540 80.420 ;
        RECT 123.710 80.355 124.240 80.720 ;
        RECT 123.710 79.655 123.880 80.355 ;
        RECT 124.410 80.275 124.580 80.890 ;
        RECT 124.750 80.535 124.920 81.335 ;
        RECT 125.090 80.835 125.340 81.165 ;
        RECT 125.565 80.865 126.450 81.035 ;
        RECT 124.410 80.185 124.920 80.275 ;
        RECT 122.960 79.375 123.185 79.505 ;
        RECT 123.355 79.435 123.880 79.655 ;
        RECT 124.050 80.015 124.920 80.185 ;
        RECT 122.595 78.785 122.845 79.245 ;
        RECT 123.015 79.235 123.185 79.375 ;
        RECT 124.050 79.235 124.220 80.015 ;
        RECT 124.750 79.945 124.920 80.015 ;
        RECT 124.430 79.765 124.630 79.795 ;
        RECT 125.090 79.765 125.260 80.835 ;
        RECT 125.430 79.945 125.620 80.665 ;
        RECT 124.430 79.465 125.260 79.765 ;
        RECT 125.790 79.735 126.110 80.695 ;
        RECT 123.015 79.065 123.350 79.235 ;
        RECT 123.545 79.065 124.220 79.235 ;
        RECT 124.540 78.785 124.910 79.285 ;
        RECT 125.090 79.235 125.260 79.465 ;
        RECT 125.645 79.405 126.110 79.735 ;
        RECT 126.280 80.025 126.450 80.865 ;
        RECT 126.630 80.835 126.945 81.335 ;
        RECT 127.175 80.605 127.515 81.165 ;
        RECT 126.620 80.230 127.515 80.605 ;
        RECT 127.685 80.325 127.855 81.335 ;
        RECT 127.325 80.025 127.515 80.230 ;
        RECT 128.025 80.275 128.355 81.120 ;
        RECT 128.025 80.195 128.415 80.275 ;
        RECT 128.585 80.195 128.865 81.335 ;
        RECT 128.200 80.145 128.415 80.195 ;
        RECT 129.035 80.185 129.365 81.165 ;
        RECT 129.535 80.195 129.795 81.335 ;
        RECT 126.280 79.695 127.155 80.025 ;
        RECT 127.325 79.695 128.075 80.025 ;
        RECT 126.280 79.235 126.450 79.695 ;
        RECT 127.325 79.525 127.525 79.695 ;
        RECT 128.245 79.565 128.415 80.145 ;
        RECT 128.595 79.755 128.930 80.025 ;
        RECT 129.100 79.585 129.270 80.185 ;
        RECT 129.440 79.775 129.775 80.025 ;
        RECT 130.885 79.615 131.405 81.165 ;
        RECT 131.575 80.610 131.905 81.335 ;
        RECT 132.815 80.665 132.985 81.165 ;
        RECT 133.155 80.835 133.485 81.335 ;
        RECT 132.815 80.495 133.420 80.665 ;
        RECT 128.190 79.525 128.415 79.565 ;
        RECT 125.090 79.065 125.495 79.235 ;
        RECT 125.665 79.065 126.450 79.235 ;
        RECT 126.725 78.785 126.935 79.315 ;
        RECT 127.195 79.000 127.525 79.525 ;
        RECT 128.035 79.440 128.415 79.525 ;
        RECT 127.695 78.785 127.865 79.395 ;
        RECT 128.035 79.005 128.365 79.440 ;
        RECT 128.585 78.785 128.895 79.585 ;
        RECT 129.100 78.955 129.795 79.585 ;
        RECT 131.065 78.785 131.405 79.445 ;
        RECT 131.575 78.955 132.095 80.440 ;
        RECT 132.725 79.685 132.970 80.325 ;
        RECT 133.250 80.100 133.420 80.495 ;
        RECT 133.655 80.385 133.880 81.165 ;
        RECT 133.250 79.770 133.480 80.100 ;
        RECT 133.250 79.505 133.420 79.770 ;
        RECT 132.815 79.335 133.420 79.505 ;
        RECT 132.815 79.045 132.985 79.335 ;
        RECT 133.155 78.785 133.485 79.165 ;
        RECT 133.655 79.045 133.825 80.385 ;
        RECT 134.070 80.365 134.425 81.115 ;
        RECT 134.595 80.535 134.885 81.335 ;
        RECT 135.385 80.955 136.245 81.125 ;
        RECT 135.935 80.805 136.245 80.955 ;
        RECT 136.415 80.875 136.735 81.335 ;
        RECT 135.935 80.790 136.260 80.805 ;
        RECT 136.030 80.785 136.260 80.790 ;
        RECT 136.030 80.765 136.270 80.785 ;
        RECT 136.030 80.745 136.285 80.765 ;
        RECT 136.045 80.735 136.285 80.745 ;
        RECT 136.070 80.710 136.285 80.735 ;
        RECT 134.070 80.195 134.755 80.365 ;
        RECT 134.075 79.655 134.405 80.025 ;
        RECT 134.585 79.935 134.755 80.195 ;
        RECT 135.085 80.055 135.420 80.705 ;
        RECT 135.590 80.260 135.925 80.610 ;
        RECT 134.585 79.485 134.960 79.935 ;
        RECT 135.590 79.740 135.905 80.260 ;
        RECT 136.095 80.150 136.285 80.710 ;
        RECT 136.935 80.565 137.180 81.135 ;
        RECT 136.455 80.235 137.180 80.565 ;
        RECT 137.360 80.270 137.645 81.335 ;
        RECT 137.815 80.370 138.075 81.155 ;
        RECT 134.150 79.465 134.960 79.485 ;
        RECT 134.150 79.315 134.755 79.465 ;
        RECT 135.200 79.435 135.905 79.740 ;
        RECT 136.075 80.025 136.285 80.150 ;
        RECT 137.010 80.025 137.180 80.235 ;
        RECT 136.075 79.695 136.840 80.025 ;
        RECT 137.010 79.695 137.735 80.025 ;
        RECT 134.150 79.045 134.345 79.315 ;
        RECT 136.075 79.235 136.245 79.695 ;
        RECT 137.010 79.420 137.180 79.695 ;
        RECT 137.905 79.445 138.075 80.370 ;
        RECT 138.705 80.170 138.995 81.335 ;
        RECT 139.165 80.245 140.835 81.335 ;
        RECT 141.025 80.745 141.265 81.135 ;
        RECT 141.435 80.925 141.785 81.335 ;
        RECT 141.025 80.545 141.775 80.745 ;
        RECT 139.165 79.555 139.915 80.075 ;
        RECT 140.085 79.725 140.835 80.245 ;
        RECT 134.515 78.785 134.845 79.145 ;
        RECT 135.405 79.065 136.245 79.235 ;
        RECT 136.415 78.785 136.685 79.245 ;
        RECT 136.935 78.960 137.180 79.420 ;
        RECT 137.395 78.785 137.620 79.415 ;
        RECT 137.815 79.115 138.075 79.445 ;
        RECT 138.705 78.785 138.995 79.510 ;
        RECT 139.165 78.785 140.835 79.555 ;
        RECT 141.025 79.025 141.255 80.365 ;
        RECT 141.435 79.865 141.775 80.545 ;
        RECT 141.955 80.045 142.285 81.155 ;
        RECT 142.455 80.685 142.635 81.155 ;
        RECT 142.805 80.855 143.135 81.335 ;
        RECT 143.310 80.685 143.480 81.155 ;
        RECT 142.455 80.485 143.480 80.685 ;
        RECT 141.435 78.965 141.665 79.865 ;
        RECT 141.955 79.745 142.500 80.045 ;
        RECT 141.865 78.785 142.110 79.565 ;
        RECT 142.280 79.515 142.500 79.745 ;
        RECT 142.670 79.695 143.095 80.315 ;
        RECT 143.290 79.695 143.550 80.315 ;
        RECT 143.745 80.195 144.030 81.335 ;
        RECT 143.760 79.515 144.020 80.025 ;
        RECT 142.280 79.325 144.020 79.515 ;
        RECT 142.280 78.965 142.710 79.325 ;
        RECT 143.290 78.785 144.020 79.155 ;
        RECT 144.220 78.965 144.500 81.155 ;
        RECT 145.235 80.665 145.405 81.165 ;
        RECT 145.575 80.835 145.905 81.335 ;
        RECT 145.235 80.495 145.900 80.665 ;
        RECT 145.150 79.675 145.500 80.325 ;
        RECT 145.670 79.505 145.900 80.495 ;
        RECT 145.235 79.335 145.900 79.505 ;
        RECT 145.235 79.045 145.405 79.335 ;
        RECT 145.575 78.785 145.905 79.165 ;
        RECT 146.075 79.045 146.260 81.165 ;
        RECT 146.500 80.875 146.765 81.335 ;
        RECT 146.935 80.740 147.185 81.165 ;
        RECT 147.395 80.890 148.500 81.060 ;
        RECT 146.880 80.610 147.185 80.740 ;
        RECT 146.430 79.415 146.710 80.365 ;
        RECT 146.880 79.505 147.050 80.610 ;
        RECT 147.220 79.825 147.460 80.420 ;
        RECT 147.630 80.355 148.160 80.720 ;
        RECT 147.630 79.655 147.800 80.355 ;
        RECT 148.330 80.275 148.500 80.890 ;
        RECT 148.670 80.535 148.840 81.335 ;
        RECT 149.010 80.835 149.260 81.165 ;
        RECT 149.485 80.865 150.370 81.035 ;
        RECT 148.330 80.185 148.840 80.275 ;
        RECT 146.880 79.375 147.105 79.505 ;
        RECT 147.275 79.435 147.800 79.655 ;
        RECT 147.970 80.015 148.840 80.185 ;
        RECT 146.515 78.785 146.765 79.245 ;
        RECT 146.935 79.235 147.105 79.375 ;
        RECT 147.970 79.235 148.140 80.015 ;
        RECT 148.670 79.945 148.840 80.015 ;
        RECT 148.350 79.765 148.550 79.795 ;
        RECT 149.010 79.765 149.180 80.835 ;
        RECT 149.350 79.945 149.540 80.665 ;
        RECT 148.350 79.465 149.180 79.765 ;
        RECT 149.710 79.735 150.030 80.695 ;
        RECT 146.935 79.065 147.270 79.235 ;
        RECT 147.465 79.065 148.140 79.235 ;
        RECT 148.460 78.785 148.830 79.285 ;
        RECT 149.010 79.235 149.180 79.465 ;
        RECT 149.565 79.405 150.030 79.735 ;
        RECT 150.200 80.025 150.370 80.865 ;
        RECT 150.550 80.835 150.865 81.335 ;
        RECT 151.095 80.605 151.435 81.165 ;
        RECT 150.540 80.230 151.435 80.605 ;
        RECT 151.605 80.325 151.775 81.335 ;
        RECT 151.245 80.025 151.435 80.230 ;
        RECT 151.945 80.275 152.275 81.120 ;
        RECT 151.945 80.195 152.335 80.275 ;
        RECT 152.505 80.245 155.095 81.335 ;
        RECT 152.120 80.145 152.335 80.195 ;
        RECT 150.200 79.695 151.075 80.025 ;
        RECT 151.245 79.695 151.995 80.025 ;
        RECT 150.200 79.235 150.370 79.695 ;
        RECT 151.245 79.525 151.445 79.695 ;
        RECT 152.165 79.565 152.335 80.145 ;
        RECT 152.110 79.525 152.335 79.565 ;
        RECT 149.010 79.065 149.415 79.235 ;
        RECT 149.585 79.065 150.370 79.235 ;
        RECT 150.645 78.785 150.855 79.315 ;
        RECT 151.115 79.000 151.445 79.525 ;
        RECT 151.955 79.440 152.335 79.525 ;
        RECT 152.505 79.555 153.715 80.075 ;
        RECT 153.885 79.725 155.095 80.245 ;
        RECT 155.725 80.245 156.935 81.335 ;
        RECT 155.725 79.705 156.245 80.245 ;
        RECT 151.615 78.785 151.785 79.395 ;
        RECT 151.955 79.005 152.285 79.440 ;
        RECT 152.505 78.785 155.095 79.555 ;
        RECT 156.415 79.535 156.935 80.075 ;
        RECT 155.725 78.785 156.935 79.535 ;
        RECT 22.700 78.615 157.020 78.785 ;
        RECT 22.785 77.865 23.995 78.615 ;
        RECT 24.165 77.865 25.375 78.615 ;
        RECT 25.635 78.065 25.805 78.355 ;
        RECT 25.975 78.235 26.305 78.615 ;
        RECT 25.635 77.895 26.240 78.065 ;
        RECT 22.785 77.325 23.305 77.865 ;
        RECT 23.475 77.155 23.995 77.695 ;
        RECT 24.165 77.325 24.685 77.865 ;
        RECT 24.855 77.155 25.375 77.695 ;
        RECT 22.785 76.065 23.995 77.155 ;
        RECT 24.165 76.065 25.375 77.155 ;
        RECT 25.545 77.075 25.790 77.715 ;
        RECT 26.070 77.630 26.240 77.895 ;
        RECT 26.070 77.300 26.300 77.630 ;
        RECT 26.070 76.905 26.240 77.300 ;
        RECT 25.635 76.735 26.240 76.905 ;
        RECT 26.475 77.015 26.645 78.355 ;
        RECT 26.970 78.085 27.165 78.355 ;
        RECT 27.335 78.255 27.665 78.615 ;
        RECT 28.225 78.165 29.065 78.335 ;
        RECT 26.970 77.935 27.575 78.085 ;
        RECT 26.970 77.915 27.780 77.935 ;
        RECT 26.895 77.375 27.225 77.745 ;
        RECT 27.405 77.465 27.780 77.915 ;
        RECT 28.020 77.660 28.725 77.965 ;
        RECT 27.405 77.205 27.575 77.465 ;
        RECT 26.890 77.035 27.575 77.205 ;
        RECT 25.635 76.235 25.805 76.735 ;
        RECT 25.975 76.065 26.305 76.565 ;
        RECT 26.475 76.235 26.700 77.015 ;
        RECT 26.890 76.285 27.245 77.035 ;
        RECT 27.415 76.065 27.705 76.865 ;
        RECT 27.905 76.695 28.240 77.345 ;
        RECT 28.410 77.140 28.725 77.660 ;
        RECT 28.895 77.705 29.065 78.165 ;
        RECT 29.235 78.155 29.505 78.615 ;
        RECT 29.755 77.980 30.000 78.440 ;
        RECT 30.215 77.985 30.440 78.615 ;
        RECT 29.830 77.705 30.000 77.980 ;
        RECT 30.635 77.955 30.895 78.285 ;
        RECT 28.895 77.375 29.660 77.705 ;
        RECT 29.830 77.375 30.555 77.705 ;
        RECT 28.895 77.250 29.105 77.375 ;
        RECT 28.410 76.790 28.745 77.140 ;
        RECT 28.915 76.690 29.105 77.250 ;
        RECT 29.830 77.165 30.000 77.375 ;
        RECT 29.275 76.835 30.000 77.165 ;
        RECT 28.890 76.665 29.105 76.690 ;
        RECT 28.865 76.655 29.105 76.665 ;
        RECT 28.850 76.635 29.105 76.655 ;
        RECT 28.850 76.615 29.090 76.635 ;
        RECT 28.850 76.610 29.080 76.615 ;
        RECT 28.755 76.595 29.080 76.610 ;
        RECT 28.755 76.445 29.065 76.595 ;
        RECT 28.205 76.275 29.065 76.445 ;
        RECT 29.235 76.065 29.555 76.525 ;
        RECT 29.755 76.265 30.000 76.835 ;
        RECT 30.180 76.065 30.465 77.130 ;
        RECT 30.725 77.030 30.895 77.955 ;
        RECT 31.065 77.865 32.275 78.615 ;
        RECT 31.065 77.325 31.585 77.865 ;
        RECT 31.755 77.155 32.275 77.695 ;
        RECT 30.635 76.245 30.895 77.030 ;
        RECT 31.065 76.065 32.275 77.155 ;
        RECT 32.445 76.960 32.965 78.445 ;
        RECT 33.135 77.955 33.475 78.615 ;
        RECT 34.745 77.815 35.440 78.445 ;
        RECT 35.645 77.815 35.955 78.615 ;
        RECT 36.125 78.070 41.470 78.615 ;
        RECT 32.635 76.065 32.965 76.790 ;
        RECT 33.135 76.235 33.655 77.785 ;
        RECT 34.765 77.375 35.100 77.625 ;
        RECT 35.270 77.215 35.440 77.815 ;
        RECT 35.610 77.375 35.945 77.645 ;
        RECT 37.710 77.240 38.050 78.070 ;
        RECT 41.645 77.845 43.315 78.615 ;
        RECT 43.575 78.065 43.745 78.445 ;
        RECT 43.925 78.235 44.255 78.615 ;
        RECT 43.575 77.895 44.240 78.065 ;
        RECT 44.435 77.940 44.695 78.445 ;
        RECT 34.745 76.065 35.005 77.205 ;
        RECT 35.175 76.235 35.505 77.215 ;
        RECT 35.675 76.065 35.955 77.205 ;
        RECT 39.530 76.500 39.880 77.750 ;
        RECT 41.645 77.325 42.395 77.845 ;
        RECT 42.565 77.155 43.315 77.675 ;
        RECT 43.505 77.345 43.835 77.715 ;
        RECT 44.070 77.640 44.240 77.895 ;
        RECT 44.070 77.310 44.355 77.640 ;
        RECT 44.070 77.165 44.240 77.310 ;
        RECT 36.125 76.065 41.470 76.500 ;
        RECT 41.645 76.065 43.315 77.155 ;
        RECT 43.575 76.995 44.240 77.165 ;
        RECT 44.525 77.140 44.695 77.940 ;
        RECT 43.575 76.235 43.745 76.995 ;
        RECT 43.925 76.065 44.255 76.825 ;
        RECT 44.425 76.235 44.695 77.140 ;
        RECT 44.865 77.940 45.125 78.445 ;
        RECT 45.305 78.235 45.635 78.615 ;
        RECT 45.815 78.065 45.985 78.445 ;
        RECT 44.865 77.140 45.035 77.940 ;
        RECT 45.320 77.895 45.985 78.065 ;
        RECT 45.320 77.640 45.490 77.895 ;
        RECT 46.245 77.845 47.915 78.615 ;
        RECT 48.545 77.890 48.835 78.615 ;
        RECT 49.005 77.965 49.265 78.445 ;
        RECT 49.435 78.155 49.765 78.615 ;
        RECT 49.955 77.975 50.155 78.395 ;
        RECT 45.205 77.310 45.490 77.640 ;
        RECT 45.725 77.345 46.055 77.715 ;
        RECT 46.245 77.325 46.995 77.845 ;
        RECT 45.320 77.165 45.490 77.310 ;
        RECT 44.865 76.235 45.135 77.140 ;
        RECT 45.320 76.995 45.985 77.165 ;
        RECT 47.165 77.155 47.915 77.675 ;
        RECT 45.305 76.065 45.635 76.825 ;
        RECT 45.815 76.235 45.985 76.995 ;
        RECT 46.245 76.065 47.915 77.155 ;
        RECT 48.545 76.065 48.835 77.230 ;
        RECT 49.005 76.935 49.175 77.965 ;
        RECT 49.345 77.275 49.575 77.705 ;
        RECT 49.745 77.455 50.155 77.975 ;
        RECT 50.325 78.130 51.115 78.395 ;
        RECT 50.325 77.275 50.580 78.130 ;
        RECT 51.295 77.795 51.625 78.215 ;
        RECT 51.795 77.795 52.055 78.615 ;
        RECT 52.390 78.105 52.630 78.615 ;
        RECT 52.810 78.105 53.090 78.435 ;
        RECT 53.320 78.105 53.535 78.615 ;
        RECT 51.295 77.705 51.545 77.795 ;
        RECT 50.750 77.455 51.545 77.705 ;
        RECT 49.345 77.105 51.135 77.275 ;
        RECT 49.005 76.235 49.280 76.935 ;
        RECT 49.450 76.810 50.165 77.105 ;
        RECT 50.385 76.745 50.715 76.935 ;
        RECT 49.490 76.065 49.705 76.610 ;
        RECT 49.875 76.235 50.350 76.575 ;
        RECT 50.520 76.570 50.715 76.745 ;
        RECT 50.885 76.740 51.135 77.105 ;
        RECT 50.520 76.065 51.135 76.570 ;
        RECT 51.375 76.235 51.545 77.455 ;
        RECT 51.715 76.745 52.055 77.625 ;
        RECT 52.285 77.375 52.640 77.935 ;
        RECT 52.810 77.205 52.980 78.105 ;
        RECT 53.150 77.375 53.415 77.935 ;
        RECT 53.705 77.875 54.320 78.445 ;
        RECT 54.530 78.215 54.865 78.615 ;
        RECT 55.035 78.045 55.240 78.445 ;
        RECT 55.450 78.135 55.725 78.615 ;
        RECT 55.935 78.115 56.195 78.445 ;
        RECT 53.665 77.205 53.835 77.705 ;
        RECT 52.410 77.035 53.835 77.205 ;
        RECT 52.410 76.860 52.800 77.035 ;
        RECT 51.795 76.065 52.055 76.575 ;
        RECT 53.285 76.065 53.615 76.865 ;
        RECT 54.005 76.855 54.320 77.875 ;
        RECT 53.785 76.235 54.320 76.855 ;
        RECT 54.555 77.875 55.240 78.045 ;
        RECT 54.555 76.845 54.895 77.875 ;
        RECT 55.065 77.205 55.315 77.705 ;
        RECT 55.495 77.375 55.855 77.955 ;
        RECT 56.025 77.205 56.195 78.115 ;
        RECT 56.915 78.065 57.085 78.355 ;
        RECT 57.255 78.235 57.585 78.615 ;
        RECT 56.915 77.895 57.520 78.065 ;
        RECT 55.065 77.035 56.195 77.205 ;
        RECT 56.825 77.075 57.070 77.715 ;
        RECT 57.350 77.630 57.520 77.895 ;
        RECT 57.350 77.300 57.580 77.630 ;
        RECT 54.555 76.670 55.220 76.845 ;
        RECT 54.530 76.065 54.865 76.490 ;
        RECT 55.035 76.265 55.220 76.670 ;
        RECT 55.425 76.065 55.755 76.845 ;
        RECT 55.925 76.265 56.195 77.035 ;
        RECT 57.350 76.905 57.520 77.300 ;
        RECT 56.915 76.735 57.520 76.905 ;
        RECT 57.755 77.015 57.925 78.355 ;
        RECT 58.250 78.085 58.445 78.355 ;
        RECT 58.615 78.255 58.945 78.615 ;
        RECT 59.505 78.165 60.345 78.335 ;
        RECT 58.250 77.935 58.855 78.085 ;
        RECT 58.250 77.915 59.060 77.935 ;
        RECT 58.175 77.375 58.505 77.745 ;
        RECT 58.685 77.465 59.060 77.915 ;
        RECT 59.300 77.660 60.005 77.965 ;
        RECT 58.685 77.205 58.855 77.465 ;
        RECT 58.170 77.035 58.855 77.205 ;
        RECT 56.915 76.235 57.085 76.735 ;
        RECT 57.255 76.065 57.585 76.565 ;
        RECT 57.755 76.235 57.980 77.015 ;
        RECT 58.170 76.285 58.525 77.035 ;
        RECT 58.695 76.065 58.985 76.865 ;
        RECT 59.185 76.695 59.520 77.345 ;
        RECT 59.690 77.140 60.005 77.660 ;
        RECT 60.175 77.705 60.345 78.165 ;
        RECT 60.515 78.155 60.785 78.615 ;
        RECT 61.035 77.980 61.280 78.440 ;
        RECT 61.495 77.985 61.720 78.615 ;
        RECT 61.110 77.705 61.280 77.980 ;
        RECT 61.915 77.955 62.175 78.285 ;
        RECT 62.525 77.955 62.865 78.615 ;
        RECT 60.175 77.375 60.940 77.705 ;
        RECT 61.110 77.375 61.835 77.705 ;
        RECT 60.175 77.250 60.385 77.375 ;
        RECT 59.690 76.790 60.025 77.140 ;
        RECT 60.195 76.690 60.385 77.250 ;
        RECT 61.110 77.165 61.280 77.375 ;
        RECT 60.555 76.835 61.280 77.165 ;
        RECT 60.170 76.665 60.385 76.690 ;
        RECT 60.145 76.655 60.385 76.665 ;
        RECT 60.130 76.635 60.385 76.655 ;
        RECT 60.130 76.615 60.370 76.635 ;
        RECT 60.130 76.610 60.360 76.615 ;
        RECT 60.035 76.595 60.360 76.610 ;
        RECT 60.035 76.445 60.345 76.595 ;
        RECT 59.485 76.275 60.345 76.445 ;
        RECT 60.515 76.065 60.835 76.525 ;
        RECT 61.035 76.265 61.280 76.835 ;
        RECT 61.460 76.065 61.745 77.130 ;
        RECT 62.005 77.030 62.175 77.955 ;
        RECT 61.915 76.245 62.175 77.030 ;
        RECT 62.345 76.235 62.865 77.785 ;
        RECT 63.035 76.960 63.555 78.445 ;
        RECT 63.725 77.845 66.315 78.615 ;
        RECT 67.125 77.955 67.465 78.615 ;
        RECT 63.725 77.325 64.935 77.845 ;
        RECT 65.105 77.155 66.315 77.675 ;
        RECT 63.035 76.065 63.365 76.790 ;
        RECT 63.725 76.065 66.315 77.155 ;
        RECT 66.945 76.235 67.465 77.785 ;
        RECT 67.635 76.960 68.155 78.445 ;
        RECT 68.505 77.955 68.845 78.615 ;
        RECT 67.635 76.065 67.965 76.790 ;
        RECT 68.325 76.235 68.845 77.785 ;
        RECT 69.015 76.960 69.535 78.445 ;
        RECT 69.705 77.845 72.295 78.615 ;
        RECT 73.015 78.065 73.185 78.445 ;
        RECT 73.365 78.235 73.695 78.615 ;
        RECT 73.015 77.895 73.680 78.065 ;
        RECT 73.875 77.940 74.135 78.445 ;
        RECT 69.705 77.325 70.915 77.845 ;
        RECT 71.085 77.155 72.295 77.675 ;
        RECT 72.945 77.345 73.275 77.715 ;
        RECT 73.510 77.640 73.680 77.895 ;
        RECT 73.510 77.310 73.795 77.640 ;
        RECT 73.510 77.165 73.680 77.310 ;
        RECT 69.015 76.065 69.345 76.790 ;
        RECT 69.705 76.065 72.295 77.155 ;
        RECT 73.015 76.995 73.680 77.165 ;
        RECT 73.965 77.140 74.135 77.940 ;
        RECT 74.305 77.890 74.595 78.615 ;
        RECT 75.225 77.815 75.535 78.615 ;
        RECT 75.740 77.815 76.435 78.445 ;
        RECT 75.235 77.375 75.570 77.645 ;
        RECT 73.015 76.235 73.185 76.995 ;
        RECT 73.365 76.065 73.695 76.825 ;
        RECT 73.865 76.235 74.135 77.140 ;
        RECT 74.305 76.065 74.595 77.230 ;
        RECT 75.740 77.215 75.910 77.815 ;
        RECT 76.625 77.805 76.865 78.615 ;
        RECT 77.035 77.805 77.365 78.445 ;
        RECT 77.535 77.805 77.805 78.615 ;
        RECT 78.315 78.215 78.645 78.615 ;
        RECT 78.815 78.045 79.145 78.385 ;
        RECT 80.195 78.215 80.525 78.615 ;
        RECT 78.160 77.875 80.525 78.045 ;
        RECT 80.695 77.890 81.025 78.400 ;
        RECT 76.080 77.375 76.415 77.625 ;
        RECT 76.605 77.375 76.955 77.625 ;
        RECT 75.225 76.065 75.505 77.205 ;
        RECT 75.675 76.235 76.005 77.215 ;
        RECT 77.125 77.205 77.295 77.805 ;
        RECT 77.465 77.375 77.815 77.625 ;
        RECT 76.175 76.065 76.435 77.205 ;
        RECT 76.615 77.035 77.295 77.205 ;
        RECT 76.615 76.250 76.945 77.035 ;
        RECT 77.475 76.065 77.805 77.205 ;
        RECT 78.160 76.875 78.330 77.875 ;
        RECT 80.355 77.705 80.525 77.875 ;
        RECT 78.500 77.045 78.745 77.705 ;
        RECT 78.960 77.045 79.225 77.705 ;
        RECT 79.420 77.045 79.705 77.705 ;
        RECT 79.880 77.375 80.185 77.705 ;
        RECT 80.355 77.375 80.665 77.705 ;
        RECT 79.880 77.045 80.095 77.375 ;
        RECT 78.160 76.705 78.615 76.875 ;
        RECT 78.285 76.275 78.615 76.705 ;
        RECT 78.795 76.705 80.085 76.875 ;
        RECT 78.795 76.285 79.045 76.705 ;
        RECT 79.275 76.065 79.605 76.535 ;
        RECT 79.835 76.285 80.085 76.705 ;
        RECT 80.275 76.065 80.525 77.205 ;
        RECT 80.835 77.125 81.025 77.890 ;
        RECT 80.695 76.275 81.025 77.125 ;
        RECT 81.205 78.115 81.465 78.445 ;
        RECT 81.675 78.135 81.950 78.615 ;
        RECT 81.205 77.205 81.375 78.115 ;
        RECT 82.160 78.045 82.365 78.445 ;
        RECT 82.535 78.215 82.870 78.615 ;
        RECT 83.045 78.115 83.305 78.445 ;
        RECT 83.515 78.135 83.790 78.615 ;
        RECT 81.545 77.375 81.905 77.955 ;
        RECT 82.160 77.875 82.845 78.045 ;
        RECT 82.085 77.205 82.335 77.705 ;
        RECT 81.205 77.035 82.335 77.205 ;
        RECT 81.205 76.265 81.475 77.035 ;
        RECT 82.505 76.845 82.845 77.875 ;
        RECT 81.645 76.065 81.975 76.845 ;
        RECT 82.180 76.670 82.845 76.845 ;
        RECT 83.045 77.205 83.215 78.115 ;
        RECT 84.000 78.045 84.205 78.445 ;
        RECT 84.375 78.215 84.710 78.615 ;
        RECT 85.895 78.065 86.065 78.445 ;
        RECT 86.245 78.235 86.575 78.615 ;
        RECT 83.385 77.375 83.745 77.955 ;
        RECT 84.000 77.875 84.685 78.045 ;
        RECT 85.895 77.895 86.560 78.065 ;
        RECT 86.755 77.940 87.015 78.445 ;
        RECT 87.365 77.955 87.705 78.615 ;
        RECT 83.925 77.205 84.175 77.705 ;
        RECT 83.045 77.035 84.175 77.205 ;
        RECT 82.180 76.265 82.365 76.670 ;
        RECT 82.535 76.065 82.870 76.490 ;
        RECT 83.045 76.265 83.315 77.035 ;
        RECT 84.345 76.845 84.685 77.875 ;
        RECT 85.825 77.345 86.155 77.715 ;
        RECT 86.390 77.640 86.560 77.895 ;
        RECT 86.390 77.310 86.675 77.640 ;
        RECT 86.390 77.165 86.560 77.310 ;
        RECT 83.485 76.065 83.815 76.845 ;
        RECT 84.020 76.670 84.685 76.845 ;
        RECT 85.895 76.995 86.560 77.165 ;
        RECT 86.845 77.140 87.015 77.940 ;
        RECT 84.020 76.265 84.205 76.670 ;
        RECT 84.375 76.065 84.710 76.490 ;
        RECT 85.895 76.235 86.065 76.995 ;
        RECT 86.245 76.065 86.575 76.825 ;
        RECT 86.745 76.235 87.015 77.140 ;
        RECT 87.185 76.235 87.705 77.785 ;
        RECT 87.875 76.960 88.395 78.445 ;
        RECT 89.485 76.960 90.005 78.445 ;
        RECT 90.175 77.955 90.515 78.615 ;
        RECT 90.955 78.065 91.125 78.355 ;
        RECT 91.295 78.235 91.625 78.615 ;
        RECT 90.955 77.895 91.560 78.065 ;
        RECT 87.875 76.065 88.205 76.790 ;
        RECT 89.675 76.065 90.005 76.790 ;
        RECT 90.175 76.235 90.695 77.785 ;
        RECT 90.865 77.075 91.110 77.715 ;
        RECT 91.390 77.630 91.560 77.895 ;
        RECT 91.390 77.300 91.620 77.630 ;
        RECT 91.390 76.905 91.560 77.300 ;
        RECT 90.955 76.735 91.560 76.905 ;
        RECT 91.795 77.015 91.965 78.355 ;
        RECT 92.290 78.085 92.485 78.355 ;
        RECT 92.655 78.255 92.985 78.615 ;
        RECT 93.545 78.165 94.385 78.335 ;
        RECT 92.290 77.935 92.895 78.085 ;
        RECT 92.290 77.915 93.100 77.935 ;
        RECT 92.215 77.375 92.545 77.745 ;
        RECT 92.725 77.465 93.100 77.915 ;
        RECT 93.340 77.660 94.045 77.965 ;
        RECT 92.725 77.205 92.895 77.465 ;
        RECT 92.210 77.035 92.895 77.205 ;
        RECT 90.955 76.235 91.125 76.735 ;
        RECT 91.295 76.065 91.625 76.565 ;
        RECT 91.795 76.235 92.020 77.015 ;
        RECT 92.210 76.285 92.565 77.035 ;
        RECT 92.735 76.065 93.025 76.865 ;
        RECT 93.225 76.695 93.560 77.345 ;
        RECT 93.730 77.140 94.045 77.660 ;
        RECT 94.215 77.705 94.385 78.165 ;
        RECT 94.555 78.155 94.825 78.615 ;
        RECT 95.075 77.980 95.320 78.440 ;
        RECT 95.535 77.985 95.760 78.615 ;
        RECT 95.150 77.705 95.320 77.980 ;
        RECT 95.955 77.955 96.215 78.285 ;
        RECT 94.215 77.375 94.980 77.705 ;
        RECT 95.150 77.375 95.875 77.705 ;
        RECT 94.215 77.250 94.425 77.375 ;
        RECT 93.730 76.790 94.065 77.140 ;
        RECT 94.235 76.690 94.425 77.250 ;
        RECT 95.150 77.165 95.320 77.375 ;
        RECT 94.595 76.835 95.320 77.165 ;
        RECT 94.210 76.665 94.425 76.690 ;
        RECT 94.185 76.655 94.425 76.665 ;
        RECT 94.170 76.635 94.425 76.655 ;
        RECT 94.170 76.615 94.410 76.635 ;
        RECT 94.170 76.610 94.400 76.615 ;
        RECT 94.075 76.595 94.400 76.610 ;
        RECT 94.075 76.445 94.385 76.595 ;
        RECT 93.525 76.275 94.385 76.445 ;
        RECT 94.555 76.065 94.875 76.525 ;
        RECT 95.075 76.265 95.320 76.835 ;
        RECT 95.500 76.065 95.785 77.130 ;
        RECT 96.045 77.030 96.215 77.955 ;
        RECT 96.385 77.845 99.895 78.615 ;
        RECT 100.065 77.890 100.355 78.615 ;
        RECT 100.525 77.865 101.735 78.615 ;
        RECT 102.085 77.955 102.425 78.615 ;
        RECT 96.385 77.325 98.035 77.845 ;
        RECT 98.205 77.155 99.895 77.675 ;
        RECT 100.525 77.325 101.045 77.865 ;
        RECT 95.955 76.245 96.215 77.030 ;
        RECT 96.385 76.065 99.895 77.155 ;
        RECT 100.065 76.065 100.355 77.230 ;
        RECT 101.215 77.155 101.735 77.695 ;
        RECT 100.525 76.065 101.735 77.155 ;
        RECT 101.905 76.235 102.425 77.785 ;
        RECT 102.595 76.960 103.115 78.445 ;
        RECT 103.285 78.070 108.630 78.615 ;
        RECT 104.870 77.240 105.210 78.070 ;
        RECT 108.895 78.065 109.065 78.355 ;
        RECT 109.235 78.235 109.565 78.615 ;
        RECT 108.895 77.895 109.500 78.065 ;
        RECT 102.595 76.065 102.925 76.790 ;
        RECT 106.690 76.500 107.040 77.750 ;
        RECT 108.805 77.075 109.050 77.715 ;
        RECT 109.330 77.630 109.500 77.895 ;
        RECT 109.330 77.300 109.560 77.630 ;
        RECT 109.330 76.905 109.500 77.300 ;
        RECT 108.895 76.735 109.500 76.905 ;
        RECT 109.735 77.015 109.905 78.355 ;
        RECT 110.230 78.085 110.425 78.355 ;
        RECT 110.595 78.255 110.925 78.615 ;
        RECT 111.485 78.165 112.325 78.335 ;
        RECT 110.230 77.935 110.835 78.085 ;
        RECT 110.230 77.915 111.040 77.935 ;
        RECT 110.155 77.375 110.485 77.745 ;
        RECT 110.665 77.465 111.040 77.915 ;
        RECT 111.280 77.660 111.985 77.965 ;
        RECT 110.665 77.205 110.835 77.465 ;
        RECT 110.150 77.035 110.835 77.205 ;
        RECT 103.285 76.065 108.630 76.500 ;
        RECT 108.895 76.235 109.065 76.735 ;
        RECT 109.235 76.065 109.565 76.565 ;
        RECT 109.735 76.235 109.960 77.015 ;
        RECT 110.150 76.285 110.505 77.035 ;
        RECT 110.675 76.065 110.965 76.865 ;
        RECT 111.165 76.695 111.500 77.345 ;
        RECT 111.670 77.140 111.985 77.660 ;
        RECT 112.155 77.705 112.325 78.165 ;
        RECT 112.495 78.155 112.765 78.615 ;
        RECT 113.015 77.980 113.260 78.440 ;
        RECT 113.475 77.985 113.700 78.615 ;
        RECT 113.090 77.705 113.260 77.980 ;
        RECT 113.895 77.955 114.155 78.285 ;
        RECT 112.155 77.375 112.920 77.705 ;
        RECT 113.090 77.375 113.815 77.705 ;
        RECT 112.155 77.250 112.365 77.375 ;
        RECT 111.670 76.790 112.005 77.140 ;
        RECT 112.175 76.690 112.365 77.250 ;
        RECT 113.090 77.165 113.260 77.375 ;
        RECT 112.535 76.835 113.260 77.165 ;
        RECT 112.150 76.665 112.365 76.690 ;
        RECT 112.125 76.655 112.365 76.665 ;
        RECT 112.110 76.635 112.365 76.655 ;
        RECT 112.110 76.615 112.350 76.635 ;
        RECT 112.110 76.610 112.340 76.615 ;
        RECT 112.015 76.595 112.340 76.610 ;
        RECT 112.015 76.445 112.325 76.595 ;
        RECT 111.465 76.275 112.325 76.445 ;
        RECT 112.495 76.065 112.815 76.525 ;
        RECT 113.015 76.265 113.260 76.835 ;
        RECT 113.440 76.065 113.725 77.130 ;
        RECT 113.985 77.030 114.155 77.955 ;
        RECT 114.875 78.065 115.045 78.445 ;
        RECT 115.225 78.235 115.555 78.615 ;
        RECT 114.875 77.895 115.540 78.065 ;
        RECT 115.735 77.940 115.995 78.445 ;
        RECT 114.805 77.345 115.135 77.715 ;
        RECT 115.370 77.640 115.540 77.895 ;
        RECT 115.370 77.310 115.655 77.640 ;
        RECT 115.370 77.165 115.540 77.310 ;
        RECT 113.895 76.245 114.155 77.030 ;
        RECT 114.875 76.995 115.540 77.165 ;
        RECT 115.825 77.140 115.995 77.940 ;
        RECT 116.255 78.065 116.425 78.355 ;
        RECT 116.595 78.235 116.925 78.615 ;
        RECT 116.255 77.895 116.860 78.065 ;
        RECT 114.875 76.235 115.045 76.995 ;
        RECT 115.225 76.065 115.555 76.825 ;
        RECT 115.725 76.235 115.995 77.140 ;
        RECT 116.165 77.075 116.410 77.715 ;
        RECT 116.690 77.630 116.860 77.895 ;
        RECT 116.690 77.300 116.920 77.630 ;
        RECT 116.690 76.905 116.860 77.300 ;
        RECT 116.255 76.735 116.860 76.905 ;
        RECT 117.095 77.015 117.265 78.355 ;
        RECT 117.590 78.085 117.785 78.355 ;
        RECT 117.955 78.255 118.285 78.615 ;
        RECT 118.845 78.165 119.685 78.335 ;
        RECT 117.590 77.935 118.195 78.085 ;
        RECT 117.590 77.915 118.400 77.935 ;
        RECT 117.515 77.375 117.845 77.745 ;
        RECT 118.025 77.465 118.400 77.915 ;
        RECT 118.640 77.660 119.345 77.965 ;
        RECT 118.025 77.205 118.195 77.465 ;
        RECT 117.510 77.035 118.195 77.205 ;
        RECT 116.255 76.235 116.425 76.735 ;
        RECT 116.595 76.065 116.925 76.565 ;
        RECT 117.095 76.235 117.320 77.015 ;
        RECT 117.510 76.285 117.865 77.035 ;
        RECT 118.035 76.065 118.325 76.865 ;
        RECT 118.525 76.695 118.860 77.345 ;
        RECT 119.030 77.140 119.345 77.660 ;
        RECT 119.515 77.705 119.685 78.165 ;
        RECT 119.855 78.155 120.125 78.615 ;
        RECT 120.375 77.980 120.620 78.440 ;
        RECT 120.835 77.985 121.060 78.615 ;
        RECT 120.450 77.705 120.620 77.980 ;
        RECT 121.255 77.955 121.515 78.285 ;
        RECT 119.515 77.375 120.280 77.705 ;
        RECT 120.450 77.375 121.175 77.705 ;
        RECT 119.515 77.250 119.725 77.375 ;
        RECT 119.030 76.790 119.365 77.140 ;
        RECT 119.535 76.690 119.725 77.250 ;
        RECT 120.450 77.165 120.620 77.375 ;
        RECT 119.895 76.835 120.620 77.165 ;
        RECT 119.510 76.665 119.725 76.690 ;
        RECT 119.485 76.655 119.725 76.665 ;
        RECT 119.470 76.635 119.725 76.655 ;
        RECT 119.470 76.615 119.710 76.635 ;
        RECT 119.470 76.610 119.700 76.615 ;
        RECT 119.375 76.595 119.700 76.610 ;
        RECT 119.375 76.445 119.685 76.595 ;
        RECT 118.825 76.275 119.685 76.445 ;
        RECT 119.855 76.065 120.175 76.525 ;
        RECT 120.375 76.265 120.620 76.835 ;
        RECT 120.800 76.065 121.085 77.130 ;
        RECT 121.345 77.030 121.515 77.955 ;
        RECT 121.685 77.845 125.195 78.615 ;
        RECT 125.825 77.890 126.115 78.615 ;
        RECT 126.285 77.845 128.875 78.615 ;
        RECT 129.135 78.065 129.305 78.445 ;
        RECT 129.485 78.235 129.815 78.615 ;
        RECT 129.135 77.895 129.800 78.065 ;
        RECT 129.995 77.940 130.255 78.445 ;
        RECT 121.685 77.325 123.335 77.845 ;
        RECT 123.505 77.155 125.195 77.675 ;
        RECT 126.285 77.325 127.495 77.845 ;
        RECT 121.255 76.245 121.515 77.030 ;
        RECT 121.685 76.065 125.195 77.155 ;
        RECT 125.825 76.065 126.115 77.230 ;
        RECT 127.665 77.155 128.875 77.675 ;
        RECT 129.065 77.345 129.395 77.715 ;
        RECT 129.630 77.640 129.800 77.895 ;
        RECT 129.630 77.310 129.915 77.640 ;
        RECT 129.630 77.165 129.800 77.310 ;
        RECT 126.285 76.065 128.875 77.155 ;
        RECT 129.135 76.995 129.800 77.165 ;
        RECT 130.085 77.140 130.255 77.940 ;
        RECT 130.515 78.065 130.685 78.355 ;
        RECT 130.855 78.235 131.185 78.615 ;
        RECT 130.515 77.895 131.120 78.065 ;
        RECT 129.135 76.235 129.305 76.995 ;
        RECT 129.485 76.065 129.815 76.825 ;
        RECT 129.985 76.235 130.255 77.140 ;
        RECT 130.425 77.075 130.670 77.715 ;
        RECT 130.950 77.630 131.120 77.895 ;
        RECT 130.950 77.300 131.180 77.630 ;
        RECT 130.950 76.905 131.120 77.300 ;
        RECT 130.515 76.735 131.120 76.905 ;
        RECT 131.355 77.015 131.525 78.355 ;
        RECT 131.850 78.085 132.045 78.355 ;
        RECT 132.215 78.255 132.545 78.615 ;
        RECT 133.105 78.165 133.945 78.335 ;
        RECT 131.850 77.935 132.455 78.085 ;
        RECT 131.850 77.915 132.660 77.935 ;
        RECT 131.775 77.375 132.105 77.745 ;
        RECT 132.285 77.465 132.660 77.915 ;
        RECT 132.900 77.660 133.605 77.965 ;
        RECT 132.285 77.205 132.455 77.465 ;
        RECT 131.770 77.035 132.455 77.205 ;
        RECT 130.515 76.235 130.685 76.735 ;
        RECT 130.855 76.065 131.185 76.565 ;
        RECT 131.355 76.235 131.580 77.015 ;
        RECT 131.770 76.285 132.125 77.035 ;
        RECT 132.295 76.065 132.585 76.865 ;
        RECT 132.785 76.695 133.120 77.345 ;
        RECT 133.290 77.140 133.605 77.660 ;
        RECT 133.775 77.705 133.945 78.165 ;
        RECT 134.115 78.155 134.385 78.615 ;
        RECT 134.635 77.980 134.880 78.440 ;
        RECT 135.095 77.985 135.320 78.615 ;
        RECT 134.710 77.705 134.880 77.980 ;
        RECT 135.515 77.955 135.775 78.285 ;
        RECT 133.775 77.375 134.540 77.705 ;
        RECT 134.710 77.375 135.435 77.705 ;
        RECT 133.775 77.250 133.985 77.375 ;
        RECT 133.290 76.790 133.625 77.140 ;
        RECT 133.795 76.690 133.985 77.250 ;
        RECT 134.710 77.165 134.880 77.375 ;
        RECT 134.155 76.835 134.880 77.165 ;
        RECT 133.770 76.665 133.985 76.690 ;
        RECT 133.745 76.655 133.985 76.665 ;
        RECT 133.730 76.635 133.985 76.655 ;
        RECT 133.730 76.615 133.970 76.635 ;
        RECT 133.730 76.610 133.960 76.615 ;
        RECT 133.635 76.595 133.960 76.610 ;
        RECT 133.635 76.445 133.945 76.595 ;
        RECT 133.085 76.275 133.945 76.445 ;
        RECT 134.115 76.065 134.435 76.525 ;
        RECT 134.635 76.265 134.880 76.835 ;
        RECT 135.060 76.065 135.345 77.130 ;
        RECT 135.605 77.030 135.775 77.955 ;
        RECT 135.515 76.245 135.775 77.030 ;
        RECT 135.945 77.940 136.205 78.445 ;
        RECT 136.385 78.235 136.715 78.615 ;
        RECT 136.895 78.065 137.065 78.445 ;
        RECT 135.945 77.140 136.115 77.940 ;
        RECT 136.400 77.895 137.065 78.065 ;
        RECT 136.400 77.640 136.570 77.895 ;
        RECT 137.325 77.845 139.915 78.615 ;
        RECT 136.285 77.310 136.570 77.640 ;
        RECT 136.805 77.345 137.135 77.715 ;
        RECT 137.325 77.325 138.535 77.845 ;
        RECT 140.085 77.795 140.345 78.615 ;
        RECT 140.515 77.795 140.845 78.215 ;
        RECT 141.025 78.130 141.815 78.395 ;
        RECT 140.595 77.705 140.845 77.795 ;
        RECT 136.400 77.165 136.570 77.310 ;
        RECT 135.945 76.235 136.215 77.140 ;
        RECT 136.400 76.995 137.065 77.165 ;
        RECT 138.705 77.155 139.915 77.675 ;
        RECT 136.385 76.065 136.715 76.825 ;
        RECT 136.895 76.235 137.065 76.995 ;
        RECT 137.325 76.065 139.915 77.155 ;
        RECT 140.085 76.745 140.425 77.625 ;
        RECT 140.595 77.455 141.390 77.705 ;
        RECT 140.085 76.065 140.345 76.575 ;
        RECT 140.595 76.235 140.765 77.455 ;
        RECT 141.560 77.275 141.815 78.130 ;
        RECT 141.985 77.975 142.185 78.395 ;
        RECT 142.375 78.155 142.705 78.615 ;
        RECT 141.985 77.455 142.395 77.975 ;
        RECT 142.875 77.965 143.135 78.445 ;
        RECT 142.565 77.275 142.795 77.705 ;
        RECT 141.005 77.105 142.795 77.275 ;
        RECT 141.005 76.740 141.255 77.105 ;
        RECT 141.425 76.745 141.755 76.935 ;
        RECT 141.975 76.810 142.690 77.105 ;
        RECT 142.965 76.935 143.135 77.965 ;
        RECT 143.305 77.845 144.975 78.615 ;
        RECT 145.640 77.875 146.255 78.445 ;
        RECT 146.425 78.105 146.640 78.615 ;
        RECT 146.870 78.105 147.150 78.435 ;
        RECT 147.330 78.105 147.570 78.615 ;
        RECT 143.305 77.325 144.055 77.845 ;
        RECT 144.225 77.155 144.975 77.675 ;
        RECT 141.425 76.570 141.620 76.745 ;
        RECT 141.005 76.065 141.620 76.570 ;
        RECT 141.790 76.235 142.265 76.575 ;
        RECT 142.435 76.065 142.650 76.610 ;
        RECT 142.860 76.235 143.135 76.935 ;
        RECT 143.305 76.065 144.975 77.155 ;
        RECT 145.640 76.855 145.955 77.875 ;
        RECT 146.125 77.205 146.295 77.705 ;
        RECT 146.545 77.375 146.810 77.935 ;
        RECT 146.980 77.205 147.150 78.105 ;
        RECT 147.320 77.375 147.675 77.935 ;
        RECT 147.905 77.845 151.415 78.615 ;
        RECT 151.585 77.890 151.875 78.615 ;
        RECT 152.045 77.845 155.555 78.615 ;
        RECT 155.725 77.865 156.935 78.615 ;
        RECT 147.905 77.325 149.555 77.845 ;
        RECT 146.125 77.035 147.550 77.205 ;
        RECT 149.725 77.155 151.415 77.675 ;
        RECT 152.045 77.325 153.695 77.845 ;
        RECT 145.640 76.235 146.175 76.855 ;
        RECT 146.345 76.065 146.675 76.865 ;
        RECT 147.160 76.860 147.550 77.035 ;
        RECT 147.905 76.065 151.415 77.155 ;
        RECT 151.585 76.065 151.875 77.230 ;
        RECT 153.865 77.155 155.555 77.675 ;
        RECT 152.045 76.065 155.555 77.155 ;
        RECT 155.725 77.155 156.245 77.695 ;
        RECT 156.415 77.325 156.935 77.865 ;
        RECT 155.725 76.065 156.935 77.155 ;
        RECT 22.700 75.895 157.020 76.065 ;
        RECT 22.785 74.805 23.995 75.895 ;
        RECT 24.165 74.805 25.835 75.895 ;
        RECT 26.655 75.170 26.985 75.895 ;
        RECT 22.785 74.095 23.305 74.635 ;
        RECT 23.475 74.265 23.995 74.805 ;
        RECT 24.165 74.115 24.915 74.635 ;
        RECT 25.085 74.285 25.835 74.805 ;
        RECT 22.785 73.345 23.995 74.095 ;
        RECT 24.165 73.345 25.835 74.115 ;
        RECT 26.465 73.515 26.985 75.000 ;
        RECT 27.155 74.175 27.675 75.725 ;
        RECT 27.935 75.225 28.105 75.725 ;
        RECT 28.275 75.395 28.605 75.895 ;
        RECT 27.935 75.055 28.540 75.225 ;
        RECT 27.845 74.245 28.090 74.885 ;
        RECT 28.370 74.660 28.540 75.055 ;
        RECT 28.775 74.945 29.000 75.725 ;
        RECT 28.370 74.330 28.600 74.660 ;
        RECT 28.370 74.065 28.540 74.330 ;
        RECT 27.155 73.345 27.495 74.005 ;
        RECT 27.935 73.895 28.540 74.065 ;
        RECT 27.935 73.605 28.105 73.895 ;
        RECT 28.275 73.345 28.605 73.725 ;
        RECT 28.775 73.605 28.945 74.945 ;
        RECT 29.190 74.925 29.545 75.675 ;
        RECT 29.715 75.095 30.005 75.895 ;
        RECT 30.505 75.515 31.365 75.685 ;
        RECT 31.055 75.365 31.365 75.515 ;
        RECT 31.535 75.435 31.855 75.895 ;
        RECT 31.055 75.350 31.380 75.365 ;
        RECT 31.150 75.345 31.380 75.350 ;
        RECT 31.150 75.325 31.390 75.345 ;
        RECT 31.150 75.305 31.405 75.325 ;
        RECT 31.165 75.295 31.405 75.305 ;
        RECT 31.190 75.270 31.405 75.295 ;
        RECT 29.190 74.755 29.875 74.925 ;
        RECT 29.195 74.215 29.525 74.585 ;
        RECT 29.705 74.495 29.875 74.755 ;
        RECT 30.205 74.615 30.540 75.265 ;
        RECT 30.710 74.820 31.045 75.170 ;
        RECT 29.705 74.045 30.080 74.495 ;
        RECT 30.710 74.300 31.025 74.820 ;
        RECT 31.215 74.710 31.405 75.270 ;
        RECT 32.055 75.125 32.300 75.695 ;
        RECT 31.575 74.795 32.300 75.125 ;
        RECT 32.480 74.830 32.765 75.895 ;
        RECT 32.935 74.930 33.195 75.715 ;
        RECT 29.270 74.025 30.080 74.045 ;
        RECT 29.270 73.875 29.875 74.025 ;
        RECT 30.320 73.995 31.025 74.300 ;
        RECT 31.195 74.585 31.405 74.710 ;
        RECT 32.130 74.585 32.300 74.795 ;
        RECT 31.195 74.255 31.960 74.585 ;
        RECT 32.130 74.255 32.855 74.585 ;
        RECT 29.270 73.605 29.465 73.875 ;
        RECT 31.195 73.795 31.365 74.255 ;
        RECT 32.130 73.980 32.300 74.255 ;
        RECT 33.025 74.005 33.195 74.930 ;
        RECT 34.375 74.965 34.545 75.725 ;
        RECT 34.725 75.135 35.055 75.895 ;
        RECT 34.375 74.795 35.040 74.965 ;
        RECT 35.225 74.820 35.495 75.725 ;
        RECT 34.870 74.650 35.040 74.795 ;
        RECT 34.305 74.245 34.635 74.615 ;
        RECT 34.870 74.320 35.155 74.650 ;
        RECT 34.870 74.065 35.040 74.320 ;
        RECT 29.635 73.345 29.965 73.705 ;
        RECT 30.525 73.625 31.365 73.795 ;
        RECT 31.535 73.345 31.805 73.805 ;
        RECT 32.055 73.520 32.300 73.980 ;
        RECT 32.515 73.345 32.740 73.975 ;
        RECT 32.935 73.675 33.195 74.005 ;
        RECT 34.375 73.895 35.040 74.065 ;
        RECT 35.325 74.020 35.495 74.820 ;
        RECT 35.665 74.730 35.955 75.895 ;
        RECT 36.215 75.225 36.385 75.725 ;
        RECT 36.555 75.395 36.885 75.895 ;
        RECT 36.215 75.055 36.820 75.225 ;
        RECT 36.125 74.245 36.370 74.885 ;
        RECT 36.650 74.660 36.820 75.055 ;
        RECT 37.055 74.945 37.280 75.725 ;
        RECT 36.650 74.330 36.880 74.660 ;
        RECT 34.375 73.515 34.545 73.895 ;
        RECT 34.725 73.345 35.055 73.725 ;
        RECT 35.235 73.515 35.495 74.020 ;
        RECT 35.665 73.345 35.955 74.070 ;
        RECT 36.650 74.065 36.820 74.330 ;
        RECT 36.215 73.895 36.820 74.065 ;
        RECT 36.215 73.605 36.385 73.895 ;
        RECT 36.555 73.345 36.885 73.725 ;
        RECT 37.055 73.605 37.225 74.945 ;
        RECT 37.470 74.925 37.825 75.675 ;
        RECT 37.995 75.095 38.285 75.895 ;
        RECT 38.785 75.515 39.645 75.685 ;
        RECT 39.335 75.365 39.645 75.515 ;
        RECT 39.815 75.435 40.135 75.895 ;
        RECT 39.335 75.350 39.660 75.365 ;
        RECT 39.430 75.345 39.660 75.350 ;
        RECT 39.430 75.325 39.670 75.345 ;
        RECT 39.430 75.305 39.685 75.325 ;
        RECT 39.445 75.295 39.685 75.305 ;
        RECT 39.470 75.270 39.685 75.295 ;
        RECT 37.470 74.755 38.155 74.925 ;
        RECT 37.475 74.215 37.805 74.585 ;
        RECT 37.985 74.495 38.155 74.755 ;
        RECT 38.485 74.615 38.820 75.265 ;
        RECT 38.990 74.820 39.325 75.170 ;
        RECT 37.985 74.045 38.360 74.495 ;
        RECT 38.990 74.300 39.305 74.820 ;
        RECT 39.495 74.710 39.685 75.270 ;
        RECT 40.335 75.125 40.580 75.695 ;
        RECT 39.855 74.795 40.580 75.125 ;
        RECT 40.760 74.830 41.045 75.895 ;
        RECT 41.215 74.930 41.475 75.715 ;
        RECT 37.550 74.025 38.360 74.045 ;
        RECT 37.550 73.875 38.155 74.025 ;
        RECT 38.600 73.995 39.305 74.300 ;
        RECT 39.475 74.585 39.685 74.710 ;
        RECT 40.410 74.585 40.580 74.795 ;
        RECT 39.475 74.255 40.240 74.585 ;
        RECT 40.410 74.255 41.135 74.585 ;
        RECT 37.550 73.605 37.745 73.875 ;
        RECT 39.475 73.795 39.645 74.255 ;
        RECT 40.410 73.980 40.580 74.255 ;
        RECT 41.305 74.005 41.475 74.930 ;
        RECT 41.655 74.755 41.985 75.895 ;
        RECT 42.515 74.925 42.845 75.710 ;
        RECT 43.025 75.460 48.370 75.895 ;
        RECT 42.165 74.755 42.845 74.925 ;
        RECT 41.645 74.335 41.995 74.585 ;
        RECT 42.165 74.155 42.335 74.755 ;
        RECT 42.505 74.335 42.855 74.585 ;
        RECT 37.915 73.345 38.245 73.705 ;
        RECT 38.805 73.625 39.645 73.795 ;
        RECT 39.815 73.345 40.085 73.805 ;
        RECT 40.335 73.520 40.580 73.980 ;
        RECT 40.795 73.345 41.020 73.975 ;
        RECT 41.215 73.675 41.475 74.005 ;
        RECT 41.655 73.345 41.925 74.155 ;
        RECT 42.095 73.515 42.425 74.155 ;
        RECT 42.595 73.345 42.835 74.155 ;
        RECT 44.610 73.890 44.950 74.720 ;
        RECT 46.430 74.210 46.780 75.460 ;
        RECT 48.545 74.805 50.215 75.895 ;
        RECT 48.545 74.115 49.295 74.635 ;
        RECT 49.465 74.285 50.215 74.805 ;
        RECT 50.385 74.755 50.665 75.895 ;
        RECT 50.835 74.745 51.165 75.725 ;
        RECT 51.335 74.755 51.595 75.895 ;
        RECT 51.765 74.805 55.275 75.895 ;
        RECT 55.550 75.435 55.720 75.895 ;
        RECT 55.890 75.265 56.220 75.725 ;
        RECT 50.395 74.315 50.730 74.585 ;
        RECT 50.900 74.145 51.070 74.745 ;
        RECT 51.240 74.335 51.575 74.585 ;
        RECT 43.025 73.345 48.370 73.890 ;
        RECT 48.545 73.345 50.215 74.115 ;
        RECT 50.385 73.345 50.695 74.145 ;
        RECT 50.900 73.515 51.595 74.145 ;
        RECT 51.765 74.115 53.415 74.635 ;
        RECT 53.585 74.285 55.275 74.805 ;
        RECT 55.445 75.095 56.220 75.265 ;
        RECT 56.390 75.095 56.560 75.895 ;
        RECT 51.765 73.345 55.275 74.115 ;
        RECT 55.445 74.085 55.875 75.095 ;
        RECT 57.145 74.925 57.505 75.100 ;
        RECT 56.045 74.755 57.505 74.925 ;
        RECT 57.750 74.945 58.015 75.715 ;
        RECT 58.185 75.175 58.515 75.895 ;
        RECT 58.705 75.355 58.965 75.715 ;
        RECT 59.135 75.525 59.465 75.895 ;
        RECT 59.635 75.355 59.895 75.715 ;
        RECT 58.705 75.125 59.895 75.355 ;
        RECT 60.465 74.945 60.755 75.715 ;
        RECT 56.045 74.255 56.215 74.755 ;
        RECT 55.445 73.915 56.140 74.085 ;
        RECT 56.385 74.025 56.795 74.585 ;
        RECT 55.470 73.345 55.800 73.745 ;
        RECT 55.970 73.645 56.140 73.915 ;
        RECT 56.965 73.855 57.145 74.755 ;
        RECT 57.315 74.195 57.510 74.585 ;
        RECT 57.315 74.025 57.515 74.195 ;
        RECT 56.310 73.345 56.625 73.855 ;
        RECT 56.855 73.515 57.145 73.855 ;
        RECT 57.315 73.345 57.555 73.855 ;
        RECT 57.750 73.525 58.085 74.945 ;
        RECT 58.260 74.765 60.755 74.945 ;
        RECT 58.260 74.075 58.485 74.765 ;
        RECT 61.425 74.730 61.715 75.895 ;
        RECT 61.920 75.105 62.455 75.725 ;
        RECT 58.685 74.255 58.965 74.585 ;
        RECT 59.145 74.255 59.720 74.585 ;
        RECT 59.900 74.255 60.335 74.585 ;
        RECT 60.515 74.255 60.785 74.585 ;
        RECT 61.920 74.085 62.235 75.105 ;
        RECT 62.625 75.095 62.955 75.895 ;
        RECT 63.440 74.925 63.830 75.100 ;
        RECT 62.405 74.755 63.830 74.925 ;
        RECT 64.195 74.925 64.525 75.710 ;
        RECT 64.195 74.755 64.875 74.925 ;
        RECT 65.055 74.755 65.385 75.895 ;
        RECT 65.565 74.805 66.775 75.895 ;
        RECT 67.035 75.225 67.205 75.725 ;
        RECT 67.375 75.395 67.705 75.895 ;
        RECT 67.035 75.055 67.640 75.225 ;
        RECT 62.405 74.255 62.575 74.755 ;
        RECT 58.260 73.885 60.745 74.075 ;
        RECT 58.265 73.345 59.010 73.715 ;
        RECT 59.575 73.525 59.830 73.885 ;
        RECT 60.010 73.345 60.340 73.715 ;
        RECT 60.520 73.525 60.745 73.885 ;
        RECT 61.425 73.345 61.715 74.070 ;
        RECT 61.920 73.515 62.535 74.085 ;
        RECT 62.825 74.025 63.090 74.585 ;
        RECT 63.260 73.855 63.430 74.755 ;
        RECT 63.600 74.025 63.955 74.585 ;
        RECT 64.185 74.335 64.535 74.585 ;
        RECT 64.705 74.155 64.875 74.755 ;
        RECT 65.045 74.335 65.395 74.585 ;
        RECT 62.705 73.345 62.920 73.855 ;
        RECT 63.150 73.525 63.430 73.855 ;
        RECT 63.610 73.345 63.850 73.855 ;
        RECT 64.205 73.345 64.445 74.155 ;
        RECT 64.615 73.515 64.945 74.155 ;
        RECT 65.115 73.345 65.385 74.155 ;
        RECT 65.565 74.095 66.085 74.635 ;
        RECT 66.255 74.265 66.775 74.805 ;
        RECT 66.945 74.245 67.190 74.885 ;
        RECT 67.470 74.660 67.640 75.055 ;
        RECT 67.875 74.945 68.100 75.725 ;
        RECT 67.470 74.330 67.700 74.660 ;
        RECT 65.565 73.345 66.775 74.095 ;
        RECT 67.470 74.065 67.640 74.330 ;
        RECT 67.035 73.895 67.640 74.065 ;
        RECT 67.035 73.605 67.205 73.895 ;
        RECT 67.375 73.345 67.705 73.725 ;
        RECT 67.875 73.605 68.045 74.945 ;
        RECT 68.290 74.925 68.645 75.675 ;
        RECT 68.815 75.095 69.105 75.895 ;
        RECT 69.605 75.515 70.465 75.685 ;
        RECT 70.155 75.365 70.465 75.515 ;
        RECT 70.635 75.435 70.955 75.895 ;
        RECT 70.155 75.350 70.480 75.365 ;
        RECT 70.250 75.345 70.480 75.350 ;
        RECT 70.250 75.325 70.490 75.345 ;
        RECT 70.250 75.305 70.505 75.325 ;
        RECT 70.265 75.295 70.505 75.305 ;
        RECT 70.290 75.270 70.505 75.295 ;
        RECT 68.290 74.755 68.975 74.925 ;
        RECT 68.295 74.215 68.625 74.585 ;
        RECT 68.805 74.495 68.975 74.755 ;
        RECT 69.305 74.615 69.640 75.265 ;
        RECT 69.810 74.820 70.145 75.170 ;
        RECT 68.805 74.045 69.180 74.495 ;
        RECT 69.810 74.300 70.125 74.820 ;
        RECT 70.315 74.710 70.505 75.270 ;
        RECT 71.155 75.125 71.400 75.695 ;
        RECT 70.675 74.795 71.400 75.125 ;
        RECT 71.580 74.830 71.865 75.895 ;
        RECT 72.035 74.930 72.295 75.715 ;
        RECT 68.370 74.025 69.180 74.045 ;
        RECT 68.370 73.875 68.975 74.025 ;
        RECT 69.420 73.995 70.125 74.300 ;
        RECT 70.295 74.585 70.505 74.710 ;
        RECT 71.230 74.585 71.400 74.795 ;
        RECT 70.295 74.255 71.060 74.585 ;
        RECT 71.230 74.255 71.955 74.585 ;
        RECT 68.370 73.605 68.565 73.875 ;
        RECT 70.295 73.795 70.465 74.255 ;
        RECT 71.230 73.980 71.400 74.255 ;
        RECT 72.125 74.005 72.295 74.930 ;
        RECT 72.475 74.925 72.805 75.710 ;
        RECT 72.475 74.755 73.155 74.925 ;
        RECT 73.335 74.755 73.665 75.895 ;
        RECT 73.845 74.805 75.055 75.895 ;
        RECT 72.465 74.335 72.815 74.585 ;
        RECT 72.985 74.155 73.155 74.755 ;
        RECT 73.325 74.335 73.675 74.585 ;
        RECT 68.735 73.345 69.065 73.705 ;
        RECT 69.625 73.625 70.465 73.795 ;
        RECT 70.635 73.345 70.905 73.805 ;
        RECT 71.155 73.520 71.400 73.980 ;
        RECT 71.615 73.345 71.840 73.975 ;
        RECT 72.035 73.675 72.295 74.005 ;
        RECT 72.485 73.345 72.725 74.155 ;
        RECT 72.895 73.515 73.225 74.155 ;
        RECT 73.395 73.345 73.665 74.155 ;
        RECT 73.845 74.095 74.365 74.635 ;
        RECT 74.535 74.265 75.055 74.805 ;
        RECT 75.225 75.025 75.500 75.725 ;
        RECT 75.710 75.350 75.925 75.895 ;
        RECT 76.095 75.385 76.570 75.725 ;
        RECT 76.740 75.390 77.355 75.895 ;
        RECT 76.740 75.215 76.935 75.390 ;
        RECT 73.845 73.345 75.055 74.095 ;
        RECT 75.225 73.995 75.395 75.025 ;
        RECT 75.670 74.855 76.385 75.150 ;
        RECT 76.605 75.025 76.935 75.215 ;
        RECT 77.105 74.855 77.355 75.220 ;
        RECT 75.565 74.685 77.355 74.855 ;
        RECT 75.565 74.255 75.795 74.685 ;
        RECT 75.225 73.515 75.485 73.995 ;
        RECT 75.965 73.985 76.375 74.505 ;
        RECT 75.655 73.345 75.985 73.805 ;
        RECT 76.175 73.565 76.375 73.985 ;
        RECT 76.545 73.830 76.800 74.685 ;
        RECT 77.595 74.505 77.765 75.725 ;
        RECT 78.015 75.385 78.275 75.895 ;
        RECT 76.970 74.255 77.765 74.505 ;
        RECT 77.935 74.335 78.275 75.215 ;
        RECT 78.445 74.805 81.955 75.895 ;
        RECT 77.515 74.165 77.765 74.255 ;
        RECT 76.545 73.565 77.335 73.830 ;
        RECT 77.515 73.745 77.845 74.165 ;
        RECT 78.015 73.345 78.275 74.165 ;
        RECT 78.445 74.115 80.095 74.635 ;
        RECT 80.265 74.285 81.955 74.805 ;
        RECT 83.055 74.755 83.385 75.895 ;
        RECT 83.915 74.925 84.245 75.710 ;
        RECT 83.565 74.755 84.245 74.925 ;
        RECT 84.425 74.805 85.635 75.895 ;
        RECT 83.045 74.335 83.395 74.585 ;
        RECT 83.565 74.155 83.735 74.755 ;
        RECT 83.905 74.335 84.255 74.585 ;
        RECT 78.445 73.345 81.955 74.115 ;
        RECT 83.055 73.345 83.325 74.155 ;
        RECT 83.495 73.515 83.825 74.155 ;
        RECT 83.995 73.345 84.235 74.155 ;
        RECT 84.425 74.095 84.945 74.635 ;
        RECT 85.115 74.265 85.635 74.805 ;
        RECT 85.845 74.755 86.075 75.895 ;
        RECT 86.245 74.745 86.575 75.725 ;
        RECT 86.745 74.755 86.955 75.895 ;
        RECT 85.825 74.335 86.155 74.585 ;
        RECT 84.425 73.345 85.635 74.095 ;
        RECT 85.845 73.345 86.075 74.165 ;
        RECT 86.325 74.145 86.575 74.745 ;
        RECT 87.185 74.730 87.475 75.895 ;
        RECT 88.110 74.755 88.385 75.725 ;
        RECT 88.595 75.095 88.875 75.895 ;
        RECT 89.045 75.385 90.235 75.675 ;
        RECT 89.045 75.045 90.215 75.215 ;
        RECT 89.045 74.925 89.215 75.045 ;
        RECT 88.555 74.755 89.215 74.925 ;
        RECT 86.245 73.515 86.575 74.145 ;
        RECT 86.745 73.345 86.955 74.165 ;
        RECT 87.185 73.345 87.475 74.070 ;
        RECT 88.110 74.020 88.280 74.755 ;
        RECT 88.555 74.585 88.725 74.755 ;
        RECT 89.525 74.585 89.720 74.875 ;
        RECT 89.890 74.755 90.215 75.045 ;
        RECT 90.495 74.965 90.665 75.725 ;
        RECT 90.845 75.135 91.175 75.895 ;
        RECT 90.495 74.795 91.160 74.965 ;
        RECT 91.345 74.820 91.615 75.725 ;
        RECT 90.990 74.650 91.160 74.795 ;
        RECT 88.450 74.255 88.725 74.585 ;
        RECT 88.895 74.255 89.720 74.585 ;
        RECT 89.890 74.255 90.235 74.585 ;
        RECT 88.555 74.085 88.725 74.255 ;
        RECT 90.425 74.245 90.755 74.615 ;
        RECT 90.990 74.320 91.275 74.650 ;
        RECT 88.110 73.675 88.385 74.020 ;
        RECT 88.555 73.915 90.220 74.085 ;
        RECT 90.990 74.065 91.160 74.320 ;
        RECT 88.575 73.345 88.955 73.745 ;
        RECT 89.125 73.565 89.295 73.915 ;
        RECT 89.465 73.345 89.795 73.745 ;
        RECT 89.965 73.565 90.220 73.915 ;
        RECT 90.495 73.895 91.160 74.065 ;
        RECT 91.445 74.020 91.615 74.820 ;
        RECT 91.785 74.805 94.375 75.895 ;
        RECT 90.495 73.515 90.665 73.895 ;
        RECT 90.845 73.345 91.175 73.725 ;
        RECT 91.355 73.515 91.615 74.020 ;
        RECT 91.785 74.115 92.995 74.635 ;
        RECT 93.165 74.285 94.375 74.805 ;
        RECT 95.015 74.755 95.345 75.895 ;
        RECT 95.875 74.925 96.205 75.710 ;
        RECT 96.585 75.225 96.865 75.895 ;
        RECT 97.035 75.005 97.335 75.555 ;
        RECT 97.535 75.175 97.865 75.895 ;
        RECT 98.055 75.175 98.515 75.725 ;
        RECT 99.145 75.385 100.335 75.675 ;
        RECT 95.525 74.755 96.205 74.925 ;
        RECT 95.005 74.335 95.355 74.585 ;
        RECT 95.525 74.155 95.695 74.755 ;
        RECT 96.400 74.585 96.665 74.945 ;
        RECT 97.035 74.835 97.975 75.005 ;
        RECT 97.805 74.585 97.975 74.835 ;
        RECT 95.865 74.335 96.215 74.585 ;
        RECT 96.400 74.335 97.075 74.585 ;
        RECT 97.295 74.335 97.635 74.585 ;
        RECT 97.805 74.255 98.095 74.585 ;
        RECT 97.805 74.165 97.975 74.255 ;
        RECT 91.785 73.345 94.375 74.115 ;
        RECT 95.015 73.345 95.285 74.155 ;
        RECT 95.455 73.515 95.785 74.155 ;
        RECT 95.955 73.345 96.195 74.155 ;
        RECT 96.585 73.975 97.975 74.165 ;
        RECT 96.585 73.615 96.915 73.975 ;
        RECT 98.265 73.805 98.515 75.175 ;
        RECT 99.165 75.045 100.335 75.215 ;
        RECT 100.505 75.095 100.785 75.895 ;
        RECT 99.165 74.755 99.490 75.045 ;
        RECT 100.165 74.925 100.335 75.045 ;
        RECT 99.660 74.585 99.855 74.875 ;
        RECT 100.165 74.755 100.825 74.925 ;
        RECT 100.995 74.755 101.270 75.725 ;
        RECT 101.535 75.225 101.705 75.725 ;
        RECT 101.875 75.395 102.205 75.895 ;
        RECT 101.535 75.055 102.140 75.225 ;
        RECT 100.655 74.585 100.825 74.755 ;
        RECT 99.145 74.255 99.490 74.585 ;
        RECT 99.660 74.255 100.485 74.585 ;
        RECT 100.655 74.255 100.930 74.585 ;
        RECT 100.655 74.085 100.825 74.255 ;
        RECT 97.535 73.345 97.785 73.805 ;
        RECT 97.955 73.515 98.515 73.805 ;
        RECT 99.160 73.915 100.825 74.085 ;
        RECT 101.100 74.020 101.270 74.755 ;
        RECT 101.445 74.245 101.690 74.885 ;
        RECT 101.970 74.660 102.140 75.055 ;
        RECT 102.375 74.945 102.600 75.725 ;
        RECT 101.970 74.330 102.200 74.660 ;
        RECT 101.970 74.065 102.140 74.330 ;
        RECT 99.160 73.565 99.415 73.915 ;
        RECT 99.585 73.345 99.915 73.745 ;
        RECT 100.085 73.565 100.255 73.915 ;
        RECT 100.425 73.345 100.805 73.745 ;
        RECT 100.995 73.675 101.270 74.020 ;
        RECT 101.535 73.895 102.140 74.065 ;
        RECT 101.535 73.605 101.705 73.895 ;
        RECT 101.875 73.345 102.205 73.725 ;
        RECT 102.375 73.605 102.545 74.945 ;
        RECT 102.790 74.925 103.145 75.675 ;
        RECT 103.315 75.095 103.605 75.895 ;
        RECT 104.105 75.515 104.965 75.685 ;
        RECT 104.655 75.365 104.965 75.515 ;
        RECT 105.135 75.435 105.455 75.895 ;
        RECT 104.655 75.350 104.980 75.365 ;
        RECT 104.750 75.345 104.980 75.350 ;
        RECT 104.750 75.325 104.990 75.345 ;
        RECT 104.750 75.305 105.005 75.325 ;
        RECT 104.765 75.295 105.005 75.305 ;
        RECT 104.790 75.270 105.005 75.295 ;
        RECT 102.790 74.755 103.475 74.925 ;
        RECT 102.795 74.215 103.125 74.585 ;
        RECT 103.305 74.495 103.475 74.755 ;
        RECT 103.805 74.615 104.140 75.265 ;
        RECT 104.310 74.820 104.645 75.170 ;
        RECT 103.305 74.045 103.680 74.495 ;
        RECT 104.310 74.300 104.625 74.820 ;
        RECT 104.815 74.710 105.005 75.270 ;
        RECT 105.655 75.125 105.900 75.695 ;
        RECT 105.175 74.795 105.900 75.125 ;
        RECT 106.080 74.830 106.365 75.895 ;
        RECT 106.535 74.930 106.795 75.715 ;
        RECT 102.870 74.025 103.680 74.045 ;
        RECT 102.870 73.875 103.475 74.025 ;
        RECT 103.920 73.995 104.625 74.300 ;
        RECT 104.795 74.585 105.005 74.710 ;
        RECT 105.730 74.585 105.900 74.795 ;
        RECT 104.795 74.255 105.560 74.585 ;
        RECT 105.730 74.255 106.455 74.585 ;
        RECT 102.870 73.605 103.065 73.875 ;
        RECT 104.795 73.795 104.965 74.255 ;
        RECT 105.730 73.980 105.900 74.255 ;
        RECT 106.625 74.005 106.795 74.930 ;
        RECT 107.150 74.925 107.540 75.100 ;
        RECT 108.025 75.095 108.355 75.895 ;
        RECT 108.525 75.105 109.060 75.725 ;
        RECT 109.725 75.385 109.985 75.895 ;
        RECT 107.150 74.755 108.575 74.925 ;
        RECT 107.025 74.025 107.380 74.585 ;
        RECT 103.235 73.345 103.565 73.705 ;
        RECT 104.125 73.625 104.965 73.795 ;
        RECT 105.135 73.345 105.405 73.805 ;
        RECT 105.655 73.520 105.900 73.980 ;
        RECT 106.115 73.345 106.340 73.975 ;
        RECT 106.535 73.675 106.795 74.005 ;
        RECT 107.550 73.855 107.720 74.755 ;
        RECT 107.890 74.025 108.155 74.585 ;
        RECT 108.405 74.255 108.575 74.755 ;
        RECT 108.745 74.085 109.060 75.105 ;
        RECT 109.725 74.335 110.065 75.215 ;
        RECT 110.235 74.505 110.405 75.725 ;
        RECT 110.645 75.390 111.260 75.895 ;
        RECT 110.645 74.855 110.895 75.220 ;
        RECT 111.065 75.215 111.260 75.390 ;
        RECT 111.430 75.385 111.905 75.725 ;
        RECT 112.075 75.350 112.290 75.895 ;
        RECT 111.065 75.025 111.395 75.215 ;
        RECT 111.615 74.855 112.330 75.150 ;
        RECT 112.500 75.025 112.775 75.725 ;
        RECT 110.645 74.685 112.435 74.855 ;
        RECT 110.235 74.255 111.030 74.505 ;
        RECT 110.235 74.165 110.485 74.255 ;
        RECT 107.130 73.345 107.370 73.855 ;
        RECT 107.550 73.525 107.830 73.855 ;
        RECT 108.060 73.345 108.275 73.855 ;
        RECT 108.445 73.515 109.060 74.085 ;
        RECT 109.725 73.345 109.985 74.165 ;
        RECT 110.155 73.745 110.485 74.165 ;
        RECT 111.200 73.830 111.455 74.685 ;
        RECT 110.665 73.565 111.455 73.830 ;
        RECT 111.625 73.985 112.035 74.505 ;
        RECT 112.205 74.255 112.435 74.685 ;
        RECT 112.605 73.995 112.775 75.025 ;
        RECT 112.945 74.730 113.235 75.895 ;
        RECT 113.405 74.755 113.665 75.895 ;
        RECT 113.835 74.745 114.165 75.725 ;
        RECT 114.335 74.755 114.615 75.895 ;
        RECT 114.795 74.835 115.125 75.685 ;
        RECT 113.425 74.335 113.760 74.585 ;
        RECT 113.930 74.145 114.100 74.745 ;
        RECT 114.270 74.315 114.605 74.585 ;
        RECT 111.625 73.565 111.825 73.985 ;
        RECT 112.015 73.345 112.345 73.805 ;
        RECT 112.515 73.515 112.775 73.995 ;
        RECT 112.945 73.345 113.235 74.070 ;
        RECT 113.405 73.515 114.100 74.145 ;
        RECT 114.305 73.345 114.615 74.145 ;
        RECT 114.795 74.070 114.985 74.835 ;
        RECT 115.295 74.755 115.545 75.895 ;
        RECT 115.735 75.255 115.985 75.675 ;
        RECT 116.215 75.425 116.545 75.895 ;
        RECT 116.775 75.255 117.025 75.675 ;
        RECT 115.735 75.085 117.025 75.255 ;
        RECT 117.205 75.255 117.535 75.685 ;
        RECT 117.205 75.085 117.660 75.255 ;
        RECT 115.725 74.585 115.940 74.915 ;
        RECT 115.155 74.255 115.465 74.585 ;
        RECT 115.635 74.255 115.940 74.585 ;
        RECT 116.115 74.255 116.400 74.915 ;
        RECT 116.595 74.255 116.860 74.915 ;
        RECT 117.075 74.255 117.320 74.915 ;
        RECT 115.295 74.085 115.465 74.255 ;
        RECT 117.490 74.085 117.660 75.085 ;
        RECT 118.015 74.925 118.345 75.710 ;
        RECT 118.015 74.755 118.695 74.925 ;
        RECT 118.875 74.755 119.205 75.895 ;
        RECT 119.385 74.805 122.895 75.895 ;
        RECT 118.005 74.335 118.355 74.585 ;
        RECT 118.525 74.155 118.695 74.755 ;
        RECT 118.865 74.335 119.215 74.585 ;
        RECT 114.795 73.560 115.125 74.070 ;
        RECT 115.295 73.915 117.660 74.085 ;
        RECT 115.295 73.345 115.625 73.745 ;
        RECT 116.675 73.575 117.005 73.915 ;
        RECT 117.175 73.345 117.505 73.745 ;
        RECT 118.025 73.345 118.265 74.155 ;
        RECT 118.435 73.515 118.765 74.155 ;
        RECT 118.935 73.345 119.205 74.155 ;
        RECT 119.385 74.115 121.035 74.635 ;
        RECT 121.205 74.285 122.895 74.805 ;
        RECT 123.075 74.755 123.405 75.895 ;
        RECT 123.935 74.925 124.265 75.710 ;
        RECT 123.585 74.755 124.265 74.925 ;
        RECT 124.445 74.805 127.035 75.895 ;
        RECT 123.065 74.335 123.415 74.585 ;
        RECT 123.585 74.155 123.755 74.755 ;
        RECT 123.925 74.335 124.275 74.585 ;
        RECT 119.385 73.345 122.895 74.115 ;
        RECT 123.075 73.345 123.345 74.155 ;
        RECT 123.515 73.515 123.845 74.155 ;
        RECT 124.015 73.345 124.255 74.155 ;
        RECT 124.445 74.115 125.655 74.635 ;
        RECT 125.825 74.285 127.035 74.805 ;
        RECT 127.705 74.755 127.935 75.895 ;
        RECT 128.105 74.745 128.435 75.725 ;
        RECT 128.605 74.755 128.815 75.895 ;
        RECT 129.045 74.805 130.715 75.895 ;
        RECT 130.885 75.385 132.075 75.675 ;
        RECT 127.685 74.335 128.015 74.585 ;
        RECT 124.445 73.345 127.035 74.115 ;
        RECT 127.705 73.345 127.935 74.165 ;
        RECT 128.185 74.145 128.435 74.745 ;
        RECT 128.105 73.515 128.435 74.145 ;
        RECT 128.605 73.345 128.815 74.165 ;
        RECT 129.045 74.115 129.795 74.635 ;
        RECT 129.965 74.285 130.715 74.805 ;
        RECT 130.905 75.045 132.075 75.215 ;
        RECT 132.245 75.095 132.525 75.895 ;
        RECT 130.905 74.755 131.230 75.045 ;
        RECT 131.905 74.925 132.075 75.045 ;
        RECT 131.400 74.585 131.595 74.875 ;
        RECT 131.905 74.755 132.565 74.925 ;
        RECT 132.735 74.755 133.010 75.725 ;
        RECT 133.185 74.805 134.855 75.895 ;
        RECT 132.395 74.585 132.565 74.755 ;
        RECT 130.885 74.255 131.230 74.585 ;
        RECT 131.400 74.255 132.225 74.585 ;
        RECT 132.395 74.255 132.670 74.585 ;
        RECT 129.045 73.345 130.715 74.115 ;
        RECT 132.395 74.085 132.565 74.255 ;
        RECT 130.900 73.915 132.565 74.085 ;
        RECT 132.840 74.020 133.010 74.755 ;
        RECT 130.900 73.565 131.155 73.915 ;
        RECT 131.325 73.345 131.655 73.745 ;
        RECT 131.825 73.565 131.995 73.915 ;
        RECT 132.165 73.345 132.545 73.745 ;
        RECT 132.735 73.675 133.010 74.020 ;
        RECT 133.185 74.115 133.935 74.635 ;
        RECT 134.105 74.285 134.855 74.805 ;
        RECT 135.035 74.755 135.365 75.895 ;
        RECT 135.895 74.925 136.225 75.710 ;
        RECT 135.545 74.755 136.225 74.925 ;
        RECT 137.415 74.965 137.585 75.725 ;
        RECT 137.765 75.135 138.095 75.895 ;
        RECT 137.415 74.795 138.080 74.965 ;
        RECT 138.265 74.820 138.535 75.725 ;
        RECT 135.025 74.335 135.375 74.585 ;
        RECT 135.545 74.155 135.715 74.755 ;
        RECT 137.910 74.650 138.080 74.795 ;
        RECT 135.885 74.335 136.235 74.585 ;
        RECT 137.345 74.245 137.675 74.615 ;
        RECT 137.910 74.320 138.195 74.650 ;
        RECT 133.185 73.345 134.855 74.115 ;
        RECT 135.035 73.345 135.305 74.155 ;
        RECT 135.475 73.515 135.805 74.155 ;
        RECT 135.975 73.345 136.215 74.155 ;
        RECT 137.910 74.065 138.080 74.320 ;
        RECT 137.415 73.895 138.080 74.065 ;
        RECT 138.365 74.020 138.535 74.820 ;
        RECT 138.705 74.730 138.995 75.895 ;
        RECT 140.275 75.170 140.605 75.895 ;
        RECT 137.415 73.515 137.585 73.895 ;
        RECT 137.765 73.345 138.095 73.725 ;
        RECT 138.275 73.515 138.535 74.020 ;
        RECT 138.705 73.345 138.995 74.070 ;
        RECT 140.085 73.515 140.605 75.000 ;
        RECT 140.775 74.175 141.295 75.725 ;
        RECT 141.555 75.225 141.725 75.725 ;
        RECT 141.895 75.395 142.225 75.895 ;
        RECT 141.555 75.055 142.160 75.225 ;
        RECT 141.465 74.245 141.710 74.885 ;
        RECT 141.990 74.660 142.160 75.055 ;
        RECT 142.395 74.945 142.620 75.725 ;
        RECT 141.990 74.330 142.220 74.660 ;
        RECT 141.990 74.065 142.160 74.330 ;
        RECT 140.775 73.345 141.115 74.005 ;
        RECT 141.555 73.895 142.160 74.065 ;
        RECT 141.555 73.605 141.725 73.895 ;
        RECT 141.895 73.345 142.225 73.725 ;
        RECT 142.395 73.605 142.565 74.945 ;
        RECT 142.810 74.925 143.165 75.675 ;
        RECT 143.335 75.095 143.625 75.895 ;
        RECT 144.125 75.515 144.985 75.685 ;
        RECT 144.675 75.365 144.985 75.515 ;
        RECT 145.155 75.435 145.475 75.895 ;
        RECT 144.675 75.350 145.000 75.365 ;
        RECT 144.770 75.345 145.000 75.350 ;
        RECT 144.770 75.325 145.010 75.345 ;
        RECT 144.770 75.305 145.025 75.325 ;
        RECT 144.785 75.295 145.025 75.305 ;
        RECT 144.810 75.270 145.025 75.295 ;
        RECT 142.810 74.755 143.495 74.925 ;
        RECT 142.815 74.215 143.145 74.585 ;
        RECT 143.325 74.495 143.495 74.755 ;
        RECT 143.825 74.615 144.160 75.265 ;
        RECT 144.330 74.820 144.665 75.170 ;
        RECT 143.325 74.045 143.700 74.495 ;
        RECT 144.330 74.300 144.645 74.820 ;
        RECT 144.835 74.710 145.025 75.270 ;
        RECT 145.675 75.125 145.920 75.695 ;
        RECT 145.195 74.795 145.920 75.125 ;
        RECT 146.100 74.830 146.385 75.895 ;
        RECT 146.555 74.930 146.815 75.715 ;
        RECT 146.985 75.460 152.330 75.895 ;
        RECT 142.890 74.025 143.700 74.045 ;
        RECT 142.890 73.875 143.495 74.025 ;
        RECT 143.940 73.995 144.645 74.300 ;
        RECT 144.815 74.585 145.025 74.710 ;
        RECT 145.750 74.585 145.920 74.795 ;
        RECT 144.815 74.255 145.580 74.585 ;
        RECT 145.750 74.255 146.475 74.585 ;
        RECT 142.890 73.605 143.085 73.875 ;
        RECT 144.815 73.795 144.985 74.255 ;
        RECT 145.750 73.980 145.920 74.255 ;
        RECT 146.645 74.005 146.815 74.930 ;
        RECT 143.255 73.345 143.585 73.705 ;
        RECT 144.145 73.625 144.985 73.795 ;
        RECT 145.155 73.345 145.425 73.805 ;
        RECT 145.675 73.520 145.920 73.980 ;
        RECT 146.135 73.345 146.360 73.975 ;
        RECT 146.555 73.675 146.815 74.005 ;
        RECT 148.570 73.890 148.910 74.720 ;
        RECT 150.390 74.210 150.740 75.460 ;
        RECT 152.505 74.805 155.095 75.895 ;
        RECT 152.505 74.115 153.715 74.635 ;
        RECT 153.885 74.285 155.095 74.805 ;
        RECT 155.725 74.805 156.935 75.895 ;
        RECT 155.725 74.265 156.245 74.805 ;
        RECT 146.985 73.345 152.330 73.890 ;
        RECT 152.505 73.345 155.095 74.115 ;
        RECT 156.415 74.095 156.935 74.635 ;
        RECT 155.725 73.345 156.935 74.095 ;
        RECT 22.700 73.175 157.020 73.345 ;
        RECT 22.785 72.425 23.995 73.175 ;
        RECT 24.165 72.630 29.510 73.175 ;
        RECT 29.685 72.630 35.030 73.175 ;
        RECT 22.785 71.885 23.305 72.425 ;
        RECT 23.475 71.715 23.995 72.255 ;
        RECT 25.750 71.800 26.090 72.630 ;
        RECT 22.785 70.625 23.995 71.715 ;
        RECT 27.570 71.060 27.920 72.310 ;
        RECT 31.270 71.800 31.610 72.630 ;
        RECT 35.205 72.405 37.795 73.175 ;
        RECT 33.090 71.060 33.440 72.310 ;
        RECT 35.205 71.885 36.415 72.405 ;
        RECT 38.005 72.355 38.235 73.175 ;
        RECT 38.405 72.375 38.735 73.005 ;
        RECT 36.585 71.715 37.795 72.235 ;
        RECT 37.985 71.935 38.315 72.185 ;
        RECT 38.485 71.775 38.735 72.375 ;
        RECT 38.905 72.355 39.115 73.175 ;
        RECT 39.365 72.445 39.655 73.175 ;
        RECT 39.355 71.935 39.655 72.265 ;
        RECT 39.835 72.245 40.065 72.885 ;
        RECT 40.245 72.625 40.555 72.995 ;
        RECT 40.735 72.805 41.405 73.175 ;
        RECT 40.245 72.425 41.475 72.625 ;
        RECT 39.835 71.935 40.360 72.245 ;
        RECT 40.540 71.935 41.005 72.245 ;
        RECT 24.165 70.625 29.510 71.060 ;
        RECT 29.685 70.625 35.030 71.060 ;
        RECT 35.205 70.625 37.795 71.715 ;
        RECT 38.005 70.625 38.235 71.765 ;
        RECT 38.405 70.795 38.735 71.775 ;
        RECT 38.905 70.625 39.115 71.765 ;
        RECT 41.185 71.755 41.475 72.425 ;
        RECT 39.365 71.515 40.525 71.755 ;
        RECT 39.365 70.805 39.625 71.515 ;
        RECT 39.795 70.625 40.125 71.335 ;
        RECT 40.295 70.805 40.525 71.515 ;
        RECT 40.705 71.535 41.475 71.755 ;
        RECT 40.705 70.805 40.975 71.535 ;
        RECT 41.155 70.625 41.495 71.355 ;
        RECT 41.665 70.805 41.925 72.995 ;
        RECT 43.040 72.605 43.295 72.955 ;
        RECT 43.465 72.775 43.795 73.175 ;
        RECT 43.965 72.605 44.135 72.955 ;
        RECT 44.305 72.775 44.685 73.175 ;
        RECT 43.040 72.435 44.705 72.605 ;
        RECT 44.875 72.500 45.150 72.845 ;
        RECT 44.535 72.265 44.705 72.435 ;
        RECT 43.025 71.935 43.370 72.265 ;
        RECT 43.540 71.935 44.365 72.265 ;
        RECT 44.535 71.935 44.810 72.265 ;
        RECT 43.045 71.475 43.370 71.765 ;
        RECT 43.540 71.645 43.735 71.935 ;
        RECT 44.535 71.765 44.705 71.935 ;
        RECT 44.980 71.765 45.150 72.500 ;
        RECT 45.325 72.405 47.915 73.175 ;
        RECT 48.545 72.450 48.835 73.175 ;
        RECT 49.005 72.425 50.215 73.175 ;
        RECT 45.325 71.885 46.535 72.405 ;
        RECT 44.045 71.595 44.705 71.765 ;
        RECT 44.045 71.475 44.215 71.595 ;
        RECT 43.045 71.305 44.215 71.475 ;
        RECT 43.025 70.845 44.215 71.135 ;
        RECT 44.385 70.625 44.665 71.425 ;
        RECT 44.875 70.795 45.150 71.765 ;
        RECT 46.705 71.715 47.915 72.235 ;
        RECT 49.005 71.885 49.525 72.425 ;
        RECT 50.395 72.365 50.665 73.175 ;
        RECT 50.835 72.365 51.165 73.005 ;
        RECT 51.335 72.365 51.575 73.175 ;
        RECT 52.230 72.500 52.505 72.845 ;
        RECT 52.695 72.775 53.075 73.175 ;
        RECT 53.245 72.605 53.415 72.955 ;
        RECT 53.585 72.775 53.915 73.175 ;
        RECT 54.085 72.605 54.340 72.955 ;
        RECT 45.325 70.625 47.915 71.715 ;
        RECT 48.545 70.625 48.835 71.790 ;
        RECT 49.695 71.715 50.215 72.255 ;
        RECT 50.385 71.935 50.735 72.185 ;
        RECT 50.905 71.765 51.075 72.365 ;
        RECT 51.245 71.935 51.595 72.185 ;
        RECT 52.230 71.765 52.400 72.500 ;
        RECT 52.675 72.435 54.340 72.605 ;
        RECT 52.675 72.265 52.845 72.435 ;
        RECT 54.565 72.355 54.795 73.175 ;
        RECT 54.965 72.375 55.295 73.005 ;
        RECT 52.570 71.935 52.845 72.265 ;
        RECT 53.015 71.935 53.840 72.265 ;
        RECT 54.010 71.935 54.355 72.265 ;
        RECT 54.545 71.935 54.875 72.185 ;
        RECT 52.675 71.765 52.845 71.935 ;
        RECT 49.005 70.625 50.215 71.715 ;
        RECT 50.395 70.625 50.725 71.765 ;
        RECT 50.905 71.595 51.585 71.765 ;
        RECT 51.255 70.810 51.585 71.595 ;
        RECT 52.230 70.795 52.505 71.765 ;
        RECT 52.675 71.595 53.335 71.765 ;
        RECT 53.645 71.645 53.840 71.935 ;
        RECT 55.045 71.775 55.295 72.375 ;
        RECT 55.465 72.355 55.675 73.175 ;
        RECT 55.905 72.425 57.115 73.175 ;
        RECT 55.905 71.885 56.425 72.425 ;
        RECT 57.295 72.365 57.565 73.175 ;
        RECT 57.735 72.365 58.065 73.005 ;
        RECT 58.235 72.365 58.475 73.175 ;
        RECT 58.665 72.405 60.335 73.175 ;
        RECT 53.165 71.475 53.335 71.595 ;
        RECT 54.010 71.475 54.335 71.765 ;
        RECT 52.715 70.625 52.995 71.425 ;
        RECT 53.165 71.305 54.335 71.475 ;
        RECT 53.165 70.845 54.355 71.135 ;
        RECT 54.565 70.625 54.795 71.765 ;
        RECT 54.965 70.795 55.295 71.775 ;
        RECT 55.465 70.625 55.675 71.765 ;
        RECT 56.595 71.715 57.115 72.255 ;
        RECT 57.285 71.935 57.635 72.185 ;
        RECT 57.805 71.765 57.975 72.365 ;
        RECT 58.145 71.935 58.495 72.185 ;
        RECT 58.665 71.885 59.415 72.405 ;
        RECT 60.965 72.375 61.275 73.175 ;
        RECT 61.480 72.375 62.175 73.005 ;
        RECT 62.345 72.405 64.935 73.175 ;
        RECT 65.655 72.625 65.825 72.915 ;
        RECT 65.995 72.795 66.325 73.175 ;
        RECT 65.655 72.455 66.260 72.625 ;
        RECT 55.905 70.625 57.115 71.715 ;
        RECT 57.295 70.625 57.625 71.765 ;
        RECT 57.805 71.595 58.485 71.765 ;
        RECT 59.585 71.715 60.335 72.235 ;
        RECT 60.975 71.935 61.310 72.205 ;
        RECT 61.480 71.775 61.650 72.375 ;
        RECT 61.820 71.935 62.155 72.185 ;
        RECT 62.345 71.885 63.555 72.405 ;
        RECT 58.155 70.810 58.485 71.595 ;
        RECT 58.665 70.625 60.335 71.715 ;
        RECT 60.965 70.625 61.245 71.765 ;
        RECT 61.415 70.795 61.745 71.775 ;
        RECT 61.915 70.625 62.175 71.765 ;
        RECT 63.725 71.715 64.935 72.235 ;
        RECT 62.345 70.625 64.935 71.715 ;
        RECT 65.565 71.635 65.810 72.275 ;
        RECT 66.090 72.190 66.260 72.455 ;
        RECT 66.090 71.860 66.320 72.190 ;
        RECT 66.090 71.465 66.260 71.860 ;
        RECT 65.655 71.295 66.260 71.465 ;
        RECT 66.495 71.575 66.665 72.915 ;
        RECT 66.990 72.645 67.185 72.915 ;
        RECT 67.355 72.815 67.685 73.175 ;
        RECT 68.245 72.725 69.085 72.895 ;
        RECT 66.990 72.495 67.595 72.645 ;
        RECT 66.990 72.475 67.800 72.495 ;
        RECT 66.915 71.935 67.245 72.305 ;
        RECT 67.425 72.025 67.800 72.475 ;
        RECT 68.040 72.220 68.745 72.525 ;
        RECT 67.425 71.765 67.595 72.025 ;
        RECT 66.910 71.595 67.595 71.765 ;
        RECT 65.655 70.795 65.825 71.295 ;
        RECT 65.995 70.625 66.325 71.125 ;
        RECT 66.495 70.795 66.720 71.575 ;
        RECT 66.910 70.845 67.265 71.595 ;
        RECT 67.435 70.625 67.725 71.425 ;
        RECT 67.925 71.255 68.260 71.905 ;
        RECT 68.430 71.700 68.745 72.220 ;
        RECT 68.915 72.265 69.085 72.725 ;
        RECT 69.255 72.715 69.525 73.175 ;
        RECT 69.775 72.540 70.020 73.000 ;
        RECT 70.235 72.545 70.460 73.175 ;
        RECT 69.850 72.265 70.020 72.540 ;
        RECT 70.655 72.515 70.915 72.845 ;
        RECT 68.915 71.935 69.680 72.265 ;
        RECT 69.850 71.935 70.575 72.265 ;
        RECT 68.915 71.810 69.125 71.935 ;
        RECT 68.430 71.350 68.765 71.700 ;
        RECT 68.935 71.250 69.125 71.810 ;
        RECT 69.850 71.725 70.020 71.935 ;
        RECT 69.295 71.395 70.020 71.725 ;
        RECT 68.910 71.225 69.125 71.250 ;
        RECT 68.885 71.215 69.125 71.225 ;
        RECT 68.870 71.195 69.125 71.215 ;
        RECT 68.870 71.175 69.110 71.195 ;
        RECT 68.870 71.170 69.100 71.175 ;
        RECT 68.775 71.155 69.100 71.170 ;
        RECT 68.775 71.005 69.085 71.155 ;
        RECT 68.225 70.835 69.085 71.005 ;
        RECT 69.255 70.625 69.575 71.085 ;
        RECT 69.775 70.825 70.020 71.395 ;
        RECT 70.200 70.625 70.485 71.690 ;
        RECT 70.745 71.590 70.915 72.515 ;
        RECT 71.085 72.405 73.675 73.175 ;
        RECT 74.305 72.450 74.595 73.175 ;
        RECT 71.085 71.885 72.295 72.405 ;
        RECT 74.765 72.375 75.075 73.175 ;
        RECT 75.280 72.375 75.975 73.005 ;
        RECT 76.145 72.405 78.735 73.175 ;
        RECT 79.370 72.670 79.705 73.175 ;
        RECT 79.875 72.605 80.115 72.980 ;
        RECT 80.395 72.845 80.565 72.990 ;
        RECT 80.395 72.650 80.770 72.845 ;
        RECT 81.130 72.680 81.525 73.175 ;
        RECT 72.465 71.715 73.675 72.235 ;
        RECT 74.775 71.935 75.110 72.205 ;
        RECT 70.655 70.805 70.915 71.590 ;
        RECT 71.085 70.625 73.675 71.715 ;
        RECT 74.305 70.625 74.595 71.790 ;
        RECT 75.280 71.775 75.450 72.375 ;
        RECT 75.620 71.935 75.955 72.185 ;
        RECT 76.145 71.885 77.355 72.405 ;
        RECT 74.765 70.625 75.045 71.765 ;
        RECT 75.215 70.795 75.545 71.775 ;
        RECT 75.715 70.625 75.975 71.765 ;
        RECT 77.525 71.715 78.735 72.235 ;
        RECT 76.145 70.625 78.735 71.715 ;
        RECT 79.425 71.645 79.725 72.495 ;
        RECT 79.895 72.455 80.115 72.605 ;
        RECT 79.895 72.125 80.430 72.455 ;
        RECT 80.600 72.315 80.770 72.650 ;
        RECT 81.695 72.485 81.935 73.005 ;
        RECT 79.895 71.475 80.130 72.125 ;
        RECT 80.600 71.955 81.585 72.315 ;
        RECT 79.455 71.245 80.130 71.475 ;
        RECT 80.300 71.935 81.585 71.955 ;
        RECT 80.300 71.785 81.160 71.935 ;
        RECT 79.455 70.815 79.625 71.245 ;
        RECT 79.795 70.625 80.125 71.075 ;
        RECT 80.300 70.840 80.585 71.785 ;
        RECT 81.760 71.680 81.935 72.485 ;
        RECT 82.325 72.545 82.655 72.905 ;
        RECT 83.275 72.715 83.525 73.175 ;
        RECT 83.695 72.715 84.255 73.005 ;
        RECT 82.325 72.355 83.715 72.545 ;
        RECT 83.545 72.265 83.715 72.355 ;
        RECT 80.760 71.305 81.455 71.615 ;
        RECT 80.765 70.625 81.450 71.095 ;
        RECT 81.630 70.895 81.935 71.680 ;
        RECT 82.140 71.935 82.815 72.185 ;
        RECT 83.035 71.935 83.375 72.185 ;
        RECT 83.545 71.935 83.835 72.265 ;
        RECT 82.140 71.575 82.405 71.935 ;
        RECT 83.545 71.685 83.715 71.935 ;
        RECT 82.775 71.515 83.715 71.685 ;
        RECT 82.325 70.625 82.605 71.295 ;
        RECT 82.775 70.965 83.075 71.515 ;
        RECT 84.005 71.345 84.255 72.715 ;
        RECT 84.425 72.405 87.015 73.175 ;
        RECT 87.195 72.675 87.525 73.175 ;
        RECT 87.725 72.605 87.895 72.955 ;
        RECT 88.095 72.775 88.425 73.175 ;
        RECT 88.595 72.605 88.765 72.955 ;
        RECT 88.935 72.775 89.315 73.175 ;
        RECT 84.425 71.885 85.635 72.405 ;
        RECT 85.805 71.715 87.015 72.235 ;
        RECT 87.190 71.935 87.540 72.505 ;
        RECT 87.725 72.435 89.335 72.605 ;
        RECT 89.505 72.500 89.775 72.845 ;
        RECT 89.945 72.630 95.290 73.175 ;
        RECT 96.385 72.795 97.275 72.965 ;
        RECT 89.165 72.265 89.335 72.435 ;
        RECT 83.275 70.625 83.605 71.345 ;
        RECT 83.795 70.795 84.255 71.345 ;
        RECT 84.425 70.625 87.015 71.715 ;
        RECT 87.190 71.475 87.510 71.765 ;
        RECT 87.710 71.645 88.420 72.265 ;
        RECT 88.590 71.935 88.995 72.265 ;
        RECT 89.165 71.935 89.435 72.265 ;
        RECT 89.165 71.765 89.335 71.935 ;
        RECT 89.605 71.765 89.775 72.500 ;
        RECT 91.530 71.800 91.870 72.630 ;
        RECT 88.610 71.595 89.335 71.765 ;
        RECT 88.610 71.475 88.780 71.595 ;
        RECT 87.190 71.305 88.780 71.475 ;
        RECT 87.190 70.845 88.845 71.135 ;
        RECT 89.015 70.625 89.295 71.425 ;
        RECT 89.505 70.795 89.775 71.765 ;
        RECT 93.350 71.060 93.700 72.310 ;
        RECT 96.385 72.240 96.935 72.625 ;
        RECT 97.105 72.070 97.275 72.795 ;
        RECT 96.385 72.000 97.275 72.070 ;
        RECT 97.445 72.470 97.665 72.955 ;
        RECT 97.835 72.635 98.085 73.175 ;
        RECT 98.255 72.525 98.515 73.005 ;
        RECT 97.445 72.045 97.775 72.470 ;
        RECT 96.385 71.975 97.280 72.000 ;
        RECT 96.385 71.960 97.290 71.975 ;
        RECT 96.385 71.945 97.295 71.960 ;
        RECT 96.385 71.940 97.305 71.945 ;
        RECT 96.385 71.930 97.310 71.940 ;
        RECT 96.385 71.920 97.315 71.930 ;
        RECT 96.385 71.915 97.325 71.920 ;
        RECT 96.385 71.905 97.335 71.915 ;
        RECT 96.385 71.900 97.345 71.905 ;
        RECT 96.385 71.450 96.645 71.900 ;
        RECT 97.010 71.895 97.345 71.900 ;
        RECT 97.010 71.890 97.360 71.895 ;
        RECT 97.010 71.880 97.375 71.890 ;
        RECT 97.010 71.875 97.400 71.880 ;
        RECT 97.945 71.875 98.175 72.270 ;
        RECT 97.010 71.870 98.175 71.875 ;
        RECT 97.040 71.835 98.175 71.870 ;
        RECT 97.075 71.810 98.175 71.835 ;
        RECT 97.105 71.780 98.175 71.810 ;
        RECT 97.125 71.750 98.175 71.780 ;
        RECT 97.145 71.720 98.175 71.750 ;
        RECT 97.215 71.710 98.175 71.720 ;
        RECT 97.240 71.700 98.175 71.710 ;
        RECT 97.260 71.685 98.175 71.700 ;
        RECT 97.280 71.670 98.175 71.685 ;
        RECT 97.285 71.660 98.070 71.670 ;
        RECT 97.300 71.625 98.070 71.660 ;
        RECT 96.815 71.305 97.145 71.550 ;
        RECT 97.315 71.375 98.070 71.625 ;
        RECT 98.345 71.495 98.515 72.525 ;
        RECT 98.775 72.625 98.945 73.005 ;
        RECT 99.125 72.795 99.455 73.175 ;
        RECT 98.775 72.455 99.440 72.625 ;
        RECT 99.635 72.500 99.895 73.005 ;
        RECT 98.705 71.905 99.035 72.275 ;
        RECT 99.270 72.200 99.440 72.455 ;
        RECT 99.270 71.870 99.555 72.200 ;
        RECT 99.270 71.725 99.440 71.870 ;
        RECT 96.815 71.280 97.000 71.305 ;
        RECT 96.385 71.180 97.000 71.280 ;
        RECT 89.945 70.625 95.290 71.060 ;
        RECT 96.385 70.625 96.990 71.180 ;
        RECT 97.165 70.795 97.645 71.135 ;
        RECT 97.815 70.625 98.070 71.170 ;
        RECT 98.240 70.795 98.515 71.495 ;
        RECT 98.775 71.555 99.440 71.725 ;
        RECT 99.725 71.700 99.895 72.500 ;
        RECT 100.065 72.450 100.355 73.175 ;
        RECT 101.535 72.625 101.705 73.005 ;
        RECT 101.885 72.795 102.215 73.175 ;
        RECT 101.535 72.455 102.200 72.625 ;
        RECT 102.395 72.500 102.655 73.005 ;
        RECT 103.005 72.515 103.345 73.175 ;
        RECT 101.465 71.905 101.795 72.275 ;
        RECT 102.030 72.200 102.200 72.455 ;
        RECT 102.030 71.870 102.315 72.200 ;
        RECT 98.775 70.795 98.945 71.555 ;
        RECT 99.125 70.625 99.455 71.385 ;
        RECT 99.625 70.795 99.895 71.700 ;
        RECT 100.065 70.625 100.355 71.790 ;
        RECT 102.030 71.725 102.200 71.870 ;
        RECT 101.535 71.555 102.200 71.725 ;
        RECT 102.485 71.700 102.655 72.500 ;
        RECT 101.535 70.795 101.705 71.555 ;
        RECT 101.885 70.625 102.215 71.385 ;
        RECT 102.385 70.795 102.655 71.700 ;
        RECT 102.825 70.795 103.345 72.345 ;
        RECT 103.515 71.520 104.035 73.005 ;
        RECT 104.205 72.405 107.715 73.175 ;
        RECT 108.805 72.675 109.065 73.005 ;
        RECT 109.275 72.695 109.550 73.175 ;
        RECT 104.205 71.885 105.855 72.405 ;
        RECT 106.025 71.715 107.715 72.235 ;
        RECT 103.515 70.625 103.845 71.350 ;
        RECT 104.205 70.625 107.715 71.715 ;
        RECT 108.805 71.765 108.975 72.675 ;
        RECT 109.760 72.605 109.965 73.005 ;
        RECT 110.135 72.775 110.470 73.175 ;
        RECT 110.645 72.675 110.905 73.005 ;
        RECT 111.115 72.695 111.390 73.175 ;
        RECT 109.145 71.935 109.505 72.515 ;
        RECT 109.760 72.435 110.445 72.605 ;
        RECT 109.685 71.765 109.935 72.265 ;
        RECT 108.805 71.595 109.935 71.765 ;
        RECT 108.805 70.825 109.075 71.595 ;
        RECT 110.105 71.405 110.445 72.435 ;
        RECT 109.245 70.625 109.575 71.405 ;
        RECT 109.780 71.230 110.445 71.405 ;
        RECT 110.645 71.765 110.815 72.675 ;
        RECT 111.600 72.605 111.805 73.005 ;
        RECT 111.975 72.775 112.310 73.175 ;
        RECT 110.985 71.935 111.345 72.515 ;
        RECT 111.600 72.435 112.285 72.605 ;
        RECT 111.525 71.765 111.775 72.265 ;
        RECT 110.645 71.595 111.775 71.765 ;
        RECT 109.780 70.825 109.965 71.230 ;
        RECT 110.135 70.625 110.470 71.050 ;
        RECT 110.645 70.825 110.915 71.595 ;
        RECT 111.945 71.405 112.285 72.435 ;
        RECT 112.485 72.425 113.695 73.175 ;
        RECT 112.485 71.885 113.005 72.425 ;
        RECT 113.865 72.375 114.175 73.175 ;
        RECT 114.380 72.375 115.075 73.005 ;
        RECT 115.245 72.405 116.915 73.175 ;
        RECT 117.550 72.670 117.885 73.175 ;
        RECT 118.055 72.605 118.295 72.980 ;
        RECT 118.575 72.845 118.745 72.990 ;
        RECT 118.575 72.650 118.950 72.845 ;
        RECT 119.310 72.680 119.705 73.175 ;
        RECT 113.175 71.715 113.695 72.255 ;
        RECT 113.875 71.935 114.210 72.205 ;
        RECT 114.380 71.775 114.550 72.375 ;
        RECT 114.720 71.935 115.055 72.185 ;
        RECT 115.245 71.885 115.995 72.405 ;
        RECT 111.085 70.625 111.415 71.405 ;
        RECT 111.620 71.230 112.285 71.405 ;
        RECT 111.620 70.825 111.805 71.230 ;
        RECT 111.975 70.625 112.310 71.050 ;
        RECT 112.485 70.625 113.695 71.715 ;
        RECT 113.865 70.625 114.145 71.765 ;
        RECT 114.315 70.795 114.645 71.775 ;
        RECT 114.815 70.625 115.075 71.765 ;
        RECT 116.165 71.715 116.915 72.235 ;
        RECT 115.245 70.625 116.915 71.715 ;
        RECT 117.605 71.645 117.905 72.495 ;
        RECT 118.075 72.455 118.295 72.605 ;
        RECT 118.075 72.125 118.610 72.455 ;
        RECT 118.780 72.315 118.950 72.650 ;
        RECT 119.875 72.485 120.115 73.005 ;
        RECT 118.075 71.475 118.310 72.125 ;
        RECT 118.780 71.955 119.765 72.315 ;
        RECT 117.635 71.245 118.310 71.475 ;
        RECT 118.480 71.935 119.765 71.955 ;
        RECT 118.480 71.785 119.340 71.935 ;
        RECT 117.635 70.815 117.805 71.245 ;
        RECT 117.975 70.625 118.305 71.075 ;
        RECT 118.480 70.840 118.765 71.785 ;
        RECT 119.940 71.680 120.115 72.485 ;
        RECT 118.940 71.305 119.635 71.615 ;
        RECT 118.945 70.625 119.630 71.095 ;
        RECT 119.810 70.895 120.115 71.680 ;
        RECT 120.330 72.420 120.565 72.750 ;
        RECT 120.735 72.435 121.065 73.175 ;
        RECT 121.300 72.795 122.495 73.005 ;
        RECT 120.330 71.765 120.500 72.420 ;
        RECT 121.300 72.355 121.575 72.795 ;
        RECT 121.745 72.455 122.075 72.625 ;
        RECT 121.750 72.355 122.075 72.455 ;
        RECT 122.245 72.565 122.495 72.795 ;
        RECT 122.665 72.735 122.835 73.175 ;
        RECT 123.005 72.565 123.355 73.005 ;
        RECT 122.245 72.355 123.355 72.565 ;
        RECT 123.545 72.365 123.785 73.175 ;
        RECT 123.955 72.365 124.285 73.005 ;
        RECT 124.455 72.365 124.725 73.175 ;
        RECT 125.825 72.450 126.115 73.175 ;
        RECT 126.755 72.675 127.085 73.175 ;
        RECT 127.285 72.605 127.455 72.955 ;
        RECT 127.655 72.775 127.985 73.175 ;
        RECT 128.155 72.605 128.325 72.955 ;
        RECT 128.495 72.775 128.875 73.175 ;
        RECT 120.675 71.935 121.020 72.265 ;
        RECT 121.250 71.765 121.580 72.185 ;
        RECT 120.330 71.595 121.580 71.765 ;
        RECT 120.330 71.400 120.630 71.595 ;
        RECT 121.750 71.425 122.030 72.355 ;
        RECT 122.210 71.985 123.355 72.185 ;
        RECT 122.210 71.605 122.400 71.985 ;
        RECT 123.525 71.935 123.875 72.185 ;
        RECT 124.045 71.765 124.215 72.365 ;
        RECT 124.385 71.935 124.735 72.185 ;
        RECT 126.750 71.935 127.100 72.505 ;
        RECT 127.285 72.435 128.895 72.605 ;
        RECT 129.065 72.500 129.335 72.845 ;
        RECT 129.505 72.630 134.850 73.175 ;
        RECT 128.725 72.265 128.895 72.435 ;
        RECT 122.580 71.425 122.855 71.765 ;
        RECT 120.800 70.625 121.055 71.425 ;
        RECT 121.255 71.255 122.855 71.425 ;
        RECT 121.255 70.795 121.585 71.255 ;
        RECT 121.755 70.625 122.330 71.085 ;
        RECT 122.500 70.795 122.855 71.255 ;
        RECT 123.025 70.625 123.355 71.765 ;
        RECT 123.535 71.595 124.215 71.765 ;
        RECT 123.535 70.810 123.865 71.595 ;
        RECT 124.395 70.625 124.725 71.765 ;
        RECT 125.825 70.625 126.115 71.790 ;
        RECT 126.750 71.475 127.070 71.765 ;
        RECT 127.270 71.645 127.980 72.265 ;
        RECT 128.150 71.935 128.555 72.265 ;
        RECT 128.725 71.935 128.995 72.265 ;
        RECT 128.725 71.765 128.895 71.935 ;
        RECT 129.165 71.765 129.335 72.500 ;
        RECT 131.090 71.800 131.430 72.630 ;
        RECT 135.025 72.425 136.235 73.175 ;
        RECT 136.605 72.545 136.935 72.905 ;
        RECT 137.555 72.715 137.805 73.175 ;
        RECT 137.975 72.715 138.535 73.005 ;
        RECT 138.705 72.795 139.595 72.965 ;
        RECT 128.170 71.595 128.895 71.765 ;
        RECT 128.170 71.475 128.340 71.595 ;
        RECT 126.750 71.305 128.340 71.475 ;
        RECT 126.750 70.845 128.405 71.135 ;
        RECT 128.575 70.625 128.855 71.425 ;
        RECT 129.065 70.795 129.335 71.765 ;
        RECT 132.910 71.060 133.260 72.310 ;
        RECT 135.025 71.885 135.545 72.425 ;
        RECT 136.605 72.355 137.995 72.545 ;
        RECT 137.825 72.265 137.995 72.355 ;
        RECT 135.715 71.715 136.235 72.255 ;
        RECT 129.505 70.625 134.850 71.060 ;
        RECT 135.025 70.625 136.235 71.715 ;
        RECT 136.420 71.935 137.095 72.185 ;
        RECT 137.315 71.935 137.655 72.185 ;
        RECT 137.825 71.935 138.115 72.265 ;
        RECT 136.420 71.575 136.685 71.935 ;
        RECT 137.825 71.685 137.995 71.935 ;
        RECT 137.055 71.515 137.995 71.685 ;
        RECT 136.605 70.625 136.885 71.295 ;
        RECT 137.055 70.965 137.355 71.515 ;
        RECT 138.285 71.345 138.535 72.715 ;
        RECT 138.705 72.240 139.255 72.625 ;
        RECT 139.425 72.070 139.595 72.795 ;
        RECT 138.705 72.000 139.595 72.070 ;
        RECT 139.765 72.470 139.985 72.955 ;
        RECT 140.155 72.635 140.405 73.175 ;
        RECT 140.575 72.525 140.835 73.005 ;
        RECT 139.765 72.045 140.095 72.470 ;
        RECT 138.705 71.975 139.600 72.000 ;
        RECT 138.705 71.960 139.610 71.975 ;
        RECT 138.705 71.945 139.615 71.960 ;
        RECT 138.705 71.940 139.625 71.945 ;
        RECT 138.705 71.930 139.630 71.940 ;
        RECT 138.705 71.920 139.635 71.930 ;
        RECT 138.705 71.915 139.645 71.920 ;
        RECT 138.705 71.905 139.655 71.915 ;
        RECT 138.705 71.900 139.665 71.905 ;
        RECT 138.705 71.450 138.965 71.900 ;
        RECT 139.330 71.895 139.665 71.900 ;
        RECT 139.330 71.890 139.680 71.895 ;
        RECT 139.330 71.880 139.695 71.890 ;
        RECT 139.330 71.875 139.720 71.880 ;
        RECT 140.265 71.875 140.495 72.270 ;
        RECT 139.330 71.870 140.495 71.875 ;
        RECT 139.360 71.835 140.495 71.870 ;
        RECT 139.395 71.810 140.495 71.835 ;
        RECT 139.425 71.780 140.495 71.810 ;
        RECT 139.445 71.750 140.495 71.780 ;
        RECT 139.465 71.720 140.495 71.750 ;
        RECT 139.535 71.710 140.495 71.720 ;
        RECT 139.560 71.700 140.495 71.710 ;
        RECT 139.580 71.685 140.495 71.700 ;
        RECT 139.600 71.670 140.495 71.685 ;
        RECT 139.605 71.660 140.390 71.670 ;
        RECT 139.620 71.625 140.390 71.660 ;
        RECT 137.555 70.625 137.885 71.345 ;
        RECT 138.075 70.795 138.535 71.345 ;
        RECT 139.135 71.305 139.465 71.550 ;
        RECT 139.635 71.375 140.390 71.625 ;
        RECT 140.665 71.495 140.835 72.525 ;
        RECT 141.005 71.520 141.525 73.005 ;
        RECT 141.695 72.515 142.035 73.175 ;
        RECT 142.475 72.625 142.645 72.915 ;
        RECT 142.815 72.795 143.145 73.175 ;
        RECT 142.475 72.455 143.080 72.625 ;
        RECT 139.135 71.280 139.320 71.305 ;
        RECT 138.705 71.180 139.320 71.280 ;
        RECT 138.705 70.625 139.310 71.180 ;
        RECT 139.485 70.795 139.965 71.135 ;
        RECT 140.135 70.625 140.390 71.170 ;
        RECT 140.560 70.795 140.835 71.495 ;
        RECT 141.195 70.625 141.525 71.350 ;
        RECT 141.695 70.795 142.215 72.345 ;
        RECT 142.385 71.635 142.630 72.275 ;
        RECT 142.910 72.190 143.080 72.455 ;
        RECT 142.910 71.860 143.140 72.190 ;
        RECT 142.910 71.465 143.080 71.860 ;
        RECT 142.475 71.295 143.080 71.465 ;
        RECT 143.315 71.575 143.485 72.915 ;
        RECT 143.810 72.645 144.005 72.915 ;
        RECT 144.175 72.815 144.505 73.175 ;
        RECT 145.065 72.725 145.905 72.895 ;
        RECT 143.810 72.495 144.415 72.645 ;
        RECT 143.810 72.475 144.620 72.495 ;
        RECT 143.735 71.935 144.065 72.305 ;
        RECT 144.245 72.025 144.620 72.475 ;
        RECT 144.860 72.220 145.565 72.525 ;
        RECT 144.245 71.765 144.415 72.025 ;
        RECT 143.730 71.595 144.415 71.765 ;
        RECT 142.475 70.795 142.645 71.295 ;
        RECT 142.815 70.625 143.145 71.125 ;
        RECT 143.315 70.795 143.540 71.575 ;
        RECT 143.730 70.845 144.085 71.595 ;
        RECT 144.255 70.625 144.545 71.425 ;
        RECT 144.745 71.255 145.080 71.905 ;
        RECT 145.250 71.700 145.565 72.220 ;
        RECT 145.735 72.265 145.905 72.725 ;
        RECT 146.075 72.715 146.345 73.175 ;
        RECT 146.595 72.540 146.840 73.000 ;
        RECT 147.055 72.545 147.280 73.175 ;
        RECT 146.670 72.265 146.840 72.540 ;
        RECT 147.475 72.515 147.735 72.845 ;
        RECT 145.735 71.935 146.500 72.265 ;
        RECT 146.670 71.935 147.395 72.265 ;
        RECT 145.735 71.810 145.945 71.935 ;
        RECT 145.250 71.350 145.585 71.700 ;
        RECT 145.755 71.250 145.945 71.810 ;
        RECT 146.670 71.725 146.840 71.935 ;
        RECT 146.115 71.395 146.840 71.725 ;
        RECT 145.730 71.225 145.945 71.250 ;
        RECT 145.705 71.215 145.945 71.225 ;
        RECT 145.690 71.195 145.945 71.215 ;
        RECT 145.690 71.175 145.930 71.195 ;
        RECT 145.690 71.170 145.920 71.175 ;
        RECT 145.595 71.155 145.920 71.170 ;
        RECT 145.595 71.005 145.905 71.155 ;
        RECT 145.045 70.835 145.905 71.005 ;
        RECT 146.075 70.625 146.395 71.085 ;
        RECT 146.595 70.825 146.840 71.395 ;
        RECT 147.020 70.625 147.305 71.690 ;
        RECT 147.565 71.590 147.735 72.515 ;
        RECT 147.905 72.405 151.415 73.175 ;
        RECT 151.585 72.450 151.875 73.175 ;
        RECT 152.045 72.405 155.555 73.175 ;
        RECT 155.725 72.425 156.935 73.175 ;
        RECT 147.905 71.885 149.555 72.405 ;
        RECT 149.725 71.715 151.415 72.235 ;
        RECT 152.045 71.885 153.695 72.405 ;
        RECT 147.475 70.805 147.735 71.590 ;
        RECT 147.905 70.625 151.415 71.715 ;
        RECT 151.585 70.625 151.875 71.790 ;
        RECT 153.865 71.715 155.555 72.235 ;
        RECT 152.045 70.625 155.555 71.715 ;
        RECT 155.725 71.715 156.245 72.255 ;
        RECT 156.415 71.885 156.935 72.425 ;
        RECT 155.725 70.625 156.935 71.715 ;
        RECT 22.700 70.455 157.020 70.625 ;
        RECT 22.785 69.365 23.995 70.455 ;
        RECT 24.165 70.020 29.510 70.455 ;
        RECT 29.685 70.020 35.030 70.455 ;
        RECT 22.785 68.655 23.305 69.195 ;
        RECT 23.475 68.825 23.995 69.365 ;
        RECT 22.785 67.905 23.995 68.655 ;
        RECT 25.750 68.450 26.090 69.280 ;
        RECT 27.570 68.770 27.920 70.020 ;
        RECT 31.270 68.450 31.610 69.280 ;
        RECT 33.090 68.770 33.440 70.020 ;
        RECT 35.665 69.290 35.955 70.455 ;
        RECT 36.595 69.315 36.925 70.455 ;
        RECT 37.455 69.485 37.785 70.270 ;
        RECT 37.105 69.315 37.785 69.485 ;
        RECT 37.965 69.365 39.635 70.455 ;
        RECT 40.265 69.945 41.455 70.235 ;
        RECT 36.585 68.895 36.935 69.145 ;
        RECT 37.105 68.715 37.275 69.315 ;
        RECT 37.445 68.895 37.795 69.145 ;
        RECT 24.165 67.905 29.510 68.450 ;
        RECT 29.685 67.905 35.030 68.450 ;
        RECT 35.665 67.905 35.955 68.630 ;
        RECT 36.595 67.905 36.865 68.715 ;
        RECT 37.035 68.075 37.365 68.715 ;
        RECT 37.535 67.905 37.775 68.715 ;
        RECT 37.965 68.675 38.715 69.195 ;
        RECT 38.885 68.845 39.635 69.365 ;
        RECT 40.285 69.605 41.455 69.775 ;
        RECT 41.625 69.655 41.905 70.455 ;
        RECT 40.285 69.315 40.610 69.605 ;
        RECT 41.285 69.485 41.455 69.605 ;
        RECT 40.780 69.145 40.975 69.435 ;
        RECT 41.285 69.315 41.945 69.485 ;
        RECT 42.115 69.315 42.390 70.285 ;
        RECT 41.775 69.145 41.945 69.315 ;
        RECT 40.265 68.815 40.610 69.145 ;
        RECT 40.780 68.815 41.605 69.145 ;
        RECT 41.775 68.815 42.050 69.145 ;
        RECT 37.965 67.905 39.635 68.675 ;
        RECT 41.775 68.645 41.945 68.815 ;
        RECT 40.280 68.475 41.945 68.645 ;
        RECT 42.220 68.580 42.390 69.315 ;
        RECT 40.280 68.125 40.535 68.475 ;
        RECT 40.705 67.905 41.035 68.305 ;
        RECT 41.205 68.125 41.375 68.475 ;
        RECT 41.545 67.905 41.925 68.305 ;
        RECT 42.115 68.235 42.390 68.580 ;
        RECT 42.570 69.505 42.835 70.275 ;
        RECT 43.005 69.735 43.335 70.455 ;
        RECT 43.525 69.915 43.785 70.275 ;
        RECT 43.955 70.085 44.285 70.455 ;
        RECT 44.455 69.915 44.715 70.275 ;
        RECT 43.525 69.685 44.715 69.915 ;
        RECT 45.285 69.505 45.575 70.275 ;
        RECT 42.570 68.085 42.905 69.505 ;
        RECT 43.080 69.325 45.575 69.505 ;
        RECT 45.795 69.485 46.125 70.270 ;
        RECT 43.080 68.635 43.305 69.325 ;
        RECT 45.795 69.315 46.475 69.485 ;
        RECT 46.655 69.315 46.985 70.455 ;
        RECT 47.165 69.315 47.495 70.455 ;
        RECT 47.665 69.825 48.020 70.285 ;
        RECT 48.190 69.995 48.765 70.455 ;
        RECT 48.935 69.825 49.265 70.285 ;
        RECT 47.665 69.655 49.265 69.825 ;
        RECT 49.465 69.655 49.720 70.455 ;
        RECT 51.805 69.995 52.020 70.455 ;
        RECT 52.190 69.825 52.520 70.285 ;
        RECT 47.665 69.315 47.940 69.655 ;
        RECT 43.505 68.815 43.785 69.145 ;
        RECT 43.965 68.815 44.540 69.145 ;
        RECT 44.720 68.815 45.155 69.145 ;
        RECT 45.335 68.815 45.605 69.145 ;
        RECT 45.785 68.895 46.135 69.145 ;
        RECT 46.305 68.715 46.475 69.315 ;
        RECT 46.645 68.895 46.995 69.145 ;
        RECT 48.120 69.095 48.310 69.475 ;
        RECT 47.165 68.925 48.315 69.095 ;
        RECT 47.165 68.895 48.310 68.925 ;
        RECT 48.490 68.725 48.770 69.655 ;
        RECT 49.890 69.485 50.190 69.680 ;
        RECT 48.940 69.315 50.190 69.485 ;
        RECT 48.940 68.895 49.270 69.315 ;
        RECT 49.500 68.815 49.845 69.145 ;
        RECT 43.080 68.445 45.565 68.635 ;
        RECT 43.085 67.905 43.830 68.275 ;
        RECT 44.395 68.085 44.650 68.445 ;
        RECT 44.830 67.905 45.160 68.275 ;
        RECT 45.340 68.085 45.565 68.445 ;
        RECT 45.805 67.905 46.045 68.715 ;
        RECT 46.215 68.075 46.545 68.715 ;
        RECT 46.715 67.905 46.985 68.715 ;
        RECT 47.165 68.515 48.275 68.725 ;
        RECT 47.165 68.075 47.515 68.515 ;
        RECT 47.685 67.905 47.855 68.345 ;
        RECT 48.025 68.285 48.275 68.515 ;
        RECT 48.445 68.625 48.770 68.725 ;
        RECT 48.445 68.455 48.775 68.625 ;
        RECT 48.945 68.285 49.220 68.725 ;
        RECT 50.020 68.660 50.190 69.315 ;
        RECT 48.025 68.075 49.220 68.285 ;
        RECT 49.455 67.905 49.785 68.645 ;
        RECT 49.955 68.330 50.190 68.660 ;
        RECT 51.350 69.655 52.520 69.825 ;
        RECT 52.690 69.655 52.940 70.455 ;
        RECT 51.350 68.365 51.720 69.655 ;
        RECT 53.150 69.485 53.430 69.645 ;
        RECT 52.095 69.315 53.430 69.485 ;
        RECT 53.615 69.485 53.945 70.270 ;
        RECT 53.615 69.315 54.295 69.485 ;
        RECT 54.475 69.315 54.805 70.455 ;
        RECT 54.985 69.365 58.495 70.455 ;
        RECT 52.095 69.145 52.265 69.315 ;
        RECT 51.890 68.895 52.265 69.145 ;
        RECT 52.435 68.895 52.910 69.135 ;
        RECT 53.080 68.895 53.430 69.135 ;
        RECT 53.605 68.895 53.955 69.145 ;
        RECT 52.095 68.725 52.265 68.895 ;
        RECT 52.095 68.555 53.430 68.725 ;
        RECT 54.125 68.715 54.295 69.315 ;
        RECT 54.465 68.895 54.815 69.145 ;
        RECT 51.350 68.075 52.100 68.365 ;
        RECT 52.610 67.905 52.940 68.365 ;
        RECT 53.160 68.345 53.430 68.555 ;
        RECT 53.625 67.905 53.865 68.715 ;
        RECT 54.035 68.075 54.365 68.715 ;
        RECT 54.535 67.905 54.805 68.715 ;
        RECT 54.985 68.675 56.635 69.195 ;
        RECT 56.805 68.845 58.495 69.365 ;
        RECT 59.125 69.315 59.385 70.455 ;
        RECT 59.555 69.305 59.885 70.285 ;
        RECT 60.055 69.315 60.335 70.455 ;
        RECT 59.145 68.895 59.480 69.145 ;
        RECT 59.650 68.705 59.820 69.305 ;
        RECT 61.425 69.290 61.715 70.455 ;
        RECT 59.990 68.875 60.325 69.145 ;
        RECT 61.885 68.735 62.405 70.285 ;
        RECT 62.575 69.730 62.905 70.455 ;
        RECT 54.985 67.905 58.495 68.675 ;
        RECT 59.125 68.075 59.820 68.705 ;
        RECT 60.025 67.905 60.335 68.705 ;
        RECT 61.425 67.905 61.715 68.630 ;
        RECT 62.065 67.905 62.405 68.565 ;
        RECT 62.575 68.075 63.095 69.560 ;
        RECT 63.265 69.365 66.775 70.455 ;
        RECT 63.265 68.675 64.915 69.195 ;
        RECT 65.085 68.845 66.775 69.365 ;
        RECT 67.900 69.665 68.435 70.285 ;
        RECT 63.265 67.905 66.775 68.675 ;
        RECT 67.900 68.645 68.215 69.665 ;
        RECT 68.605 69.655 68.935 70.455 ;
        RECT 69.420 69.485 69.810 69.660 ;
        RECT 68.385 69.315 69.810 69.485 ;
        RECT 70.165 69.315 70.435 70.285 ;
        RECT 70.645 69.655 70.925 70.455 ;
        RECT 71.105 69.905 72.300 70.235 ;
        RECT 71.430 69.485 71.850 69.735 ;
        RECT 70.605 69.315 71.850 69.485 ;
        RECT 68.385 68.815 68.555 69.315 ;
        RECT 67.900 68.075 68.515 68.645 ;
        RECT 68.805 68.585 69.070 69.145 ;
        RECT 69.240 68.415 69.410 69.315 ;
        RECT 69.580 68.585 69.935 69.145 ;
        RECT 70.165 68.580 70.335 69.315 ;
        RECT 70.605 69.145 70.775 69.315 ;
        RECT 72.075 69.145 72.245 69.705 ;
        RECT 72.495 69.315 72.750 70.455 ;
        RECT 73.420 69.655 73.670 70.455 ;
        RECT 73.840 69.825 74.170 70.285 ;
        RECT 74.340 69.995 74.555 70.455 ;
        RECT 73.840 69.655 75.010 69.825 ;
        RECT 72.930 69.485 73.210 69.645 ;
        RECT 72.930 69.315 74.265 69.485 ;
        RECT 74.095 69.145 74.265 69.315 ;
        RECT 70.545 68.815 70.775 69.145 ;
        RECT 71.505 68.815 72.245 69.145 ;
        RECT 72.415 68.895 72.750 69.145 ;
        RECT 72.930 68.895 73.280 69.135 ;
        RECT 73.450 68.895 73.925 69.135 ;
        RECT 74.095 68.895 74.470 69.145 ;
        RECT 70.605 68.645 70.775 68.815 ;
        RECT 71.995 68.725 72.245 68.815 ;
        RECT 74.095 68.725 74.265 68.895 ;
        RECT 68.685 67.905 68.900 68.415 ;
        RECT 69.130 68.085 69.410 68.415 ;
        RECT 69.590 67.905 69.830 68.415 ;
        RECT 70.165 68.235 70.435 68.580 ;
        RECT 70.605 68.475 71.345 68.645 ;
        RECT 71.995 68.555 72.730 68.725 ;
        RECT 70.625 67.905 71.005 68.305 ;
        RECT 71.175 68.125 71.345 68.475 ;
        RECT 71.515 67.905 72.250 68.385 ;
        RECT 72.420 68.085 72.730 68.555 ;
        RECT 72.930 68.555 74.265 68.725 ;
        RECT 72.930 68.345 73.200 68.555 ;
        RECT 74.640 68.365 75.010 69.655 ;
        RECT 75.225 69.365 76.895 70.455 ;
        RECT 73.420 67.905 73.750 68.365 ;
        RECT 74.260 68.075 75.010 68.365 ;
        RECT 75.225 68.675 75.975 69.195 ;
        RECT 76.145 68.845 76.895 69.365 ;
        RECT 77.525 69.315 77.855 70.455 ;
        RECT 78.025 69.825 78.380 70.285 ;
        RECT 78.550 69.995 79.125 70.455 ;
        RECT 79.295 69.825 79.625 70.285 ;
        RECT 78.025 69.655 79.625 69.825 ;
        RECT 79.825 69.655 80.080 70.455 ;
        RECT 78.025 69.315 78.300 69.655 ;
        RECT 78.480 69.095 78.670 69.475 ;
        RECT 77.525 68.895 78.670 69.095 ;
        RECT 78.850 68.755 79.130 69.655 ;
        RECT 80.250 69.485 80.550 69.680 ;
        RECT 79.300 69.315 80.550 69.485 ;
        RECT 80.745 69.365 81.955 70.455 ;
        RECT 79.300 68.895 79.630 69.315 ;
        RECT 79.860 68.815 80.205 69.145 ;
        RECT 78.850 68.725 79.135 68.755 ;
        RECT 75.225 67.905 76.895 68.675 ;
        RECT 77.525 68.515 78.635 68.725 ;
        RECT 77.525 68.075 77.875 68.515 ;
        RECT 78.045 67.905 78.215 68.345 ;
        RECT 78.385 68.285 78.635 68.515 ;
        RECT 78.805 68.455 79.135 68.725 ;
        RECT 79.305 68.285 79.580 68.725 ;
        RECT 80.380 68.660 80.550 69.315 ;
        RECT 78.385 68.075 79.580 68.285 ;
        RECT 79.815 67.905 80.145 68.645 ;
        RECT 80.315 68.330 80.550 68.660 ;
        RECT 80.745 68.655 81.265 69.195 ;
        RECT 81.435 68.825 81.955 69.365 ;
        RECT 82.130 69.315 82.450 70.455 ;
        RECT 82.630 69.145 82.825 70.195 ;
        RECT 83.005 69.605 83.335 70.285 ;
        RECT 83.535 69.655 83.790 70.455 ;
        RECT 83.005 69.325 83.355 69.605 ;
        RECT 83.975 69.485 84.305 70.270 ;
        RECT 82.190 69.095 82.450 69.145 ;
        RECT 82.185 68.925 82.450 69.095 ;
        RECT 82.190 68.815 82.450 68.925 ;
        RECT 82.630 68.815 83.015 69.145 ;
        RECT 83.185 68.945 83.355 69.325 ;
        RECT 83.545 69.115 83.790 69.475 ;
        RECT 83.975 69.315 84.655 69.485 ;
        RECT 84.835 69.315 85.165 70.455 ;
        RECT 85.815 69.315 86.145 70.455 ;
        RECT 86.675 69.485 87.005 70.270 ;
        RECT 86.325 69.315 87.005 69.485 ;
        RECT 83.185 68.775 83.705 68.945 ;
        RECT 83.965 68.895 84.315 69.145 ;
        RECT 80.745 67.905 81.955 68.655 ;
        RECT 82.130 68.435 83.345 68.605 ;
        RECT 82.130 68.085 82.420 68.435 ;
        RECT 82.615 67.905 82.945 68.265 ;
        RECT 83.115 68.130 83.345 68.435 ;
        RECT 83.535 68.415 83.705 68.775 ;
        RECT 84.485 68.715 84.655 69.315 ;
        RECT 84.825 68.895 85.175 69.145 ;
        RECT 85.805 68.895 86.155 69.145 ;
        RECT 86.325 68.715 86.495 69.315 ;
        RECT 87.185 69.290 87.475 70.455 ;
        RECT 87.655 69.315 87.985 70.455 ;
        RECT 88.515 69.485 88.845 70.270 ;
        RECT 89.525 69.995 89.740 70.455 ;
        RECT 89.910 69.825 90.240 70.285 ;
        RECT 88.165 69.315 88.845 69.485 ;
        RECT 89.070 69.655 90.240 69.825 ;
        RECT 90.410 69.655 90.660 70.455 ;
        RECT 86.665 68.895 87.015 69.145 ;
        RECT 87.645 68.895 87.995 69.145 ;
        RECT 88.165 68.715 88.335 69.315 ;
        RECT 88.505 68.895 88.855 69.145 ;
        RECT 83.535 68.245 83.735 68.415 ;
        RECT 83.535 68.210 83.705 68.245 ;
        RECT 83.985 67.905 84.225 68.715 ;
        RECT 84.395 68.075 84.725 68.715 ;
        RECT 84.895 67.905 85.165 68.715 ;
        RECT 85.815 67.905 86.085 68.715 ;
        RECT 86.255 68.075 86.585 68.715 ;
        RECT 86.755 67.905 86.995 68.715 ;
        RECT 87.185 67.905 87.475 68.630 ;
        RECT 87.655 67.905 87.925 68.715 ;
        RECT 88.095 68.075 88.425 68.715 ;
        RECT 88.595 67.905 88.835 68.715 ;
        RECT 89.070 68.365 89.440 69.655 ;
        RECT 90.870 69.485 91.150 69.645 ;
        RECT 89.815 69.315 91.150 69.485 ;
        RECT 91.335 69.485 91.665 70.270 ;
        RECT 91.335 69.315 92.015 69.485 ;
        RECT 92.195 69.315 92.525 70.455 ;
        RECT 93.625 69.945 93.885 70.455 ;
        RECT 89.815 69.145 89.985 69.315 ;
        RECT 89.610 68.895 89.985 69.145 ;
        RECT 90.155 68.895 90.630 69.135 ;
        RECT 90.800 68.895 91.150 69.135 ;
        RECT 91.325 68.895 91.675 69.145 ;
        RECT 89.815 68.725 89.985 68.895 ;
        RECT 89.815 68.555 91.150 68.725 ;
        RECT 91.845 68.715 92.015 69.315 ;
        RECT 92.185 68.895 92.535 69.145 ;
        RECT 93.625 68.895 93.965 69.775 ;
        RECT 94.135 69.065 94.305 70.285 ;
        RECT 94.545 69.950 95.160 70.455 ;
        RECT 94.545 69.415 94.795 69.780 ;
        RECT 94.965 69.775 95.160 69.950 ;
        RECT 95.330 69.945 95.805 70.285 ;
        RECT 95.975 69.910 96.190 70.455 ;
        RECT 94.965 69.585 95.295 69.775 ;
        RECT 95.515 69.415 96.230 69.710 ;
        RECT 96.400 69.585 96.675 70.285 ;
        RECT 96.845 69.945 97.105 70.455 ;
        RECT 94.545 69.245 96.335 69.415 ;
        RECT 94.135 68.815 94.930 69.065 ;
        RECT 94.135 68.725 94.385 68.815 ;
        RECT 89.070 68.075 89.820 68.365 ;
        RECT 90.330 67.905 90.660 68.365 ;
        RECT 90.880 68.345 91.150 68.555 ;
        RECT 91.345 67.905 91.585 68.715 ;
        RECT 91.755 68.075 92.085 68.715 ;
        RECT 92.255 67.905 92.525 68.715 ;
        RECT 93.625 67.905 93.885 68.725 ;
        RECT 94.055 68.305 94.385 68.725 ;
        RECT 95.100 68.390 95.355 69.245 ;
        RECT 94.565 68.125 95.355 68.390 ;
        RECT 95.525 68.545 95.935 69.065 ;
        RECT 96.105 68.815 96.335 69.245 ;
        RECT 96.505 68.555 96.675 69.585 ;
        RECT 96.845 68.895 97.185 69.775 ;
        RECT 97.355 69.065 97.525 70.285 ;
        RECT 97.765 69.950 98.380 70.455 ;
        RECT 97.765 69.415 98.015 69.780 ;
        RECT 98.185 69.775 98.380 69.950 ;
        RECT 98.550 69.945 99.025 70.285 ;
        RECT 99.195 69.910 99.410 70.455 ;
        RECT 98.185 69.585 98.515 69.775 ;
        RECT 98.735 69.415 99.450 69.710 ;
        RECT 99.620 69.585 99.895 70.285 ;
        RECT 97.765 69.245 99.555 69.415 ;
        RECT 97.355 68.815 98.150 69.065 ;
        RECT 97.355 68.725 97.605 68.815 ;
        RECT 95.525 68.125 95.725 68.545 ;
        RECT 95.915 67.905 96.245 68.365 ;
        RECT 96.415 68.075 96.675 68.555 ;
        RECT 96.845 67.905 97.105 68.725 ;
        RECT 97.275 68.305 97.605 68.725 ;
        RECT 98.320 68.390 98.575 69.245 ;
        RECT 97.785 68.125 98.575 68.390 ;
        RECT 98.745 68.545 99.155 69.065 ;
        RECT 99.325 68.815 99.555 69.245 ;
        RECT 99.725 68.555 99.895 69.585 ;
        RECT 100.615 69.525 100.785 70.285 ;
        RECT 100.965 69.695 101.295 70.455 ;
        RECT 100.615 69.355 101.280 69.525 ;
        RECT 101.465 69.380 101.735 70.285 ;
        RECT 101.995 69.785 102.165 70.285 ;
        RECT 102.335 69.955 102.665 70.455 ;
        RECT 101.995 69.615 102.600 69.785 ;
        RECT 101.110 69.210 101.280 69.355 ;
        RECT 100.545 68.805 100.875 69.175 ;
        RECT 101.110 68.880 101.395 69.210 ;
        RECT 101.110 68.625 101.280 68.880 ;
        RECT 98.745 68.125 98.945 68.545 ;
        RECT 99.135 67.905 99.465 68.365 ;
        RECT 99.635 68.075 99.895 68.555 ;
        RECT 100.615 68.455 101.280 68.625 ;
        RECT 101.565 68.580 101.735 69.380 ;
        RECT 101.905 68.805 102.150 69.445 ;
        RECT 102.430 69.220 102.600 69.615 ;
        RECT 102.835 69.505 103.060 70.285 ;
        RECT 102.430 68.890 102.660 69.220 ;
        RECT 102.430 68.625 102.600 68.890 ;
        RECT 100.615 68.075 100.785 68.455 ;
        RECT 100.965 67.905 101.295 68.285 ;
        RECT 101.475 68.075 101.735 68.580 ;
        RECT 101.995 68.455 102.600 68.625 ;
        RECT 101.995 68.165 102.165 68.455 ;
        RECT 102.335 67.905 102.665 68.285 ;
        RECT 102.835 68.165 103.005 69.505 ;
        RECT 103.250 69.485 103.605 70.235 ;
        RECT 103.775 69.655 104.065 70.455 ;
        RECT 104.565 70.075 105.425 70.245 ;
        RECT 105.115 69.925 105.425 70.075 ;
        RECT 105.595 69.995 105.915 70.455 ;
        RECT 105.115 69.910 105.440 69.925 ;
        RECT 105.210 69.905 105.440 69.910 ;
        RECT 105.210 69.885 105.450 69.905 ;
        RECT 105.210 69.865 105.465 69.885 ;
        RECT 105.225 69.855 105.465 69.865 ;
        RECT 105.250 69.830 105.465 69.855 ;
        RECT 103.250 69.315 103.935 69.485 ;
        RECT 103.255 68.775 103.585 69.145 ;
        RECT 103.765 69.055 103.935 69.315 ;
        RECT 104.265 69.175 104.600 69.825 ;
        RECT 104.770 69.380 105.105 69.730 ;
        RECT 103.765 68.605 104.140 69.055 ;
        RECT 104.770 68.860 105.085 69.380 ;
        RECT 105.275 69.270 105.465 69.830 ;
        RECT 106.115 69.685 106.360 70.255 ;
        RECT 105.635 69.355 106.360 69.685 ;
        RECT 106.540 69.390 106.825 70.455 ;
        RECT 106.995 69.490 107.255 70.275 ;
        RECT 103.330 68.585 104.140 68.605 ;
        RECT 103.330 68.435 103.935 68.585 ;
        RECT 104.380 68.555 105.085 68.860 ;
        RECT 105.255 69.145 105.465 69.270 ;
        RECT 106.190 69.145 106.360 69.355 ;
        RECT 105.255 68.815 106.020 69.145 ;
        RECT 106.190 68.815 106.915 69.145 ;
        RECT 103.330 68.165 103.525 68.435 ;
        RECT 105.255 68.355 105.425 68.815 ;
        RECT 106.190 68.540 106.360 68.815 ;
        RECT 107.085 68.565 107.255 69.490 ;
        RECT 107.430 69.315 107.685 70.455 ;
        RECT 107.880 69.905 109.075 70.235 ;
        RECT 107.935 69.145 108.105 69.705 ;
        RECT 108.330 69.485 108.750 69.735 ;
        RECT 109.255 69.655 109.535 70.455 ;
        RECT 108.330 69.315 109.575 69.485 ;
        RECT 109.745 69.315 110.015 70.285 ;
        RECT 109.405 69.145 109.575 69.315 ;
        RECT 109.785 69.265 110.015 69.315 ;
        RECT 107.430 68.895 107.765 69.145 ;
        RECT 107.935 68.815 108.675 69.145 ;
        RECT 109.405 68.815 109.635 69.145 ;
        RECT 107.935 68.725 108.185 68.815 ;
        RECT 103.695 67.905 104.025 68.265 ;
        RECT 104.585 68.185 105.425 68.355 ;
        RECT 105.595 67.905 105.865 68.365 ;
        RECT 106.115 68.080 106.360 68.540 ;
        RECT 106.575 67.905 106.800 68.535 ;
        RECT 106.995 68.235 107.255 68.565 ;
        RECT 107.450 68.555 108.185 68.725 ;
        RECT 109.405 68.645 109.575 68.815 ;
        RECT 107.450 68.085 107.760 68.555 ;
        RECT 108.835 68.475 109.575 68.645 ;
        RECT 109.845 68.580 110.015 69.265 ;
        RECT 107.930 67.905 108.665 68.385 ;
        RECT 108.835 68.125 109.005 68.475 ;
        RECT 109.175 67.905 109.555 68.305 ;
        RECT 109.745 68.235 110.015 68.580 ;
        RECT 110.220 69.665 110.755 70.285 ;
        RECT 110.220 68.645 110.535 69.665 ;
        RECT 110.925 69.655 111.255 70.455 ;
        RECT 111.740 69.485 112.130 69.660 ;
        RECT 110.705 69.315 112.130 69.485 ;
        RECT 110.705 68.815 110.875 69.315 ;
        RECT 110.220 68.075 110.835 68.645 ;
        RECT 111.125 68.585 111.390 69.145 ;
        RECT 111.560 68.415 111.730 69.315 ;
        RECT 112.945 69.290 113.235 70.455 ;
        RECT 113.900 69.655 114.150 70.455 ;
        RECT 114.320 69.825 114.650 70.285 ;
        RECT 114.820 69.995 115.035 70.455 ;
        RECT 114.320 69.655 115.490 69.825 ;
        RECT 113.410 69.485 113.690 69.645 ;
        RECT 113.410 69.315 114.745 69.485 ;
        RECT 114.575 69.145 114.745 69.315 ;
        RECT 111.900 68.585 112.255 69.145 ;
        RECT 113.410 68.895 113.760 69.135 ;
        RECT 113.930 68.895 114.405 69.135 ;
        RECT 114.575 68.895 114.950 69.145 ;
        RECT 114.575 68.725 114.745 68.895 ;
        RECT 111.005 67.905 111.220 68.415 ;
        RECT 111.450 68.085 111.730 68.415 ;
        RECT 111.910 67.905 112.150 68.415 ;
        RECT 112.945 67.905 113.235 68.630 ;
        RECT 113.410 68.555 114.745 68.725 ;
        RECT 113.410 68.345 113.680 68.555 ;
        RECT 115.120 68.365 115.490 69.655 ;
        RECT 115.705 69.365 117.375 70.455 ;
        RECT 118.205 69.785 118.485 70.455 ;
        RECT 118.655 69.565 118.955 70.115 ;
        RECT 119.155 69.735 119.485 70.455 ;
        RECT 119.675 69.735 120.135 70.285 ;
        RECT 113.900 67.905 114.230 68.365 ;
        RECT 114.740 68.075 115.490 68.365 ;
        RECT 115.705 68.675 116.455 69.195 ;
        RECT 116.625 68.845 117.375 69.365 ;
        RECT 118.020 69.145 118.285 69.505 ;
        RECT 118.655 69.395 119.595 69.565 ;
        RECT 119.425 69.145 119.595 69.395 ;
        RECT 118.020 68.895 118.695 69.145 ;
        RECT 118.915 68.895 119.255 69.145 ;
        RECT 119.425 68.815 119.715 69.145 ;
        RECT 119.425 68.725 119.595 68.815 ;
        RECT 115.705 67.905 117.375 68.675 ;
        RECT 118.205 68.535 119.595 68.725 ;
        RECT 118.205 68.175 118.535 68.535 ;
        RECT 119.885 68.365 120.135 69.735 ;
        RECT 120.305 69.365 121.975 70.455 ;
        RECT 119.155 67.905 119.405 68.365 ;
        RECT 119.575 68.075 120.135 68.365 ;
        RECT 120.305 68.675 121.055 69.195 ;
        RECT 121.225 68.845 121.975 69.365 ;
        RECT 122.610 69.315 122.930 70.455 ;
        RECT 123.110 69.145 123.305 70.195 ;
        RECT 123.485 69.605 123.815 70.285 ;
        RECT 124.015 69.655 124.270 70.455 ;
        RECT 123.485 69.325 123.835 69.605 ;
        RECT 122.670 69.095 122.930 69.145 ;
        RECT 122.665 68.925 122.930 69.095 ;
        RECT 122.670 68.815 122.930 68.925 ;
        RECT 123.110 68.815 123.495 69.145 ;
        RECT 123.665 68.945 123.835 69.325 ;
        RECT 124.025 69.115 124.270 69.475 ;
        RECT 124.445 69.365 127.955 70.455 ;
        RECT 128.620 69.655 128.870 70.455 ;
        RECT 129.040 69.825 129.370 70.285 ;
        RECT 129.540 69.995 129.755 70.455 ;
        RECT 129.040 69.655 130.210 69.825 ;
        RECT 123.665 68.775 124.185 68.945 ;
        RECT 120.305 67.905 121.975 68.675 ;
        RECT 122.610 68.435 123.825 68.605 ;
        RECT 122.610 68.085 122.900 68.435 ;
        RECT 123.095 67.905 123.425 68.265 ;
        RECT 123.595 68.130 123.825 68.435 ;
        RECT 124.015 68.210 124.185 68.775 ;
        RECT 124.445 68.675 126.095 69.195 ;
        RECT 126.265 68.845 127.955 69.365 ;
        RECT 128.130 69.485 128.410 69.645 ;
        RECT 128.130 69.315 129.465 69.485 ;
        RECT 129.295 69.145 129.465 69.315 ;
        RECT 128.130 68.895 128.480 69.135 ;
        RECT 128.650 68.895 129.125 69.135 ;
        RECT 129.295 68.895 129.670 69.145 ;
        RECT 129.295 68.725 129.465 68.895 ;
        RECT 124.445 67.905 127.955 68.675 ;
        RECT 128.130 68.555 129.465 68.725 ;
        RECT 128.130 68.345 128.400 68.555 ;
        RECT 129.840 68.365 130.210 69.655 ;
        RECT 130.435 69.315 130.765 70.455 ;
        RECT 131.295 69.485 131.625 70.270 ;
        RECT 130.945 69.315 131.625 69.485 ;
        RECT 131.815 69.485 132.145 70.270 ;
        RECT 131.815 69.315 132.495 69.485 ;
        RECT 132.675 69.315 133.005 70.455 ;
        RECT 133.185 69.945 133.445 70.455 ;
        RECT 130.425 68.895 130.775 69.145 ;
        RECT 130.945 68.715 131.115 69.315 ;
        RECT 131.285 68.895 131.635 69.145 ;
        RECT 131.805 68.895 132.155 69.145 ;
        RECT 132.325 68.715 132.495 69.315 ;
        RECT 132.665 68.895 133.015 69.145 ;
        RECT 133.185 68.895 133.525 69.775 ;
        RECT 133.695 69.065 133.865 70.285 ;
        RECT 134.105 69.950 134.720 70.455 ;
        RECT 134.105 69.415 134.355 69.780 ;
        RECT 134.525 69.775 134.720 69.950 ;
        RECT 134.890 69.945 135.365 70.285 ;
        RECT 135.535 69.910 135.750 70.455 ;
        RECT 134.525 69.585 134.855 69.775 ;
        RECT 135.075 69.415 135.790 69.710 ;
        RECT 135.960 69.585 136.235 70.285 ;
        RECT 134.105 69.245 135.895 69.415 ;
        RECT 133.695 68.815 134.490 69.065 ;
        RECT 133.695 68.725 133.945 68.815 ;
        RECT 128.620 67.905 128.950 68.365 ;
        RECT 129.460 68.075 130.210 68.365 ;
        RECT 130.435 67.905 130.705 68.715 ;
        RECT 130.875 68.075 131.205 68.715 ;
        RECT 131.375 67.905 131.615 68.715 ;
        RECT 131.825 67.905 132.065 68.715 ;
        RECT 132.235 68.075 132.565 68.715 ;
        RECT 132.735 67.905 133.005 68.715 ;
        RECT 133.185 67.905 133.445 68.725 ;
        RECT 133.615 68.305 133.945 68.725 ;
        RECT 134.660 68.390 134.915 69.245 ;
        RECT 134.125 68.125 134.915 68.390 ;
        RECT 135.085 68.545 135.495 69.065 ;
        RECT 135.665 68.815 135.895 69.245 ;
        RECT 136.065 68.555 136.235 69.585 ;
        RECT 137.415 69.525 137.585 70.285 ;
        RECT 137.765 69.695 138.095 70.455 ;
        RECT 137.415 69.355 138.080 69.525 ;
        RECT 138.265 69.380 138.535 70.285 ;
        RECT 137.910 69.210 138.080 69.355 ;
        RECT 137.345 68.805 137.675 69.175 ;
        RECT 137.910 68.880 138.195 69.210 ;
        RECT 137.910 68.625 138.080 68.880 ;
        RECT 135.085 68.125 135.285 68.545 ;
        RECT 135.475 67.905 135.805 68.365 ;
        RECT 135.975 68.075 136.235 68.555 ;
        RECT 137.415 68.455 138.080 68.625 ;
        RECT 138.365 68.580 138.535 69.380 ;
        RECT 138.705 69.290 138.995 70.455 ;
        RECT 139.165 69.945 140.355 70.235 ;
        RECT 139.185 69.605 140.355 69.775 ;
        RECT 140.525 69.655 140.805 70.455 ;
        RECT 139.185 69.315 139.510 69.605 ;
        RECT 140.185 69.485 140.355 69.605 ;
        RECT 139.680 69.145 139.875 69.435 ;
        RECT 140.185 69.315 140.845 69.485 ;
        RECT 141.015 69.315 141.290 70.285 ;
        RECT 141.465 69.945 142.655 70.235 ;
        RECT 141.485 69.605 142.655 69.775 ;
        RECT 142.825 69.655 143.105 70.455 ;
        RECT 141.485 69.315 141.810 69.605 ;
        RECT 142.485 69.485 142.655 69.605 ;
        RECT 140.675 69.145 140.845 69.315 ;
        RECT 139.165 68.815 139.510 69.145 ;
        RECT 139.680 68.815 140.505 69.145 ;
        RECT 140.675 68.815 140.950 69.145 ;
        RECT 140.675 68.645 140.845 68.815 ;
        RECT 137.415 68.075 137.585 68.455 ;
        RECT 137.765 67.905 138.095 68.285 ;
        RECT 138.275 68.075 138.535 68.580 ;
        RECT 138.705 67.905 138.995 68.630 ;
        RECT 139.180 68.475 140.845 68.645 ;
        RECT 141.120 68.580 141.290 69.315 ;
        RECT 141.980 69.145 142.175 69.435 ;
        RECT 142.485 69.315 143.145 69.485 ;
        RECT 143.315 69.315 143.590 70.285 ;
        RECT 142.975 69.145 143.145 69.315 ;
        RECT 141.465 68.815 141.810 69.145 ;
        RECT 141.980 68.815 142.805 69.145 ;
        RECT 142.975 68.815 143.250 69.145 ;
        RECT 142.975 68.645 143.145 68.815 ;
        RECT 139.180 68.125 139.435 68.475 ;
        RECT 139.605 67.905 139.935 68.305 ;
        RECT 140.105 68.125 140.275 68.475 ;
        RECT 140.445 67.905 140.825 68.305 ;
        RECT 141.015 68.235 141.290 68.580 ;
        RECT 141.480 68.475 143.145 68.645 ;
        RECT 143.420 68.580 143.590 69.315 ;
        RECT 141.480 68.125 141.735 68.475 ;
        RECT 141.905 67.905 142.235 68.305 ;
        RECT 142.405 68.125 142.575 68.475 ;
        RECT 142.745 67.905 143.125 68.305 ;
        RECT 143.315 68.235 143.590 68.580 ;
        RECT 143.765 69.380 144.035 70.285 ;
        RECT 144.205 69.695 144.535 70.455 ;
        RECT 144.715 69.525 144.885 70.285 ;
        RECT 143.765 68.580 143.935 69.380 ;
        RECT 144.220 69.355 144.885 69.525 ;
        RECT 145.235 69.525 145.405 70.285 ;
        RECT 145.585 69.695 145.915 70.455 ;
        RECT 145.235 69.355 145.900 69.525 ;
        RECT 146.085 69.380 146.355 70.285 ;
        RECT 146.525 70.020 151.870 70.455 ;
        RECT 144.220 69.210 144.390 69.355 ;
        RECT 144.105 68.880 144.390 69.210 ;
        RECT 145.730 69.210 145.900 69.355 ;
        RECT 144.220 68.625 144.390 68.880 ;
        RECT 144.625 68.805 144.955 69.175 ;
        RECT 145.165 68.805 145.495 69.175 ;
        RECT 145.730 68.880 146.015 69.210 ;
        RECT 145.730 68.625 145.900 68.880 ;
        RECT 143.765 68.075 144.025 68.580 ;
        RECT 144.220 68.455 144.885 68.625 ;
        RECT 144.205 67.905 144.535 68.285 ;
        RECT 144.715 68.075 144.885 68.455 ;
        RECT 145.235 68.455 145.900 68.625 ;
        RECT 146.185 68.580 146.355 69.380 ;
        RECT 145.235 68.075 145.405 68.455 ;
        RECT 145.585 67.905 145.915 68.285 ;
        RECT 146.095 68.075 146.355 68.580 ;
        RECT 148.110 68.450 148.450 69.280 ;
        RECT 149.930 68.770 150.280 70.020 ;
        RECT 152.045 69.365 155.555 70.455 ;
        RECT 152.045 68.675 153.695 69.195 ;
        RECT 153.865 68.845 155.555 69.365 ;
        RECT 155.725 69.365 156.935 70.455 ;
        RECT 155.725 68.825 156.245 69.365 ;
        RECT 146.525 67.905 151.870 68.450 ;
        RECT 152.045 67.905 155.555 68.675 ;
        RECT 156.415 68.655 156.935 69.195 ;
        RECT 155.725 67.905 156.935 68.655 ;
        RECT 22.700 67.735 157.020 67.905 ;
        RECT 22.785 66.985 23.995 67.735 ;
        RECT 24.165 67.190 29.510 67.735 ;
        RECT 22.785 66.445 23.305 66.985 ;
        RECT 23.475 66.275 23.995 66.815 ;
        RECT 25.750 66.360 26.090 67.190 ;
        RECT 22.785 65.185 23.995 66.275 ;
        RECT 27.570 65.620 27.920 66.870 ;
        RECT 30.145 66.080 30.665 67.565 ;
        RECT 30.835 67.075 31.175 67.735 ;
        RECT 31.615 67.185 31.785 67.475 ;
        RECT 31.955 67.355 32.285 67.735 ;
        RECT 31.615 67.015 32.220 67.185 ;
        RECT 24.165 65.185 29.510 65.620 ;
        RECT 30.335 65.185 30.665 65.910 ;
        RECT 30.835 65.355 31.355 66.905 ;
        RECT 31.525 66.195 31.770 66.835 ;
        RECT 32.050 66.750 32.220 67.015 ;
        RECT 32.050 66.420 32.280 66.750 ;
        RECT 32.050 66.025 32.220 66.420 ;
        RECT 31.615 65.855 32.220 66.025 ;
        RECT 32.455 66.135 32.625 67.475 ;
        RECT 32.995 67.205 33.165 67.475 ;
        RECT 33.335 67.375 33.665 67.735 ;
        RECT 34.300 67.285 34.960 67.455 ;
        RECT 32.995 67.055 33.600 67.205 ;
        RECT 32.995 67.035 33.800 67.055 ;
        RECT 32.920 66.495 33.250 66.865 ;
        RECT 33.430 66.725 33.800 67.035 ;
        RECT 34.175 66.785 34.555 67.115 ;
        RECT 33.430 66.325 33.600 66.725 ;
        RECT 32.915 66.155 33.600 66.325 ;
        RECT 31.615 65.355 31.785 65.855 ;
        RECT 31.955 65.185 32.285 65.685 ;
        RECT 32.455 65.355 32.680 66.135 ;
        RECT 32.915 65.405 33.245 66.155 ;
        RECT 33.415 65.185 33.730 65.985 ;
        RECT 33.930 65.815 34.215 66.465 ;
        RECT 34.385 66.405 34.555 66.785 ;
        RECT 34.790 66.825 34.960 67.285 ;
        RECT 35.200 66.995 35.530 67.735 ;
        RECT 35.800 66.995 36.020 67.405 ;
        RECT 36.200 66.995 36.485 67.735 ;
        RECT 36.655 67.135 36.905 67.405 ;
        RECT 37.075 67.270 37.335 67.735 ;
        RECT 36.655 66.995 36.940 67.135 ;
        RECT 35.850 66.825 36.020 66.995 ;
        RECT 36.770 66.825 36.940 66.995 ;
        RECT 37.515 66.925 37.785 67.735 ;
        RECT 37.955 66.925 38.285 67.565 ;
        RECT 38.455 66.925 38.695 67.735 ;
        RECT 38.885 66.965 42.395 67.735 ;
        RECT 34.790 66.655 35.660 66.825 ;
        RECT 34.940 66.495 35.660 66.655 ;
        RECT 35.850 66.495 36.600 66.825 ;
        RECT 36.770 66.495 37.335 66.825 ;
        RECT 37.505 66.495 37.855 66.745 ;
        RECT 34.385 65.825 34.725 66.405 ;
        RECT 34.940 65.565 35.110 66.495 ;
        RECT 35.850 66.285 36.020 66.495 ;
        RECT 36.770 66.325 36.940 66.495 ;
        RECT 38.025 66.325 38.195 66.925 ;
        RECT 38.365 66.495 38.715 66.745 ;
        RECT 38.885 66.445 40.535 66.965 ;
        RECT 42.585 66.925 42.825 67.735 ;
        RECT 42.995 66.925 43.325 67.565 ;
        RECT 43.495 66.925 43.765 67.735 ;
        RECT 35.300 65.955 36.020 66.285 ;
        RECT 34.360 65.395 35.110 65.565 ;
        RECT 35.280 65.185 35.580 65.685 ;
        RECT 35.800 65.385 36.020 65.955 ;
        RECT 36.200 65.185 36.485 66.325 ;
        RECT 36.655 66.180 36.940 66.325 ;
        RECT 36.655 65.365 36.905 66.180 ;
        RECT 37.075 65.185 37.335 66.065 ;
        RECT 37.515 65.185 37.845 66.325 ;
        RECT 38.025 66.155 38.705 66.325 ;
        RECT 40.705 66.275 42.395 66.795 ;
        RECT 42.565 66.495 42.915 66.745 ;
        RECT 43.085 66.325 43.255 66.925 ;
        RECT 44.005 66.915 44.215 67.735 ;
        RECT 44.385 66.935 44.715 67.565 ;
        RECT 43.425 66.495 43.775 66.745 ;
        RECT 44.385 66.335 44.635 66.935 ;
        RECT 44.885 66.915 45.115 67.735 ;
        RECT 45.325 66.965 46.995 67.735 ;
        RECT 44.805 66.495 45.135 66.745 ;
        RECT 45.325 66.445 46.075 66.965 ;
        RECT 47.175 66.925 47.445 67.735 ;
        RECT 47.615 66.925 47.945 67.565 ;
        RECT 48.115 66.925 48.355 67.735 ;
        RECT 48.545 67.010 48.835 67.735 ;
        RECT 49.005 67.270 49.265 67.735 ;
        RECT 49.435 67.135 49.685 67.405 ;
        RECT 49.400 66.995 49.685 67.135 ;
        RECT 49.855 66.995 50.140 67.735 ;
        RECT 50.320 66.995 50.540 67.405 ;
        RECT 50.810 66.995 51.140 67.735 ;
        RECT 51.380 67.285 52.040 67.455 ;
        RECT 52.675 67.375 53.005 67.735 ;
        RECT 38.375 65.370 38.705 66.155 ;
        RECT 38.885 65.185 42.395 66.275 ;
        RECT 42.575 66.155 43.255 66.325 ;
        RECT 42.575 65.370 42.905 66.155 ;
        RECT 43.435 65.185 43.765 66.325 ;
        RECT 44.005 65.185 44.215 66.325 ;
        RECT 44.385 65.355 44.715 66.335 ;
        RECT 44.885 65.185 45.115 66.325 ;
        RECT 46.245 66.275 46.995 66.795 ;
        RECT 47.165 66.495 47.515 66.745 ;
        RECT 47.685 66.325 47.855 66.925 ;
        RECT 49.400 66.825 49.570 66.995 ;
        RECT 50.320 66.825 50.490 66.995 ;
        RECT 51.380 66.825 51.550 67.285 ;
        RECT 53.175 67.205 53.345 67.475 ;
        RECT 48.025 66.495 48.375 66.745 ;
        RECT 49.005 66.495 49.570 66.825 ;
        RECT 49.740 66.495 50.490 66.825 ;
        RECT 50.680 66.655 51.550 66.825 ;
        RECT 51.785 66.785 52.165 67.115 ;
        RECT 52.740 67.055 53.345 67.205 ;
        RECT 52.540 67.035 53.345 67.055 ;
        RECT 50.680 66.495 51.400 66.655 ;
        RECT 45.325 65.185 46.995 66.275 ;
        RECT 47.175 65.185 47.505 66.325 ;
        RECT 47.685 66.155 48.365 66.325 ;
        RECT 48.035 65.370 48.365 66.155 ;
        RECT 48.545 65.185 48.835 66.350 ;
        RECT 49.400 66.325 49.570 66.495 ;
        RECT 49.400 66.180 49.685 66.325 ;
        RECT 49.005 65.185 49.265 66.065 ;
        RECT 49.435 65.365 49.685 66.180 ;
        RECT 49.855 65.185 50.140 66.325 ;
        RECT 50.320 66.285 50.490 66.495 ;
        RECT 50.320 65.955 51.040 66.285 ;
        RECT 50.320 65.385 50.540 65.955 ;
        RECT 50.760 65.185 51.060 65.685 ;
        RECT 51.230 65.565 51.400 66.495 ;
        RECT 51.785 66.405 51.955 66.785 ;
        RECT 52.540 66.725 52.910 67.035 ;
        RECT 51.615 65.825 51.955 66.405 ;
        RECT 52.125 65.815 52.410 66.465 ;
        RECT 52.740 66.325 52.910 66.725 ;
        RECT 53.090 66.495 53.420 66.865 ;
        RECT 52.740 66.155 53.425 66.325 ;
        RECT 51.230 65.395 51.980 65.565 ;
        RECT 52.610 65.185 52.925 65.985 ;
        RECT 53.095 65.405 53.425 66.155 ;
        RECT 53.715 66.135 53.885 67.475 ;
        RECT 54.055 67.355 54.385 67.735 ;
        RECT 54.555 67.185 54.725 67.475 ;
        RECT 54.120 67.015 54.725 67.185 ;
        RECT 55.165 67.075 55.505 67.735 ;
        RECT 54.120 66.750 54.290 67.015 ;
        RECT 54.060 66.420 54.290 66.750 ;
        RECT 53.660 65.355 53.885 66.135 ;
        RECT 54.120 66.025 54.290 66.420 ;
        RECT 54.570 66.195 54.815 66.835 ;
        RECT 54.120 65.855 54.725 66.025 ;
        RECT 54.055 65.185 54.385 65.685 ;
        RECT 54.555 65.355 54.725 65.855 ;
        RECT 54.985 65.355 55.505 66.905 ;
        RECT 55.675 66.080 56.195 67.565 ;
        RECT 56.375 66.925 56.645 67.735 ;
        RECT 56.815 66.925 57.145 67.565 ;
        RECT 57.315 66.925 57.555 67.735 ;
        RECT 57.755 66.925 58.025 67.735 ;
        RECT 58.195 66.925 58.525 67.565 ;
        RECT 58.695 66.925 58.935 67.735 ;
        RECT 59.135 66.925 59.405 67.735 ;
        RECT 59.575 66.925 59.905 67.565 ;
        RECT 60.075 66.925 60.315 67.735 ;
        RECT 60.595 67.185 60.765 67.475 ;
        RECT 60.935 67.355 61.265 67.735 ;
        RECT 60.595 67.015 61.200 67.185 ;
        RECT 56.365 66.495 56.715 66.745 ;
        RECT 56.885 66.325 57.055 66.925 ;
        RECT 57.225 66.495 57.575 66.745 ;
        RECT 57.745 66.495 58.095 66.745 ;
        RECT 58.265 66.325 58.435 66.925 ;
        RECT 58.605 66.495 58.955 66.745 ;
        RECT 59.125 66.495 59.475 66.745 ;
        RECT 59.645 66.325 59.815 66.925 ;
        RECT 59.985 66.495 60.335 66.745 ;
        RECT 55.675 65.185 56.005 65.910 ;
        RECT 56.375 65.185 56.705 66.325 ;
        RECT 56.885 66.155 57.565 66.325 ;
        RECT 57.235 65.370 57.565 66.155 ;
        RECT 57.755 65.185 58.085 66.325 ;
        RECT 58.265 66.155 58.945 66.325 ;
        RECT 58.615 65.370 58.945 66.155 ;
        RECT 59.135 65.185 59.465 66.325 ;
        RECT 59.645 66.155 60.325 66.325 ;
        RECT 60.505 66.195 60.750 66.835 ;
        RECT 61.030 66.750 61.200 67.015 ;
        RECT 61.030 66.420 61.260 66.750 ;
        RECT 59.995 65.370 60.325 66.155 ;
        RECT 61.030 66.025 61.200 66.420 ;
        RECT 60.595 65.855 61.200 66.025 ;
        RECT 61.435 66.135 61.605 67.475 ;
        RECT 61.975 67.205 62.145 67.475 ;
        RECT 62.315 67.375 62.645 67.735 ;
        RECT 63.280 67.285 63.940 67.455 ;
        RECT 61.975 67.055 62.580 67.205 ;
        RECT 61.975 67.035 62.780 67.055 ;
        RECT 61.900 66.495 62.230 66.865 ;
        RECT 62.410 66.725 62.780 67.035 ;
        RECT 63.155 66.785 63.535 67.115 ;
        RECT 62.410 66.325 62.580 66.725 ;
        RECT 61.895 66.155 62.580 66.325 ;
        RECT 60.595 65.355 60.765 65.855 ;
        RECT 60.935 65.185 61.265 65.685 ;
        RECT 61.435 65.355 61.660 66.135 ;
        RECT 61.895 65.405 62.225 66.155 ;
        RECT 62.395 65.185 62.710 65.985 ;
        RECT 62.910 65.815 63.195 66.465 ;
        RECT 63.365 66.405 63.535 66.785 ;
        RECT 63.770 66.825 63.940 67.285 ;
        RECT 64.180 66.995 64.510 67.735 ;
        RECT 64.780 66.995 65.000 67.405 ;
        RECT 65.180 66.995 65.465 67.735 ;
        RECT 65.635 67.135 65.885 67.405 ;
        RECT 66.055 67.270 66.315 67.735 ;
        RECT 65.635 66.995 65.920 67.135 ;
        RECT 64.830 66.825 65.000 66.995 ;
        RECT 65.750 66.825 65.920 66.995 ;
        RECT 66.485 66.965 68.155 67.735 ;
        RECT 63.770 66.655 64.640 66.825 ;
        RECT 63.920 66.495 64.640 66.655 ;
        RECT 64.830 66.495 65.580 66.825 ;
        RECT 65.750 66.495 66.315 66.825 ;
        RECT 63.365 65.825 63.705 66.405 ;
        RECT 63.920 65.565 64.090 66.495 ;
        RECT 64.830 66.285 65.000 66.495 ;
        RECT 65.750 66.325 65.920 66.495 ;
        RECT 66.485 66.445 67.235 66.965 ;
        RECT 68.345 66.925 68.585 67.735 ;
        RECT 68.755 66.925 69.085 67.565 ;
        RECT 69.255 66.925 69.525 67.735 ;
        RECT 69.715 66.925 69.985 67.735 ;
        RECT 70.155 66.925 70.485 67.565 ;
        RECT 70.655 66.925 70.895 67.735 ;
        RECT 71.105 66.925 71.345 67.735 ;
        RECT 71.515 66.925 71.845 67.565 ;
        RECT 72.015 66.925 72.285 67.735 ;
        RECT 72.465 66.965 74.135 67.735 ;
        RECT 74.305 67.010 74.595 67.735 ;
        RECT 64.280 65.955 65.000 66.285 ;
        RECT 63.340 65.395 64.090 65.565 ;
        RECT 64.260 65.185 64.560 65.685 ;
        RECT 64.780 65.385 65.000 65.955 ;
        RECT 65.180 65.185 65.465 66.325 ;
        RECT 65.635 66.180 65.920 66.325 ;
        RECT 67.405 66.275 68.155 66.795 ;
        RECT 68.325 66.495 68.675 66.745 ;
        RECT 68.845 66.325 69.015 66.925 ;
        RECT 69.185 66.495 69.535 66.745 ;
        RECT 69.705 66.495 70.055 66.745 ;
        RECT 70.225 66.325 70.395 66.925 ;
        RECT 70.565 66.495 70.915 66.745 ;
        RECT 71.085 66.495 71.435 66.745 ;
        RECT 71.605 66.325 71.775 66.925 ;
        RECT 71.945 66.495 72.295 66.745 ;
        RECT 72.465 66.445 73.215 66.965 ;
        RECT 74.775 66.925 75.045 67.735 ;
        RECT 75.215 66.925 75.545 67.565 ;
        RECT 75.715 66.925 75.955 67.735 ;
        RECT 76.615 66.925 76.885 67.735 ;
        RECT 77.055 66.925 77.385 67.565 ;
        RECT 77.555 66.925 77.795 67.735 ;
        RECT 77.995 66.925 78.265 67.735 ;
        RECT 78.435 66.925 78.765 67.565 ;
        RECT 78.935 66.925 79.175 67.735 ;
        RECT 79.365 66.965 81.035 67.735 ;
        RECT 81.845 67.075 82.185 67.735 ;
        RECT 65.635 65.365 65.885 66.180 ;
        RECT 66.055 65.185 66.315 66.065 ;
        RECT 66.485 65.185 68.155 66.275 ;
        RECT 68.335 66.155 69.015 66.325 ;
        RECT 68.335 65.370 68.665 66.155 ;
        RECT 69.195 65.185 69.525 66.325 ;
        RECT 69.715 65.185 70.045 66.325 ;
        RECT 70.225 66.155 70.905 66.325 ;
        RECT 70.575 65.370 70.905 66.155 ;
        RECT 71.095 66.155 71.775 66.325 ;
        RECT 71.095 65.370 71.425 66.155 ;
        RECT 71.955 65.185 72.285 66.325 ;
        RECT 73.385 66.275 74.135 66.795 ;
        RECT 74.765 66.495 75.115 66.745 ;
        RECT 72.465 65.185 74.135 66.275 ;
        RECT 74.305 65.185 74.595 66.350 ;
        RECT 75.285 66.325 75.455 66.925 ;
        RECT 75.625 66.495 75.975 66.745 ;
        RECT 76.605 66.495 76.955 66.745 ;
        RECT 77.125 66.325 77.295 66.925 ;
        RECT 77.465 66.495 77.815 66.745 ;
        RECT 77.985 66.495 78.335 66.745 ;
        RECT 78.505 66.325 78.675 66.925 ;
        RECT 78.845 66.495 79.195 66.745 ;
        RECT 79.365 66.445 80.115 66.965 ;
        RECT 74.775 65.185 75.105 66.325 ;
        RECT 75.285 66.155 75.965 66.325 ;
        RECT 75.635 65.370 75.965 66.155 ;
        RECT 76.615 65.185 76.945 66.325 ;
        RECT 77.125 66.155 77.805 66.325 ;
        RECT 77.475 65.370 77.805 66.155 ;
        RECT 77.995 65.185 78.325 66.325 ;
        RECT 78.505 66.155 79.185 66.325 ;
        RECT 80.285 66.275 81.035 66.795 ;
        RECT 78.855 65.370 79.185 66.155 ;
        RECT 79.365 65.185 81.035 66.275 ;
        RECT 81.665 65.355 82.185 66.905 ;
        RECT 82.355 66.080 82.875 67.565 ;
        RECT 83.045 67.190 88.390 67.735 ;
        RECT 84.630 66.360 84.970 67.190 ;
        RECT 89.495 66.925 89.765 67.735 ;
        RECT 89.935 66.925 90.265 67.565 ;
        RECT 90.435 66.925 90.675 67.735 ;
        RECT 90.865 67.190 96.210 67.735 ;
        RECT 82.355 65.185 82.685 65.910 ;
        RECT 86.450 65.620 86.800 66.870 ;
        RECT 89.485 66.495 89.835 66.745 ;
        RECT 90.005 66.325 90.175 66.925 ;
        RECT 90.345 66.495 90.695 66.745 ;
        RECT 92.450 66.360 92.790 67.190 ;
        RECT 96.565 67.075 96.905 67.735 ;
        RECT 83.045 65.185 88.390 65.620 ;
        RECT 89.495 65.185 89.825 66.325 ;
        RECT 90.005 66.155 90.685 66.325 ;
        RECT 90.355 65.370 90.685 66.155 ;
        RECT 94.270 65.620 94.620 66.870 ;
        RECT 90.865 65.185 96.210 65.620 ;
        RECT 96.385 65.355 96.905 66.905 ;
        RECT 97.075 66.080 97.595 67.565 ;
        RECT 97.780 67.165 98.035 67.515 ;
        RECT 98.205 67.335 98.535 67.735 ;
        RECT 98.705 67.165 98.875 67.515 ;
        RECT 99.045 67.335 99.425 67.735 ;
        RECT 97.780 66.995 99.445 67.165 ;
        RECT 99.615 67.060 99.890 67.405 ;
        RECT 99.275 66.825 99.445 66.995 ;
        RECT 97.765 66.495 98.110 66.825 ;
        RECT 98.280 66.495 99.105 66.825 ;
        RECT 99.275 66.495 99.550 66.825 ;
        RECT 97.785 66.035 98.110 66.325 ;
        RECT 98.280 66.205 98.475 66.495 ;
        RECT 99.275 66.325 99.445 66.495 ;
        RECT 99.720 66.325 99.890 67.060 ;
        RECT 100.065 67.010 100.355 67.735 ;
        RECT 100.615 67.185 100.785 67.565 ;
        RECT 100.965 67.355 101.295 67.735 ;
        RECT 100.615 67.015 101.280 67.185 ;
        RECT 101.475 67.060 101.735 67.565 ;
        RECT 100.545 66.465 100.875 66.835 ;
        RECT 101.110 66.760 101.280 67.015 ;
        RECT 101.110 66.430 101.395 66.760 ;
        RECT 98.785 66.155 99.445 66.325 ;
        RECT 98.785 66.035 98.955 66.155 ;
        RECT 97.075 65.185 97.405 65.910 ;
        RECT 97.785 65.865 98.955 66.035 ;
        RECT 97.765 65.405 98.955 65.695 ;
        RECT 99.125 65.185 99.405 65.985 ;
        RECT 99.615 65.355 99.890 66.325 ;
        RECT 100.065 65.185 100.355 66.350 ;
        RECT 101.110 66.285 101.280 66.430 ;
        RECT 100.615 66.115 101.280 66.285 ;
        RECT 101.565 66.260 101.735 67.060 ;
        RECT 101.995 67.185 102.165 67.565 ;
        RECT 102.345 67.355 102.675 67.735 ;
        RECT 101.995 67.015 102.660 67.185 ;
        RECT 102.855 67.060 103.115 67.565 ;
        RECT 101.925 66.465 102.255 66.835 ;
        RECT 102.490 66.760 102.660 67.015 ;
        RECT 102.490 66.430 102.775 66.760 ;
        RECT 102.490 66.285 102.660 66.430 ;
        RECT 100.615 65.355 100.785 66.115 ;
        RECT 100.965 65.185 101.295 65.945 ;
        RECT 101.465 65.355 101.735 66.260 ;
        RECT 101.995 66.115 102.660 66.285 ;
        RECT 102.945 66.260 103.115 67.060 ;
        RECT 103.285 66.965 106.795 67.735 ;
        RECT 106.965 66.985 108.175 67.735 ;
        RECT 103.285 66.445 104.935 66.965 ;
        RECT 105.105 66.275 106.795 66.795 ;
        RECT 106.965 66.445 107.485 66.985 ;
        RECT 108.365 66.925 108.605 67.735 ;
        RECT 108.775 66.925 109.105 67.565 ;
        RECT 109.275 66.925 109.545 67.735 ;
        RECT 109.735 66.925 110.005 67.735 ;
        RECT 110.175 66.925 110.505 67.565 ;
        RECT 110.675 66.925 110.915 67.735 ;
        RECT 111.105 66.965 112.775 67.735 ;
        RECT 107.655 66.275 108.175 66.815 ;
        RECT 108.345 66.495 108.695 66.745 ;
        RECT 108.865 66.325 109.035 66.925 ;
        RECT 109.205 66.495 109.555 66.745 ;
        RECT 109.725 66.495 110.075 66.745 ;
        RECT 110.245 66.325 110.415 66.925 ;
        RECT 110.585 66.495 110.935 66.745 ;
        RECT 111.105 66.445 111.855 66.965 ;
        RECT 112.955 66.925 113.225 67.735 ;
        RECT 113.395 66.925 113.725 67.565 ;
        RECT 113.895 66.925 114.135 67.735 ;
        RECT 114.335 66.925 114.605 67.735 ;
        RECT 114.775 66.925 115.105 67.565 ;
        RECT 115.275 66.925 115.515 67.735 ;
        RECT 115.705 66.965 118.295 67.735 ;
        RECT 101.995 65.355 102.165 66.115 ;
        RECT 102.345 65.185 102.675 65.945 ;
        RECT 102.845 65.355 103.115 66.260 ;
        RECT 103.285 65.185 106.795 66.275 ;
        RECT 106.965 65.185 108.175 66.275 ;
        RECT 108.355 66.155 109.035 66.325 ;
        RECT 108.355 65.370 108.685 66.155 ;
        RECT 109.215 65.185 109.545 66.325 ;
        RECT 109.735 65.185 110.065 66.325 ;
        RECT 110.245 66.155 110.925 66.325 ;
        RECT 112.025 66.275 112.775 66.795 ;
        RECT 112.945 66.495 113.295 66.745 ;
        RECT 113.465 66.325 113.635 66.925 ;
        RECT 113.805 66.495 114.155 66.745 ;
        RECT 114.325 66.495 114.675 66.745 ;
        RECT 114.845 66.325 115.015 66.925 ;
        RECT 115.185 66.495 115.535 66.745 ;
        RECT 115.705 66.445 116.915 66.965 ;
        RECT 118.935 66.925 119.205 67.735 ;
        RECT 119.375 66.925 119.705 67.565 ;
        RECT 119.875 66.925 120.115 67.735 ;
        RECT 120.315 66.925 120.585 67.735 ;
        RECT 120.755 66.925 121.085 67.565 ;
        RECT 121.255 66.925 121.495 67.735 ;
        RECT 121.685 66.985 122.895 67.735 ;
        RECT 110.595 65.370 110.925 66.155 ;
        RECT 111.105 65.185 112.775 66.275 ;
        RECT 112.955 65.185 113.285 66.325 ;
        RECT 113.465 66.155 114.145 66.325 ;
        RECT 113.815 65.370 114.145 66.155 ;
        RECT 114.335 65.185 114.665 66.325 ;
        RECT 114.845 66.155 115.525 66.325 ;
        RECT 117.085 66.275 118.295 66.795 ;
        RECT 118.925 66.495 119.275 66.745 ;
        RECT 119.445 66.325 119.615 66.925 ;
        RECT 119.785 66.495 120.135 66.745 ;
        RECT 120.305 66.495 120.655 66.745 ;
        RECT 120.825 66.325 120.995 66.925 ;
        RECT 121.165 66.495 121.515 66.745 ;
        RECT 121.685 66.445 122.205 66.985 ;
        RECT 123.075 66.925 123.345 67.735 ;
        RECT 123.515 66.925 123.845 67.565 ;
        RECT 124.015 66.925 124.255 67.735 ;
        RECT 124.445 66.985 125.655 67.735 ;
        RECT 125.825 67.010 126.115 67.735 ;
        RECT 115.195 65.370 115.525 66.155 ;
        RECT 115.705 65.185 118.295 66.275 ;
        RECT 118.935 65.185 119.265 66.325 ;
        RECT 119.445 66.155 120.125 66.325 ;
        RECT 119.795 65.370 120.125 66.155 ;
        RECT 120.315 65.185 120.645 66.325 ;
        RECT 120.825 66.155 121.505 66.325 ;
        RECT 122.375 66.275 122.895 66.815 ;
        RECT 123.065 66.495 123.415 66.745 ;
        RECT 123.585 66.325 123.755 66.925 ;
        RECT 123.925 66.495 124.275 66.745 ;
        RECT 124.445 66.445 124.965 66.985 ;
        RECT 126.285 66.965 128.875 67.735 ;
        RECT 121.175 65.370 121.505 66.155 ;
        RECT 121.685 65.185 122.895 66.275 ;
        RECT 123.075 65.185 123.405 66.325 ;
        RECT 123.585 66.155 124.265 66.325 ;
        RECT 125.135 66.275 125.655 66.815 ;
        RECT 126.285 66.445 127.495 66.965 ;
        RECT 129.515 66.925 129.785 67.735 ;
        RECT 129.955 66.925 130.285 67.565 ;
        RECT 130.455 66.925 130.695 67.735 ;
        RECT 130.895 66.925 131.165 67.735 ;
        RECT 131.335 66.925 131.665 67.565 ;
        RECT 131.835 66.925 132.075 67.735 ;
        RECT 123.935 65.370 124.265 66.155 ;
        RECT 124.445 65.185 125.655 66.275 ;
        RECT 125.825 65.185 126.115 66.350 ;
        RECT 127.665 66.275 128.875 66.795 ;
        RECT 129.505 66.495 129.855 66.745 ;
        RECT 130.025 66.325 130.195 66.925 ;
        RECT 130.365 66.495 130.715 66.745 ;
        RECT 130.885 66.495 131.235 66.745 ;
        RECT 131.405 66.325 131.575 66.925 ;
        RECT 133.185 66.915 133.445 67.735 ;
        RECT 133.615 66.915 133.945 67.335 ;
        RECT 134.125 67.250 134.915 67.515 ;
        RECT 133.695 66.825 133.945 66.915 ;
        RECT 131.745 66.495 132.095 66.745 ;
        RECT 126.285 65.185 128.875 66.275 ;
        RECT 129.515 65.185 129.845 66.325 ;
        RECT 130.025 66.155 130.705 66.325 ;
        RECT 130.375 65.370 130.705 66.155 ;
        RECT 130.895 65.185 131.225 66.325 ;
        RECT 131.405 66.155 132.085 66.325 ;
        RECT 131.755 65.370 132.085 66.155 ;
        RECT 133.185 65.865 133.525 66.745 ;
        RECT 133.695 66.575 134.490 66.825 ;
        RECT 133.185 65.185 133.445 65.695 ;
        RECT 133.695 65.355 133.865 66.575 ;
        RECT 134.660 66.395 134.915 67.250 ;
        RECT 135.085 67.095 135.285 67.515 ;
        RECT 135.475 67.275 135.805 67.735 ;
        RECT 135.085 66.575 135.495 67.095 ;
        RECT 135.975 67.085 136.235 67.565 ;
        RECT 135.665 66.395 135.895 66.825 ;
        RECT 134.105 66.225 135.895 66.395 ;
        RECT 134.105 65.860 134.355 66.225 ;
        RECT 134.525 65.865 134.855 66.055 ;
        RECT 135.075 65.930 135.790 66.225 ;
        RECT 136.065 66.055 136.235 67.085 ;
        RECT 136.405 66.985 137.615 67.735 ;
        RECT 137.875 67.185 138.045 67.565 ;
        RECT 138.225 67.355 138.555 67.735 ;
        RECT 137.875 67.015 138.540 67.185 ;
        RECT 138.735 67.060 138.995 67.565 ;
        RECT 139.165 67.190 144.510 67.735 ;
        RECT 144.685 67.190 150.030 67.735 ;
        RECT 136.405 66.445 136.925 66.985 ;
        RECT 137.095 66.275 137.615 66.815 ;
        RECT 137.805 66.465 138.135 66.835 ;
        RECT 138.370 66.760 138.540 67.015 ;
        RECT 138.370 66.430 138.655 66.760 ;
        RECT 138.370 66.285 138.540 66.430 ;
        RECT 134.525 65.690 134.720 65.865 ;
        RECT 134.105 65.185 134.720 65.690 ;
        RECT 134.890 65.355 135.365 65.695 ;
        RECT 135.535 65.185 135.750 65.730 ;
        RECT 135.960 65.355 136.235 66.055 ;
        RECT 136.405 65.185 137.615 66.275 ;
        RECT 137.875 66.115 138.540 66.285 ;
        RECT 138.825 66.260 138.995 67.060 ;
        RECT 140.750 66.360 141.090 67.190 ;
        RECT 137.875 65.355 138.045 66.115 ;
        RECT 138.225 65.185 138.555 65.945 ;
        RECT 138.725 65.355 138.995 66.260 ;
        RECT 142.570 65.620 142.920 66.870 ;
        RECT 146.270 66.360 146.610 67.190 ;
        RECT 150.205 66.985 151.415 67.735 ;
        RECT 151.585 67.010 151.875 67.735 ;
        RECT 148.090 65.620 148.440 66.870 ;
        RECT 150.205 66.445 150.725 66.985 ;
        RECT 152.045 66.965 155.555 67.735 ;
        RECT 155.725 66.985 156.935 67.735 ;
        RECT 150.895 66.275 151.415 66.815 ;
        RECT 152.045 66.445 153.695 66.965 ;
        RECT 139.165 65.185 144.510 65.620 ;
        RECT 144.685 65.185 150.030 65.620 ;
        RECT 150.205 65.185 151.415 66.275 ;
        RECT 151.585 65.185 151.875 66.350 ;
        RECT 153.865 66.275 155.555 66.795 ;
        RECT 152.045 65.185 155.555 66.275 ;
        RECT 155.725 66.275 156.245 66.815 ;
        RECT 156.415 66.445 156.935 66.985 ;
        RECT 155.725 65.185 156.935 66.275 ;
        RECT 22.700 65.015 157.020 65.185 ;
        RECT 22.785 63.925 23.995 65.015 ;
        RECT 24.715 64.345 24.885 64.845 ;
        RECT 25.055 64.515 25.385 65.015 ;
        RECT 24.715 64.175 25.320 64.345 ;
        RECT 22.785 63.215 23.305 63.755 ;
        RECT 23.475 63.385 23.995 63.925 ;
        RECT 24.625 63.365 24.870 64.005 ;
        RECT 25.150 63.780 25.320 64.175 ;
        RECT 25.555 64.065 25.780 64.845 ;
        RECT 25.150 63.450 25.380 63.780 ;
        RECT 22.785 62.465 23.995 63.215 ;
        RECT 25.150 63.185 25.320 63.450 ;
        RECT 24.715 63.015 25.320 63.185 ;
        RECT 24.715 62.725 24.885 63.015 ;
        RECT 25.055 62.465 25.385 62.845 ;
        RECT 25.555 62.725 25.725 64.065 ;
        RECT 26.015 64.045 26.345 64.795 ;
        RECT 26.515 64.215 26.830 65.015 ;
        RECT 27.460 64.635 28.210 64.805 ;
        RECT 26.015 63.875 26.700 64.045 ;
        RECT 26.020 63.335 26.350 63.705 ;
        RECT 26.530 63.475 26.700 63.875 ;
        RECT 27.030 63.735 27.315 64.385 ;
        RECT 27.485 63.795 27.825 64.375 ;
        RECT 26.530 63.165 26.900 63.475 ;
        RECT 27.485 63.415 27.655 63.795 ;
        RECT 28.040 63.705 28.210 64.635 ;
        RECT 28.380 64.515 28.680 65.015 ;
        RECT 28.900 64.245 29.120 64.815 ;
        RECT 28.400 63.915 29.120 64.245 ;
        RECT 28.950 63.705 29.120 63.915 ;
        RECT 29.300 63.875 29.585 65.015 ;
        RECT 29.755 64.020 30.005 64.835 ;
        RECT 30.175 64.135 30.435 65.015 ;
        RECT 29.755 63.875 30.040 64.020 ;
        RECT 29.870 63.705 30.040 63.875 ;
        RECT 28.040 63.545 28.760 63.705 ;
        RECT 26.095 63.145 26.900 63.165 ;
        RECT 26.095 62.995 26.700 63.145 ;
        RECT 27.275 63.085 27.655 63.415 ;
        RECT 27.890 63.375 28.760 63.545 ;
        RECT 28.950 63.375 29.700 63.705 ;
        RECT 29.870 63.375 30.435 63.705 ;
        RECT 26.095 62.725 26.265 62.995 ;
        RECT 27.890 62.915 28.060 63.375 ;
        RECT 28.950 63.205 29.120 63.375 ;
        RECT 29.870 63.205 30.040 63.375 ;
        RECT 30.605 63.295 31.125 64.845 ;
        RECT 31.295 64.290 31.625 65.015 ;
        RECT 26.435 62.465 26.765 62.825 ;
        RECT 27.400 62.745 28.060 62.915 ;
        RECT 28.300 62.465 28.630 63.205 ;
        RECT 28.900 62.795 29.120 63.205 ;
        RECT 29.300 62.465 29.585 63.205 ;
        RECT 29.755 63.065 30.040 63.205 ;
        RECT 29.755 62.795 30.005 63.065 ;
        RECT 30.175 62.465 30.435 62.930 ;
        RECT 30.785 62.465 31.125 63.125 ;
        RECT 31.295 62.635 31.815 64.120 ;
        RECT 31.985 63.925 33.655 65.015 ;
        RECT 31.985 63.235 32.735 63.755 ;
        RECT 32.905 63.405 33.655 63.925 ;
        RECT 33.835 64.045 34.165 64.830 ;
        RECT 33.835 63.875 34.515 64.045 ;
        RECT 34.695 63.875 35.025 65.015 ;
        RECT 33.825 63.455 34.175 63.705 ;
        RECT 34.345 63.275 34.515 63.875 ;
        RECT 35.665 63.850 35.955 65.015 ;
        RECT 36.135 63.875 36.465 65.015 ;
        RECT 36.995 64.045 37.325 64.830 ;
        RECT 36.645 63.875 37.325 64.045 ;
        RECT 37.515 63.875 37.845 65.015 ;
        RECT 38.375 64.045 38.705 64.830 ;
        RECT 38.025 63.875 38.705 64.045 ;
        RECT 38.885 63.925 40.095 65.015 ;
        RECT 40.455 64.290 40.785 65.015 ;
        RECT 34.685 63.455 35.035 63.705 ;
        RECT 36.125 63.455 36.475 63.705 ;
        RECT 36.645 63.275 36.815 63.875 ;
        RECT 36.985 63.455 37.335 63.705 ;
        RECT 37.505 63.455 37.855 63.705 ;
        RECT 38.025 63.275 38.195 63.875 ;
        RECT 38.365 63.455 38.715 63.705 ;
        RECT 31.985 62.465 33.655 63.235 ;
        RECT 33.845 62.465 34.085 63.275 ;
        RECT 34.255 62.635 34.585 63.275 ;
        RECT 34.755 62.465 35.025 63.275 ;
        RECT 35.665 62.465 35.955 63.190 ;
        RECT 36.135 62.465 36.405 63.275 ;
        RECT 36.575 62.635 36.905 63.275 ;
        RECT 37.075 62.465 37.315 63.275 ;
        RECT 37.515 62.465 37.785 63.275 ;
        RECT 37.955 62.635 38.285 63.275 ;
        RECT 38.455 62.465 38.695 63.275 ;
        RECT 38.885 63.215 39.405 63.755 ;
        RECT 39.575 63.385 40.095 63.925 ;
        RECT 38.885 62.465 40.095 63.215 ;
        RECT 40.265 62.635 40.785 64.120 ;
        RECT 40.955 63.295 41.475 64.845 ;
        RECT 41.655 64.045 41.985 64.830 ;
        RECT 41.655 63.875 42.335 64.045 ;
        RECT 42.515 63.875 42.845 65.015 ;
        RECT 43.035 63.875 43.365 65.015 ;
        RECT 43.895 64.045 44.225 64.830 ;
        RECT 45.415 64.345 45.585 64.845 ;
        RECT 45.755 64.515 46.085 65.015 ;
        RECT 45.415 64.175 46.020 64.345 ;
        RECT 43.545 63.875 44.225 64.045 ;
        RECT 41.645 63.455 41.995 63.705 ;
        RECT 42.165 63.275 42.335 63.875 ;
        RECT 42.505 63.455 42.855 63.705 ;
        RECT 43.025 63.455 43.375 63.705 ;
        RECT 43.545 63.275 43.715 63.875 ;
        RECT 43.885 63.455 44.235 63.705 ;
        RECT 45.325 63.365 45.570 64.005 ;
        RECT 45.850 63.780 46.020 64.175 ;
        RECT 46.255 64.065 46.480 64.845 ;
        RECT 45.850 63.450 46.080 63.780 ;
        RECT 40.955 62.465 41.295 63.125 ;
        RECT 41.665 62.465 41.905 63.275 ;
        RECT 42.075 62.635 42.405 63.275 ;
        RECT 42.575 62.465 42.845 63.275 ;
        RECT 43.035 62.465 43.305 63.275 ;
        RECT 43.475 62.635 43.805 63.275 ;
        RECT 43.975 62.465 44.215 63.275 ;
        RECT 45.850 63.185 46.020 63.450 ;
        RECT 45.415 63.015 46.020 63.185 ;
        RECT 45.415 62.725 45.585 63.015 ;
        RECT 45.755 62.465 46.085 62.845 ;
        RECT 46.255 62.725 46.425 64.065 ;
        RECT 46.715 64.045 47.045 64.795 ;
        RECT 47.215 64.215 47.530 65.015 ;
        RECT 48.160 64.635 48.910 64.805 ;
        RECT 46.715 63.875 47.400 64.045 ;
        RECT 46.720 63.335 47.050 63.705 ;
        RECT 47.230 63.475 47.400 63.875 ;
        RECT 47.730 63.735 48.015 64.385 ;
        RECT 48.185 63.795 48.525 64.375 ;
        RECT 47.230 63.165 47.600 63.475 ;
        RECT 48.185 63.415 48.355 63.795 ;
        RECT 48.740 63.705 48.910 64.635 ;
        RECT 49.080 64.515 49.380 65.015 ;
        RECT 49.600 64.245 49.820 64.815 ;
        RECT 49.100 63.915 49.820 64.245 ;
        RECT 49.650 63.705 49.820 63.915 ;
        RECT 50.000 63.875 50.285 65.015 ;
        RECT 50.455 64.020 50.705 64.835 ;
        RECT 50.875 64.135 51.135 65.015 ;
        RECT 51.395 64.345 51.565 64.845 ;
        RECT 51.735 64.515 52.065 65.015 ;
        RECT 51.395 64.175 52.000 64.345 ;
        RECT 50.455 63.875 50.740 64.020 ;
        RECT 50.570 63.705 50.740 63.875 ;
        RECT 48.740 63.545 49.460 63.705 ;
        RECT 46.795 63.145 47.600 63.165 ;
        RECT 46.795 62.995 47.400 63.145 ;
        RECT 47.975 63.085 48.355 63.415 ;
        RECT 48.590 63.375 49.460 63.545 ;
        RECT 49.650 63.375 50.400 63.705 ;
        RECT 50.570 63.375 51.135 63.705 ;
        RECT 46.795 62.725 46.965 62.995 ;
        RECT 48.590 62.915 48.760 63.375 ;
        RECT 49.650 63.205 49.820 63.375 ;
        RECT 50.570 63.205 50.740 63.375 ;
        RECT 51.305 63.365 51.550 64.005 ;
        RECT 51.830 63.780 52.000 64.175 ;
        RECT 52.235 64.065 52.460 64.845 ;
        RECT 51.830 63.450 52.060 63.780 ;
        RECT 47.135 62.465 47.465 62.825 ;
        RECT 48.100 62.745 48.760 62.915 ;
        RECT 49.000 62.465 49.330 63.205 ;
        RECT 49.600 62.795 49.820 63.205 ;
        RECT 50.000 62.465 50.285 63.205 ;
        RECT 50.455 63.065 50.740 63.205 ;
        RECT 51.830 63.185 52.000 63.450 ;
        RECT 50.455 62.795 50.705 63.065 ;
        RECT 51.395 63.015 52.000 63.185 ;
        RECT 50.875 62.465 51.135 62.930 ;
        RECT 51.395 62.725 51.565 63.015 ;
        RECT 51.735 62.465 52.065 62.845 ;
        RECT 52.235 62.725 52.405 64.065 ;
        RECT 52.695 64.045 53.025 64.795 ;
        RECT 53.195 64.215 53.510 65.015 ;
        RECT 54.140 64.635 54.890 64.805 ;
        RECT 52.695 63.875 53.380 64.045 ;
        RECT 52.700 63.335 53.030 63.705 ;
        RECT 53.210 63.475 53.380 63.875 ;
        RECT 53.710 63.735 53.995 64.385 ;
        RECT 54.165 63.795 54.505 64.375 ;
        RECT 53.210 63.165 53.580 63.475 ;
        RECT 54.165 63.415 54.335 63.795 ;
        RECT 54.720 63.705 54.890 64.635 ;
        RECT 55.060 64.515 55.360 65.015 ;
        RECT 55.580 64.245 55.800 64.815 ;
        RECT 55.080 63.915 55.800 64.245 ;
        RECT 55.630 63.705 55.800 63.915 ;
        RECT 55.980 63.875 56.265 65.015 ;
        RECT 56.435 64.020 56.685 64.835 ;
        RECT 56.855 64.135 57.115 65.015 ;
        RECT 56.435 63.875 56.720 64.020 ;
        RECT 56.550 63.705 56.720 63.875 ;
        RECT 54.720 63.545 55.440 63.705 ;
        RECT 52.775 63.145 53.580 63.165 ;
        RECT 52.775 62.995 53.380 63.145 ;
        RECT 53.955 63.085 54.335 63.415 ;
        RECT 54.570 63.375 55.440 63.545 ;
        RECT 55.630 63.375 56.380 63.705 ;
        RECT 56.550 63.375 57.115 63.705 ;
        RECT 52.775 62.725 52.945 62.995 ;
        RECT 54.570 62.915 54.740 63.375 ;
        RECT 55.630 63.205 55.800 63.375 ;
        RECT 56.550 63.205 56.720 63.375 ;
        RECT 57.285 63.295 57.805 64.845 ;
        RECT 57.975 64.290 58.305 65.015 ;
        RECT 53.115 62.465 53.445 62.825 ;
        RECT 54.080 62.745 54.740 62.915 ;
        RECT 54.980 62.465 55.310 63.205 ;
        RECT 55.580 62.795 55.800 63.205 ;
        RECT 55.980 62.465 56.265 63.205 ;
        RECT 56.435 63.065 56.720 63.205 ;
        RECT 56.435 62.795 56.685 63.065 ;
        RECT 56.855 62.465 57.115 62.930 ;
        RECT 57.465 62.465 57.805 63.125 ;
        RECT 57.975 62.635 58.495 64.120 ;
        RECT 58.665 63.925 61.255 65.015 ;
        RECT 58.665 63.235 59.875 63.755 ;
        RECT 60.045 63.405 61.255 63.925 ;
        RECT 61.425 63.850 61.715 65.015 ;
        RECT 61.885 63.925 64.475 65.015 ;
        RECT 65.195 64.345 65.365 64.845 ;
        RECT 65.535 64.515 65.865 65.015 ;
        RECT 65.195 64.175 65.800 64.345 ;
        RECT 61.885 63.235 63.095 63.755 ;
        RECT 63.265 63.405 64.475 63.925 ;
        RECT 65.105 63.365 65.350 64.005 ;
        RECT 65.630 63.780 65.800 64.175 ;
        RECT 66.035 64.065 66.260 64.845 ;
        RECT 65.630 63.450 65.860 63.780 ;
        RECT 58.665 62.465 61.255 63.235 ;
        RECT 61.425 62.465 61.715 63.190 ;
        RECT 61.885 62.465 64.475 63.235 ;
        RECT 65.630 63.185 65.800 63.450 ;
        RECT 65.195 63.015 65.800 63.185 ;
        RECT 65.195 62.725 65.365 63.015 ;
        RECT 65.535 62.465 65.865 62.845 ;
        RECT 66.035 62.725 66.205 64.065 ;
        RECT 66.495 64.045 66.825 64.795 ;
        RECT 66.995 64.215 67.310 65.015 ;
        RECT 67.940 64.635 68.690 64.805 ;
        RECT 66.495 63.875 67.180 64.045 ;
        RECT 66.500 63.335 66.830 63.705 ;
        RECT 67.010 63.475 67.180 63.875 ;
        RECT 67.510 63.735 67.795 64.385 ;
        RECT 67.965 63.795 68.305 64.375 ;
        RECT 67.010 63.165 67.380 63.475 ;
        RECT 67.965 63.415 68.135 63.795 ;
        RECT 68.520 63.705 68.690 64.635 ;
        RECT 68.860 64.515 69.160 65.015 ;
        RECT 69.380 64.245 69.600 64.815 ;
        RECT 68.880 63.915 69.600 64.245 ;
        RECT 69.430 63.705 69.600 63.915 ;
        RECT 69.780 63.875 70.065 65.015 ;
        RECT 70.235 64.020 70.485 64.835 ;
        RECT 70.655 64.135 70.915 65.015 ;
        RECT 70.235 63.875 70.520 64.020 ;
        RECT 71.085 63.925 72.755 65.015 ;
        RECT 73.575 64.290 73.905 65.015 ;
        RECT 70.350 63.705 70.520 63.875 ;
        RECT 68.520 63.545 69.240 63.705 ;
        RECT 66.575 63.145 67.380 63.165 ;
        RECT 66.575 62.995 67.180 63.145 ;
        RECT 67.755 63.085 68.135 63.415 ;
        RECT 68.370 63.375 69.240 63.545 ;
        RECT 69.430 63.375 70.180 63.705 ;
        RECT 70.350 63.375 70.915 63.705 ;
        RECT 66.575 62.725 66.745 62.995 ;
        RECT 68.370 62.915 68.540 63.375 ;
        RECT 69.430 63.205 69.600 63.375 ;
        RECT 70.350 63.205 70.520 63.375 ;
        RECT 66.915 62.465 67.245 62.825 ;
        RECT 67.880 62.745 68.540 62.915 ;
        RECT 68.780 62.465 69.110 63.205 ;
        RECT 69.380 62.795 69.600 63.205 ;
        RECT 69.780 62.465 70.065 63.205 ;
        RECT 70.235 63.065 70.520 63.205 ;
        RECT 71.085 63.235 71.835 63.755 ;
        RECT 72.005 63.405 72.755 63.925 ;
        RECT 70.235 62.795 70.485 63.065 ;
        RECT 70.655 62.465 70.915 62.930 ;
        RECT 71.085 62.465 72.755 63.235 ;
        RECT 73.385 62.635 73.905 64.120 ;
        RECT 74.075 63.295 74.595 64.845 ;
        RECT 75.225 63.295 75.745 64.845 ;
        RECT 75.915 64.290 76.245 65.015 ;
        RECT 76.795 64.290 77.125 65.015 ;
        RECT 74.075 62.465 74.415 63.125 ;
        RECT 75.405 62.465 75.745 63.125 ;
        RECT 75.915 62.635 76.435 64.120 ;
        RECT 76.605 62.635 77.125 64.120 ;
        RECT 77.295 63.295 77.815 64.845 ;
        RECT 78.075 64.345 78.245 64.845 ;
        RECT 78.415 64.515 78.745 65.015 ;
        RECT 78.075 64.175 78.680 64.345 ;
        RECT 77.985 63.365 78.230 64.005 ;
        RECT 78.510 63.780 78.680 64.175 ;
        RECT 78.915 64.065 79.140 64.845 ;
        RECT 78.510 63.450 78.740 63.780 ;
        RECT 78.510 63.185 78.680 63.450 ;
        RECT 77.295 62.465 77.635 63.125 ;
        RECT 78.075 63.015 78.680 63.185 ;
        RECT 78.075 62.725 78.245 63.015 ;
        RECT 78.415 62.465 78.745 62.845 ;
        RECT 78.915 62.725 79.085 64.065 ;
        RECT 79.375 64.045 79.705 64.795 ;
        RECT 79.875 64.215 80.190 65.015 ;
        RECT 80.820 64.635 81.570 64.805 ;
        RECT 79.375 63.875 80.060 64.045 ;
        RECT 79.380 63.335 79.710 63.705 ;
        RECT 79.890 63.475 80.060 63.875 ;
        RECT 80.390 63.735 80.675 64.385 ;
        RECT 80.845 63.795 81.185 64.375 ;
        RECT 79.890 63.165 80.260 63.475 ;
        RECT 80.845 63.415 81.015 63.795 ;
        RECT 81.400 63.705 81.570 64.635 ;
        RECT 81.740 64.515 82.040 65.015 ;
        RECT 82.260 64.245 82.480 64.815 ;
        RECT 81.760 63.915 82.480 64.245 ;
        RECT 82.310 63.705 82.480 63.915 ;
        RECT 82.660 63.875 82.945 65.015 ;
        RECT 83.115 64.020 83.365 64.835 ;
        RECT 83.535 64.135 83.795 65.015 ;
        RECT 83.975 64.045 84.305 64.830 ;
        RECT 83.115 63.875 83.400 64.020 ;
        RECT 83.975 63.875 84.655 64.045 ;
        RECT 84.835 63.875 85.165 65.015 ;
        RECT 85.355 64.045 85.685 64.830 ;
        RECT 85.355 63.875 86.035 64.045 ;
        RECT 86.215 63.875 86.545 65.015 ;
        RECT 83.230 63.705 83.400 63.875 ;
        RECT 81.400 63.545 82.120 63.705 ;
        RECT 79.455 63.145 80.260 63.165 ;
        RECT 79.455 62.995 80.060 63.145 ;
        RECT 80.635 63.085 81.015 63.415 ;
        RECT 81.250 63.375 82.120 63.545 ;
        RECT 82.310 63.375 83.060 63.705 ;
        RECT 83.230 63.375 83.795 63.705 ;
        RECT 83.965 63.455 84.315 63.705 ;
        RECT 79.455 62.725 79.625 62.995 ;
        RECT 81.250 62.915 81.420 63.375 ;
        RECT 82.310 63.205 82.480 63.375 ;
        RECT 83.230 63.205 83.400 63.375 ;
        RECT 84.485 63.275 84.655 63.875 ;
        RECT 84.825 63.455 85.175 63.705 ;
        RECT 85.345 63.455 85.695 63.705 ;
        RECT 85.865 63.275 86.035 63.875 ;
        RECT 87.185 63.850 87.475 65.015 ;
        RECT 86.205 63.455 86.555 63.705 ;
        RECT 87.645 63.295 88.165 64.845 ;
        RECT 88.335 64.290 88.665 65.015 ;
        RECT 79.795 62.465 80.125 62.825 ;
        RECT 80.760 62.745 81.420 62.915 ;
        RECT 81.660 62.465 81.990 63.205 ;
        RECT 82.260 62.795 82.480 63.205 ;
        RECT 82.660 62.465 82.945 63.205 ;
        RECT 83.115 63.065 83.400 63.205 ;
        RECT 83.115 62.795 83.365 63.065 ;
        RECT 83.535 62.465 83.795 62.930 ;
        RECT 83.985 62.465 84.225 63.275 ;
        RECT 84.395 62.635 84.725 63.275 ;
        RECT 84.895 62.465 85.165 63.275 ;
        RECT 85.365 62.465 85.605 63.275 ;
        RECT 85.775 62.635 86.105 63.275 ;
        RECT 86.275 62.465 86.545 63.275 ;
        RECT 87.185 62.465 87.475 63.190 ;
        RECT 87.825 62.465 88.165 63.125 ;
        RECT 88.335 62.635 88.855 64.120 ;
        RECT 89.025 63.925 90.235 65.015 ;
        RECT 89.025 63.215 89.545 63.755 ;
        RECT 89.715 63.385 90.235 63.925 ;
        RECT 90.405 63.295 90.925 64.845 ;
        RECT 91.095 64.290 91.425 65.015 ;
        RECT 89.025 62.465 90.235 63.215 ;
        RECT 90.585 62.465 90.925 63.125 ;
        RECT 91.095 62.635 91.615 64.120 ;
        RECT 92.705 63.295 93.225 64.845 ;
        RECT 93.395 64.290 93.725 65.015 ;
        RECT 92.885 62.465 93.225 63.125 ;
        RECT 93.395 62.635 93.915 64.120 ;
        RECT 94.085 63.925 95.755 65.015 ;
        RECT 96.015 64.345 96.185 64.845 ;
        RECT 96.355 64.515 96.685 65.015 ;
        RECT 96.015 64.175 96.620 64.345 ;
        RECT 94.085 63.235 94.835 63.755 ;
        RECT 95.005 63.405 95.755 63.925 ;
        RECT 95.925 63.365 96.170 64.005 ;
        RECT 96.450 63.780 96.620 64.175 ;
        RECT 96.855 64.065 97.080 64.845 ;
        RECT 96.450 63.450 96.680 63.780 ;
        RECT 94.085 62.465 95.755 63.235 ;
        RECT 96.450 63.185 96.620 63.450 ;
        RECT 96.015 63.015 96.620 63.185 ;
        RECT 96.015 62.725 96.185 63.015 ;
        RECT 96.355 62.465 96.685 62.845 ;
        RECT 96.855 62.725 97.025 64.065 ;
        RECT 97.315 64.045 97.645 64.795 ;
        RECT 97.815 64.215 98.130 65.015 ;
        RECT 98.760 64.635 99.510 64.805 ;
        RECT 97.315 63.875 98.000 64.045 ;
        RECT 97.320 63.335 97.650 63.705 ;
        RECT 97.830 63.475 98.000 63.875 ;
        RECT 98.330 63.735 98.615 64.385 ;
        RECT 98.785 63.795 99.125 64.375 ;
        RECT 97.830 63.165 98.200 63.475 ;
        RECT 98.785 63.415 98.955 63.795 ;
        RECT 99.340 63.705 99.510 64.635 ;
        RECT 99.680 64.515 99.980 65.015 ;
        RECT 100.200 64.245 100.420 64.815 ;
        RECT 99.700 63.915 100.420 64.245 ;
        RECT 100.250 63.705 100.420 63.915 ;
        RECT 100.600 63.875 100.885 65.015 ;
        RECT 101.055 64.020 101.305 64.835 ;
        RECT 101.475 64.135 101.735 65.015 ;
        RECT 101.055 63.875 101.340 64.020 ;
        RECT 101.170 63.705 101.340 63.875 ;
        RECT 99.340 63.545 100.060 63.705 ;
        RECT 97.395 63.145 98.200 63.165 ;
        RECT 97.395 62.995 98.000 63.145 ;
        RECT 98.575 63.085 98.955 63.415 ;
        RECT 99.190 63.375 100.060 63.545 ;
        RECT 100.250 63.375 101.000 63.705 ;
        RECT 101.170 63.375 101.735 63.705 ;
        RECT 97.395 62.725 97.565 62.995 ;
        RECT 99.190 62.915 99.360 63.375 ;
        RECT 100.250 63.205 100.420 63.375 ;
        RECT 101.170 63.205 101.340 63.375 ;
        RECT 101.905 63.295 102.425 64.845 ;
        RECT 102.595 64.290 102.925 65.015 ;
        RECT 103.475 64.290 103.805 65.015 ;
        RECT 97.735 62.465 98.065 62.825 ;
        RECT 98.700 62.745 99.360 62.915 ;
        RECT 99.600 62.465 99.930 63.205 ;
        RECT 100.200 62.795 100.420 63.205 ;
        RECT 100.600 62.465 100.885 63.205 ;
        RECT 101.055 63.065 101.340 63.205 ;
        RECT 101.055 62.795 101.305 63.065 ;
        RECT 101.475 62.465 101.735 62.930 ;
        RECT 102.085 62.465 102.425 63.125 ;
        RECT 102.595 62.635 103.115 64.120 ;
        RECT 103.285 62.635 103.805 64.120 ;
        RECT 103.975 63.295 104.495 64.845 ;
        RECT 104.665 63.925 106.335 65.015 ;
        RECT 104.665 63.235 105.415 63.755 ;
        RECT 105.585 63.405 106.335 63.925 ;
        RECT 106.965 63.295 107.485 64.845 ;
        RECT 107.655 64.290 107.985 65.015 ;
        RECT 108.535 64.290 108.865 65.015 ;
        RECT 103.975 62.465 104.315 63.125 ;
        RECT 104.665 62.465 106.335 63.235 ;
        RECT 107.145 62.465 107.485 63.125 ;
        RECT 107.655 62.635 108.175 64.120 ;
        RECT 108.345 62.635 108.865 64.120 ;
        RECT 109.035 63.295 109.555 64.845 ;
        RECT 109.725 63.925 112.315 65.015 ;
        RECT 109.725 63.235 110.935 63.755 ;
        RECT 111.105 63.405 112.315 63.925 ;
        RECT 112.945 63.850 113.235 65.015 ;
        RECT 113.405 63.295 113.925 64.845 ;
        RECT 114.095 64.290 114.425 65.015 ;
        RECT 114.975 64.290 115.305 65.015 ;
        RECT 109.035 62.465 109.375 63.125 ;
        RECT 109.725 62.465 112.315 63.235 ;
        RECT 112.945 62.465 113.235 63.190 ;
        RECT 113.585 62.465 113.925 63.125 ;
        RECT 114.095 62.635 114.615 64.120 ;
        RECT 114.785 62.635 115.305 64.120 ;
        RECT 115.475 63.295 115.995 64.845 ;
        RECT 116.355 64.290 116.685 65.015 ;
        RECT 115.475 62.465 115.815 63.125 ;
        RECT 116.165 62.635 116.685 64.120 ;
        RECT 116.855 63.295 117.375 64.845 ;
        RECT 117.635 64.345 117.805 64.845 ;
        RECT 117.975 64.515 118.305 65.015 ;
        RECT 117.635 64.175 118.240 64.345 ;
        RECT 117.545 63.365 117.790 64.005 ;
        RECT 118.070 63.780 118.240 64.175 ;
        RECT 118.475 64.065 118.700 64.845 ;
        RECT 118.070 63.450 118.300 63.780 ;
        RECT 118.070 63.185 118.240 63.450 ;
        RECT 116.855 62.465 117.195 63.125 ;
        RECT 117.635 63.015 118.240 63.185 ;
        RECT 117.635 62.725 117.805 63.015 ;
        RECT 117.975 62.465 118.305 62.845 ;
        RECT 118.475 62.725 118.645 64.065 ;
        RECT 118.935 64.045 119.265 64.795 ;
        RECT 119.435 64.215 119.750 65.015 ;
        RECT 120.380 64.635 121.130 64.805 ;
        RECT 118.935 63.875 119.620 64.045 ;
        RECT 118.940 63.335 119.270 63.705 ;
        RECT 119.450 63.475 119.620 63.875 ;
        RECT 119.950 63.735 120.235 64.385 ;
        RECT 120.405 63.795 120.745 64.375 ;
        RECT 119.450 63.165 119.820 63.475 ;
        RECT 120.405 63.415 120.575 63.795 ;
        RECT 120.960 63.705 121.130 64.635 ;
        RECT 121.300 64.515 121.600 65.015 ;
        RECT 121.820 64.245 122.040 64.815 ;
        RECT 121.320 63.915 122.040 64.245 ;
        RECT 121.870 63.705 122.040 63.915 ;
        RECT 122.220 63.875 122.505 65.015 ;
        RECT 122.675 64.020 122.925 64.835 ;
        RECT 123.095 64.135 123.355 65.015 ;
        RECT 122.675 63.875 122.960 64.020 ;
        RECT 124.455 63.875 124.785 65.015 ;
        RECT 125.315 64.045 125.645 64.830 ;
        RECT 125.915 64.345 126.085 64.845 ;
        RECT 126.255 64.515 126.585 65.015 ;
        RECT 125.915 64.175 126.520 64.345 ;
        RECT 124.965 63.875 125.645 64.045 ;
        RECT 122.790 63.705 122.960 63.875 ;
        RECT 120.960 63.545 121.680 63.705 ;
        RECT 119.015 63.145 119.820 63.165 ;
        RECT 119.015 62.995 119.620 63.145 ;
        RECT 120.195 63.085 120.575 63.415 ;
        RECT 120.810 63.375 121.680 63.545 ;
        RECT 121.870 63.375 122.620 63.705 ;
        RECT 122.790 63.375 123.355 63.705 ;
        RECT 124.445 63.455 124.795 63.705 ;
        RECT 119.015 62.725 119.185 62.995 ;
        RECT 120.810 62.915 120.980 63.375 ;
        RECT 121.870 63.205 122.040 63.375 ;
        RECT 122.790 63.205 122.960 63.375 ;
        RECT 124.965 63.275 125.135 63.875 ;
        RECT 125.305 63.455 125.655 63.705 ;
        RECT 125.825 63.365 126.070 64.005 ;
        RECT 126.350 63.780 126.520 64.175 ;
        RECT 126.755 64.065 126.980 64.845 ;
        RECT 126.350 63.450 126.580 63.780 ;
        RECT 119.355 62.465 119.685 62.825 ;
        RECT 120.320 62.745 120.980 62.915 ;
        RECT 121.220 62.465 121.550 63.205 ;
        RECT 121.820 62.795 122.040 63.205 ;
        RECT 122.220 62.465 122.505 63.205 ;
        RECT 122.675 63.065 122.960 63.205 ;
        RECT 122.675 62.795 122.925 63.065 ;
        RECT 123.095 62.465 123.355 62.930 ;
        RECT 124.455 62.465 124.725 63.275 ;
        RECT 124.895 62.635 125.225 63.275 ;
        RECT 125.395 62.465 125.635 63.275 ;
        RECT 126.350 63.185 126.520 63.450 ;
        RECT 125.915 63.015 126.520 63.185 ;
        RECT 125.915 62.725 126.085 63.015 ;
        RECT 126.255 62.465 126.585 62.845 ;
        RECT 126.755 62.725 126.925 64.065 ;
        RECT 127.215 64.045 127.545 64.795 ;
        RECT 127.715 64.215 128.030 65.015 ;
        RECT 128.660 64.635 129.410 64.805 ;
        RECT 127.215 63.875 127.900 64.045 ;
        RECT 127.220 63.335 127.550 63.705 ;
        RECT 127.730 63.475 127.900 63.875 ;
        RECT 128.230 63.735 128.515 64.385 ;
        RECT 128.685 63.795 129.025 64.375 ;
        RECT 127.730 63.165 128.100 63.475 ;
        RECT 128.685 63.415 128.855 63.795 ;
        RECT 129.240 63.705 129.410 64.635 ;
        RECT 129.580 64.515 129.880 65.015 ;
        RECT 130.100 64.245 130.320 64.815 ;
        RECT 129.600 63.915 130.320 64.245 ;
        RECT 130.150 63.705 130.320 63.915 ;
        RECT 130.500 63.875 130.785 65.015 ;
        RECT 130.955 64.020 131.205 64.835 ;
        RECT 131.375 64.135 131.635 65.015 ;
        RECT 130.955 63.875 131.240 64.020 ;
        RECT 131.070 63.705 131.240 63.875 ;
        RECT 129.240 63.545 129.960 63.705 ;
        RECT 127.295 63.145 128.100 63.165 ;
        RECT 127.295 62.995 127.900 63.145 ;
        RECT 128.475 63.085 128.855 63.415 ;
        RECT 129.090 63.375 129.960 63.545 ;
        RECT 130.150 63.375 130.900 63.705 ;
        RECT 131.070 63.375 131.635 63.705 ;
        RECT 127.295 62.725 127.465 62.995 ;
        RECT 129.090 62.915 129.260 63.375 ;
        RECT 130.150 63.205 130.320 63.375 ;
        RECT 131.070 63.205 131.240 63.375 ;
        RECT 131.805 63.295 132.325 64.845 ;
        RECT 132.495 64.290 132.825 65.015 ;
        RECT 127.635 62.465 127.965 62.825 ;
        RECT 128.600 62.745 129.260 62.915 ;
        RECT 129.500 62.465 129.830 63.205 ;
        RECT 130.100 62.795 130.320 63.205 ;
        RECT 130.500 62.465 130.785 63.205 ;
        RECT 130.955 63.065 131.240 63.205 ;
        RECT 130.955 62.795 131.205 63.065 ;
        RECT 131.375 62.465 131.635 62.930 ;
        RECT 131.985 62.465 132.325 63.125 ;
        RECT 132.495 62.635 133.015 64.120 ;
        RECT 133.185 63.295 133.705 64.845 ;
        RECT 133.875 64.290 134.205 65.015 ;
        RECT 134.755 64.290 135.085 65.015 ;
        RECT 133.365 62.465 133.705 63.125 ;
        RECT 133.875 62.635 134.395 64.120 ;
        RECT 134.565 62.635 135.085 64.120 ;
        RECT 135.255 63.295 135.775 64.845 ;
        RECT 135.945 63.925 137.155 65.015 ;
        RECT 137.515 64.290 137.845 65.015 ;
        RECT 135.945 63.215 136.465 63.755 ;
        RECT 136.635 63.385 137.155 63.925 ;
        RECT 135.255 62.465 135.595 63.125 ;
        RECT 135.945 62.465 137.155 63.215 ;
        RECT 137.325 62.635 137.845 64.120 ;
        RECT 138.015 63.295 138.535 64.845 ;
        RECT 138.705 63.850 138.995 65.015 ;
        RECT 139.715 64.345 139.885 64.845 ;
        RECT 140.055 64.515 140.385 65.015 ;
        RECT 139.715 64.175 140.320 64.345 ;
        RECT 139.625 63.365 139.870 64.005 ;
        RECT 140.150 63.780 140.320 64.175 ;
        RECT 140.555 64.065 140.780 64.845 ;
        RECT 140.150 63.450 140.380 63.780 ;
        RECT 138.015 62.465 138.355 63.125 ;
        RECT 138.705 62.465 138.995 63.190 ;
        RECT 140.150 63.185 140.320 63.450 ;
        RECT 139.715 63.015 140.320 63.185 ;
        RECT 139.715 62.725 139.885 63.015 ;
        RECT 140.055 62.465 140.385 62.845 ;
        RECT 140.555 62.725 140.725 64.065 ;
        RECT 141.015 64.045 141.345 64.795 ;
        RECT 141.515 64.215 141.830 65.015 ;
        RECT 142.460 64.635 143.210 64.805 ;
        RECT 141.015 63.875 141.700 64.045 ;
        RECT 141.020 63.335 141.350 63.705 ;
        RECT 141.530 63.475 141.700 63.875 ;
        RECT 142.030 63.735 142.315 64.385 ;
        RECT 142.485 63.795 142.825 64.375 ;
        RECT 141.530 63.165 141.900 63.475 ;
        RECT 142.485 63.415 142.655 63.795 ;
        RECT 143.040 63.705 143.210 64.635 ;
        RECT 143.380 64.515 143.680 65.015 ;
        RECT 143.900 64.245 144.120 64.815 ;
        RECT 143.400 63.915 144.120 64.245 ;
        RECT 143.950 63.705 144.120 63.915 ;
        RECT 144.300 63.875 144.585 65.015 ;
        RECT 144.755 64.020 145.005 64.835 ;
        RECT 145.175 64.135 145.435 65.015 ;
        RECT 144.755 63.875 145.040 64.020 ;
        RECT 144.870 63.705 145.040 63.875 ;
        RECT 143.040 63.545 143.760 63.705 ;
        RECT 141.095 63.145 141.900 63.165 ;
        RECT 141.095 62.995 141.700 63.145 ;
        RECT 142.275 63.085 142.655 63.415 ;
        RECT 142.890 63.375 143.760 63.545 ;
        RECT 143.950 63.375 144.700 63.705 ;
        RECT 144.870 63.375 145.435 63.705 ;
        RECT 141.095 62.725 141.265 62.995 ;
        RECT 142.890 62.915 143.060 63.375 ;
        RECT 143.950 63.205 144.120 63.375 ;
        RECT 144.870 63.205 145.040 63.375 ;
        RECT 145.605 63.295 146.125 64.845 ;
        RECT 146.295 64.290 146.625 65.015 ;
        RECT 141.435 62.465 141.765 62.825 ;
        RECT 142.400 62.745 143.060 62.915 ;
        RECT 143.300 62.465 143.630 63.205 ;
        RECT 143.900 62.795 144.120 63.205 ;
        RECT 144.300 62.465 144.585 63.205 ;
        RECT 144.755 63.065 145.040 63.205 ;
        RECT 144.755 62.795 145.005 63.065 ;
        RECT 145.175 62.465 145.435 62.930 ;
        RECT 145.785 62.465 146.125 63.125 ;
        RECT 146.295 62.635 146.815 64.120 ;
        RECT 146.985 63.295 147.505 64.845 ;
        RECT 147.675 64.290 148.005 65.015 ;
        RECT 148.365 64.580 153.710 65.015 ;
        RECT 147.165 62.465 147.505 63.125 ;
        RECT 147.675 62.635 148.195 64.120 ;
        RECT 149.950 63.010 150.290 63.840 ;
        RECT 151.770 63.330 152.120 64.580 ;
        RECT 153.885 63.925 155.555 65.015 ;
        RECT 153.885 63.235 154.635 63.755 ;
        RECT 154.805 63.405 155.555 63.925 ;
        RECT 155.725 63.925 156.935 65.015 ;
        RECT 155.725 63.385 156.245 63.925 ;
        RECT 148.365 62.465 153.710 63.010 ;
        RECT 153.885 62.465 155.555 63.235 ;
        RECT 156.415 63.215 156.935 63.755 ;
        RECT 155.725 62.465 156.935 63.215 ;
        RECT 22.700 62.295 157.020 62.465 ;
        RECT 22.785 61.545 23.995 62.295 ;
        RECT 24.715 61.745 24.885 62.035 ;
        RECT 25.055 61.915 25.385 62.295 ;
        RECT 24.715 61.575 25.320 61.745 ;
        RECT 22.785 61.005 23.305 61.545 ;
        RECT 23.475 60.835 23.995 61.375 ;
        RECT 22.785 59.745 23.995 60.835 ;
        RECT 24.625 60.755 24.870 61.395 ;
        RECT 25.150 61.310 25.320 61.575 ;
        RECT 25.150 60.980 25.380 61.310 ;
        RECT 25.150 60.585 25.320 60.980 ;
        RECT 24.715 60.415 25.320 60.585 ;
        RECT 25.555 60.695 25.725 62.035 ;
        RECT 26.095 61.765 26.265 62.035 ;
        RECT 26.435 61.935 26.765 62.295 ;
        RECT 27.400 61.845 28.060 62.015 ;
        RECT 26.095 61.615 26.700 61.765 ;
        RECT 26.095 61.595 26.900 61.615 ;
        RECT 26.020 61.055 26.350 61.425 ;
        RECT 26.530 61.285 26.900 61.595 ;
        RECT 27.275 61.345 27.655 61.675 ;
        RECT 26.530 60.885 26.700 61.285 ;
        RECT 26.015 60.715 26.700 60.885 ;
        RECT 24.715 59.915 24.885 60.415 ;
        RECT 25.055 59.745 25.385 60.245 ;
        RECT 25.555 59.915 25.780 60.695 ;
        RECT 26.015 59.965 26.345 60.715 ;
        RECT 26.515 59.745 26.830 60.545 ;
        RECT 27.030 60.375 27.315 61.025 ;
        RECT 27.485 60.965 27.655 61.345 ;
        RECT 27.890 61.385 28.060 61.845 ;
        RECT 28.300 61.555 28.630 62.295 ;
        RECT 28.900 61.555 29.120 61.965 ;
        RECT 29.300 61.555 29.585 62.295 ;
        RECT 29.755 61.695 30.005 61.965 ;
        RECT 30.175 61.830 30.435 62.295 ;
        RECT 30.605 61.830 30.865 62.295 ;
        RECT 31.035 61.695 31.285 61.965 ;
        RECT 29.755 61.555 30.040 61.695 ;
        RECT 28.950 61.385 29.120 61.555 ;
        RECT 29.870 61.385 30.040 61.555 ;
        RECT 31.000 61.555 31.285 61.695 ;
        RECT 31.455 61.555 31.740 62.295 ;
        RECT 31.920 61.555 32.140 61.965 ;
        RECT 32.410 61.555 32.740 62.295 ;
        RECT 32.980 61.845 33.640 62.015 ;
        RECT 34.275 61.935 34.605 62.295 ;
        RECT 31.000 61.385 31.170 61.555 ;
        RECT 31.920 61.385 32.090 61.555 ;
        RECT 32.980 61.385 33.150 61.845 ;
        RECT 34.775 61.765 34.945 62.035 ;
        RECT 27.890 61.215 28.760 61.385 ;
        RECT 28.040 61.055 28.760 61.215 ;
        RECT 28.950 61.055 29.700 61.385 ;
        RECT 29.870 61.055 30.435 61.385 ;
        RECT 30.605 61.055 31.170 61.385 ;
        RECT 31.340 61.055 32.090 61.385 ;
        RECT 32.280 61.215 33.150 61.385 ;
        RECT 33.385 61.345 33.765 61.675 ;
        RECT 34.340 61.615 34.945 61.765 ;
        RECT 34.140 61.595 34.945 61.615 ;
        RECT 32.280 61.055 33.000 61.215 ;
        RECT 27.485 60.385 27.825 60.965 ;
        RECT 28.040 60.125 28.210 61.055 ;
        RECT 28.950 60.845 29.120 61.055 ;
        RECT 29.870 60.885 30.040 61.055 ;
        RECT 28.400 60.515 29.120 60.845 ;
        RECT 27.460 59.955 28.210 60.125 ;
        RECT 28.380 59.745 28.680 60.245 ;
        RECT 28.900 59.945 29.120 60.515 ;
        RECT 29.300 59.745 29.585 60.885 ;
        RECT 29.755 60.740 30.040 60.885 ;
        RECT 31.000 60.885 31.170 61.055 ;
        RECT 31.000 60.740 31.285 60.885 ;
        RECT 29.755 59.925 30.005 60.740 ;
        RECT 30.175 59.745 30.435 60.625 ;
        RECT 30.605 59.745 30.865 60.625 ;
        RECT 31.035 59.925 31.285 60.740 ;
        RECT 31.455 59.745 31.740 60.885 ;
        RECT 31.920 60.845 32.090 61.055 ;
        RECT 31.920 60.515 32.640 60.845 ;
        RECT 31.920 59.945 32.140 60.515 ;
        RECT 32.360 59.745 32.660 60.245 ;
        RECT 32.830 60.125 33.000 61.055 ;
        RECT 33.385 60.965 33.555 61.345 ;
        RECT 34.140 61.285 34.510 61.595 ;
        RECT 33.215 60.385 33.555 60.965 ;
        RECT 33.725 60.375 34.010 61.025 ;
        RECT 34.340 60.885 34.510 61.285 ;
        RECT 34.690 61.055 35.020 61.425 ;
        RECT 34.340 60.715 35.025 60.885 ;
        RECT 32.830 59.955 33.580 60.125 ;
        RECT 34.210 59.745 34.525 60.545 ;
        RECT 34.695 59.965 35.025 60.715 ;
        RECT 35.315 60.695 35.485 62.035 ;
        RECT 35.655 61.915 35.985 62.295 ;
        RECT 36.155 61.745 36.325 62.035 ;
        RECT 35.720 61.575 36.325 61.745 ;
        RECT 36.675 61.745 36.845 62.035 ;
        RECT 37.015 61.915 37.345 62.295 ;
        RECT 36.675 61.575 37.280 61.745 ;
        RECT 35.720 61.310 35.890 61.575 ;
        RECT 35.660 60.980 35.890 61.310 ;
        RECT 35.260 59.915 35.485 60.695 ;
        RECT 35.720 60.585 35.890 60.980 ;
        RECT 36.170 60.755 36.415 61.395 ;
        RECT 36.585 60.755 36.830 61.395 ;
        RECT 37.110 61.310 37.280 61.575 ;
        RECT 37.110 60.980 37.340 61.310 ;
        RECT 37.110 60.585 37.280 60.980 ;
        RECT 35.720 60.415 36.325 60.585 ;
        RECT 35.655 59.745 35.985 60.245 ;
        RECT 36.155 59.915 36.325 60.415 ;
        RECT 36.675 60.415 37.280 60.585 ;
        RECT 37.515 60.695 37.685 62.035 ;
        RECT 38.055 61.765 38.225 62.035 ;
        RECT 38.395 61.935 38.725 62.295 ;
        RECT 39.360 61.845 40.020 62.015 ;
        RECT 38.055 61.615 38.660 61.765 ;
        RECT 38.055 61.595 38.860 61.615 ;
        RECT 37.980 61.055 38.310 61.425 ;
        RECT 38.490 61.285 38.860 61.595 ;
        RECT 39.235 61.345 39.615 61.675 ;
        RECT 38.490 60.885 38.660 61.285 ;
        RECT 37.975 60.715 38.660 60.885 ;
        RECT 36.675 59.915 36.845 60.415 ;
        RECT 37.015 59.745 37.345 60.245 ;
        RECT 37.515 59.915 37.740 60.695 ;
        RECT 37.975 59.965 38.305 60.715 ;
        RECT 38.475 59.745 38.790 60.545 ;
        RECT 38.990 60.375 39.275 61.025 ;
        RECT 39.445 60.965 39.615 61.345 ;
        RECT 39.850 61.385 40.020 61.845 ;
        RECT 40.260 61.555 40.590 62.295 ;
        RECT 40.860 61.555 41.080 61.965 ;
        RECT 41.260 61.555 41.545 62.295 ;
        RECT 41.715 61.695 41.965 61.965 ;
        RECT 42.135 61.830 42.395 62.295 ;
        RECT 42.655 61.745 42.825 62.035 ;
        RECT 42.995 61.915 43.325 62.295 ;
        RECT 41.715 61.555 42.000 61.695 ;
        RECT 42.655 61.575 43.260 61.745 ;
        RECT 40.910 61.385 41.080 61.555 ;
        RECT 41.830 61.385 42.000 61.555 ;
        RECT 39.850 61.215 40.720 61.385 ;
        RECT 40.000 61.055 40.720 61.215 ;
        RECT 40.910 61.055 41.660 61.385 ;
        RECT 41.830 61.055 42.395 61.385 ;
        RECT 39.445 60.385 39.785 60.965 ;
        RECT 40.000 60.125 40.170 61.055 ;
        RECT 40.910 60.845 41.080 61.055 ;
        RECT 41.830 60.885 42.000 61.055 ;
        RECT 40.360 60.515 41.080 60.845 ;
        RECT 39.420 59.955 40.170 60.125 ;
        RECT 40.340 59.745 40.640 60.245 ;
        RECT 40.860 59.945 41.080 60.515 ;
        RECT 41.260 59.745 41.545 60.885 ;
        RECT 41.715 60.740 42.000 60.885 ;
        RECT 42.565 60.755 42.810 61.395 ;
        RECT 43.090 61.310 43.260 61.575 ;
        RECT 43.090 60.980 43.320 61.310 ;
        RECT 41.715 59.925 41.965 60.740 ;
        RECT 42.135 59.745 42.395 60.625 ;
        RECT 43.090 60.585 43.260 60.980 ;
        RECT 42.655 60.415 43.260 60.585 ;
        RECT 43.495 60.695 43.665 62.035 ;
        RECT 44.035 61.765 44.205 62.035 ;
        RECT 44.375 61.935 44.705 62.295 ;
        RECT 45.340 61.845 46.000 62.015 ;
        RECT 44.035 61.615 44.640 61.765 ;
        RECT 44.035 61.595 44.840 61.615 ;
        RECT 43.960 61.055 44.290 61.425 ;
        RECT 44.470 61.285 44.840 61.595 ;
        RECT 45.215 61.345 45.595 61.675 ;
        RECT 44.470 60.885 44.640 61.285 ;
        RECT 43.955 60.715 44.640 60.885 ;
        RECT 42.655 59.915 42.825 60.415 ;
        RECT 42.995 59.745 43.325 60.245 ;
        RECT 43.495 59.915 43.720 60.695 ;
        RECT 43.955 59.965 44.285 60.715 ;
        RECT 44.455 59.745 44.770 60.545 ;
        RECT 44.970 60.375 45.255 61.025 ;
        RECT 45.425 60.965 45.595 61.345 ;
        RECT 45.830 61.385 46.000 61.845 ;
        RECT 46.240 61.555 46.570 62.295 ;
        RECT 46.840 61.555 47.060 61.965 ;
        RECT 47.240 61.555 47.525 62.295 ;
        RECT 47.695 61.695 47.945 61.965 ;
        RECT 48.115 61.830 48.375 62.295 ;
        RECT 47.695 61.555 47.980 61.695 ;
        RECT 48.545 61.570 48.835 62.295 ;
        RECT 46.890 61.385 47.060 61.555 ;
        RECT 47.810 61.385 47.980 61.555 ;
        RECT 45.830 61.215 46.700 61.385 ;
        RECT 45.980 61.055 46.700 61.215 ;
        RECT 46.890 61.055 47.640 61.385 ;
        RECT 47.810 61.055 48.375 61.385 ;
        RECT 45.425 60.385 45.765 60.965 ;
        RECT 45.980 60.125 46.150 61.055 ;
        RECT 46.890 60.845 47.060 61.055 ;
        RECT 47.810 60.885 47.980 61.055 ;
        RECT 46.340 60.515 47.060 60.845 ;
        RECT 45.400 59.955 46.150 60.125 ;
        RECT 46.320 59.745 46.620 60.245 ;
        RECT 46.840 59.945 47.060 60.515 ;
        RECT 47.240 59.745 47.525 60.885 ;
        RECT 47.695 60.740 47.980 60.885 ;
        RECT 47.695 59.925 47.945 60.740 ;
        RECT 48.115 59.745 48.375 60.625 ;
        RECT 48.545 59.745 48.835 60.910 ;
        RECT 49.005 60.640 49.525 62.125 ;
        RECT 49.695 61.635 50.035 62.295 ;
        RECT 50.565 61.635 50.905 62.295 ;
        RECT 49.195 59.745 49.525 60.470 ;
        RECT 49.695 59.915 50.215 61.465 ;
        RECT 50.385 59.915 50.905 61.465 ;
        RECT 51.075 60.640 51.595 62.125 ;
        RECT 52.225 60.640 52.745 62.125 ;
        RECT 52.915 61.635 53.255 62.295 ;
        RECT 53.695 61.745 53.865 62.035 ;
        RECT 54.035 61.915 54.365 62.295 ;
        RECT 53.695 61.575 54.300 61.745 ;
        RECT 51.075 59.745 51.405 60.470 ;
        RECT 52.415 59.745 52.745 60.470 ;
        RECT 52.915 59.915 53.435 61.465 ;
        RECT 53.605 60.755 53.850 61.395 ;
        RECT 54.130 61.310 54.300 61.575 ;
        RECT 54.130 60.980 54.360 61.310 ;
        RECT 54.130 60.585 54.300 60.980 ;
        RECT 53.695 60.415 54.300 60.585 ;
        RECT 54.535 60.695 54.705 62.035 ;
        RECT 55.075 61.765 55.245 62.035 ;
        RECT 55.415 61.935 55.745 62.295 ;
        RECT 56.380 61.845 57.040 62.015 ;
        RECT 55.075 61.615 55.680 61.765 ;
        RECT 55.075 61.595 55.880 61.615 ;
        RECT 55.000 61.055 55.330 61.425 ;
        RECT 55.510 61.285 55.880 61.595 ;
        RECT 56.255 61.345 56.635 61.675 ;
        RECT 55.510 60.885 55.680 61.285 ;
        RECT 54.995 60.715 55.680 60.885 ;
        RECT 53.695 59.915 53.865 60.415 ;
        RECT 54.035 59.745 54.365 60.245 ;
        RECT 54.535 59.915 54.760 60.695 ;
        RECT 54.995 59.965 55.325 60.715 ;
        RECT 55.495 59.745 55.810 60.545 ;
        RECT 56.010 60.375 56.295 61.025 ;
        RECT 56.465 60.965 56.635 61.345 ;
        RECT 56.870 61.385 57.040 61.845 ;
        RECT 57.280 61.555 57.610 62.295 ;
        RECT 57.880 61.555 58.100 61.965 ;
        RECT 58.280 61.555 58.565 62.295 ;
        RECT 58.735 61.695 58.985 61.965 ;
        RECT 59.155 61.830 59.415 62.295 ;
        RECT 59.675 61.745 59.845 62.035 ;
        RECT 60.015 61.915 60.345 62.295 ;
        RECT 58.735 61.555 59.020 61.695 ;
        RECT 59.675 61.575 60.280 61.745 ;
        RECT 57.930 61.385 58.100 61.555 ;
        RECT 58.850 61.385 59.020 61.555 ;
        RECT 56.870 61.215 57.740 61.385 ;
        RECT 57.020 61.055 57.740 61.215 ;
        RECT 57.930 61.055 58.680 61.385 ;
        RECT 58.850 61.055 59.415 61.385 ;
        RECT 56.465 60.385 56.805 60.965 ;
        RECT 57.020 60.125 57.190 61.055 ;
        RECT 57.930 60.845 58.100 61.055 ;
        RECT 58.850 60.885 59.020 61.055 ;
        RECT 57.380 60.515 58.100 60.845 ;
        RECT 56.440 59.955 57.190 60.125 ;
        RECT 57.360 59.745 57.660 60.245 ;
        RECT 57.880 59.945 58.100 60.515 ;
        RECT 58.280 59.745 58.565 60.885 ;
        RECT 58.735 60.740 59.020 60.885 ;
        RECT 59.585 60.755 59.830 61.395 ;
        RECT 60.110 61.310 60.280 61.575 ;
        RECT 60.110 60.980 60.340 61.310 ;
        RECT 58.735 59.925 58.985 60.740 ;
        RECT 59.155 59.745 59.415 60.625 ;
        RECT 60.110 60.585 60.280 60.980 ;
        RECT 59.675 60.415 60.280 60.585 ;
        RECT 60.515 60.695 60.685 62.035 ;
        RECT 61.055 61.765 61.225 62.035 ;
        RECT 61.395 61.935 61.725 62.295 ;
        RECT 62.360 61.845 63.020 62.015 ;
        RECT 61.055 61.615 61.660 61.765 ;
        RECT 61.055 61.595 61.860 61.615 ;
        RECT 60.980 61.055 61.310 61.425 ;
        RECT 61.490 61.285 61.860 61.595 ;
        RECT 62.235 61.345 62.615 61.675 ;
        RECT 61.490 60.885 61.660 61.285 ;
        RECT 60.975 60.715 61.660 60.885 ;
        RECT 59.675 59.915 59.845 60.415 ;
        RECT 60.015 59.745 60.345 60.245 ;
        RECT 60.515 59.915 60.740 60.695 ;
        RECT 60.975 59.965 61.305 60.715 ;
        RECT 61.475 59.745 61.790 60.545 ;
        RECT 61.990 60.375 62.275 61.025 ;
        RECT 62.445 60.965 62.615 61.345 ;
        RECT 62.850 61.385 63.020 61.845 ;
        RECT 63.260 61.555 63.590 62.295 ;
        RECT 63.860 61.555 64.080 61.965 ;
        RECT 64.260 61.555 64.545 62.295 ;
        RECT 64.715 61.695 64.965 61.965 ;
        RECT 65.135 61.830 65.395 62.295 ;
        RECT 64.715 61.555 65.000 61.695 ;
        RECT 63.910 61.385 64.080 61.555 ;
        RECT 64.830 61.385 65.000 61.555 ;
        RECT 62.850 61.215 63.720 61.385 ;
        RECT 63.000 61.055 63.720 61.215 ;
        RECT 63.910 61.055 64.660 61.385 ;
        RECT 64.830 61.055 65.395 61.385 ;
        RECT 62.445 60.385 62.785 60.965 ;
        RECT 63.000 60.125 63.170 61.055 ;
        RECT 63.910 60.845 64.080 61.055 ;
        RECT 64.830 60.885 65.000 61.055 ;
        RECT 63.360 60.515 64.080 60.845 ;
        RECT 62.420 59.955 63.170 60.125 ;
        RECT 63.340 59.745 63.640 60.245 ;
        RECT 63.860 59.945 64.080 60.515 ;
        RECT 64.260 59.745 64.545 60.885 ;
        RECT 64.715 60.740 65.000 60.885 ;
        RECT 64.715 59.925 64.965 60.740 ;
        RECT 65.565 60.640 66.085 62.125 ;
        RECT 66.255 61.635 66.595 62.295 ;
        RECT 65.135 59.745 65.395 60.625 ;
        RECT 65.755 59.745 66.085 60.470 ;
        RECT 66.255 59.915 66.775 61.465 ;
        RECT 66.945 60.640 67.465 62.125 ;
        RECT 67.635 61.635 67.975 62.295 ;
        RECT 68.415 61.745 68.585 62.035 ;
        RECT 68.755 61.915 69.085 62.295 ;
        RECT 68.415 61.575 69.020 61.745 ;
        RECT 67.135 59.745 67.465 60.470 ;
        RECT 67.635 59.915 68.155 61.465 ;
        RECT 68.325 60.755 68.570 61.395 ;
        RECT 68.850 61.310 69.020 61.575 ;
        RECT 68.850 60.980 69.080 61.310 ;
        RECT 68.850 60.585 69.020 60.980 ;
        RECT 68.415 60.415 69.020 60.585 ;
        RECT 69.255 60.695 69.425 62.035 ;
        RECT 69.795 61.765 69.965 62.035 ;
        RECT 70.135 61.935 70.465 62.295 ;
        RECT 71.100 61.845 71.760 62.015 ;
        RECT 69.795 61.615 70.400 61.765 ;
        RECT 69.795 61.595 70.600 61.615 ;
        RECT 69.720 61.055 70.050 61.425 ;
        RECT 70.230 61.285 70.600 61.595 ;
        RECT 70.975 61.345 71.355 61.675 ;
        RECT 70.230 60.885 70.400 61.285 ;
        RECT 69.715 60.715 70.400 60.885 ;
        RECT 68.415 59.915 68.585 60.415 ;
        RECT 68.755 59.745 69.085 60.245 ;
        RECT 69.255 59.915 69.480 60.695 ;
        RECT 69.715 59.965 70.045 60.715 ;
        RECT 70.215 59.745 70.530 60.545 ;
        RECT 70.730 60.375 71.015 61.025 ;
        RECT 71.185 60.965 71.355 61.345 ;
        RECT 71.590 61.385 71.760 61.845 ;
        RECT 72.000 61.555 72.330 62.295 ;
        RECT 72.600 61.555 72.820 61.965 ;
        RECT 73.000 61.555 73.285 62.295 ;
        RECT 73.455 61.695 73.705 61.965 ;
        RECT 73.875 61.830 74.135 62.295 ;
        RECT 73.455 61.555 73.740 61.695 ;
        RECT 74.305 61.570 74.595 62.295 ;
        RECT 74.855 61.745 75.025 62.035 ;
        RECT 75.195 61.915 75.525 62.295 ;
        RECT 74.855 61.575 75.460 61.745 ;
        RECT 72.650 61.385 72.820 61.555 ;
        RECT 73.570 61.385 73.740 61.555 ;
        RECT 71.590 61.215 72.460 61.385 ;
        RECT 71.740 61.055 72.460 61.215 ;
        RECT 72.650 61.055 73.400 61.385 ;
        RECT 73.570 61.055 74.135 61.385 ;
        RECT 71.185 60.385 71.525 60.965 ;
        RECT 71.740 60.125 71.910 61.055 ;
        RECT 72.650 60.845 72.820 61.055 ;
        RECT 73.570 60.885 73.740 61.055 ;
        RECT 72.100 60.515 72.820 60.845 ;
        RECT 71.160 59.955 71.910 60.125 ;
        RECT 72.080 59.745 72.380 60.245 ;
        RECT 72.600 59.945 72.820 60.515 ;
        RECT 73.000 59.745 73.285 60.885 ;
        RECT 73.455 60.740 73.740 60.885 ;
        RECT 73.455 59.925 73.705 60.740 ;
        RECT 73.875 59.745 74.135 60.625 ;
        RECT 74.305 59.745 74.595 60.910 ;
        RECT 74.765 60.755 75.010 61.395 ;
        RECT 75.290 61.310 75.460 61.575 ;
        RECT 75.290 60.980 75.520 61.310 ;
        RECT 75.290 60.585 75.460 60.980 ;
        RECT 74.855 60.415 75.460 60.585 ;
        RECT 75.695 60.695 75.865 62.035 ;
        RECT 76.235 61.765 76.405 62.035 ;
        RECT 76.575 61.935 76.905 62.295 ;
        RECT 77.540 61.845 78.200 62.015 ;
        RECT 76.235 61.615 76.840 61.765 ;
        RECT 76.235 61.595 77.040 61.615 ;
        RECT 76.160 61.055 76.490 61.425 ;
        RECT 76.670 61.285 77.040 61.595 ;
        RECT 77.415 61.345 77.795 61.675 ;
        RECT 76.670 60.885 76.840 61.285 ;
        RECT 76.155 60.715 76.840 60.885 ;
        RECT 74.855 59.915 75.025 60.415 ;
        RECT 75.195 59.745 75.525 60.245 ;
        RECT 75.695 59.915 75.920 60.695 ;
        RECT 76.155 59.965 76.485 60.715 ;
        RECT 76.655 59.745 76.970 60.545 ;
        RECT 77.170 60.375 77.455 61.025 ;
        RECT 77.625 60.965 77.795 61.345 ;
        RECT 78.030 61.385 78.200 61.845 ;
        RECT 78.440 61.555 78.770 62.295 ;
        RECT 79.040 61.555 79.260 61.965 ;
        RECT 79.440 61.555 79.725 62.295 ;
        RECT 79.895 61.695 80.145 61.965 ;
        RECT 80.315 61.830 80.575 62.295 ;
        RECT 80.745 61.830 81.005 62.295 ;
        RECT 81.175 61.695 81.425 61.965 ;
        RECT 79.895 61.555 80.180 61.695 ;
        RECT 79.090 61.385 79.260 61.555 ;
        RECT 80.010 61.385 80.180 61.555 ;
        RECT 81.140 61.555 81.425 61.695 ;
        RECT 81.595 61.555 81.880 62.295 ;
        RECT 82.060 61.555 82.280 61.965 ;
        RECT 82.550 61.555 82.880 62.295 ;
        RECT 83.120 61.845 83.780 62.015 ;
        RECT 84.415 61.935 84.745 62.295 ;
        RECT 81.140 61.385 81.310 61.555 ;
        RECT 82.060 61.385 82.230 61.555 ;
        RECT 83.120 61.385 83.290 61.845 ;
        RECT 84.915 61.765 85.085 62.035 ;
        RECT 78.030 61.215 78.900 61.385 ;
        RECT 78.180 61.055 78.900 61.215 ;
        RECT 79.090 61.055 79.840 61.385 ;
        RECT 80.010 61.055 80.575 61.385 ;
        RECT 80.745 61.055 81.310 61.385 ;
        RECT 81.480 61.055 82.230 61.385 ;
        RECT 82.420 61.215 83.290 61.385 ;
        RECT 83.525 61.345 83.905 61.675 ;
        RECT 84.480 61.615 85.085 61.765 ;
        RECT 84.280 61.595 85.085 61.615 ;
        RECT 82.420 61.055 83.140 61.215 ;
        RECT 77.625 60.385 77.965 60.965 ;
        RECT 78.180 60.125 78.350 61.055 ;
        RECT 79.090 60.845 79.260 61.055 ;
        RECT 80.010 60.885 80.180 61.055 ;
        RECT 78.540 60.515 79.260 60.845 ;
        RECT 77.600 59.955 78.350 60.125 ;
        RECT 78.520 59.745 78.820 60.245 ;
        RECT 79.040 59.945 79.260 60.515 ;
        RECT 79.440 59.745 79.725 60.885 ;
        RECT 79.895 60.740 80.180 60.885 ;
        RECT 81.140 60.885 81.310 61.055 ;
        RECT 81.140 60.740 81.425 60.885 ;
        RECT 79.895 59.925 80.145 60.740 ;
        RECT 80.315 59.745 80.575 60.625 ;
        RECT 80.745 59.745 81.005 60.625 ;
        RECT 81.175 59.925 81.425 60.740 ;
        RECT 81.595 59.745 81.880 60.885 ;
        RECT 82.060 60.845 82.230 61.055 ;
        RECT 82.060 60.515 82.780 60.845 ;
        RECT 82.060 59.945 82.280 60.515 ;
        RECT 82.500 59.745 82.800 60.245 ;
        RECT 82.970 60.125 83.140 61.055 ;
        RECT 83.525 60.965 83.695 61.345 ;
        RECT 84.280 61.285 84.650 61.595 ;
        RECT 83.355 60.385 83.695 60.965 ;
        RECT 83.865 60.375 84.150 61.025 ;
        RECT 84.480 60.885 84.650 61.285 ;
        RECT 84.830 61.055 85.160 61.425 ;
        RECT 84.480 60.715 85.165 60.885 ;
        RECT 82.970 59.955 83.720 60.125 ;
        RECT 84.350 59.745 84.665 60.545 ;
        RECT 84.835 59.965 85.165 60.715 ;
        RECT 85.455 60.695 85.625 62.035 ;
        RECT 85.795 61.915 86.125 62.295 ;
        RECT 86.295 61.745 86.465 62.035 ;
        RECT 85.860 61.575 86.465 61.745 ;
        RECT 86.815 61.745 86.985 62.035 ;
        RECT 87.155 61.915 87.485 62.295 ;
        RECT 86.815 61.575 87.420 61.745 ;
        RECT 85.860 61.310 86.030 61.575 ;
        RECT 85.800 60.980 86.030 61.310 ;
        RECT 85.400 59.915 85.625 60.695 ;
        RECT 85.860 60.585 86.030 60.980 ;
        RECT 86.310 60.755 86.555 61.395 ;
        RECT 86.725 60.755 86.970 61.395 ;
        RECT 87.250 61.310 87.420 61.575 ;
        RECT 87.250 60.980 87.480 61.310 ;
        RECT 87.250 60.585 87.420 60.980 ;
        RECT 85.860 60.415 86.465 60.585 ;
        RECT 85.795 59.745 86.125 60.245 ;
        RECT 86.295 59.915 86.465 60.415 ;
        RECT 86.815 60.415 87.420 60.585 ;
        RECT 87.655 60.695 87.825 62.035 ;
        RECT 88.195 61.765 88.365 62.035 ;
        RECT 88.535 61.935 88.865 62.295 ;
        RECT 89.500 61.845 90.160 62.015 ;
        RECT 88.195 61.615 88.800 61.765 ;
        RECT 88.195 61.595 89.000 61.615 ;
        RECT 88.120 61.055 88.450 61.425 ;
        RECT 88.630 61.285 89.000 61.595 ;
        RECT 89.375 61.345 89.755 61.675 ;
        RECT 88.630 60.885 88.800 61.285 ;
        RECT 88.115 60.715 88.800 60.885 ;
        RECT 86.815 59.915 86.985 60.415 ;
        RECT 87.155 59.745 87.485 60.245 ;
        RECT 87.655 59.915 87.880 60.695 ;
        RECT 88.115 59.965 88.445 60.715 ;
        RECT 88.615 59.745 88.930 60.545 ;
        RECT 89.130 60.375 89.415 61.025 ;
        RECT 89.585 60.965 89.755 61.345 ;
        RECT 89.990 61.385 90.160 61.845 ;
        RECT 90.400 61.555 90.730 62.295 ;
        RECT 91.000 61.555 91.220 61.965 ;
        RECT 91.400 61.555 91.685 62.295 ;
        RECT 91.855 61.695 92.105 61.965 ;
        RECT 92.275 61.830 92.535 62.295 ;
        RECT 92.795 61.745 92.965 62.035 ;
        RECT 93.135 61.915 93.465 62.295 ;
        RECT 91.855 61.555 92.140 61.695 ;
        RECT 92.795 61.575 93.400 61.745 ;
        RECT 91.050 61.385 91.220 61.555 ;
        RECT 91.970 61.385 92.140 61.555 ;
        RECT 89.990 61.215 90.860 61.385 ;
        RECT 90.140 61.055 90.860 61.215 ;
        RECT 91.050 61.055 91.800 61.385 ;
        RECT 91.970 61.055 92.535 61.385 ;
        RECT 89.585 60.385 89.925 60.965 ;
        RECT 90.140 60.125 90.310 61.055 ;
        RECT 91.050 60.845 91.220 61.055 ;
        RECT 91.970 60.885 92.140 61.055 ;
        RECT 90.500 60.515 91.220 60.845 ;
        RECT 89.560 59.955 90.310 60.125 ;
        RECT 90.480 59.745 90.780 60.245 ;
        RECT 91.000 59.945 91.220 60.515 ;
        RECT 91.400 59.745 91.685 60.885 ;
        RECT 91.855 60.740 92.140 60.885 ;
        RECT 92.705 60.755 92.950 61.395 ;
        RECT 93.230 61.310 93.400 61.575 ;
        RECT 93.230 60.980 93.460 61.310 ;
        RECT 91.855 59.925 92.105 60.740 ;
        RECT 92.275 59.745 92.535 60.625 ;
        RECT 93.230 60.585 93.400 60.980 ;
        RECT 92.795 60.415 93.400 60.585 ;
        RECT 93.635 60.695 93.805 62.035 ;
        RECT 94.175 61.765 94.345 62.035 ;
        RECT 94.515 61.935 94.845 62.295 ;
        RECT 95.480 61.845 96.140 62.015 ;
        RECT 94.175 61.615 94.780 61.765 ;
        RECT 94.175 61.595 94.980 61.615 ;
        RECT 94.100 61.055 94.430 61.425 ;
        RECT 94.610 61.285 94.980 61.595 ;
        RECT 95.355 61.345 95.735 61.675 ;
        RECT 94.610 60.885 94.780 61.285 ;
        RECT 94.095 60.715 94.780 60.885 ;
        RECT 92.795 59.915 92.965 60.415 ;
        RECT 93.135 59.745 93.465 60.245 ;
        RECT 93.635 59.915 93.860 60.695 ;
        RECT 94.095 59.965 94.425 60.715 ;
        RECT 94.595 59.745 94.910 60.545 ;
        RECT 95.110 60.375 95.395 61.025 ;
        RECT 95.565 60.965 95.735 61.345 ;
        RECT 95.970 61.385 96.140 61.845 ;
        RECT 96.380 61.555 96.710 62.295 ;
        RECT 96.980 61.555 97.200 61.965 ;
        RECT 97.380 61.555 97.665 62.295 ;
        RECT 97.835 61.695 98.085 61.965 ;
        RECT 98.255 61.830 98.515 62.295 ;
        RECT 97.835 61.555 98.120 61.695 ;
        RECT 97.030 61.385 97.200 61.555 ;
        RECT 97.950 61.385 98.120 61.555 ;
        RECT 95.970 61.215 96.840 61.385 ;
        RECT 96.120 61.055 96.840 61.215 ;
        RECT 97.030 61.055 97.780 61.385 ;
        RECT 97.950 61.055 98.515 61.385 ;
        RECT 95.565 60.385 95.905 60.965 ;
        RECT 96.120 60.125 96.290 61.055 ;
        RECT 97.030 60.845 97.200 61.055 ;
        RECT 97.950 60.885 98.120 61.055 ;
        RECT 96.480 60.515 97.200 60.845 ;
        RECT 95.540 59.955 96.290 60.125 ;
        RECT 96.460 59.745 96.760 60.245 ;
        RECT 96.980 59.945 97.200 60.515 ;
        RECT 97.380 59.745 97.665 60.885 ;
        RECT 97.835 60.740 98.120 60.885 ;
        RECT 97.835 59.925 98.085 60.740 ;
        RECT 98.685 60.640 99.205 62.125 ;
        RECT 99.375 61.635 99.715 62.295 ;
        RECT 100.065 61.570 100.355 62.295 ;
        RECT 100.615 61.745 100.785 62.035 ;
        RECT 100.955 61.915 101.285 62.295 ;
        RECT 100.615 61.575 101.220 61.745 ;
        RECT 98.255 59.745 98.515 60.625 ;
        RECT 98.875 59.745 99.205 60.470 ;
        RECT 99.375 59.915 99.895 61.465 ;
        RECT 100.065 59.745 100.355 60.910 ;
        RECT 100.525 60.755 100.770 61.395 ;
        RECT 101.050 61.310 101.220 61.575 ;
        RECT 101.050 60.980 101.280 61.310 ;
        RECT 101.050 60.585 101.220 60.980 ;
        RECT 100.615 60.415 101.220 60.585 ;
        RECT 101.455 60.695 101.625 62.035 ;
        RECT 101.995 61.765 102.165 62.035 ;
        RECT 102.335 61.935 102.665 62.295 ;
        RECT 103.300 61.845 103.960 62.015 ;
        RECT 101.995 61.615 102.600 61.765 ;
        RECT 101.995 61.595 102.800 61.615 ;
        RECT 101.920 61.055 102.250 61.425 ;
        RECT 102.430 61.285 102.800 61.595 ;
        RECT 103.175 61.345 103.555 61.675 ;
        RECT 102.430 60.885 102.600 61.285 ;
        RECT 101.915 60.715 102.600 60.885 ;
        RECT 100.615 59.915 100.785 60.415 ;
        RECT 100.955 59.745 101.285 60.245 ;
        RECT 101.455 59.915 101.680 60.695 ;
        RECT 101.915 59.965 102.245 60.715 ;
        RECT 102.415 59.745 102.730 60.545 ;
        RECT 102.930 60.375 103.215 61.025 ;
        RECT 103.385 60.965 103.555 61.345 ;
        RECT 103.790 61.385 103.960 61.845 ;
        RECT 104.200 61.555 104.530 62.295 ;
        RECT 104.800 61.555 105.020 61.965 ;
        RECT 105.200 61.555 105.485 62.295 ;
        RECT 105.655 61.695 105.905 61.965 ;
        RECT 106.075 61.830 106.335 62.295 ;
        RECT 106.595 61.745 106.765 62.035 ;
        RECT 106.935 61.915 107.265 62.295 ;
        RECT 105.655 61.555 105.940 61.695 ;
        RECT 106.595 61.575 107.200 61.745 ;
        RECT 104.850 61.385 105.020 61.555 ;
        RECT 105.770 61.385 105.940 61.555 ;
        RECT 103.790 61.215 104.660 61.385 ;
        RECT 103.940 61.055 104.660 61.215 ;
        RECT 104.850 61.055 105.600 61.385 ;
        RECT 105.770 61.055 106.335 61.385 ;
        RECT 103.385 60.385 103.725 60.965 ;
        RECT 103.940 60.125 104.110 61.055 ;
        RECT 104.850 60.845 105.020 61.055 ;
        RECT 105.770 60.885 105.940 61.055 ;
        RECT 104.300 60.515 105.020 60.845 ;
        RECT 103.360 59.955 104.110 60.125 ;
        RECT 104.280 59.745 104.580 60.245 ;
        RECT 104.800 59.945 105.020 60.515 ;
        RECT 105.200 59.745 105.485 60.885 ;
        RECT 105.655 60.740 105.940 60.885 ;
        RECT 106.505 60.755 106.750 61.395 ;
        RECT 107.030 61.310 107.200 61.575 ;
        RECT 107.030 60.980 107.260 61.310 ;
        RECT 105.655 59.925 105.905 60.740 ;
        RECT 106.075 59.745 106.335 60.625 ;
        RECT 107.030 60.585 107.200 60.980 ;
        RECT 106.595 60.415 107.200 60.585 ;
        RECT 107.435 60.695 107.605 62.035 ;
        RECT 107.975 61.765 108.145 62.035 ;
        RECT 108.315 61.935 108.645 62.295 ;
        RECT 109.280 61.845 109.940 62.015 ;
        RECT 107.975 61.615 108.580 61.765 ;
        RECT 107.975 61.595 108.780 61.615 ;
        RECT 107.900 61.055 108.230 61.425 ;
        RECT 108.410 61.285 108.780 61.595 ;
        RECT 109.155 61.345 109.535 61.675 ;
        RECT 108.410 60.885 108.580 61.285 ;
        RECT 107.895 60.715 108.580 60.885 ;
        RECT 106.595 59.915 106.765 60.415 ;
        RECT 106.935 59.745 107.265 60.245 ;
        RECT 107.435 59.915 107.660 60.695 ;
        RECT 107.895 59.965 108.225 60.715 ;
        RECT 108.395 59.745 108.710 60.545 ;
        RECT 108.910 60.375 109.195 61.025 ;
        RECT 109.365 60.965 109.535 61.345 ;
        RECT 109.770 61.385 109.940 61.845 ;
        RECT 110.180 61.555 110.510 62.295 ;
        RECT 110.780 61.555 111.000 61.965 ;
        RECT 111.180 61.555 111.465 62.295 ;
        RECT 111.635 61.695 111.885 61.965 ;
        RECT 112.055 61.830 112.315 62.295 ;
        RECT 112.575 61.745 112.745 62.035 ;
        RECT 112.915 61.915 113.245 62.295 ;
        RECT 111.635 61.555 111.920 61.695 ;
        RECT 112.575 61.575 113.180 61.745 ;
        RECT 110.830 61.385 111.000 61.555 ;
        RECT 111.750 61.385 111.920 61.555 ;
        RECT 109.770 61.215 110.640 61.385 ;
        RECT 109.920 61.055 110.640 61.215 ;
        RECT 110.830 61.055 111.580 61.385 ;
        RECT 111.750 61.055 112.315 61.385 ;
        RECT 109.365 60.385 109.705 60.965 ;
        RECT 109.920 60.125 110.090 61.055 ;
        RECT 110.830 60.845 111.000 61.055 ;
        RECT 111.750 60.885 111.920 61.055 ;
        RECT 110.280 60.515 111.000 60.845 ;
        RECT 109.340 59.955 110.090 60.125 ;
        RECT 110.260 59.745 110.560 60.245 ;
        RECT 110.780 59.945 111.000 60.515 ;
        RECT 111.180 59.745 111.465 60.885 ;
        RECT 111.635 60.740 111.920 60.885 ;
        RECT 112.485 60.755 112.730 61.395 ;
        RECT 113.010 61.310 113.180 61.575 ;
        RECT 113.010 60.980 113.240 61.310 ;
        RECT 111.635 59.925 111.885 60.740 ;
        RECT 112.055 59.745 112.315 60.625 ;
        RECT 113.010 60.585 113.180 60.980 ;
        RECT 112.575 60.415 113.180 60.585 ;
        RECT 113.415 60.695 113.585 62.035 ;
        RECT 113.955 61.765 114.125 62.035 ;
        RECT 114.295 61.935 114.625 62.295 ;
        RECT 115.260 61.845 115.920 62.015 ;
        RECT 113.955 61.615 114.560 61.765 ;
        RECT 113.955 61.595 114.760 61.615 ;
        RECT 113.880 61.055 114.210 61.425 ;
        RECT 114.390 61.285 114.760 61.595 ;
        RECT 115.135 61.345 115.515 61.675 ;
        RECT 114.390 60.885 114.560 61.285 ;
        RECT 113.875 60.715 114.560 60.885 ;
        RECT 112.575 59.915 112.745 60.415 ;
        RECT 112.915 59.745 113.245 60.245 ;
        RECT 113.415 59.915 113.640 60.695 ;
        RECT 113.875 59.965 114.205 60.715 ;
        RECT 114.375 59.745 114.690 60.545 ;
        RECT 114.890 60.375 115.175 61.025 ;
        RECT 115.345 60.965 115.515 61.345 ;
        RECT 115.750 61.385 115.920 61.845 ;
        RECT 116.160 61.555 116.490 62.295 ;
        RECT 116.760 61.555 116.980 61.965 ;
        RECT 117.160 61.555 117.445 62.295 ;
        RECT 117.615 61.695 117.865 61.965 ;
        RECT 118.035 61.830 118.295 62.295 ;
        RECT 118.555 61.745 118.725 62.035 ;
        RECT 118.895 61.915 119.225 62.295 ;
        RECT 117.615 61.555 117.900 61.695 ;
        RECT 118.555 61.575 119.160 61.745 ;
        RECT 116.810 61.385 116.980 61.555 ;
        RECT 117.730 61.385 117.900 61.555 ;
        RECT 115.750 61.215 116.620 61.385 ;
        RECT 115.900 61.055 116.620 61.215 ;
        RECT 116.810 61.055 117.560 61.385 ;
        RECT 117.730 61.055 118.295 61.385 ;
        RECT 115.345 60.385 115.685 60.965 ;
        RECT 115.900 60.125 116.070 61.055 ;
        RECT 116.810 60.845 116.980 61.055 ;
        RECT 117.730 60.885 117.900 61.055 ;
        RECT 116.260 60.515 116.980 60.845 ;
        RECT 115.320 59.955 116.070 60.125 ;
        RECT 116.240 59.745 116.540 60.245 ;
        RECT 116.760 59.945 116.980 60.515 ;
        RECT 117.160 59.745 117.445 60.885 ;
        RECT 117.615 60.740 117.900 60.885 ;
        RECT 118.465 60.755 118.710 61.395 ;
        RECT 118.990 61.310 119.160 61.575 ;
        RECT 118.990 60.980 119.220 61.310 ;
        RECT 117.615 59.925 117.865 60.740 ;
        RECT 118.035 59.745 118.295 60.625 ;
        RECT 118.990 60.585 119.160 60.980 ;
        RECT 118.555 60.415 119.160 60.585 ;
        RECT 119.395 60.695 119.565 62.035 ;
        RECT 119.935 61.765 120.105 62.035 ;
        RECT 120.275 61.935 120.605 62.295 ;
        RECT 121.240 61.845 121.900 62.015 ;
        RECT 119.935 61.615 120.540 61.765 ;
        RECT 119.935 61.595 120.740 61.615 ;
        RECT 119.860 61.055 120.190 61.425 ;
        RECT 120.370 61.285 120.740 61.595 ;
        RECT 121.115 61.345 121.495 61.675 ;
        RECT 120.370 60.885 120.540 61.285 ;
        RECT 119.855 60.715 120.540 60.885 ;
        RECT 118.555 59.915 118.725 60.415 ;
        RECT 118.895 59.745 119.225 60.245 ;
        RECT 119.395 59.915 119.620 60.695 ;
        RECT 119.855 59.965 120.185 60.715 ;
        RECT 120.355 59.745 120.670 60.545 ;
        RECT 120.870 60.375 121.155 61.025 ;
        RECT 121.325 60.965 121.495 61.345 ;
        RECT 121.730 61.385 121.900 61.845 ;
        RECT 122.140 61.555 122.470 62.295 ;
        RECT 122.740 61.555 122.960 61.965 ;
        RECT 123.140 61.555 123.425 62.295 ;
        RECT 123.595 61.695 123.845 61.965 ;
        RECT 124.015 61.830 124.275 62.295 ;
        RECT 123.595 61.555 123.880 61.695 ;
        RECT 124.625 61.635 124.965 62.295 ;
        RECT 122.790 61.385 122.960 61.555 ;
        RECT 123.710 61.385 123.880 61.555 ;
        RECT 121.730 61.215 122.600 61.385 ;
        RECT 121.880 61.055 122.600 61.215 ;
        RECT 122.790 61.055 123.540 61.385 ;
        RECT 123.710 61.055 124.275 61.385 ;
        RECT 121.325 60.385 121.665 60.965 ;
        RECT 121.880 60.125 122.050 61.055 ;
        RECT 122.790 60.845 122.960 61.055 ;
        RECT 123.710 60.885 123.880 61.055 ;
        RECT 122.240 60.515 122.960 60.845 ;
        RECT 121.300 59.955 122.050 60.125 ;
        RECT 122.220 59.745 122.520 60.245 ;
        RECT 122.740 59.945 122.960 60.515 ;
        RECT 123.140 59.745 123.425 60.885 ;
        RECT 123.595 60.740 123.880 60.885 ;
        RECT 123.595 59.925 123.845 60.740 ;
        RECT 124.015 59.745 124.275 60.625 ;
        RECT 124.445 59.915 124.965 61.465 ;
        RECT 125.135 60.640 125.655 62.125 ;
        RECT 125.825 61.570 126.115 62.295 ;
        RECT 126.375 61.745 126.545 62.035 ;
        RECT 126.715 61.915 127.045 62.295 ;
        RECT 126.375 61.575 126.980 61.745 ;
        RECT 125.135 59.745 125.465 60.470 ;
        RECT 125.825 59.745 126.115 60.910 ;
        RECT 126.285 60.755 126.530 61.395 ;
        RECT 126.810 61.310 126.980 61.575 ;
        RECT 126.810 60.980 127.040 61.310 ;
        RECT 126.810 60.585 126.980 60.980 ;
        RECT 126.375 60.415 126.980 60.585 ;
        RECT 127.215 60.695 127.385 62.035 ;
        RECT 127.755 61.765 127.925 62.035 ;
        RECT 128.095 61.935 128.425 62.295 ;
        RECT 129.060 61.845 129.720 62.015 ;
        RECT 127.755 61.615 128.360 61.765 ;
        RECT 127.755 61.595 128.560 61.615 ;
        RECT 127.680 61.055 128.010 61.425 ;
        RECT 128.190 61.285 128.560 61.595 ;
        RECT 128.935 61.345 129.315 61.675 ;
        RECT 128.190 60.885 128.360 61.285 ;
        RECT 127.675 60.715 128.360 60.885 ;
        RECT 126.375 59.915 126.545 60.415 ;
        RECT 126.715 59.745 127.045 60.245 ;
        RECT 127.215 59.915 127.440 60.695 ;
        RECT 127.675 59.965 128.005 60.715 ;
        RECT 128.175 59.745 128.490 60.545 ;
        RECT 128.690 60.375 128.975 61.025 ;
        RECT 129.145 60.965 129.315 61.345 ;
        RECT 129.550 61.385 129.720 61.845 ;
        RECT 129.960 61.555 130.290 62.295 ;
        RECT 130.560 61.555 130.780 61.965 ;
        RECT 130.960 61.555 131.245 62.295 ;
        RECT 131.415 61.695 131.665 61.965 ;
        RECT 131.835 61.830 132.095 62.295 ;
        RECT 132.355 61.745 132.525 62.035 ;
        RECT 132.695 61.915 133.025 62.295 ;
        RECT 131.415 61.555 131.700 61.695 ;
        RECT 132.355 61.575 132.960 61.745 ;
        RECT 130.610 61.385 130.780 61.555 ;
        RECT 131.530 61.385 131.700 61.555 ;
        RECT 129.550 61.215 130.420 61.385 ;
        RECT 129.700 61.055 130.420 61.215 ;
        RECT 130.610 61.055 131.360 61.385 ;
        RECT 131.530 61.055 132.095 61.385 ;
        RECT 129.145 60.385 129.485 60.965 ;
        RECT 129.700 60.125 129.870 61.055 ;
        RECT 130.610 60.845 130.780 61.055 ;
        RECT 131.530 60.885 131.700 61.055 ;
        RECT 130.060 60.515 130.780 60.845 ;
        RECT 129.120 59.955 129.870 60.125 ;
        RECT 130.040 59.745 130.340 60.245 ;
        RECT 130.560 59.945 130.780 60.515 ;
        RECT 130.960 59.745 131.245 60.885 ;
        RECT 131.415 60.740 131.700 60.885 ;
        RECT 132.265 60.755 132.510 61.395 ;
        RECT 132.790 61.310 132.960 61.575 ;
        RECT 132.790 60.980 133.020 61.310 ;
        RECT 131.415 59.925 131.665 60.740 ;
        RECT 131.835 59.745 132.095 60.625 ;
        RECT 132.790 60.585 132.960 60.980 ;
        RECT 132.355 60.415 132.960 60.585 ;
        RECT 133.195 60.695 133.365 62.035 ;
        RECT 133.735 61.765 133.905 62.035 ;
        RECT 134.075 61.935 134.405 62.295 ;
        RECT 135.040 61.845 135.700 62.015 ;
        RECT 133.735 61.615 134.340 61.765 ;
        RECT 133.735 61.595 134.540 61.615 ;
        RECT 133.660 61.055 133.990 61.425 ;
        RECT 134.170 61.285 134.540 61.595 ;
        RECT 134.915 61.345 135.295 61.675 ;
        RECT 134.170 60.885 134.340 61.285 ;
        RECT 133.655 60.715 134.340 60.885 ;
        RECT 132.355 59.915 132.525 60.415 ;
        RECT 132.695 59.745 133.025 60.245 ;
        RECT 133.195 59.915 133.420 60.695 ;
        RECT 133.655 59.965 133.985 60.715 ;
        RECT 134.155 59.745 134.470 60.545 ;
        RECT 134.670 60.375 134.955 61.025 ;
        RECT 135.125 60.965 135.295 61.345 ;
        RECT 135.530 61.385 135.700 61.845 ;
        RECT 135.940 61.555 136.270 62.295 ;
        RECT 136.540 61.555 136.760 61.965 ;
        RECT 136.940 61.555 137.225 62.295 ;
        RECT 137.395 61.695 137.645 61.965 ;
        RECT 137.815 61.830 138.075 62.295 ;
        RECT 138.335 61.745 138.505 62.035 ;
        RECT 138.675 61.915 139.005 62.295 ;
        RECT 137.395 61.555 137.680 61.695 ;
        RECT 138.335 61.575 138.940 61.745 ;
        RECT 136.590 61.385 136.760 61.555 ;
        RECT 137.510 61.385 137.680 61.555 ;
        RECT 135.530 61.215 136.400 61.385 ;
        RECT 135.680 61.055 136.400 61.215 ;
        RECT 136.590 61.055 137.340 61.385 ;
        RECT 137.510 61.055 138.075 61.385 ;
        RECT 135.125 60.385 135.465 60.965 ;
        RECT 135.680 60.125 135.850 61.055 ;
        RECT 136.590 60.845 136.760 61.055 ;
        RECT 137.510 60.885 137.680 61.055 ;
        RECT 136.040 60.515 136.760 60.845 ;
        RECT 135.100 59.955 135.850 60.125 ;
        RECT 136.020 59.745 136.320 60.245 ;
        RECT 136.540 59.945 136.760 60.515 ;
        RECT 136.940 59.745 137.225 60.885 ;
        RECT 137.395 60.740 137.680 60.885 ;
        RECT 138.245 60.755 138.490 61.395 ;
        RECT 138.770 61.310 138.940 61.575 ;
        RECT 138.770 60.980 139.000 61.310 ;
        RECT 137.395 59.925 137.645 60.740 ;
        RECT 137.815 59.745 138.075 60.625 ;
        RECT 138.770 60.585 138.940 60.980 ;
        RECT 138.335 60.415 138.940 60.585 ;
        RECT 139.175 60.695 139.345 62.035 ;
        RECT 139.715 61.765 139.885 62.035 ;
        RECT 140.055 61.935 140.385 62.295 ;
        RECT 141.020 61.845 141.680 62.015 ;
        RECT 139.715 61.615 140.320 61.765 ;
        RECT 139.715 61.595 140.520 61.615 ;
        RECT 139.640 61.055 139.970 61.425 ;
        RECT 140.150 61.285 140.520 61.595 ;
        RECT 140.895 61.345 141.275 61.675 ;
        RECT 140.150 60.885 140.320 61.285 ;
        RECT 139.635 60.715 140.320 60.885 ;
        RECT 138.335 59.915 138.505 60.415 ;
        RECT 138.675 59.745 139.005 60.245 ;
        RECT 139.175 59.915 139.400 60.695 ;
        RECT 139.635 59.965 139.965 60.715 ;
        RECT 140.135 59.745 140.450 60.545 ;
        RECT 140.650 60.375 140.935 61.025 ;
        RECT 141.105 60.965 141.275 61.345 ;
        RECT 141.510 61.385 141.680 61.845 ;
        RECT 141.920 61.555 142.250 62.295 ;
        RECT 142.520 61.555 142.740 61.965 ;
        RECT 142.920 61.555 143.205 62.295 ;
        RECT 143.375 61.695 143.625 61.965 ;
        RECT 143.795 61.830 144.055 62.295 ;
        RECT 144.315 61.745 144.485 62.035 ;
        RECT 144.655 61.915 144.985 62.295 ;
        RECT 143.375 61.555 143.660 61.695 ;
        RECT 144.315 61.575 144.920 61.745 ;
        RECT 142.570 61.385 142.740 61.555 ;
        RECT 143.490 61.385 143.660 61.555 ;
        RECT 141.510 61.215 142.380 61.385 ;
        RECT 141.660 61.055 142.380 61.215 ;
        RECT 142.570 61.055 143.320 61.385 ;
        RECT 143.490 61.055 144.055 61.385 ;
        RECT 141.105 60.385 141.445 60.965 ;
        RECT 141.660 60.125 141.830 61.055 ;
        RECT 142.570 60.845 142.740 61.055 ;
        RECT 143.490 60.885 143.660 61.055 ;
        RECT 142.020 60.515 142.740 60.845 ;
        RECT 141.080 59.955 141.830 60.125 ;
        RECT 142.000 59.745 142.300 60.245 ;
        RECT 142.520 59.945 142.740 60.515 ;
        RECT 142.920 59.745 143.205 60.885 ;
        RECT 143.375 60.740 143.660 60.885 ;
        RECT 144.225 60.755 144.470 61.395 ;
        RECT 144.750 61.310 144.920 61.575 ;
        RECT 144.750 60.980 144.980 61.310 ;
        RECT 143.375 59.925 143.625 60.740 ;
        RECT 143.795 59.745 144.055 60.625 ;
        RECT 144.750 60.585 144.920 60.980 ;
        RECT 144.315 60.415 144.920 60.585 ;
        RECT 145.155 60.695 145.325 62.035 ;
        RECT 145.695 61.765 145.865 62.035 ;
        RECT 146.035 61.935 146.365 62.295 ;
        RECT 147.000 61.845 147.660 62.015 ;
        RECT 145.695 61.615 146.300 61.765 ;
        RECT 145.695 61.595 146.500 61.615 ;
        RECT 145.620 61.055 145.950 61.425 ;
        RECT 146.130 61.285 146.500 61.595 ;
        RECT 146.875 61.345 147.255 61.675 ;
        RECT 146.130 60.885 146.300 61.285 ;
        RECT 145.615 60.715 146.300 60.885 ;
        RECT 144.315 59.915 144.485 60.415 ;
        RECT 144.655 59.745 144.985 60.245 ;
        RECT 145.155 59.915 145.380 60.695 ;
        RECT 145.615 59.965 145.945 60.715 ;
        RECT 146.115 59.745 146.430 60.545 ;
        RECT 146.630 60.375 146.915 61.025 ;
        RECT 147.085 60.965 147.255 61.345 ;
        RECT 147.490 61.385 147.660 61.845 ;
        RECT 147.900 61.555 148.230 62.295 ;
        RECT 148.500 61.555 148.720 61.965 ;
        RECT 148.900 61.555 149.185 62.295 ;
        RECT 149.355 61.695 149.605 61.965 ;
        RECT 149.775 61.830 150.035 62.295 ;
        RECT 149.355 61.555 149.640 61.695 ;
        RECT 148.550 61.385 148.720 61.555 ;
        RECT 149.470 61.385 149.640 61.555 ;
        RECT 150.205 61.545 151.415 62.295 ;
        RECT 151.585 61.570 151.875 62.295 ;
        RECT 147.490 61.215 148.360 61.385 ;
        RECT 147.640 61.055 148.360 61.215 ;
        RECT 148.550 61.055 149.300 61.385 ;
        RECT 149.470 61.055 150.035 61.385 ;
        RECT 147.085 60.385 147.425 60.965 ;
        RECT 147.640 60.125 147.810 61.055 ;
        RECT 148.550 60.845 148.720 61.055 ;
        RECT 149.470 60.885 149.640 61.055 ;
        RECT 150.205 61.005 150.725 61.545 ;
        RECT 152.045 61.525 155.555 62.295 ;
        RECT 155.725 61.545 156.935 62.295 ;
        RECT 148.000 60.515 148.720 60.845 ;
        RECT 147.060 59.955 147.810 60.125 ;
        RECT 147.980 59.745 148.280 60.245 ;
        RECT 148.500 59.945 148.720 60.515 ;
        RECT 148.900 59.745 149.185 60.885 ;
        RECT 149.355 60.740 149.640 60.885 ;
        RECT 150.895 60.835 151.415 61.375 ;
        RECT 152.045 61.005 153.695 61.525 ;
        RECT 149.355 59.925 149.605 60.740 ;
        RECT 149.775 59.745 150.035 60.625 ;
        RECT 150.205 59.745 151.415 60.835 ;
        RECT 151.585 59.745 151.875 60.910 ;
        RECT 153.865 60.835 155.555 61.355 ;
        RECT 152.045 59.745 155.555 60.835 ;
        RECT 155.725 60.835 156.245 61.375 ;
        RECT 156.415 61.005 156.935 61.545 ;
        RECT 155.725 59.745 156.935 60.835 ;
        RECT 22.700 59.575 157.020 59.745 ;
        RECT 22.785 58.485 23.995 59.575 ;
        RECT 22.785 57.775 23.305 58.315 ;
        RECT 23.475 57.945 23.995 58.485 ;
        RECT 25.085 57.855 25.605 59.405 ;
        RECT 25.775 58.850 26.105 59.575 ;
        RECT 22.785 57.025 23.995 57.775 ;
        RECT 25.265 57.025 25.605 57.685 ;
        RECT 25.775 57.195 26.295 58.680 ;
        RECT 26.925 57.855 27.445 59.405 ;
        RECT 27.615 58.850 27.945 59.575 ;
        RECT 27.105 57.025 27.445 57.685 ;
        RECT 27.615 57.195 28.135 58.680 ;
        RECT 28.305 58.485 29.515 59.575 ;
        RECT 29.775 58.905 29.945 59.405 ;
        RECT 30.115 59.075 30.445 59.575 ;
        RECT 29.775 58.735 30.380 58.905 ;
        RECT 28.305 57.775 28.825 58.315 ;
        RECT 28.995 57.945 29.515 58.485 ;
        RECT 29.685 57.925 29.930 58.565 ;
        RECT 30.210 58.340 30.380 58.735 ;
        RECT 30.615 58.625 30.840 59.405 ;
        RECT 30.210 58.010 30.440 58.340 ;
        RECT 28.305 57.025 29.515 57.775 ;
        RECT 30.210 57.745 30.380 58.010 ;
        RECT 29.775 57.575 30.380 57.745 ;
        RECT 29.775 57.285 29.945 57.575 ;
        RECT 30.115 57.025 30.445 57.405 ;
        RECT 30.615 57.285 30.785 58.625 ;
        RECT 31.075 58.605 31.405 59.355 ;
        RECT 31.575 58.775 31.890 59.575 ;
        RECT 32.520 59.195 33.270 59.365 ;
        RECT 31.075 58.435 31.760 58.605 ;
        RECT 31.080 57.895 31.410 58.265 ;
        RECT 31.590 58.035 31.760 58.435 ;
        RECT 32.090 58.295 32.375 58.945 ;
        RECT 32.545 58.355 32.885 58.935 ;
        RECT 31.590 57.725 31.960 58.035 ;
        RECT 32.545 57.975 32.715 58.355 ;
        RECT 33.100 58.265 33.270 59.195 ;
        RECT 33.440 59.075 33.740 59.575 ;
        RECT 33.960 58.805 34.180 59.375 ;
        RECT 33.460 58.475 34.180 58.805 ;
        RECT 34.010 58.265 34.180 58.475 ;
        RECT 34.360 58.435 34.645 59.575 ;
        RECT 34.815 58.580 35.065 59.395 ;
        RECT 35.235 58.695 35.495 59.575 ;
        RECT 34.815 58.435 35.100 58.580 ;
        RECT 34.930 58.265 35.100 58.435 ;
        RECT 35.665 58.410 35.955 59.575 ;
        RECT 33.100 58.105 33.820 58.265 ;
        RECT 31.155 57.705 31.960 57.725 ;
        RECT 31.155 57.555 31.760 57.705 ;
        RECT 32.335 57.645 32.715 57.975 ;
        RECT 32.950 57.935 33.820 58.105 ;
        RECT 34.010 57.935 34.760 58.265 ;
        RECT 34.930 57.935 35.495 58.265 ;
        RECT 31.155 57.285 31.325 57.555 ;
        RECT 32.950 57.475 33.120 57.935 ;
        RECT 34.010 57.765 34.180 57.935 ;
        RECT 34.930 57.765 35.100 57.935 ;
        RECT 37.045 57.855 37.565 59.405 ;
        RECT 37.735 58.850 38.065 59.575 ;
        RECT 31.495 57.025 31.825 57.385 ;
        RECT 32.460 57.305 33.120 57.475 ;
        RECT 33.360 57.025 33.690 57.765 ;
        RECT 33.960 57.355 34.180 57.765 ;
        RECT 34.360 57.025 34.645 57.765 ;
        RECT 34.815 57.625 35.100 57.765 ;
        RECT 34.815 57.355 35.065 57.625 ;
        RECT 35.235 57.025 35.495 57.490 ;
        RECT 35.665 57.025 35.955 57.750 ;
        RECT 37.225 57.025 37.565 57.685 ;
        RECT 37.735 57.195 38.255 58.680 ;
        RECT 38.425 57.855 38.945 59.405 ;
        RECT 39.115 58.850 39.445 59.575 ;
        RECT 38.605 57.025 38.945 57.685 ;
        RECT 39.115 57.195 39.635 58.680 ;
        RECT 39.805 58.485 41.015 59.575 ;
        RECT 41.275 58.905 41.445 59.405 ;
        RECT 41.615 59.075 41.945 59.575 ;
        RECT 41.275 58.735 41.880 58.905 ;
        RECT 39.805 57.775 40.325 58.315 ;
        RECT 40.495 57.945 41.015 58.485 ;
        RECT 41.185 57.925 41.430 58.565 ;
        RECT 41.710 58.340 41.880 58.735 ;
        RECT 42.115 58.625 42.340 59.405 ;
        RECT 41.710 58.010 41.940 58.340 ;
        RECT 39.805 57.025 41.015 57.775 ;
        RECT 41.710 57.745 41.880 58.010 ;
        RECT 41.275 57.575 41.880 57.745 ;
        RECT 41.275 57.285 41.445 57.575 ;
        RECT 41.615 57.025 41.945 57.405 ;
        RECT 42.115 57.285 42.285 58.625 ;
        RECT 42.575 58.605 42.905 59.355 ;
        RECT 43.075 58.775 43.390 59.575 ;
        RECT 44.020 59.195 44.770 59.365 ;
        RECT 42.575 58.435 43.260 58.605 ;
        RECT 42.580 57.895 42.910 58.265 ;
        RECT 43.090 58.035 43.260 58.435 ;
        RECT 43.590 58.295 43.875 58.945 ;
        RECT 44.045 58.355 44.385 58.935 ;
        RECT 43.090 57.725 43.460 58.035 ;
        RECT 44.045 57.975 44.215 58.355 ;
        RECT 44.600 58.265 44.770 59.195 ;
        RECT 44.940 59.075 45.240 59.575 ;
        RECT 45.460 58.805 45.680 59.375 ;
        RECT 44.960 58.475 45.680 58.805 ;
        RECT 45.510 58.265 45.680 58.475 ;
        RECT 45.860 58.435 46.145 59.575 ;
        RECT 46.315 58.580 46.565 59.395 ;
        RECT 46.735 58.695 46.995 59.575 ;
        RECT 46.315 58.435 46.600 58.580 ;
        RECT 46.430 58.265 46.600 58.435 ;
        RECT 44.600 58.105 45.320 58.265 ;
        RECT 42.655 57.705 43.460 57.725 ;
        RECT 42.655 57.555 43.260 57.705 ;
        RECT 43.835 57.645 44.215 57.975 ;
        RECT 44.450 57.935 45.320 58.105 ;
        RECT 45.510 57.935 46.260 58.265 ;
        RECT 46.430 57.935 46.995 58.265 ;
        RECT 42.655 57.285 42.825 57.555 ;
        RECT 44.450 57.475 44.620 57.935 ;
        RECT 45.510 57.765 45.680 57.935 ;
        RECT 46.430 57.765 46.600 57.935 ;
        RECT 47.165 57.855 47.685 59.405 ;
        RECT 47.855 58.850 48.185 59.575 ;
        RECT 42.995 57.025 43.325 57.385 ;
        RECT 43.960 57.305 44.620 57.475 ;
        RECT 44.860 57.025 45.190 57.765 ;
        RECT 45.460 57.355 45.680 57.765 ;
        RECT 45.860 57.025 46.145 57.765 ;
        RECT 46.315 57.625 46.600 57.765 ;
        RECT 46.315 57.355 46.565 57.625 ;
        RECT 46.735 57.025 46.995 57.490 ;
        RECT 47.345 57.025 47.685 57.685 ;
        RECT 47.855 57.195 48.375 58.680 ;
        RECT 48.545 58.410 48.835 59.575 ;
        RECT 49.005 58.485 52.515 59.575 ;
        RECT 53.695 58.905 53.865 59.405 ;
        RECT 54.035 59.075 54.365 59.575 ;
        RECT 53.695 58.735 54.300 58.905 ;
        RECT 49.005 57.795 50.655 58.315 ;
        RECT 50.825 57.965 52.515 58.485 ;
        RECT 53.605 57.925 53.850 58.565 ;
        RECT 54.130 58.340 54.300 58.735 ;
        RECT 54.535 58.625 54.760 59.405 ;
        RECT 54.130 58.010 54.360 58.340 ;
        RECT 48.545 57.025 48.835 57.750 ;
        RECT 49.005 57.025 52.515 57.795 ;
        RECT 54.130 57.745 54.300 58.010 ;
        RECT 53.695 57.575 54.300 57.745 ;
        RECT 53.695 57.285 53.865 57.575 ;
        RECT 54.035 57.025 54.365 57.405 ;
        RECT 54.535 57.285 54.705 58.625 ;
        RECT 54.995 58.605 55.325 59.355 ;
        RECT 55.495 58.775 55.810 59.575 ;
        RECT 56.440 59.195 57.190 59.365 ;
        RECT 54.995 58.435 55.680 58.605 ;
        RECT 55.000 57.895 55.330 58.265 ;
        RECT 55.510 58.035 55.680 58.435 ;
        RECT 56.010 58.295 56.295 58.945 ;
        RECT 56.465 58.355 56.805 58.935 ;
        RECT 55.510 57.725 55.880 58.035 ;
        RECT 56.465 57.975 56.635 58.355 ;
        RECT 57.020 58.265 57.190 59.195 ;
        RECT 57.360 59.075 57.660 59.575 ;
        RECT 57.880 58.805 58.100 59.375 ;
        RECT 57.380 58.475 58.100 58.805 ;
        RECT 57.930 58.265 58.100 58.475 ;
        RECT 58.280 58.435 58.565 59.575 ;
        RECT 58.735 58.580 58.985 59.395 ;
        RECT 59.155 58.695 59.415 59.575 ;
        RECT 58.735 58.435 59.020 58.580 ;
        RECT 58.850 58.265 59.020 58.435 ;
        RECT 57.020 58.105 57.740 58.265 ;
        RECT 55.075 57.705 55.880 57.725 ;
        RECT 55.075 57.555 55.680 57.705 ;
        RECT 56.255 57.645 56.635 57.975 ;
        RECT 56.870 57.935 57.740 58.105 ;
        RECT 57.930 57.935 58.680 58.265 ;
        RECT 58.850 57.935 59.415 58.265 ;
        RECT 55.075 57.285 55.245 57.555 ;
        RECT 56.870 57.475 57.040 57.935 ;
        RECT 57.930 57.765 58.100 57.935 ;
        RECT 58.850 57.765 59.020 57.935 ;
        RECT 59.585 57.855 60.105 59.405 ;
        RECT 60.275 58.850 60.605 59.575 ;
        RECT 55.415 57.025 55.745 57.385 ;
        RECT 56.380 57.305 57.040 57.475 ;
        RECT 57.280 57.025 57.610 57.765 ;
        RECT 57.880 57.355 58.100 57.765 ;
        RECT 58.280 57.025 58.565 57.765 ;
        RECT 58.735 57.625 59.020 57.765 ;
        RECT 58.735 57.355 58.985 57.625 ;
        RECT 59.155 57.025 59.415 57.490 ;
        RECT 59.765 57.025 60.105 57.685 ;
        RECT 60.275 57.195 60.795 58.680 ;
        RECT 61.425 58.410 61.715 59.575 ;
        RECT 61.885 58.485 64.475 59.575 ;
        RECT 61.885 57.795 63.095 58.315 ;
        RECT 63.265 57.965 64.475 58.485 ;
        RECT 65.105 57.855 65.625 59.405 ;
        RECT 65.795 58.850 66.125 59.575 ;
        RECT 67.035 58.905 67.205 59.405 ;
        RECT 67.375 59.075 67.705 59.575 ;
        RECT 67.035 58.735 67.640 58.905 ;
        RECT 61.425 57.025 61.715 57.750 ;
        RECT 61.885 57.025 64.475 57.795 ;
        RECT 65.285 57.025 65.625 57.685 ;
        RECT 65.795 57.195 66.315 58.680 ;
        RECT 66.945 57.925 67.190 58.565 ;
        RECT 67.470 58.340 67.640 58.735 ;
        RECT 67.875 58.625 68.100 59.405 ;
        RECT 67.470 58.010 67.700 58.340 ;
        RECT 67.470 57.745 67.640 58.010 ;
        RECT 67.035 57.575 67.640 57.745 ;
        RECT 67.035 57.285 67.205 57.575 ;
        RECT 67.375 57.025 67.705 57.405 ;
        RECT 67.875 57.285 68.045 58.625 ;
        RECT 68.335 58.605 68.665 59.355 ;
        RECT 68.835 58.775 69.150 59.575 ;
        RECT 69.780 59.195 70.530 59.365 ;
        RECT 68.335 58.435 69.020 58.605 ;
        RECT 68.340 57.895 68.670 58.265 ;
        RECT 68.850 58.035 69.020 58.435 ;
        RECT 69.350 58.295 69.635 58.945 ;
        RECT 69.805 58.355 70.145 58.935 ;
        RECT 68.850 57.725 69.220 58.035 ;
        RECT 69.805 57.975 69.975 58.355 ;
        RECT 70.360 58.265 70.530 59.195 ;
        RECT 70.700 59.075 71.000 59.575 ;
        RECT 71.220 58.805 71.440 59.375 ;
        RECT 70.720 58.475 71.440 58.805 ;
        RECT 71.270 58.265 71.440 58.475 ;
        RECT 71.620 58.435 71.905 59.575 ;
        RECT 72.075 58.580 72.325 59.395 ;
        RECT 72.495 58.695 72.755 59.575 ;
        RECT 72.075 58.435 72.360 58.580 ;
        RECT 72.925 58.485 74.135 59.575 ;
        RECT 72.190 58.265 72.360 58.435 ;
        RECT 70.360 58.105 71.080 58.265 ;
        RECT 68.415 57.705 69.220 57.725 ;
        RECT 68.415 57.555 69.020 57.705 ;
        RECT 69.595 57.645 69.975 57.975 ;
        RECT 70.210 57.935 71.080 58.105 ;
        RECT 71.270 57.935 72.020 58.265 ;
        RECT 72.190 57.935 72.755 58.265 ;
        RECT 68.415 57.285 68.585 57.555 ;
        RECT 70.210 57.475 70.380 57.935 ;
        RECT 71.270 57.765 71.440 57.935 ;
        RECT 72.190 57.765 72.360 57.935 ;
        RECT 68.755 57.025 69.085 57.385 ;
        RECT 69.720 57.305 70.380 57.475 ;
        RECT 70.620 57.025 70.950 57.765 ;
        RECT 71.220 57.355 71.440 57.765 ;
        RECT 71.620 57.025 71.905 57.765 ;
        RECT 72.075 57.625 72.360 57.765 ;
        RECT 72.925 57.775 73.445 58.315 ;
        RECT 73.615 57.945 74.135 58.485 ;
        RECT 74.305 58.410 74.595 59.575 ;
        RECT 74.855 58.905 75.025 59.405 ;
        RECT 75.195 59.075 75.525 59.575 ;
        RECT 74.855 58.735 75.460 58.905 ;
        RECT 74.765 57.925 75.010 58.565 ;
        RECT 75.290 58.340 75.460 58.735 ;
        RECT 75.695 58.625 75.920 59.405 ;
        RECT 75.290 58.010 75.520 58.340 ;
        RECT 72.075 57.355 72.325 57.625 ;
        RECT 72.495 57.025 72.755 57.490 ;
        RECT 72.925 57.025 74.135 57.775 ;
        RECT 74.305 57.025 74.595 57.750 ;
        RECT 75.290 57.745 75.460 58.010 ;
        RECT 74.855 57.575 75.460 57.745 ;
        RECT 74.855 57.285 75.025 57.575 ;
        RECT 75.195 57.025 75.525 57.405 ;
        RECT 75.695 57.285 75.865 58.625 ;
        RECT 76.155 58.605 76.485 59.355 ;
        RECT 76.655 58.775 76.970 59.575 ;
        RECT 77.600 59.195 78.350 59.365 ;
        RECT 76.155 58.435 76.840 58.605 ;
        RECT 76.160 57.895 76.490 58.265 ;
        RECT 76.670 58.035 76.840 58.435 ;
        RECT 77.170 58.295 77.455 58.945 ;
        RECT 77.625 58.355 77.965 58.935 ;
        RECT 76.670 57.725 77.040 58.035 ;
        RECT 77.625 57.975 77.795 58.355 ;
        RECT 78.180 58.265 78.350 59.195 ;
        RECT 78.520 59.075 78.820 59.575 ;
        RECT 79.040 58.805 79.260 59.375 ;
        RECT 78.540 58.475 79.260 58.805 ;
        RECT 79.090 58.265 79.260 58.475 ;
        RECT 79.440 58.435 79.725 59.575 ;
        RECT 79.895 58.580 80.145 59.395 ;
        RECT 80.315 58.695 80.575 59.575 ;
        RECT 81.295 58.905 81.465 59.405 ;
        RECT 81.635 59.075 81.965 59.575 ;
        RECT 81.295 58.735 81.900 58.905 ;
        RECT 79.895 58.435 80.180 58.580 ;
        RECT 80.010 58.265 80.180 58.435 ;
        RECT 78.180 58.105 78.900 58.265 ;
        RECT 76.235 57.705 77.040 57.725 ;
        RECT 76.235 57.555 76.840 57.705 ;
        RECT 77.415 57.645 77.795 57.975 ;
        RECT 78.030 57.935 78.900 58.105 ;
        RECT 79.090 57.935 79.840 58.265 ;
        RECT 80.010 57.935 80.575 58.265 ;
        RECT 76.235 57.285 76.405 57.555 ;
        RECT 78.030 57.475 78.200 57.935 ;
        RECT 79.090 57.765 79.260 57.935 ;
        RECT 80.010 57.765 80.180 57.935 ;
        RECT 81.205 57.925 81.450 58.565 ;
        RECT 81.730 58.340 81.900 58.735 ;
        RECT 82.135 58.625 82.360 59.405 ;
        RECT 81.730 58.010 81.960 58.340 ;
        RECT 76.575 57.025 76.905 57.385 ;
        RECT 77.540 57.305 78.200 57.475 ;
        RECT 78.440 57.025 78.770 57.765 ;
        RECT 79.040 57.355 79.260 57.765 ;
        RECT 79.440 57.025 79.725 57.765 ;
        RECT 79.895 57.625 80.180 57.765 ;
        RECT 81.730 57.745 81.900 58.010 ;
        RECT 79.895 57.355 80.145 57.625 ;
        RECT 81.295 57.575 81.900 57.745 ;
        RECT 80.315 57.025 80.575 57.490 ;
        RECT 81.295 57.285 81.465 57.575 ;
        RECT 81.635 57.025 81.965 57.405 ;
        RECT 82.135 57.285 82.305 58.625 ;
        RECT 82.595 58.605 82.925 59.355 ;
        RECT 83.095 58.775 83.410 59.575 ;
        RECT 84.040 59.195 84.790 59.365 ;
        RECT 82.595 58.435 83.280 58.605 ;
        RECT 82.600 57.895 82.930 58.265 ;
        RECT 83.110 58.035 83.280 58.435 ;
        RECT 83.610 58.295 83.895 58.945 ;
        RECT 84.065 58.355 84.405 58.935 ;
        RECT 83.110 57.725 83.480 58.035 ;
        RECT 84.065 57.975 84.235 58.355 ;
        RECT 84.620 58.265 84.790 59.195 ;
        RECT 84.960 59.075 85.260 59.575 ;
        RECT 85.480 58.805 85.700 59.375 ;
        RECT 84.980 58.475 85.700 58.805 ;
        RECT 85.530 58.265 85.700 58.475 ;
        RECT 85.880 58.435 86.165 59.575 ;
        RECT 86.335 58.580 86.585 59.395 ;
        RECT 86.755 58.695 87.015 59.575 ;
        RECT 86.335 58.435 86.620 58.580 ;
        RECT 86.450 58.265 86.620 58.435 ;
        RECT 87.185 58.410 87.475 59.575 ;
        RECT 84.620 58.105 85.340 58.265 ;
        RECT 82.675 57.705 83.480 57.725 ;
        RECT 82.675 57.555 83.280 57.705 ;
        RECT 83.855 57.645 84.235 57.975 ;
        RECT 84.470 57.935 85.340 58.105 ;
        RECT 85.530 57.935 86.280 58.265 ;
        RECT 86.450 57.935 87.015 58.265 ;
        RECT 82.675 57.285 82.845 57.555 ;
        RECT 84.470 57.475 84.640 57.935 ;
        RECT 85.530 57.765 85.700 57.935 ;
        RECT 86.450 57.765 86.620 57.935 ;
        RECT 88.105 57.855 88.625 59.405 ;
        RECT 88.795 58.850 89.125 59.575 ;
        RECT 90.035 58.905 90.205 59.405 ;
        RECT 90.375 59.075 90.705 59.575 ;
        RECT 90.035 58.735 90.640 58.905 ;
        RECT 83.015 57.025 83.345 57.385 ;
        RECT 83.980 57.305 84.640 57.475 ;
        RECT 84.880 57.025 85.210 57.765 ;
        RECT 85.480 57.355 85.700 57.765 ;
        RECT 85.880 57.025 86.165 57.765 ;
        RECT 86.335 57.625 86.620 57.765 ;
        RECT 86.335 57.355 86.585 57.625 ;
        RECT 86.755 57.025 87.015 57.490 ;
        RECT 87.185 57.025 87.475 57.750 ;
        RECT 88.285 57.025 88.625 57.685 ;
        RECT 88.795 57.195 89.315 58.680 ;
        RECT 89.945 57.925 90.190 58.565 ;
        RECT 90.470 58.340 90.640 58.735 ;
        RECT 90.875 58.625 91.100 59.405 ;
        RECT 90.470 58.010 90.700 58.340 ;
        RECT 90.470 57.745 90.640 58.010 ;
        RECT 90.035 57.575 90.640 57.745 ;
        RECT 90.035 57.285 90.205 57.575 ;
        RECT 90.375 57.025 90.705 57.405 ;
        RECT 90.875 57.285 91.045 58.625 ;
        RECT 91.335 58.605 91.665 59.355 ;
        RECT 91.835 58.775 92.150 59.575 ;
        RECT 92.780 59.195 93.530 59.365 ;
        RECT 91.335 58.435 92.020 58.605 ;
        RECT 91.340 57.895 91.670 58.265 ;
        RECT 91.850 58.035 92.020 58.435 ;
        RECT 92.350 58.295 92.635 58.945 ;
        RECT 92.805 58.355 93.145 58.935 ;
        RECT 91.850 57.725 92.220 58.035 ;
        RECT 92.805 57.975 92.975 58.355 ;
        RECT 93.360 58.265 93.530 59.195 ;
        RECT 93.700 59.075 94.000 59.575 ;
        RECT 94.220 58.805 94.440 59.375 ;
        RECT 93.720 58.475 94.440 58.805 ;
        RECT 94.270 58.265 94.440 58.475 ;
        RECT 94.620 58.435 94.905 59.575 ;
        RECT 95.075 58.580 95.325 59.395 ;
        RECT 95.495 58.695 95.755 59.575 ;
        RECT 95.075 58.435 95.360 58.580 ;
        RECT 95.925 58.485 99.435 59.575 ;
        RECT 95.190 58.265 95.360 58.435 ;
        RECT 93.360 58.105 94.080 58.265 ;
        RECT 91.415 57.705 92.220 57.725 ;
        RECT 91.415 57.555 92.020 57.705 ;
        RECT 92.595 57.645 92.975 57.975 ;
        RECT 93.210 57.935 94.080 58.105 ;
        RECT 94.270 57.935 95.020 58.265 ;
        RECT 95.190 57.935 95.755 58.265 ;
        RECT 91.415 57.285 91.585 57.555 ;
        RECT 93.210 57.475 93.380 57.935 ;
        RECT 94.270 57.765 94.440 57.935 ;
        RECT 95.190 57.765 95.360 57.935 ;
        RECT 91.755 57.025 92.085 57.385 ;
        RECT 92.720 57.305 93.380 57.475 ;
        RECT 93.620 57.025 93.950 57.765 ;
        RECT 94.220 57.355 94.440 57.765 ;
        RECT 94.620 57.025 94.905 57.765 ;
        RECT 95.075 57.625 95.360 57.765 ;
        RECT 95.925 57.795 97.575 58.315 ;
        RECT 97.745 57.965 99.435 58.485 ;
        RECT 100.065 58.410 100.355 59.575 ;
        RECT 101.075 58.905 101.245 59.405 ;
        RECT 101.415 59.075 101.745 59.575 ;
        RECT 101.075 58.735 101.680 58.905 ;
        RECT 100.985 57.925 101.230 58.565 ;
        RECT 101.510 58.340 101.680 58.735 ;
        RECT 101.915 58.625 102.140 59.405 ;
        RECT 101.510 58.010 101.740 58.340 ;
        RECT 95.075 57.355 95.325 57.625 ;
        RECT 95.495 57.025 95.755 57.490 ;
        RECT 95.925 57.025 99.435 57.795 ;
        RECT 100.065 57.025 100.355 57.750 ;
        RECT 101.510 57.745 101.680 58.010 ;
        RECT 101.075 57.575 101.680 57.745 ;
        RECT 101.075 57.285 101.245 57.575 ;
        RECT 101.415 57.025 101.745 57.405 ;
        RECT 101.915 57.285 102.085 58.625 ;
        RECT 102.375 58.605 102.705 59.355 ;
        RECT 102.875 58.775 103.190 59.575 ;
        RECT 103.820 59.195 104.570 59.365 ;
        RECT 102.375 58.435 103.060 58.605 ;
        RECT 102.380 57.895 102.710 58.265 ;
        RECT 102.890 58.035 103.060 58.435 ;
        RECT 103.390 58.295 103.675 58.945 ;
        RECT 103.845 58.355 104.185 58.935 ;
        RECT 102.890 57.725 103.260 58.035 ;
        RECT 103.845 57.975 104.015 58.355 ;
        RECT 104.400 58.265 104.570 59.195 ;
        RECT 104.740 59.075 105.040 59.575 ;
        RECT 105.260 58.805 105.480 59.375 ;
        RECT 104.760 58.475 105.480 58.805 ;
        RECT 105.310 58.265 105.480 58.475 ;
        RECT 105.660 58.435 105.945 59.575 ;
        RECT 106.115 58.580 106.365 59.395 ;
        RECT 106.535 58.695 106.795 59.575 ;
        RECT 107.055 58.905 107.225 59.405 ;
        RECT 107.395 59.075 107.725 59.575 ;
        RECT 107.055 58.735 107.660 58.905 ;
        RECT 106.115 58.435 106.400 58.580 ;
        RECT 106.230 58.265 106.400 58.435 ;
        RECT 104.400 58.105 105.120 58.265 ;
        RECT 102.455 57.705 103.260 57.725 ;
        RECT 102.455 57.555 103.060 57.705 ;
        RECT 103.635 57.645 104.015 57.975 ;
        RECT 104.250 57.935 105.120 58.105 ;
        RECT 105.310 57.935 106.060 58.265 ;
        RECT 106.230 57.935 106.795 58.265 ;
        RECT 102.455 57.285 102.625 57.555 ;
        RECT 104.250 57.475 104.420 57.935 ;
        RECT 105.310 57.765 105.480 57.935 ;
        RECT 106.230 57.765 106.400 57.935 ;
        RECT 106.965 57.925 107.210 58.565 ;
        RECT 107.490 58.340 107.660 58.735 ;
        RECT 107.895 58.625 108.120 59.405 ;
        RECT 107.490 58.010 107.720 58.340 ;
        RECT 102.795 57.025 103.125 57.385 ;
        RECT 103.760 57.305 104.420 57.475 ;
        RECT 104.660 57.025 104.990 57.765 ;
        RECT 105.260 57.355 105.480 57.765 ;
        RECT 105.660 57.025 105.945 57.765 ;
        RECT 106.115 57.625 106.400 57.765 ;
        RECT 107.490 57.745 107.660 58.010 ;
        RECT 106.115 57.355 106.365 57.625 ;
        RECT 107.055 57.575 107.660 57.745 ;
        RECT 106.535 57.025 106.795 57.490 ;
        RECT 107.055 57.285 107.225 57.575 ;
        RECT 107.395 57.025 107.725 57.405 ;
        RECT 107.895 57.285 108.065 58.625 ;
        RECT 108.355 58.605 108.685 59.355 ;
        RECT 108.855 58.775 109.170 59.575 ;
        RECT 109.800 59.195 110.550 59.365 ;
        RECT 108.355 58.435 109.040 58.605 ;
        RECT 108.360 57.895 108.690 58.265 ;
        RECT 108.870 58.035 109.040 58.435 ;
        RECT 109.370 58.295 109.655 58.945 ;
        RECT 109.825 58.355 110.165 58.935 ;
        RECT 108.870 57.725 109.240 58.035 ;
        RECT 109.825 57.975 109.995 58.355 ;
        RECT 110.380 58.265 110.550 59.195 ;
        RECT 110.720 59.075 111.020 59.575 ;
        RECT 111.240 58.805 111.460 59.375 ;
        RECT 110.740 58.475 111.460 58.805 ;
        RECT 111.290 58.265 111.460 58.475 ;
        RECT 111.640 58.435 111.925 59.575 ;
        RECT 112.095 58.580 112.345 59.395 ;
        RECT 112.515 58.695 112.775 59.575 ;
        RECT 112.095 58.435 112.380 58.580 ;
        RECT 112.210 58.265 112.380 58.435 ;
        RECT 112.945 58.410 113.235 59.575 ;
        RECT 113.495 58.905 113.665 59.405 ;
        RECT 113.835 59.075 114.165 59.575 ;
        RECT 113.495 58.735 114.100 58.905 ;
        RECT 110.380 58.105 111.100 58.265 ;
        RECT 108.435 57.705 109.240 57.725 ;
        RECT 108.435 57.555 109.040 57.705 ;
        RECT 109.615 57.645 109.995 57.975 ;
        RECT 110.230 57.935 111.100 58.105 ;
        RECT 111.290 57.935 112.040 58.265 ;
        RECT 112.210 57.935 112.775 58.265 ;
        RECT 108.435 57.285 108.605 57.555 ;
        RECT 110.230 57.475 110.400 57.935 ;
        RECT 111.290 57.765 111.460 57.935 ;
        RECT 112.210 57.765 112.380 57.935 ;
        RECT 113.405 57.925 113.650 58.565 ;
        RECT 113.930 58.340 114.100 58.735 ;
        RECT 114.335 58.625 114.560 59.405 ;
        RECT 113.930 58.010 114.160 58.340 ;
        RECT 108.775 57.025 109.105 57.385 ;
        RECT 109.740 57.305 110.400 57.475 ;
        RECT 110.640 57.025 110.970 57.765 ;
        RECT 111.240 57.355 111.460 57.765 ;
        RECT 111.640 57.025 111.925 57.765 ;
        RECT 112.095 57.625 112.380 57.765 ;
        RECT 112.095 57.355 112.345 57.625 ;
        RECT 112.515 57.025 112.775 57.490 ;
        RECT 112.945 57.025 113.235 57.750 ;
        RECT 113.930 57.745 114.100 58.010 ;
        RECT 113.495 57.575 114.100 57.745 ;
        RECT 113.495 57.285 113.665 57.575 ;
        RECT 113.835 57.025 114.165 57.405 ;
        RECT 114.335 57.285 114.505 58.625 ;
        RECT 114.795 58.605 115.125 59.355 ;
        RECT 115.295 58.775 115.610 59.575 ;
        RECT 116.240 59.195 116.990 59.365 ;
        RECT 114.795 58.435 115.480 58.605 ;
        RECT 114.800 57.895 115.130 58.265 ;
        RECT 115.310 58.035 115.480 58.435 ;
        RECT 115.810 58.295 116.095 58.945 ;
        RECT 116.265 58.355 116.605 58.935 ;
        RECT 115.310 57.725 115.680 58.035 ;
        RECT 116.265 57.975 116.435 58.355 ;
        RECT 116.820 58.265 116.990 59.195 ;
        RECT 117.160 59.075 117.460 59.575 ;
        RECT 117.680 58.805 117.900 59.375 ;
        RECT 117.180 58.475 117.900 58.805 ;
        RECT 117.730 58.265 117.900 58.475 ;
        RECT 118.080 58.435 118.365 59.575 ;
        RECT 118.535 58.580 118.785 59.395 ;
        RECT 118.955 58.695 119.215 59.575 ;
        RECT 119.935 58.905 120.105 59.405 ;
        RECT 120.275 59.075 120.605 59.575 ;
        RECT 119.935 58.735 120.540 58.905 ;
        RECT 118.535 58.435 118.820 58.580 ;
        RECT 118.650 58.265 118.820 58.435 ;
        RECT 116.820 58.105 117.540 58.265 ;
        RECT 114.875 57.705 115.680 57.725 ;
        RECT 114.875 57.555 115.480 57.705 ;
        RECT 116.055 57.645 116.435 57.975 ;
        RECT 116.670 57.935 117.540 58.105 ;
        RECT 117.730 57.935 118.480 58.265 ;
        RECT 118.650 57.935 119.215 58.265 ;
        RECT 114.875 57.285 115.045 57.555 ;
        RECT 116.670 57.475 116.840 57.935 ;
        RECT 117.730 57.765 117.900 57.935 ;
        RECT 118.650 57.765 118.820 57.935 ;
        RECT 119.845 57.925 120.090 58.565 ;
        RECT 120.370 58.340 120.540 58.735 ;
        RECT 120.775 58.625 121.000 59.405 ;
        RECT 120.370 58.010 120.600 58.340 ;
        RECT 115.215 57.025 115.545 57.385 ;
        RECT 116.180 57.305 116.840 57.475 ;
        RECT 117.080 57.025 117.410 57.765 ;
        RECT 117.680 57.355 117.900 57.765 ;
        RECT 118.080 57.025 118.365 57.765 ;
        RECT 118.535 57.625 118.820 57.765 ;
        RECT 120.370 57.745 120.540 58.010 ;
        RECT 118.535 57.355 118.785 57.625 ;
        RECT 119.935 57.575 120.540 57.745 ;
        RECT 118.955 57.025 119.215 57.490 ;
        RECT 119.935 57.285 120.105 57.575 ;
        RECT 120.275 57.025 120.605 57.405 ;
        RECT 120.775 57.285 120.945 58.625 ;
        RECT 121.235 58.605 121.565 59.355 ;
        RECT 121.735 58.775 122.050 59.575 ;
        RECT 122.680 59.195 123.430 59.365 ;
        RECT 121.235 58.435 121.920 58.605 ;
        RECT 121.240 57.895 121.570 58.265 ;
        RECT 121.750 58.035 121.920 58.435 ;
        RECT 122.250 58.295 122.535 58.945 ;
        RECT 122.705 58.355 123.045 58.935 ;
        RECT 121.750 57.725 122.120 58.035 ;
        RECT 122.705 57.975 122.875 58.355 ;
        RECT 123.260 58.265 123.430 59.195 ;
        RECT 123.600 59.075 123.900 59.575 ;
        RECT 124.120 58.805 124.340 59.375 ;
        RECT 123.620 58.475 124.340 58.805 ;
        RECT 124.170 58.265 124.340 58.475 ;
        RECT 124.520 58.435 124.805 59.575 ;
        RECT 124.975 58.580 125.225 59.395 ;
        RECT 125.395 58.695 125.655 59.575 ;
        RECT 124.975 58.435 125.260 58.580 ;
        RECT 125.090 58.265 125.260 58.435 ;
        RECT 125.825 58.410 126.115 59.575 ;
        RECT 123.260 58.105 123.980 58.265 ;
        RECT 121.315 57.705 122.120 57.725 ;
        RECT 121.315 57.555 121.920 57.705 ;
        RECT 122.495 57.645 122.875 57.975 ;
        RECT 123.110 57.935 123.980 58.105 ;
        RECT 124.170 57.935 124.920 58.265 ;
        RECT 125.090 57.935 125.655 58.265 ;
        RECT 121.315 57.285 121.485 57.555 ;
        RECT 123.110 57.475 123.280 57.935 ;
        RECT 124.170 57.765 124.340 57.935 ;
        RECT 125.090 57.765 125.260 57.935 ;
        RECT 126.285 57.855 126.805 59.405 ;
        RECT 126.975 58.850 127.305 59.575 ;
        RECT 121.655 57.025 121.985 57.385 ;
        RECT 122.620 57.305 123.280 57.475 ;
        RECT 123.520 57.025 123.850 57.765 ;
        RECT 124.120 57.355 124.340 57.765 ;
        RECT 124.520 57.025 124.805 57.765 ;
        RECT 124.975 57.625 125.260 57.765 ;
        RECT 124.975 57.355 125.225 57.625 ;
        RECT 125.395 57.025 125.655 57.490 ;
        RECT 125.825 57.025 126.115 57.750 ;
        RECT 126.465 57.025 126.805 57.685 ;
        RECT 126.975 57.195 127.495 58.680 ;
        RECT 127.665 57.855 128.185 59.405 ;
        RECT 128.355 58.850 128.685 59.575 ;
        RECT 127.845 57.025 128.185 57.685 ;
        RECT 128.355 57.195 128.875 58.680 ;
        RECT 129.045 58.485 130.715 59.575 ;
        RECT 130.975 58.905 131.145 59.405 ;
        RECT 131.315 59.075 131.645 59.575 ;
        RECT 130.975 58.735 131.580 58.905 ;
        RECT 129.045 57.795 129.795 58.315 ;
        RECT 129.965 57.965 130.715 58.485 ;
        RECT 130.885 57.925 131.130 58.565 ;
        RECT 131.410 58.340 131.580 58.735 ;
        RECT 131.815 58.625 132.040 59.405 ;
        RECT 131.410 58.010 131.640 58.340 ;
        RECT 129.045 57.025 130.715 57.795 ;
        RECT 131.410 57.745 131.580 58.010 ;
        RECT 130.975 57.575 131.580 57.745 ;
        RECT 130.975 57.285 131.145 57.575 ;
        RECT 131.315 57.025 131.645 57.405 ;
        RECT 131.815 57.285 131.985 58.625 ;
        RECT 132.275 58.605 132.605 59.355 ;
        RECT 132.775 58.775 133.090 59.575 ;
        RECT 133.720 59.195 134.470 59.365 ;
        RECT 132.275 58.435 132.960 58.605 ;
        RECT 132.280 57.895 132.610 58.265 ;
        RECT 132.790 58.035 132.960 58.435 ;
        RECT 133.290 58.295 133.575 58.945 ;
        RECT 133.745 58.355 134.085 58.935 ;
        RECT 132.790 57.725 133.160 58.035 ;
        RECT 133.745 57.975 133.915 58.355 ;
        RECT 134.300 58.265 134.470 59.195 ;
        RECT 134.640 59.075 134.940 59.575 ;
        RECT 135.160 58.805 135.380 59.375 ;
        RECT 134.660 58.475 135.380 58.805 ;
        RECT 135.210 58.265 135.380 58.475 ;
        RECT 135.560 58.435 135.845 59.575 ;
        RECT 136.015 58.580 136.265 59.395 ;
        RECT 136.435 58.695 136.695 59.575 ;
        RECT 137.515 58.850 137.845 59.575 ;
        RECT 136.015 58.435 136.300 58.580 ;
        RECT 136.130 58.265 136.300 58.435 ;
        RECT 134.300 58.105 135.020 58.265 ;
        RECT 132.355 57.705 133.160 57.725 ;
        RECT 132.355 57.555 132.960 57.705 ;
        RECT 133.535 57.645 133.915 57.975 ;
        RECT 134.150 57.935 135.020 58.105 ;
        RECT 135.210 57.935 135.960 58.265 ;
        RECT 136.130 57.935 136.695 58.265 ;
        RECT 132.355 57.285 132.525 57.555 ;
        RECT 134.150 57.475 134.320 57.935 ;
        RECT 135.210 57.765 135.380 57.935 ;
        RECT 136.130 57.765 136.300 57.935 ;
        RECT 132.695 57.025 133.025 57.385 ;
        RECT 133.660 57.305 134.320 57.475 ;
        RECT 134.560 57.025 134.890 57.765 ;
        RECT 135.160 57.355 135.380 57.765 ;
        RECT 135.560 57.025 135.845 57.765 ;
        RECT 136.015 57.625 136.300 57.765 ;
        RECT 136.015 57.355 136.265 57.625 ;
        RECT 136.435 57.025 136.695 57.490 ;
        RECT 137.325 57.195 137.845 58.680 ;
        RECT 138.015 57.855 138.535 59.405 ;
        RECT 138.705 58.410 138.995 59.575 ;
        RECT 139.255 58.905 139.425 59.405 ;
        RECT 139.595 59.075 139.925 59.575 ;
        RECT 139.255 58.735 139.860 58.905 ;
        RECT 139.165 57.925 139.410 58.565 ;
        RECT 139.690 58.340 139.860 58.735 ;
        RECT 140.095 58.625 140.320 59.405 ;
        RECT 139.690 58.010 139.920 58.340 ;
        RECT 138.015 57.025 138.355 57.685 ;
        RECT 138.705 57.025 138.995 57.750 ;
        RECT 139.690 57.745 139.860 58.010 ;
        RECT 139.255 57.575 139.860 57.745 ;
        RECT 139.255 57.285 139.425 57.575 ;
        RECT 139.595 57.025 139.925 57.405 ;
        RECT 140.095 57.285 140.265 58.625 ;
        RECT 140.555 58.605 140.885 59.355 ;
        RECT 141.055 58.775 141.370 59.575 ;
        RECT 142.000 59.195 142.750 59.365 ;
        RECT 140.555 58.435 141.240 58.605 ;
        RECT 140.560 57.895 140.890 58.265 ;
        RECT 141.070 58.035 141.240 58.435 ;
        RECT 141.570 58.295 141.855 58.945 ;
        RECT 142.025 58.355 142.365 58.935 ;
        RECT 141.070 57.725 141.440 58.035 ;
        RECT 142.025 57.975 142.195 58.355 ;
        RECT 142.580 58.265 142.750 59.195 ;
        RECT 142.920 59.075 143.220 59.575 ;
        RECT 143.440 58.805 143.660 59.375 ;
        RECT 142.940 58.475 143.660 58.805 ;
        RECT 143.490 58.265 143.660 58.475 ;
        RECT 143.840 58.435 144.125 59.575 ;
        RECT 144.295 58.580 144.545 59.395 ;
        RECT 144.715 58.695 144.975 59.575 ;
        RECT 145.235 58.905 145.405 59.405 ;
        RECT 145.575 59.075 145.905 59.575 ;
        RECT 145.235 58.735 145.840 58.905 ;
        RECT 144.295 58.435 144.580 58.580 ;
        RECT 144.410 58.265 144.580 58.435 ;
        RECT 142.580 58.105 143.300 58.265 ;
        RECT 140.635 57.705 141.440 57.725 ;
        RECT 140.635 57.555 141.240 57.705 ;
        RECT 141.815 57.645 142.195 57.975 ;
        RECT 142.430 57.935 143.300 58.105 ;
        RECT 143.490 57.935 144.240 58.265 ;
        RECT 144.410 57.935 144.975 58.265 ;
        RECT 140.635 57.285 140.805 57.555 ;
        RECT 142.430 57.475 142.600 57.935 ;
        RECT 143.490 57.765 143.660 57.935 ;
        RECT 144.410 57.765 144.580 57.935 ;
        RECT 145.145 57.925 145.390 58.565 ;
        RECT 145.670 58.340 145.840 58.735 ;
        RECT 146.075 58.625 146.300 59.405 ;
        RECT 145.670 58.010 145.900 58.340 ;
        RECT 140.975 57.025 141.305 57.385 ;
        RECT 141.940 57.305 142.600 57.475 ;
        RECT 142.840 57.025 143.170 57.765 ;
        RECT 143.440 57.355 143.660 57.765 ;
        RECT 143.840 57.025 144.125 57.765 ;
        RECT 144.295 57.625 144.580 57.765 ;
        RECT 145.670 57.745 145.840 58.010 ;
        RECT 144.295 57.355 144.545 57.625 ;
        RECT 145.235 57.575 145.840 57.745 ;
        RECT 144.715 57.025 144.975 57.490 ;
        RECT 145.235 57.285 145.405 57.575 ;
        RECT 145.575 57.025 145.905 57.405 ;
        RECT 146.075 57.285 146.245 58.625 ;
        RECT 146.535 58.605 146.865 59.355 ;
        RECT 147.035 58.775 147.350 59.575 ;
        RECT 147.980 59.195 148.730 59.365 ;
        RECT 146.535 58.435 147.220 58.605 ;
        RECT 146.540 57.895 146.870 58.265 ;
        RECT 147.050 58.035 147.220 58.435 ;
        RECT 147.550 58.295 147.835 58.945 ;
        RECT 148.005 58.355 148.345 58.935 ;
        RECT 147.050 57.725 147.420 58.035 ;
        RECT 148.005 57.975 148.175 58.355 ;
        RECT 148.560 58.265 148.730 59.195 ;
        RECT 148.900 59.075 149.200 59.575 ;
        RECT 149.420 58.805 149.640 59.375 ;
        RECT 148.920 58.475 149.640 58.805 ;
        RECT 149.470 58.265 149.640 58.475 ;
        RECT 149.820 58.435 150.105 59.575 ;
        RECT 150.275 58.580 150.525 59.395 ;
        RECT 150.695 58.695 150.955 59.575 ;
        RECT 150.275 58.435 150.560 58.580 ;
        RECT 150.390 58.265 150.560 58.435 ;
        RECT 151.585 58.410 151.875 59.575 ;
        RECT 152.045 58.485 155.555 59.575 ;
        RECT 148.560 58.105 149.280 58.265 ;
        RECT 146.615 57.705 147.420 57.725 ;
        RECT 146.615 57.555 147.220 57.705 ;
        RECT 147.795 57.645 148.175 57.975 ;
        RECT 148.410 57.935 149.280 58.105 ;
        RECT 149.470 57.935 150.220 58.265 ;
        RECT 150.390 57.935 150.955 58.265 ;
        RECT 146.615 57.285 146.785 57.555 ;
        RECT 148.410 57.475 148.580 57.935 ;
        RECT 149.470 57.765 149.640 57.935 ;
        RECT 150.390 57.765 150.560 57.935 ;
        RECT 146.955 57.025 147.285 57.385 ;
        RECT 147.920 57.305 148.580 57.475 ;
        RECT 148.820 57.025 149.150 57.765 ;
        RECT 149.420 57.355 149.640 57.765 ;
        RECT 149.820 57.025 150.105 57.765 ;
        RECT 150.275 57.625 150.560 57.765 ;
        RECT 152.045 57.795 153.695 58.315 ;
        RECT 153.865 57.965 155.555 58.485 ;
        RECT 155.725 58.485 156.935 59.575 ;
        RECT 155.725 57.945 156.245 58.485 ;
        RECT 150.275 57.355 150.525 57.625 ;
        RECT 150.695 57.025 150.955 57.490 ;
        RECT 151.585 57.025 151.875 57.750 ;
        RECT 152.045 57.025 155.555 57.795 ;
        RECT 156.415 57.775 156.935 58.315 ;
        RECT 155.725 57.025 156.935 57.775 ;
        RECT 22.700 56.855 157.020 57.025 ;
        RECT 114.100 49.650 116.700 49.820 ;
        RECT 114.100 48.800 114.270 49.650 ;
        RECT 114.900 49.140 115.900 49.310 ;
        RECT 74.220 48.250 76.820 48.420 ;
        RECT 33.000 47.410 35.600 47.580 ;
        RECT 33.000 46.560 33.170 47.410 ;
        RECT 33.800 46.900 34.800 47.070 ;
        RECT 32.980 44.760 33.180 46.560 ;
        RECT 33.000 34.010 33.170 44.760 ;
        RECT 33.570 34.690 33.740 46.730 ;
        RECT 34.860 34.690 35.030 46.730 ;
        RECT 33.800 34.350 34.800 34.520 ;
        RECT 35.430 34.010 35.600 47.410 ;
        RECT 74.220 47.400 74.390 48.250 ;
        RECT 75.020 47.740 76.020 47.910 ;
        RECT 74.200 45.600 74.400 47.400 ;
        RECT 33.000 33.840 35.600 34.010 ;
        RECT 40.000 38.410 42.600 38.580 ;
        RECT 40.000 34.010 40.170 38.410 ;
        RECT 40.800 37.900 41.800 38.070 ;
        RECT 42.430 38.060 42.600 38.410 ;
        RECT 40.570 34.690 40.740 37.730 ;
        RECT 41.860 34.690 42.030 37.730 ;
        RECT 42.430 36.510 42.630 38.060 ;
        RECT 43.700 37.960 46.300 38.130 ;
        RECT 43.700 37.660 43.870 37.960 ;
        RECT 43.680 36.510 43.880 37.660 ;
        RECT 44.500 37.450 45.500 37.620 ;
        RECT 40.800 34.350 41.800 34.520 ;
        RECT 42.430 34.010 42.600 36.510 ;
        RECT 43.700 34.440 43.870 36.510 ;
        RECT 44.270 35.120 44.440 37.280 ;
        RECT 45.560 35.120 45.730 37.280 ;
        RECT 44.500 34.780 45.500 34.950 ;
        RECT 46.130 34.440 46.300 37.960 ;
        RECT 43.700 34.270 46.300 34.440 ;
        RECT 46.710 34.760 49.950 34.930 ;
        RECT 40.000 33.840 42.600 34.010 ;
        RECT 46.710 33.910 46.880 34.760 ;
        RECT 49.780 34.410 49.950 34.760 ;
        RECT 50.410 34.760 53.150 34.930 ;
        RECT 50.410 34.410 50.580 34.760 ;
        RECT 47.560 34.190 49.100 34.360 ;
        RECT 35.000 32.910 37.600 33.080 ;
        RECT 35.000 31.960 35.170 32.910 ;
        RECT 35.800 32.400 36.800 32.570 ;
        RECT 34.980 30.160 35.180 31.960 ;
        RECT 35.000 23.030 35.170 30.160 ;
        RECT 35.570 23.710 35.740 32.230 ;
        RECT 36.860 23.710 37.030 32.230 ;
        RECT 35.800 23.370 36.800 23.540 ;
        RECT 37.430 23.030 37.600 32.910 ;
        RECT 46.680 32.860 46.880 33.910 ;
        RECT 47.220 33.130 47.390 34.130 ;
        RECT 49.270 33.130 49.440 34.130 ;
        RECT 47.560 32.900 49.100 33.070 ;
        RECT 46.710 32.500 46.880 32.860 ;
        RECT 49.780 32.860 49.980 34.410 ;
        RECT 50.380 32.860 50.580 34.410 ;
        RECT 51.260 34.190 52.300 34.360 ;
        RECT 50.920 33.130 51.090 34.130 ;
        RECT 52.470 33.130 52.640 34.130 ;
        RECT 51.260 32.900 52.300 33.070 ;
        RECT 49.780 32.500 49.950 32.860 ;
        RECT 46.710 32.330 49.950 32.500 ;
        RECT 50.410 32.500 50.580 32.860 ;
        RECT 52.980 32.500 53.150 34.760 ;
        RECT 74.220 34.850 74.390 45.600 ;
        RECT 74.790 35.530 74.960 47.570 ;
        RECT 76.080 35.530 76.250 47.570 ;
        RECT 75.020 35.190 76.020 35.360 ;
        RECT 76.650 34.850 76.820 48.250 ;
        RECT 114.080 47.000 114.280 48.800 ;
        RECT 74.220 34.680 76.820 34.850 ;
        RECT 81.220 39.250 83.820 39.420 ;
        RECT 81.220 34.850 81.390 39.250 ;
        RECT 82.020 38.740 83.020 38.910 ;
        RECT 83.650 38.900 83.820 39.250 ;
        RECT 81.790 35.530 81.960 38.570 ;
        RECT 83.080 35.530 83.250 38.570 ;
        RECT 83.650 37.350 83.850 38.900 ;
        RECT 84.920 38.800 87.520 38.970 ;
        RECT 84.920 38.500 85.090 38.800 ;
        RECT 84.900 37.350 85.100 38.500 ;
        RECT 85.720 38.290 86.720 38.460 ;
        RECT 82.020 35.190 83.020 35.360 ;
        RECT 83.650 34.850 83.820 37.350 ;
        RECT 84.920 35.280 85.090 37.350 ;
        RECT 85.490 35.960 85.660 38.120 ;
        RECT 86.780 35.960 86.950 38.120 ;
        RECT 85.720 35.620 86.720 35.790 ;
        RECT 87.350 35.280 87.520 38.800 ;
        RECT 114.100 36.250 114.270 47.000 ;
        RECT 114.670 36.930 114.840 48.970 ;
        RECT 115.960 36.930 116.130 48.970 ;
        RECT 114.900 36.590 115.900 36.760 ;
        RECT 116.530 36.250 116.700 49.650 ;
        RECT 114.100 36.080 116.700 36.250 ;
        RECT 121.100 40.650 123.700 40.820 ;
        RECT 121.100 36.250 121.270 40.650 ;
        RECT 121.900 40.140 122.900 40.310 ;
        RECT 123.530 40.300 123.700 40.650 ;
        RECT 121.670 36.930 121.840 39.970 ;
        RECT 122.960 36.930 123.130 39.970 ;
        RECT 123.530 38.750 123.730 40.300 ;
        RECT 124.800 40.200 127.400 40.370 ;
        RECT 124.800 39.900 124.970 40.200 ;
        RECT 124.780 38.750 124.980 39.900 ;
        RECT 125.600 39.690 126.600 39.860 ;
        RECT 121.900 36.590 122.900 36.760 ;
        RECT 123.530 36.250 123.700 38.750 ;
        RECT 124.800 36.680 124.970 38.750 ;
        RECT 125.370 37.360 125.540 39.520 ;
        RECT 126.660 37.360 126.830 39.520 ;
        RECT 125.600 37.020 126.600 37.190 ;
        RECT 127.230 36.680 127.400 40.200 ;
        RECT 124.800 36.510 127.400 36.680 ;
        RECT 127.810 37.000 131.050 37.170 ;
        RECT 121.100 36.080 123.700 36.250 ;
        RECT 127.810 36.150 127.980 37.000 ;
        RECT 130.880 36.650 131.050 37.000 ;
        RECT 131.510 37.000 134.250 37.170 ;
        RECT 131.510 36.650 131.680 37.000 ;
        RECT 128.660 36.430 130.200 36.600 ;
        RECT 84.920 35.110 87.520 35.280 ;
        RECT 87.930 35.600 91.170 35.770 ;
        RECT 81.220 34.680 83.820 34.850 ;
        RECT 87.930 34.750 88.100 35.600 ;
        RECT 91.000 35.250 91.170 35.600 ;
        RECT 91.630 35.600 94.370 35.770 ;
        RECT 91.630 35.250 91.800 35.600 ;
        RECT 88.780 35.030 90.320 35.200 ;
        RECT 76.220 33.750 78.820 33.920 ;
        RECT 76.220 32.800 76.390 33.750 ;
        RECT 77.020 33.240 78.020 33.410 ;
        RECT 50.410 32.330 53.150 32.500 ;
        RECT 50.410 31.810 53.150 31.980 ;
        RECT 50.410 30.460 50.580 31.810 ;
        RECT 51.260 31.240 52.300 31.410 ;
        RECT 50.330 29.360 50.580 30.460 ;
        RECT 50.920 29.680 51.090 31.180 ;
        RECT 52.470 29.680 52.640 31.180 ;
        RECT 51.260 29.450 52.300 29.620 ;
        RECT 50.410 29.050 50.580 29.360 ;
        RECT 52.980 29.050 53.150 31.810 ;
        RECT 76.200 31.000 76.400 32.800 ;
        RECT 50.410 28.880 53.150 29.050 ;
        RECT 50.430 28.230 50.830 28.310 ;
        RECT 49.980 28.060 53.700 28.230 ;
        RECT 49.980 27.860 50.150 28.060 ;
        RECT 49.980 27.410 50.230 27.860 ;
        RECT 50.780 27.550 52.900 27.720 ;
        RECT 49.980 25.660 50.150 27.410 ;
        RECT 50.550 26.340 50.720 27.380 ;
        RECT 52.960 26.340 53.130 27.380 ;
        RECT 50.780 26.000 52.900 26.170 ;
        RECT 53.530 25.660 53.700 28.060 ;
        RECT 49.980 25.490 53.700 25.660 ;
        RECT 35.000 22.860 37.600 23.030 ;
        RECT 50.150 24.510 54.750 24.680 ;
        RECT 50.150 22.110 50.320 24.510 ;
        RECT 50.950 24.000 53.950 24.170 ;
        RECT 50.720 22.790 50.890 23.830 ;
        RECT 54.010 22.790 54.180 23.830 ;
        RECT 50.950 22.450 53.950 22.620 ;
        RECT 54.580 22.110 54.750 24.510 ;
        RECT 76.220 23.870 76.390 31.000 ;
        RECT 76.790 24.550 76.960 33.070 ;
        RECT 78.080 24.550 78.250 33.070 ;
        RECT 77.020 24.210 78.020 24.380 ;
        RECT 78.650 23.870 78.820 33.750 ;
        RECT 87.900 33.700 88.100 34.750 ;
        RECT 88.440 33.970 88.610 34.970 ;
        RECT 90.490 33.970 90.660 34.970 ;
        RECT 88.780 33.740 90.320 33.910 ;
        RECT 87.930 33.340 88.100 33.700 ;
        RECT 91.000 33.700 91.200 35.250 ;
        RECT 91.600 33.700 91.800 35.250 ;
        RECT 92.480 35.030 93.520 35.200 ;
        RECT 92.140 33.970 92.310 34.970 ;
        RECT 93.690 33.970 93.860 34.970 ;
        RECT 92.480 33.740 93.520 33.910 ;
        RECT 91.000 33.340 91.170 33.700 ;
        RECT 87.930 33.170 91.170 33.340 ;
        RECT 91.630 33.340 91.800 33.700 ;
        RECT 94.200 33.340 94.370 35.600 ;
        RECT 116.100 35.150 118.700 35.320 ;
        RECT 116.100 34.200 116.270 35.150 ;
        RECT 116.900 34.640 117.900 34.810 ;
        RECT 91.630 33.170 94.370 33.340 ;
        RECT 91.630 32.650 94.370 32.820 ;
        RECT 91.630 31.300 91.800 32.650 ;
        RECT 92.480 32.080 93.520 32.250 ;
        RECT 91.550 30.200 91.800 31.300 ;
        RECT 92.140 30.520 92.310 32.020 ;
        RECT 93.690 30.520 93.860 32.020 ;
        RECT 92.480 30.290 93.520 30.460 ;
        RECT 91.630 29.890 91.800 30.200 ;
        RECT 94.200 29.890 94.370 32.650 ;
        RECT 116.080 32.400 116.280 34.200 ;
        RECT 91.630 29.720 94.370 29.890 ;
        RECT 91.650 29.070 92.050 29.150 ;
        RECT 91.200 28.900 94.920 29.070 ;
        RECT 91.200 28.700 91.370 28.900 ;
        RECT 91.200 28.250 91.450 28.700 ;
        RECT 92.000 28.390 94.120 28.560 ;
        RECT 91.200 26.500 91.370 28.250 ;
        RECT 91.770 27.180 91.940 28.220 ;
        RECT 94.180 27.180 94.350 28.220 ;
        RECT 92.000 26.840 94.120 27.010 ;
        RECT 94.750 26.500 94.920 28.900 ;
        RECT 91.200 26.330 94.920 26.500 ;
        RECT 76.220 23.700 78.820 23.870 ;
        RECT 91.370 25.350 95.970 25.520 ;
        RECT 91.370 22.950 91.540 25.350 ;
        RECT 92.170 24.840 95.170 25.010 ;
        RECT 91.940 23.630 92.110 24.670 ;
        RECT 95.230 23.630 95.400 24.670 ;
        RECT 92.170 23.290 95.170 23.460 ;
        RECT 95.800 22.950 95.970 25.350 ;
        RECT 116.100 25.270 116.270 32.400 ;
        RECT 116.670 25.950 116.840 34.470 ;
        RECT 117.960 25.950 118.130 34.470 ;
        RECT 116.900 25.610 117.900 25.780 ;
        RECT 118.530 25.270 118.700 35.150 ;
        RECT 127.780 35.100 127.980 36.150 ;
        RECT 128.320 35.370 128.490 36.370 ;
        RECT 130.370 35.370 130.540 36.370 ;
        RECT 128.660 35.140 130.200 35.310 ;
        RECT 127.810 34.740 127.980 35.100 ;
        RECT 130.880 35.100 131.080 36.650 ;
        RECT 131.480 35.100 131.680 36.650 ;
        RECT 132.360 36.430 133.400 36.600 ;
        RECT 132.020 35.370 132.190 36.370 ;
        RECT 133.570 35.370 133.740 36.370 ;
        RECT 132.360 35.140 133.400 35.310 ;
        RECT 130.880 34.740 131.050 35.100 ;
        RECT 127.810 34.570 131.050 34.740 ;
        RECT 131.510 34.740 131.680 35.100 ;
        RECT 134.080 34.740 134.250 37.000 ;
        RECT 131.510 34.570 134.250 34.740 ;
        RECT 131.510 34.050 134.250 34.220 ;
        RECT 131.510 32.700 131.680 34.050 ;
        RECT 132.360 33.480 133.400 33.650 ;
        RECT 131.430 31.600 131.680 32.700 ;
        RECT 132.020 31.920 132.190 33.420 ;
        RECT 133.570 31.920 133.740 33.420 ;
        RECT 132.360 31.690 133.400 31.860 ;
        RECT 131.510 31.290 131.680 31.600 ;
        RECT 134.080 31.290 134.250 34.050 ;
        RECT 131.510 31.120 134.250 31.290 ;
        RECT 131.530 30.470 131.930 30.550 ;
        RECT 131.080 30.300 134.800 30.470 ;
        RECT 131.080 30.100 131.250 30.300 ;
        RECT 131.080 29.650 131.330 30.100 ;
        RECT 131.880 29.790 134.000 29.960 ;
        RECT 131.080 27.900 131.250 29.650 ;
        RECT 131.650 28.580 131.820 29.620 ;
        RECT 134.060 28.580 134.230 29.620 ;
        RECT 131.880 28.240 134.000 28.410 ;
        RECT 134.630 27.900 134.800 30.300 ;
        RECT 131.080 27.730 134.800 27.900 ;
        RECT 116.100 25.100 118.700 25.270 ;
        RECT 131.250 26.750 135.850 26.920 ;
        RECT 131.250 24.350 131.420 26.750 ;
        RECT 132.050 26.240 135.050 26.410 ;
        RECT 131.820 25.030 131.990 26.070 ;
        RECT 135.110 25.030 135.280 26.070 ;
        RECT 132.050 24.690 135.050 24.860 ;
        RECT 135.680 24.350 135.850 26.750 ;
        RECT 117.600 24.150 120.200 24.320 ;
        RECT 131.250 24.180 135.850 24.350 ;
        RECT 131.560 24.150 134.320 24.180 ;
        RECT 117.600 23.200 117.770 24.150 ;
        RECT 118.400 23.640 119.400 23.810 ;
        RECT 36.500 21.910 39.100 22.080 ;
        RECT 50.150 21.940 54.750 22.110 ;
        RECT 77.720 22.750 80.320 22.920 ;
        RECT 91.370 22.780 95.970 22.950 ;
        RECT 91.680 22.750 94.440 22.780 ;
        RECT 50.460 21.910 53.220 21.940 ;
        RECT 36.500 20.960 36.670 21.910 ;
        RECT 37.300 21.400 38.300 21.570 ;
        RECT 36.480 19.060 36.680 20.960 ;
        RECT 36.500 14.510 36.670 19.060 ;
        RECT 37.070 15.190 37.240 21.230 ;
        RECT 38.360 15.190 38.530 21.230 ;
        RECT 37.300 14.850 38.300 15.020 ;
        RECT 38.930 14.510 39.100 21.910 ;
        RECT 77.720 21.800 77.890 22.750 ;
        RECT 78.520 22.240 79.520 22.410 ;
        RECT 50.120 20.930 55.960 21.100 ;
        RECT 50.120 18.530 50.290 20.930 ;
        RECT 50.920 20.420 55.160 20.590 ;
        RECT 50.690 19.210 50.860 20.250 ;
        RECT 55.220 19.210 55.390 20.250 ;
        RECT 50.920 18.870 55.160 19.040 ;
        RECT 55.790 18.530 55.960 20.930 ;
        RECT 77.700 19.900 77.900 21.800 ;
        RECT 50.120 18.360 55.960 18.530 ;
        RECT 50.460 18.330 53.220 18.360 ;
        RECT 49.990 17.350 57.590 17.520 ;
        RECT 49.990 14.950 50.160 17.350 ;
        RECT 50.790 16.840 56.790 17.010 ;
        RECT 50.560 15.630 50.730 16.670 ;
        RECT 56.850 15.630 57.020 16.670 ;
        RECT 50.790 15.290 56.790 15.460 ;
        RECT 57.420 14.950 57.590 17.350 ;
        RECT 77.720 15.350 77.890 19.900 ;
        RECT 78.290 16.030 78.460 22.070 ;
        RECT 79.580 16.030 79.750 22.070 ;
        RECT 78.520 15.690 79.520 15.860 ;
        RECT 80.150 15.350 80.320 22.750 ;
        RECT 91.340 21.770 97.180 21.940 ;
        RECT 91.340 19.370 91.510 21.770 ;
        RECT 92.140 21.260 96.380 21.430 ;
        RECT 91.910 20.050 92.080 21.090 ;
        RECT 96.440 20.050 96.610 21.090 ;
        RECT 92.140 19.710 96.380 19.880 ;
        RECT 97.010 19.370 97.180 21.770 ;
        RECT 117.580 21.300 117.780 23.200 ;
        RECT 91.340 19.200 97.180 19.370 ;
        RECT 91.680 19.170 94.440 19.200 ;
        RECT 91.210 18.190 98.810 18.360 ;
        RECT 91.210 15.790 91.380 18.190 ;
        RECT 92.010 17.680 98.010 17.850 ;
        RECT 91.780 16.470 91.950 17.510 ;
        RECT 98.070 16.470 98.240 17.510 ;
        RECT 92.010 16.130 98.010 16.300 ;
        RECT 98.640 15.790 98.810 18.190 ;
        RECT 117.600 16.750 117.770 21.300 ;
        RECT 118.170 17.430 118.340 23.470 ;
        RECT 119.460 17.430 119.630 23.470 ;
        RECT 118.400 17.090 119.400 17.260 ;
        RECT 120.030 16.750 120.200 24.150 ;
        RECT 131.220 23.170 137.060 23.340 ;
        RECT 131.220 20.770 131.390 23.170 ;
        RECT 132.020 22.660 136.260 22.830 ;
        RECT 131.790 21.450 131.960 22.490 ;
        RECT 136.320 21.450 136.490 22.490 ;
        RECT 132.020 21.110 136.260 21.280 ;
        RECT 136.890 20.770 137.060 23.170 ;
        RECT 131.220 20.600 137.060 20.770 ;
        RECT 131.560 20.570 134.320 20.600 ;
        RECT 131.090 19.590 138.690 19.760 ;
        RECT 131.090 17.190 131.260 19.590 ;
        RECT 131.890 19.080 137.890 19.250 ;
        RECT 131.660 17.870 131.830 18.910 ;
        RECT 137.950 17.870 138.120 18.910 ;
        RECT 131.890 17.530 137.890 17.700 ;
        RECT 138.520 17.190 138.690 19.590 ;
        RECT 131.090 17.020 138.690 17.190 ;
        RECT 131.560 16.990 134.320 17.020 ;
        RECT 117.600 16.580 120.200 16.750 ;
        RECT 131.110 16.010 141.190 16.180 ;
        RECT 91.210 15.620 98.810 15.790 ;
        RECT 119.600 15.650 122.200 15.820 ;
        RECT 91.680 15.590 94.440 15.620 ;
        RECT 77.720 15.180 80.320 15.350 ;
        RECT 119.600 15.000 119.770 15.650 ;
        RECT 120.400 15.140 121.400 15.310 ;
        RECT 49.990 14.780 57.590 14.950 ;
        RECT 50.460 14.750 53.220 14.780 ;
        RECT 36.500 14.340 39.100 14.510 ;
        RECT 91.230 14.610 101.310 14.780 ;
        RECT 79.720 14.250 82.320 14.420 ;
        RECT 50.010 13.770 60.090 13.940 ;
        RECT 38.500 13.410 41.100 13.580 ;
        RECT 38.500 12.760 38.670 13.410 ;
        RECT 39.300 12.900 40.300 13.070 ;
        RECT 38.480 10.960 38.680 12.760 ;
        RECT 38.500 7.770 38.670 10.960 ;
        RECT 39.070 8.450 39.240 12.730 ;
        RECT 40.360 8.450 40.530 12.730 ;
        RECT 39.300 8.110 40.300 8.280 ;
        RECT 40.930 7.770 41.100 13.410 ;
        RECT 50.010 11.370 50.180 13.770 ;
        RECT 50.810 13.260 59.290 13.430 ;
        RECT 50.580 12.050 50.750 13.090 ;
        RECT 59.350 12.050 59.520 13.090 ;
        RECT 50.810 11.710 59.290 11.880 ;
        RECT 59.920 11.370 60.090 13.770 ;
        RECT 79.720 13.600 79.890 14.250 ;
        RECT 80.520 13.740 81.520 13.910 ;
        RECT 79.700 11.800 79.900 13.600 ;
        RECT 50.010 11.200 60.090 11.370 ;
        RECT 50.460 11.170 53.220 11.200 ;
        RECT 38.500 7.600 41.100 7.770 ;
        RECT 50.020 10.190 63.620 10.360 ;
        RECT 50.020 7.790 50.190 10.190 ;
        RECT 50.820 9.680 62.820 9.850 ;
        RECT 50.590 8.470 50.760 9.510 ;
        RECT 62.880 8.470 63.050 9.510 ;
        RECT 50.820 8.130 62.820 8.300 ;
        RECT 60.380 7.790 63.130 7.810 ;
        RECT 63.450 7.790 63.620 10.190 ;
        RECT 79.720 8.610 79.890 11.800 ;
        RECT 80.290 9.290 80.460 13.570 ;
        RECT 81.580 9.290 81.750 13.570 ;
        RECT 80.520 8.950 81.520 9.120 ;
        RECT 82.150 8.610 82.320 14.250 ;
        RECT 91.230 12.210 91.400 14.610 ;
        RECT 92.030 14.100 100.510 14.270 ;
        RECT 91.800 12.890 91.970 13.930 ;
        RECT 100.570 12.890 100.740 13.930 ;
        RECT 92.030 12.550 100.510 12.720 ;
        RECT 101.140 12.210 101.310 14.610 ;
        RECT 119.580 13.200 119.780 15.000 ;
        RECT 91.230 12.040 101.310 12.210 ;
        RECT 91.680 12.010 94.440 12.040 ;
        RECT 79.720 8.440 82.320 8.610 ;
        RECT 91.240 11.030 104.840 11.200 ;
        RECT 91.240 8.630 91.410 11.030 ;
        RECT 92.040 10.520 104.040 10.690 ;
        RECT 91.810 9.310 91.980 10.350 ;
        RECT 104.100 9.310 104.270 10.350 ;
        RECT 92.040 8.970 104.040 9.140 ;
        RECT 101.600 8.630 104.350 8.650 ;
        RECT 104.670 8.630 104.840 11.030 ;
        RECT 119.600 10.010 119.770 13.200 ;
        RECT 120.170 10.690 120.340 14.970 ;
        RECT 121.460 10.690 121.630 14.970 ;
        RECT 120.400 10.350 121.400 10.520 ;
        RECT 122.030 10.010 122.200 15.650 ;
        RECT 131.110 13.610 131.280 16.010 ;
        RECT 131.910 15.500 140.390 15.670 ;
        RECT 131.680 14.290 131.850 15.330 ;
        RECT 140.450 14.290 140.620 15.330 ;
        RECT 131.910 13.950 140.390 14.120 ;
        RECT 141.020 13.610 141.190 16.010 ;
        RECT 131.110 13.440 141.190 13.610 ;
        RECT 131.560 13.410 134.320 13.440 ;
        RECT 119.600 9.840 122.200 10.010 ;
        RECT 131.120 12.430 144.720 12.600 ;
        RECT 131.120 10.030 131.290 12.430 ;
        RECT 131.920 11.920 143.920 12.090 ;
        RECT 131.690 10.710 131.860 11.750 ;
        RECT 143.980 10.710 144.150 11.750 ;
        RECT 131.920 10.370 143.920 10.540 ;
        RECT 141.480 10.030 144.230 10.050 ;
        RECT 144.550 10.030 144.720 12.430 ;
        RECT 131.120 9.860 144.720 10.030 ;
        RECT 141.480 9.850 144.230 9.860 ;
        RECT 91.240 8.460 104.840 8.630 ;
        RECT 101.600 8.450 104.350 8.460 ;
        RECT 50.020 7.620 63.620 7.790 ;
        RECT 60.380 7.610 63.130 7.620 ;
      LAYER met1 ;
        RECT 103.270 209.840 103.590 209.900 ;
        RECT 117.070 209.840 117.390 209.900 ;
        RECT 103.270 209.700 117.390 209.840 ;
        RECT 103.270 209.640 103.590 209.700 ;
        RECT 117.070 209.640 117.390 209.700 ;
        RECT 22.700 209.020 157.820 209.500 ;
        RECT 61.885 208.635 62.175 208.865 ;
        RECT 79.825 208.820 80.115 208.865 ;
        RECT 117.070 208.820 117.390 208.880 ;
        RECT 152.505 208.820 152.795 208.865 ;
        RECT 79.825 208.680 89.700 208.820 ;
        RECT 79.825 208.635 80.115 208.680 ;
        RECT 61.960 208.480 62.100 208.635 ;
        RECT 70.610 208.525 70.930 208.540 ;
        RECT 49.080 208.340 62.100 208.480 ;
        RECT 48.070 208.140 48.390 208.200 ;
        RECT 49.080 208.185 49.220 208.340 ;
        RECT 70.545 208.295 70.930 208.525 ;
        RECT 71.545 208.480 71.835 208.525 ;
        RECT 71.545 208.340 72.680 208.480 ;
        RECT 71.545 208.295 71.835 208.340 ;
        RECT 70.610 208.280 70.930 208.295 ;
        RECT 49.005 208.140 49.295 208.185 ;
        RECT 48.070 208.000 49.295 208.140 ;
        RECT 48.070 207.940 48.390 208.000 ;
        RECT 49.005 207.955 49.295 208.000 ;
        RECT 51.765 207.955 52.055 208.185 ;
        RECT 52.685 208.140 52.975 208.185 ;
        RECT 54.985 208.140 55.275 208.185 ;
        RECT 57.285 208.140 57.575 208.185 ;
        RECT 52.685 208.000 54.280 208.140 ;
        RECT 52.685 207.955 52.975 208.000 ;
        RECT 51.840 207.800 51.980 207.955 ;
        RECT 51.840 207.660 53.360 207.800 ;
        RECT 51.750 207.460 52.070 207.520 ;
        RECT 53.220 207.505 53.360 207.660 ;
        RECT 50.460 207.320 52.070 207.460 ;
        RECT 50.460 207.165 50.600 207.320 ;
        RECT 51.750 207.260 52.070 207.320 ;
        RECT 53.145 207.275 53.435 207.505 ;
        RECT 54.140 207.460 54.280 208.000 ;
        RECT 54.985 208.000 57.575 208.140 ;
        RECT 54.985 207.955 55.275 208.000 ;
        RECT 57.285 207.955 57.575 208.000 ;
        RECT 57.730 208.140 58.050 208.200 ;
        RECT 62.805 208.140 63.095 208.185 ;
        RECT 57.730 208.000 63.095 208.140 ;
        RECT 57.730 207.940 58.050 208.000 ;
        RECT 62.805 207.955 63.095 208.000 ;
        RECT 63.710 208.140 64.030 208.200 ;
        RECT 64.185 208.140 64.475 208.185 ;
        RECT 63.710 208.000 64.475 208.140 ;
        RECT 63.710 207.940 64.030 208.000 ;
        RECT 64.185 207.955 64.475 208.000 ;
        RECT 71.070 208.140 71.390 208.200 ;
        RECT 72.005 208.140 72.295 208.185 ;
        RECT 71.070 208.000 72.295 208.140 ;
        RECT 71.070 207.940 71.390 208.000 ;
        RECT 72.005 207.955 72.295 208.000 ;
        RECT 54.510 207.600 54.830 207.860 ;
        RECT 60.030 207.600 60.350 207.860 ;
        RECT 72.540 207.800 72.680 208.340 ;
        RECT 78.430 208.140 78.750 208.200 ;
        RECT 78.905 208.140 79.195 208.185 ;
        RECT 78.430 208.000 79.195 208.140 ;
        RECT 78.430 207.940 78.750 208.000 ;
        RECT 78.905 207.955 79.195 208.000 ;
        RECT 80.270 208.140 80.590 208.200 ;
        RECT 80.745 208.140 81.035 208.185 ;
        RECT 80.270 208.000 81.035 208.140 ;
        RECT 80.270 207.940 80.590 208.000 ;
        RECT 80.745 207.955 81.035 208.000 ;
        RECT 81.665 208.140 81.955 208.185 ;
        RECT 82.585 208.140 82.875 208.185 ;
        RECT 81.665 208.000 82.875 208.140 ;
        RECT 81.665 207.955 81.955 208.000 ;
        RECT 82.585 207.955 82.875 208.000 ;
        RECT 63.800 207.660 72.680 207.800 ;
        RECT 63.800 207.520 63.940 207.660 ;
        RECT 63.710 207.460 64.030 207.520 ;
        RECT 54.140 207.320 64.030 207.460 ;
        RECT 63.710 207.260 64.030 207.320 ;
        RECT 65.105 207.460 65.395 207.505 ;
        RECT 76.130 207.460 76.450 207.520 ;
        RECT 65.105 207.320 76.450 207.460 ;
        RECT 80.820 207.460 80.960 207.955 ;
        RECT 83.490 207.800 83.810 207.860 ;
        RECT 89.560 207.845 89.700 208.680 ;
        RECT 109.340 208.680 112.240 208.820 ;
        RECT 100.510 208.480 100.830 208.540 ;
        RECT 109.340 208.525 109.480 208.680 ;
        RECT 100.510 208.340 103.960 208.480 ;
        RECT 100.510 208.280 100.830 208.340 ;
        RECT 90.850 207.940 91.170 208.200 ;
        RECT 91.325 207.955 91.615 208.185 ;
        RECT 93.150 208.140 93.470 208.200 ;
        RECT 93.625 208.140 93.915 208.185 ;
        RECT 93.150 208.000 93.915 208.140 ;
        RECT 85.345 207.800 85.635 207.845 ;
        RECT 83.490 207.660 85.635 207.800 ;
        RECT 83.490 207.600 83.810 207.660 ;
        RECT 85.345 207.615 85.635 207.660 ;
        RECT 89.485 207.800 89.775 207.845 ;
        RECT 90.940 207.800 91.080 207.940 ;
        RECT 89.485 207.660 91.080 207.800 ;
        RECT 91.400 207.800 91.540 207.955 ;
        RECT 93.150 207.940 93.470 208.000 ;
        RECT 93.625 207.955 93.915 208.000 ;
        RECT 103.270 207.940 103.590 208.200 ;
        RECT 103.820 208.185 103.960 208.340 ;
        RECT 109.265 208.295 109.555 208.525 ;
        RECT 109.710 208.480 110.030 208.540 ;
        RECT 111.565 208.480 111.855 208.525 ;
        RECT 109.710 208.340 111.855 208.480 ;
        RECT 112.100 208.480 112.240 208.680 ;
        RECT 117.070 208.680 152.795 208.820 ;
        RECT 117.070 208.620 117.390 208.680 ;
        RECT 152.505 208.635 152.795 208.680 ;
        RECT 114.325 208.480 114.615 208.525 ;
        RECT 115.690 208.480 116.010 208.540 ;
        RECT 112.100 208.340 116.010 208.480 ;
        RECT 109.710 208.280 110.030 208.340 ;
        RECT 111.565 208.295 111.855 208.340 ;
        RECT 114.325 208.295 114.615 208.340 ;
        RECT 115.690 208.280 116.010 208.340 ;
        RECT 116.610 208.480 116.930 208.540 ;
        RECT 122.145 208.480 122.435 208.525 ;
        RECT 116.610 208.340 122.435 208.480 ;
        RECT 116.610 208.280 116.930 208.340 ;
        RECT 122.145 208.295 122.435 208.340 ;
        RECT 123.985 208.480 124.275 208.525 ;
        RECT 124.430 208.480 124.750 208.540 ;
        RECT 123.985 208.340 124.750 208.480 ;
        RECT 123.985 208.295 124.275 208.340 ;
        RECT 124.430 208.280 124.750 208.340 ;
        RECT 130.410 208.480 130.730 208.540 ;
        RECT 131.345 208.480 131.635 208.525 ;
        RECT 130.410 208.340 131.635 208.480 ;
        RECT 130.410 208.280 130.730 208.340 ;
        RECT 131.345 208.295 131.635 208.340 ;
        RECT 103.745 207.955 104.035 208.185 ;
        RECT 108.330 207.940 108.650 208.200 ;
        RECT 108.790 207.940 109.110 208.200 ;
        RECT 110.170 207.940 110.490 208.200 ;
        RECT 113.405 207.955 113.695 208.185 ;
        RECT 113.850 208.140 114.170 208.200 ;
        RECT 114.785 208.140 115.075 208.185 ;
        RECT 113.850 208.000 115.075 208.140 ;
        RECT 91.400 207.660 100.740 207.800 ;
        RECT 89.485 207.615 89.775 207.660 ;
        RECT 100.600 207.505 100.740 207.660 ;
        RECT 101.905 207.615 102.195 207.845 ;
        RECT 113.480 207.800 113.620 207.955 ;
        RECT 113.850 207.940 114.170 208.000 ;
        RECT 114.785 207.955 115.075 208.000 ;
        RECT 115.230 207.940 115.550 208.200 ;
        RECT 134.550 207.940 134.870 208.200 ;
        RECT 137.310 208.140 137.630 208.200 ;
        RECT 139.165 208.140 139.455 208.185 ;
        RECT 137.310 208.000 139.455 208.140 ;
        RECT 137.310 207.940 137.630 208.000 ;
        RECT 139.165 207.955 139.455 208.000 ;
        RECT 152.030 208.140 152.350 208.200 ;
        RECT 153.425 208.140 153.715 208.185 ;
        RECT 152.030 208.000 153.715 208.140 ;
        RECT 152.030 207.940 152.350 208.000 ;
        RECT 153.425 207.955 153.715 208.000 ;
        RECT 117.545 207.800 117.835 207.845 ;
        RECT 113.480 207.660 117.835 207.800 ;
        RECT 117.545 207.615 117.835 207.660 ;
        RECT 120.765 207.800 121.055 207.845 ;
        RECT 122.130 207.800 122.450 207.860 ;
        RECT 120.765 207.660 122.450 207.800 ;
        RECT 120.765 207.615 121.055 207.660 ;
        RECT 90.500 207.460 90.790 207.505 ;
        RECT 80.820 207.320 90.790 207.460 ;
        RECT 65.105 207.275 65.395 207.320 ;
        RECT 76.130 207.260 76.450 207.320 ;
        RECT 90.500 207.275 90.790 207.320 ;
        RECT 100.525 207.275 100.815 207.505 ;
        RECT 50.385 206.935 50.675 207.165 ;
        RECT 51.290 206.920 51.610 207.180 ;
        RECT 52.225 207.120 52.515 207.165 ;
        RECT 54.510 207.120 54.830 207.180 ;
        RECT 52.225 206.980 54.830 207.120 ;
        RECT 52.225 206.935 52.515 206.980 ;
        RECT 54.510 206.920 54.830 206.980 ;
        RECT 68.310 207.120 68.630 207.180 ;
        RECT 69.705 207.120 69.995 207.165 ;
        RECT 68.310 206.980 69.995 207.120 ;
        RECT 68.310 206.920 68.630 206.980 ;
        RECT 69.705 206.935 69.995 206.980 ;
        RECT 70.625 207.120 70.915 207.165 ;
        RECT 71.530 207.120 71.850 207.180 ;
        RECT 70.625 206.980 71.850 207.120 ;
        RECT 70.625 206.935 70.915 206.980 ;
        RECT 71.530 206.920 71.850 206.980 ;
        RECT 72.925 207.120 73.215 207.165 ;
        RECT 75.210 207.120 75.530 207.180 ;
        RECT 72.925 206.980 75.530 207.120 ;
        RECT 72.925 206.935 73.215 206.980 ;
        RECT 75.210 206.920 75.530 206.980 ;
        RECT 78.430 207.120 78.750 207.180 ;
        RECT 81.205 207.120 81.495 207.165 ;
        RECT 78.430 206.980 81.495 207.120 ;
        RECT 78.430 206.920 78.750 206.980 ;
        RECT 81.205 206.935 81.495 206.980 ;
        RECT 88.090 206.920 88.410 207.180 ;
        RECT 89.930 206.920 90.250 207.180 ;
        RECT 93.610 207.120 93.930 207.180 ;
        RECT 94.545 207.120 94.835 207.165 ;
        RECT 101.980 207.120 102.120 207.615 ;
        RECT 122.130 207.600 122.450 207.660 ;
        RECT 137.770 207.800 138.090 207.860 ;
        RECT 140.545 207.800 140.835 207.845 ;
        RECT 137.770 207.660 140.835 207.800 ;
        RECT 137.770 207.600 138.090 207.660 ;
        RECT 140.545 207.615 140.835 207.660 ;
        RECT 117.070 207.460 117.390 207.520 ;
        RECT 123.065 207.460 123.355 207.505 ;
        RECT 115.780 207.320 116.840 207.460 ;
        RECT 93.610 206.980 102.120 207.120 ;
        RECT 102.825 207.120 103.115 207.165 ;
        RECT 103.730 207.120 104.050 207.180 ;
        RECT 104.665 207.120 104.955 207.165 ;
        RECT 102.825 206.980 104.955 207.120 ;
        RECT 93.610 206.920 93.930 206.980 ;
        RECT 94.545 206.935 94.835 206.980 ;
        RECT 102.825 206.935 103.115 206.980 ;
        RECT 103.730 206.920 104.050 206.980 ;
        RECT 104.665 206.935 104.955 206.980 ;
        RECT 107.425 207.120 107.715 207.165 ;
        RECT 107.870 207.120 108.190 207.180 ;
        RECT 107.425 206.980 108.190 207.120 ;
        RECT 107.425 206.935 107.715 206.980 ;
        RECT 107.870 206.920 108.190 206.980 ;
        RECT 108.790 207.120 109.110 207.180 ;
        RECT 111.105 207.120 111.395 207.165 ;
        RECT 108.790 206.980 111.395 207.120 ;
        RECT 108.790 206.920 109.110 206.980 ;
        RECT 111.105 206.935 111.395 206.980 ;
        RECT 113.390 207.120 113.710 207.180 ;
        RECT 115.780 207.120 115.920 207.320 ;
        RECT 113.390 206.980 115.920 207.120 ;
        RECT 113.390 206.920 113.710 206.980 ;
        RECT 116.150 206.920 116.470 207.180 ;
        RECT 116.700 207.120 116.840 207.320 ;
        RECT 117.070 207.320 123.355 207.460 ;
        RECT 117.070 207.260 117.390 207.320 ;
        RECT 123.065 207.275 123.355 207.320 ;
        RECT 121.685 207.120 121.975 207.165 ;
        RECT 116.700 206.980 121.975 207.120 ;
        RECT 121.685 206.935 121.975 206.980 ;
        RECT 130.885 207.120 131.175 207.165 ;
        RECT 131.790 207.120 132.110 207.180 ;
        RECT 130.885 206.980 132.110 207.120 ;
        RECT 130.885 206.935 131.175 206.980 ;
        RECT 131.790 206.920 132.110 206.980 ;
        RECT 132.710 207.120 133.030 207.180 ;
        RECT 133.645 207.120 133.935 207.165 ;
        RECT 132.710 206.980 133.935 207.120 ;
        RECT 132.710 206.920 133.030 206.980 ;
        RECT 133.645 206.935 133.935 206.980 ;
        RECT 22.700 206.300 157.020 206.780 ;
        RECT 60.030 205.900 60.350 206.160 ;
        RECT 75.685 206.100 75.975 206.145 ;
        RECT 80.270 206.100 80.590 206.160 ;
        RECT 75.685 205.960 80.590 206.100 ;
        RECT 75.685 205.915 75.975 205.960 ;
        RECT 80.270 205.900 80.590 205.960 ;
        RECT 83.490 205.900 83.810 206.160 ;
        RECT 31.050 205.760 31.340 205.805 ;
        RECT 32.620 205.760 32.910 205.805 ;
        RECT 34.720 205.760 35.010 205.805 ;
        RECT 31.050 205.620 35.010 205.760 ;
        RECT 31.050 205.575 31.340 205.620 ;
        RECT 32.620 205.575 32.910 205.620 ;
        RECT 34.720 205.575 35.010 205.620 ;
        RECT 36.610 205.760 36.900 205.805 ;
        RECT 38.710 205.760 39.000 205.805 ;
        RECT 40.280 205.760 40.570 205.805 ;
        RECT 36.610 205.620 40.570 205.760 ;
        RECT 36.610 205.575 36.900 205.620 ;
        RECT 38.710 205.575 39.000 205.620 ;
        RECT 40.280 205.575 40.570 205.620 ;
        RECT 41.630 205.760 41.950 205.820 ;
        RECT 43.025 205.760 43.315 205.805 ;
        RECT 41.630 205.620 43.315 205.760 ;
        RECT 41.630 205.560 41.950 205.620 ;
        RECT 43.025 205.575 43.315 205.620 ;
        RECT 44.430 205.760 44.720 205.805 ;
        RECT 46.530 205.760 46.820 205.805 ;
        RECT 48.100 205.760 48.390 205.805 ;
        RECT 44.430 205.620 48.390 205.760 ;
        RECT 44.430 205.575 44.720 205.620 ;
        RECT 46.530 205.575 46.820 205.620 ;
        RECT 48.100 205.575 48.390 205.620 ;
        RECT 53.630 205.760 53.920 205.805 ;
        RECT 55.730 205.760 56.020 205.805 ;
        RECT 57.300 205.760 57.590 205.805 ;
        RECT 53.630 205.620 57.590 205.760 ;
        RECT 53.630 205.575 53.920 205.620 ;
        RECT 55.730 205.575 56.020 205.620 ;
        RECT 57.300 205.575 57.590 205.620 ;
        RECT 67.890 205.760 68.180 205.805 ;
        RECT 69.990 205.760 70.280 205.805 ;
        RECT 71.560 205.760 71.850 205.805 ;
        RECT 67.890 205.620 71.850 205.760 ;
        RECT 67.890 205.575 68.180 205.620 ;
        RECT 69.990 205.575 70.280 205.620 ;
        RECT 71.560 205.575 71.850 205.620 ;
        RECT 77.090 205.760 77.380 205.805 ;
        RECT 79.190 205.760 79.480 205.805 ;
        RECT 80.760 205.760 81.050 205.805 ;
        RECT 77.090 205.620 81.050 205.760 ;
        RECT 77.090 205.575 77.380 205.620 ;
        RECT 79.190 205.575 79.480 205.620 ;
        RECT 80.760 205.575 81.050 205.620 ;
        RECT 92.230 205.760 92.520 205.805 ;
        RECT 93.800 205.760 94.090 205.805 ;
        RECT 95.900 205.760 96.190 205.805 ;
        RECT 92.230 205.620 96.190 205.760 ;
        RECT 92.230 205.575 92.520 205.620 ;
        RECT 93.800 205.575 94.090 205.620 ;
        RECT 95.900 205.575 96.190 205.620 ;
        RECT 100.050 205.560 100.370 205.820 ;
        RECT 102.810 205.760 103.100 205.805 ;
        RECT 104.380 205.760 104.670 205.805 ;
        RECT 106.480 205.760 106.770 205.805 ;
        RECT 102.810 205.620 106.770 205.760 ;
        RECT 102.810 205.575 103.100 205.620 ;
        RECT 104.380 205.575 104.670 205.620 ;
        RECT 106.480 205.575 106.770 205.620 ;
        RECT 109.265 205.760 109.555 205.805 ;
        RECT 110.170 205.760 110.490 205.820 ;
        RECT 109.265 205.620 110.490 205.760 ;
        RECT 109.265 205.575 109.555 205.620 ;
        RECT 110.170 205.560 110.490 205.620 ;
        RECT 114.810 205.760 115.100 205.805 ;
        RECT 116.910 205.760 117.200 205.805 ;
        RECT 118.480 205.760 118.770 205.805 ;
        RECT 114.810 205.620 118.770 205.760 ;
        RECT 114.810 205.575 115.100 205.620 ;
        RECT 116.910 205.575 117.200 205.620 ;
        RECT 118.480 205.575 118.770 205.620 ;
        RECT 121.225 205.575 121.515 205.805 ;
        RECT 125.825 205.760 126.115 205.805 ;
        RECT 127.650 205.760 127.970 205.820 ;
        RECT 125.825 205.620 127.970 205.760 ;
        RECT 125.825 205.575 126.115 205.620 ;
        RECT 30.615 205.420 30.905 205.465 ;
        RECT 33.135 205.420 33.425 205.465 ;
        RECT 34.325 205.420 34.615 205.465 ;
        RECT 30.615 205.280 34.615 205.420 ;
        RECT 30.615 205.235 30.905 205.280 ;
        RECT 33.135 205.235 33.425 205.280 ;
        RECT 34.325 205.235 34.615 205.280 ;
        RECT 37.005 205.420 37.295 205.465 ;
        RECT 38.195 205.420 38.485 205.465 ;
        RECT 40.715 205.420 41.005 205.465 ;
        RECT 37.005 205.280 41.005 205.420 ;
        RECT 37.005 205.235 37.295 205.280 ;
        RECT 38.195 205.235 38.485 205.280 ;
        RECT 40.715 205.235 41.005 205.280 ;
        RECT 44.825 205.420 45.115 205.465 ;
        RECT 46.015 205.420 46.305 205.465 ;
        RECT 48.535 205.420 48.825 205.465 ;
        RECT 44.825 205.280 48.825 205.420 ;
        RECT 44.825 205.235 45.115 205.280 ;
        RECT 46.015 205.235 46.305 205.280 ;
        RECT 48.535 205.235 48.825 205.280 ;
        RECT 52.210 205.420 52.530 205.480 ;
        RECT 53.145 205.420 53.435 205.465 ;
        RECT 52.210 205.280 53.435 205.420 ;
        RECT 52.210 205.220 52.530 205.280 ;
        RECT 53.145 205.235 53.435 205.280 ;
        RECT 54.025 205.420 54.315 205.465 ;
        RECT 55.215 205.420 55.505 205.465 ;
        RECT 57.735 205.420 58.025 205.465 ;
        RECT 54.025 205.280 58.025 205.420 ;
        RECT 54.025 205.235 54.315 205.280 ;
        RECT 55.215 205.235 55.505 205.280 ;
        RECT 57.735 205.235 58.025 205.280 ;
        RECT 62.330 205.420 62.650 205.480 ;
        RECT 67.405 205.420 67.695 205.465 ;
        RECT 62.330 205.280 67.695 205.420 ;
        RECT 62.330 205.220 62.650 205.280 ;
        RECT 67.405 205.235 67.695 205.280 ;
        RECT 68.285 205.420 68.575 205.465 ;
        RECT 69.475 205.420 69.765 205.465 ;
        RECT 71.995 205.420 72.285 205.465 ;
        RECT 76.590 205.420 76.910 205.480 ;
        RECT 68.285 205.280 72.285 205.420 ;
        RECT 68.285 205.235 68.575 205.280 ;
        RECT 69.475 205.235 69.765 205.280 ;
        RECT 71.995 205.235 72.285 205.280 ;
        RECT 74.840 205.280 76.910 205.420 ;
        RECT 35.205 205.080 35.495 205.125 ;
        RECT 36.110 205.080 36.430 205.140 ;
        RECT 35.205 204.940 36.430 205.080 ;
        RECT 35.205 204.895 35.495 204.940 ;
        RECT 36.110 204.880 36.430 204.940 ;
        RECT 43.945 205.080 44.235 205.125 ;
        RECT 47.610 205.080 47.930 205.140 ;
        RECT 52.300 205.080 52.440 205.220 ;
        RECT 54.510 205.125 54.830 205.140 ;
        RECT 43.945 204.940 52.440 205.080 ;
        RECT 43.945 204.895 44.235 204.940 ;
        RECT 47.610 204.880 47.930 204.940 ;
        RECT 52.685 204.895 52.975 205.125 ;
        RECT 54.480 205.080 54.830 205.125 ;
        RECT 54.315 204.940 54.830 205.080 ;
        RECT 54.480 204.895 54.830 204.940 ;
        RECT 33.810 204.785 34.130 204.800 ;
        RECT 33.810 204.555 34.160 204.785 ;
        RECT 37.460 204.555 37.750 204.785 ;
        RECT 41.630 204.740 41.950 204.800 ;
        RECT 45.170 204.740 45.460 204.785 ;
        RECT 41.630 204.600 45.460 204.740 ;
        RECT 33.810 204.540 34.130 204.555 ;
        RECT 28.305 204.400 28.595 204.445 ;
        RECT 34.730 204.400 35.050 204.460 ;
        RECT 28.305 204.260 35.050 204.400 ;
        RECT 28.305 204.215 28.595 204.260 ;
        RECT 34.730 204.200 35.050 204.260 ;
        RECT 37.030 204.400 37.350 204.460 ;
        RECT 37.580 204.400 37.720 204.555 ;
        RECT 41.630 204.540 41.950 204.600 ;
        RECT 45.170 204.555 45.460 204.600 ;
        RECT 48.990 204.740 49.310 204.800 ;
        RECT 52.760 204.740 52.900 204.895 ;
        RECT 54.510 204.880 54.830 204.895 ;
        RECT 61.410 205.080 61.730 205.140 ;
        RECT 61.885 205.080 62.175 205.125 ;
        RECT 61.410 204.940 62.175 205.080 ;
        RECT 61.410 204.880 61.730 204.940 ;
        RECT 61.885 204.895 62.175 204.940 ;
        RECT 62.805 204.895 63.095 205.125 ;
        RECT 48.990 204.600 52.900 204.740 ;
        RECT 62.880 204.740 63.020 204.895 ;
        RECT 64.170 204.880 64.490 205.140 ;
        RECT 65.550 204.880 65.870 205.140 ;
        RECT 66.025 205.080 66.315 205.125 ;
        RECT 66.930 205.080 67.250 205.140 ;
        RECT 66.025 204.940 67.250 205.080 ;
        RECT 67.480 205.080 67.620 205.235 ;
        RECT 74.840 205.080 74.980 205.280 ;
        RECT 76.590 205.220 76.910 205.280 ;
        RECT 77.485 205.420 77.775 205.465 ;
        RECT 78.675 205.420 78.965 205.465 ;
        RECT 81.195 205.420 81.485 205.465 ;
        RECT 77.485 205.280 81.485 205.420 ;
        RECT 77.485 205.235 77.775 205.280 ;
        RECT 78.675 205.235 78.965 205.280 ;
        RECT 81.195 205.235 81.485 205.280 ;
        RECT 91.795 205.420 92.085 205.465 ;
        RECT 94.315 205.420 94.605 205.465 ;
        RECT 95.505 205.420 95.795 205.465 ;
        RECT 91.795 205.280 95.795 205.420 ;
        RECT 91.795 205.235 92.085 205.280 ;
        RECT 94.315 205.235 94.605 205.280 ;
        RECT 95.505 205.235 95.795 205.280 ;
        RECT 102.375 205.420 102.665 205.465 ;
        RECT 104.895 205.420 105.185 205.465 ;
        RECT 106.085 205.420 106.375 205.465 ;
        RECT 102.375 205.280 106.375 205.420 ;
        RECT 102.375 205.235 102.665 205.280 ;
        RECT 104.895 205.235 105.185 205.280 ;
        RECT 106.085 205.235 106.375 205.280 ;
        RECT 115.205 205.420 115.495 205.465 ;
        RECT 116.395 205.420 116.685 205.465 ;
        RECT 118.915 205.420 119.205 205.465 ;
        RECT 115.205 205.280 119.205 205.420 ;
        RECT 121.300 205.420 121.440 205.575 ;
        RECT 127.650 205.560 127.970 205.620 ;
        RECT 129.505 205.760 129.795 205.805 ;
        RECT 131.830 205.760 132.120 205.805 ;
        RECT 133.930 205.760 134.220 205.805 ;
        RECT 135.500 205.760 135.790 205.805 ;
        RECT 129.505 205.620 130.410 205.760 ;
        RECT 129.505 205.575 129.795 205.620 ;
        RECT 122.130 205.420 122.450 205.480 ;
        RECT 121.300 205.280 122.450 205.420 ;
        RECT 115.205 205.235 115.495 205.280 ;
        RECT 116.395 205.235 116.685 205.280 ;
        RECT 118.915 205.235 119.205 205.280 ;
        RECT 122.130 205.220 122.450 205.280 ;
        RECT 124.445 205.420 124.735 205.465 ;
        RECT 129.030 205.420 129.350 205.480 ;
        RECT 124.445 205.280 129.350 205.420 ;
        RECT 124.445 205.235 124.735 205.280 ;
        RECT 129.030 205.220 129.350 205.280 ;
        RECT 67.480 204.940 74.980 205.080 ;
        RECT 66.025 204.895 66.315 204.940 ;
        RECT 66.930 204.880 67.250 204.940 ;
        RECT 75.210 204.880 75.530 205.140 ;
        RECT 76.130 204.880 76.450 205.140 ;
        RECT 85.345 205.080 85.635 205.125 ;
        RECT 85.790 205.080 86.110 205.140 ;
        RECT 85.345 204.940 86.110 205.080 ;
        RECT 85.345 204.895 85.635 204.940 ;
        RECT 85.790 204.880 86.110 204.940 ;
        RECT 88.550 204.880 88.870 205.140 ;
        RECT 96.385 204.895 96.675 205.125 ;
        RECT 96.830 205.080 97.150 205.140 ;
        RECT 97.765 205.080 98.055 205.125 ;
        RECT 96.830 204.940 98.055 205.080 ;
        RECT 68.630 204.740 68.920 204.785 ;
        RECT 62.880 204.600 65.320 204.740 ;
        RECT 48.990 204.540 49.310 204.600 ;
        RECT 37.030 204.260 37.720 204.400 ;
        RECT 50.370 204.400 50.690 204.460 ;
        RECT 50.845 204.400 51.135 204.445 ;
        RECT 50.370 204.260 51.135 204.400 ;
        RECT 37.030 204.200 37.350 204.260 ;
        RECT 50.370 204.200 50.690 204.260 ;
        RECT 50.845 204.215 51.135 204.260 ;
        RECT 51.750 204.200 52.070 204.460 ;
        RECT 62.790 204.200 63.110 204.460 ;
        RECT 63.250 204.200 63.570 204.460 ;
        RECT 65.180 204.445 65.320 204.600 ;
        RECT 67.020 204.600 68.920 204.740 ;
        RECT 65.105 204.400 65.395 204.445 ;
        RECT 66.470 204.400 66.790 204.460 ;
        RECT 67.020 204.445 67.160 204.600 ;
        RECT 68.630 204.555 68.920 204.600 ;
        RECT 77.050 204.740 77.370 204.800 ;
        RECT 77.830 204.740 78.120 204.785 ;
        RECT 89.930 204.740 90.250 204.800 ;
        RECT 77.050 204.600 78.120 204.740 ;
        RECT 77.050 204.540 77.370 204.600 ;
        RECT 77.830 204.555 78.120 204.600 ;
        RECT 86.340 204.600 90.250 204.740 ;
        RECT 65.105 204.260 66.790 204.400 ;
        RECT 65.105 204.215 65.395 204.260 ;
        RECT 66.470 204.200 66.790 204.260 ;
        RECT 66.945 204.215 67.235 204.445 ;
        RECT 72.910 204.400 73.230 204.460 ;
        RECT 74.290 204.400 74.610 204.460 ;
        RECT 72.910 204.260 74.610 204.400 ;
        RECT 72.910 204.200 73.230 204.260 ;
        RECT 74.290 204.200 74.610 204.260 ;
        RECT 85.790 204.400 86.110 204.460 ;
        RECT 86.340 204.445 86.480 204.600 ;
        RECT 89.930 204.540 90.250 204.600 ;
        RECT 95.160 204.740 95.450 204.785 ;
        RECT 96.460 204.740 96.600 204.895 ;
        RECT 96.830 204.880 97.150 204.940 ;
        RECT 97.765 204.895 98.055 204.940 ;
        RECT 98.685 205.080 98.975 205.125 ;
        RECT 100.510 205.080 100.830 205.140 ;
        RECT 106.965 205.080 107.255 205.125 ;
        RECT 98.685 204.940 100.830 205.080 ;
        RECT 98.685 204.895 98.975 204.940 ;
        RECT 100.510 204.880 100.830 204.940 ;
        RECT 104.280 204.940 107.255 205.080 ;
        RECT 104.280 204.800 104.420 204.940 ;
        RECT 106.965 204.895 107.255 204.940 ;
        RECT 112.470 204.880 112.790 205.140 ;
        RECT 114.325 205.080 114.615 205.125 ;
        RECT 114.325 204.940 116.840 205.080 ;
        RECT 114.325 204.895 114.615 204.940 ;
        RECT 116.700 204.800 116.840 204.940 ;
        RECT 122.605 204.895 122.895 205.125 ;
        RECT 127.205 205.080 127.495 205.125 ;
        RECT 130.270 205.080 130.410 205.620 ;
        RECT 131.830 205.620 135.790 205.760 ;
        RECT 131.830 205.575 132.120 205.620 ;
        RECT 133.930 205.575 134.220 205.620 ;
        RECT 135.500 205.575 135.790 205.620 ;
        RECT 138.230 205.760 138.550 205.820 ;
        RECT 140.545 205.760 140.835 205.805 ;
        RECT 138.230 205.620 140.835 205.760 ;
        RECT 138.230 205.560 138.550 205.620 ;
        RECT 140.545 205.575 140.835 205.620 ;
        RECT 143.290 205.760 143.580 205.805 ;
        RECT 144.860 205.760 145.150 205.805 ;
        RECT 146.960 205.760 147.250 205.805 ;
        RECT 143.290 205.620 147.250 205.760 ;
        RECT 143.290 205.575 143.580 205.620 ;
        RECT 144.860 205.575 145.150 205.620 ;
        RECT 146.960 205.575 147.250 205.620 ;
        RECT 132.225 205.420 132.515 205.465 ;
        RECT 133.415 205.420 133.705 205.465 ;
        RECT 135.935 205.420 136.225 205.465 ;
        RECT 141.910 205.420 142.230 205.480 ;
        RECT 132.225 205.280 136.225 205.420 ;
        RECT 132.225 205.235 132.515 205.280 ;
        RECT 133.415 205.235 133.705 205.280 ;
        RECT 135.935 205.235 136.225 205.280 ;
        RECT 138.780 205.280 142.230 205.420 ;
        RECT 127.205 204.940 130.410 205.080 ;
        RECT 127.205 204.895 127.495 204.940 ;
        RECT 104.190 204.740 104.510 204.800 ;
        RECT 105.630 204.740 105.920 204.785 ;
        RECT 95.160 204.600 96.140 204.740 ;
        RECT 96.460 204.600 104.510 204.740 ;
        RECT 95.160 204.555 95.450 204.600 ;
        RECT 86.265 204.400 86.555 204.445 ;
        RECT 85.790 204.260 86.555 204.400 ;
        RECT 85.790 204.200 86.110 204.260 ;
        RECT 86.265 204.215 86.555 204.260 ;
        RECT 87.630 204.200 87.950 204.460 ;
        RECT 89.485 204.400 89.775 204.445 ;
        RECT 92.690 204.400 93.010 204.460 ;
        RECT 89.485 204.260 93.010 204.400 ;
        RECT 96.000 204.400 96.140 204.600 ;
        RECT 104.190 204.540 104.510 204.600 ;
        RECT 104.740 204.600 105.920 204.740 ;
        RECT 96.845 204.400 97.135 204.445 ;
        RECT 96.000 204.260 97.135 204.400 ;
        RECT 89.485 204.215 89.775 204.260 ;
        RECT 92.690 204.200 93.010 204.260 ;
        RECT 96.845 204.215 97.135 204.260 ;
        RECT 99.605 204.400 99.895 204.445 ;
        RECT 104.740 204.400 104.880 204.600 ;
        RECT 105.630 204.555 105.920 204.600 ;
        RECT 115.660 204.740 115.950 204.785 ;
        RECT 116.150 204.740 116.470 204.800 ;
        RECT 115.660 204.600 116.470 204.740 ;
        RECT 115.660 204.555 115.950 204.600 ;
        RECT 116.150 204.540 116.470 204.600 ;
        RECT 116.610 204.540 116.930 204.800 ;
        RECT 122.680 204.740 122.820 204.895 ;
        RECT 122.680 204.600 127.420 204.740 ;
        RECT 127.280 204.460 127.420 204.600 ;
        RECT 127.650 204.540 127.970 204.800 ;
        RECT 130.270 204.740 130.410 204.940 ;
        RECT 131.330 204.880 131.650 205.140 ;
        RECT 132.710 205.125 133.030 205.140 ;
        RECT 132.680 205.080 133.030 205.125 ;
        RECT 132.515 204.940 133.030 205.080 ;
        RECT 132.680 204.895 133.030 204.940 ;
        RECT 132.710 204.880 133.030 204.895 ;
        RECT 138.780 204.740 138.920 205.280 ;
        RECT 141.910 205.220 142.230 205.280 ;
        RECT 142.855 205.420 143.145 205.465 ;
        RECT 145.375 205.420 145.665 205.465 ;
        RECT 146.565 205.420 146.855 205.465 ;
        RECT 142.855 205.280 146.855 205.420 ;
        RECT 142.855 205.235 143.145 205.280 ;
        RECT 145.375 205.235 145.665 205.280 ;
        RECT 146.565 205.235 146.855 205.280 ;
        RECT 139.165 205.080 139.455 205.125 ;
        RECT 140.530 205.080 140.850 205.140 ;
        RECT 139.165 204.940 140.850 205.080 ;
        RECT 139.165 204.895 139.455 204.940 ;
        RECT 140.530 204.880 140.850 204.940 ;
        RECT 147.430 204.880 147.750 205.140 ;
        RECT 146.110 204.740 146.400 204.785 ;
        RECT 130.270 204.600 138.920 204.740 ;
        RECT 140.160 204.600 146.400 204.740 ;
        RECT 99.605 204.260 104.880 204.400 ;
        RECT 124.905 204.400 125.195 204.445 ;
        RECT 126.730 204.400 127.050 204.460 ;
        RECT 124.905 204.260 127.050 204.400 ;
        RECT 99.605 204.215 99.895 204.260 ;
        RECT 124.905 204.215 125.195 204.260 ;
        RECT 126.730 204.200 127.050 204.260 ;
        RECT 127.190 204.200 127.510 204.460 ;
        RECT 129.950 204.200 130.270 204.460 ;
        RECT 135.930 204.400 136.250 204.460 ;
        RECT 140.160 204.445 140.300 204.600 ;
        RECT 146.110 204.555 146.400 204.600 ;
        RECT 138.245 204.400 138.535 204.445 ;
        RECT 135.930 204.260 138.535 204.400 ;
        RECT 135.930 204.200 136.250 204.260 ;
        RECT 138.245 204.215 138.535 204.260 ;
        RECT 140.085 204.215 140.375 204.445 ;
        RECT 22.700 203.580 157.820 204.060 ;
        RECT 24.625 203.380 24.915 203.425 ;
        RECT 26.910 203.380 27.230 203.440 ;
        RECT 24.625 203.240 27.230 203.380 ;
        RECT 24.625 203.195 24.915 203.240 ;
        RECT 26.910 203.180 27.230 203.240 ;
        RECT 41.630 203.180 41.950 203.440 ;
        RECT 65.550 203.380 65.870 203.440 ;
        RECT 66.945 203.380 67.235 203.425 ;
        RECT 65.550 203.240 67.235 203.380 ;
        RECT 65.550 203.180 65.870 203.240 ;
        RECT 66.945 203.195 67.235 203.240 ;
        RECT 70.610 203.180 70.930 203.440 ;
        RECT 71.530 203.380 71.850 203.440 ;
        RECT 72.925 203.380 73.215 203.425 ;
        RECT 71.530 203.240 73.215 203.380 ;
        RECT 71.530 203.180 71.850 203.240 ;
        RECT 72.925 203.195 73.215 203.240 ;
        RECT 75.210 203.380 75.530 203.440 ;
        RECT 79.365 203.380 79.655 203.425 ;
        RECT 75.210 203.240 79.655 203.380 ;
        RECT 75.210 203.180 75.530 203.240 ;
        RECT 79.365 203.195 79.655 203.240 ;
        RECT 79.825 203.380 80.115 203.425 ;
        RECT 83.490 203.380 83.810 203.440 ;
        RECT 79.825 203.240 83.810 203.380 ;
        RECT 79.825 203.195 80.115 203.240 ;
        RECT 83.490 203.180 83.810 203.240 ;
        RECT 92.690 203.380 93.010 203.440 ;
        RECT 95.450 203.380 95.770 203.440 ;
        RECT 92.690 203.240 96.600 203.380 ;
        RECT 92.690 203.180 93.010 203.240 ;
        RECT 95.450 203.180 95.770 203.240 ;
        RECT 36.110 203.040 36.430 203.100 ;
        RECT 37.490 203.040 37.810 203.100 ;
        RECT 43.025 203.040 43.315 203.085 ;
        RECT 47.610 203.040 47.930 203.100 ;
        RECT 64.630 203.040 64.950 203.100 ;
        RECT 76.130 203.040 76.450 203.100 ;
        RECT 77.985 203.040 78.275 203.085 ;
        RECT 36.110 202.900 47.930 203.040 ;
        RECT 36.110 202.840 36.430 202.900 ;
        RECT 37.490 202.840 37.810 202.900 ;
        RECT 43.025 202.855 43.315 202.900 ;
        RECT 47.610 202.840 47.930 202.900 ;
        RECT 48.620 202.900 64.950 203.040 ;
        RECT 30.245 202.700 30.535 202.745 ;
        RECT 31.525 202.700 31.815 202.745 ;
        RECT 36.200 202.700 36.340 202.840 ;
        RECT 30.245 202.560 31.280 202.700 ;
        RECT 30.245 202.515 30.535 202.560 ;
        RECT 26.935 202.360 27.225 202.405 ;
        RECT 29.455 202.360 29.745 202.405 ;
        RECT 30.645 202.360 30.935 202.405 ;
        RECT 26.935 202.220 30.935 202.360 ;
        RECT 31.140 202.360 31.280 202.560 ;
        RECT 31.525 202.560 36.340 202.700 ;
        RECT 36.570 202.700 36.890 202.760 ;
        RECT 38.885 202.700 39.175 202.745 ;
        RECT 36.570 202.560 39.175 202.700 ;
        RECT 31.525 202.515 31.815 202.560 ;
        RECT 36.570 202.500 36.890 202.560 ;
        RECT 38.885 202.515 39.175 202.560 ;
        RECT 39.805 202.515 40.095 202.745 ;
        RECT 39.880 202.360 40.020 202.515 ;
        RECT 40.710 202.500 41.030 202.760 ;
        RECT 46.705 202.700 46.995 202.745 ;
        RECT 48.620 202.700 48.760 202.900 ;
        RECT 64.630 202.840 64.950 202.900 ;
        RECT 71.620 202.900 73.140 203.040 ;
        RECT 46.705 202.560 48.760 202.700 ;
        RECT 46.705 202.515 46.995 202.560 ;
        RECT 49.910 202.500 50.230 202.760 ;
        RECT 51.290 202.500 51.610 202.760 ;
        RECT 52.670 202.500 52.990 202.760 ;
        RECT 54.970 202.500 55.290 202.760 ;
        RECT 61.380 202.700 61.670 202.745 ;
        RECT 63.250 202.700 63.570 202.760 ;
        RECT 71.620 202.745 71.760 202.900 ;
        RECT 73.000 202.760 73.140 202.900 ;
        RECT 76.130 202.900 78.275 203.040 ;
        RECT 76.130 202.840 76.450 202.900 ;
        RECT 77.985 202.855 78.275 202.900 ;
        RECT 84.840 203.040 85.130 203.085 ;
        RECT 87.630 203.040 87.950 203.100 ;
        RECT 84.840 202.900 87.950 203.040 ;
        RECT 84.840 202.855 85.130 202.900 ;
        RECT 87.630 202.840 87.950 202.900 ;
        RECT 91.785 203.040 92.075 203.085 ;
        RECT 91.785 202.900 93.380 203.040 ;
        RECT 91.785 202.855 92.075 202.900 ;
        RECT 61.380 202.560 63.570 202.700 ;
        RECT 61.380 202.515 61.670 202.560 ;
        RECT 63.250 202.500 63.570 202.560 ;
        RECT 71.545 202.515 71.835 202.745 ;
        RECT 72.465 202.515 72.755 202.745 ;
        RECT 48.990 202.360 49.310 202.420 ;
        RECT 31.140 202.220 32.660 202.360 ;
        RECT 39.880 202.220 49.310 202.360 ;
        RECT 26.935 202.175 27.225 202.220 ;
        RECT 29.455 202.175 29.745 202.220 ;
        RECT 30.645 202.175 30.935 202.220 ;
        RECT 27.370 202.020 27.660 202.065 ;
        RECT 28.940 202.020 29.230 202.065 ;
        RECT 31.040 202.020 31.330 202.065 ;
        RECT 27.370 201.880 31.330 202.020 ;
        RECT 27.370 201.835 27.660 201.880 ;
        RECT 28.940 201.835 29.230 201.880 ;
        RECT 31.040 201.835 31.330 201.880 ;
        RECT 32.520 201.740 32.660 202.220 ;
        RECT 48.990 202.160 49.310 202.220 ;
        RECT 54.050 202.160 54.370 202.420 ;
        RECT 60.045 202.175 60.335 202.405 ;
        RECT 60.925 202.360 61.215 202.405 ;
        RECT 62.115 202.360 62.405 202.405 ;
        RECT 64.635 202.360 64.925 202.405 ;
        RECT 60.925 202.220 64.925 202.360 ;
        RECT 60.925 202.175 61.215 202.220 ;
        RECT 62.115 202.175 62.405 202.220 ;
        RECT 64.635 202.175 64.925 202.220 ;
        RECT 70.150 202.360 70.470 202.420 ;
        RECT 72.540 202.360 72.680 202.515 ;
        RECT 72.910 202.500 73.230 202.760 ;
        RECT 73.845 202.515 74.135 202.745 ;
        RECT 76.605 202.700 76.895 202.745 ;
        RECT 80.285 202.700 80.575 202.745 ;
        RECT 76.605 202.560 82.110 202.700 ;
        RECT 76.605 202.515 76.895 202.560 ;
        RECT 80.285 202.515 80.575 202.560 ;
        RECT 73.920 202.360 74.060 202.515 ;
        RECT 70.150 202.220 74.060 202.360 ;
        RECT 81.970 202.360 82.110 202.560 ;
        RECT 92.690 202.500 93.010 202.760 ;
        RECT 93.240 202.700 93.380 202.900 ;
        RECT 95.910 202.840 96.230 203.100 ;
        RECT 96.460 203.040 96.600 203.240 ;
        RECT 96.830 203.180 97.150 203.440 ;
        RECT 100.510 203.180 100.830 203.440 ;
        RECT 112.470 203.380 112.790 203.440 ;
        RECT 113.405 203.380 113.695 203.425 ;
        RECT 127.650 203.380 127.970 203.440 ;
        RECT 138.230 203.380 138.550 203.440 ;
        RECT 112.470 203.240 127.970 203.380 ;
        RECT 112.470 203.180 112.790 203.240 ;
        RECT 113.405 203.195 113.695 203.240 ;
        RECT 127.650 203.180 127.970 203.240 ;
        RECT 131.420 203.240 138.550 203.380 ;
        RECT 96.460 202.900 98.900 203.040 ;
        RECT 98.760 202.745 98.900 202.900 ;
        RECT 101.445 202.855 101.735 203.085 ;
        RECT 103.730 203.040 104.050 203.100 ;
        RECT 104.205 203.040 104.495 203.085 ;
        RECT 126.730 203.040 127.050 203.100 ;
        RECT 131.420 203.085 131.560 203.240 ;
        RECT 138.230 203.180 138.550 203.240 ;
        RECT 140.530 203.180 140.850 203.440 ;
        RECT 131.345 203.040 131.635 203.085 ;
        RECT 103.730 202.900 104.495 203.040 ;
        RECT 98.225 202.700 98.515 202.745 ;
        RECT 93.240 202.560 98.515 202.700 ;
        RECT 96.000 202.420 96.140 202.560 ;
        RECT 98.225 202.515 98.515 202.560 ;
        RECT 98.685 202.515 98.975 202.745 ;
        RECT 82.570 202.360 82.890 202.420 ;
        RECT 81.970 202.220 82.890 202.360 ;
        RECT 32.430 201.680 32.750 201.740 ;
        RECT 32.905 201.680 33.195 201.725 ;
        RECT 32.430 201.540 33.195 201.680 ;
        RECT 32.430 201.480 32.750 201.540 ;
        RECT 32.905 201.495 33.195 201.540 ;
        RECT 37.950 201.680 38.270 201.740 ;
        RECT 39.345 201.680 39.635 201.725 ;
        RECT 37.950 201.540 39.635 201.680 ;
        RECT 60.120 201.680 60.260 202.175 ;
        RECT 70.150 202.160 70.470 202.220 ;
        RECT 82.570 202.160 82.890 202.220 ;
        RECT 83.030 202.360 83.350 202.420 ;
        RECT 83.505 202.360 83.795 202.405 ;
        RECT 83.030 202.220 83.795 202.360 ;
        RECT 83.030 202.160 83.350 202.220 ;
        RECT 83.505 202.175 83.795 202.220 ;
        RECT 84.385 202.360 84.675 202.405 ;
        RECT 85.575 202.360 85.865 202.405 ;
        RECT 88.095 202.360 88.385 202.405 ;
        RECT 84.385 202.220 88.385 202.360 ;
        RECT 84.385 202.175 84.675 202.220 ;
        RECT 85.575 202.175 85.865 202.220 ;
        RECT 88.095 202.175 88.385 202.220 ;
        RECT 95.910 202.160 96.230 202.420 ;
        RECT 96.830 202.360 97.150 202.420 ;
        RECT 101.520 202.360 101.660 202.855 ;
        RECT 103.730 202.840 104.050 202.900 ;
        RECT 104.205 202.855 104.495 202.900 ;
        RECT 106.580 202.900 114.080 203.040 ;
        RECT 106.580 202.405 106.720 202.900 ;
        RECT 107.870 202.745 108.190 202.760 ;
        RECT 113.940 202.745 114.080 202.900 ;
        RECT 126.730 202.900 129.720 203.040 ;
        RECT 126.730 202.840 127.050 202.900 ;
        RECT 107.840 202.700 108.190 202.745 ;
        RECT 107.675 202.560 108.190 202.700 ;
        RECT 107.840 202.515 108.190 202.560 ;
        RECT 113.865 202.515 114.155 202.745 ;
        RECT 114.310 202.700 114.630 202.760 ;
        RECT 115.145 202.700 115.435 202.745 ;
        RECT 114.310 202.560 115.435 202.700 ;
        RECT 107.870 202.500 108.190 202.515 ;
        RECT 114.310 202.500 114.630 202.560 ;
        RECT 115.145 202.515 115.435 202.560 ;
        RECT 122.130 202.700 122.450 202.760 ;
        RECT 127.190 202.700 127.510 202.760 ;
        RECT 122.130 202.560 126.960 202.700 ;
        RECT 122.130 202.500 122.450 202.560 ;
        RECT 126.820 202.405 126.960 202.560 ;
        RECT 127.190 202.560 128.340 202.700 ;
        RECT 127.190 202.500 127.510 202.560 ;
        RECT 106.505 202.360 106.795 202.405 ;
        RECT 96.830 202.220 101.660 202.360 ;
        RECT 104.280 202.220 106.795 202.360 ;
        RECT 96.830 202.160 97.150 202.220 ;
        RECT 104.280 202.080 104.420 202.220 ;
        RECT 106.505 202.175 106.795 202.220 ;
        RECT 107.385 202.360 107.675 202.405 ;
        RECT 108.575 202.360 108.865 202.405 ;
        RECT 111.095 202.360 111.385 202.405 ;
        RECT 107.385 202.220 111.385 202.360 ;
        RECT 107.385 202.175 107.675 202.220 ;
        RECT 108.575 202.175 108.865 202.220 ;
        RECT 111.095 202.175 111.385 202.220 ;
        RECT 114.745 202.360 115.035 202.405 ;
        RECT 115.935 202.360 116.225 202.405 ;
        RECT 118.455 202.360 118.745 202.405 ;
        RECT 123.985 202.360 124.275 202.405 ;
        RECT 114.745 202.220 118.745 202.360 ;
        RECT 114.745 202.175 115.035 202.220 ;
        RECT 115.935 202.175 116.225 202.220 ;
        RECT 118.455 202.175 118.745 202.220 ;
        RECT 120.840 202.220 124.275 202.360 ;
        RECT 60.530 202.020 60.820 202.065 ;
        RECT 62.630 202.020 62.920 202.065 ;
        RECT 64.200 202.020 64.490 202.065 ;
        RECT 60.530 201.880 64.490 202.020 ;
        RECT 60.530 201.835 60.820 201.880 ;
        RECT 62.630 201.835 62.920 201.880 ;
        RECT 64.200 201.835 64.490 201.880 ;
        RECT 83.990 202.020 84.280 202.065 ;
        RECT 86.090 202.020 86.380 202.065 ;
        RECT 87.660 202.020 87.950 202.065 ;
        RECT 83.990 201.880 87.950 202.020 ;
        RECT 83.990 201.835 84.280 201.880 ;
        RECT 86.090 201.835 86.380 201.880 ;
        RECT 87.660 201.835 87.950 201.880 ;
        RECT 94.085 202.020 94.375 202.065 ;
        RECT 96.370 202.020 96.690 202.080 ;
        RECT 97.305 202.020 97.595 202.065 ;
        RECT 94.085 201.880 97.595 202.020 ;
        RECT 94.085 201.835 94.375 201.880 ;
        RECT 96.370 201.820 96.690 201.880 ;
        RECT 97.305 201.835 97.595 201.880 ;
        RECT 102.810 202.020 103.130 202.080 ;
        RECT 103.285 202.020 103.575 202.065 ;
        RECT 102.810 201.880 103.575 202.020 ;
        RECT 102.810 201.820 103.130 201.880 ;
        RECT 103.285 201.835 103.575 201.880 ;
        RECT 104.190 201.820 104.510 202.080 ;
        RECT 106.990 202.020 107.280 202.065 ;
        RECT 109.090 202.020 109.380 202.065 ;
        RECT 110.660 202.020 110.950 202.065 ;
        RECT 106.990 201.880 110.950 202.020 ;
        RECT 106.990 201.835 107.280 201.880 ;
        RECT 109.090 201.835 109.380 201.880 ;
        RECT 110.660 201.835 110.950 201.880 ;
        RECT 114.350 202.020 114.640 202.065 ;
        RECT 116.450 202.020 116.740 202.065 ;
        RECT 118.020 202.020 118.310 202.065 ;
        RECT 114.350 201.880 118.310 202.020 ;
        RECT 114.350 201.835 114.640 201.880 ;
        RECT 116.450 201.835 116.740 201.880 ;
        RECT 118.020 201.835 118.310 201.880 ;
        RECT 120.290 202.020 120.610 202.080 ;
        RECT 120.840 202.065 120.980 202.220 ;
        RECT 123.985 202.175 124.275 202.220 ;
        RECT 126.745 202.175 127.035 202.405 ;
        RECT 127.665 202.175 127.955 202.405 ;
        RECT 128.200 202.360 128.340 202.560 ;
        RECT 129.030 202.500 129.350 202.760 ;
        RECT 129.580 202.745 129.720 202.900 ;
        RECT 130.270 202.900 131.635 203.040 ;
        RECT 129.505 202.515 129.795 202.745 ;
        RECT 130.270 202.360 130.410 202.900 ;
        RECT 131.345 202.855 131.635 202.900 ;
        RECT 132.250 202.840 132.570 203.100 ;
        RECT 132.725 203.040 133.015 203.085 ;
        RECT 133.630 203.040 133.950 203.100 ;
        RECT 132.725 202.900 133.950 203.040 ;
        RECT 132.725 202.855 133.015 202.900 ;
        RECT 133.630 202.840 133.950 202.900 ;
        RECT 135.485 203.040 135.775 203.085 ;
        RECT 139.625 203.040 139.915 203.085 ;
        RECT 145.130 203.040 145.450 203.100 ;
        RECT 135.485 202.900 145.450 203.040 ;
        RECT 135.485 202.855 135.775 202.900 ;
        RECT 139.625 202.855 139.915 202.900 ;
        RECT 145.130 202.840 145.450 202.900 ;
        RECT 133.170 202.500 133.490 202.760 ;
        RECT 134.105 202.700 134.395 202.745 ;
        RECT 137.310 202.700 137.630 202.760 ;
        RECT 137.785 202.700 138.075 202.745 ;
        RECT 134.105 202.560 138.075 202.700 ;
        RECT 134.105 202.515 134.395 202.560 ;
        RECT 137.310 202.500 137.630 202.560 ;
        RECT 137.785 202.515 138.075 202.560 ;
        RECT 143.765 202.700 144.055 202.745 ;
        RECT 152.045 202.700 152.335 202.745 ;
        RECT 143.765 202.560 152.335 202.700 ;
        RECT 143.765 202.515 144.055 202.560 ;
        RECT 152.045 202.515 152.335 202.560 ;
        RECT 128.200 202.220 130.410 202.360 ;
        RECT 141.450 202.360 141.770 202.420 ;
        RECT 142.370 202.360 142.690 202.420 ;
        RECT 143.305 202.360 143.595 202.405 ;
        RECT 141.450 202.220 143.595 202.360 ;
        RECT 120.765 202.020 121.055 202.065 ;
        RECT 120.290 201.880 121.055 202.020 ;
        RECT 127.740 202.020 127.880 202.175 ;
        RECT 141.450 202.160 141.770 202.220 ;
        RECT 142.370 202.160 142.690 202.220 ;
        RECT 143.305 202.175 143.595 202.220 ;
        RECT 154.790 202.160 155.110 202.420 ;
        RECT 132.710 202.020 133.030 202.080 ;
        RECT 136.850 202.020 137.170 202.080 ;
        RECT 137.325 202.020 137.615 202.065 ;
        RECT 127.740 201.880 130.180 202.020 ;
        RECT 120.290 201.820 120.610 201.880 ;
        RECT 120.765 201.835 121.055 201.880 ;
        RECT 130.040 201.740 130.180 201.880 ;
        RECT 132.710 201.880 136.160 202.020 ;
        RECT 132.710 201.820 133.030 201.880 ;
        RECT 61.870 201.680 62.190 201.740 ;
        RECT 60.120 201.540 62.190 201.680 ;
        RECT 37.950 201.480 38.270 201.540 ;
        RECT 39.345 201.495 39.635 201.540 ;
        RECT 61.870 201.480 62.190 201.540 ;
        RECT 81.190 201.480 81.510 201.740 ;
        RECT 86.710 201.680 87.030 201.740 ;
        RECT 90.405 201.680 90.695 201.725 ;
        RECT 86.710 201.540 90.695 201.680 ;
        RECT 86.710 201.480 87.030 201.540 ;
        RECT 90.405 201.495 90.695 201.540 ;
        RECT 93.625 201.680 93.915 201.725 ;
        RECT 95.925 201.680 96.215 201.725 ;
        RECT 93.625 201.540 96.215 201.680 ;
        RECT 93.625 201.495 93.915 201.540 ;
        RECT 95.925 201.495 96.215 201.540 ;
        RECT 98.210 201.680 98.530 201.740 ;
        RECT 101.445 201.680 101.735 201.725 ;
        RECT 98.210 201.540 101.735 201.680 ;
        RECT 98.210 201.480 98.530 201.540 ;
        RECT 101.445 201.495 101.735 201.540 ;
        RECT 104.650 201.480 104.970 201.740 ;
        RECT 121.210 201.480 121.530 201.740 ;
        RECT 127.190 201.680 127.510 201.740 ;
        RECT 128.585 201.680 128.875 201.725 ;
        RECT 127.190 201.540 128.875 201.680 ;
        RECT 127.190 201.480 127.510 201.540 ;
        RECT 128.585 201.495 128.875 201.540 ;
        RECT 129.950 201.480 130.270 201.740 ;
        RECT 130.870 201.480 131.190 201.740 ;
        RECT 134.550 201.480 134.870 201.740 ;
        RECT 135.470 201.480 135.790 201.740 ;
        RECT 136.020 201.680 136.160 201.880 ;
        RECT 136.850 201.880 137.615 202.020 ;
        RECT 136.850 201.820 137.170 201.880 ;
        RECT 137.325 201.835 137.615 201.880 ;
        RECT 145.605 202.020 145.895 202.065 ;
        RECT 146.970 202.020 147.290 202.080 ;
        RECT 145.605 201.880 147.290 202.020 ;
        RECT 145.605 201.835 145.895 201.880 ;
        RECT 146.970 201.820 147.290 201.880 ;
        RECT 137.770 201.680 138.090 201.740 ;
        RECT 136.020 201.540 138.090 201.680 ;
        RECT 137.770 201.480 138.090 201.540 ;
        RECT 138.690 201.680 139.010 201.740 ;
        RECT 139.625 201.680 139.915 201.725 ;
        RECT 138.690 201.540 139.915 201.680 ;
        RECT 138.690 201.480 139.010 201.540 ;
        RECT 139.625 201.495 139.915 201.540 ;
        RECT 22.700 200.860 157.020 201.340 ;
        RECT 49.925 200.660 50.215 200.705 ;
        RECT 54.970 200.660 55.290 200.720 ;
        RECT 49.925 200.520 55.290 200.660 ;
        RECT 49.925 200.475 50.215 200.520 ;
        RECT 54.970 200.460 55.290 200.520 ;
        RECT 62.790 200.460 63.110 200.720 ;
        RECT 77.050 200.460 77.370 200.720 ;
        RECT 98.210 200.460 98.530 200.720 ;
        RECT 101.445 200.660 101.735 200.705 ;
        RECT 103.270 200.660 103.590 200.720 ;
        RECT 101.445 200.520 103.590 200.660 ;
        RECT 101.445 200.475 101.735 200.520 ;
        RECT 103.270 200.460 103.590 200.520 ;
        RECT 113.405 200.660 113.695 200.705 ;
        RECT 114.310 200.660 114.630 200.720 ;
        RECT 113.405 200.520 114.630 200.660 ;
        RECT 113.405 200.475 113.695 200.520 ;
        RECT 114.310 200.460 114.630 200.520 ;
        RECT 121.670 200.460 121.990 200.720 ;
        RECT 127.190 200.460 127.510 200.720 ;
        RECT 132.725 200.475 133.015 200.705 ;
        RECT 37.990 200.320 38.280 200.365 ;
        RECT 40.090 200.320 40.380 200.365 ;
        RECT 41.660 200.320 41.950 200.365 ;
        RECT 48.530 200.320 48.850 200.380 ;
        RECT 37.990 200.180 41.950 200.320 ;
        RECT 37.990 200.135 38.280 200.180 ;
        RECT 40.090 200.135 40.380 200.180 ;
        RECT 41.660 200.135 41.950 200.180 ;
        RECT 46.320 200.180 48.850 200.320 ;
        RECT 37.490 199.780 37.810 200.040 ;
        RECT 38.385 199.980 38.675 200.025 ;
        RECT 39.575 199.980 39.865 200.025 ;
        RECT 42.095 199.980 42.385 200.025 ;
        RECT 38.385 199.840 42.385 199.980 ;
        RECT 38.385 199.795 38.675 199.840 ;
        RECT 39.575 199.795 39.865 199.840 ;
        RECT 42.095 199.795 42.385 199.840 ;
        RECT 37.950 199.640 38.270 199.700 ;
        RECT 38.785 199.640 39.075 199.685 ;
        RECT 37.950 199.500 39.075 199.640 ;
        RECT 37.950 199.440 38.270 199.500 ;
        RECT 38.785 199.455 39.075 199.500 ;
        RECT 45.785 199.640 46.075 199.685 ;
        RECT 46.320 199.640 46.460 200.180 ;
        RECT 48.530 200.120 48.850 200.180 ;
        RECT 49.465 200.320 49.755 200.365 ;
        RECT 51.750 200.320 52.070 200.380 ;
        RECT 49.465 200.180 52.070 200.320 ;
        RECT 49.465 200.135 49.755 200.180 ;
        RECT 51.750 200.120 52.070 200.180 ;
        RECT 61.885 200.320 62.175 200.365 ;
        RECT 64.170 200.320 64.490 200.380 ;
        RECT 61.885 200.180 64.490 200.320 ;
        RECT 61.885 200.135 62.175 200.180 ;
        RECT 64.170 200.120 64.490 200.180 ;
        RECT 64.645 200.320 64.935 200.365 ;
        RECT 65.105 200.320 65.395 200.365 ;
        RECT 70.150 200.320 70.470 200.380 ;
        RECT 64.645 200.180 70.470 200.320 ;
        RECT 64.645 200.135 64.935 200.180 ;
        RECT 65.105 200.135 65.395 200.180 ;
        RECT 70.150 200.120 70.470 200.180 ;
        RECT 82.570 200.320 82.890 200.380 ;
        RECT 105.570 200.320 105.890 200.380 ;
        RECT 127.650 200.320 127.970 200.380 ;
        RECT 128.125 200.320 128.415 200.365 ;
        RECT 82.570 200.180 127.420 200.320 ;
        RECT 82.570 200.120 82.890 200.180 ;
        RECT 105.570 200.120 105.890 200.180 ;
        RECT 71.530 199.980 71.850 200.040 ;
        RECT 81.650 199.980 81.970 200.040 ;
        RECT 88.090 199.980 88.410 200.040 ;
        RECT 45.785 199.500 46.460 199.640 ;
        RECT 46.780 199.840 51.060 199.980 ;
        RECT 45.785 199.455 46.075 199.500 ;
        RECT 46.780 199.360 46.920 199.840 ;
        RECT 47.165 199.455 47.455 199.685 ;
        RECT 47.625 199.640 47.915 199.685 ;
        RECT 48.070 199.640 48.390 199.700 ;
        RECT 47.625 199.500 48.390 199.640 ;
        RECT 47.625 199.455 47.915 199.500 ;
        RECT 46.690 199.300 47.010 199.360 ;
        RECT 44.480 199.160 47.010 199.300 ;
        RECT 47.240 199.300 47.380 199.455 ;
        RECT 48.070 199.440 48.390 199.500 ;
        RECT 48.530 199.640 48.850 199.700 ;
        RECT 50.370 199.640 50.690 199.700 ;
        RECT 50.920 199.685 51.060 199.840 ;
        RECT 70.240 199.840 71.850 199.980 ;
        RECT 48.530 199.500 50.690 199.640 ;
        RECT 48.530 199.440 48.850 199.500 ;
        RECT 50.370 199.440 50.690 199.500 ;
        RECT 50.845 199.455 51.135 199.685 ;
        RECT 65.105 199.455 65.395 199.685 ;
        RECT 66.025 199.640 66.315 199.685 ;
        RECT 66.470 199.640 66.790 199.700 ;
        RECT 66.025 199.500 66.790 199.640 ;
        RECT 66.025 199.455 66.315 199.500 ;
        RECT 51.765 199.300 52.055 199.345 ;
        RECT 53.130 199.300 53.450 199.360 ;
        RECT 47.240 199.160 47.840 199.300 ;
        RECT 44.480 199.005 44.620 199.160 ;
        RECT 46.690 199.100 47.010 199.160 ;
        RECT 47.700 199.020 47.840 199.160 ;
        RECT 51.765 199.160 53.450 199.300 ;
        RECT 51.765 199.115 52.055 199.160 ;
        RECT 53.130 199.100 53.450 199.160 ;
        RECT 61.410 199.300 61.730 199.360 ;
        RECT 65.180 199.300 65.320 199.455 ;
        RECT 66.470 199.440 66.790 199.500 ;
        RECT 67.865 199.640 68.155 199.685 ;
        RECT 69.690 199.640 70.010 199.700 ;
        RECT 70.240 199.685 70.380 199.840 ;
        RECT 71.530 199.780 71.850 199.840 ;
        RECT 78.060 199.840 88.410 199.980 ;
        RECT 67.865 199.500 70.010 199.640 ;
        RECT 67.865 199.455 68.155 199.500 ;
        RECT 69.690 199.440 70.010 199.500 ;
        RECT 70.165 199.455 70.455 199.685 ;
        RECT 71.070 199.440 71.390 199.700 ;
        RECT 78.060 199.685 78.200 199.840 ;
        RECT 81.650 199.780 81.970 199.840 ;
        RECT 88.090 199.780 88.410 199.840 ;
        RECT 93.610 199.980 93.930 200.040 ;
        RECT 112.470 199.980 112.790 200.040 ;
        RECT 114.770 199.980 115.090 200.040 ;
        RECT 121.210 199.980 121.530 200.040 ;
        RECT 93.610 199.840 112.790 199.980 ;
        RECT 93.610 199.780 93.930 199.840 ;
        RECT 112.470 199.780 112.790 199.840 ;
        RECT 114.400 199.840 115.090 199.980 ;
        RECT 77.985 199.455 78.275 199.685 ;
        RECT 78.430 199.440 78.750 199.700 ;
        RECT 85.805 199.640 86.095 199.685 ;
        RECT 86.710 199.640 87.030 199.700 ;
        RECT 85.805 199.500 87.030 199.640 ;
        RECT 85.805 199.455 86.095 199.500 ;
        RECT 86.710 199.440 87.030 199.500 ;
        RECT 96.370 199.440 96.690 199.700 ;
        RECT 97.290 199.640 97.610 199.700 ;
        RECT 100.050 199.640 100.370 199.700 ;
        RECT 97.290 199.500 100.370 199.640 ;
        RECT 97.290 199.440 97.610 199.500 ;
        RECT 100.050 199.440 100.370 199.500 ;
        RECT 102.810 199.440 103.130 199.700 ;
        RECT 103.730 199.440 104.050 199.700 ;
        RECT 114.400 199.685 114.540 199.840 ;
        RECT 114.770 199.780 115.090 199.840 ;
        RECT 116.240 199.840 121.530 199.980 ;
        RECT 104.205 199.455 104.495 199.685 ;
        RECT 114.325 199.455 114.615 199.685 ;
        RECT 115.245 199.640 115.535 199.685 ;
        RECT 115.690 199.640 116.010 199.700 ;
        RECT 116.240 199.685 116.380 199.840 ;
        RECT 121.210 199.780 121.530 199.840 ;
        RECT 122.605 199.980 122.895 200.025 ;
        RECT 124.430 199.980 124.750 200.040 ;
        RECT 122.605 199.840 124.750 199.980 ;
        RECT 122.605 199.795 122.895 199.840 ;
        RECT 124.430 199.780 124.750 199.840 ;
        RECT 126.730 199.780 127.050 200.040 ;
        RECT 127.280 199.980 127.420 200.180 ;
        RECT 127.650 200.180 128.415 200.320 ;
        RECT 132.800 200.320 132.940 200.475 ;
        RECT 135.470 200.460 135.790 200.720 ;
        RECT 137.770 200.660 138.090 200.720 ;
        RECT 154.345 200.660 154.635 200.705 ;
        RECT 154.790 200.660 155.110 200.720 ;
        RECT 137.400 200.520 155.110 200.660 ;
        RECT 133.630 200.320 133.950 200.380 ;
        RECT 136.390 200.320 136.710 200.380 ;
        RECT 132.800 200.180 136.710 200.320 ;
        RECT 127.650 200.120 127.970 200.180 ;
        RECT 128.125 200.135 128.415 200.180 ;
        RECT 133.630 200.120 133.950 200.180 ;
        RECT 132.710 199.980 133.030 200.040 ;
        RECT 127.280 199.840 133.030 199.980 ;
        RECT 132.710 199.780 133.030 199.840 ;
        RECT 115.245 199.500 116.010 199.640 ;
        RECT 115.245 199.455 115.535 199.500 ;
        RECT 61.410 199.160 65.320 199.300 ;
        RECT 61.410 199.100 61.730 199.160 ;
        RECT 74.750 199.100 75.070 199.360 ;
        RECT 75.670 199.100 75.990 199.360 ;
        RECT 77.065 199.300 77.355 199.345 ;
        RECT 80.730 199.300 81.050 199.360 ;
        RECT 77.065 199.160 81.050 199.300 ;
        RECT 77.065 199.115 77.355 199.160 ;
        RECT 80.730 199.100 81.050 199.160 ;
        RECT 84.885 199.300 85.175 199.345 ;
        RECT 85.330 199.300 85.650 199.360 ;
        RECT 84.885 199.160 85.650 199.300 ;
        RECT 84.885 199.115 85.175 199.160 ;
        RECT 85.330 199.100 85.650 199.160 ;
        RECT 99.130 199.300 99.450 199.360 ;
        RECT 100.525 199.300 100.815 199.345 ;
        RECT 99.130 199.160 100.815 199.300 ;
        RECT 99.130 199.100 99.450 199.160 ;
        RECT 100.525 199.115 100.815 199.160 ;
        RECT 103.270 199.100 103.590 199.360 ;
        RECT 104.280 199.300 104.420 199.455 ;
        RECT 115.690 199.440 116.010 199.500 ;
        RECT 116.165 199.455 116.455 199.685 ;
        RECT 120.290 199.440 120.610 199.700 ;
        RECT 126.270 199.440 126.590 199.700 ;
        RECT 132.250 199.640 132.570 199.700 ;
        RECT 134.550 199.640 134.870 199.700 ;
        RECT 131.880 199.500 134.870 199.640 ;
        RECT 103.820 199.160 104.420 199.300 ;
        RECT 114.785 199.300 115.075 199.345 ;
        RECT 117.070 199.300 117.390 199.360 ;
        RECT 114.785 199.160 117.390 199.300 ;
        RECT 44.405 198.775 44.695 199.005 ;
        RECT 44.850 198.760 45.170 199.020 ;
        RECT 47.610 198.760 47.930 199.020 ;
        RECT 48.070 198.960 48.390 199.020 ;
        RECT 50.385 198.960 50.675 199.005 ;
        RECT 48.070 198.820 50.675 198.960 ;
        RECT 48.070 198.760 48.390 198.820 ;
        RECT 50.385 198.775 50.675 198.820 ;
        RECT 62.790 198.960 63.110 199.020 ;
        RECT 63.710 198.960 64.030 199.020 ;
        RECT 62.790 198.820 64.030 198.960 ;
        RECT 62.790 198.760 63.110 198.820 ;
        RECT 63.710 198.760 64.030 198.820 ;
        RECT 66.930 198.760 67.250 199.020 ;
        RECT 70.610 198.760 70.930 199.020 ;
        RECT 76.590 198.760 76.910 199.020 ;
        RECT 86.250 198.960 86.570 199.020 ;
        RECT 101.430 199.005 101.750 199.020 ;
        RECT 86.725 198.960 87.015 199.005 ;
        RECT 86.250 198.820 87.015 198.960 ;
        RECT 86.250 198.760 86.570 198.820 ;
        RECT 86.725 198.775 87.015 198.820 ;
        RECT 101.430 198.775 101.815 199.005 ;
        RECT 102.365 198.960 102.655 199.005 ;
        RECT 103.820 198.960 103.960 199.160 ;
        RECT 114.785 199.115 115.075 199.160 ;
        RECT 117.070 199.100 117.390 199.160 ;
        RECT 121.670 199.300 121.990 199.360 ;
        RECT 131.880 199.345 132.020 199.500 ;
        RECT 132.250 199.440 132.570 199.500 ;
        RECT 134.550 199.440 134.870 199.500 ;
        RECT 135.025 199.640 135.315 199.685 ;
        RECT 135.560 199.640 135.700 200.180 ;
        RECT 136.390 200.120 136.710 200.180 ;
        RECT 135.025 199.500 135.700 199.640 ;
        RECT 135.930 199.640 136.250 199.700 ;
        RECT 136.405 199.640 136.695 199.685 ;
        RECT 135.930 199.500 136.695 199.640 ;
        RECT 135.025 199.455 135.315 199.500 ;
        RECT 135.930 199.440 136.250 199.500 ;
        RECT 136.405 199.455 136.695 199.500 ;
        RECT 137.400 199.345 137.540 200.520 ;
        RECT 137.770 200.460 138.090 200.520 ;
        RECT 154.345 200.475 154.635 200.520 ;
        RECT 154.790 200.460 155.110 200.520 ;
        RECT 140.570 200.320 140.860 200.365 ;
        RECT 142.670 200.320 142.960 200.365 ;
        RECT 144.240 200.320 144.530 200.365 ;
        RECT 140.570 200.180 144.530 200.320 ;
        RECT 140.570 200.135 140.860 200.180 ;
        RECT 142.670 200.135 142.960 200.180 ;
        RECT 144.240 200.135 144.530 200.180 ;
        RECT 147.930 200.320 148.220 200.365 ;
        RECT 150.030 200.320 150.320 200.365 ;
        RECT 151.600 200.320 151.890 200.365 ;
        RECT 147.930 200.180 151.890 200.320 ;
        RECT 147.930 200.135 148.220 200.180 ;
        RECT 150.030 200.135 150.320 200.180 ;
        RECT 151.600 200.135 151.890 200.180 ;
        RECT 140.070 199.780 140.390 200.040 ;
        RECT 140.965 199.980 141.255 200.025 ;
        RECT 142.155 199.980 142.445 200.025 ;
        RECT 144.675 199.980 144.965 200.025 ;
        RECT 140.965 199.840 144.965 199.980 ;
        RECT 140.965 199.795 141.255 199.840 ;
        RECT 142.155 199.795 142.445 199.840 ;
        RECT 144.675 199.795 144.965 199.840 ;
        RECT 148.325 199.980 148.615 200.025 ;
        RECT 149.515 199.980 149.805 200.025 ;
        RECT 152.035 199.980 152.325 200.025 ;
        RECT 148.325 199.840 152.325 199.980 ;
        RECT 148.325 199.795 148.615 199.840 ;
        RECT 149.515 199.795 149.805 199.840 ;
        RECT 152.035 199.795 152.325 199.840 ;
        RECT 137.785 199.640 138.075 199.685 ;
        RECT 140.530 199.640 140.850 199.700 ;
        RECT 137.785 199.500 140.850 199.640 ;
        RECT 137.785 199.455 138.075 199.500 ;
        RECT 140.530 199.440 140.850 199.500 ;
        RECT 147.430 199.640 147.750 199.700 ;
        RECT 150.650 199.640 150.970 199.700 ;
        RECT 147.430 199.500 150.970 199.640 ;
        RECT 147.430 199.440 147.750 199.500 ;
        RECT 150.650 199.440 150.970 199.500 ;
        RECT 141.450 199.345 141.770 199.360 ;
        RECT 131.805 199.300 132.095 199.345 ;
        RECT 121.670 199.160 132.095 199.300 ;
        RECT 121.670 199.100 121.990 199.160 ;
        RECT 131.805 199.115 132.095 199.160 ;
        RECT 133.720 199.160 137.080 199.300 ;
        RECT 102.365 198.820 103.960 198.960 ;
        RECT 102.365 198.775 102.655 198.820 ;
        RECT 101.430 198.760 101.750 198.775 ;
        RECT 105.110 198.760 105.430 199.020 ;
        RECT 132.710 199.005 133.030 199.020 ;
        RECT 133.720 199.005 133.860 199.160 ;
        RECT 136.940 199.020 137.080 199.160 ;
        RECT 137.325 199.115 137.615 199.345 ;
        RECT 141.420 199.115 141.770 199.345 ;
        RECT 141.450 199.100 141.770 199.115 ;
        RECT 141.910 199.300 142.230 199.360 ;
        RECT 147.890 199.300 148.210 199.360 ;
        RECT 148.670 199.300 148.960 199.345 ;
        RECT 141.910 199.160 147.200 199.300 ;
        RECT 141.910 199.100 142.230 199.160 ;
        RECT 132.710 198.775 133.095 199.005 ;
        RECT 133.645 198.775 133.935 199.005 ;
        RECT 132.710 198.760 133.030 198.775 ;
        RECT 134.550 198.760 134.870 199.020 ;
        RECT 136.850 198.760 137.170 199.020 ;
        RECT 147.060 199.005 147.200 199.160 ;
        RECT 147.890 199.160 148.960 199.300 ;
        RECT 147.890 199.100 148.210 199.160 ;
        RECT 148.670 199.115 148.960 199.160 ;
        RECT 146.985 198.775 147.275 199.005 ;
        RECT 22.700 198.140 157.820 198.620 ;
        RECT 35.190 197.940 35.510 198.000 ;
        RECT 36.570 197.940 36.890 198.000 ;
        RECT 40.710 197.940 41.030 198.000 ;
        RECT 42.105 197.940 42.395 197.985 ;
        RECT 35.190 197.800 40.020 197.940 ;
        RECT 35.190 197.740 35.510 197.800 ;
        RECT 36.570 197.740 36.890 197.800 ;
        RECT 37.490 197.600 37.810 197.660 ;
        RECT 39.880 197.600 40.020 197.800 ;
        RECT 40.710 197.800 42.395 197.940 ;
        RECT 40.710 197.740 41.030 197.800 ;
        RECT 42.105 197.755 42.395 197.800 ;
        RECT 42.945 197.940 43.235 197.985 ;
        RECT 44.850 197.940 45.170 198.000 ;
        RECT 42.945 197.800 45.170 197.940 ;
        RECT 42.945 197.755 43.235 197.800 ;
        RECT 44.850 197.740 45.170 197.800 ;
        RECT 48.990 197.740 49.310 198.000 ;
        RECT 54.050 197.940 54.370 198.000 ;
        RECT 71.530 197.940 71.850 198.000 ;
        RECT 86.265 197.940 86.555 197.985 ;
        RECT 54.050 197.800 63.480 197.940 ;
        RECT 54.050 197.740 54.370 197.800 ;
        RECT 60.490 197.645 60.810 197.660 ;
        RECT 43.945 197.600 44.235 197.645 ;
        RECT 37.490 197.460 39.560 197.600 ;
        RECT 39.880 197.460 44.235 197.600 ;
        RECT 37.490 197.400 37.810 197.460 ;
        RECT 37.950 197.305 38.270 197.320 ;
        RECT 39.420 197.305 39.560 197.460 ;
        RECT 43.945 197.415 44.235 197.460 ;
        RECT 60.425 197.415 60.810 197.645 ;
        RECT 61.425 197.600 61.715 197.645 ;
        RECT 62.790 197.600 63.110 197.660 ;
        RECT 61.425 197.460 63.110 197.600 ;
        RECT 61.425 197.415 61.715 197.460 ;
        RECT 60.490 197.400 60.810 197.415 ;
        RECT 62.790 197.400 63.110 197.460 ;
        RECT 37.950 197.075 38.300 197.305 ;
        RECT 39.345 197.075 39.635 197.305 ;
        RECT 46.690 197.260 47.010 197.320 ;
        RECT 53.590 197.305 53.910 197.320 ;
        RECT 50.845 197.260 51.135 197.305 ;
        RECT 46.690 197.120 51.135 197.260 ;
        RECT 37.950 197.060 38.270 197.075 ;
        RECT 46.690 197.060 47.010 197.120 ;
        RECT 50.845 197.075 51.135 197.120 ;
        RECT 53.560 197.075 53.910 197.305 ;
        RECT 53.590 197.060 53.910 197.075 ;
        RECT 59.110 197.260 59.430 197.320 ;
        RECT 63.340 197.305 63.480 197.800 ;
        RECT 71.530 197.800 72.680 197.940 ;
        RECT 71.530 197.740 71.850 197.800 ;
        RECT 65.980 197.600 66.270 197.645 ;
        RECT 66.930 197.600 67.250 197.660 ;
        RECT 65.980 197.460 67.250 197.600 ;
        RECT 72.540 197.600 72.680 197.800 ;
        RECT 81.970 197.800 86.555 197.940 ;
        RECT 77.510 197.600 77.830 197.660 ;
        RECT 77.985 197.600 78.275 197.645 ;
        RECT 81.970 197.600 82.110 197.800 ;
        RECT 86.265 197.755 86.555 197.800 ;
        RECT 87.185 197.940 87.475 197.985 ;
        RECT 88.550 197.940 88.870 198.000 ;
        RECT 95.910 197.985 96.230 198.000 ;
        RECT 87.185 197.800 88.870 197.940 ;
        RECT 87.185 197.755 87.475 197.800 ;
        RECT 72.540 197.460 73.200 197.600 ;
        RECT 65.980 197.415 66.270 197.460 ;
        RECT 66.930 197.400 67.250 197.460 ;
        RECT 61.885 197.260 62.175 197.305 ;
        RECT 59.110 197.120 62.175 197.260 ;
        RECT 59.110 197.060 59.430 197.120 ;
        RECT 61.885 197.075 62.175 197.120 ;
        RECT 62.345 197.075 62.635 197.305 ;
        RECT 63.265 197.260 63.555 197.305 ;
        RECT 68.770 197.260 69.090 197.320 ;
        RECT 73.060 197.305 73.200 197.460 ;
        RECT 77.510 197.460 82.110 197.600 ;
        RECT 86.340 197.600 86.480 197.755 ;
        RECT 88.550 197.740 88.870 197.800 ;
        RECT 90.940 197.800 95.680 197.940 ;
        RECT 90.940 197.645 91.080 197.800 ;
        RECT 90.865 197.600 91.155 197.645 ;
        RECT 86.340 197.460 91.155 197.600 ;
        RECT 77.510 197.400 77.830 197.460 ;
        RECT 77.985 197.415 78.275 197.460 ;
        RECT 90.865 197.415 91.155 197.460 ;
        RECT 95.005 197.415 95.295 197.645 ;
        RECT 95.540 197.600 95.680 197.800 ;
        RECT 95.910 197.755 96.295 197.985 ;
        RECT 96.845 197.940 97.135 197.985 ;
        RECT 101.430 197.940 101.750 198.000 ;
        RECT 102.365 197.940 102.655 197.985 ;
        RECT 96.845 197.800 100.740 197.940 ;
        RECT 96.845 197.755 97.135 197.800 ;
        RECT 95.910 197.740 96.230 197.755 ;
        RECT 99.130 197.600 99.450 197.660 ;
        RECT 100.600 197.645 100.740 197.800 ;
        RECT 101.430 197.800 102.655 197.940 ;
        RECT 101.430 197.740 101.750 197.800 ;
        RECT 102.365 197.755 102.655 197.800 ;
        RECT 138.690 197.740 139.010 198.000 ;
        RECT 141.005 197.940 141.295 197.985 ;
        RECT 141.450 197.940 141.770 198.000 ;
        RECT 141.005 197.800 141.770 197.940 ;
        RECT 141.005 197.755 141.295 197.800 ;
        RECT 141.450 197.740 141.770 197.800 ;
        RECT 147.890 197.740 148.210 198.000 ;
        RECT 95.540 197.460 99.450 197.600 ;
        RECT 63.265 197.120 69.090 197.260 ;
        RECT 63.265 197.075 63.555 197.120 ;
        RECT 34.755 196.920 35.045 196.965 ;
        RECT 37.275 196.920 37.565 196.965 ;
        RECT 38.465 196.920 38.755 196.965 ;
        RECT 34.755 196.780 38.755 196.920 ;
        RECT 34.755 196.735 35.045 196.780 ;
        RECT 37.275 196.735 37.565 196.780 ;
        RECT 38.465 196.735 38.755 196.780 ;
        RECT 51.305 196.735 51.595 196.965 ;
        RECT 35.190 196.580 35.480 196.625 ;
        RECT 36.760 196.580 37.050 196.625 ;
        RECT 38.860 196.580 39.150 196.625 ;
        RECT 35.190 196.440 39.150 196.580 ;
        RECT 35.190 196.395 35.480 196.440 ;
        RECT 36.760 196.395 37.050 196.440 ;
        RECT 38.860 196.395 39.150 196.440 ;
        RECT 32.445 196.240 32.735 196.285 ;
        RECT 34.270 196.240 34.590 196.300 ;
        RECT 32.445 196.100 34.590 196.240 ;
        RECT 32.445 196.055 32.735 196.100 ;
        RECT 34.270 196.040 34.590 196.100 ;
        RECT 43.025 196.240 43.315 196.285 ;
        RECT 48.070 196.240 48.390 196.300 ;
        RECT 43.025 196.100 48.390 196.240 ;
        RECT 51.380 196.240 51.520 196.735 ;
        RECT 52.210 196.720 52.530 196.980 ;
        RECT 53.105 196.920 53.395 196.965 ;
        RECT 54.295 196.920 54.585 196.965 ;
        RECT 56.815 196.920 57.105 196.965 ;
        RECT 53.105 196.780 57.105 196.920 ;
        RECT 53.105 196.735 53.395 196.780 ;
        RECT 54.295 196.735 54.585 196.780 ;
        RECT 56.815 196.735 57.105 196.780 ;
        RECT 60.030 196.920 60.350 196.980 ;
        RECT 62.420 196.920 62.560 197.075 ;
        RECT 68.770 197.060 69.090 197.120 ;
        RECT 71.945 197.075 72.235 197.305 ;
        RECT 72.925 197.075 73.215 197.305 ;
        RECT 74.765 197.075 75.055 197.305 ;
        RECT 84.425 197.260 84.715 197.305 ;
        RECT 84.870 197.260 85.190 197.320 ;
        RECT 92.245 197.260 92.535 197.305 ;
        RECT 84.425 197.120 92.535 197.260 ;
        RECT 84.425 197.075 84.715 197.120 ;
        RECT 60.030 196.780 62.560 196.920 ;
        RECT 60.030 196.720 60.350 196.780 ;
        RECT 64.645 196.735 64.935 196.965 ;
        RECT 65.525 196.920 65.815 196.965 ;
        RECT 66.715 196.920 67.005 196.965 ;
        RECT 69.235 196.920 69.525 196.965 ;
        RECT 65.525 196.780 69.525 196.920 ;
        RECT 65.525 196.735 65.815 196.780 ;
        RECT 66.715 196.735 67.005 196.780 ;
        RECT 69.235 196.735 69.525 196.780 ;
        RECT 71.070 196.920 71.390 196.980 ;
        RECT 72.035 196.920 72.175 197.075 ;
        RECT 74.840 196.920 74.980 197.075 ;
        RECT 84.870 197.060 85.190 197.120 ;
        RECT 92.245 197.075 92.535 197.120 ;
        RECT 93.150 197.060 93.470 197.320 ;
        RECT 95.080 197.260 95.220 197.415 ;
        RECT 99.130 197.400 99.450 197.460 ;
        RECT 100.525 197.600 100.815 197.645 ;
        RECT 102.810 197.600 103.130 197.660 ;
        RECT 130.885 197.600 131.175 197.645 ;
        RECT 144.210 197.600 144.530 197.660 ;
        RECT 100.525 197.460 103.130 197.600 ;
        RECT 100.525 197.415 100.815 197.460 ;
        RECT 102.810 197.400 103.130 197.460 ;
        RECT 104.280 197.460 113.620 197.600 ;
        RECT 97.290 197.260 97.610 197.320 ;
        RECT 95.080 197.120 97.610 197.260 ;
        RECT 97.290 197.060 97.610 197.120 ;
        RECT 97.765 197.260 98.055 197.305 ;
        RECT 98.670 197.260 98.990 197.320 ;
        RECT 97.765 197.120 98.990 197.260 ;
        RECT 97.765 197.075 98.055 197.120 ;
        RECT 71.070 196.780 72.175 196.920 ;
        RECT 72.540 196.780 74.980 196.920 ;
        RECT 89.025 196.920 89.315 196.965 ;
        RECT 89.470 196.920 89.790 196.980 ;
        RECT 95.910 196.920 96.230 196.980 ;
        RECT 89.025 196.780 96.230 196.920 ;
        RECT 52.710 196.580 53.000 196.625 ;
        RECT 54.810 196.580 55.100 196.625 ;
        RECT 56.380 196.580 56.670 196.625 ;
        RECT 52.710 196.440 56.670 196.580 ;
        RECT 52.710 196.395 53.000 196.440 ;
        RECT 54.810 196.395 55.100 196.440 ;
        RECT 56.380 196.395 56.670 196.440 ;
        RECT 57.270 196.580 57.590 196.640 ;
        RECT 59.585 196.580 59.875 196.625 ;
        RECT 57.270 196.440 59.875 196.580 ;
        RECT 57.270 196.380 57.590 196.440 ;
        RECT 59.585 196.395 59.875 196.440 ;
        RECT 61.410 196.580 61.730 196.640 ;
        RECT 61.885 196.580 62.175 196.625 ;
        RECT 61.410 196.440 62.175 196.580 ;
        RECT 61.410 196.380 61.730 196.440 ;
        RECT 61.885 196.395 62.175 196.440 ;
        RECT 62.330 196.580 62.650 196.640 ;
        RECT 64.720 196.580 64.860 196.735 ;
        RECT 71.070 196.720 71.390 196.780 ;
        RECT 62.330 196.440 64.860 196.580 ;
        RECT 65.130 196.580 65.420 196.625 ;
        RECT 67.230 196.580 67.520 196.625 ;
        RECT 68.800 196.580 69.090 196.625 ;
        RECT 65.130 196.440 69.090 196.580 ;
        RECT 62.330 196.380 62.650 196.440 ;
        RECT 65.130 196.395 65.420 196.440 ;
        RECT 67.230 196.395 67.520 196.440 ;
        RECT 68.800 196.395 69.090 196.440 ;
        RECT 71.530 196.580 71.850 196.640 ;
        RECT 72.540 196.580 72.680 196.780 ;
        RECT 89.025 196.735 89.315 196.780 ;
        RECT 89.470 196.720 89.790 196.780 ;
        RECT 95.910 196.720 96.230 196.780 ;
        RECT 96.830 196.920 97.150 196.980 ;
        RECT 97.840 196.920 97.980 197.075 ;
        RECT 98.670 197.060 98.990 197.120 ;
        RECT 96.830 196.780 97.980 196.920 ;
        RECT 96.830 196.720 97.150 196.780 ;
        RECT 71.530 196.440 72.680 196.580 ;
        RECT 72.925 196.580 73.215 196.625 ;
        RECT 74.750 196.580 75.070 196.640 ;
        RECT 72.925 196.440 75.070 196.580 ;
        RECT 71.530 196.380 71.850 196.440 ;
        RECT 72.925 196.395 73.215 196.440 ;
        RECT 74.750 196.380 75.070 196.440 ;
        RECT 76.130 196.380 76.450 196.640 ;
        RECT 94.085 196.580 94.375 196.625 ;
        RECT 90.940 196.440 94.375 196.580 ;
        RECT 53.130 196.240 53.450 196.300 ;
        RECT 51.380 196.100 53.450 196.240 ;
        RECT 43.025 196.055 43.315 196.100 ;
        RECT 48.070 196.040 48.390 196.100 ;
        RECT 53.130 196.040 53.450 196.100 ;
        RECT 59.110 196.040 59.430 196.300 ;
        RECT 60.505 196.240 60.795 196.285 ;
        RECT 61.500 196.240 61.640 196.380 ;
        RECT 60.505 196.100 61.640 196.240 ;
        RECT 71.070 196.240 71.390 196.300 ;
        RECT 75.210 196.240 75.530 196.300 ;
        RECT 71.070 196.100 75.530 196.240 ;
        RECT 60.505 196.055 60.795 196.100 ;
        RECT 71.070 196.040 71.390 196.100 ;
        RECT 75.210 196.040 75.530 196.100 ;
        RECT 76.590 196.240 76.910 196.300 ;
        RECT 77.985 196.240 78.275 196.285 ;
        RECT 76.590 196.100 78.275 196.240 ;
        RECT 76.590 196.040 76.910 196.100 ;
        RECT 77.985 196.055 78.275 196.100 ;
        RECT 78.890 196.040 79.210 196.300 ;
        RECT 86.250 196.040 86.570 196.300 ;
        RECT 90.940 196.285 91.080 196.440 ;
        RECT 94.085 196.395 94.375 196.440 ;
        RECT 98.685 196.580 98.975 196.625 ;
        RECT 99.220 196.580 99.360 197.400 ;
        RECT 104.280 197.320 104.420 197.460 ;
        RECT 101.445 197.075 101.735 197.305 ;
        RECT 103.745 197.260 104.035 197.305 ;
        RECT 104.190 197.260 104.510 197.320 ;
        RECT 105.110 197.305 105.430 197.320 ;
        RECT 105.080 197.260 105.430 197.305 ;
        RECT 103.745 197.120 104.510 197.260 ;
        RECT 104.915 197.120 105.430 197.260 ;
        RECT 103.745 197.075 104.035 197.120 ;
        RECT 98.685 196.440 99.360 196.580 ;
        RECT 98.685 196.395 98.975 196.440 ;
        RECT 90.865 196.055 91.155 196.285 ;
        RECT 91.310 196.240 91.630 196.300 ;
        RECT 91.785 196.240 92.075 196.285 ;
        RECT 91.310 196.100 92.075 196.240 ;
        RECT 91.310 196.040 91.630 196.100 ;
        RECT 91.785 196.055 92.075 196.100 ;
        RECT 95.450 196.240 95.770 196.300 ;
        RECT 95.925 196.240 96.215 196.285 ;
        RECT 95.450 196.100 96.215 196.240 ;
        RECT 101.520 196.240 101.660 197.075 ;
        RECT 104.190 197.060 104.510 197.120 ;
        RECT 105.080 197.075 105.430 197.120 ;
        RECT 105.110 197.060 105.430 197.075 ;
        RECT 107.870 197.260 108.190 197.320 ;
        RECT 111.565 197.260 111.855 197.305 ;
        RECT 107.870 197.120 111.855 197.260 ;
        RECT 107.870 197.060 108.190 197.120 ;
        RECT 111.565 197.075 111.855 197.120 ;
        RECT 112.010 197.060 112.330 197.320 ;
        RECT 113.480 197.305 113.620 197.460 ;
        RECT 130.885 197.460 144.530 197.600 ;
        RECT 130.885 197.415 131.175 197.460 ;
        RECT 144.210 197.400 144.530 197.460 ;
        RECT 113.405 197.075 113.695 197.305 ;
        RECT 113.850 197.260 114.170 197.320 ;
        RECT 114.685 197.260 114.975 197.305 ;
        RECT 113.850 197.120 114.975 197.260 ;
        RECT 113.850 197.060 114.170 197.120 ;
        RECT 114.685 197.075 114.975 197.120 ;
        RECT 116.610 197.260 116.930 197.320 ;
        RECT 126.745 197.260 127.035 197.305 ;
        RECT 131.330 197.260 131.650 197.320 ;
        RECT 116.610 197.120 131.650 197.260 ;
        RECT 116.610 197.060 116.930 197.120 ;
        RECT 126.745 197.075 127.035 197.120 ;
        RECT 131.330 197.060 131.650 197.120 ;
        RECT 132.265 197.075 132.555 197.305 ;
        RECT 133.185 197.260 133.475 197.305 ;
        RECT 134.550 197.260 134.870 197.320 ;
        RECT 133.185 197.120 134.870 197.260 ;
        RECT 133.185 197.075 133.475 197.120 ;
        RECT 104.625 196.920 104.915 196.965 ;
        RECT 105.815 196.920 106.105 196.965 ;
        RECT 108.335 196.920 108.625 196.965 ;
        RECT 104.625 196.780 108.625 196.920 ;
        RECT 104.625 196.735 104.915 196.780 ;
        RECT 105.815 196.735 106.105 196.780 ;
        RECT 108.335 196.735 108.625 196.780 ;
        RECT 114.285 196.920 114.575 196.965 ;
        RECT 115.475 196.920 115.765 196.965 ;
        RECT 117.995 196.920 118.285 196.965 ;
        RECT 114.285 196.780 118.285 196.920 ;
        RECT 114.285 196.735 114.575 196.780 ;
        RECT 115.475 196.735 115.765 196.780 ;
        RECT 117.995 196.735 118.285 196.780 ;
        RECT 118.450 196.920 118.770 196.980 ;
        RECT 120.765 196.920 121.055 196.965 ;
        RECT 118.450 196.780 121.055 196.920 ;
        RECT 118.450 196.720 118.770 196.780 ;
        RECT 120.765 196.735 121.055 196.780 ;
        RECT 123.525 196.920 123.815 196.965 ;
        RECT 128.110 196.920 128.430 196.980 ;
        RECT 132.340 196.920 132.480 197.075 ;
        RECT 134.550 197.060 134.870 197.120 ;
        RECT 136.850 197.060 137.170 197.320 ;
        RECT 137.785 197.260 138.075 197.305 ;
        RECT 138.230 197.260 138.550 197.320 ;
        RECT 137.785 197.120 138.550 197.260 ;
        RECT 137.785 197.075 138.075 197.120 ;
        RECT 138.230 197.060 138.550 197.120 ;
        RECT 140.085 197.260 140.375 197.305 ;
        RECT 141.450 197.260 141.770 197.320 ;
        RECT 140.085 197.120 141.770 197.260 ;
        RECT 140.085 197.075 140.375 197.120 ;
        RECT 141.450 197.060 141.770 197.120 ;
        RECT 146.970 197.060 147.290 197.320 ;
        RECT 147.905 197.075 148.195 197.305 ;
        RECT 123.525 196.780 132.480 196.920 ;
        RECT 145.130 196.920 145.450 196.980 ;
        RECT 147.980 196.920 148.120 197.075 ;
        RECT 145.130 196.780 148.120 196.920 ;
        RECT 123.525 196.735 123.815 196.780 ;
        RECT 104.230 196.580 104.520 196.625 ;
        RECT 106.330 196.580 106.620 196.625 ;
        RECT 107.900 196.580 108.190 196.625 ;
        RECT 104.230 196.440 108.190 196.580 ;
        RECT 104.230 196.395 104.520 196.440 ;
        RECT 106.330 196.395 106.620 196.440 ;
        RECT 107.900 196.395 108.190 196.440 ;
        RECT 113.890 196.580 114.180 196.625 ;
        RECT 115.990 196.580 116.280 196.625 ;
        RECT 117.560 196.580 117.850 196.625 ;
        RECT 113.890 196.440 117.850 196.580 ;
        RECT 113.890 196.395 114.180 196.440 ;
        RECT 115.990 196.395 116.280 196.440 ;
        RECT 117.560 196.395 117.850 196.440 ;
        RECT 120.305 196.580 120.595 196.625 ;
        RECT 123.600 196.580 123.740 196.735 ;
        RECT 128.110 196.720 128.430 196.780 ;
        RECT 145.130 196.720 145.450 196.780 ;
        RECT 131.790 196.580 132.110 196.640 ;
        RECT 120.305 196.440 123.740 196.580 ;
        RECT 130.270 196.440 132.110 196.580 ;
        RECT 120.305 196.395 120.595 196.440 ;
        RECT 103.730 196.240 104.050 196.300 ;
        RECT 109.250 196.240 109.570 196.300 ;
        RECT 110.645 196.240 110.935 196.285 ;
        RECT 101.520 196.100 110.935 196.240 ;
        RECT 95.450 196.040 95.770 196.100 ;
        RECT 95.925 196.055 96.215 196.100 ;
        RECT 103.730 196.040 104.050 196.100 ;
        RECT 109.250 196.040 109.570 196.100 ;
        RECT 110.645 196.055 110.935 196.100 ;
        RECT 114.770 196.240 115.090 196.300 ;
        RECT 130.270 196.240 130.410 196.440 ;
        RECT 131.790 196.380 132.110 196.440 ;
        RECT 114.770 196.100 130.410 196.240 ;
        RECT 114.770 196.040 115.090 196.100 ;
        RECT 131.330 196.040 131.650 196.300 ;
        RECT 22.700 195.420 157.020 195.900 ;
        RECT 37.045 195.220 37.335 195.265 ;
        RECT 37.950 195.220 38.270 195.280 ;
        RECT 37.045 195.080 38.270 195.220 ;
        RECT 37.045 195.035 37.335 195.080 ;
        RECT 37.950 195.020 38.270 195.080 ;
        RECT 50.370 195.020 50.690 195.280 ;
        RECT 53.590 195.220 53.910 195.280 ;
        RECT 54.525 195.220 54.815 195.265 ;
        RECT 53.590 195.080 54.815 195.220 ;
        RECT 53.590 195.020 53.910 195.080 ;
        RECT 54.525 195.035 54.815 195.080 ;
        RECT 60.490 195.020 60.810 195.280 ;
        RECT 69.690 195.020 70.010 195.280 ;
        RECT 70.610 195.020 70.930 195.280 ;
        RECT 84.870 195.020 85.190 195.280 ;
        RECT 86.710 195.220 87.030 195.280 ;
        RECT 88.565 195.220 88.855 195.265 ;
        RECT 86.710 195.080 88.855 195.220 ;
        RECT 86.710 195.020 87.030 195.080 ;
        RECT 88.565 195.035 88.855 195.080 ;
        RECT 89.470 195.020 89.790 195.280 ;
        RECT 89.945 195.220 90.235 195.265 ;
        RECT 93.150 195.220 93.470 195.280 ;
        RECT 89.945 195.080 93.470 195.220 ;
        RECT 89.945 195.035 90.235 195.080 ;
        RECT 72.465 194.880 72.755 194.925 ;
        RECT 74.750 194.880 75.070 194.940 ;
        RECT 72.465 194.740 75.070 194.880 ;
        RECT 72.465 194.695 72.755 194.740 ;
        RECT 74.750 194.680 75.070 194.740 ;
        RECT 75.670 194.680 75.990 194.940 ;
        RECT 77.090 194.880 77.380 194.925 ;
        RECT 79.190 194.880 79.480 194.925 ;
        RECT 80.760 194.880 81.050 194.925 ;
        RECT 77.090 194.740 81.050 194.880 ;
        RECT 77.090 194.695 77.380 194.740 ;
        RECT 79.190 194.695 79.480 194.740 ;
        RECT 80.760 194.695 81.050 194.740 ;
        RECT 71.530 194.540 71.850 194.600 ;
        RECT 71.530 194.400 74.980 194.540 ;
        RECT 71.530 194.340 71.850 194.400 ;
        RECT 36.110 194.000 36.430 194.260 ;
        RECT 40.265 194.200 40.555 194.245 ;
        RECT 40.710 194.200 41.030 194.260 ;
        RECT 40.265 194.060 41.030 194.200 ;
        RECT 40.265 194.015 40.555 194.060 ;
        RECT 40.710 194.000 41.030 194.060 ;
        RECT 46.690 194.200 47.010 194.260 ;
        RECT 47.625 194.200 47.915 194.245 ;
        RECT 46.690 194.060 47.915 194.200 ;
        RECT 46.690 194.000 47.010 194.060 ;
        RECT 47.625 194.015 47.915 194.060 ;
        RECT 48.530 194.200 48.850 194.260 ;
        RECT 49.005 194.200 49.295 194.245 ;
        RECT 48.530 194.060 49.295 194.200 ;
        RECT 48.530 194.000 48.850 194.060 ;
        RECT 49.005 194.015 49.295 194.060 ;
        RECT 52.225 194.200 52.515 194.245 ;
        RECT 54.050 194.200 54.370 194.260 ;
        RECT 52.225 194.060 54.370 194.200 ;
        RECT 52.225 194.015 52.515 194.060 ;
        RECT 54.050 194.000 54.370 194.060 ;
        RECT 55.445 194.200 55.735 194.245 ;
        RECT 57.270 194.200 57.590 194.260 ;
        RECT 55.445 194.060 57.590 194.200 ;
        RECT 55.445 194.015 55.735 194.060 ;
        RECT 57.270 194.000 57.590 194.060 ;
        RECT 58.205 194.015 58.495 194.245 ;
        RECT 59.110 194.200 59.430 194.260 ;
        RECT 59.585 194.200 59.875 194.245 ;
        RECT 61.870 194.200 62.190 194.260 ;
        RECT 68.325 194.200 68.615 194.245 ;
        RECT 59.110 194.060 61.640 194.200 ;
        RECT 33.825 193.675 34.115 193.905 ;
        RECT 34.745 193.860 35.035 193.905 ;
        RECT 35.650 193.860 35.970 193.920 ;
        RECT 34.745 193.720 35.970 193.860 ;
        RECT 34.745 193.675 35.035 193.720 ;
        RECT 32.905 193.520 33.195 193.565 ;
        RECT 33.350 193.520 33.670 193.580 ;
        RECT 32.905 193.380 33.670 193.520 ;
        RECT 33.900 193.520 34.040 193.675 ;
        RECT 35.650 193.660 35.970 193.720 ;
        RECT 48.085 193.860 48.375 193.905 ;
        RECT 50.830 193.860 51.150 193.920 ;
        RECT 48.085 193.720 51.150 193.860 ;
        RECT 48.085 193.675 48.375 193.720 ;
        RECT 50.830 193.660 51.150 193.720 ;
        RECT 53.130 193.860 53.450 193.920 ;
        RECT 58.280 193.860 58.420 194.015 ;
        RECT 59.110 194.000 59.430 194.060 ;
        RECT 59.585 194.015 59.875 194.060 ;
        RECT 53.130 193.720 58.420 193.860 ;
        RECT 58.665 193.860 58.955 193.905 ;
        RECT 60.030 193.860 60.350 193.920 ;
        RECT 58.665 193.720 60.350 193.860 ;
        RECT 61.500 193.860 61.640 194.060 ;
        RECT 61.870 194.060 68.615 194.200 ;
        RECT 61.870 194.000 62.190 194.060 ;
        RECT 68.325 194.015 68.615 194.060 ;
        RECT 70.150 194.200 70.470 194.260 ;
        RECT 73.845 194.200 74.135 194.245 ;
        RECT 70.150 194.060 74.135 194.200 ;
        RECT 70.150 194.000 70.470 194.060 ;
        RECT 73.845 194.015 74.135 194.060 ;
        RECT 74.290 194.000 74.610 194.260 ;
        RECT 74.840 194.245 74.980 194.400 ;
        RECT 76.590 194.340 76.910 194.600 ;
        RECT 86.800 194.585 86.940 195.020 ;
        RECT 77.485 194.540 77.775 194.585 ;
        RECT 78.675 194.540 78.965 194.585 ;
        RECT 81.195 194.540 81.485 194.585 ;
        RECT 77.485 194.400 81.485 194.540 ;
        RECT 77.485 194.355 77.775 194.400 ;
        RECT 78.675 194.355 78.965 194.400 ;
        RECT 81.195 194.355 81.485 194.400 ;
        RECT 86.725 194.355 87.015 194.585 ;
        RECT 74.765 194.015 75.055 194.245 ;
        RECT 76.130 194.200 76.450 194.260 ;
        RECT 85.330 194.200 85.650 194.260 ;
        RECT 85.805 194.200 86.095 194.245 ;
        RECT 75.300 194.060 86.095 194.200 ;
        RECT 62.330 193.860 62.650 193.920 ;
        RECT 61.500 193.720 62.650 193.860 ;
        RECT 53.130 193.660 53.450 193.720 ;
        RECT 58.665 193.675 58.955 193.720 ;
        RECT 60.030 193.660 60.350 193.720 ;
        RECT 62.330 193.660 62.650 193.720 ;
        RECT 64.630 193.860 64.950 193.920 ;
        RECT 71.530 193.860 71.850 193.920 ;
        RECT 64.630 193.720 71.850 193.860 ;
        RECT 64.630 193.660 64.950 193.720 ;
        RECT 71.530 193.660 71.850 193.720 ;
        RECT 72.925 193.860 73.215 193.905 ;
        RECT 75.300 193.860 75.440 194.060 ;
        RECT 76.130 194.000 76.450 194.060 ;
        RECT 85.330 194.000 85.650 194.060 ;
        RECT 85.805 194.015 86.095 194.060 ;
        RECT 77.970 193.905 78.290 193.920 ;
        RECT 72.925 193.720 75.440 193.860 ;
        RECT 72.925 193.675 73.215 193.720 ;
        RECT 77.940 193.675 78.290 193.905 ;
        RECT 77.970 193.660 78.290 193.675 ;
        RECT 34.270 193.520 34.590 193.580 ;
        RECT 36.570 193.520 36.890 193.580 ;
        RECT 33.900 193.380 36.890 193.520 ;
        RECT 32.905 193.335 33.195 193.380 ;
        RECT 33.350 193.320 33.670 193.380 ;
        RECT 34.270 193.320 34.590 193.380 ;
        RECT 36.570 193.320 36.890 193.380 ;
        RECT 39.330 193.320 39.650 193.580 ;
        RECT 49.450 193.520 49.770 193.580 ;
        RECT 51.305 193.520 51.595 193.565 ;
        RECT 49.450 193.380 51.595 193.520 ;
        RECT 49.450 193.320 49.770 193.380 ;
        RECT 51.305 193.335 51.595 193.380 ;
        RECT 53.590 193.320 53.910 193.580 ;
        RECT 62.790 193.520 63.110 193.580 ;
        RECT 70.625 193.520 70.915 193.565 ;
        RECT 77.510 193.520 77.830 193.580 ;
        RECT 62.790 193.380 77.830 193.520 ;
        RECT 62.790 193.320 63.110 193.380 ;
        RECT 70.625 193.335 70.915 193.380 ;
        RECT 77.510 193.320 77.830 193.380 ;
        RECT 83.490 193.320 83.810 193.580 ;
        RECT 85.880 193.520 86.020 194.015 ;
        RECT 87.645 193.860 87.935 193.905 ;
        RECT 88.090 193.860 88.410 193.920 ;
        RECT 90.020 193.860 90.160 195.035 ;
        RECT 93.150 195.020 93.470 195.080 ;
        RECT 112.010 195.020 112.330 195.280 ;
        RECT 113.405 195.220 113.695 195.265 ;
        RECT 113.850 195.220 114.170 195.280 ;
        RECT 113.405 195.080 114.170 195.220 ;
        RECT 113.405 195.035 113.695 195.080 ;
        RECT 113.850 195.020 114.170 195.080 ;
        RECT 120.290 195.220 120.610 195.280 ;
        RECT 121.225 195.220 121.515 195.265 ;
        RECT 120.290 195.080 121.515 195.220 ;
        RECT 120.290 195.020 120.610 195.080 ;
        RECT 121.225 195.035 121.515 195.080 ;
        RECT 125.365 195.220 125.655 195.265 ;
        RECT 126.270 195.220 126.590 195.280 ;
        RECT 125.365 195.080 126.590 195.220 ;
        RECT 125.365 195.035 125.655 195.080 ;
        RECT 126.270 195.020 126.590 195.080 ;
        RECT 128.110 195.020 128.430 195.280 ;
        RECT 130.410 195.220 130.730 195.280 ;
        RECT 133.170 195.220 133.490 195.280 ;
        RECT 130.410 195.080 133.490 195.220 ;
        RECT 130.410 195.020 130.730 195.080 ;
        RECT 133.170 195.020 133.490 195.080 ;
        RECT 140.085 195.220 140.375 195.265 ;
        RECT 140.990 195.220 141.310 195.280 ;
        RECT 140.085 195.080 141.310 195.220 ;
        RECT 140.085 195.035 140.375 195.080 ;
        RECT 140.990 195.020 141.310 195.080 ;
        RECT 141.450 195.020 141.770 195.280 ;
        RECT 142.385 195.035 142.675 195.265 ;
        RECT 92.690 194.880 92.980 194.925 ;
        RECT 94.260 194.880 94.550 194.925 ;
        RECT 96.360 194.880 96.650 194.925 ;
        RECT 92.690 194.740 96.650 194.880 ;
        RECT 92.690 194.695 92.980 194.740 ;
        RECT 94.260 194.695 94.550 194.740 ;
        RECT 96.360 194.695 96.650 194.740 ;
        RECT 101.930 194.880 102.220 194.925 ;
        RECT 104.030 194.880 104.320 194.925 ;
        RECT 105.600 194.880 105.890 194.925 ;
        RECT 101.930 194.740 105.890 194.880 ;
        RECT 101.930 194.695 102.220 194.740 ;
        RECT 104.030 194.695 104.320 194.740 ;
        RECT 105.600 194.695 105.890 194.740 ;
        RECT 108.345 194.695 108.635 194.925 ;
        RECT 124.430 194.880 124.750 194.940 ;
        RECT 130.870 194.880 131.190 194.940 ;
        RECT 124.430 194.740 127.420 194.880 ;
        RECT 92.255 194.540 92.545 194.585 ;
        RECT 94.775 194.540 95.065 194.585 ;
        RECT 95.965 194.540 96.255 194.585 ;
        RECT 92.255 194.400 96.255 194.540 ;
        RECT 92.255 194.355 92.545 194.400 ;
        RECT 94.775 194.355 95.065 194.400 ;
        RECT 95.965 194.355 96.255 194.400 ;
        RECT 96.845 194.540 97.135 194.585 ;
        RECT 102.325 194.540 102.615 194.585 ;
        RECT 103.515 194.540 103.805 194.585 ;
        RECT 106.035 194.540 106.325 194.585 ;
        RECT 96.845 194.400 101.660 194.540 ;
        RECT 96.845 194.355 97.135 194.400 ;
        RECT 98.210 194.000 98.530 194.260 ;
        RECT 101.520 194.245 101.660 194.400 ;
        RECT 102.325 194.400 106.325 194.540 ;
        RECT 108.420 194.540 108.560 194.695 ;
        RECT 124.430 194.680 124.750 194.740 ;
        RECT 127.280 194.585 127.420 194.740 ;
        RECT 127.740 194.740 131.190 194.880 ;
        RECT 108.805 194.540 109.095 194.585 ;
        RECT 108.420 194.400 109.095 194.540 ;
        RECT 102.325 194.355 102.615 194.400 ;
        RECT 103.515 194.355 103.805 194.400 ;
        RECT 106.035 194.355 106.325 194.400 ;
        RECT 108.805 194.355 109.095 194.400 ;
        RECT 123.065 194.540 123.355 194.585 ;
        RECT 126.745 194.540 127.035 194.585 ;
        RECT 123.065 194.400 127.035 194.540 ;
        RECT 123.065 194.355 123.355 194.400 ;
        RECT 126.745 194.355 127.035 194.400 ;
        RECT 127.205 194.355 127.495 194.585 ;
        RECT 101.445 194.200 101.735 194.245 ;
        RECT 104.190 194.200 104.510 194.260 ;
        RECT 105.110 194.200 105.430 194.260 ;
        RECT 101.445 194.060 105.430 194.200 ;
        RECT 101.445 194.015 101.735 194.060 ;
        RECT 104.190 194.000 104.510 194.060 ;
        RECT 105.110 194.000 105.430 194.060 ;
        RECT 112.010 194.200 112.330 194.260 ;
        RECT 114.310 194.200 114.630 194.260 ;
        RECT 112.010 194.060 114.630 194.200 ;
        RECT 112.010 194.000 112.330 194.060 ;
        RECT 114.310 194.000 114.630 194.060 ;
        RECT 114.770 194.000 115.090 194.260 ;
        RECT 115.245 194.200 115.535 194.245 ;
        RECT 115.690 194.200 116.010 194.260 ;
        RECT 115.245 194.060 116.010 194.200 ;
        RECT 115.245 194.015 115.535 194.060 ;
        RECT 87.645 193.720 90.160 193.860 ;
        RECT 92.230 193.860 92.550 193.920 ;
        RECT 95.510 193.860 95.800 193.905 ;
        RECT 92.230 193.720 95.800 193.860 ;
        RECT 87.645 193.675 87.935 193.720 ;
        RECT 88.090 193.660 88.410 193.720 ;
        RECT 92.230 193.660 92.550 193.720 ;
        RECT 95.510 193.675 95.800 193.720 ;
        RECT 100.985 193.860 101.275 193.905 ;
        RECT 102.670 193.860 102.960 193.905 ;
        RECT 100.985 193.720 102.960 193.860 ;
        RECT 100.985 193.675 101.275 193.720 ;
        RECT 102.670 193.675 102.960 193.720 ;
        RECT 111.550 193.860 111.870 193.920 ;
        RECT 115.320 193.860 115.460 194.015 ;
        RECT 115.690 194.000 116.010 194.060 ;
        RECT 116.165 194.200 116.455 194.245 ;
        RECT 118.450 194.200 118.770 194.260 ;
        RECT 116.165 194.060 118.770 194.200 ;
        RECT 116.165 194.015 116.455 194.060 ;
        RECT 118.450 194.000 118.770 194.060 ;
        RECT 120.765 194.200 121.055 194.245 ;
        RECT 121.670 194.200 121.990 194.260 ;
        RECT 120.765 194.060 121.990 194.200 ;
        RECT 120.765 194.015 121.055 194.060 ;
        RECT 121.670 194.000 121.990 194.060 ;
        RECT 123.985 194.200 124.275 194.245 ;
        RECT 123.985 194.060 126.500 194.200 ;
        RECT 123.985 194.015 124.275 194.060 ;
        RECT 126.360 193.920 126.500 194.060 ;
        RECT 111.550 193.720 115.460 193.860 ;
        RECT 111.550 193.660 111.870 193.720 ;
        RECT 124.430 193.660 124.750 193.920 ;
        RECT 125.365 193.675 125.655 193.905 ;
        RECT 88.645 193.520 88.935 193.565 ;
        RECT 85.880 193.380 88.935 193.520 ;
        RECT 125.440 193.520 125.580 193.675 ;
        RECT 126.270 193.660 126.590 193.920 ;
        RECT 127.190 193.520 127.510 193.580 ;
        RECT 127.740 193.520 127.880 194.740 ;
        RECT 130.870 194.680 131.190 194.740 ;
        RECT 137.770 194.880 138.090 194.940 ;
        RECT 142.460 194.880 142.600 195.035 ;
        RECT 137.770 194.740 142.600 194.880 ;
        RECT 137.770 194.680 138.090 194.740 ;
        RECT 134.550 194.540 134.870 194.600 ;
        RECT 130.270 194.400 134.870 194.540 ;
        RECT 128.585 194.200 128.875 194.245 ;
        RECT 130.270 194.200 130.410 194.400 ;
        RECT 134.550 194.340 134.870 194.400 ;
        RECT 135.485 194.540 135.775 194.585 ;
        RECT 142.830 194.540 143.150 194.600 ;
        RECT 135.485 194.400 143.150 194.540 ;
        RECT 135.485 194.355 135.775 194.400 ;
        RECT 142.830 194.340 143.150 194.400 ;
        RECT 128.585 194.060 130.410 194.200 ;
        RECT 128.585 194.015 128.875 194.060 ;
        RECT 130.885 194.015 131.175 194.245 ;
        RECT 131.805 194.200 132.095 194.245 ;
        RECT 133.630 194.200 133.950 194.260 ;
        RECT 131.805 194.060 133.950 194.200 ;
        RECT 131.805 194.015 132.095 194.060 ;
        RECT 130.960 193.860 131.100 194.015 ;
        RECT 133.630 194.000 133.950 194.060 ;
        RECT 135.010 194.000 135.330 194.260 ;
        RECT 135.945 194.200 136.235 194.245 ;
        RECT 137.770 194.200 138.090 194.260 ;
        RECT 135.945 194.060 138.090 194.200 ;
        RECT 135.945 194.015 136.235 194.060 ;
        RECT 137.770 194.000 138.090 194.060 ;
        RECT 138.245 194.200 138.535 194.245 ;
        RECT 138.245 194.060 141.680 194.200 ;
        RECT 138.245 194.015 138.535 194.060 ;
        RECT 133.170 193.860 133.490 193.920 ;
        RECT 130.960 193.720 133.490 193.860 ;
        RECT 133.170 193.660 133.490 193.720 ;
        RECT 136.405 193.860 136.695 193.905 ;
        RECT 136.850 193.860 137.170 193.920 ;
        RECT 136.405 193.720 137.170 193.860 ;
        RECT 136.405 193.675 136.695 193.720 ;
        RECT 136.850 193.660 137.170 193.720 ;
        RECT 137.325 193.860 137.615 193.905 ;
        RECT 138.690 193.860 139.010 193.920 ;
        RECT 139.925 193.860 140.215 193.905 ;
        RECT 137.325 193.720 138.000 193.860 ;
        RECT 137.325 193.675 137.615 193.720 ;
        RECT 125.440 193.380 127.880 193.520 ;
        RECT 130.870 193.520 131.190 193.580 ;
        RECT 131.345 193.520 131.635 193.565 ;
        RECT 130.870 193.380 131.635 193.520 ;
        RECT 137.860 193.520 138.000 193.720 ;
        RECT 138.690 193.720 140.215 193.860 ;
        RECT 138.690 193.660 139.010 193.720 ;
        RECT 139.925 193.675 140.215 193.720 ;
        RECT 140.990 193.660 141.310 193.920 ;
        RECT 141.540 193.860 141.680 194.060 ;
        RECT 145.590 194.000 145.910 194.260 ;
        RECT 142.225 193.860 142.515 193.905 ;
        RECT 141.540 193.720 142.515 193.860 ;
        RECT 142.225 193.675 142.515 193.720 ;
        RECT 143.305 193.860 143.595 193.905 ;
        RECT 145.130 193.860 145.450 193.920 ;
        RECT 143.305 193.720 145.450 193.860 ;
        RECT 143.305 193.675 143.595 193.720 ;
        RECT 145.130 193.660 145.450 193.720 ;
        RECT 138.230 193.520 138.550 193.580 ;
        RECT 137.860 193.380 138.550 193.520 ;
        RECT 88.645 193.335 88.935 193.380 ;
        RECT 127.190 193.320 127.510 193.380 ;
        RECT 130.870 193.320 131.190 193.380 ;
        RECT 131.345 193.335 131.635 193.380 ;
        RECT 138.230 193.320 138.550 193.380 ;
        RECT 139.150 193.320 139.470 193.580 ;
        RECT 146.510 193.320 146.830 193.580 ;
        RECT 22.700 192.700 157.820 193.180 ;
        RECT 34.285 192.500 34.575 192.545 ;
        RECT 36.110 192.500 36.430 192.560 ;
        RECT 34.285 192.360 36.430 192.500 ;
        RECT 34.285 192.315 34.575 192.360 ;
        RECT 36.110 192.300 36.430 192.360 ;
        RECT 50.370 192.500 50.690 192.560 ;
        RECT 51.765 192.500 52.055 192.545 ;
        RECT 54.510 192.500 54.830 192.560 ;
        RECT 50.370 192.360 54.830 192.500 ;
        RECT 50.370 192.300 50.690 192.360 ;
        RECT 51.765 192.315 52.055 192.360 ;
        RECT 54.510 192.300 54.830 192.360 ;
        RECT 60.030 192.500 60.350 192.560 ;
        RECT 60.030 192.360 63.020 192.500 ;
        RECT 60.030 192.300 60.350 192.360 ;
        RECT 33.365 191.975 33.655 192.205 ;
        RECT 38.840 192.160 39.130 192.205 ;
        RECT 39.330 192.160 39.650 192.220 ;
        RECT 38.840 192.020 39.650 192.160 ;
        RECT 38.840 191.975 39.130 192.020 ;
        RECT 29.210 191.820 29.530 191.880 ;
        RECT 33.440 191.820 33.580 191.975 ;
        RECT 39.330 191.960 39.650 192.020 ;
        RECT 46.245 192.160 46.535 192.205 ;
        RECT 48.530 192.160 48.850 192.220 ;
        RECT 54.050 192.160 54.370 192.220 ;
        RECT 62.880 192.205 63.020 192.360 ;
        RECT 77.970 192.300 78.290 192.560 ;
        RECT 92.230 192.300 92.550 192.560 ;
        RECT 98.210 192.500 98.530 192.560 ;
        RECT 101.905 192.500 102.195 192.545 ;
        RECT 126.730 192.500 127.050 192.560 ;
        RECT 137.325 192.500 137.615 192.545 ;
        RECT 137.770 192.500 138.090 192.560 ;
        RECT 98.210 192.360 102.195 192.500 ;
        RECT 98.210 192.300 98.530 192.360 ;
        RECT 101.905 192.315 102.195 192.360 ;
        RECT 108.420 192.360 127.050 192.500 ;
        RECT 46.245 192.020 48.850 192.160 ;
        RECT 46.245 191.975 46.535 192.020 ;
        RECT 48.530 191.960 48.850 192.020 ;
        RECT 49.080 192.020 54.370 192.160 ;
        RECT 29.210 191.680 33.580 191.820 ;
        RECT 35.665 191.820 35.955 191.865 ;
        RECT 36.110 191.820 36.430 191.880 ;
        RECT 35.665 191.680 36.430 191.820 ;
        RECT 29.210 191.620 29.530 191.680 ;
        RECT 35.665 191.635 35.955 191.680 ;
        RECT 36.110 191.620 36.430 191.680 ;
        RECT 37.505 191.820 37.795 191.865 ;
        RECT 37.950 191.820 38.270 191.880 ;
        RECT 37.505 191.680 38.270 191.820 ;
        RECT 37.505 191.635 37.795 191.680 ;
        RECT 37.950 191.620 38.270 191.680 ;
        RECT 46.690 191.620 47.010 191.880 ;
        RECT 47.165 191.820 47.455 191.865 ;
        RECT 49.080 191.820 49.220 192.020 ;
        RECT 54.050 191.960 54.370 192.020 ;
        RECT 62.805 191.975 63.095 192.205 ;
        RECT 75.670 192.160 75.990 192.220 ;
        RECT 83.490 192.160 83.810 192.220 ;
        RECT 75.670 192.020 83.810 192.160 ;
        RECT 75.670 191.960 75.990 192.020 ;
        RECT 47.165 191.680 49.220 191.820 ;
        RECT 47.165 191.635 47.455 191.680 ;
        RECT 49.450 191.620 49.770 191.880 ;
        RECT 50.830 191.820 51.150 191.880 ;
        RECT 51.305 191.820 51.595 191.865 ;
        RECT 50.830 191.680 51.595 191.820 ;
        RECT 50.830 191.620 51.150 191.680 ;
        RECT 51.305 191.635 51.595 191.680 ;
        RECT 54.970 191.820 55.290 191.880 ;
        RECT 57.330 191.820 57.620 191.865 ;
        RECT 54.970 191.680 57.620 191.820 ;
        RECT 54.970 191.620 55.290 191.680 ;
        RECT 57.330 191.635 57.620 191.680 ;
        RECT 73.385 191.820 73.675 191.865 ;
        RECT 74.290 191.820 74.610 191.880 ;
        RECT 73.385 191.680 74.610 191.820 ;
        RECT 73.385 191.635 73.675 191.680 ;
        RECT 74.290 191.620 74.610 191.680 ;
        RECT 78.890 191.620 79.210 191.880 ;
        RECT 80.360 191.865 80.500 192.020 ;
        RECT 83.490 191.960 83.810 192.020 ;
        RECT 102.365 192.160 102.655 192.205 ;
        RECT 103.730 192.160 104.050 192.220 ;
        RECT 107.870 192.160 108.190 192.220 ;
        RECT 102.365 192.020 108.190 192.160 ;
        RECT 102.365 191.975 102.655 192.020 ;
        RECT 103.730 191.960 104.050 192.020 ;
        RECT 107.870 191.960 108.190 192.020 ;
        RECT 80.285 191.635 80.575 191.865 ;
        RECT 85.805 191.820 86.095 191.865 ;
        RECT 86.710 191.820 87.030 191.880 ;
        RECT 85.805 191.680 87.030 191.820 ;
        RECT 85.805 191.635 86.095 191.680 ;
        RECT 86.710 191.620 87.030 191.680 ;
        RECT 88.090 191.820 88.410 191.880 ;
        RECT 88.565 191.820 88.855 191.865 ;
        RECT 88.090 191.680 88.855 191.820 ;
        RECT 88.090 191.620 88.410 191.680 ;
        RECT 88.565 191.635 88.855 191.680 ;
        RECT 91.310 191.620 91.630 191.880 ;
        RECT 94.545 191.820 94.835 191.865 ;
        RECT 95.450 191.820 95.770 191.880 ;
        RECT 94.545 191.680 95.770 191.820 ;
        RECT 94.545 191.635 94.835 191.680 ;
        RECT 95.450 191.620 95.770 191.680 ;
        RECT 97.290 191.820 97.610 191.880 ;
        RECT 98.225 191.820 98.515 191.865 ;
        RECT 97.290 191.680 98.515 191.820 ;
        RECT 97.290 191.620 97.610 191.680 ;
        RECT 98.225 191.635 98.515 191.680 ;
        RECT 99.130 191.820 99.450 191.880 ;
        RECT 100.525 191.820 100.815 191.865 ;
        RECT 99.130 191.680 100.815 191.820 ;
        RECT 99.130 191.620 99.450 191.680 ;
        RECT 100.525 191.635 100.815 191.680 ;
        RECT 102.825 191.820 103.115 191.865 ;
        RECT 103.270 191.820 103.590 191.880 ;
        RECT 108.420 191.820 108.560 192.360 ;
        RECT 126.730 192.300 127.050 192.360 ;
        RECT 127.740 192.360 128.340 192.500 ;
        RECT 127.205 192.160 127.495 192.205 ;
        RECT 109.340 192.020 113.620 192.160 ;
        RECT 102.825 191.680 103.590 191.820 ;
        RECT 102.825 191.635 103.115 191.680 ;
        RECT 103.270 191.620 103.590 191.680 ;
        RECT 103.820 191.680 108.560 191.820 ;
        RECT 35.190 191.480 35.510 191.540 ;
        RECT 30.220 191.340 35.510 191.480 ;
        RECT 30.220 191.200 30.360 191.340 ;
        RECT 35.190 191.280 35.510 191.340 ;
        RECT 36.570 191.280 36.890 191.540 ;
        RECT 38.385 191.480 38.675 191.525 ;
        RECT 39.575 191.480 39.865 191.525 ;
        RECT 42.095 191.480 42.385 191.525 ;
        RECT 38.385 191.340 42.385 191.480 ;
        RECT 38.385 191.295 38.675 191.340 ;
        RECT 39.575 191.295 39.865 191.340 ;
        RECT 42.095 191.295 42.385 191.340 ;
        RECT 48.070 191.480 48.390 191.540 ;
        RECT 49.925 191.480 50.215 191.525 ;
        RECT 48.070 191.340 50.215 191.480 ;
        RECT 48.070 191.280 48.390 191.340 ;
        RECT 49.925 191.295 50.215 191.340 ;
        RECT 54.075 191.480 54.365 191.525 ;
        RECT 56.595 191.480 56.885 191.525 ;
        RECT 57.785 191.480 58.075 191.525 ;
        RECT 54.075 191.340 58.075 191.480 ;
        RECT 54.075 191.295 54.365 191.340 ;
        RECT 56.595 191.295 56.885 191.340 ;
        RECT 57.785 191.295 58.075 191.340 ;
        RECT 58.665 191.480 58.955 191.525 ;
        RECT 61.870 191.480 62.190 191.540 ;
        RECT 58.665 191.340 62.190 191.480 ;
        RECT 58.665 191.295 58.955 191.340 ;
        RECT 61.870 191.280 62.190 191.340 ;
        RECT 62.330 191.480 62.650 191.540 ;
        RECT 67.865 191.480 68.155 191.525 ;
        RECT 62.330 191.340 68.155 191.480 ;
        RECT 62.330 191.280 62.650 191.340 ;
        RECT 67.865 191.295 68.155 191.340 ;
        RECT 68.770 191.480 69.090 191.540 ;
        RECT 103.820 191.480 103.960 191.680 ;
        RECT 108.790 191.620 109.110 191.880 ;
        RECT 109.340 191.865 109.480 192.020 ;
        RECT 113.480 191.880 113.620 192.020 ;
        RECT 126.360 192.020 127.495 192.160 ;
        RECT 109.265 191.635 109.555 191.865 ;
        RECT 109.710 191.820 110.030 191.880 ;
        RECT 110.545 191.820 110.835 191.865 ;
        RECT 109.710 191.680 110.835 191.820 ;
        RECT 109.710 191.620 110.030 191.680 ;
        RECT 110.545 191.635 110.835 191.680 ;
        RECT 113.390 191.820 113.710 191.880 ;
        RECT 116.610 191.820 116.930 191.880 ;
        RECT 113.390 191.680 116.930 191.820 ;
        RECT 113.390 191.620 113.710 191.680 ;
        RECT 116.610 191.620 116.930 191.680 ;
        RECT 117.070 191.820 117.390 191.880 ;
        RECT 117.905 191.820 118.195 191.865 ;
        RECT 117.070 191.680 118.195 191.820 ;
        RECT 117.070 191.620 117.390 191.680 ;
        RECT 117.905 191.635 118.195 191.680 ;
        RECT 68.770 191.340 103.960 191.480 ;
        RECT 68.770 191.280 69.090 191.340 ;
        RECT 105.110 191.280 105.430 191.540 ;
        RECT 110.145 191.480 110.435 191.525 ;
        RECT 111.335 191.480 111.625 191.525 ;
        RECT 113.855 191.480 114.145 191.525 ;
        RECT 110.145 191.340 114.145 191.480 ;
        RECT 110.145 191.295 110.435 191.340 ;
        RECT 111.335 191.295 111.625 191.340 ;
        RECT 113.855 191.295 114.145 191.340 ;
        RECT 117.505 191.480 117.795 191.525 ;
        RECT 118.695 191.480 118.985 191.525 ;
        RECT 121.215 191.480 121.505 191.525 ;
        RECT 117.505 191.340 121.505 191.480 ;
        RECT 126.360 191.480 126.500 192.020 ;
        RECT 127.205 191.975 127.495 192.020 ;
        RECT 126.745 191.820 127.035 191.865 ;
        RECT 127.740 191.820 127.880 192.360 ;
        RECT 128.200 192.160 128.340 192.360 ;
        RECT 137.325 192.360 138.090 192.500 ;
        RECT 137.325 192.315 137.615 192.360 ;
        RECT 137.770 192.300 138.090 192.360 ;
        RECT 140.990 192.500 141.310 192.560 ;
        RECT 144.225 192.500 144.515 192.545 ;
        RECT 140.990 192.360 144.515 192.500 ;
        RECT 140.990 192.300 141.310 192.360 ;
        RECT 144.225 192.315 144.515 192.360 ;
        RECT 130.410 192.160 130.730 192.220 ;
        RECT 131.805 192.160 132.095 192.205 ;
        RECT 138.230 192.160 138.550 192.220 ;
        RECT 140.530 192.160 140.850 192.220 ;
        RECT 128.200 192.020 132.095 192.160 ;
        RECT 130.410 191.960 130.730 192.020 ;
        RECT 131.805 191.975 132.095 192.020 ;
        RECT 136.940 192.020 140.850 192.160 ;
        RECT 126.745 191.680 127.880 191.820 ;
        RECT 126.745 191.635 127.035 191.680 ;
        RECT 128.125 191.635 128.415 191.865 ;
        RECT 129.505 191.820 129.795 191.865 ;
        RECT 130.870 191.820 131.190 191.880 ;
        RECT 129.505 191.680 131.190 191.820 ;
        RECT 129.505 191.635 129.795 191.680 ;
        RECT 127.650 191.480 127.970 191.540 ;
        RECT 126.360 191.340 127.970 191.480 ;
        RECT 128.200 191.480 128.340 191.635 ;
        RECT 130.870 191.620 131.190 191.680 ;
        RECT 133.170 191.620 133.490 191.880 ;
        RECT 133.630 191.620 133.950 191.880 ;
        RECT 134.090 191.620 134.410 191.880 ;
        RECT 135.010 191.620 135.330 191.880 ;
        RECT 136.940 191.865 137.080 192.020 ;
        RECT 138.230 191.960 138.550 192.020 ;
        RECT 140.530 191.960 140.850 192.020 ;
        RECT 136.865 191.635 137.155 191.865 ;
        RECT 137.310 191.820 137.630 191.880 ;
        RECT 137.785 191.820 138.075 191.865 ;
        RECT 137.310 191.680 138.075 191.820 ;
        RECT 137.310 191.620 137.630 191.680 ;
        RECT 137.785 191.635 138.075 191.680 ;
        RECT 139.165 191.820 139.455 191.865 ;
        RECT 141.080 191.820 141.220 192.300 ;
        RECT 142.845 192.160 143.135 192.205 ;
        RECT 145.130 192.160 145.450 192.220 ;
        RECT 142.845 192.020 145.450 192.160 ;
        RECT 142.845 191.975 143.135 192.020 ;
        RECT 145.130 191.960 145.450 192.020 ;
        RECT 146.510 192.160 146.830 192.220 ;
        RECT 149.790 192.160 150.080 192.205 ;
        RECT 146.510 192.020 150.080 192.160 ;
        RECT 146.510 191.960 146.830 192.020 ;
        RECT 149.790 191.975 150.080 192.020 ;
        RECT 139.165 191.680 141.220 191.820 ;
        RECT 150.650 191.820 150.970 191.880 ;
        RECT 151.125 191.820 151.415 191.865 ;
        RECT 150.650 191.680 151.415 191.820 ;
        RECT 139.165 191.635 139.455 191.680 ;
        RECT 150.650 191.620 150.970 191.680 ;
        RECT 151.125 191.635 151.415 191.680 ;
        RECT 129.965 191.480 130.255 191.525 ;
        RECT 128.200 191.340 130.255 191.480 ;
        RECT 135.100 191.480 135.240 191.620 ;
        RECT 138.705 191.480 138.995 191.525 ;
        RECT 135.100 191.340 138.995 191.480 ;
        RECT 117.505 191.295 117.795 191.340 ;
        RECT 118.695 191.295 118.985 191.340 ;
        RECT 121.215 191.295 121.505 191.340 ;
        RECT 127.650 191.280 127.970 191.340 ;
        RECT 129.965 191.295 130.255 191.340 ;
        RECT 138.705 191.295 138.995 191.340 ;
        RECT 146.535 191.480 146.825 191.525 ;
        RECT 149.055 191.480 149.345 191.525 ;
        RECT 150.245 191.480 150.535 191.525 ;
        RECT 146.535 191.340 150.535 191.480 ;
        RECT 146.535 191.295 146.825 191.340 ;
        RECT 149.055 191.295 149.345 191.340 ;
        RECT 150.245 191.295 150.535 191.340 ;
        RECT 30.130 190.940 30.450 191.200 ;
        RECT 31.525 191.140 31.815 191.185 ;
        RECT 37.990 191.140 38.280 191.185 ;
        RECT 40.090 191.140 40.380 191.185 ;
        RECT 41.660 191.140 41.950 191.185 ;
        RECT 31.525 191.000 34.960 191.140 ;
        RECT 31.525 190.955 31.815 191.000 ;
        RECT 33.350 190.600 33.670 190.860 ;
        RECT 34.820 190.845 34.960 191.000 ;
        RECT 37.990 191.000 41.950 191.140 ;
        RECT 37.990 190.955 38.280 191.000 ;
        RECT 40.090 190.955 40.380 191.000 ;
        RECT 41.660 190.955 41.950 191.000 ;
        RECT 45.325 190.955 45.615 191.185 ;
        RECT 54.510 191.140 54.800 191.185 ;
        RECT 56.080 191.140 56.370 191.185 ;
        RECT 58.180 191.140 58.470 191.185 ;
        RECT 54.510 191.000 58.470 191.140 ;
        RECT 54.510 190.955 54.800 191.000 ;
        RECT 56.080 190.955 56.370 191.000 ;
        RECT 58.180 190.955 58.470 191.000 ;
        RECT 64.645 191.140 64.935 191.185 ;
        RECT 64.645 191.000 66.240 191.140 ;
        RECT 64.645 190.955 64.935 191.000 ;
        RECT 34.745 190.800 35.035 190.845 ;
        RECT 35.650 190.800 35.970 190.860 ;
        RECT 34.745 190.660 35.970 190.800 ;
        RECT 34.745 190.615 35.035 190.660 ;
        RECT 35.650 190.600 35.970 190.660 ;
        RECT 44.390 190.800 44.710 190.860 ;
        RECT 45.400 190.800 45.540 190.955 ;
        RECT 44.390 190.660 45.540 190.800 ;
        RECT 45.770 190.800 46.090 190.860 ;
        RECT 48.085 190.800 48.375 190.845 ;
        RECT 45.770 190.660 48.375 190.800 ;
        RECT 44.390 190.600 44.710 190.660 ;
        RECT 45.770 190.600 46.090 190.660 ;
        RECT 48.085 190.615 48.375 190.660 ;
        RECT 48.990 190.600 49.310 190.860 ;
        RECT 50.830 190.600 51.150 190.860 ;
        RECT 65.090 190.600 65.410 190.860 ;
        RECT 65.550 190.600 65.870 190.860 ;
        RECT 66.100 190.800 66.240 191.000 ;
        RECT 66.470 190.940 66.790 191.200 ;
        RECT 104.190 191.140 104.510 191.200 ;
        RECT 105.570 191.140 105.890 191.200 ;
        RECT 104.190 191.000 105.890 191.140 ;
        RECT 104.190 190.940 104.510 191.000 ;
        RECT 105.570 190.940 105.890 191.000 ;
        RECT 109.750 191.140 110.040 191.185 ;
        RECT 111.850 191.140 112.140 191.185 ;
        RECT 113.420 191.140 113.710 191.185 ;
        RECT 109.750 191.000 113.710 191.140 ;
        RECT 109.750 190.955 110.040 191.000 ;
        RECT 111.850 190.955 112.140 191.000 ;
        RECT 113.420 190.955 113.710 191.000 ;
        RECT 117.110 191.140 117.400 191.185 ;
        RECT 119.210 191.140 119.500 191.185 ;
        RECT 120.780 191.140 121.070 191.185 ;
        RECT 117.110 191.000 121.070 191.140 ;
        RECT 117.110 190.955 117.400 191.000 ;
        RECT 119.210 190.955 119.500 191.000 ;
        RECT 120.780 190.955 121.070 191.000 ;
        RECT 125.810 191.140 126.130 191.200 ;
        RECT 125.810 191.000 128.800 191.140 ;
        RECT 125.810 190.940 126.130 191.000 ;
        RECT 69.230 190.800 69.550 190.860 ;
        RECT 66.100 190.660 69.550 190.800 ;
        RECT 69.230 190.600 69.550 190.660 ;
        RECT 72.925 190.800 73.215 190.845 ;
        RECT 74.290 190.800 74.610 190.860 ;
        RECT 72.925 190.660 74.610 190.800 ;
        RECT 72.925 190.615 73.215 190.660 ;
        RECT 74.290 190.600 74.610 190.660 ;
        RECT 79.810 190.600 80.130 190.860 ;
        RECT 84.870 190.800 85.190 190.860 ;
        RECT 85.345 190.800 85.635 190.845 ;
        RECT 84.870 190.660 85.635 190.800 ;
        RECT 84.870 190.600 85.190 190.660 ;
        RECT 85.345 190.615 85.635 190.660 ;
        RECT 88.105 190.800 88.395 190.845 ;
        RECT 89.010 190.800 89.330 190.860 ;
        RECT 88.105 190.660 89.330 190.800 ;
        RECT 88.105 190.615 88.395 190.660 ;
        RECT 89.010 190.600 89.330 190.660 ;
        RECT 94.085 190.800 94.375 190.845 ;
        RECT 94.530 190.800 94.850 190.860 ;
        RECT 94.085 190.660 94.850 190.800 ;
        RECT 94.085 190.615 94.375 190.660 ;
        RECT 94.530 190.600 94.850 190.660 ;
        RECT 97.765 190.800 98.055 190.845 ;
        RECT 98.210 190.800 98.530 190.860 ;
        RECT 97.765 190.660 98.530 190.800 ;
        RECT 97.765 190.615 98.055 190.660 ;
        RECT 98.210 190.600 98.530 190.660 ;
        RECT 116.150 190.600 116.470 190.860 ;
        RECT 123.510 190.600 123.830 190.860 ;
        RECT 127.650 190.800 127.970 190.860 ;
        RECT 128.660 190.845 128.800 191.000 ;
        RECT 128.125 190.800 128.415 190.845 ;
        RECT 127.650 190.660 128.415 190.800 ;
        RECT 127.650 190.600 127.970 190.660 ;
        RECT 128.125 190.615 128.415 190.660 ;
        RECT 128.585 190.615 128.875 190.845 ;
        RECT 130.040 190.800 130.180 191.295 ;
        RECT 132.265 191.140 132.555 191.185 ;
        RECT 130.960 191.000 132.555 191.140 ;
        RECT 130.960 190.800 131.100 191.000 ;
        RECT 132.265 190.955 132.555 191.000 ;
        RECT 139.150 191.140 139.470 191.200 ;
        RECT 141.005 191.140 141.295 191.185 ;
        RECT 139.150 191.000 141.295 191.140 ;
        RECT 139.150 190.940 139.470 191.000 ;
        RECT 141.005 190.955 141.295 191.000 ;
        RECT 143.765 191.140 144.055 191.185 ;
        RECT 145.590 191.140 145.910 191.200 ;
        RECT 143.765 191.000 145.910 191.140 ;
        RECT 143.765 190.955 144.055 191.000 ;
        RECT 145.590 190.940 145.910 191.000 ;
        RECT 146.970 191.140 147.260 191.185 ;
        RECT 148.540 191.140 148.830 191.185 ;
        RECT 150.640 191.140 150.930 191.185 ;
        RECT 146.970 191.000 150.930 191.140 ;
        RECT 146.970 190.955 147.260 191.000 ;
        RECT 148.540 190.955 148.830 191.000 ;
        RECT 150.640 190.955 150.930 191.000 ;
        RECT 130.040 190.660 131.100 190.800 ;
        RECT 131.330 190.600 131.650 190.860 ;
        RECT 142.830 190.600 143.150 190.860 ;
        RECT 22.700 189.980 157.020 190.460 ;
        RECT 32.445 189.780 32.735 189.825 ;
        RECT 33.810 189.780 34.130 189.840 ;
        RECT 32.445 189.640 34.130 189.780 ;
        RECT 32.445 189.595 32.735 189.640 ;
        RECT 33.810 189.580 34.130 189.640 ;
        RECT 39.805 189.595 40.095 189.825 ;
        RECT 24.650 189.440 24.940 189.485 ;
        RECT 26.750 189.440 27.040 189.485 ;
        RECT 28.320 189.440 28.610 189.485 ;
        RECT 24.650 189.300 28.610 189.440 ;
        RECT 39.880 189.440 40.020 189.595 ;
        RECT 40.710 189.580 41.030 189.840 ;
        RECT 48.070 189.580 48.390 189.840 ;
        RECT 48.530 189.780 48.850 189.840 ;
        RECT 49.005 189.780 49.295 189.825 ;
        RECT 57.745 189.780 58.035 189.825 ;
        RECT 48.530 189.640 49.295 189.780 ;
        RECT 48.530 189.580 48.850 189.640 ;
        RECT 49.005 189.595 49.295 189.640 ;
        RECT 53.220 189.640 58.035 189.780 ;
        RECT 42.565 189.440 42.855 189.485 ;
        RECT 45.770 189.440 46.090 189.500 ;
        RECT 39.880 189.300 42.855 189.440 ;
        RECT 24.650 189.255 24.940 189.300 ;
        RECT 26.750 189.255 27.040 189.300 ;
        RECT 28.320 189.255 28.610 189.300 ;
        RECT 42.565 189.255 42.855 189.300 ;
        RECT 43.100 189.300 46.090 189.440 ;
        RECT 25.045 189.100 25.335 189.145 ;
        RECT 26.235 189.100 26.525 189.145 ;
        RECT 28.755 189.100 29.045 189.145 ;
        RECT 25.045 188.960 29.045 189.100 ;
        RECT 25.045 188.915 25.335 188.960 ;
        RECT 26.235 188.915 26.525 188.960 ;
        RECT 28.755 188.915 29.045 188.960 ;
        RECT 35.190 189.100 35.510 189.160 ;
        RECT 36.110 189.100 36.430 189.160 ;
        RECT 37.965 189.100 38.255 189.145 ;
        RECT 43.100 189.100 43.240 189.300 ;
        RECT 45.770 189.240 46.090 189.300 ;
        RECT 35.190 188.960 43.240 189.100 ;
        RECT 43.945 189.100 44.235 189.145 ;
        RECT 46.690 189.100 47.010 189.160 ;
        RECT 43.945 188.960 47.010 189.100 ;
        RECT 35.190 188.900 35.510 188.960 ;
        RECT 36.110 188.900 36.430 188.960 ;
        RECT 37.965 188.915 38.255 188.960 ;
        RECT 43.945 188.915 44.235 188.960 ;
        RECT 46.690 188.900 47.010 188.960 ;
        RECT 24.150 188.560 24.470 188.820 ;
        RECT 31.970 188.760 32.290 188.820 ;
        RECT 34.285 188.760 34.575 188.805 ;
        RECT 31.970 188.620 34.575 188.760 ;
        RECT 31.970 188.560 32.290 188.620 ;
        RECT 34.285 188.575 34.575 188.620 ;
        RECT 43.485 188.575 43.775 188.805 ;
        RECT 44.405 188.575 44.695 188.805 ;
        RECT 25.530 188.465 25.850 188.480 ;
        RECT 25.500 188.235 25.850 188.465 ;
        RECT 25.530 188.220 25.850 188.235 ;
        RECT 27.370 188.420 27.690 188.480 ;
        RECT 29.210 188.420 29.530 188.480 ;
        RECT 32.445 188.420 32.735 188.465 ;
        RECT 39.805 188.420 40.095 188.465 ;
        RECT 27.370 188.280 40.095 188.420 ;
        RECT 27.370 188.220 27.690 188.280 ;
        RECT 29.210 188.220 29.530 188.280 ;
        RECT 32.445 188.235 32.735 188.280 ;
        RECT 39.805 188.235 40.095 188.280 ;
        RECT 31.050 187.880 31.370 188.140 ;
        RECT 31.510 187.880 31.830 188.140 ;
        RECT 43.560 188.080 43.700 188.575 ;
        RECT 44.480 188.420 44.620 188.575 ;
        RECT 44.850 188.560 45.170 188.820 ;
        RECT 48.620 188.760 48.760 189.580 ;
        RECT 53.220 189.440 53.360 189.640 ;
        RECT 57.745 189.595 58.035 189.640 ;
        RECT 63.725 189.780 64.015 189.825 ;
        RECT 66.470 189.780 66.790 189.840 ;
        RECT 70.150 189.780 70.470 189.840 ;
        RECT 63.725 189.640 70.470 189.780 ;
        RECT 63.725 189.595 64.015 189.640 ;
        RECT 66.470 189.580 66.790 189.640 ;
        RECT 70.150 189.580 70.470 189.640 ;
        RECT 92.705 189.780 92.995 189.825 ;
        RECT 101.430 189.780 101.750 189.840 ;
        RECT 92.705 189.640 101.750 189.780 ;
        RECT 92.705 189.595 92.995 189.640 ;
        RECT 101.430 189.580 101.750 189.640 ;
        RECT 108.805 189.780 109.095 189.825 ;
        RECT 109.710 189.780 110.030 189.840 ;
        RECT 108.805 189.640 110.030 189.780 ;
        RECT 108.805 189.595 109.095 189.640 ;
        RECT 109.710 189.580 110.030 189.640 ;
        RECT 112.485 189.780 112.775 189.825 ;
        RECT 117.070 189.780 117.390 189.840 ;
        RECT 112.485 189.640 117.390 189.780 ;
        RECT 112.485 189.595 112.775 189.640 ;
        RECT 117.070 189.580 117.390 189.640 ;
        RECT 127.190 189.580 127.510 189.840 ;
        RECT 129.045 189.780 129.335 189.825 ;
        RECT 130.410 189.780 130.730 189.840 ;
        RECT 129.045 189.640 130.730 189.780 ;
        RECT 129.045 189.595 129.335 189.640 ;
        RECT 130.410 189.580 130.730 189.640 ;
        RECT 133.630 189.780 133.950 189.840 ;
        RECT 135.945 189.780 136.235 189.825 ;
        RECT 133.630 189.640 136.235 189.780 ;
        RECT 133.630 189.580 133.950 189.640 ;
        RECT 135.945 189.595 136.235 189.640 ;
        RECT 141.005 189.780 141.295 189.825 ;
        RECT 145.605 189.780 145.895 189.825 ;
        RECT 141.005 189.640 145.895 189.780 ;
        RECT 141.005 189.595 141.295 189.640 ;
        RECT 145.605 189.595 145.895 189.640 ;
        RECT 51.380 189.300 53.360 189.440 ;
        RECT 51.380 189.100 51.520 189.300 ;
        RECT 65.550 189.240 65.870 189.500 ;
        RECT 71.545 189.255 71.835 189.485 ;
        RECT 95.465 189.440 95.755 189.485 ;
        RECT 97.750 189.440 98.070 189.500 ;
        RECT 111.550 189.440 111.870 189.500 ;
        RECT 128.125 189.440 128.415 189.485 ;
        RECT 132.250 189.440 132.570 189.500 ;
        RECT 95.465 189.300 98.070 189.440 ;
        RECT 95.465 189.255 95.755 189.300 ;
        RECT 50.920 188.960 51.520 189.100 ;
        RECT 51.750 189.100 52.070 189.160 ;
        RECT 51.750 188.960 52.900 189.100 ;
        RECT 45.400 188.620 48.760 188.760 ;
        RECT 45.400 188.420 45.540 188.620 ;
        RECT 50.370 188.560 50.690 188.820 ;
        RECT 50.920 188.805 51.060 188.960 ;
        RECT 51.750 188.900 52.070 188.960 ;
        RECT 52.760 188.805 52.900 188.960 ;
        RECT 54.510 188.900 54.830 189.160 ;
        RECT 65.640 189.100 65.780 189.240 ;
        RECT 65.180 188.960 65.780 189.100 ;
        RECT 50.845 188.575 51.135 188.805 ;
        RECT 52.225 188.760 52.515 188.805 ;
        RECT 51.380 188.620 52.515 188.760 ;
        RECT 44.480 188.280 45.540 188.420 ;
        RECT 48.530 188.420 48.850 188.480 ;
        RECT 51.380 188.420 51.520 188.620 ;
        RECT 52.225 188.575 52.515 188.620 ;
        RECT 52.685 188.575 52.975 188.805 ;
        RECT 60.490 188.560 60.810 188.820 ;
        RECT 62.330 188.560 62.650 188.820 ;
        RECT 65.180 188.805 65.320 188.960 ;
        RECT 65.105 188.575 65.395 188.805 ;
        RECT 65.550 188.760 65.870 188.820 ;
        RECT 67.635 188.760 67.925 188.805 ;
        RECT 65.550 188.620 66.065 188.760 ;
        RECT 67.635 188.620 68.540 188.760 ;
        RECT 65.550 188.560 65.870 188.620 ;
        RECT 67.635 188.575 67.925 188.620 ;
        RECT 48.530 188.280 51.520 188.420 ;
        RECT 51.765 188.420 52.055 188.465 ;
        RECT 54.510 188.420 54.830 188.480 ;
        RECT 51.765 188.280 54.830 188.420 ;
        RECT 48.530 188.220 48.850 188.280 ;
        RECT 51.765 188.235 52.055 188.280 ;
        RECT 54.510 188.220 54.830 188.280 ;
        RECT 66.485 188.235 66.775 188.465 ;
        RECT 47.610 188.080 47.930 188.140 ;
        RECT 49.450 188.080 49.770 188.140 ;
        RECT 43.560 187.940 49.770 188.080 ;
        RECT 47.610 187.880 47.930 187.940 ;
        RECT 49.450 187.880 49.770 187.940 ;
        RECT 50.370 188.080 50.690 188.140 ;
        RECT 51.290 188.080 51.610 188.140 ;
        RECT 50.370 187.940 51.610 188.080 ;
        RECT 50.370 187.880 50.690 187.940 ;
        RECT 51.290 187.880 51.610 187.940 ;
        RECT 53.605 188.080 53.895 188.125 ;
        RECT 54.050 188.080 54.370 188.140 ;
        RECT 53.605 187.940 54.370 188.080 ;
        RECT 53.605 187.895 53.895 187.940 ;
        RECT 54.050 187.880 54.370 187.940 ;
        RECT 57.270 187.880 57.590 188.140 ;
        RECT 64.645 188.080 64.935 188.125 ;
        RECT 66.560 188.080 66.700 188.235 ;
        RECT 66.930 188.220 67.250 188.480 ;
        RECT 68.400 188.420 68.540 188.620 ;
        RECT 68.770 188.560 69.090 188.820 ;
        RECT 70.165 188.760 70.455 188.805 ;
        RECT 71.620 188.760 71.760 189.255 ;
        RECT 97.750 189.240 98.070 189.300 ;
        RECT 107.040 189.300 111.870 189.440 ;
        RECT 78.445 189.100 78.735 189.145 ;
        RECT 83.950 189.100 84.270 189.160 ;
        RECT 78.445 188.960 84.270 189.100 ;
        RECT 78.445 188.915 78.735 188.960 ;
        RECT 70.165 188.620 71.760 188.760 ;
        RECT 70.165 188.575 70.455 188.620 ;
        RECT 72.450 188.560 72.770 188.820 ;
        RECT 72.925 188.760 73.215 188.805 ;
        RECT 73.830 188.760 74.150 188.820 ;
        RECT 72.925 188.620 74.150 188.760 ;
        RECT 72.925 188.575 73.215 188.620 ;
        RECT 73.830 188.560 74.150 188.620 ;
        RECT 74.305 188.760 74.595 188.805 ;
        RECT 75.210 188.760 75.530 188.820 ;
        RECT 74.305 188.620 75.530 188.760 ;
        RECT 74.305 188.575 74.595 188.620 ;
        RECT 75.210 188.560 75.530 188.620 ;
        RECT 75.670 188.760 75.990 188.820 ;
        RECT 77.065 188.760 77.355 188.805 ;
        RECT 75.670 188.620 77.355 188.760 ;
        RECT 75.670 188.560 75.990 188.620 ;
        RECT 77.065 188.575 77.355 188.620 ;
        RECT 77.525 188.575 77.815 188.805 ;
        RECT 78.905 188.760 79.195 188.805 ;
        RECT 79.810 188.760 80.130 188.820 ;
        RECT 80.820 188.805 80.960 188.960 ;
        RECT 83.950 188.900 84.270 188.960 ;
        RECT 85.805 188.915 86.095 189.145 ;
        RECT 104.650 189.100 104.970 189.160 ;
        RECT 86.340 188.960 89.240 189.100 ;
        RECT 78.905 188.620 80.130 188.760 ;
        RECT 78.905 188.575 79.195 188.620 ;
        RECT 70.610 188.420 70.930 188.480 ;
        RECT 68.400 188.280 70.930 188.420 ;
        RECT 70.610 188.220 70.930 188.280 ;
        RECT 73.385 188.235 73.675 188.465 ;
        RECT 75.300 188.420 75.440 188.560 ;
        RECT 77.600 188.420 77.740 188.575 ;
        RECT 79.810 188.560 80.130 188.620 ;
        RECT 80.745 188.575 81.035 188.805 ;
        RECT 81.665 188.760 81.955 188.805 ;
        RECT 84.410 188.760 84.730 188.820 ;
        RECT 81.665 188.620 84.730 188.760 ;
        RECT 81.665 188.575 81.955 188.620 ;
        RECT 84.410 188.560 84.730 188.620 ;
        RECT 84.870 188.560 85.190 188.820 ;
        RECT 75.300 188.280 77.740 188.420 ;
        RECT 81.205 188.420 81.495 188.465 ;
        RECT 84.960 188.420 85.100 188.560 ;
        RECT 81.205 188.280 85.100 188.420 ;
        RECT 85.880 188.420 86.020 188.915 ;
        RECT 86.340 188.805 86.480 188.960 ;
        RECT 89.100 188.820 89.240 188.960 ;
        RECT 90.480 188.960 94.760 189.100 ;
        RECT 86.265 188.575 86.555 188.805 ;
        RECT 88.565 188.575 88.855 188.805 ;
        RECT 86.710 188.420 87.030 188.480 ;
        RECT 88.640 188.420 88.780 188.575 ;
        RECT 89.010 188.560 89.330 188.820 ;
        RECT 90.480 188.805 90.620 188.960 ;
        RECT 94.620 188.820 94.760 188.960 ;
        RECT 96.000 188.960 98.440 189.100 ;
        RECT 90.405 188.575 90.695 188.805 ;
        RECT 91.310 188.560 91.630 188.820 ;
        RECT 94.070 188.760 94.390 188.820 ;
        RECT 92.320 188.620 94.390 188.760 ;
        RECT 85.880 188.280 88.780 188.420 ;
        RECT 89.485 188.420 89.775 188.465 ;
        RECT 92.320 188.420 92.460 188.620 ;
        RECT 94.070 188.560 94.390 188.620 ;
        RECT 94.530 188.560 94.850 188.820 ;
        RECT 96.000 188.805 96.140 188.960 ;
        RECT 98.300 188.820 98.440 188.960 ;
        RECT 104.650 188.960 106.720 189.100 ;
        RECT 104.650 188.900 104.970 188.960 ;
        RECT 95.925 188.575 96.215 188.805 ;
        RECT 97.750 188.560 98.070 188.820 ;
        RECT 98.210 188.560 98.530 188.820 ;
        RECT 99.130 188.560 99.450 188.820 ;
        RECT 99.605 188.760 99.895 188.805 ;
        RECT 105.570 188.760 105.890 188.820 ;
        RECT 99.605 188.620 105.890 188.760 ;
        RECT 99.605 188.575 99.895 188.620 ;
        RECT 105.570 188.560 105.890 188.620 ;
        RECT 106.045 188.575 106.335 188.805 ;
        RECT 89.485 188.280 92.460 188.420 ;
        RECT 92.705 188.420 92.995 188.465 ;
        RECT 96.845 188.420 97.135 188.465 ;
        RECT 92.705 188.280 97.135 188.420 ;
        RECT 81.205 188.235 81.495 188.280 ;
        RECT 64.645 187.940 66.700 188.080 ;
        RECT 68.325 188.080 68.615 188.125 ;
        RECT 69.245 188.080 69.535 188.125 ;
        RECT 68.325 187.940 69.535 188.080 ;
        RECT 64.645 187.895 64.935 187.940 ;
        RECT 68.325 187.895 68.615 187.940 ;
        RECT 69.245 187.895 69.535 187.940 ;
        RECT 71.070 187.880 71.390 188.140 ;
        RECT 73.460 188.080 73.600 188.235 ;
        RECT 86.710 188.220 87.030 188.280 ;
        RECT 89.485 188.235 89.775 188.280 ;
        RECT 92.705 188.235 92.995 188.280 ;
        RECT 96.845 188.235 97.135 188.280 ;
        RECT 75.670 188.080 75.990 188.140 ;
        RECT 73.460 187.940 75.990 188.080 ;
        RECT 75.670 187.880 75.990 187.940 ;
        RECT 76.145 188.080 76.435 188.125 ;
        RECT 77.050 188.080 77.370 188.140 ;
        RECT 76.145 187.940 77.370 188.080 ;
        RECT 76.145 187.895 76.435 187.940 ;
        RECT 77.050 187.880 77.370 187.940 ;
        RECT 77.970 188.080 78.290 188.140 ;
        RECT 82.585 188.080 82.875 188.125 ;
        RECT 77.970 187.940 82.875 188.080 ;
        RECT 77.970 187.880 78.290 187.940 ;
        RECT 82.585 187.895 82.875 187.940 ;
        RECT 83.490 187.880 83.810 188.140 ;
        RECT 84.870 188.080 85.190 188.140 ;
        RECT 87.645 188.080 87.935 188.125 ;
        RECT 84.870 187.940 87.935 188.080 ;
        RECT 84.870 187.880 85.190 187.940 ;
        RECT 87.645 187.895 87.935 187.940 ;
        RECT 91.785 188.080 92.075 188.125 ;
        RECT 93.165 188.080 93.455 188.125 ;
        RECT 91.785 187.940 93.455 188.080 ;
        RECT 91.785 187.895 92.075 187.940 ;
        RECT 93.165 187.895 93.455 187.940 ;
        RECT 98.210 188.080 98.530 188.140 ;
        RECT 103.730 188.080 104.050 188.140 ;
        RECT 98.210 187.940 104.050 188.080 ;
        RECT 106.120 188.080 106.260 188.575 ;
        RECT 106.580 188.420 106.720 188.960 ;
        RECT 107.040 188.805 107.180 189.300 ;
        RECT 111.550 189.240 111.870 189.300 ;
        RECT 120.840 189.300 127.880 189.440 ;
        RECT 118.925 189.100 119.215 189.145 ;
        RECT 109.800 188.960 119.215 189.100 ;
        RECT 106.965 188.575 107.255 188.805 ;
        RECT 107.885 188.760 108.175 188.805 ;
        RECT 108.790 188.760 109.110 188.820 ;
        RECT 109.800 188.805 109.940 188.960 ;
        RECT 118.925 188.915 119.215 188.960 ;
        RECT 107.885 188.620 109.110 188.760 ;
        RECT 107.885 188.575 108.175 188.620 ;
        RECT 108.790 188.560 109.110 188.620 ;
        RECT 109.725 188.575 110.015 188.805 ;
        RECT 110.630 188.560 110.950 188.820 ;
        RECT 111.565 188.760 111.855 188.805 ;
        RECT 112.010 188.760 112.330 188.820 ;
        RECT 111.565 188.620 112.330 188.760 ;
        RECT 111.565 188.575 111.855 188.620 ;
        RECT 112.010 188.560 112.330 188.620 ;
        RECT 116.150 188.760 116.470 188.820 ;
        RECT 116.625 188.760 116.915 188.805 ;
        RECT 120.840 188.760 120.980 189.300 ;
        RECT 126.270 188.900 126.590 189.160 ;
        RECT 116.150 188.620 120.980 188.760 ;
        RECT 116.150 188.560 116.470 188.620 ;
        RECT 116.625 188.575 116.915 188.620 ;
        RECT 122.145 188.575 122.435 188.805 ;
        RECT 107.410 188.420 107.730 188.480 ;
        RECT 106.580 188.280 107.730 188.420 ;
        RECT 107.410 188.220 107.730 188.280 ;
        RECT 111.090 188.220 111.410 188.480 ;
        RECT 113.405 188.080 113.695 188.125 ;
        RECT 106.120 187.940 113.695 188.080 ;
        RECT 122.220 188.080 122.360 188.575 ;
        RECT 124.430 188.560 124.750 188.820 ;
        RECT 125.350 188.560 125.670 188.820 ;
        RECT 125.810 188.560 126.130 188.820 ;
        RECT 127.205 188.575 127.495 188.805 ;
        RECT 127.740 188.760 127.880 189.300 ;
        RECT 128.125 189.300 132.570 189.440 ;
        RECT 128.125 189.255 128.415 189.300 ;
        RECT 132.250 189.240 132.570 189.300 ;
        RECT 148.390 189.440 148.680 189.485 ;
        RECT 150.490 189.440 150.780 189.485 ;
        RECT 152.060 189.440 152.350 189.485 ;
        RECT 148.390 189.300 152.350 189.440 ;
        RECT 148.390 189.255 148.680 189.300 ;
        RECT 150.490 189.255 150.780 189.300 ;
        RECT 152.060 189.255 152.350 189.300 ;
        RECT 129.490 189.100 129.810 189.160 ;
        RECT 133.170 189.100 133.490 189.160 ;
        RECT 148.785 189.100 149.075 189.145 ;
        RECT 149.975 189.100 150.265 189.145 ;
        RECT 152.495 189.100 152.785 189.145 ;
        RECT 129.490 188.960 133.490 189.100 ;
        RECT 129.490 188.900 129.810 188.960 ;
        RECT 133.170 188.900 133.490 188.960 ;
        RECT 139.240 188.960 142.600 189.100 ;
        RECT 129.965 188.760 130.255 188.805 ;
        RECT 130.410 188.760 130.730 188.820 ;
        RECT 127.740 188.620 129.720 188.760 ;
        RECT 124.905 188.420 125.195 188.465 ;
        RECT 127.280 188.420 127.420 188.575 ;
        RECT 129.030 188.420 129.350 188.480 ;
        RECT 124.905 188.280 129.350 188.420 ;
        RECT 129.580 188.420 129.720 188.620 ;
        RECT 129.965 188.620 130.730 188.760 ;
        RECT 129.965 188.575 130.255 188.620 ;
        RECT 130.410 188.560 130.730 188.620 ;
        RECT 130.885 188.760 131.175 188.805 ;
        RECT 134.090 188.760 134.410 188.820 ;
        RECT 130.885 188.620 134.410 188.760 ;
        RECT 130.885 188.575 131.175 188.620 ;
        RECT 130.960 188.420 131.100 188.575 ;
        RECT 134.090 188.560 134.410 188.620 ;
        RECT 136.405 188.575 136.695 188.805 ;
        RECT 138.690 188.760 139.010 188.820 ;
        RECT 139.240 188.805 139.380 188.960 ;
        RECT 142.460 188.805 142.600 188.960 ;
        RECT 148.785 188.960 152.785 189.100 ;
        RECT 148.785 188.915 149.075 188.960 ;
        RECT 149.975 188.915 150.265 188.960 ;
        RECT 152.495 188.915 152.785 188.960 ;
        RECT 139.165 188.760 139.455 188.805 ;
        RECT 138.690 188.620 139.455 188.760 ;
        RECT 129.580 188.280 131.100 188.420 ;
        RECT 136.480 188.420 136.620 188.575 ;
        RECT 138.690 188.560 139.010 188.620 ;
        RECT 139.165 188.575 139.455 188.620 ;
        RECT 141.925 188.575 142.215 188.805 ;
        RECT 142.385 188.575 142.675 188.805 ;
        RECT 143.305 188.760 143.595 188.805 ;
        RECT 143.765 188.760 144.055 188.805 ;
        RECT 145.130 188.760 145.450 188.820 ;
        RECT 143.305 188.620 145.450 188.760 ;
        RECT 143.305 188.575 143.595 188.620 ;
        RECT 143.765 188.575 144.055 188.620 ;
        RECT 140.070 188.420 140.390 188.480 ;
        RECT 142.000 188.420 142.140 188.575 ;
        RECT 145.130 188.560 145.450 188.620 ;
        RECT 146.510 188.760 146.830 188.820 ;
        RECT 147.905 188.760 148.195 188.805 ;
        RECT 150.650 188.760 150.970 188.820 ;
        RECT 146.510 188.620 150.970 188.760 ;
        RECT 146.510 188.560 146.830 188.620 ;
        RECT 147.905 188.575 148.195 188.620 ;
        RECT 150.650 188.560 150.970 188.620 ;
        RECT 149.270 188.465 149.590 188.480 ;
        RECT 136.480 188.280 148.580 188.420 ;
        RECT 124.905 188.235 125.195 188.280 ;
        RECT 129.030 188.220 129.350 188.280 ;
        RECT 140.070 188.220 140.390 188.280 ;
        RECT 123.510 188.080 123.830 188.140 ;
        RECT 129.490 188.080 129.810 188.140 ;
        RECT 122.220 187.940 129.810 188.080 ;
        RECT 98.210 187.880 98.530 187.940 ;
        RECT 103.730 187.880 104.050 187.940 ;
        RECT 113.405 187.895 113.695 187.940 ;
        RECT 123.510 187.880 123.830 187.940 ;
        RECT 129.490 187.880 129.810 187.940 ;
        RECT 130.410 188.080 130.730 188.140 ;
        RECT 135.010 188.080 135.330 188.140 ;
        RECT 130.410 187.940 135.330 188.080 ;
        RECT 130.410 187.880 130.730 187.940 ;
        RECT 135.010 187.880 135.330 187.940 ;
        RECT 145.590 187.880 145.910 188.140 ;
        RECT 146.525 188.080 146.815 188.125 ;
        RECT 147.890 188.080 148.210 188.140 ;
        RECT 146.525 187.940 148.210 188.080 ;
        RECT 148.440 188.080 148.580 188.280 ;
        RECT 149.240 188.235 149.590 188.465 ;
        RECT 149.270 188.220 149.590 188.235 ;
        RECT 154.805 188.080 155.095 188.125 ;
        RECT 148.440 187.940 155.095 188.080 ;
        RECT 146.525 187.895 146.815 187.940 ;
        RECT 147.890 187.880 148.210 187.940 ;
        RECT 154.805 187.895 155.095 187.940 ;
        RECT 22.700 187.260 157.820 187.740 ;
        RECT 25.530 186.860 25.850 187.120 ;
        RECT 31.050 187.060 31.370 187.120 ;
        RECT 31.050 186.920 33.580 187.060 ;
        RECT 31.050 186.860 31.370 186.920 ;
        RECT 33.440 186.765 33.580 186.920 ;
        RECT 33.810 186.860 34.130 187.120 ;
        RECT 47.625 187.060 47.915 187.105 ;
        RECT 48.070 187.060 48.390 187.120 ;
        RECT 47.625 186.920 48.390 187.060 ;
        RECT 47.625 186.875 47.915 186.920 ;
        RECT 48.070 186.860 48.390 186.920 ;
        RECT 50.830 187.060 51.150 187.120 ;
        RECT 60.045 187.060 60.335 187.105 ;
        RECT 60.490 187.060 60.810 187.120 ;
        RECT 67.865 187.060 68.155 187.105 ;
        RECT 50.830 186.920 60.810 187.060 ;
        RECT 50.830 186.860 51.150 186.920 ;
        RECT 60.045 186.875 60.335 186.920 ;
        RECT 60.490 186.860 60.810 186.920 ;
        RECT 61.960 186.920 68.155 187.060 ;
        RECT 61.960 186.765 62.100 186.920 ;
        RECT 67.865 186.875 68.155 186.920 ;
        RECT 77.050 186.860 77.370 187.120 ;
        RECT 85.805 187.060 86.095 187.105 ;
        RECT 91.310 187.060 91.630 187.120 ;
        RECT 102.810 187.060 103.130 187.120 ;
        RECT 85.805 186.920 91.630 187.060 ;
        RECT 85.805 186.875 86.095 186.920 ;
        RECT 91.310 186.860 91.630 186.920 ;
        RECT 98.760 186.920 103.130 187.060 ;
        RECT 32.365 186.720 32.655 186.765 ;
        RECT 33.365 186.720 33.655 186.765 ;
        RECT 34.745 186.720 35.035 186.765 ;
        RECT 32.365 186.580 33.120 186.720 ;
        RECT 32.365 186.535 32.655 186.580 ;
        RECT 26.465 186.380 26.755 186.425 ;
        RECT 31.510 186.380 31.830 186.440 ;
        RECT 26.465 186.240 31.830 186.380 ;
        RECT 32.980 186.380 33.120 186.580 ;
        RECT 33.365 186.580 36.340 186.720 ;
        RECT 33.365 186.535 33.655 186.580 ;
        RECT 34.745 186.535 35.035 186.580 ;
        RECT 35.190 186.380 35.510 186.440 ;
        RECT 32.980 186.240 35.510 186.380 ;
        RECT 26.465 186.195 26.755 186.240 ;
        RECT 31.510 186.180 31.830 186.240 ;
        RECT 35.190 186.180 35.510 186.240 ;
        RECT 35.650 186.180 35.970 186.440 ;
        RECT 36.200 186.425 36.340 186.580 ;
        RECT 61.885 186.535 62.175 186.765 ;
        RECT 62.965 186.720 63.255 186.765 ;
        RECT 69.690 186.720 70.010 186.780 ;
        RECT 72.765 186.720 73.055 186.765 ;
        RECT 62.420 186.580 73.055 186.720 ;
        RECT 36.125 186.195 36.415 186.425 ;
        RECT 36.585 186.380 36.875 186.425 ;
        RECT 41.630 186.380 41.950 186.440 ;
        RECT 36.585 186.240 41.950 186.380 ;
        RECT 36.585 186.195 36.875 186.240 ;
        RECT 41.630 186.180 41.950 186.240 ;
        RECT 46.705 186.380 46.995 186.425 ;
        RECT 47.150 186.380 47.470 186.440 ;
        RECT 46.705 186.240 47.470 186.380 ;
        RECT 46.705 186.195 46.995 186.240 ;
        RECT 47.150 186.180 47.470 186.240 ;
        RECT 48.085 186.380 48.375 186.425 ;
        RECT 48.990 186.380 49.310 186.440 ;
        RECT 48.085 186.240 49.310 186.380 ;
        RECT 48.085 186.195 48.375 186.240 ;
        RECT 48.990 186.180 49.310 186.240 ;
        RECT 49.465 186.195 49.755 186.425 ;
        RECT 37.490 186.040 37.810 186.100 ;
        RECT 39.805 186.040 40.095 186.085 ;
        RECT 37.490 185.900 40.095 186.040 ;
        RECT 47.240 186.040 47.380 186.180 ;
        RECT 49.540 186.040 49.680 186.195 ;
        RECT 50.370 186.180 50.690 186.440 ;
        RECT 50.830 186.180 51.150 186.440 ;
        RECT 52.210 186.380 52.530 186.440 ;
        RECT 53.145 186.380 53.435 186.425 ;
        RECT 54.425 186.380 54.715 186.425 ;
        RECT 52.210 186.240 53.435 186.380 ;
        RECT 52.210 186.180 52.530 186.240 ;
        RECT 53.145 186.195 53.435 186.240 ;
        RECT 53.680 186.240 54.715 186.380 ;
        RECT 53.680 186.040 53.820 186.240 ;
        RECT 54.425 186.195 54.715 186.240 ;
        RECT 61.410 186.380 61.730 186.440 ;
        RECT 62.420 186.380 62.560 186.580 ;
        RECT 62.965 186.535 63.255 186.580 ;
        RECT 69.690 186.520 70.010 186.580 ;
        RECT 72.765 186.535 73.055 186.580 ;
        RECT 73.845 186.720 74.135 186.765 ;
        RECT 78.430 186.720 78.750 186.780 ;
        RECT 73.845 186.580 78.750 186.720 ;
        RECT 73.845 186.535 74.135 186.580 ;
        RECT 78.430 186.520 78.750 186.580 ;
        RECT 78.905 186.720 79.195 186.765 ;
        RECT 83.965 186.720 84.255 186.765 ;
        RECT 78.905 186.580 84.255 186.720 ;
        RECT 78.905 186.535 79.195 186.580 ;
        RECT 83.965 186.535 84.255 186.580 ;
        RECT 65.105 186.380 65.395 186.425 ;
        RECT 61.410 186.240 62.560 186.380 ;
        RECT 63.800 186.240 65.395 186.380 ;
        RECT 61.410 186.180 61.730 186.240 ;
        RECT 47.240 185.900 49.680 186.040 ;
        RECT 53.220 185.900 53.820 186.040 ;
        RECT 54.025 186.040 54.315 186.085 ;
        RECT 55.215 186.040 55.505 186.085 ;
        RECT 57.735 186.040 58.025 186.085 ;
        RECT 54.025 185.900 58.025 186.040 ;
        RECT 37.490 185.840 37.810 185.900 ;
        RECT 39.805 185.855 40.095 185.900 ;
        RECT 31.525 185.700 31.815 185.745 ;
        RECT 31.970 185.700 32.290 185.760 ;
        RECT 36.570 185.700 36.890 185.760 ;
        RECT 40.710 185.700 41.030 185.760 ;
        RECT 41.185 185.700 41.475 185.745 ;
        RECT 31.525 185.560 32.290 185.700 ;
        RECT 31.525 185.515 31.815 185.560 ;
        RECT 31.970 185.500 32.290 185.560 ;
        RECT 33.670 185.560 41.475 185.700 ;
        RECT 32.445 185.360 32.735 185.405 ;
        RECT 33.670 185.360 33.810 185.560 ;
        RECT 36.570 185.500 36.890 185.560 ;
        RECT 40.710 185.500 41.030 185.560 ;
        RECT 41.185 185.515 41.475 185.560 ;
        RECT 51.750 185.500 52.070 185.760 ;
        RECT 32.445 185.220 33.810 185.360 ;
        RECT 42.105 185.360 42.395 185.405 ;
        RECT 43.010 185.360 43.330 185.420 ;
        RECT 42.105 185.220 43.330 185.360 ;
        RECT 32.445 185.175 32.735 185.220 ;
        RECT 42.105 185.175 42.395 185.220 ;
        RECT 43.010 185.160 43.330 185.220 ;
        RECT 44.850 185.360 45.170 185.420 ;
        RECT 45.785 185.360 46.075 185.405 ;
        RECT 44.850 185.220 46.075 185.360 ;
        RECT 53.220 185.360 53.360 185.900 ;
        RECT 54.025 185.855 54.315 185.900 ;
        RECT 55.215 185.855 55.505 185.900 ;
        RECT 57.735 185.855 58.025 185.900 ;
        RECT 63.800 185.745 63.940 186.240 ;
        RECT 65.105 186.195 65.395 186.240 ;
        RECT 66.010 186.180 66.330 186.440 ;
        RECT 66.485 186.380 66.775 186.425 ;
        RECT 67.850 186.380 68.170 186.440 ;
        RECT 66.485 186.240 68.170 186.380 ;
        RECT 66.485 186.195 66.775 186.240 ;
        RECT 67.850 186.180 68.170 186.240 ;
        RECT 70.150 186.380 70.470 186.440 ;
        RECT 70.625 186.380 70.915 186.425 ;
        RECT 70.150 186.240 70.915 186.380 ;
        RECT 70.150 186.180 70.470 186.240 ;
        RECT 70.625 186.195 70.915 186.240 ;
        RECT 71.070 186.380 71.390 186.440 ;
        RECT 76.605 186.380 76.895 186.425 ;
        RECT 71.070 186.240 76.895 186.380 ;
        RECT 71.070 186.180 71.390 186.240 ;
        RECT 76.605 186.195 76.895 186.240 ;
        RECT 77.970 186.180 78.290 186.440 ;
        RECT 80.270 186.180 80.590 186.440 ;
        RECT 81.205 186.195 81.495 186.425 ;
        RECT 81.665 186.380 81.955 186.425 ;
        RECT 82.110 186.380 82.430 186.440 ;
        RECT 81.665 186.240 82.430 186.380 ;
        RECT 81.665 186.195 81.955 186.240 ;
        RECT 77.050 186.040 77.370 186.100 ;
        RECT 81.280 186.040 81.420 186.195 ;
        RECT 82.110 186.180 82.430 186.240 ;
        RECT 83.490 186.180 83.810 186.440 ;
        RECT 84.870 186.180 85.190 186.440 ;
        RECT 93.610 186.380 93.930 186.440 ;
        RECT 88.180 186.240 93.930 186.380 ;
        RECT 88.180 186.040 88.320 186.240 ;
        RECT 93.610 186.180 93.930 186.240 ;
        RECT 98.210 186.180 98.530 186.440 ;
        RECT 98.760 186.425 98.900 186.920 ;
        RECT 102.810 186.860 103.130 186.920 ;
        RECT 103.270 187.060 103.590 187.120 ;
        RECT 128.110 187.060 128.430 187.120 ;
        RECT 132.710 187.060 133.030 187.120 ;
        RECT 103.270 186.920 133.030 187.060 ;
        RECT 103.270 186.860 103.590 186.920 ;
        RECT 128.110 186.860 128.430 186.920 ;
        RECT 132.710 186.860 133.030 186.920 ;
        RECT 138.690 187.060 139.010 187.120 ;
        RECT 139.955 187.060 140.245 187.105 ;
        RECT 138.690 186.920 140.245 187.060 ;
        RECT 138.690 186.860 139.010 186.920 ;
        RECT 139.955 186.875 140.245 186.920 ;
        RECT 148.825 187.060 149.115 187.105 ;
        RECT 149.270 187.060 149.590 187.120 ;
        RECT 148.825 186.920 149.590 187.060 ;
        RECT 148.825 186.875 149.115 186.920 ;
        RECT 149.270 186.860 149.590 186.920 ;
        RECT 99.605 186.720 99.895 186.765 ;
        RECT 118.005 186.720 118.295 186.765 ;
        RECT 99.605 186.580 100.740 186.720 ;
        RECT 99.605 186.535 99.895 186.580 ;
        RECT 100.600 186.425 100.740 186.580 ;
        RECT 110.260 186.580 118.295 186.720 ;
        RECT 98.685 186.195 98.975 186.425 ;
        RECT 100.525 186.195 100.815 186.425 ;
        RECT 101.430 186.180 101.750 186.440 ;
        RECT 103.270 186.180 103.590 186.440 ;
        RECT 106.505 186.380 106.795 186.425 ;
        RECT 108.805 186.380 109.095 186.425 ;
        RECT 109.250 186.380 109.570 186.440 ;
        RECT 110.260 186.425 110.400 186.580 ;
        RECT 118.005 186.535 118.295 186.580 ;
        RECT 122.145 186.720 122.435 186.765 ;
        RECT 125.350 186.720 125.670 186.780 ;
        RECT 126.285 186.720 126.575 186.765 ;
        RECT 141.005 186.720 141.295 186.765 ;
        RECT 144.225 186.720 144.515 186.765 ;
        RECT 122.145 186.580 126.575 186.720 ;
        RECT 122.145 186.535 122.435 186.580 ;
        RECT 125.350 186.520 125.670 186.580 ;
        RECT 126.285 186.535 126.575 186.580 ;
        RECT 126.820 186.580 144.900 186.720 ;
        RECT 106.505 186.240 109.570 186.380 ;
        RECT 106.505 186.195 106.795 186.240 ;
        RECT 108.805 186.195 109.095 186.240 ;
        RECT 109.250 186.180 109.570 186.240 ;
        RECT 110.185 186.195 110.475 186.425 ;
        RECT 111.090 186.180 111.410 186.440 ;
        RECT 111.565 186.195 111.855 186.425 ;
        RECT 77.050 185.900 88.320 186.040 ;
        RECT 99.605 186.040 99.895 186.085 ;
        RECT 104.650 186.040 104.970 186.100 ;
        RECT 105.125 186.040 105.415 186.085 ;
        RECT 108.345 186.040 108.635 186.085 ;
        RECT 99.605 185.900 103.960 186.040 ;
        RECT 77.050 185.840 77.370 185.900 ;
        RECT 99.605 185.855 99.895 185.900 ;
        RECT 53.630 185.700 53.920 185.745 ;
        RECT 55.730 185.700 56.020 185.745 ;
        RECT 57.300 185.700 57.590 185.745 ;
        RECT 53.630 185.560 57.590 185.700 ;
        RECT 53.630 185.515 53.920 185.560 ;
        RECT 55.730 185.515 56.020 185.560 ;
        RECT 57.300 185.515 57.590 185.560 ;
        RECT 63.725 185.515 64.015 185.745 ;
        RECT 71.070 185.700 71.390 185.760 ;
        RECT 72.450 185.700 72.770 185.760 ;
        RECT 71.070 185.560 72.770 185.700 ;
        RECT 71.070 185.500 71.390 185.560 ;
        RECT 72.450 185.500 72.770 185.560 ;
        RECT 100.050 185.700 100.370 185.760 ;
        RECT 103.820 185.745 103.960 185.900 ;
        RECT 104.650 185.900 108.635 186.040 ;
        RECT 104.650 185.840 104.970 185.900 ;
        RECT 105.125 185.855 105.415 185.900 ;
        RECT 108.345 185.855 108.635 185.900 ;
        RECT 109.710 186.040 110.030 186.100 ;
        RECT 111.640 186.040 111.780 186.195 ;
        RECT 112.010 186.180 112.330 186.440 ;
        RECT 123.050 186.180 123.370 186.440 ;
        RECT 123.525 186.195 123.815 186.425 ;
        RECT 109.710 185.900 114.080 186.040 ;
        RECT 109.710 185.840 110.030 185.900 ;
        RECT 101.445 185.700 101.735 185.745 ;
        RECT 100.050 185.560 101.735 185.700 ;
        RECT 100.050 185.500 100.370 185.560 ;
        RECT 101.445 185.515 101.735 185.560 ;
        RECT 103.745 185.515 104.035 185.745 ;
        RECT 105.570 185.700 105.890 185.760 ;
        RECT 106.965 185.700 107.255 185.745 ;
        RECT 105.570 185.560 107.255 185.700 ;
        RECT 105.570 185.500 105.890 185.560 ;
        RECT 106.965 185.515 107.255 185.560 ;
        RECT 111.090 185.700 111.410 185.760 ;
        RECT 113.405 185.700 113.695 185.745 ;
        RECT 111.090 185.560 113.695 185.700 ;
        RECT 113.940 185.700 114.080 185.900 ;
        RECT 116.610 185.840 116.930 186.100 ;
        RECT 121.225 186.040 121.515 186.085 ;
        RECT 121.670 186.040 121.990 186.100 ;
        RECT 121.225 185.900 121.990 186.040 ;
        RECT 121.225 185.855 121.515 185.900 ;
        RECT 121.670 185.840 121.990 185.900 ;
        RECT 123.600 186.040 123.740 186.195 ;
        RECT 124.890 186.180 125.210 186.440 ;
        RECT 126.820 186.040 126.960 186.580 ;
        RECT 141.005 186.535 141.295 186.580 ;
        RECT 144.225 186.535 144.515 186.580 ;
        RECT 127.650 186.180 127.970 186.440 ;
        RECT 129.030 186.180 129.350 186.440 ;
        RECT 135.485 186.380 135.775 186.425 ;
        RECT 138.690 186.380 139.010 186.440 ;
        RECT 135.485 186.240 139.010 186.380 ;
        RECT 135.485 186.195 135.775 186.240 ;
        RECT 138.690 186.180 139.010 186.240 ;
        RECT 123.600 185.900 126.960 186.040 ;
        RECT 118.450 185.700 118.770 185.760 ;
        RECT 113.940 185.560 118.770 185.700 ;
        RECT 111.090 185.500 111.410 185.560 ;
        RECT 113.405 185.515 113.695 185.560 ;
        RECT 118.450 185.500 118.770 185.560 ;
        RECT 54.050 185.360 54.370 185.420 ;
        RECT 53.220 185.220 54.370 185.360 ;
        RECT 44.850 185.160 45.170 185.220 ;
        RECT 45.785 185.175 46.075 185.220 ;
        RECT 54.050 185.160 54.370 185.220 ;
        RECT 62.790 185.160 63.110 185.420 ;
        RECT 63.250 185.360 63.570 185.420 ;
        RECT 64.185 185.360 64.475 185.405 ;
        RECT 63.250 185.220 64.475 185.360 ;
        RECT 63.250 185.160 63.570 185.220 ;
        RECT 64.185 185.175 64.475 185.220 ;
        RECT 68.310 185.360 68.630 185.420 ;
        RECT 72.005 185.360 72.295 185.405 ;
        RECT 68.310 185.220 72.295 185.360 ;
        RECT 68.310 185.160 68.630 185.220 ;
        RECT 72.005 185.175 72.295 185.220 ;
        RECT 72.925 185.360 73.215 185.405 ;
        RECT 74.750 185.360 75.070 185.420 ;
        RECT 72.925 185.220 75.070 185.360 ;
        RECT 72.925 185.175 73.215 185.220 ;
        RECT 74.750 185.160 75.070 185.220 ;
        RECT 79.350 185.160 79.670 185.420 ;
        RECT 101.890 185.360 102.210 185.420 ;
        RECT 104.665 185.360 104.955 185.405 ;
        RECT 101.890 185.220 104.955 185.360 ;
        RECT 101.890 185.160 102.210 185.220 ;
        RECT 104.665 185.175 104.955 185.220 ;
        RECT 112.930 185.160 113.250 185.420 ;
        RECT 120.750 185.360 121.070 185.420 ;
        RECT 123.600 185.360 123.740 185.900 ;
        RECT 127.190 185.840 127.510 186.100 ;
        RECT 131.330 186.040 131.650 186.100 ;
        RECT 127.740 185.900 131.650 186.040 ;
        RECT 144.760 186.040 144.900 186.580 ;
        RECT 145.130 186.520 145.450 186.780 ;
        RECT 147.890 186.180 148.210 186.440 ;
        RECT 145.130 186.040 145.450 186.100 ;
        RECT 144.760 185.900 145.450 186.040 ;
        RECT 126.745 185.700 127.035 185.745 ;
        RECT 127.740 185.700 127.880 185.900 ;
        RECT 131.330 185.840 131.650 185.900 ;
        RECT 145.130 185.840 145.450 185.900 ;
        RECT 126.745 185.560 127.880 185.700 ;
        RECT 128.125 185.700 128.415 185.745 ;
        RECT 130.870 185.700 131.190 185.760 ;
        RECT 128.125 185.560 131.190 185.700 ;
        RECT 126.745 185.515 127.035 185.560 ;
        RECT 128.125 185.515 128.415 185.560 ;
        RECT 130.870 185.500 131.190 185.560 ;
        RECT 139.165 185.700 139.455 185.745 ;
        RECT 141.450 185.700 141.770 185.760 ;
        RECT 139.165 185.560 141.770 185.700 ;
        RECT 139.165 185.515 139.455 185.560 ;
        RECT 141.450 185.500 141.770 185.560 ;
        RECT 120.750 185.220 123.740 185.360 ;
        RECT 120.750 185.160 121.070 185.220 ;
        RECT 124.430 185.160 124.750 185.420 ;
        RECT 136.405 185.360 136.695 185.405 ;
        RECT 136.850 185.360 137.170 185.420 ;
        RECT 136.405 185.220 137.170 185.360 ;
        RECT 136.405 185.175 136.695 185.220 ;
        RECT 136.850 185.160 137.170 185.220 ;
        RECT 140.070 185.160 140.390 185.420 ;
        RECT 143.290 185.160 143.610 185.420 ;
        RECT 22.700 184.540 157.020 185.020 ;
        RECT 54.970 184.140 55.290 184.400 ;
        RECT 60.045 184.340 60.335 184.385 ;
        RECT 62.790 184.340 63.110 184.400 ;
        RECT 68.770 184.340 69.090 184.400 ;
        RECT 69.705 184.340 69.995 184.385 ;
        RECT 60.045 184.200 68.540 184.340 ;
        RECT 60.045 184.155 60.335 184.200 ;
        RECT 62.790 184.140 63.110 184.200 ;
        RECT 33.810 184.000 34.130 184.060 ;
        RECT 31.600 183.860 34.130 184.000 ;
        RECT 31.600 183.365 31.740 183.860 ;
        RECT 33.810 183.800 34.130 183.860 ;
        RECT 62.370 184.000 62.660 184.045 ;
        RECT 64.470 184.000 64.760 184.045 ;
        RECT 66.040 184.000 66.330 184.045 ;
        RECT 62.370 183.860 66.330 184.000 ;
        RECT 68.400 184.000 68.540 184.200 ;
        RECT 68.770 184.200 69.995 184.340 ;
        RECT 68.770 184.140 69.090 184.200 ;
        RECT 69.705 184.155 69.995 184.200 ;
        RECT 71.070 184.340 71.390 184.400 ;
        RECT 72.005 184.340 72.295 184.385 ;
        RECT 71.070 184.200 72.295 184.340 ;
        RECT 71.070 184.140 71.390 184.200 ;
        RECT 72.005 184.155 72.295 184.200 ;
        RECT 78.430 184.340 78.750 184.400 ;
        RECT 79.365 184.340 79.655 184.385 ;
        RECT 94.070 184.340 94.390 184.400 ;
        RECT 94.545 184.340 94.835 184.385 ;
        RECT 78.430 184.200 79.655 184.340 ;
        RECT 78.430 184.140 78.750 184.200 ;
        RECT 79.365 184.155 79.655 184.200 ;
        RECT 81.970 184.200 93.840 184.340 ;
        RECT 74.750 184.000 75.070 184.060 ;
        RECT 68.400 183.860 75.070 184.000 ;
        RECT 62.370 183.815 62.660 183.860 ;
        RECT 64.470 183.815 64.760 183.860 ;
        RECT 66.040 183.815 66.330 183.860 ;
        RECT 74.750 183.800 75.070 183.860 ;
        RECT 75.210 184.000 75.530 184.060 ;
        RECT 81.970 184.000 82.110 184.200 ;
        RECT 75.210 183.860 82.110 184.000 ;
        RECT 88.130 184.000 88.420 184.045 ;
        RECT 90.230 184.000 90.520 184.045 ;
        RECT 91.800 184.000 92.090 184.045 ;
        RECT 88.130 183.860 92.090 184.000 ;
        RECT 93.700 184.000 93.840 184.200 ;
        RECT 94.070 184.200 94.835 184.340 ;
        RECT 94.070 184.140 94.390 184.200 ;
        RECT 94.545 184.155 94.835 184.200 ;
        RECT 99.130 184.340 99.450 184.400 ;
        RECT 101.890 184.340 102.210 184.400 ;
        RECT 99.130 184.200 102.210 184.340 ;
        RECT 99.130 184.140 99.450 184.200 ;
        RECT 101.890 184.140 102.210 184.200 ;
        RECT 122.145 184.340 122.435 184.385 ;
        RECT 123.970 184.340 124.290 184.400 ;
        RECT 122.145 184.200 124.290 184.340 ;
        RECT 122.145 184.155 122.435 184.200 ;
        RECT 123.970 184.140 124.290 184.200 ;
        RECT 124.890 184.340 125.210 184.400 ;
        RECT 129.950 184.340 130.270 184.400 ;
        RECT 131.345 184.340 131.635 184.385 ;
        RECT 124.890 184.200 131.635 184.340 ;
        RECT 124.890 184.140 125.210 184.200 ;
        RECT 129.950 184.140 130.270 184.200 ;
        RECT 131.345 184.155 131.635 184.200 ;
        RECT 138.690 184.340 139.010 184.400 ;
        RECT 139.165 184.340 139.455 184.385 ;
        RECT 138.690 184.200 139.455 184.340 ;
        RECT 138.690 184.140 139.010 184.200 ;
        RECT 139.165 184.155 139.455 184.200 ;
        RECT 140.070 184.140 140.390 184.400 ;
        RECT 143.290 184.140 143.610 184.400 ;
        RECT 144.685 184.340 144.975 184.385 ;
        RECT 145.130 184.340 145.450 184.400 ;
        RECT 144.685 184.200 145.450 184.340 ;
        RECT 144.685 184.155 144.975 184.200 ;
        RECT 145.130 184.140 145.450 184.200 ;
        RECT 103.270 184.000 103.590 184.060 ;
        RECT 93.700 183.860 103.590 184.000 ;
        RECT 75.210 183.800 75.530 183.860 ;
        RECT 88.130 183.815 88.420 183.860 ;
        RECT 90.230 183.815 90.520 183.860 ;
        RECT 91.800 183.815 92.090 183.860 ;
        RECT 103.270 183.800 103.590 183.860 ;
        RECT 113.890 184.000 114.180 184.045 ;
        RECT 115.990 184.000 116.280 184.045 ;
        RECT 117.560 184.000 117.850 184.045 ;
        RECT 113.890 183.860 117.850 184.000 ;
        RECT 113.890 183.815 114.180 183.860 ;
        RECT 115.990 183.815 116.280 183.860 ;
        RECT 117.560 183.815 117.850 183.860 ;
        RECT 123.525 184.000 123.815 184.045 ;
        RECT 127.190 184.000 127.510 184.060 ;
        RECT 123.525 183.860 127.510 184.000 ;
        RECT 123.525 183.815 123.815 183.860 ;
        RECT 31.970 183.660 32.290 183.720 ;
        RECT 31.970 183.520 33.120 183.660 ;
        RECT 31.970 183.460 32.290 183.520 ;
        RECT 32.980 183.365 33.120 183.520 ;
        RECT 33.350 183.460 33.670 183.720 ;
        RECT 44.850 183.460 45.170 183.720 ;
        RECT 54.510 183.660 54.830 183.720 ;
        RECT 62.765 183.660 63.055 183.705 ;
        RECT 63.955 183.660 64.245 183.705 ;
        RECT 66.475 183.660 66.765 183.705 ;
        RECT 54.510 183.520 57.040 183.660 ;
        RECT 54.510 183.460 54.830 183.520 ;
        RECT 31.525 183.135 31.815 183.365 ;
        RECT 32.445 183.135 32.735 183.365 ;
        RECT 32.905 183.135 33.195 183.365 ;
        RECT 33.440 183.320 33.580 183.460 ;
        RECT 33.825 183.320 34.115 183.365 ;
        RECT 33.440 183.180 34.115 183.320 ;
        RECT 33.825 183.135 34.115 183.180 ;
        RECT 32.520 182.980 32.660 183.135 ;
        RECT 34.270 183.120 34.590 183.380 ;
        RECT 42.090 183.320 42.410 183.380 ;
        RECT 44.405 183.320 44.695 183.365 ;
        RECT 42.090 183.180 44.695 183.320 ;
        RECT 42.090 183.120 42.410 183.180 ;
        RECT 44.405 183.135 44.695 183.180 ;
        RECT 45.310 183.120 45.630 183.380 ;
        RECT 45.770 183.120 46.090 183.380 ;
        RECT 51.290 183.320 51.610 183.380 ;
        RECT 54.970 183.320 55.290 183.380 ;
        RECT 56.900 183.365 57.040 183.520 ;
        RECT 62.765 183.520 66.765 183.660 ;
        RECT 62.765 183.475 63.055 183.520 ;
        RECT 63.955 183.475 64.245 183.520 ;
        RECT 66.475 183.475 66.765 183.520 ;
        RECT 66.930 183.660 67.250 183.720 ;
        RECT 74.290 183.660 74.610 183.720 ;
        RECT 66.930 183.520 71.300 183.660 ;
        RECT 66.930 183.460 67.250 183.520 ;
        RECT 55.905 183.320 56.195 183.365 ;
        RECT 51.290 183.180 56.195 183.320 ;
        RECT 51.290 183.120 51.610 183.180 ;
        RECT 54.970 183.120 55.290 183.180 ;
        RECT 55.905 183.135 56.195 183.180 ;
        RECT 56.825 183.135 57.115 183.365 ;
        RECT 57.270 183.320 57.590 183.380 ;
        RECT 57.745 183.320 58.035 183.365 ;
        RECT 61.410 183.320 61.730 183.380 ;
        RECT 57.270 183.180 58.035 183.320 ;
        RECT 57.270 183.120 57.590 183.180 ;
        RECT 57.745 183.135 58.035 183.180 ;
        RECT 60.120 183.180 61.730 183.320 ;
        RECT 33.365 182.980 33.655 183.025 ;
        RECT 32.520 182.840 33.655 182.980 ;
        RECT 32.980 182.700 33.120 182.840 ;
        RECT 33.365 182.795 33.655 182.840 ;
        RECT 36.110 182.780 36.430 183.040 ;
        RECT 37.950 182.980 38.270 183.040 ;
        RECT 39.805 182.980 40.095 183.025 ;
        RECT 37.950 182.840 40.095 182.980 ;
        RECT 37.950 182.780 38.270 182.840 ;
        RECT 39.805 182.795 40.095 182.840 ;
        RECT 56.365 182.795 56.655 183.025 ;
        RECT 29.210 182.640 29.530 182.700 ;
        RECT 31.525 182.640 31.815 182.685 ;
        RECT 29.210 182.500 31.815 182.640 ;
        RECT 29.210 182.440 29.530 182.500 ;
        RECT 31.525 182.455 31.815 182.500 ;
        RECT 32.890 182.440 33.210 182.700 ;
        RECT 35.190 182.440 35.510 182.700 ;
        RECT 41.170 182.640 41.490 182.700 ;
        RECT 43.485 182.640 43.775 182.685 ;
        RECT 41.170 182.500 43.775 182.640 ;
        RECT 56.440 182.640 56.580 182.795 ;
        RECT 59.110 182.780 59.430 183.040 ;
        RECT 60.120 183.025 60.260 183.180 ;
        RECT 61.410 183.120 61.730 183.180 ;
        RECT 61.870 183.120 62.190 183.380 ;
        RECT 63.250 183.365 63.570 183.380 ;
        RECT 63.220 183.320 63.570 183.365 ;
        RECT 63.055 183.180 63.570 183.320 ;
        RECT 63.220 183.135 63.570 183.180 ;
        RECT 63.250 183.120 63.570 183.135 ;
        RECT 70.610 183.120 70.930 183.380 ;
        RECT 71.160 183.365 71.300 183.520 ;
        RECT 72.540 183.520 74.610 183.660 ;
        RECT 72.540 183.365 72.680 183.520 ;
        RECT 74.290 183.460 74.610 183.520 ;
        RECT 75.670 183.660 75.990 183.720 ;
        RECT 78.445 183.660 78.735 183.705 ;
        RECT 83.030 183.660 83.350 183.720 ;
        RECT 87.645 183.660 87.935 183.705 ;
        RECT 75.670 183.520 87.935 183.660 ;
        RECT 75.670 183.460 75.990 183.520 ;
        RECT 78.445 183.475 78.735 183.520 ;
        RECT 83.030 183.460 83.350 183.520 ;
        RECT 87.645 183.475 87.935 183.520 ;
        RECT 88.525 183.660 88.815 183.705 ;
        RECT 89.715 183.660 90.005 183.705 ;
        RECT 92.235 183.660 92.525 183.705 ;
        RECT 88.525 183.520 92.525 183.660 ;
        RECT 88.525 183.475 88.815 183.520 ;
        RECT 89.715 183.475 90.005 183.520 ;
        RECT 92.235 183.475 92.525 183.520 ;
        RECT 94.070 183.660 94.390 183.720 ;
        RECT 96.845 183.660 97.135 183.705 ;
        RECT 94.070 183.520 97.135 183.660 ;
        RECT 94.070 183.460 94.390 183.520 ;
        RECT 96.845 183.475 97.135 183.520 ;
        RECT 98.670 183.660 98.990 183.720 ;
        RECT 99.145 183.660 99.435 183.705 ;
        RECT 98.670 183.520 99.435 183.660 ;
        RECT 98.670 183.460 98.990 183.520 ;
        RECT 99.145 183.475 99.435 183.520 ;
        RECT 103.730 183.460 104.050 183.720 ;
        RECT 112.010 183.660 112.330 183.720 ;
        RECT 109.340 183.520 112.330 183.660 ;
        RECT 109.340 183.380 109.480 183.520 ;
        RECT 112.010 183.460 112.330 183.520 ;
        RECT 113.390 183.460 113.710 183.720 ;
        RECT 114.285 183.660 114.575 183.705 ;
        RECT 115.475 183.660 115.765 183.705 ;
        RECT 117.995 183.660 118.285 183.705 ;
        RECT 114.285 183.520 118.285 183.660 ;
        RECT 114.285 183.475 114.575 183.520 ;
        RECT 115.475 183.475 115.765 183.520 ;
        RECT 117.995 183.475 118.285 183.520 ;
        RECT 71.085 183.135 71.375 183.365 ;
        RECT 72.465 183.135 72.755 183.365 ;
        RECT 76.130 183.320 76.450 183.380 ;
        RECT 82.125 183.320 82.415 183.365 ;
        RECT 76.130 183.180 82.415 183.320 ;
        RECT 76.130 183.120 76.450 183.180 ;
        RECT 82.125 183.135 82.415 183.180 ;
        RECT 83.950 183.120 84.270 183.380 ;
        RECT 95.925 183.320 96.215 183.365 ;
        RECT 97.290 183.320 97.610 183.380 ;
        RECT 95.925 183.180 97.610 183.320 ;
        RECT 95.925 183.135 96.215 183.180 ;
        RECT 97.290 183.120 97.610 183.180 ;
        RECT 98.225 183.320 98.515 183.365 ;
        RECT 100.050 183.320 100.370 183.380 ;
        RECT 98.225 183.180 100.370 183.320 ;
        RECT 98.225 183.135 98.515 183.180 ;
        RECT 100.050 183.120 100.370 183.180 ;
        RECT 102.810 183.120 103.130 183.380 ;
        RECT 109.250 183.120 109.570 183.380 ;
        RECT 110.185 183.320 110.475 183.365 ;
        RECT 110.630 183.320 110.950 183.380 ;
        RECT 110.185 183.180 110.950 183.320 ;
        RECT 110.185 183.135 110.475 183.180 ;
        RECT 110.630 183.120 110.950 183.180 ;
        RECT 111.090 183.120 111.410 183.380 ;
        RECT 112.930 183.320 113.250 183.380 ;
        RECT 114.685 183.320 114.975 183.365 ;
        RECT 112.930 183.180 114.975 183.320 ;
        RECT 112.930 183.120 113.250 183.180 ;
        RECT 114.685 183.135 114.975 183.180 ;
        RECT 120.765 183.320 121.055 183.365 ;
        RECT 121.210 183.320 121.530 183.380 ;
        RECT 123.050 183.320 123.370 183.380 ;
        RECT 120.765 183.180 123.370 183.320 ;
        RECT 120.765 183.135 121.055 183.180 ;
        RECT 121.210 183.120 121.530 183.180 ;
        RECT 123.050 183.120 123.370 183.180 ;
        RECT 60.120 182.840 60.415 183.025 ;
        RECT 66.010 182.980 66.330 183.040 ;
        RECT 60.125 182.795 60.415 182.840 ;
        RECT 60.580 182.840 66.330 182.980 ;
        RECT 59.570 182.640 59.890 182.700 ;
        RECT 60.580 182.640 60.720 182.840 ;
        RECT 66.010 182.780 66.330 182.840 ;
        RECT 69.230 182.980 69.550 183.040 ;
        RECT 71.530 182.980 71.850 183.040 ;
        RECT 74.305 182.980 74.595 183.025 ;
        RECT 69.230 182.840 74.595 182.980 ;
        RECT 69.230 182.780 69.550 182.840 ;
        RECT 71.530 182.780 71.850 182.840 ;
        RECT 74.305 182.795 74.595 182.840 ;
        RECT 88.090 182.980 88.410 183.040 ;
        RECT 88.870 182.980 89.160 183.025 ;
        RECT 88.090 182.840 89.160 182.980 ;
        RECT 88.090 182.780 88.410 182.840 ;
        RECT 88.870 182.795 89.160 182.840 ;
        RECT 109.710 182.780 110.030 183.040 ;
        RECT 121.670 182.980 121.990 183.040 ;
        RECT 120.380 182.840 121.990 182.980 ;
        RECT 56.440 182.500 60.720 182.640 ;
        RECT 60.965 182.640 61.255 182.685 ;
        RECT 66.930 182.640 67.250 182.700 ;
        RECT 60.965 182.500 67.250 182.640 ;
        RECT 41.170 182.440 41.490 182.500 ;
        RECT 43.485 182.455 43.775 182.500 ;
        RECT 59.570 182.440 59.890 182.500 ;
        RECT 60.965 182.455 61.255 182.500 ;
        RECT 66.930 182.440 67.250 182.500 ;
        RECT 68.785 182.640 69.075 182.685 ;
        RECT 70.150 182.640 70.470 182.700 ;
        RECT 68.785 182.500 70.470 182.640 ;
        RECT 68.785 182.455 69.075 182.500 ;
        RECT 70.150 182.440 70.470 182.500 ;
        RECT 84.870 182.640 85.190 182.700 ;
        RECT 86.725 182.640 87.015 182.685 ;
        RECT 84.870 182.500 87.015 182.640 ;
        RECT 84.870 182.440 85.190 182.500 ;
        RECT 86.725 182.455 87.015 182.500 ;
        RECT 94.990 182.440 95.310 182.700 ;
        RECT 108.330 182.440 108.650 182.700 ;
        RECT 120.380 182.685 120.520 182.840 ;
        RECT 121.670 182.780 121.990 182.840 ;
        RECT 122.145 182.980 122.435 183.025 ;
        RECT 123.600 182.980 123.740 183.815 ;
        RECT 127.190 183.800 127.510 183.860 ;
        RECT 134.090 184.000 134.380 184.045 ;
        RECT 135.660 184.000 135.950 184.045 ;
        RECT 137.760 184.000 138.050 184.045 ;
        RECT 134.090 183.860 138.050 184.000 ;
        RECT 134.090 183.815 134.380 183.860 ;
        RECT 135.660 183.815 135.950 183.860 ;
        RECT 137.760 183.815 138.050 183.860 ;
        RECT 141.450 183.800 141.770 184.060 ;
        RECT 147.430 184.000 147.720 184.045 ;
        RECT 149.000 184.000 149.290 184.045 ;
        RECT 151.100 184.000 151.390 184.045 ;
        RECT 147.430 183.860 151.390 184.000 ;
        RECT 147.430 183.815 147.720 183.860 ;
        RECT 149.000 183.815 149.290 183.860 ;
        RECT 151.100 183.815 151.390 183.860 ;
        RECT 126.285 183.660 126.575 183.705 ;
        RECT 124.520 183.520 126.575 183.660 ;
        RECT 124.520 183.380 124.660 183.520 ;
        RECT 126.285 183.475 126.575 183.520 ;
        RECT 133.655 183.660 133.945 183.705 ;
        RECT 136.175 183.660 136.465 183.705 ;
        RECT 137.365 183.660 137.655 183.705 ;
        RECT 133.655 183.520 137.655 183.660 ;
        RECT 133.655 183.475 133.945 183.520 ;
        RECT 136.175 183.475 136.465 183.520 ;
        RECT 137.365 183.475 137.655 183.520 ;
        RECT 138.245 183.660 138.535 183.705 ;
        RECT 146.510 183.660 146.830 183.720 ;
        RECT 138.245 183.520 146.830 183.660 ;
        RECT 138.245 183.475 138.535 183.520 ;
        RECT 146.510 183.460 146.830 183.520 ;
        RECT 146.995 183.660 147.285 183.705 ;
        RECT 149.515 183.660 149.805 183.705 ;
        RECT 150.705 183.660 150.995 183.705 ;
        RECT 146.995 183.520 150.995 183.660 ;
        RECT 146.995 183.475 147.285 183.520 ;
        RECT 149.515 183.475 149.805 183.520 ;
        RECT 150.705 183.475 150.995 183.520 ;
        RECT 124.430 183.120 124.750 183.380 ;
        RECT 124.890 183.120 125.210 183.380 ;
        RECT 136.850 183.365 137.170 183.380 ;
        RECT 125.825 183.135 126.115 183.365 ;
        RECT 136.850 183.320 137.200 183.365 ;
        RECT 145.590 183.320 145.910 183.380 ;
        RECT 136.850 183.180 137.365 183.320 ;
        RECT 141.080 183.180 145.910 183.320 ;
        RECT 146.600 183.320 146.740 183.460 ;
        RECT 151.585 183.320 151.875 183.365 ;
        RECT 146.600 183.180 151.875 183.320 ;
        RECT 136.850 183.135 137.200 183.180 ;
        RECT 122.145 182.840 123.740 182.980 ;
        RECT 122.145 182.795 122.435 182.840 ;
        RECT 120.305 182.455 120.595 182.685 ;
        RECT 120.750 182.640 121.070 182.700 ;
        RECT 121.225 182.640 121.515 182.685 ;
        RECT 120.750 182.500 121.515 182.640 ;
        RECT 121.760 182.640 121.900 182.780 ;
        RECT 125.900 182.640 126.040 183.135 ;
        RECT 136.850 183.120 137.170 183.135 ;
        RECT 141.080 183.025 141.220 183.180 ;
        RECT 145.590 183.120 145.910 183.180 ;
        RECT 151.585 183.135 151.875 183.180 ;
        RECT 141.005 182.795 141.295 183.025 ;
        RECT 145.130 182.980 145.450 183.040 ;
        RECT 144.300 182.840 145.450 182.980 ;
        RECT 121.760 182.500 126.040 182.640 ;
        RECT 136.850 182.640 137.170 182.700 ;
        RECT 139.955 182.640 140.245 182.685 ;
        RECT 136.850 182.500 140.245 182.640 ;
        RECT 120.750 182.440 121.070 182.500 ;
        RECT 121.225 182.455 121.515 182.500 ;
        RECT 136.850 182.440 137.170 182.500 ;
        RECT 139.955 182.455 140.245 182.500 ;
        RECT 143.290 182.440 143.610 182.700 ;
        RECT 144.300 182.685 144.440 182.840 ;
        RECT 145.130 182.780 145.450 182.840 ;
        RECT 146.050 182.980 146.370 183.040 ;
        RECT 150.250 182.980 150.540 183.025 ;
        RECT 146.050 182.840 150.540 182.980 ;
        RECT 146.050 182.780 146.370 182.840 ;
        RECT 150.250 182.795 150.540 182.840 ;
        RECT 144.225 182.455 144.515 182.685 ;
        RECT 22.700 181.820 157.820 182.300 ;
        RECT 33.350 181.620 33.670 181.680 ;
        RECT 40.725 181.620 41.015 181.665 ;
        RECT 32.980 181.480 41.015 181.620 ;
        RECT 25.160 181.140 26.220 181.280 ;
        RECT 24.150 180.940 24.470 181.000 ;
        RECT 25.160 180.940 25.300 181.140 ;
        RECT 25.530 180.985 25.850 181.000 ;
        RECT 24.150 180.800 25.300 180.940 ;
        RECT 24.150 180.740 24.470 180.800 ;
        RECT 25.500 180.755 25.850 180.985 ;
        RECT 26.080 180.940 26.220 181.140 ;
        RECT 31.525 180.940 31.815 180.985 ;
        RECT 31.970 180.940 32.290 181.000 ;
        RECT 26.080 180.800 30.360 180.940 ;
        RECT 25.530 180.740 25.850 180.755 ;
        RECT 25.045 180.600 25.335 180.645 ;
        RECT 26.235 180.600 26.525 180.645 ;
        RECT 28.755 180.600 29.045 180.645 ;
        RECT 25.045 180.460 29.045 180.600 ;
        RECT 25.045 180.415 25.335 180.460 ;
        RECT 26.235 180.415 26.525 180.460 ;
        RECT 28.755 180.415 29.045 180.460 ;
        RECT 24.650 180.260 24.940 180.305 ;
        RECT 26.750 180.260 27.040 180.305 ;
        RECT 28.320 180.260 28.610 180.305 ;
        RECT 24.650 180.120 28.610 180.260 ;
        RECT 30.220 180.260 30.360 180.800 ;
        RECT 31.525 180.800 32.290 180.940 ;
        RECT 31.525 180.755 31.815 180.800 ;
        RECT 31.970 180.740 32.290 180.800 ;
        RECT 32.445 180.940 32.735 180.985 ;
        RECT 32.980 180.940 33.120 181.480 ;
        RECT 33.350 181.420 33.670 181.480 ;
        RECT 40.725 181.435 41.015 181.480 ;
        RECT 42.090 181.420 42.410 181.680 ;
        RECT 47.610 181.620 47.930 181.680 ;
        RECT 48.085 181.620 48.375 181.665 ;
        RECT 47.610 181.480 48.375 181.620 ;
        RECT 47.610 181.420 47.930 181.480 ;
        RECT 48.085 181.435 48.375 181.480 ;
        RECT 59.110 181.620 59.430 181.680 ;
        RECT 69.705 181.620 69.995 181.665 ;
        RECT 59.110 181.480 69.995 181.620 ;
        RECT 59.110 181.420 59.430 181.480 ;
        RECT 69.705 181.435 69.995 181.480 ;
        RECT 70.150 181.620 70.470 181.680 ;
        RECT 80.270 181.620 80.590 181.680 ;
        RECT 83.045 181.620 83.335 181.665 ;
        RECT 70.150 181.480 80.040 181.620 ;
        RECT 70.150 181.420 70.470 181.480 ;
        RECT 37.950 181.280 38.270 181.340 ;
        RECT 33.900 181.140 38.270 181.280 ;
        RECT 33.900 180.985 34.040 181.140 ;
        RECT 37.950 181.080 38.270 181.140 ;
        RECT 54.510 181.280 54.830 181.340 ;
        RECT 59.585 181.280 59.875 181.325 ;
        RECT 54.510 181.140 59.875 181.280 ;
        RECT 54.510 181.080 54.830 181.140 ;
        RECT 59.585 181.095 59.875 181.140 ;
        RECT 61.410 181.280 61.730 181.340 ;
        RECT 67.405 181.280 67.695 181.325 ;
        RECT 75.210 181.280 75.530 181.340 ;
        RECT 61.410 181.140 75.530 181.280 ;
        RECT 61.410 181.080 61.730 181.140 ;
        RECT 67.405 181.095 67.695 181.140 ;
        RECT 75.210 181.080 75.530 181.140 ;
        RECT 77.020 181.280 77.310 181.325 ;
        RECT 79.350 181.280 79.670 181.340 ;
        RECT 77.020 181.140 79.670 181.280 ;
        RECT 79.900 181.280 80.040 181.480 ;
        RECT 80.270 181.480 83.335 181.620 ;
        RECT 80.270 181.420 80.590 181.480 ;
        RECT 83.045 181.435 83.335 181.480 ;
        RECT 88.090 181.620 88.410 181.680 ;
        RECT 89.485 181.620 89.775 181.665 ;
        RECT 88.090 181.480 89.775 181.620 ;
        RECT 88.090 181.420 88.410 181.480 ;
        RECT 89.485 181.435 89.775 181.480 ;
        RECT 91.785 181.435 92.075 181.665 ;
        RECT 94.085 181.620 94.375 181.665 ;
        RECT 94.990 181.620 95.310 181.680 ;
        RECT 94.085 181.480 95.310 181.620 ;
        RECT 94.085 181.435 94.375 181.480 ;
        RECT 83.805 181.280 84.095 181.325 ;
        RECT 79.900 181.140 84.640 181.280 ;
        RECT 77.020 181.095 77.310 181.140 ;
        RECT 79.350 181.080 79.670 181.140 ;
        RECT 83.805 181.095 84.095 181.140 ;
        RECT 35.190 180.985 35.510 181.000 ;
        RECT 32.445 180.800 33.120 180.940 ;
        RECT 32.445 180.755 32.735 180.800 ;
        RECT 33.825 180.755 34.115 180.985 ;
        RECT 35.160 180.940 35.510 180.985 ;
        RECT 34.995 180.800 35.510 180.940 ;
        RECT 35.160 180.755 35.510 180.800 ;
        RECT 30.590 180.600 30.910 180.660 ;
        RECT 32.520 180.600 32.660 180.755 ;
        RECT 30.590 180.460 32.660 180.600 ;
        RECT 30.590 180.400 30.910 180.460 ;
        RECT 33.900 180.260 34.040 180.755 ;
        RECT 35.190 180.740 35.510 180.755 ;
        RECT 44.850 180.740 45.170 181.000 ;
        RECT 45.310 180.740 45.630 181.000 ;
        RECT 54.970 180.740 55.290 181.000 ;
        RECT 56.365 180.940 56.655 180.985 ;
        RECT 58.190 180.940 58.510 181.000 ;
        RECT 56.365 180.800 58.510 180.940 ;
        RECT 56.365 180.755 56.655 180.800 ;
        RECT 58.190 180.740 58.510 180.800 ;
        RECT 58.665 180.755 58.955 180.985 ;
        RECT 59.125 180.755 59.415 180.985 ;
        RECT 60.505 180.940 60.795 180.985 ;
        RECT 62.345 180.940 62.635 180.985 ;
        RECT 60.505 180.800 62.635 180.940 ;
        RECT 60.505 180.755 60.795 180.800 ;
        RECT 62.345 180.755 62.635 180.800 ;
        RECT 66.945 180.940 67.235 180.985 ;
        RECT 67.850 180.940 68.170 181.000 ;
        RECT 66.945 180.800 68.170 180.940 ;
        RECT 66.945 180.755 67.235 180.800 ;
        RECT 34.705 180.600 34.995 180.645 ;
        RECT 35.895 180.600 36.185 180.645 ;
        RECT 38.415 180.600 38.705 180.645 ;
        RECT 34.705 180.460 38.705 180.600 ;
        RECT 34.705 180.415 34.995 180.460 ;
        RECT 35.895 180.415 36.185 180.460 ;
        RECT 38.415 180.415 38.705 180.460 ;
        RECT 43.485 180.600 43.775 180.645 ;
        RECT 44.390 180.600 44.710 180.660 ;
        RECT 43.485 180.460 44.710 180.600 ;
        RECT 43.485 180.415 43.775 180.460 ;
        RECT 44.390 180.400 44.710 180.460 ;
        RECT 46.690 180.400 47.010 180.660 ;
        RECT 54.510 180.400 54.830 180.660 ;
        RECT 55.060 180.600 55.200 180.740 ;
        RECT 58.740 180.600 58.880 180.755 ;
        RECT 55.060 180.460 58.880 180.600 ;
        RECT 59.200 180.600 59.340 180.755 ;
        RECT 67.850 180.740 68.170 180.800 ;
        RECT 68.310 180.740 68.630 181.000 ;
        RECT 70.610 180.940 70.930 181.000 ;
        RECT 72.465 180.940 72.755 180.985 ;
        RECT 70.610 180.800 72.755 180.940 ;
        RECT 70.610 180.740 70.930 180.800 ;
        RECT 72.465 180.755 72.755 180.800 ;
        RECT 75.670 180.740 75.990 181.000 ;
        RECT 84.500 180.940 84.640 181.140 ;
        RECT 84.870 181.080 85.190 181.340 ;
        RECT 89.930 180.940 90.250 181.000 ;
        RECT 84.500 180.800 90.250 180.940 ;
        RECT 89.930 180.740 90.250 180.800 ;
        RECT 90.405 180.940 90.695 180.985 ;
        RECT 91.860 180.940 92.000 181.435 ;
        RECT 94.990 181.420 95.310 181.480 ;
        RECT 115.705 181.620 115.995 181.665 ;
        RECT 116.610 181.620 116.930 181.680 ;
        RECT 115.705 181.480 116.930 181.620 ;
        RECT 115.705 181.435 115.995 181.480 ;
        RECT 116.610 181.420 116.930 181.480 ;
        RECT 121.210 181.420 121.530 181.680 ;
        RECT 126.730 181.620 127.050 181.680 ;
        RECT 130.410 181.620 130.730 181.680 ;
        RECT 133.630 181.620 133.950 181.680 ;
        RECT 126.730 181.480 133.950 181.620 ;
        RECT 126.730 181.420 127.050 181.480 ;
        RECT 130.410 181.420 130.730 181.480 ;
        RECT 133.630 181.420 133.950 181.480 ;
        RECT 136.850 181.420 137.170 181.680 ;
        RECT 141.450 181.620 141.770 181.680 ;
        RECT 138.780 181.480 141.770 181.620 ;
        RECT 108.330 181.280 108.650 181.340 ;
        RECT 110.030 181.280 110.320 181.325 ;
        RECT 108.330 181.140 110.320 181.280 ;
        RECT 108.330 181.080 108.650 181.140 ;
        RECT 110.030 181.095 110.320 181.140 ;
        RECT 90.405 180.800 92.000 180.940 ;
        RECT 93.625 180.940 93.915 180.985 ;
        RECT 94.530 180.940 94.850 181.000 ;
        RECT 114.770 180.940 115.090 181.000 ;
        RECT 93.625 180.800 115.090 180.940 ;
        RECT 116.700 180.940 116.840 181.420 ;
        RECT 129.950 181.280 130.270 181.340 ;
        RECT 138.780 181.325 138.920 181.480 ;
        RECT 141.450 181.420 141.770 181.480 ;
        RECT 143.765 181.620 144.055 181.665 ;
        RECT 145.590 181.620 145.910 181.680 ;
        RECT 143.765 181.480 145.910 181.620 ;
        RECT 143.765 181.435 144.055 181.480 ;
        RECT 145.590 181.420 145.910 181.480 ;
        RECT 146.050 181.420 146.370 181.680 ;
        RECT 129.950 181.140 135.240 181.280 ;
        RECT 129.950 181.080 130.270 181.140 ;
        RECT 120.765 180.940 121.055 180.985 ;
        RECT 116.700 180.800 121.055 180.940 ;
        RECT 90.405 180.755 90.695 180.800 ;
        RECT 93.625 180.755 93.915 180.800 ;
        RECT 94.530 180.740 94.850 180.800 ;
        RECT 114.770 180.740 115.090 180.800 ;
        RECT 120.765 180.755 121.055 180.800 ;
        RECT 126.270 180.940 126.590 181.000 ;
        RECT 129.045 180.940 129.335 180.985 ;
        RECT 126.270 180.800 129.335 180.940 ;
        RECT 126.270 180.740 126.590 180.800 ;
        RECT 129.045 180.755 129.335 180.800 ;
        RECT 131.330 180.740 131.650 181.000 ;
        RECT 132.250 180.740 132.570 181.000 ;
        RECT 134.565 180.940 134.855 180.985 ;
        RECT 133.260 180.800 134.855 180.940 ;
        RECT 135.100 180.940 135.240 181.140 ;
        RECT 138.705 181.095 138.995 181.325 ;
        RECT 143.290 181.280 143.610 181.340 ;
        RECT 139.700 181.140 143.610 181.280 ;
        RECT 137.785 180.940 138.075 180.985 ;
        RECT 135.100 180.800 138.075 180.940 ;
        RECT 64.170 180.600 64.490 180.660 ;
        RECT 65.105 180.600 65.395 180.645 ;
        RECT 59.200 180.460 59.800 180.600 ;
        RECT 30.220 180.120 34.040 180.260 ;
        RECT 34.310 180.260 34.600 180.305 ;
        RECT 36.410 180.260 36.700 180.305 ;
        RECT 37.980 180.260 38.270 180.305 ;
        RECT 34.310 180.120 38.270 180.260 ;
        RECT 59.660 180.260 59.800 180.460 ;
        RECT 64.170 180.460 65.395 180.600 ;
        RECT 64.170 180.400 64.490 180.460 ;
        RECT 65.105 180.415 65.395 180.460 ;
        RECT 76.565 180.600 76.855 180.645 ;
        RECT 77.755 180.600 78.045 180.645 ;
        RECT 80.275 180.600 80.565 180.645 ;
        RECT 76.565 180.460 80.565 180.600 ;
        RECT 76.565 180.415 76.855 180.460 ;
        RECT 77.755 180.415 78.045 180.460 ;
        RECT 80.275 180.415 80.565 180.460 ;
        RECT 94.990 180.400 95.310 180.660 ;
        RECT 105.110 180.600 105.430 180.660 ;
        RECT 108.790 180.600 109.110 180.660 ;
        RECT 105.110 180.460 109.110 180.600 ;
        RECT 105.110 180.400 105.430 180.460 ;
        RECT 108.790 180.400 109.110 180.460 ;
        RECT 109.685 180.600 109.975 180.645 ;
        RECT 110.875 180.600 111.165 180.645 ;
        RECT 113.395 180.600 113.685 180.645 ;
        RECT 109.685 180.460 113.685 180.600 ;
        RECT 109.685 180.415 109.975 180.460 ;
        RECT 110.875 180.415 111.165 180.460 ;
        RECT 113.395 180.415 113.685 180.460 ;
        RECT 128.570 180.400 128.890 180.660 ;
        RECT 129.965 180.600 130.255 180.645 ;
        RECT 130.885 180.600 131.175 180.645 ;
        RECT 129.965 180.460 131.175 180.600 ;
        RECT 129.965 180.415 130.255 180.460 ;
        RECT 130.885 180.415 131.175 180.460 ;
        RECT 131.790 180.400 132.110 180.660 ;
        RECT 133.260 180.645 133.400 180.800 ;
        RECT 134.565 180.755 134.855 180.800 ;
        RECT 137.785 180.755 138.075 180.800 ;
        RECT 139.165 180.755 139.455 180.985 ;
        RECT 133.185 180.415 133.475 180.645 ;
        RECT 133.645 180.415 133.935 180.645 ;
        RECT 134.640 180.600 134.780 180.755 ;
        RECT 135.470 180.600 135.790 180.660 ;
        RECT 134.640 180.460 135.790 180.600 ;
        RECT 137.860 180.600 138.000 180.755 ;
        RECT 138.690 180.600 139.010 180.660 ;
        RECT 139.240 180.600 139.380 180.755 ;
        RECT 137.860 180.460 139.380 180.600 ;
        RECT 68.310 180.260 68.630 180.320 ;
        RECT 59.660 180.120 68.630 180.260 ;
        RECT 24.650 180.075 24.940 180.120 ;
        RECT 26.750 180.075 27.040 180.120 ;
        RECT 28.320 180.075 28.610 180.120 ;
        RECT 34.310 180.075 34.600 180.120 ;
        RECT 36.410 180.075 36.700 180.120 ;
        RECT 37.980 180.075 38.270 180.120 ;
        RECT 68.310 180.060 68.630 180.120 ;
        RECT 69.245 180.260 69.535 180.305 ;
        RECT 71.530 180.260 71.850 180.320 ;
        RECT 69.245 180.120 71.850 180.260 ;
        RECT 69.245 180.075 69.535 180.120 ;
        RECT 71.530 180.060 71.850 180.120 ;
        RECT 76.170 180.260 76.460 180.305 ;
        RECT 78.270 180.260 78.560 180.305 ;
        RECT 79.840 180.260 80.130 180.305 ;
        RECT 109.290 180.260 109.580 180.305 ;
        RECT 111.390 180.260 111.680 180.305 ;
        RECT 112.960 180.260 113.250 180.305 ;
        RECT 133.720 180.260 133.860 180.415 ;
        RECT 135.470 180.400 135.790 180.460 ;
        RECT 138.690 180.400 139.010 180.460 ;
        RECT 139.700 180.260 139.840 181.140 ;
        RECT 143.290 181.080 143.610 181.140 ;
        RECT 144.210 181.280 144.530 181.340 ;
        RECT 144.210 181.140 146.740 181.280 ;
        RECT 144.210 181.080 144.530 181.140 ;
        RECT 140.085 180.940 140.375 180.985 ;
        RECT 141.450 180.940 141.770 181.000 ;
        RECT 140.085 180.800 141.770 180.940 ;
        RECT 140.085 180.755 140.375 180.800 ;
        RECT 141.450 180.740 141.770 180.800 ;
        RECT 145.130 180.740 145.450 181.000 ;
        RECT 146.600 180.985 146.740 181.140 ;
        RECT 146.525 180.940 146.815 180.985 ;
        RECT 149.270 180.940 149.590 181.000 ;
        RECT 146.525 180.800 149.590 180.940 ;
        RECT 146.525 180.755 146.815 180.800 ;
        RECT 149.270 180.740 149.590 180.800 ;
        RECT 146.970 180.600 147.290 180.660 ;
        RECT 150.205 180.600 150.495 180.645 ;
        RECT 146.970 180.460 150.495 180.600 ;
        RECT 146.970 180.400 147.290 180.460 ;
        RECT 150.205 180.415 150.495 180.460 ;
        RECT 76.170 180.120 80.130 180.260 ;
        RECT 76.170 180.075 76.460 180.120 ;
        RECT 78.270 180.075 78.560 180.120 ;
        RECT 79.840 180.075 80.130 180.120 ;
        RECT 81.970 180.120 84.180 180.260 ;
        RECT 31.050 179.720 31.370 179.980 ;
        RECT 33.350 179.720 33.670 179.980 ;
        RECT 43.010 179.920 43.330 179.980 ;
        RECT 45.785 179.920 46.075 179.965 ;
        RECT 43.010 179.780 46.075 179.920 ;
        RECT 43.010 179.720 43.330 179.780 ;
        RECT 45.785 179.735 46.075 179.780 ;
        RECT 57.730 179.720 58.050 179.980 ;
        RECT 74.750 179.920 75.070 179.980 ;
        RECT 81.970 179.920 82.110 180.120 ;
        RECT 74.750 179.780 82.110 179.920 ;
        RECT 82.585 179.920 82.875 179.965 ;
        RECT 83.490 179.920 83.810 179.980 ;
        RECT 84.040 179.965 84.180 180.120 ;
        RECT 109.290 180.120 113.250 180.260 ;
        RECT 109.290 180.075 109.580 180.120 ;
        RECT 111.390 180.075 111.680 180.120 ;
        RECT 112.960 180.075 113.250 180.120 ;
        RECT 130.270 180.120 133.860 180.260 ;
        RECT 135.560 180.120 139.840 180.260 ;
        RECT 82.585 179.780 83.810 179.920 ;
        RECT 74.750 179.720 75.070 179.780 ;
        RECT 82.585 179.735 82.875 179.780 ;
        RECT 83.490 179.720 83.810 179.780 ;
        RECT 83.965 179.735 84.255 179.965 ;
        RECT 108.330 179.920 108.650 179.980 ;
        RECT 130.270 179.920 130.410 180.120 ;
        RECT 135.560 179.965 135.700 180.120 ;
        RECT 108.330 179.780 130.410 179.920 ;
        RECT 108.330 179.720 108.650 179.780 ;
        RECT 135.485 179.735 135.775 179.965 ;
        RECT 138.230 179.920 138.550 179.980 ;
        RECT 139.625 179.920 139.915 179.965 ;
        RECT 140.070 179.920 140.390 179.980 ;
        RECT 138.230 179.780 140.390 179.920 ;
        RECT 138.230 179.720 138.550 179.780 ;
        RECT 139.625 179.735 139.915 179.780 ;
        RECT 140.070 179.720 140.390 179.780 ;
        RECT 22.700 179.100 157.020 179.580 ;
        RECT 25.085 178.900 25.375 178.945 ;
        RECT 25.530 178.900 25.850 178.960 ;
        RECT 25.085 178.760 25.850 178.900 ;
        RECT 25.085 178.715 25.375 178.760 ;
        RECT 25.530 178.700 25.850 178.760 ;
        RECT 29.225 178.900 29.515 178.945 ;
        RECT 29.670 178.900 29.990 178.960 ;
        RECT 29.225 178.760 29.990 178.900 ;
        RECT 29.225 178.715 29.515 178.760 ;
        RECT 29.670 178.700 29.990 178.760 ;
        RECT 32.890 178.700 33.210 178.960 ;
        RECT 33.825 178.900 34.115 178.945 ;
        RECT 34.270 178.900 34.590 178.960 ;
        RECT 33.825 178.760 34.590 178.900 ;
        RECT 33.825 178.715 34.115 178.760 ;
        RECT 34.270 178.700 34.590 178.760 ;
        RECT 40.710 178.700 41.030 178.960 ;
        RECT 42.565 178.900 42.855 178.945 ;
        RECT 45.310 178.900 45.630 178.960 ;
        RECT 42.565 178.760 45.630 178.900 ;
        RECT 42.565 178.715 42.855 178.760 ;
        RECT 45.310 178.700 45.630 178.760 ;
        RECT 46.245 178.900 46.535 178.945 ;
        RECT 46.690 178.900 47.010 178.960 ;
        RECT 46.245 178.760 47.010 178.900 ;
        RECT 46.245 178.715 46.535 178.760 ;
        RECT 46.690 178.700 47.010 178.760 ;
        RECT 67.850 178.700 68.170 178.960 ;
        RECT 70.165 178.900 70.455 178.945 ;
        RECT 70.610 178.900 70.930 178.960 ;
        RECT 70.165 178.760 70.930 178.900 ;
        RECT 70.165 178.715 70.455 178.760 ;
        RECT 70.610 178.700 70.930 178.760 ;
        RECT 76.130 178.900 76.450 178.960 ;
        RECT 77.525 178.900 77.815 178.945 ;
        RECT 76.130 178.760 77.815 178.900 ;
        RECT 76.130 178.700 76.450 178.760 ;
        RECT 77.525 178.715 77.815 178.760 ;
        RECT 92.690 178.700 93.010 178.960 ;
        RECT 97.290 178.900 97.610 178.960 ;
        RECT 98.670 178.900 98.990 178.960 ;
        RECT 130.425 178.900 130.715 178.945 ;
        RECT 131.790 178.900 132.110 178.960 ;
        RECT 96.460 178.760 108.560 178.900 ;
        RECT 51.290 178.560 51.580 178.605 ;
        RECT 52.860 178.560 53.150 178.605 ;
        RECT 54.960 178.560 55.250 178.605 ;
        RECT 51.290 178.420 55.250 178.560 ;
        RECT 51.290 178.375 51.580 178.420 ;
        RECT 52.860 178.375 53.150 178.420 ;
        RECT 54.960 178.375 55.250 178.420 ;
        RECT 63.750 178.560 64.040 178.605 ;
        RECT 65.850 178.560 66.140 178.605 ;
        RECT 67.420 178.560 67.710 178.605 ;
        RECT 63.750 178.420 67.710 178.560 ;
        RECT 67.940 178.560 68.080 178.700 ;
        RECT 71.110 178.560 71.400 178.605 ;
        RECT 73.210 178.560 73.500 178.605 ;
        RECT 74.780 178.560 75.070 178.605 ;
        RECT 67.940 178.420 70.380 178.560 ;
        RECT 63.750 178.375 64.040 178.420 ;
        RECT 65.850 178.375 66.140 178.420 ;
        RECT 67.420 178.375 67.710 178.420 ;
        RECT 70.240 178.280 70.380 178.420 ;
        RECT 71.110 178.420 75.070 178.560 ;
        RECT 71.110 178.375 71.400 178.420 ;
        RECT 73.210 178.375 73.500 178.420 ;
        RECT 74.780 178.375 75.070 178.420 ;
        RECT 80.310 178.560 80.600 178.605 ;
        RECT 82.410 178.560 82.700 178.605 ;
        RECT 83.980 178.560 84.270 178.605 ;
        RECT 80.310 178.420 84.270 178.560 ;
        RECT 80.310 178.375 80.600 178.420 ;
        RECT 82.410 178.375 82.700 178.420 ;
        RECT 83.980 178.375 84.270 178.420 ;
        RECT 32.890 178.020 33.210 178.280 ;
        RECT 33.810 178.220 34.130 178.280 ;
        RECT 34.745 178.220 35.035 178.265 ;
        RECT 35.190 178.220 35.510 178.280 ;
        RECT 33.810 178.080 35.510 178.220 ;
        RECT 33.810 178.020 34.130 178.080 ;
        RECT 34.745 178.035 35.035 178.080 ;
        RECT 35.190 178.020 35.510 178.080 ;
        RECT 44.850 178.020 45.170 178.280 ;
        RECT 50.855 178.220 51.145 178.265 ;
        RECT 53.375 178.220 53.665 178.265 ;
        RECT 54.565 178.220 54.855 178.265 ;
        RECT 61.870 178.220 62.190 178.280 ;
        RECT 50.855 178.080 54.855 178.220 ;
        RECT 50.855 178.035 51.145 178.080 ;
        RECT 53.375 178.035 53.665 178.080 ;
        RECT 54.565 178.035 54.855 178.080 ;
        RECT 57.360 178.080 62.190 178.220 ;
        RECT 26.005 177.880 26.295 177.925 ;
        RECT 31.050 177.880 31.370 177.940 ;
        RECT 32.980 177.880 33.120 178.020 ;
        RECT 34.285 177.880 34.575 177.925 ;
        RECT 26.005 177.740 28.520 177.880 ;
        RECT 26.005 177.695 26.295 177.740 ;
        RECT 28.380 177.245 28.520 177.740 ;
        RECT 31.050 177.740 34.575 177.880 ;
        RECT 31.050 177.680 31.370 177.740 ;
        RECT 34.285 177.695 34.575 177.740 ;
        RECT 37.490 177.880 37.810 177.940 ;
        RECT 40.265 177.880 40.555 177.925 ;
        RECT 37.490 177.740 40.555 177.880 ;
        RECT 37.490 177.680 37.810 177.740 ;
        RECT 40.265 177.695 40.555 177.740 ;
        RECT 29.210 177.585 29.530 177.600 ;
        RECT 29.145 177.355 29.530 177.585 ;
        RECT 29.210 177.340 29.530 177.355 ;
        RECT 30.130 177.540 30.450 177.600 ;
        RECT 33.350 177.585 33.670 177.600 ;
        RECT 31.985 177.540 32.275 177.585 ;
        RECT 30.130 177.400 32.275 177.540 ;
        RECT 30.130 177.340 30.450 177.400 ;
        RECT 31.985 177.355 32.275 177.400 ;
        RECT 33.065 177.355 33.670 177.585 ;
        RECT 40.340 177.540 40.480 177.695 ;
        RECT 44.390 177.680 44.710 177.940 ;
        RECT 44.940 177.880 45.080 178.020 ;
        RECT 57.360 177.940 57.500 178.080 ;
        RECT 61.870 178.020 62.190 178.080 ;
        RECT 64.145 178.220 64.435 178.265 ;
        RECT 65.335 178.220 65.625 178.265 ;
        RECT 67.855 178.220 68.145 178.265 ;
        RECT 64.145 178.080 68.145 178.220 ;
        RECT 64.145 178.035 64.435 178.080 ;
        RECT 65.335 178.035 65.625 178.080 ;
        RECT 67.855 178.035 68.145 178.080 ;
        RECT 70.150 178.020 70.470 178.280 ;
        RECT 71.505 178.220 71.795 178.265 ;
        RECT 72.695 178.220 72.985 178.265 ;
        RECT 75.215 178.220 75.505 178.265 ;
        RECT 71.505 178.080 75.505 178.220 ;
        RECT 71.505 178.035 71.795 178.080 ;
        RECT 72.695 178.035 72.985 178.080 ;
        RECT 75.215 178.035 75.505 178.080 ;
        RECT 75.670 178.220 75.990 178.280 ;
        RECT 79.825 178.220 80.115 178.265 ;
        RECT 75.670 178.080 80.115 178.220 ;
        RECT 75.670 178.020 75.990 178.080 ;
        RECT 79.825 178.035 80.115 178.080 ;
        RECT 80.705 178.220 80.995 178.265 ;
        RECT 81.895 178.220 82.185 178.265 ;
        RECT 84.415 178.220 84.705 178.265 ;
        RECT 80.705 178.080 84.705 178.220 ;
        RECT 80.705 178.035 80.995 178.080 ;
        RECT 81.895 178.035 82.185 178.080 ;
        RECT 84.415 178.035 84.705 178.080 ;
        RECT 86.710 178.220 87.030 178.280 ;
        RECT 88.105 178.220 88.395 178.265 ;
        RECT 86.710 178.080 88.395 178.220 ;
        RECT 86.710 178.020 87.030 178.080 ;
        RECT 88.105 178.035 88.395 178.080 ;
        RECT 91.325 178.220 91.615 178.265 ;
        RECT 91.325 178.080 95.680 178.220 ;
        RECT 91.325 178.035 91.615 178.080 ;
        RECT 55.445 177.880 55.735 177.925 ;
        RECT 57.270 177.880 57.590 177.940 ;
        RECT 44.940 177.740 54.740 177.880 ;
        RECT 50.830 177.540 51.150 177.600 ;
        RECT 54.110 177.540 54.400 177.585 ;
        RECT 40.340 177.400 48.760 177.540 ;
        RECT 33.350 177.340 33.670 177.355 ;
        RECT 48.620 177.245 48.760 177.400 ;
        RECT 50.830 177.400 54.400 177.540 ;
        RECT 54.600 177.540 54.740 177.740 ;
        RECT 55.445 177.740 57.590 177.880 ;
        RECT 55.445 177.695 55.735 177.740 ;
        RECT 57.270 177.680 57.590 177.740 ;
        RECT 59.110 177.680 59.430 177.940 ;
        RECT 63.265 177.880 63.555 177.925 ;
        RECT 67.390 177.880 67.710 177.940 ;
        RECT 70.625 177.880 70.915 177.925 ;
        RECT 63.265 177.740 71.300 177.880 ;
        RECT 63.265 177.695 63.555 177.740 ;
        RECT 67.390 177.680 67.710 177.740 ;
        RECT 70.625 177.695 70.915 177.740 ;
        RECT 63.710 177.540 64.030 177.600 ;
        RECT 54.600 177.400 64.030 177.540 ;
        RECT 50.830 177.340 51.150 177.400 ;
        RECT 54.110 177.355 54.400 177.400 ;
        RECT 63.710 177.340 64.030 177.400 ;
        RECT 64.600 177.540 64.890 177.585 ;
        RECT 66.470 177.540 66.790 177.600 ;
        RECT 64.600 177.400 66.790 177.540 ;
        RECT 64.600 177.355 64.890 177.400 ;
        RECT 66.470 177.340 66.790 177.400 ;
        RECT 28.305 177.015 28.595 177.245 ;
        RECT 48.545 177.200 48.835 177.245 ;
        RECT 51.290 177.200 51.610 177.260 ;
        RECT 48.545 177.060 51.610 177.200 ;
        RECT 48.545 177.015 48.835 177.060 ;
        RECT 51.290 177.000 51.610 177.060 ;
        RECT 53.590 177.200 53.910 177.260 ;
        RECT 55.905 177.200 56.195 177.245 ;
        RECT 53.590 177.060 56.195 177.200 ;
        RECT 71.160 177.200 71.300 177.740 ;
        RECT 71.960 177.695 72.250 177.925 ;
        RECT 89.930 177.880 90.250 177.940 ;
        RECT 92.230 177.880 92.550 177.940 ;
        RECT 93.150 177.880 93.470 177.940 ;
        RECT 95.005 177.880 95.295 177.925 ;
        RECT 89.930 177.740 92.765 177.880 ;
        RECT 71.530 177.540 71.850 177.600 ;
        RECT 72.080 177.540 72.220 177.695 ;
        RECT 89.930 177.680 90.250 177.740 ;
        RECT 92.230 177.680 92.765 177.740 ;
        RECT 93.150 177.740 95.295 177.880 ;
        RECT 93.150 177.680 93.470 177.740 ;
        RECT 95.005 177.695 95.295 177.740 ;
        RECT 71.530 177.400 72.220 177.540 ;
        RECT 81.160 177.540 81.450 177.585 ;
        RECT 83.030 177.540 83.350 177.600 ;
        RECT 81.160 177.400 83.350 177.540 ;
        RECT 92.475 177.525 92.765 177.680 ;
        RECT 93.625 177.540 93.915 177.585 ;
        RECT 95.540 177.540 95.680 178.080 ;
        RECT 96.460 177.925 96.600 178.760 ;
        RECT 97.290 178.700 97.610 178.760 ;
        RECT 98.670 178.700 98.990 178.760 ;
        RECT 108.420 178.620 108.560 178.760 ;
        RECT 130.425 178.760 132.110 178.900 ;
        RECT 130.425 178.715 130.715 178.760 ;
        RECT 131.790 178.700 132.110 178.760 ;
        RECT 135.485 178.715 135.775 178.945 ;
        RECT 138.690 178.900 139.010 178.960 ;
        RECT 140.085 178.900 140.375 178.945 ;
        RECT 138.690 178.760 140.375 178.900 ;
        RECT 100.090 178.560 100.380 178.605 ;
        RECT 102.190 178.560 102.480 178.605 ;
        RECT 103.760 178.560 104.050 178.605 ;
        RECT 100.090 178.420 104.050 178.560 ;
        RECT 100.090 178.375 100.380 178.420 ;
        RECT 102.190 178.375 102.480 178.420 ;
        RECT 103.760 178.375 104.050 178.420 ;
        RECT 108.330 178.360 108.650 178.620 ;
        RECT 108.790 178.360 109.110 178.620 ;
        RECT 110.185 178.560 110.475 178.605 ;
        RECT 110.630 178.560 110.950 178.620 ;
        RECT 110.185 178.420 110.950 178.560 ;
        RECT 110.185 178.375 110.475 178.420 ;
        RECT 110.630 178.360 110.950 178.420 ;
        RECT 117.110 178.560 117.400 178.605 ;
        RECT 119.210 178.560 119.500 178.605 ;
        RECT 120.780 178.560 121.070 178.605 ;
        RECT 117.110 178.420 121.070 178.560 ;
        RECT 117.110 178.375 117.400 178.420 ;
        RECT 119.210 178.375 119.500 178.420 ;
        RECT 120.780 178.375 121.070 178.420 ;
        RECT 129.965 178.560 130.255 178.605 ;
        RECT 130.870 178.560 131.190 178.620 ;
        RECT 129.965 178.420 131.190 178.560 ;
        RECT 129.965 178.375 130.255 178.420 ;
        RECT 130.870 178.360 131.190 178.420 ;
        RECT 97.305 178.220 97.595 178.265 ;
        RECT 97.750 178.220 98.070 178.280 ;
        RECT 97.305 178.080 98.070 178.220 ;
        RECT 97.305 178.035 97.595 178.080 ;
        RECT 97.750 178.020 98.070 178.080 ;
        RECT 100.485 178.220 100.775 178.265 ;
        RECT 101.675 178.220 101.965 178.265 ;
        RECT 104.195 178.220 104.485 178.265 ;
        RECT 108.420 178.220 108.560 178.360 ;
        RECT 100.485 178.080 104.485 178.220 ;
        RECT 100.485 178.035 100.775 178.080 ;
        RECT 101.675 178.035 101.965 178.080 ;
        RECT 104.195 178.035 104.485 178.080 ;
        RECT 107.960 178.080 108.560 178.220 ;
        RECT 108.880 178.220 109.020 178.360 ;
        RECT 116.625 178.220 116.915 178.265 ;
        RECT 108.880 178.080 116.915 178.220 ;
        RECT 96.385 177.695 96.675 177.925 ;
        RECT 98.210 177.680 98.530 177.940 ;
        RECT 99.590 177.880 99.910 177.940 ;
        RECT 105.110 177.880 105.430 177.940 ;
        RECT 107.960 177.925 108.100 178.080 ;
        RECT 116.625 178.035 116.915 178.080 ;
        RECT 117.505 178.220 117.795 178.265 ;
        RECT 118.695 178.220 118.985 178.265 ;
        RECT 121.215 178.220 121.505 178.265 ;
        RECT 135.560 178.220 135.700 178.715 ;
        RECT 138.690 178.700 139.010 178.760 ;
        RECT 140.085 178.715 140.375 178.760 ;
        RECT 141.005 178.375 141.295 178.605 ;
        RECT 148.850 178.560 149.140 178.605 ;
        RECT 150.950 178.560 151.240 178.605 ;
        RECT 152.520 178.560 152.810 178.605 ;
        RECT 148.850 178.420 152.810 178.560 ;
        RECT 148.850 178.375 149.140 178.420 ;
        RECT 150.950 178.375 151.240 178.420 ;
        RECT 152.520 178.375 152.810 178.420 ;
        RECT 117.505 178.080 121.505 178.220 ;
        RECT 117.505 178.035 117.795 178.080 ;
        RECT 118.695 178.035 118.985 178.080 ;
        RECT 121.215 178.035 121.505 178.080 ;
        RECT 130.270 178.080 135.700 178.220 ;
        RECT 136.405 178.220 136.695 178.265 ;
        RECT 141.080 178.220 141.220 178.375 ;
        RECT 136.405 178.080 141.220 178.220 ;
        RECT 99.590 177.740 105.430 177.880 ;
        RECT 99.590 177.680 99.910 177.740 ;
        RECT 105.110 177.680 105.430 177.740 ;
        RECT 107.885 177.695 108.175 177.925 ;
        RECT 108.345 177.695 108.635 177.925 ;
        RECT 109.710 177.880 110.030 177.940 ;
        RECT 110.185 177.880 110.475 177.925 ;
        RECT 109.710 177.740 110.475 177.880 ;
        RECT 100.830 177.540 101.120 177.585 ;
        RECT 108.420 177.540 108.560 177.695 ;
        RECT 109.710 177.680 110.030 177.740 ;
        RECT 110.185 177.695 110.475 177.740 ;
        RECT 111.565 177.695 111.855 177.925 ;
        RECT 71.530 177.340 71.850 177.400 ;
        RECT 81.160 177.355 81.450 177.400 ;
        RECT 83.030 177.340 83.350 177.400 ;
        RECT 93.625 177.400 95.680 177.540 ;
        RECT 99.220 177.400 101.120 177.540 ;
        RECT 93.625 177.355 93.915 177.400 ;
        RECT 75.670 177.200 75.990 177.260 ;
        RECT 71.160 177.060 75.990 177.200 ;
        RECT 53.590 177.000 53.910 177.060 ;
        RECT 55.905 177.015 56.195 177.060 ;
        RECT 75.670 177.000 75.990 177.060 ;
        RECT 86.710 177.000 87.030 177.260 ;
        RECT 87.170 177.200 87.490 177.260 ;
        RECT 91.785 177.200 92.075 177.245 ;
        RECT 87.170 177.060 92.075 177.200 ;
        RECT 87.170 177.000 87.490 177.060 ;
        RECT 91.785 177.015 92.075 177.060 ;
        RECT 94.070 177.000 94.390 177.260 ;
        RECT 95.450 177.000 95.770 177.260 ;
        RECT 99.220 177.245 99.360 177.400 ;
        RECT 100.830 177.355 101.120 177.400 ;
        RECT 106.580 177.400 108.560 177.540 ;
        RECT 111.640 177.540 111.780 177.695 ;
        RECT 115.230 177.680 115.550 177.940 ;
        RECT 130.270 177.880 130.410 178.080 ;
        RECT 136.405 178.035 136.695 178.080 ;
        RECT 115.780 177.740 130.410 177.880 ;
        RECT 135.025 177.880 135.315 177.925 ;
        RECT 135.470 177.880 135.790 177.940 ;
        RECT 135.025 177.740 135.790 177.880 ;
        RECT 112.010 177.540 112.330 177.600 ;
        RECT 115.780 177.540 115.920 177.740 ;
        RECT 135.025 177.695 135.315 177.740 ;
        RECT 135.470 177.680 135.790 177.740 ;
        RECT 117.850 177.540 118.140 177.585 ;
        RECT 111.640 177.400 115.920 177.540 ;
        RECT 116.240 177.400 118.140 177.540 ;
        RECT 99.145 177.015 99.435 177.245 ;
        RECT 104.650 177.200 104.970 177.260 ;
        RECT 106.580 177.245 106.720 177.400 ;
        RECT 112.010 177.340 112.330 177.400 ;
        RECT 106.505 177.200 106.795 177.245 ;
        RECT 104.650 177.060 106.795 177.200 ;
        RECT 104.650 177.000 104.970 177.060 ;
        RECT 106.505 177.015 106.795 177.060 ;
        RECT 106.950 177.000 107.270 177.260 ;
        RECT 116.240 177.245 116.380 177.400 ;
        RECT 117.850 177.355 118.140 177.400 ;
        RECT 126.730 177.540 127.050 177.600 ;
        RECT 128.125 177.540 128.415 177.585 ;
        RECT 128.570 177.540 128.890 177.600 ;
        RECT 126.730 177.400 128.890 177.540 ;
        RECT 126.730 177.340 127.050 177.400 ;
        RECT 128.125 177.355 128.415 177.400 ;
        RECT 128.570 177.340 128.890 177.400 ;
        RECT 138.690 177.540 139.010 177.600 ;
        RECT 140.070 177.585 140.390 177.600 ;
        RECT 139.165 177.540 139.455 177.585 ;
        RECT 138.690 177.400 139.455 177.540 ;
        RECT 138.690 177.340 139.010 177.400 ;
        RECT 139.165 177.355 139.455 177.400 ;
        RECT 140.070 177.355 140.455 177.585 ;
        RECT 141.080 177.540 141.220 178.080 ;
        RECT 142.370 178.220 142.690 178.280 ;
        RECT 149.245 178.220 149.535 178.265 ;
        RECT 150.435 178.220 150.725 178.265 ;
        RECT 152.955 178.220 153.245 178.265 ;
        RECT 142.370 178.080 145.360 178.220 ;
        RECT 142.370 178.020 142.690 178.080 ;
        RECT 141.465 177.880 141.755 177.925 ;
        RECT 141.910 177.880 142.230 177.940 ;
        RECT 141.465 177.740 142.230 177.880 ;
        RECT 141.465 177.695 141.755 177.740 ;
        RECT 141.910 177.680 142.230 177.740 ;
        RECT 142.845 177.880 143.135 177.925 ;
        RECT 143.290 177.880 143.610 177.940 ;
        RECT 144.210 177.925 144.530 177.940 ;
        RECT 145.220 177.925 145.360 178.080 ;
        RECT 149.245 178.080 153.245 178.220 ;
        RECT 149.245 178.035 149.535 178.080 ;
        RECT 150.435 178.035 150.725 178.080 ;
        RECT 152.955 178.035 153.245 178.080 ;
        RECT 144.175 177.880 144.530 177.925 ;
        RECT 142.845 177.740 143.610 177.880 ;
        RECT 142.845 177.695 143.135 177.740 ;
        RECT 143.290 177.680 143.610 177.740 ;
        RECT 143.840 177.740 144.530 177.880 ;
        RECT 143.840 177.540 143.980 177.740 ;
        RECT 144.175 177.695 144.530 177.740 ;
        RECT 145.145 177.695 145.435 177.925 ;
        RECT 145.605 177.695 145.895 177.925 ;
        RECT 144.210 177.680 144.530 177.695 ;
        RECT 141.080 177.400 143.980 177.540 ;
        RECT 140.070 177.340 140.390 177.355 ;
        RECT 145.680 177.260 145.820 177.695 ;
        RECT 146.510 177.680 146.830 177.940 ;
        RECT 146.970 177.880 147.290 177.940 ;
        RECT 148.365 177.880 148.655 177.925 ;
        RECT 146.970 177.740 148.655 177.880 ;
        RECT 146.970 177.680 147.290 177.740 ;
        RECT 148.365 177.695 148.655 177.740 ;
        RECT 149.700 177.540 149.990 177.585 ;
        RECT 150.190 177.540 150.510 177.600 ;
        RECT 149.700 177.400 150.510 177.540 ;
        RECT 149.700 177.355 149.990 177.400 ;
        RECT 150.190 177.340 150.510 177.400 ;
        RECT 116.165 177.015 116.455 177.245 ;
        RECT 123.525 177.200 123.815 177.245 ;
        RECT 124.430 177.200 124.750 177.260 ;
        RECT 123.525 177.060 124.750 177.200 ;
        RECT 123.525 177.015 123.815 177.060 ;
        RECT 124.430 177.000 124.750 177.060 ;
        RECT 136.850 177.200 137.170 177.260 ;
        RECT 137.785 177.200 138.075 177.245 ;
        RECT 136.850 177.060 138.075 177.200 ;
        RECT 136.850 177.000 137.170 177.060 ;
        RECT 137.785 177.015 138.075 177.060 ;
        RECT 141.450 177.200 141.770 177.260 ;
        RECT 141.925 177.200 142.215 177.245 ;
        RECT 141.450 177.060 142.215 177.200 ;
        RECT 141.450 177.000 141.770 177.060 ;
        RECT 141.925 177.015 142.215 177.060 ;
        RECT 143.750 177.000 144.070 177.260 ;
        RECT 145.145 177.200 145.435 177.245 ;
        RECT 145.590 177.200 145.910 177.260 ;
        RECT 145.145 177.060 145.910 177.200 ;
        RECT 145.145 177.015 145.435 177.060 ;
        RECT 145.590 177.000 145.910 177.060 ;
        RECT 146.525 177.200 146.815 177.245 ;
        RECT 148.810 177.200 149.130 177.260 ;
        RECT 146.525 177.060 149.130 177.200 ;
        RECT 146.525 177.015 146.815 177.060 ;
        RECT 148.810 177.000 149.130 177.060 ;
        RECT 154.330 177.200 154.650 177.260 ;
        RECT 155.265 177.200 155.555 177.245 ;
        RECT 154.330 177.060 155.555 177.200 ;
        RECT 154.330 177.000 154.650 177.060 ;
        RECT 155.265 177.015 155.555 177.060 ;
        RECT 22.700 176.380 157.820 176.860 ;
        RECT 50.830 175.980 51.150 176.240 ;
        RECT 51.290 176.180 51.610 176.240 ;
        RECT 59.110 176.180 59.430 176.240 ;
        RECT 51.290 176.040 59.430 176.180 ;
        RECT 51.290 175.980 51.610 176.040 ;
        RECT 59.110 175.980 59.430 176.040 ;
        RECT 64.170 175.980 64.490 176.240 ;
        RECT 66.470 175.980 66.790 176.240 ;
        RECT 69.690 176.180 70.010 176.240 ;
        RECT 71.530 176.225 71.850 176.240 ;
        RECT 71.415 176.180 71.850 176.225 ;
        RECT 69.690 176.040 71.850 176.180 ;
        RECT 69.690 175.980 70.010 176.040 ;
        RECT 71.415 175.995 71.850 176.040 ;
        RECT 71.530 175.980 71.850 175.995 ;
        RECT 83.030 175.980 83.350 176.240 ;
        RECT 83.490 176.180 83.810 176.240 ;
        RECT 84.885 176.180 85.175 176.225 ;
        RECT 90.850 176.180 91.170 176.240 ;
        RECT 83.490 176.040 91.170 176.180 ;
        RECT 83.490 175.980 83.810 176.040 ;
        RECT 84.885 175.995 85.175 176.040 ;
        RECT 90.850 175.980 91.170 176.040 ;
        RECT 97.750 175.980 98.070 176.240 ;
        RECT 98.210 176.180 98.530 176.240 ;
        RECT 100.525 176.180 100.815 176.225 ;
        RECT 98.210 176.040 100.815 176.180 ;
        RECT 98.210 175.980 98.530 176.040 ;
        RECT 100.525 175.995 100.815 176.040 ;
        RECT 102.825 176.180 103.115 176.225 ;
        RECT 106.950 176.180 107.270 176.240 ;
        RECT 102.825 176.040 107.270 176.180 ;
        RECT 102.825 175.995 103.115 176.040 ;
        RECT 106.950 175.980 107.270 176.040 ;
        RECT 115.230 176.180 115.550 176.240 ;
        RECT 117.545 176.180 117.835 176.225 ;
        RECT 115.230 176.040 117.835 176.180 ;
        RECT 115.230 175.980 115.550 176.040 ;
        RECT 117.545 175.995 117.835 176.040 ;
        RECT 130.425 176.180 130.715 176.225 ;
        RECT 130.870 176.180 131.190 176.240 ;
        RECT 137.785 176.180 138.075 176.225 ;
        RECT 141.450 176.180 141.770 176.240 ;
        RECT 130.425 176.040 131.190 176.180 ;
        RECT 130.425 175.995 130.715 176.040 ;
        RECT 130.870 175.980 131.190 176.040 ;
        RECT 136.480 176.040 141.770 176.180 ;
        RECT 32.890 175.840 33.210 175.900 ;
        RECT 28.840 175.700 33.210 175.840 ;
        RECT 28.840 175.545 28.980 175.700 ;
        RECT 32.890 175.640 33.210 175.700 ;
        RECT 52.685 175.840 52.975 175.885 ;
        RECT 54.510 175.840 54.830 175.900 ;
        RECT 54.985 175.840 55.275 175.885 ;
        RECT 52.685 175.700 55.275 175.840 ;
        RECT 52.685 175.655 52.975 175.700 ;
        RECT 54.510 175.640 54.830 175.700 ;
        RECT 54.985 175.655 55.275 175.700 ;
        RECT 55.445 175.840 55.735 175.885 ;
        RECT 57.730 175.840 58.050 175.900 ;
        RECT 58.510 175.840 58.800 175.885 ;
        RECT 55.445 175.700 57.500 175.840 ;
        RECT 55.445 175.655 55.735 175.700 ;
        RECT 28.765 175.315 29.055 175.545 ;
        RECT 29.685 175.500 29.975 175.545 ;
        RECT 31.065 175.500 31.355 175.545 ;
        RECT 31.510 175.500 31.830 175.560 ;
        RECT 29.685 175.360 30.360 175.500 ;
        RECT 29.685 175.315 29.975 175.360 ;
        RECT 29.210 174.280 29.530 174.540 ;
        RECT 30.220 174.525 30.360 175.360 ;
        RECT 31.065 175.360 31.830 175.500 ;
        RECT 31.065 175.315 31.355 175.360 ;
        RECT 31.510 175.300 31.830 175.360 ;
        RECT 34.270 175.300 34.590 175.560 ;
        RECT 43.930 175.300 44.250 175.560 ;
        RECT 51.765 175.315 52.055 175.545 ;
        RECT 52.225 175.315 52.515 175.545 ;
        RECT 30.590 175.160 30.910 175.220 ;
        RECT 31.985 175.160 32.275 175.205 ;
        RECT 44.020 175.160 44.160 175.300 ;
        RECT 30.590 175.020 44.160 175.160 ;
        RECT 30.590 174.960 30.910 175.020 ;
        RECT 31.985 174.975 32.275 175.020 ;
        RECT 37.950 174.820 38.270 174.880 ;
        RECT 47.150 174.820 47.470 174.880 ;
        RECT 37.950 174.680 47.470 174.820 ;
        RECT 51.840 174.820 51.980 175.315 ;
        RECT 52.300 175.160 52.440 175.315 ;
        RECT 53.590 175.300 53.910 175.560 ;
        RECT 54.050 175.300 54.370 175.560 ;
        RECT 55.890 175.300 56.210 175.560 ;
        RECT 57.360 175.500 57.500 175.700 ;
        RECT 57.730 175.700 58.800 175.840 ;
        RECT 57.730 175.640 58.050 175.700 ;
        RECT 58.510 175.655 58.800 175.700 ;
        RECT 72.465 175.840 72.755 175.885 ;
        RECT 74.765 175.840 75.055 175.885 ;
        RECT 87.170 175.840 87.490 175.900 ;
        RECT 99.590 175.840 99.910 175.900 ;
        RECT 129.030 175.840 129.350 175.900 ;
        RECT 136.480 175.840 136.620 176.040 ;
        RECT 137.785 175.995 138.075 176.040 ;
        RECT 141.450 175.980 141.770 176.040 ;
        RECT 141.910 175.980 142.230 176.240 ;
        RECT 147.445 176.180 147.735 176.225 ;
        RECT 148.905 176.180 149.195 176.225 ;
        RECT 149.730 176.180 150.050 176.240 ;
        RECT 147.445 176.040 150.050 176.180 ;
        RECT 147.445 175.995 147.735 176.040 ;
        RECT 148.905 175.995 149.195 176.040 ;
        RECT 149.730 175.980 150.050 176.040 ;
        RECT 150.190 175.980 150.510 176.240 ;
        RECT 72.465 175.700 75.055 175.840 ;
        RECT 72.465 175.655 72.755 175.700 ;
        RECT 74.765 175.655 75.055 175.700 ;
        RECT 84.040 175.700 87.490 175.840 ;
        RECT 60.030 175.500 60.350 175.560 ;
        RECT 61.410 175.500 61.730 175.560 ;
        RECT 57.360 175.360 61.730 175.500 ;
        RECT 60.030 175.300 60.350 175.360 ;
        RECT 61.410 175.300 61.730 175.360 ;
        RECT 66.930 175.500 67.250 175.560 ;
        RECT 67.405 175.500 67.695 175.545 ;
        RECT 66.930 175.360 67.695 175.500 ;
        RECT 66.930 175.300 67.250 175.360 ;
        RECT 67.405 175.315 67.695 175.360 ;
        RECT 68.310 175.300 68.630 175.560 ;
        RECT 68.785 175.500 69.075 175.545 ;
        RECT 70.150 175.500 70.470 175.560 ;
        RECT 68.785 175.360 70.470 175.500 ;
        RECT 68.785 175.315 69.075 175.360 ;
        RECT 70.150 175.300 70.470 175.360 ;
        RECT 75.670 175.500 75.990 175.560 ;
        RECT 84.040 175.545 84.180 175.700 ;
        RECT 87.170 175.640 87.490 175.700 ;
        RECT 90.940 175.700 99.910 175.840 ;
        RECT 79.365 175.500 79.655 175.545 ;
        RECT 75.670 175.360 79.655 175.500 ;
        RECT 75.670 175.300 75.990 175.360 ;
        RECT 79.365 175.315 79.655 175.360 ;
        RECT 83.965 175.315 84.255 175.545 ;
        RECT 56.810 175.160 57.130 175.220 ;
        RECT 52.300 175.020 57.130 175.160 ;
        RECT 56.810 174.960 57.130 175.020 ;
        RECT 57.270 174.960 57.590 175.220 ;
        RECT 58.165 175.160 58.455 175.205 ;
        RECT 59.355 175.160 59.645 175.205 ;
        RECT 61.875 175.160 62.165 175.205 ;
        RECT 58.165 175.020 62.165 175.160 ;
        RECT 68.400 175.160 68.540 175.300 ;
        RECT 71.070 175.160 71.390 175.220 ;
        RECT 77.525 175.160 77.815 175.205 ;
        RECT 68.400 175.020 69.000 175.160 ;
        RECT 58.165 174.975 58.455 175.020 ;
        RECT 59.355 174.975 59.645 175.020 ;
        RECT 61.875 174.975 62.165 175.020 ;
        RECT 54.970 174.820 55.290 174.880 ;
        RECT 55.890 174.820 56.210 174.880 ;
        RECT 51.840 174.680 56.210 174.820 ;
        RECT 37.950 174.620 38.270 174.680 ;
        RECT 47.150 174.620 47.470 174.680 ;
        RECT 54.970 174.620 55.290 174.680 ;
        RECT 55.890 174.620 56.210 174.680 ;
        RECT 57.770 174.820 58.060 174.865 ;
        RECT 59.870 174.820 60.160 174.865 ;
        RECT 61.440 174.820 61.730 174.865 ;
        RECT 57.770 174.680 61.730 174.820 ;
        RECT 68.860 174.820 69.000 175.020 ;
        RECT 71.070 175.020 77.815 175.160 ;
        RECT 71.070 174.960 71.390 175.020 ;
        RECT 77.525 174.975 77.815 175.020 ;
        RECT 74.750 174.820 75.070 174.880 ;
        RECT 68.860 174.680 75.070 174.820 ;
        RECT 57.770 174.635 58.060 174.680 ;
        RECT 59.870 174.635 60.160 174.680 ;
        RECT 61.440 174.635 61.730 174.680 ;
        RECT 74.750 174.620 75.070 174.680 ;
        RECT 78.430 174.620 78.750 174.880 ;
        RECT 79.440 174.820 79.580 175.315 ;
        RECT 85.330 175.300 85.650 175.560 ;
        RECT 90.940 175.545 91.080 175.700 ;
        RECT 99.590 175.640 99.910 175.700 ;
        RECT 115.320 175.700 122.820 175.840 ;
        RECT 90.865 175.315 91.155 175.545 ;
        RECT 92.200 175.500 92.490 175.545 ;
        RECT 94.070 175.500 94.390 175.560 ;
        RECT 92.200 175.360 94.390 175.500 ;
        RECT 92.200 175.315 92.490 175.360 ;
        RECT 94.070 175.300 94.390 175.360 ;
        RECT 94.990 175.500 95.310 175.560 ;
        RECT 100.970 175.500 101.290 175.560 ;
        RECT 115.320 175.545 115.460 175.700 ;
        RECT 102.365 175.500 102.655 175.545 ;
        RECT 108.805 175.500 109.095 175.545 ;
        RECT 115.245 175.500 115.535 175.545 ;
        RECT 119.385 175.500 119.675 175.545 ;
        RECT 94.990 175.360 100.280 175.500 ;
        RECT 94.990 175.300 95.310 175.360 ;
        RECT 91.745 175.160 92.035 175.205 ;
        RECT 92.935 175.160 93.225 175.205 ;
        RECT 95.455 175.160 95.745 175.205 ;
        RECT 91.745 175.020 95.745 175.160 ;
        RECT 100.140 175.160 100.280 175.360 ;
        RECT 100.970 175.360 102.655 175.500 ;
        RECT 100.970 175.300 101.290 175.360 ;
        RECT 102.365 175.315 102.655 175.360 ;
        RECT 107.500 175.360 115.535 175.500 ;
        RECT 101.890 175.160 102.210 175.220 ;
        RECT 103.285 175.160 103.575 175.205 ;
        RECT 100.140 175.020 103.575 175.160 ;
        RECT 91.745 174.975 92.035 175.020 ;
        RECT 92.935 174.975 93.225 175.020 ;
        RECT 95.455 174.975 95.745 175.020 ;
        RECT 101.890 174.960 102.210 175.020 ;
        RECT 103.285 174.975 103.575 175.020 ;
        RECT 91.350 174.820 91.640 174.865 ;
        RECT 93.450 174.820 93.740 174.865 ;
        RECT 95.020 174.820 95.310 174.865 ;
        RECT 79.440 174.680 91.080 174.820 ;
        RECT 30.145 174.480 30.435 174.525 ;
        RECT 33.350 174.480 33.670 174.540 ;
        RECT 30.145 174.340 33.670 174.480 ;
        RECT 30.145 174.295 30.435 174.340 ;
        RECT 33.350 174.280 33.670 174.340 ;
        RECT 33.810 174.280 34.130 174.540 ;
        RECT 40.710 174.480 41.030 174.540 ;
        RECT 41.645 174.480 41.935 174.525 ;
        RECT 40.710 174.340 41.935 174.480 ;
        RECT 40.710 174.280 41.030 174.340 ;
        RECT 41.645 174.295 41.935 174.340 ;
        RECT 43.485 174.480 43.775 174.525 ;
        RECT 44.390 174.480 44.710 174.540 ;
        RECT 43.485 174.340 44.710 174.480 ;
        RECT 43.485 174.295 43.775 174.340 ;
        RECT 44.390 174.280 44.710 174.340 ;
        RECT 56.825 174.480 57.115 174.525 ;
        RECT 63.710 174.480 64.030 174.540 ;
        RECT 56.825 174.340 64.030 174.480 ;
        RECT 56.825 174.295 57.115 174.340 ;
        RECT 63.710 174.280 64.030 174.340 ;
        RECT 70.610 174.280 70.930 174.540 ;
        RECT 71.545 174.480 71.835 174.525 ;
        RECT 74.290 174.480 74.610 174.540 ;
        RECT 71.545 174.340 74.610 174.480 ;
        RECT 78.520 174.480 78.660 174.620 ;
        RECT 84.870 174.480 85.190 174.540 ;
        RECT 88.550 174.480 88.870 174.540 ;
        RECT 78.520 174.340 88.870 174.480 ;
        RECT 90.940 174.480 91.080 174.680 ;
        RECT 91.350 174.680 95.310 174.820 ;
        RECT 91.350 174.635 91.640 174.680 ;
        RECT 93.450 174.635 93.740 174.680 ;
        RECT 95.020 174.635 95.310 174.680 ;
        RECT 102.350 174.480 102.670 174.540 ;
        RECT 107.500 174.480 107.640 175.360 ;
        RECT 108.805 175.315 109.095 175.360 ;
        RECT 115.245 175.315 115.535 175.360 ;
        RECT 115.780 175.360 119.675 175.500 ;
        RECT 109.725 175.160 110.015 175.205 ;
        RECT 110.630 175.160 110.950 175.220 ;
        RECT 109.725 175.020 110.950 175.160 ;
        RECT 109.725 174.975 110.015 175.020 ;
        RECT 110.630 174.960 110.950 175.020 ;
        RECT 114.770 175.160 115.090 175.220 ;
        RECT 115.780 175.160 115.920 175.360 ;
        RECT 119.385 175.315 119.675 175.360 ;
        RECT 119.845 175.500 120.135 175.545 ;
        RECT 121.685 175.500 121.975 175.545 ;
        RECT 119.845 175.360 121.975 175.500 ;
        RECT 119.845 175.315 120.135 175.360 ;
        RECT 121.685 175.315 121.975 175.360 ;
        RECT 122.130 175.500 122.450 175.560 ;
        RECT 122.680 175.545 122.820 175.700 ;
        RECT 124.520 175.700 127.880 175.840 ;
        RECT 124.520 175.560 124.660 175.700 ;
        RECT 122.605 175.500 122.895 175.545 ;
        RECT 122.130 175.360 122.895 175.500 ;
        RECT 122.130 175.300 122.450 175.360 ;
        RECT 122.605 175.315 122.895 175.360 ;
        RECT 123.525 175.500 123.815 175.545 ;
        RECT 124.430 175.500 124.750 175.560 ;
        RECT 123.525 175.360 124.750 175.500 ;
        RECT 123.525 175.315 123.815 175.360 ;
        RECT 124.430 175.300 124.750 175.360 ;
        RECT 124.890 175.500 125.210 175.560 ;
        RECT 127.740 175.545 127.880 175.700 ;
        RECT 128.200 175.700 136.620 175.840 ;
        RECT 128.200 175.545 128.340 175.700 ;
        RECT 129.030 175.640 129.350 175.700 ;
        RECT 136.850 175.640 137.170 175.900 ;
        RECT 142.370 175.840 142.690 175.900 ;
        RECT 143.305 175.840 143.595 175.885 ;
        RECT 142.370 175.700 143.595 175.840 ;
        RECT 142.370 175.640 142.690 175.700 ;
        RECT 143.305 175.655 143.595 175.700 ;
        RECT 144.210 175.640 144.530 175.900 ;
        RECT 146.050 175.840 146.370 175.900 ;
        RECT 147.890 175.840 148.210 175.900 ;
        RECT 153.885 175.840 154.175 175.885 ;
        RECT 146.050 175.700 148.210 175.840 ;
        RECT 146.050 175.640 146.370 175.700 ;
        RECT 147.890 175.640 148.210 175.700 ;
        RECT 148.440 175.700 154.175 175.840 ;
        RECT 126.745 175.500 127.035 175.545 ;
        RECT 124.890 175.360 127.035 175.500 ;
        RECT 124.890 175.300 125.210 175.360 ;
        RECT 126.745 175.315 127.035 175.360 ;
        RECT 127.665 175.315 127.955 175.545 ;
        RECT 128.125 175.315 128.415 175.545 ;
        RECT 129.505 175.500 129.795 175.545 ;
        RECT 130.870 175.500 131.190 175.560 ;
        RECT 129.505 175.360 131.190 175.500 ;
        RECT 129.505 175.315 129.795 175.360 ;
        RECT 130.870 175.300 131.190 175.360 ;
        RECT 138.230 175.300 138.550 175.560 ;
        RECT 145.590 175.300 145.910 175.560 ;
        RECT 146.510 175.500 146.830 175.560 ;
        RECT 148.440 175.500 148.580 175.700 ;
        RECT 153.885 175.655 154.175 175.700 ;
        RECT 151.125 175.500 151.415 175.545 ;
        RECT 146.510 175.360 148.580 175.500 ;
        RECT 149.820 175.360 151.415 175.500 ;
        RECT 146.510 175.300 146.830 175.360 ;
        RECT 114.770 175.020 115.920 175.160 ;
        RECT 116.165 175.160 116.455 175.205 ;
        RECT 118.910 175.160 119.230 175.220 ;
        RECT 116.165 175.020 119.230 175.160 ;
        RECT 114.770 174.960 115.090 175.020 ;
        RECT 116.165 174.975 116.455 175.020 ;
        RECT 118.910 174.960 119.230 175.020 ;
        RECT 120.290 174.960 120.610 175.220 ;
        RECT 123.970 175.160 124.290 175.220 ;
        RECT 128.585 175.160 128.875 175.205 ;
        RECT 130.410 175.160 130.730 175.220 ;
        RECT 123.970 175.020 130.730 175.160 ;
        RECT 123.970 174.960 124.290 175.020 ;
        RECT 128.585 174.975 128.875 175.020 ;
        RECT 130.410 174.960 130.730 175.020 ;
        RECT 136.405 174.975 136.695 175.205 ;
        RECT 136.480 174.820 136.620 174.975 ;
        RECT 138.690 174.960 139.010 175.220 ;
        RECT 146.600 175.160 146.740 175.300 ;
        RECT 142.045 175.020 146.740 175.160 ;
        RECT 136.865 174.820 137.155 174.865 ;
        RECT 136.480 174.680 137.155 174.820 ;
        RECT 136.865 174.635 137.155 174.680 ;
        RECT 90.940 174.340 107.640 174.480 ;
        RECT 71.545 174.295 71.835 174.340 ;
        RECT 74.290 174.280 74.610 174.340 ;
        RECT 84.870 174.280 85.190 174.340 ;
        RECT 88.550 174.280 88.870 174.340 ;
        RECT 102.350 174.280 102.670 174.340 ;
        RECT 107.870 174.280 108.190 174.540 ;
        RECT 114.310 174.280 114.630 174.540 ;
        RECT 133.170 174.280 133.490 174.540 ;
        RECT 136.390 174.480 136.710 174.540 ;
        RECT 142.045 174.480 142.185 175.020 ;
        RECT 149.820 174.865 149.960 175.360 ;
        RECT 151.125 175.315 151.415 175.360 ;
        RECT 154.330 175.300 154.650 175.560 ;
        RECT 149.745 174.635 150.035 174.865 ;
        RECT 136.390 174.340 142.185 174.480 ;
        RECT 136.390 174.280 136.710 174.340 ;
        RECT 142.370 174.280 142.690 174.540 ;
        RECT 148.810 174.280 149.130 174.540 ;
        RECT 22.700 173.660 157.020 174.140 ;
        RECT 26.005 173.460 26.295 173.505 ;
        RECT 27.845 173.460 28.135 173.505 ;
        RECT 26.005 173.320 28.135 173.460 ;
        RECT 26.005 173.275 26.295 173.320 ;
        RECT 27.845 173.275 28.135 173.320 ;
        RECT 31.510 173.260 31.830 173.520 ;
        RECT 32.890 173.460 33.210 173.520 ;
        RECT 33.825 173.460 34.115 173.505 ;
        RECT 43.930 173.460 44.250 173.520 ;
        RECT 32.890 173.320 34.115 173.460 ;
        RECT 32.890 173.260 33.210 173.320 ;
        RECT 33.825 173.275 34.115 173.320 ;
        RECT 37.580 173.320 44.250 173.460 ;
        RECT 26.925 173.120 27.215 173.165 ;
        RECT 24.240 172.980 27.215 173.120 ;
        RECT 24.240 172.485 24.380 172.980 ;
        RECT 26.925 172.935 27.215 172.980 ;
        RECT 30.130 173.120 30.450 173.180 ;
        RECT 32.445 173.120 32.735 173.165 ;
        RECT 30.130 172.980 32.735 173.120 ;
        RECT 30.130 172.920 30.450 172.980 ;
        RECT 32.445 172.935 32.735 172.980 ;
        RECT 33.810 172.780 34.130 172.840 ;
        RECT 26.540 172.640 34.130 172.780 ;
        RECT 26.540 172.485 26.680 172.640 ;
        RECT 33.810 172.580 34.130 172.640 ;
        RECT 24.165 172.255 24.455 172.485 ;
        RECT 25.545 172.255 25.835 172.485 ;
        RECT 26.465 172.255 26.755 172.485 ;
        RECT 29.685 172.440 29.975 172.485 ;
        RECT 37.045 172.440 37.335 172.485 ;
        RECT 37.580 172.440 37.720 173.320 ;
        RECT 43.930 173.260 44.250 173.320 ;
        RECT 44.405 173.460 44.695 173.505 ;
        RECT 44.865 173.460 45.155 173.505 ;
        RECT 44.405 173.320 45.155 173.460 ;
        RECT 44.405 173.275 44.695 173.320 ;
        RECT 44.865 173.275 45.155 173.320 ;
        RECT 45.770 173.460 46.090 173.520 ;
        RECT 46.690 173.460 47.010 173.520 ;
        RECT 45.770 173.320 47.010 173.460 ;
        RECT 44.480 173.120 44.620 173.275 ;
        RECT 45.770 173.260 46.090 173.320 ;
        RECT 46.690 173.260 47.010 173.320 ;
        RECT 54.050 173.460 54.370 173.520 ;
        RECT 61.885 173.460 62.175 173.505 ;
        RECT 54.050 173.320 62.175 173.460 ;
        RECT 54.050 173.260 54.370 173.320 ;
        RECT 61.885 173.275 62.175 173.320 ;
        RECT 71.070 173.460 71.390 173.520 ;
        RECT 74.305 173.460 74.595 173.505 ;
        RECT 71.070 173.320 74.595 173.460 ;
        RECT 71.070 173.260 71.390 173.320 ;
        RECT 74.305 173.275 74.595 173.320 ;
        RECT 83.505 173.460 83.795 173.505 ;
        RECT 84.410 173.460 84.730 173.520 ;
        RECT 88.550 173.460 88.870 173.520 ;
        RECT 92.690 173.460 93.010 173.520 ;
        RECT 83.505 173.320 88.320 173.460 ;
        RECT 83.505 173.275 83.795 173.320 ;
        RECT 84.410 173.260 84.730 173.320 ;
        RECT 40.340 172.980 44.620 173.120 ;
        RECT 47.650 173.120 47.940 173.165 ;
        RECT 49.750 173.120 50.040 173.165 ;
        RECT 51.320 173.120 51.610 173.165 ;
        RECT 47.650 172.980 51.610 173.120 ;
        RECT 29.685 172.300 33.120 172.440 ;
        RECT 29.685 172.255 29.975 172.300 ;
        RECT 25.620 172.100 25.760 172.255 ;
        RECT 29.210 172.100 29.530 172.160 ;
        RECT 25.620 171.960 29.530 172.100 ;
        RECT 29.210 171.900 29.530 171.960 ;
        RECT 30.590 171.900 30.910 172.160 ;
        RECT 25.085 171.760 25.375 171.805 ;
        RECT 25.530 171.760 25.850 171.820 ;
        RECT 25.085 171.620 25.850 171.760 ;
        RECT 25.085 171.575 25.375 171.620 ;
        RECT 25.530 171.560 25.850 171.620 ;
        RECT 27.370 171.760 27.690 171.820 ;
        RECT 31.510 171.805 31.830 171.820 ;
        RECT 27.845 171.760 28.135 171.805 ;
        RECT 27.370 171.620 28.135 171.760 ;
        RECT 27.370 171.560 27.690 171.620 ;
        RECT 27.845 171.575 28.135 171.620 ;
        RECT 31.510 171.575 31.895 171.805 ;
        RECT 32.430 171.760 32.750 171.820 ;
        RECT 32.980 171.805 33.120 172.300 ;
        RECT 37.045 172.300 37.720 172.440 ;
        RECT 37.045 172.255 37.335 172.300 ;
        RECT 38.870 172.240 39.190 172.500 ;
        RECT 39.330 172.240 39.650 172.500 ;
        RECT 40.340 172.485 40.480 172.980 ;
        RECT 47.650 172.935 47.940 172.980 ;
        RECT 49.750 172.935 50.040 172.980 ;
        RECT 51.320 172.935 51.610 172.980 ;
        RECT 55.890 173.120 56.210 173.180 ;
        RECT 57.730 173.120 58.050 173.180 ;
        RECT 55.890 172.980 58.050 173.120 ;
        RECT 55.890 172.920 56.210 172.980 ;
        RECT 57.730 172.920 58.050 172.980 ;
        RECT 67.890 173.120 68.180 173.165 ;
        RECT 69.990 173.120 70.280 173.165 ;
        RECT 71.560 173.120 71.850 173.165 ;
        RECT 67.890 172.980 71.850 173.120 ;
        RECT 67.890 172.935 68.180 172.980 ;
        RECT 69.990 172.935 70.280 172.980 ;
        RECT 71.560 172.935 71.850 172.980 ;
        RECT 77.090 173.120 77.380 173.165 ;
        RECT 79.190 173.120 79.480 173.165 ;
        RECT 80.760 173.120 81.050 173.165 ;
        RECT 77.090 172.980 81.050 173.120 ;
        RECT 88.180 173.120 88.320 173.320 ;
        RECT 88.550 173.320 93.010 173.460 ;
        RECT 88.550 173.260 88.870 173.320 ;
        RECT 92.690 173.260 93.010 173.320 ;
        RECT 93.150 173.260 93.470 173.520 ;
        RECT 110.630 173.460 110.950 173.520 ;
        RECT 123.970 173.460 124.290 173.520 ;
        RECT 138.245 173.460 138.535 173.505 ;
        RECT 138.690 173.460 139.010 173.520 ;
        RECT 110.630 173.320 124.290 173.460 ;
        RECT 110.630 173.260 110.950 173.320 ;
        RECT 123.970 173.260 124.290 173.320 ;
        RECT 125.900 173.320 131.100 173.460 ;
        RECT 89.945 173.120 90.235 173.165 ;
        RECT 90.850 173.120 91.170 173.180 ;
        RECT 88.180 172.980 89.700 173.120 ;
        RECT 77.090 172.935 77.380 172.980 ;
        RECT 79.190 172.935 79.480 172.980 ;
        RECT 80.760 172.935 81.050 172.980 ;
        RECT 42.550 172.780 42.870 172.840 ;
        RECT 42.550 172.640 46.000 172.780 ;
        RECT 42.550 172.580 42.870 172.640 ;
        RECT 39.805 172.255 40.095 172.485 ;
        RECT 40.265 172.255 40.555 172.485 ;
        RECT 33.350 172.145 33.670 172.160 ;
        RECT 33.350 172.100 33.955 172.145 ;
        RECT 34.270 172.100 34.590 172.160 ;
        RECT 34.745 172.100 35.035 172.145 ;
        RECT 33.350 171.960 34.105 172.100 ;
        RECT 34.270 171.960 35.035 172.100 ;
        RECT 33.350 171.915 33.955 171.960 ;
        RECT 33.350 171.900 33.670 171.915 ;
        RECT 34.270 171.900 34.590 171.960 ;
        RECT 34.745 171.915 35.035 171.960 ;
        RECT 37.505 171.915 37.795 172.145 ;
        RECT 38.410 172.100 38.730 172.160 ;
        RECT 39.880 172.100 40.020 172.255 ;
        RECT 41.630 172.240 41.950 172.500 ;
        RECT 43.025 172.440 43.315 172.485 ;
        RECT 42.180 172.300 43.315 172.440 ;
        RECT 42.180 172.100 42.320 172.300 ;
        RECT 43.025 172.255 43.315 172.300 ;
        RECT 43.485 172.440 43.775 172.485 ;
        RECT 44.390 172.440 44.710 172.500 ;
        RECT 43.485 172.300 44.710 172.440 ;
        RECT 43.485 172.255 43.775 172.300 ;
        RECT 38.410 171.960 40.020 172.100 ;
        RECT 40.340 171.960 42.320 172.100 ;
        RECT 32.905 171.760 33.195 171.805 ;
        RECT 32.430 171.620 33.195 171.760 ;
        RECT 37.580 171.760 37.720 171.915 ;
        RECT 38.410 171.900 38.730 171.960 ;
        RECT 40.340 171.760 40.480 171.960 ;
        RECT 42.550 171.900 42.870 172.160 ;
        RECT 37.580 171.620 40.480 171.760 ;
        RECT 41.185 171.760 41.475 171.805 ;
        RECT 43.010 171.760 43.330 171.820 ;
        RECT 41.185 171.620 43.330 171.760 ;
        RECT 44.020 171.760 44.160 172.300 ;
        RECT 44.390 172.240 44.710 172.300 ;
        RECT 44.850 172.240 45.170 172.500 ;
        RECT 45.310 172.240 45.630 172.500 ;
        RECT 45.860 172.440 46.000 172.640 ;
        RECT 47.150 172.580 47.470 172.840 ;
        RECT 48.045 172.780 48.335 172.825 ;
        RECT 49.235 172.780 49.525 172.825 ;
        RECT 51.755 172.780 52.045 172.825 ;
        RECT 48.045 172.640 52.045 172.780 ;
        RECT 48.045 172.595 48.335 172.640 ;
        RECT 49.235 172.595 49.525 172.640 ;
        RECT 51.755 172.595 52.045 172.640 ;
        RECT 52.300 172.640 59.340 172.780 ;
        RECT 52.300 172.440 52.440 172.640 ;
        RECT 59.200 172.500 59.340 172.640 ;
        RECT 67.390 172.580 67.710 172.840 ;
        RECT 68.285 172.780 68.575 172.825 ;
        RECT 69.475 172.780 69.765 172.825 ;
        RECT 71.995 172.780 72.285 172.825 ;
        RECT 68.285 172.640 72.285 172.780 ;
        RECT 68.285 172.595 68.575 172.640 ;
        RECT 69.475 172.595 69.765 172.640 ;
        RECT 71.995 172.595 72.285 172.640 ;
        RECT 72.450 172.780 72.770 172.840 ;
        RECT 74.290 172.780 74.610 172.840 ;
        RECT 74.765 172.780 75.055 172.825 ;
        RECT 72.450 172.640 75.055 172.780 ;
        RECT 72.450 172.580 72.770 172.640 ;
        RECT 74.290 172.580 74.610 172.640 ;
        RECT 74.765 172.595 75.055 172.640 ;
        RECT 77.485 172.780 77.775 172.825 ;
        RECT 78.675 172.780 78.965 172.825 ;
        RECT 81.195 172.780 81.485 172.825 ;
        RECT 77.485 172.640 81.485 172.780 ;
        RECT 77.485 172.595 77.775 172.640 ;
        RECT 78.675 172.595 78.965 172.640 ;
        RECT 81.195 172.595 81.485 172.640 ;
        RECT 45.860 172.300 52.440 172.440 ;
        RECT 58.665 172.255 58.955 172.485 ;
        RECT 59.110 172.440 59.430 172.500 ;
        RECT 64.645 172.440 64.935 172.485 ;
        RECT 59.110 172.300 64.935 172.440 ;
        RECT 48.500 172.100 48.790 172.145 ;
        RECT 52.210 172.100 52.530 172.160 ;
        RECT 58.740 172.100 58.880 172.255 ;
        RECT 59.110 172.240 59.430 172.300 ;
        RECT 64.645 172.255 64.935 172.300 ;
        RECT 75.670 172.240 75.990 172.500 ;
        RECT 76.590 172.240 76.910 172.500 ;
        RECT 83.950 172.240 84.270 172.500 ;
        RECT 85.345 172.440 85.635 172.485 ;
        RECT 86.710 172.440 87.030 172.500 ;
        RECT 85.345 172.300 87.030 172.440 ;
        RECT 85.345 172.255 85.635 172.300 ;
        RECT 86.710 172.240 87.030 172.300 ;
        RECT 48.500 171.960 52.530 172.100 ;
        RECT 48.500 171.915 48.790 171.960 ;
        RECT 52.210 171.900 52.530 171.960 ;
        RECT 54.140 171.960 58.880 172.100 ;
        RECT 68.740 172.100 69.030 172.145 ;
        RECT 69.690 172.100 70.010 172.160 ;
        RECT 68.740 171.960 70.010 172.100 ;
        RECT 54.140 171.805 54.280 171.960 ;
        RECT 68.740 171.915 69.030 171.960 ;
        RECT 69.690 171.900 70.010 171.960 ;
        RECT 77.940 172.100 78.230 172.145 ;
        RECT 78.890 172.100 79.210 172.160 ;
        RECT 77.940 171.960 79.210 172.100 ;
        RECT 77.940 171.915 78.230 171.960 ;
        RECT 78.890 171.900 79.210 171.960 ;
        RECT 79.350 172.100 79.670 172.160 ;
        RECT 89.560 172.145 89.700 172.980 ;
        RECT 89.945 172.980 91.170 173.120 ;
        RECT 89.945 172.935 90.235 172.980 ;
        RECT 90.850 172.920 91.170 172.980 ;
        RECT 94.990 173.120 95.310 173.180 ;
        RECT 104.230 173.120 104.520 173.165 ;
        RECT 106.330 173.120 106.620 173.165 ;
        RECT 107.900 173.120 108.190 173.165 ;
        RECT 94.990 172.980 96.140 173.120 ;
        RECT 94.990 172.920 95.310 172.980 ;
        RECT 95.450 172.580 95.770 172.840 ;
        RECT 96.000 172.825 96.140 172.980 ;
        RECT 104.230 172.980 108.190 173.120 ;
        RECT 104.230 172.935 104.520 172.980 ;
        RECT 106.330 172.935 106.620 172.980 ;
        RECT 107.900 172.935 108.190 172.980 ;
        RECT 113.890 173.120 114.180 173.165 ;
        RECT 115.990 173.120 116.280 173.165 ;
        RECT 117.560 173.120 117.850 173.165 ;
        RECT 113.890 172.980 117.850 173.120 ;
        RECT 113.890 172.935 114.180 172.980 ;
        RECT 115.990 172.935 116.280 172.980 ;
        RECT 117.560 172.935 117.850 172.980 ;
        RECT 118.910 173.120 119.230 173.180 ;
        RECT 120.305 173.120 120.595 173.165 ;
        RECT 121.670 173.120 121.990 173.180 ;
        RECT 125.900 173.120 126.040 173.320 ;
        RECT 118.910 172.980 121.990 173.120 ;
        RECT 118.910 172.920 119.230 172.980 ;
        RECT 120.305 172.935 120.595 172.980 ;
        RECT 121.670 172.920 121.990 172.980 ;
        RECT 124.060 172.980 126.040 173.120 ;
        RECT 95.925 172.595 96.215 172.825 ;
        RECT 96.370 172.780 96.690 172.840 ;
        RECT 103.745 172.780 104.035 172.825 ;
        RECT 96.370 172.640 104.035 172.780 ;
        RECT 96.370 172.580 96.690 172.640 ;
        RECT 103.745 172.595 104.035 172.640 ;
        RECT 104.625 172.780 104.915 172.825 ;
        RECT 105.815 172.780 106.105 172.825 ;
        RECT 108.335 172.780 108.625 172.825 ;
        RECT 104.625 172.640 108.625 172.780 ;
        RECT 104.625 172.595 104.915 172.640 ;
        RECT 105.815 172.595 106.105 172.640 ;
        RECT 108.335 172.595 108.625 172.640 ;
        RECT 108.790 172.780 109.110 172.840 ;
        RECT 113.405 172.780 113.695 172.825 ;
        RECT 108.790 172.640 113.695 172.780 ;
        RECT 108.790 172.580 109.110 172.640 ;
        RECT 113.405 172.595 113.695 172.640 ;
        RECT 114.285 172.780 114.575 172.825 ;
        RECT 115.475 172.780 115.765 172.825 ;
        RECT 117.995 172.780 118.285 172.825 ;
        RECT 124.060 172.780 124.200 172.980 ;
        RECT 126.270 172.920 126.590 173.180 ;
        RECT 126.730 172.920 127.050 173.180 ;
        RECT 114.285 172.640 118.285 172.780 ;
        RECT 114.285 172.595 114.575 172.640 ;
        RECT 115.475 172.595 115.765 172.640 ;
        RECT 117.995 172.595 118.285 172.640 ;
        RECT 123.600 172.640 124.200 172.780 ;
        RECT 124.430 172.780 124.750 172.840 ;
        RECT 124.430 172.640 128.800 172.780 ;
        RECT 90.865 172.440 91.155 172.485 ;
        RECT 91.310 172.440 91.630 172.500 ;
        RECT 90.865 172.300 91.630 172.440 ;
        RECT 90.865 172.255 91.155 172.300 ;
        RECT 91.310 172.240 91.630 172.300 ;
        RECT 102.365 172.440 102.655 172.485 ;
        RECT 104.190 172.440 104.510 172.500 ;
        RECT 102.365 172.300 104.510 172.440 ;
        RECT 102.365 172.255 102.655 172.300 ;
        RECT 104.190 172.240 104.510 172.300 ;
        RECT 111.550 172.240 111.870 172.500 ;
        RECT 121.685 172.440 121.975 172.485 ;
        RECT 122.130 172.440 122.450 172.500 ;
        RECT 123.600 172.485 123.740 172.640 ;
        RECT 124.430 172.580 124.750 172.640 ;
        RECT 121.685 172.300 122.450 172.440 ;
        RECT 121.685 172.255 121.975 172.300 ;
        RECT 122.130 172.240 122.450 172.300 ;
        RECT 122.605 172.255 122.895 172.485 ;
        RECT 123.525 172.255 123.815 172.485 ;
        RECT 79.350 171.960 87.860 172.100 ;
        RECT 79.350 171.900 79.670 171.960 ;
        RECT 54.065 171.760 54.355 171.805 ;
        RECT 44.020 171.620 54.355 171.760 ;
        RECT 31.510 171.560 31.830 171.575 ;
        RECT 32.430 171.560 32.750 171.620 ;
        RECT 32.905 171.575 33.195 171.620 ;
        RECT 41.185 171.575 41.475 171.620 ;
        RECT 43.010 171.560 43.330 171.620 ;
        RECT 54.065 171.575 54.355 171.620 ;
        RECT 54.970 171.760 55.290 171.820 ;
        RECT 55.905 171.760 56.195 171.805 ;
        RECT 54.970 171.620 56.195 171.760 ;
        RECT 54.970 171.560 55.290 171.620 ;
        RECT 55.905 171.575 56.195 171.620 ;
        RECT 56.810 171.760 57.130 171.820 ;
        RECT 58.650 171.760 58.970 171.820 ;
        RECT 56.810 171.620 58.970 171.760 ;
        RECT 56.810 171.560 57.130 171.620 ;
        RECT 58.650 171.560 58.970 171.620 ;
        RECT 70.150 171.760 70.470 171.820 ;
        RECT 80.270 171.760 80.590 171.820 ;
        RECT 82.110 171.760 82.430 171.820 ;
        RECT 84.425 171.760 84.715 171.805 ;
        RECT 85.330 171.760 85.650 171.820 ;
        RECT 87.720 171.805 87.860 171.960 ;
        RECT 89.485 171.915 89.775 172.145 ;
        RECT 98.210 172.100 98.530 172.160 ;
        RECT 100.065 172.100 100.355 172.145 ;
        RECT 101.430 172.100 101.750 172.160 ;
        RECT 104.970 172.100 105.260 172.145 ;
        RECT 114.630 172.100 114.920 172.145 ;
        RECT 98.210 171.960 101.750 172.100 ;
        RECT 98.210 171.900 98.530 171.960 ;
        RECT 100.065 171.915 100.355 171.960 ;
        RECT 101.430 171.900 101.750 171.960 ;
        RECT 103.360 171.960 105.260 172.100 ;
        RECT 70.150 171.620 85.650 171.760 ;
        RECT 70.150 171.560 70.470 171.620 ;
        RECT 80.270 171.560 80.590 171.620 ;
        RECT 82.110 171.560 82.430 171.620 ;
        RECT 84.425 171.575 84.715 171.620 ;
        RECT 85.330 171.560 85.650 171.620 ;
        RECT 87.645 171.575 87.935 171.805 ;
        RECT 88.485 171.760 88.775 171.805 ;
        RECT 92.230 171.760 92.550 171.820 ;
        RECT 88.485 171.620 92.550 171.760 ;
        RECT 88.485 171.575 88.775 171.620 ;
        RECT 92.230 171.560 92.550 171.620 ;
        RECT 94.990 171.560 95.310 171.820 ;
        RECT 99.130 171.760 99.450 171.820 ;
        RECT 103.360 171.805 103.500 171.960 ;
        RECT 104.970 171.915 105.260 171.960 ;
        RECT 112.560 171.960 114.920 172.100 ;
        RECT 122.680 172.100 122.820 172.255 ;
        RECT 124.890 172.240 125.210 172.500 ;
        RECT 125.350 172.240 125.670 172.500 ;
        RECT 128.660 172.485 128.800 172.640 ;
        RECT 129.030 172.485 129.350 172.500 ;
        RECT 127.435 172.440 127.725 172.485 ;
        RECT 125.900 172.300 127.725 172.440 ;
        RECT 124.430 172.100 124.750 172.160 ;
        RECT 125.900 172.100 126.040 172.300 ;
        RECT 127.435 172.255 127.725 172.300 ;
        RECT 128.585 172.255 128.875 172.485 ;
        RECT 129.030 172.255 129.515 172.485 ;
        RECT 129.965 172.255 130.255 172.485 ;
        RECT 129.030 172.240 129.350 172.255 ;
        RECT 122.680 171.960 126.040 172.100 ;
        RECT 112.560 171.805 112.700 171.960 ;
        RECT 114.630 171.915 114.920 171.960 ;
        RECT 124.430 171.900 124.750 171.960 ;
        RECT 128.110 171.900 128.430 172.160 ;
        RECT 100.525 171.760 100.815 171.805 ;
        RECT 99.130 171.620 100.815 171.760 ;
        RECT 99.130 171.560 99.450 171.620 ;
        RECT 100.525 171.575 100.815 171.620 ;
        RECT 103.285 171.575 103.575 171.805 ;
        RECT 112.485 171.575 112.775 171.805 ;
        RECT 120.750 171.560 121.070 171.820 ;
        RECT 125.350 171.760 125.670 171.820 ;
        RECT 129.490 171.760 129.810 171.820 ;
        RECT 130.040 171.760 130.180 172.255 ;
        RECT 130.960 171.820 131.100 173.320 ;
        RECT 138.245 173.320 139.010 173.460 ;
        RECT 138.245 173.275 138.535 173.320 ;
        RECT 138.690 173.260 139.010 173.320 ;
        RECT 139.150 173.460 139.470 173.520 ;
        RECT 140.085 173.460 140.375 173.505 ;
        RECT 141.910 173.460 142.230 173.520 ;
        RECT 139.150 173.320 142.230 173.460 ;
        RECT 139.150 173.260 139.470 173.320 ;
        RECT 140.085 173.275 140.375 173.320 ;
        RECT 141.910 173.260 142.230 173.320 ;
        RECT 131.830 173.120 132.120 173.165 ;
        RECT 133.930 173.120 134.220 173.165 ;
        RECT 135.500 173.120 135.790 173.165 ;
        RECT 131.830 172.980 135.790 173.120 ;
        RECT 131.830 172.935 132.120 172.980 ;
        RECT 133.930 172.935 134.220 172.980 ;
        RECT 135.500 172.935 135.790 172.980 ;
        RECT 142.830 173.120 143.120 173.165 ;
        RECT 144.400 173.120 144.690 173.165 ;
        RECT 146.500 173.120 146.790 173.165 ;
        RECT 142.830 172.980 146.790 173.120 ;
        RECT 142.830 172.935 143.120 172.980 ;
        RECT 144.400 172.935 144.690 172.980 ;
        RECT 146.500 172.935 146.790 172.980 ;
        RECT 132.225 172.780 132.515 172.825 ;
        RECT 133.415 172.780 133.705 172.825 ;
        RECT 135.935 172.780 136.225 172.825 ;
        RECT 132.225 172.640 136.225 172.780 ;
        RECT 132.225 172.595 132.515 172.640 ;
        RECT 133.415 172.595 133.705 172.640 ;
        RECT 135.935 172.595 136.225 172.640 ;
        RECT 142.395 172.780 142.685 172.825 ;
        RECT 144.915 172.780 145.205 172.825 ;
        RECT 146.105 172.780 146.395 172.825 ;
        RECT 142.395 172.640 146.395 172.780 ;
        RECT 142.395 172.595 142.685 172.640 ;
        RECT 144.915 172.595 145.205 172.640 ;
        RECT 146.105 172.595 146.395 172.640 ;
        RECT 147.445 172.780 147.735 172.825 ;
        RECT 147.890 172.780 148.210 172.840 ;
        RECT 147.445 172.640 148.210 172.780 ;
        RECT 147.445 172.595 147.735 172.640 ;
        RECT 147.890 172.580 148.210 172.640 ;
        RECT 131.345 172.440 131.635 172.485 ;
        RECT 146.970 172.440 147.290 172.500 ;
        RECT 131.345 172.300 147.290 172.440 ;
        RECT 131.345 172.255 131.635 172.300 ;
        RECT 146.970 172.240 147.290 172.300 ;
        RECT 149.730 172.240 150.050 172.500 ;
        RECT 153.410 172.240 153.730 172.500 ;
        RECT 132.680 172.100 132.970 172.145 ;
        RECT 133.170 172.100 133.490 172.160 ;
        RECT 132.680 171.960 133.490 172.100 ;
        RECT 132.680 171.915 132.970 171.960 ;
        RECT 133.170 171.900 133.490 171.960 ;
        RECT 143.750 172.100 144.070 172.160 ;
        RECT 145.650 172.100 145.940 172.145 ;
        RECT 149.285 172.100 149.575 172.145 ;
        RECT 152.965 172.100 153.255 172.145 ;
        RECT 143.750 171.960 145.940 172.100 ;
        RECT 143.750 171.900 144.070 171.960 ;
        RECT 145.650 171.915 145.940 171.960 ;
        RECT 146.140 171.960 153.255 172.100 ;
        RECT 125.350 171.620 130.180 171.760 ;
        RECT 130.870 171.760 131.190 171.820 ;
        RECT 146.140 171.760 146.280 171.960 ;
        RECT 149.285 171.915 149.575 171.960 ;
        RECT 152.965 171.915 153.255 171.960 ;
        RECT 130.870 171.620 146.280 171.760 ;
        RECT 125.350 171.560 125.670 171.620 ;
        RECT 129.490 171.560 129.810 171.620 ;
        RECT 130.870 171.560 131.190 171.620 ;
        RECT 148.810 171.560 149.130 171.820 ;
        RECT 22.700 170.940 157.820 171.420 ;
        RECT 31.065 170.740 31.355 170.785 ;
        RECT 34.270 170.740 34.590 170.800 ;
        RECT 31.065 170.600 34.590 170.740 ;
        RECT 31.065 170.555 31.355 170.600 ;
        RECT 34.270 170.540 34.590 170.600 ;
        RECT 34.745 170.740 35.035 170.785 ;
        RECT 37.965 170.740 38.255 170.785 ;
        RECT 38.870 170.740 39.190 170.800 ;
        RECT 34.745 170.600 37.720 170.740 ;
        RECT 34.745 170.555 35.035 170.600 ;
        RECT 33.810 170.400 34.130 170.460 ;
        RECT 36.585 170.400 36.875 170.445 ;
        RECT 33.810 170.260 36.875 170.400 ;
        RECT 33.810 170.200 34.130 170.260 ;
        RECT 36.585 170.215 36.875 170.260 ;
        RECT 25.530 170.105 25.850 170.120 ;
        RECT 25.500 170.060 25.850 170.105 ;
        RECT 25.335 169.920 25.850 170.060 ;
        RECT 25.500 169.875 25.850 169.920 ;
        RECT 32.445 170.060 32.735 170.105 ;
        RECT 32.890 170.060 33.210 170.120 ;
        RECT 32.445 169.920 33.210 170.060 ;
        RECT 32.445 169.875 32.735 169.920 ;
        RECT 25.530 169.860 25.850 169.875 ;
        RECT 32.890 169.860 33.210 169.920 ;
        RECT 35.190 169.860 35.510 170.120 ;
        RECT 36.125 169.875 36.415 170.105 ;
        RECT 37.045 169.875 37.335 170.105 ;
        RECT 37.580 170.060 37.720 170.600 ;
        RECT 37.965 170.600 39.190 170.740 ;
        RECT 37.965 170.555 38.255 170.600 ;
        RECT 38.870 170.540 39.190 170.600 ;
        RECT 40.265 170.740 40.555 170.785 ;
        RECT 45.310 170.740 45.630 170.800 ;
        RECT 40.265 170.600 45.630 170.740 ;
        RECT 40.265 170.555 40.555 170.600 ;
        RECT 45.310 170.540 45.630 170.600 ;
        RECT 52.210 170.540 52.530 170.800 ;
        RECT 57.730 170.740 58.050 170.800 ;
        RECT 53.635 170.600 58.050 170.740 ;
        RECT 40.710 170.400 41.030 170.460 ;
        RECT 50.370 170.400 50.690 170.460 ;
        RECT 53.635 170.400 53.775 170.600 ;
        RECT 57.730 170.540 58.050 170.600 ;
        RECT 58.205 170.740 58.495 170.785 ;
        RECT 62.790 170.740 63.110 170.800 ;
        RECT 58.205 170.600 63.110 170.740 ;
        RECT 58.205 170.555 58.495 170.600 ;
        RECT 62.790 170.540 63.110 170.600 ;
        RECT 63.340 170.600 64.860 170.740 ;
        RECT 54.510 170.400 54.830 170.460 ;
        RECT 56.365 170.400 56.655 170.445 ;
        RECT 40.710 170.260 41.400 170.400 ;
        RECT 40.710 170.200 41.030 170.260 ;
        RECT 38.410 170.060 38.730 170.120 ;
        RECT 41.260 170.105 41.400 170.260 ;
        RECT 50.370 170.260 53.775 170.400 ;
        RECT 54.140 170.260 56.655 170.400 ;
        RECT 50.370 170.200 50.690 170.260 ;
        RECT 37.580 169.920 40.940 170.060 ;
        RECT 24.150 169.520 24.470 169.780 ;
        RECT 25.045 169.720 25.335 169.765 ;
        RECT 26.235 169.720 26.525 169.765 ;
        RECT 28.755 169.720 29.045 169.765 ;
        RECT 25.045 169.580 29.045 169.720 ;
        RECT 25.045 169.535 25.335 169.580 ;
        RECT 26.235 169.535 26.525 169.580 ;
        RECT 28.755 169.535 29.045 169.580 ;
        RECT 24.650 169.380 24.940 169.425 ;
        RECT 26.750 169.380 27.040 169.425 ;
        RECT 28.320 169.380 28.610 169.425 ;
        RECT 36.200 169.380 36.340 169.875 ;
        RECT 36.570 169.720 36.890 169.780 ;
        RECT 37.120 169.720 37.260 169.875 ;
        RECT 38.410 169.860 38.730 169.920 ;
        RECT 36.570 169.580 37.260 169.720 ;
        RECT 37.950 169.720 38.270 169.780 ;
        RECT 40.800 169.765 40.940 169.920 ;
        RECT 41.185 169.875 41.475 170.105 ;
        RECT 41.630 170.060 41.950 170.120 ;
        RECT 42.565 170.060 42.855 170.105 ;
        RECT 41.630 169.920 42.855 170.060 ;
        RECT 41.630 169.860 41.950 169.920 ;
        RECT 42.565 169.875 42.855 169.920 ;
        RECT 43.025 169.875 43.315 170.105 ;
        RECT 40.265 169.720 40.555 169.765 ;
        RECT 37.950 169.580 40.555 169.720 ;
        RECT 36.570 169.520 36.890 169.580 ;
        RECT 37.950 169.520 38.270 169.580 ;
        RECT 40.265 169.535 40.555 169.580 ;
        RECT 40.725 169.535 41.015 169.765 ;
        RECT 37.490 169.380 37.810 169.440 ;
        RECT 24.650 169.240 28.610 169.380 ;
        RECT 24.650 169.195 24.940 169.240 ;
        RECT 26.750 169.195 27.040 169.240 ;
        RECT 28.320 169.195 28.610 169.240 ;
        RECT 33.900 169.240 37.810 169.380 ;
        RECT 40.340 169.380 40.480 169.535 ;
        RECT 42.090 169.520 42.410 169.780 ;
        RECT 43.100 169.380 43.240 169.875 ;
        RECT 43.930 169.860 44.250 170.120 ;
        RECT 49.450 169.860 49.770 170.120 ;
        RECT 50.830 169.860 51.150 170.120 ;
        RECT 53.220 170.105 53.360 170.260 ;
        RECT 53.145 169.875 53.435 170.105 ;
        RECT 53.590 169.860 53.910 170.120 ;
        RECT 54.140 170.105 54.280 170.260 ;
        RECT 54.510 170.200 54.830 170.260 ;
        RECT 56.365 170.215 56.655 170.260 ;
        RECT 56.825 170.400 57.115 170.445 ;
        RECT 61.410 170.400 61.730 170.460 ;
        RECT 63.340 170.400 63.480 170.600 ;
        RECT 56.825 170.260 63.480 170.400 ;
        RECT 63.710 170.400 64.030 170.460 ;
        RECT 64.230 170.400 64.520 170.445 ;
        RECT 63.710 170.260 64.520 170.400 ;
        RECT 64.720 170.400 64.860 170.600 ;
        RECT 69.690 170.540 70.010 170.800 ;
        RECT 83.490 170.740 83.810 170.800 ;
        RECT 77.140 170.600 83.810 170.740 ;
        RECT 77.140 170.400 77.280 170.600 ;
        RECT 83.490 170.540 83.810 170.600 ;
        RECT 83.965 170.740 84.255 170.785 ;
        RECT 88.550 170.740 88.870 170.800 ;
        RECT 93.625 170.740 93.915 170.785 ;
        RECT 83.965 170.600 93.915 170.740 ;
        RECT 83.965 170.555 84.255 170.600 ;
        RECT 88.550 170.540 88.870 170.600 ;
        RECT 93.625 170.555 93.915 170.600 ;
        RECT 94.990 170.740 95.310 170.800 ;
        RECT 103.270 170.740 103.590 170.800 ;
        RECT 94.990 170.600 103.590 170.740 ;
        RECT 94.990 170.540 95.310 170.600 ;
        RECT 103.270 170.540 103.590 170.600 ;
        RECT 104.190 170.740 104.510 170.800 ;
        RECT 105.125 170.740 105.415 170.785 ;
        RECT 104.190 170.600 105.415 170.740 ;
        RECT 104.190 170.540 104.510 170.600 ;
        RECT 105.125 170.555 105.415 170.600 ;
        RECT 107.425 170.740 107.715 170.785 ;
        RECT 107.870 170.740 108.190 170.800 ;
        RECT 107.425 170.600 108.190 170.740 ;
        RECT 107.425 170.555 107.715 170.600 ;
        RECT 107.870 170.540 108.190 170.600 ;
        RECT 111.550 170.740 111.870 170.800 ;
        RECT 112.025 170.740 112.315 170.785 ;
        RECT 111.550 170.600 112.315 170.740 ;
        RECT 111.550 170.540 111.870 170.600 ;
        RECT 112.025 170.555 112.315 170.600 ;
        RECT 114.310 170.540 114.630 170.800 ;
        RECT 118.005 170.555 118.295 170.785 ;
        RECT 124.890 170.740 125.210 170.800 ;
        RECT 126.285 170.740 126.575 170.785 ;
        RECT 124.890 170.600 126.575 170.740 ;
        RECT 64.720 170.260 77.280 170.400 ;
        RECT 56.825 170.215 57.115 170.260 ;
        RECT 61.410 170.200 61.730 170.260 ;
        RECT 63.710 170.200 64.030 170.260 ;
        RECT 64.230 170.215 64.520 170.260 ;
        RECT 78.890 170.200 79.210 170.460 ;
        RECT 80.745 170.400 81.035 170.445 ;
        RECT 82.570 170.400 82.890 170.460 ;
        RECT 80.745 170.260 82.890 170.400 ;
        RECT 80.745 170.215 81.035 170.260 ;
        RECT 82.570 170.200 82.890 170.260 ;
        RECT 88.060 170.400 88.350 170.445 ;
        RECT 90.850 170.400 91.170 170.460 ;
        RECT 88.060 170.260 91.170 170.400 ;
        RECT 88.060 170.215 88.350 170.260 ;
        RECT 90.850 170.200 91.170 170.260 ;
        RECT 92.690 170.400 93.010 170.460 ;
        RECT 95.080 170.400 95.220 170.540 ;
        RECT 102.810 170.400 103.130 170.460 ;
        RECT 92.690 170.260 95.220 170.400 ;
        RECT 98.300 170.260 103.130 170.400 ;
        RECT 92.690 170.200 93.010 170.260 ;
        RECT 54.065 169.875 54.355 170.105 ;
        RECT 51.290 169.720 51.610 169.780 ;
        RECT 54.140 169.720 54.280 169.875 ;
        RECT 54.970 169.860 55.290 170.120 ;
        RECT 55.430 169.860 55.750 170.120 ;
        RECT 57.285 170.060 57.575 170.105 ;
        RECT 57.730 170.060 58.050 170.120 ;
        RECT 65.565 170.060 65.855 170.105 ;
        RECT 67.390 170.060 67.710 170.120 ;
        RECT 57.285 169.920 58.050 170.060 ;
        RECT 57.285 169.875 57.575 169.920 ;
        RECT 57.730 169.860 58.050 169.920 ;
        RECT 58.280 169.920 65.320 170.060 ;
        RECT 51.290 169.580 54.280 169.720 ;
        RECT 51.290 169.520 51.610 169.580 ;
        RECT 40.340 169.240 43.240 169.380 ;
        RECT 53.130 169.380 53.450 169.440 ;
        RECT 58.280 169.380 58.420 169.920 ;
        RECT 60.975 169.720 61.265 169.765 ;
        RECT 63.495 169.720 63.785 169.765 ;
        RECT 64.685 169.720 64.975 169.765 ;
        RECT 60.975 169.580 64.975 169.720 ;
        RECT 65.180 169.720 65.320 169.920 ;
        RECT 65.565 169.920 67.710 170.060 ;
        RECT 65.565 169.875 65.855 169.920 ;
        RECT 67.390 169.860 67.710 169.920 ;
        RECT 70.610 169.860 70.930 170.120 ;
        RECT 71.530 169.860 71.850 170.120 ;
        RECT 72.005 169.875 72.295 170.105 ;
        RECT 79.350 170.060 79.670 170.120 ;
        RECT 79.825 170.060 80.115 170.105 ;
        RECT 79.350 169.920 80.115 170.060 ;
        RECT 68.310 169.720 68.630 169.780 ;
        RECT 70.150 169.720 70.470 169.780 ;
        RECT 72.080 169.720 72.220 169.875 ;
        RECT 79.350 169.860 79.670 169.920 ;
        RECT 79.825 169.875 80.115 169.920 ;
        RECT 80.270 170.060 80.590 170.120 ;
        RECT 81.205 170.060 81.495 170.105 ;
        RECT 80.270 169.920 81.495 170.060 ;
        RECT 80.270 169.860 80.590 169.920 ;
        RECT 81.205 169.875 81.495 169.920 ;
        RECT 81.650 170.060 81.970 170.120 ;
        RECT 81.650 169.860 82.110 170.060 ;
        RECT 84.410 169.860 84.730 170.120 ;
        RECT 91.770 170.060 92.090 170.120 ;
        RECT 98.300 170.105 98.440 170.260 ;
        RECT 102.810 170.200 103.130 170.260 ;
        RECT 106.965 170.400 107.255 170.445 ;
        RECT 108.330 170.400 108.650 170.460 ;
        RECT 106.965 170.260 108.650 170.400 ;
        RECT 118.080 170.400 118.220 170.555 ;
        RECT 124.890 170.540 125.210 170.600 ;
        RECT 126.285 170.555 126.575 170.600 ;
        RECT 129.490 170.540 129.810 170.800 ;
        RECT 136.390 170.740 136.710 170.800 ;
        RECT 130.270 170.600 136.710 170.740 ;
        RECT 119.690 170.400 119.980 170.445 ;
        RECT 130.270 170.400 130.410 170.600 ;
        RECT 118.080 170.260 119.980 170.400 ;
        RECT 106.965 170.215 107.255 170.260 ;
        RECT 85.420 169.920 92.090 170.060 ;
        RECT 77.050 169.720 77.370 169.780 ;
        RECT 65.180 169.580 68.080 169.720 ;
        RECT 60.975 169.535 61.265 169.580 ;
        RECT 63.495 169.535 63.785 169.580 ;
        RECT 64.685 169.535 64.975 169.580 ;
        RECT 53.130 169.240 58.420 169.380 ;
        RECT 58.665 169.380 58.955 169.425 ;
        RECT 59.110 169.380 59.430 169.440 ;
        RECT 58.665 169.240 59.430 169.380 ;
        RECT 33.900 169.085 34.040 169.240 ;
        RECT 37.490 169.180 37.810 169.240 ;
        RECT 53.130 169.180 53.450 169.240 ;
        RECT 58.665 169.195 58.955 169.240 ;
        RECT 59.110 169.180 59.430 169.240 ;
        RECT 61.410 169.380 61.700 169.425 ;
        RECT 62.980 169.380 63.270 169.425 ;
        RECT 65.080 169.380 65.370 169.425 ;
        RECT 61.410 169.240 65.370 169.380 ;
        RECT 67.940 169.380 68.080 169.580 ;
        RECT 68.310 169.580 72.220 169.720 ;
        RECT 76.265 169.580 77.370 169.720 ;
        RECT 68.310 169.520 68.630 169.580 ;
        RECT 70.150 169.520 70.470 169.580 ;
        RECT 76.265 169.380 76.405 169.580 ;
        RECT 77.050 169.520 77.370 169.580 ;
        RECT 77.510 169.720 77.830 169.780 ;
        RECT 81.970 169.720 82.110 169.860 ;
        RECT 83.505 169.720 83.795 169.765 ;
        RECT 85.420 169.720 85.560 169.920 ;
        RECT 91.770 169.860 92.090 169.920 ;
        RECT 97.305 169.875 97.595 170.105 ;
        RECT 98.225 169.875 98.515 170.105 ;
        RECT 77.510 169.580 85.560 169.720 ;
        RECT 77.510 169.520 77.830 169.580 ;
        RECT 83.505 169.535 83.795 169.580 ;
        RECT 86.725 169.535 87.015 169.765 ;
        RECT 87.605 169.720 87.895 169.765 ;
        RECT 88.795 169.720 89.085 169.765 ;
        RECT 91.315 169.720 91.605 169.765 ;
        RECT 87.605 169.580 91.605 169.720 ;
        RECT 87.605 169.535 87.895 169.580 ;
        RECT 88.795 169.535 89.085 169.580 ;
        RECT 91.315 169.535 91.605 169.580 ;
        RECT 67.940 169.240 76.405 169.380 ;
        RECT 76.590 169.380 76.910 169.440 ;
        RECT 81.650 169.380 81.970 169.440 ;
        RECT 86.800 169.380 86.940 169.535 ;
        RECT 76.590 169.240 86.940 169.380 ;
        RECT 87.210 169.380 87.500 169.425 ;
        RECT 89.310 169.380 89.600 169.425 ;
        RECT 90.880 169.380 91.170 169.425 ;
        RECT 87.210 169.240 91.170 169.380 ;
        RECT 97.380 169.380 97.520 169.875 ;
        RECT 98.670 169.860 98.990 170.120 ;
        RECT 101.430 170.060 101.750 170.120 ;
        RECT 102.365 170.060 102.655 170.105 ;
        RECT 107.040 170.060 107.180 170.215 ;
        RECT 108.330 170.200 108.650 170.260 ;
        RECT 119.690 170.215 119.980 170.260 ;
        RECT 129.120 170.260 130.410 170.400 ;
        RECT 101.430 169.920 107.180 170.060 ;
        RECT 110.630 170.060 110.950 170.120 ;
        RECT 113.850 170.060 114.170 170.120 ;
        RECT 110.630 169.920 114.170 170.060 ;
        RECT 101.430 169.860 101.750 169.920 ;
        RECT 102.365 169.875 102.655 169.920 ;
        RECT 110.630 169.860 110.950 169.920 ;
        RECT 113.850 169.860 114.170 169.920 ;
        RECT 117.085 170.060 117.375 170.105 ;
        RECT 117.990 170.060 118.310 170.120 ;
        RECT 129.120 170.105 129.260 170.260 ;
        RECT 130.870 170.200 131.190 170.460 ;
        RECT 127.205 170.060 127.495 170.105 ;
        RECT 117.085 169.920 118.310 170.060 ;
        RECT 117.085 169.875 117.375 169.920 ;
        RECT 117.990 169.860 118.310 169.920 ;
        RECT 125.440 169.920 127.495 170.060 ;
        RECT 99.605 169.720 99.895 169.765 ;
        RECT 102.825 169.720 103.115 169.765 ;
        RECT 99.605 169.580 103.115 169.720 ;
        RECT 99.605 169.535 99.895 169.580 ;
        RECT 102.825 169.535 103.115 169.580 ;
        RECT 103.285 169.535 103.575 169.765 ;
        RECT 108.345 169.720 108.635 169.765 ;
        RECT 115.245 169.720 115.535 169.765 ;
        RECT 116.610 169.720 116.930 169.780 ;
        RECT 108.345 169.580 116.930 169.720 ;
        RECT 108.345 169.535 108.635 169.580 ;
        RECT 115.245 169.535 115.535 169.580 ;
        RECT 100.525 169.380 100.815 169.425 ;
        RECT 97.380 169.240 100.815 169.380 ;
        RECT 61.410 169.195 61.700 169.240 ;
        RECT 62.980 169.195 63.270 169.240 ;
        RECT 65.080 169.195 65.370 169.240 ;
        RECT 76.590 169.180 76.910 169.240 ;
        RECT 81.650 169.180 81.970 169.240 ;
        RECT 87.210 169.195 87.500 169.240 ;
        RECT 89.310 169.195 89.600 169.240 ;
        RECT 90.880 169.195 91.170 169.240 ;
        RECT 100.525 169.195 100.815 169.240 ;
        RECT 101.890 169.380 102.210 169.440 ;
        RECT 103.360 169.380 103.500 169.535 ;
        RECT 116.610 169.520 116.930 169.580 ;
        RECT 118.465 169.535 118.755 169.765 ;
        RECT 119.345 169.720 119.635 169.765 ;
        RECT 120.535 169.720 120.825 169.765 ;
        RECT 123.055 169.720 123.345 169.765 ;
        RECT 119.345 169.580 123.345 169.720 ;
        RECT 119.345 169.535 119.635 169.580 ;
        RECT 120.535 169.535 120.825 169.580 ;
        RECT 123.055 169.535 123.345 169.580 ;
        RECT 118.540 169.380 118.680 169.535 ;
        RECT 101.890 169.240 103.500 169.380 ;
        RECT 114.400 169.240 118.680 169.380 ;
        RECT 118.950 169.380 119.240 169.425 ;
        RECT 121.050 169.380 121.340 169.425 ;
        RECT 122.620 169.380 122.910 169.425 ;
        RECT 118.950 169.240 122.910 169.380 ;
        RECT 101.890 169.180 102.210 169.240 ;
        RECT 114.400 169.100 114.540 169.240 ;
        RECT 118.950 169.195 119.240 169.240 ;
        RECT 121.050 169.195 121.340 169.240 ;
        RECT 122.620 169.195 122.910 169.240 ;
        RECT 124.430 169.380 124.750 169.440 ;
        RECT 125.440 169.425 125.580 169.920 ;
        RECT 127.205 169.875 127.495 169.920 ;
        RECT 127.665 169.875 127.955 170.105 ;
        RECT 129.045 169.875 129.335 170.105 ;
        RECT 127.740 169.720 127.880 169.875 ;
        RECT 130.410 169.860 130.730 170.120 ;
        RECT 131.330 169.860 131.650 170.120 ;
        RECT 132.340 170.105 132.480 170.600 ;
        RECT 136.390 170.540 136.710 170.600 ;
        RECT 143.290 170.540 143.610 170.800 ;
        RECT 152.045 170.740 152.335 170.785 ;
        RECT 153.410 170.740 153.730 170.800 ;
        RECT 152.045 170.600 153.730 170.740 ;
        RECT 152.045 170.555 152.335 170.600 ;
        RECT 153.410 170.540 153.730 170.600 ;
        RECT 141.465 170.215 141.755 170.445 ;
        RECT 142.545 170.400 142.835 170.445 ;
        RECT 145.590 170.400 145.910 170.460 ;
        RECT 142.545 170.260 145.910 170.400 ;
        RECT 142.545 170.215 142.835 170.260 ;
        RECT 132.265 169.875 132.555 170.105 ;
        RECT 139.150 169.860 139.470 170.120 ;
        RECT 141.540 170.060 141.680 170.215 ;
        RECT 145.590 170.200 145.910 170.260 ;
        RECT 147.890 170.060 148.210 170.120 ;
        RECT 141.540 169.920 148.210 170.060 ;
        RECT 147.890 169.860 148.210 169.920 ;
        RECT 128.110 169.720 128.430 169.780 ;
        RECT 138.705 169.720 138.995 169.765 ;
        RECT 127.740 169.580 138.995 169.720 ;
        RECT 128.110 169.520 128.430 169.580 ;
        RECT 138.705 169.535 138.995 169.580 ;
        RECT 142.830 169.720 143.150 169.780 ;
        RECT 145.130 169.720 145.450 169.780 ;
        RECT 142.830 169.580 145.450 169.720 ;
        RECT 142.830 169.520 143.150 169.580 ;
        RECT 145.130 169.520 145.450 169.580 ;
        RECT 154.330 169.720 154.650 169.780 ;
        RECT 154.805 169.720 155.095 169.765 ;
        RECT 154.330 169.580 155.095 169.720 ;
        RECT 154.330 169.520 154.650 169.580 ;
        RECT 154.805 169.535 155.095 169.580 ;
        RECT 125.365 169.380 125.655 169.425 ;
        RECT 124.430 169.240 125.655 169.380 ;
        RECT 124.430 169.180 124.750 169.240 ;
        RECT 125.365 169.195 125.655 169.240 ;
        RECT 33.825 168.855 34.115 169.085 ;
        RECT 42.550 169.040 42.870 169.100 ;
        RECT 43.485 169.040 43.775 169.085 ;
        RECT 42.550 168.900 43.775 169.040 ;
        RECT 42.550 168.840 42.870 168.900 ;
        RECT 43.485 168.855 43.775 168.900 ;
        RECT 65.550 169.040 65.870 169.100 ;
        RECT 78.430 169.040 78.750 169.100 ;
        RECT 65.550 168.900 78.750 169.040 ;
        RECT 65.550 168.840 65.870 168.900 ;
        RECT 78.430 168.840 78.750 168.900 ;
        RECT 78.890 169.040 79.210 169.100 ;
        RECT 84.870 169.040 85.190 169.100 ;
        RECT 78.890 168.900 85.190 169.040 ;
        RECT 78.890 168.840 79.210 168.900 ;
        RECT 84.870 168.840 85.190 168.900 ;
        RECT 85.790 169.040 86.110 169.100 ;
        RECT 86.265 169.040 86.555 169.085 ;
        RECT 85.790 168.900 86.555 169.040 ;
        RECT 85.790 168.840 86.110 168.900 ;
        RECT 86.265 168.855 86.555 168.900 ;
        RECT 96.385 169.040 96.675 169.085 ;
        RECT 97.290 169.040 97.610 169.100 ;
        RECT 96.385 168.900 97.610 169.040 ;
        RECT 96.385 168.855 96.675 168.900 ;
        RECT 97.290 168.840 97.610 168.900 ;
        RECT 114.310 168.840 114.630 169.100 ;
        RECT 121.670 169.040 121.990 169.100 ;
        RECT 128.585 169.040 128.875 169.085 ;
        RECT 131.330 169.040 131.650 169.100 ;
        RECT 121.670 168.900 131.650 169.040 ;
        RECT 121.670 168.840 121.990 168.900 ;
        RECT 128.585 168.855 128.875 168.900 ;
        RECT 131.330 168.840 131.650 168.900 ;
        RECT 142.370 168.840 142.690 169.100 ;
        RECT 22.700 168.220 157.020 168.700 ;
        RECT 31.510 168.020 31.830 168.080 ;
        RECT 31.985 168.020 32.275 168.065 ;
        RECT 31.510 167.880 32.275 168.020 ;
        RECT 31.510 167.820 31.830 167.880 ;
        RECT 31.985 167.835 32.275 167.880 ;
        RECT 36.570 168.020 36.890 168.080 ;
        RECT 37.505 168.020 37.795 168.065 ;
        RECT 36.570 167.880 37.795 168.020 ;
        RECT 36.570 167.820 36.890 167.880 ;
        RECT 37.505 167.835 37.795 167.880 ;
        RECT 37.950 168.020 38.270 168.080 ;
        RECT 38.425 168.020 38.715 168.065 ;
        RECT 37.950 167.880 38.715 168.020 ;
        RECT 37.580 167.680 37.720 167.835 ;
        RECT 37.950 167.820 38.270 167.880 ;
        RECT 38.425 167.835 38.715 167.880 ;
        RECT 46.230 167.820 46.550 168.080 ;
        RECT 55.905 168.020 56.195 168.065 ;
        RECT 65.550 168.020 65.870 168.080 ;
        RECT 55.905 167.880 65.870 168.020 ;
        RECT 55.905 167.835 56.195 167.880 ;
        RECT 65.550 167.820 65.870 167.880 ;
        RECT 68.770 168.020 69.090 168.080 ;
        RECT 69.245 168.020 69.535 168.065 ;
        RECT 68.770 167.880 69.535 168.020 ;
        RECT 68.770 167.820 69.090 167.880 ;
        RECT 69.245 167.835 69.535 167.880 ;
        RECT 79.825 167.835 80.115 168.065 ;
        RECT 86.725 168.020 87.015 168.065 ;
        RECT 91.310 168.020 91.630 168.080 ;
        RECT 86.725 167.880 91.630 168.020 ;
        RECT 86.725 167.835 87.015 167.880 ;
        RECT 43.010 167.680 43.330 167.740 ;
        RECT 45.325 167.680 45.615 167.725 ;
        RECT 37.580 167.540 38.180 167.680 ;
        RECT 38.040 167.340 38.180 167.540 ;
        RECT 43.010 167.540 45.615 167.680 ;
        RECT 43.010 167.480 43.330 167.540 ;
        RECT 45.325 167.495 45.615 167.540 ;
        RECT 48.110 167.680 48.400 167.725 ;
        RECT 50.210 167.680 50.500 167.725 ;
        RECT 51.780 167.680 52.070 167.725 ;
        RECT 48.110 167.540 52.070 167.680 ;
        RECT 48.110 167.495 48.400 167.540 ;
        RECT 50.210 167.495 50.500 167.540 ;
        RECT 51.780 167.495 52.070 167.540 ;
        RECT 55.430 167.680 55.750 167.740 ;
        RECT 57.285 167.680 57.575 167.725 ;
        RECT 55.430 167.540 57.575 167.680 ;
        RECT 55.430 167.480 55.750 167.540 ;
        RECT 57.285 167.495 57.575 167.540 ;
        RECT 62.830 167.680 63.120 167.725 ;
        RECT 64.930 167.680 65.220 167.725 ;
        RECT 66.500 167.680 66.790 167.725 ;
        RECT 62.830 167.540 66.790 167.680 ;
        RECT 62.830 167.495 63.120 167.540 ;
        RECT 64.930 167.495 65.220 167.540 ;
        RECT 66.500 167.495 66.790 167.540 ;
        RECT 45.770 167.340 46.090 167.400 ;
        RECT 38.040 167.200 46.090 167.340 ;
        RECT 45.770 167.140 46.090 167.200 ;
        RECT 46.690 167.140 47.010 167.400 ;
        RECT 48.505 167.340 48.795 167.385 ;
        RECT 49.695 167.340 49.985 167.385 ;
        RECT 52.215 167.340 52.505 167.385 ;
        RECT 48.505 167.200 52.505 167.340 ;
        RECT 48.505 167.155 48.795 167.200 ;
        RECT 49.695 167.155 49.985 167.200 ;
        RECT 52.215 167.155 52.505 167.200 ;
        RECT 57.730 167.340 58.050 167.400 ;
        RECT 63.225 167.340 63.515 167.385 ;
        RECT 64.415 167.340 64.705 167.385 ;
        RECT 66.935 167.340 67.225 167.385 ;
        RECT 57.730 167.200 60.640 167.340 ;
        RECT 57.730 167.140 58.050 167.200 ;
        RECT 32.890 166.800 33.210 167.060 ;
        RECT 33.365 167.000 33.655 167.045 ;
        RECT 34.270 167.000 34.590 167.060 ;
        RECT 36.125 167.000 36.415 167.045 ;
        RECT 33.365 166.860 36.415 167.000 ;
        RECT 33.365 166.815 33.655 166.860 ;
        RECT 34.270 166.800 34.590 166.860 ;
        RECT 36.125 166.815 36.415 166.860 ;
        RECT 42.550 166.800 42.870 167.060 ;
        RECT 43.945 167.000 44.235 167.045 ;
        RECT 44.850 167.000 45.170 167.060 ;
        RECT 46.230 167.000 46.550 167.060 ;
        RECT 43.945 166.860 46.550 167.000 ;
        RECT 43.945 166.815 44.235 166.860 ;
        RECT 44.850 166.800 45.170 166.860 ;
        RECT 46.230 166.800 46.550 166.860 ;
        RECT 47.165 166.815 47.455 167.045 ;
        RECT 47.625 167.000 47.915 167.045 ;
        RECT 48.070 167.000 48.390 167.060 ;
        RECT 51.750 167.000 52.070 167.060 ;
        RECT 47.625 166.860 48.390 167.000 ;
        RECT 47.625 166.815 47.915 166.860 ;
        RECT 34.745 166.660 35.035 166.705 ;
        RECT 35.650 166.660 35.970 166.720 ;
        RECT 34.745 166.520 35.970 166.660 ;
        RECT 47.240 166.660 47.380 166.815 ;
        RECT 48.070 166.800 48.390 166.860 ;
        RECT 48.620 166.860 52.070 167.000 ;
        RECT 48.620 166.660 48.760 166.860 ;
        RECT 51.750 166.800 52.070 166.860 ;
        RECT 57.270 167.000 57.590 167.060 ;
        RECT 60.045 167.000 60.335 167.045 ;
        RECT 57.270 166.860 60.335 167.000 ;
        RECT 57.270 166.800 57.590 166.860 ;
        RECT 60.045 166.815 60.335 166.860 ;
        RECT 47.240 166.520 48.760 166.660 ;
        RECT 48.960 166.660 49.250 166.705 ;
        RECT 49.450 166.660 49.770 166.720 ;
        RECT 48.960 166.520 49.770 166.660 ;
        RECT 34.745 166.475 35.035 166.520 ;
        RECT 35.650 166.460 35.970 166.520 ;
        RECT 48.960 166.475 49.250 166.520 ;
        RECT 49.450 166.460 49.770 166.520 ;
        RECT 56.825 166.660 57.115 166.705 ;
        RECT 57.730 166.660 58.050 166.720 ;
        RECT 56.825 166.520 58.050 166.660 ;
        RECT 60.500 166.660 60.640 167.200 ;
        RECT 63.225 167.200 67.225 167.340 ;
        RECT 69.320 167.340 69.460 167.835 ;
        RECT 79.900 167.680 80.040 167.835 ;
        RECT 91.310 167.820 91.630 167.880 ;
        RECT 102.810 167.820 103.130 168.080 ;
        RECT 117.990 167.820 118.310 168.080 ;
        RECT 154.330 167.820 154.650 168.080 ;
        RECT 76.680 167.540 80.040 167.680 ;
        RECT 84.870 167.680 85.190 167.740 ;
        RECT 89.025 167.680 89.315 167.725 ;
        RECT 84.870 167.540 89.315 167.680 ;
        RECT 76.680 167.400 76.820 167.540 ;
        RECT 84.870 167.480 85.190 167.540 ;
        RECT 89.025 167.495 89.315 167.540 ;
        RECT 91.785 167.680 92.075 167.725 ;
        RECT 92.230 167.680 92.550 167.740 ;
        RECT 91.785 167.540 92.550 167.680 ;
        RECT 91.785 167.495 92.075 167.540 ;
        RECT 92.230 167.480 92.550 167.540 ;
        RECT 96.410 167.680 96.700 167.725 ;
        RECT 98.510 167.680 98.800 167.725 ;
        RECT 100.080 167.680 100.370 167.725 ;
        RECT 96.410 167.540 100.370 167.680 ;
        RECT 96.410 167.495 96.700 167.540 ;
        RECT 98.510 167.495 98.800 167.540 ;
        RECT 100.080 167.495 100.370 167.540 ;
        RECT 101.890 167.680 102.210 167.740 ;
        RECT 103.285 167.680 103.575 167.725 ;
        RECT 101.890 167.540 103.575 167.680 ;
        RECT 101.890 167.480 102.210 167.540 ;
        RECT 103.285 167.495 103.575 167.540 ;
        RECT 107.425 167.680 107.715 167.725 ;
        RECT 147.930 167.680 148.220 167.725 ;
        RECT 150.030 167.680 150.320 167.725 ;
        RECT 151.600 167.680 151.890 167.725 ;
        RECT 107.425 167.540 116.840 167.680 ;
        RECT 107.425 167.495 107.715 167.540 ;
        RECT 116.700 167.400 116.840 167.540 ;
        RECT 147.930 167.540 151.890 167.680 ;
        RECT 147.930 167.495 148.220 167.540 ;
        RECT 150.030 167.495 150.320 167.540 ;
        RECT 151.600 167.495 151.890 167.540 ;
        RECT 73.385 167.340 73.675 167.385 ;
        RECT 69.320 167.200 73.675 167.340 ;
        RECT 63.225 167.155 63.515 167.200 ;
        RECT 64.415 167.155 64.705 167.200 ;
        RECT 66.935 167.155 67.225 167.200 ;
        RECT 73.385 167.155 73.675 167.200 ;
        RECT 76.590 167.140 76.910 167.400 ;
        RECT 77.510 167.140 77.830 167.400 ;
        RECT 81.190 167.340 81.510 167.400 ;
        RECT 82.585 167.340 82.875 167.385 ;
        RECT 81.190 167.200 82.875 167.340 ;
        RECT 81.190 167.140 81.510 167.200 ;
        RECT 82.585 167.155 82.875 167.200 ;
        RECT 84.410 167.340 84.730 167.400 ;
        RECT 94.530 167.340 94.850 167.400 ;
        RECT 84.410 167.200 94.850 167.340 ;
        RECT 84.410 167.140 84.730 167.200 ;
        RECT 94.530 167.140 94.850 167.200 ;
        RECT 96.805 167.340 97.095 167.385 ;
        RECT 97.995 167.340 98.285 167.385 ;
        RECT 100.515 167.340 100.805 167.385 ;
        RECT 96.805 167.200 100.805 167.340 ;
        RECT 96.805 167.155 97.095 167.200 ;
        RECT 97.995 167.155 98.285 167.200 ;
        RECT 100.515 167.155 100.805 167.200 ;
        RECT 109.710 167.140 110.030 167.400 ;
        RECT 116.610 167.340 116.930 167.400 ;
        RECT 120.290 167.340 120.610 167.400 ;
        RECT 120.765 167.340 121.055 167.385 ;
        RECT 145.130 167.340 145.450 167.400 ;
        RECT 116.610 167.200 121.055 167.340 ;
        RECT 116.610 167.140 116.930 167.200 ;
        RECT 120.290 167.140 120.610 167.200 ;
        RECT 120.765 167.155 121.055 167.200 ;
        RECT 130.270 167.200 145.450 167.340 ;
        RECT 62.345 167.000 62.635 167.045 ;
        RECT 79.350 167.000 79.670 167.060 ;
        RECT 80.745 167.000 81.035 167.045 ;
        RECT 62.345 166.860 64.400 167.000 ;
        RECT 62.345 166.815 62.635 166.860 ;
        RECT 64.260 166.720 64.400 166.860 ;
        RECT 79.350 166.860 81.035 167.000 ;
        RECT 79.350 166.800 79.670 166.860 ;
        RECT 80.745 166.815 81.035 166.860 ;
        RECT 84.870 166.800 85.190 167.060 ;
        RECT 85.790 166.800 86.110 167.060 ;
        RECT 86.250 167.000 86.570 167.060 ;
        RECT 87.645 167.000 87.935 167.045 ;
        RECT 86.250 166.860 87.935 167.000 ;
        RECT 86.250 166.800 86.570 166.860 ;
        RECT 87.645 166.815 87.935 166.860 ;
        RECT 88.565 167.000 88.855 167.045 ;
        RECT 93.610 167.000 93.930 167.060 ;
        RECT 88.565 166.860 93.930 167.000 ;
        RECT 88.565 166.815 88.855 166.860 ;
        RECT 93.610 166.800 93.930 166.860 ;
        RECT 95.925 167.000 96.215 167.045 ;
        RECT 96.370 167.000 96.690 167.060 ;
        RECT 97.290 167.045 97.610 167.060 ;
        RECT 97.260 167.000 97.610 167.045 ;
        RECT 105.585 167.000 105.875 167.045 ;
        RECT 107.885 167.000 108.175 167.045 ;
        RECT 95.925 166.860 96.690 167.000 ;
        RECT 97.095 166.860 97.610 167.000 ;
        RECT 95.925 166.815 96.215 166.860 ;
        RECT 96.370 166.800 96.690 166.860 ;
        RECT 97.260 166.815 97.610 166.860 ;
        RECT 97.290 166.800 97.610 166.815 ;
        RECT 104.280 166.860 108.175 167.000 ;
        RECT 63.710 166.705 64.030 166.720 ;
        RECT 60.500 166.520 62.940 166.660 ;
        RECT 56.825 166.475 57.115 166.520 ;
        RECT 57.730 166.460 58.050 166.520 ;
        RECT 33.350 166.320 33.670 166.380 ;
        RECT 33.825 166.320 34.115 166.365 ;
        RECT 33.350 166.180 34.115 166.320 ;
        RECT 33.350 166.120 33.670 166.180 ;
        RECT 33.825 166.135 34.115 166.180 ;
        RECT 41.170 166.320 41.490 166.380 ;
        RECT 43.025 166.320 43.315 166.365 ;
        RECT 41.170 166.180 43.315 166.320 ;
        RECT 41.170 166.120 41.490 166.180 ;
        RECT 43.025 166.135 43.315 166.180 ;
        RECT 44.865 166.320 45.155 166.365 ;
        RECT 48.530 166.320 48.850 166.380 ;
        RECT 44.865 166.180 48.850 166.320 ;
        RECT 44.865 166.135 45.155 166.180 ;
        RECT 48.530 166.120 48.850 166.180 ;
        RECT 54.510 166.120 54.830 166.380 ;
        RECT 54.970 166.120 55.290 166.380 ;
        RECT 55.825 166.320 56.115 166.365 ;
        RECT 62.330 166.320 62.650 166.380 ;
        RECT 55.825 166.180 62.650 166.320 ;
        RECT 62.800 166.320 62.940 166.520 ;
        RECT 63.680 166.475 64.030 166.705 ;
        RECT 63.710 166.460 64.030 166.475 ;
        RECT 64.170 166.460 64.490 166.720 ;
        RECT 78.890 166.660 79.210 166.720 ;
        RECT 68.170 166.520 79.210 166.660 ;
        RECT 68.170 166.320 68.310 166.520 ;
        RECT 78.890 166.460 79.210 166.520 ;
        RECT 86.710 166.660 87.030 166.720 ;
        RECT 104.280 166.705 104.420 166.860 ;
        RECT 105.585 166.815 105.875 166.860 ;
        RECT 107.885 166.815 108.175 166.860 ;
        RECT 108.790 166.800 109.110 167.060 ;
        RECT 130.270 167.000 130.410 167.200 ;
        RECT 109.340 166.860 130.410 167.000 ;
        RECT 89.945 166.660 90.235 166.705 ;
        RECT 90.865 166.660 91.155 166.705 ;
        RECT 104.205 166.660 104.495 166.705 ;
        RECT 86.710 166.520 90.235 166.660 ;
        RECT 86.710 166.460 87.030 166.520 ;
        RECT 89.945 166.475 90.235 166.520 ;
        RECT 90.480 166.520 104.495 166.660 ;
        RECT 62.800 166.180 68.310 166.320 ;
        RECT 55.825 166.135 56.115 166.180 ;
        RECT 62.330 166.120 62.650 166.180 ;
        RECT 70.610 166.120 70.930 166.380 ;
        RECT 71.990 166.320 72.310 166.380 ;
        RECT 74.305 166.320 74.595 166.365 ;
        RECT 71.990 166.180 74.595 166.320 ;
        RECT 71.990 166.120 72.310 166.180 ;
        RECT 74.305 166.135 74.595 166.180 ;
        RECT 76.130 166.120 76.450 166.380 ;
        RECT 81.665 166.320 81.955 166.365 ;
        RECT 83.950 166.320 84.270 166.380 ;
        RECT 90.480 166.320 90.620 166.520 ;
        RECT 90.865 166.475 91.155 166.520 ;
        RECT 104.205 166.475 104.495 166.520 ;
        RECT 104.650 166.660 104.970 166.720 ;
        RECT 105.125 166.660 105.415 166.705 ;
        RECT 104.650 166.520 105.415 166.660 ;
        RECT 104.650 166.460 104.970 166.520 ;
        RECT 105.125 166.475 105.415 166.520 ;
        RECT 106.030 166.660 106.350 166.720 ;
        RECT 106.505 166.660 106.795 166.705 ;
        RECT 106.030 166.520 106.795 166.660 ;
        RECT 106.030 166.460 106.350 166.520 ;
        RECT 106.505 166.475 106.795 166.520 ;
        RECT 81.665 166.180 90.620 166.320 ;
        RECT 97.290 166.320 97.610 166.380 ;
        RECT 109.340 166.320 109.480 166.860 ;
        RECT 131.790 166.800 132.110 167.060 ;
        RECT 132.710 166.800 133.030 167.060 ;
        RECT 133.260 167.045 133.400 167.200 ;
        RECT 145.130 167.140 145.450 167.200 ;
        RECT 146.970 167.340 147.290 167.400 ;
        RECT 147.445 167.340 147.735 167.385 ;
        RECT 146.970 167.200 147.735 167.340 ;
        RECT 146.970 167.140 147.290 167.200 ;
        RECT 147.445 167.155 147.735 167.200 ;
        RECT 148.325 167.340 148.615 167.385 ;
        RECT 149.515 167.340 149.805 167.385 ;
        RECT 152.035 167.340 152.325 167.385 ;
        RECT 148.325 167.200 152.325 167.340 ;
        RECT 148.325 167.155 148.615 167.200 ;
        RECT 149.515 167.155 149.805 167.200 ;
        RECT 152.035 167.155 152.325 167.200 ;
        RECT 133.185 166.815 133.475 167.045 ;
        RECT 134.550 166.800 134.870 167.060 ;
        RECT 135.930 166.800 136.250 167.060 ;
        RECT 137.310 167.000 137.630 167.060 ;
        RECT 148.810 167.045 149.130 167.060 ;
        RECT 139.165 167.000 139.455 167.045 ;
        RECT 148.780 167.000 149.130 167.045 ;
        RECT 137.310 166.860 139.455 167.000 ;
        RECT 148.615 166.860 149.130 167.000 ;
        RECT 137.310 166.800 137.630 166.860 ;
        RECT 139.165 166.815 139.455 166.860 ;
        RECT 148.780 166.815 149.130 166.860 ;
        RECT 148.810 166.800 149.130 166.815 ;
        RECT 117.530 166.660 117.850 166.720 ;
        RECT 119.845 166.660 120.135 166.705 ;
        RECT 117.530 166.520 120.135 166.660 ;
        RECT 117.530 166.460 117.850 166.520 ;
        RECT 119.845 166.475 120.135 166.520 ;
        RECT 120.305 166.660 120.595 166.705 ;
        RECT 120.750 166.660 121.070 166.720 ;
        RECT 120.305 166.520 121.070 166.660 ;
        RECT 120.305 166.475 120.595 166.520 ;
        RECT 120.750 166.460 121.070 166.520 ;
        RECT 97.290 166.180 109.480 166.320 ;
        RECT 81.665 166.135 81.955 166.180 ;
        RECT 83.950 166.120 84.270 166.180 ;
        RECT 97.290 166.120 97.610 166.180 ;
        RECT 132.250 166.120 132.570 166.380 ;
        RECT 133.170 166.320 133.490 166.380 ;
        RECT 133.645 166.320 133.935 166.365 ;
        RECT 133.170 166.180 133.935 166.320 ;
        RECT 133.170 166.120 133.490 166.180 ;
        RECT 133.645 166.135 133.935 166.180 ;
        RECT 135.010 166.320 135.330 166.380 ;
        RECT 135.485 166.320 135.775 166.365 ;
        RECT 135.010 166.180 135.775 166.320 ;
        RECT 135.010 166.120 135.330 166.180 ;
        RECT 135.485 166.135 135.775 166.180 ;
        RECT 136.865 166.320 137.155 166.365 ;
        RECT 139.610 166.320 139.930 166.380 ;
        RECT 136.865 166.180 139.930 166.320 ;
        RECT 136.865 166.135 137.155 166.180 ;
        RECT 139.610 166.120 139.930 166.180 ;
        RECT 140.085 166.320 140.375 166.365 ;
        RECT 144.210 166.320 144.530 166.380 ;
        RECT 140.085 166.180 144.530 166.320 ;
        RECT 140.085 166.135 140.375 166.180 ;
        RECT 144.210 166.120 144.530 166.180 ;
        RECT 22.700 165.500 157.820 165.980 ;
        RECT 37.490 165.100 37.810 165.360 ;
        RECT 44.850 165.100 45.170 165.360 ;
        RECT 45.770 165.300 46.090 165.360 ;
        RECT 57.270 165.300 57.590 165.360 ;
        RECT 45.770 165.160 57.590 165.300 ;
        RECT 45.770 165.100 46.090 165.160 ;
        RECT 57.270 165.100 57.590 165.160 ;
        RECT 63.710 165.300 64.030 165.360 ;
        RECT 65.105 165.300 65.395 165.345 ;
        RECT 63.710 165.160 65.395 165.300 ;
        RECT 63.710 165.100 64.030 165.160 ;
        RECT 65.105 165.115 65.395 165.160 ;
        RECT 69.625 165.300 69.915 165.345 ;
        RECT 71.070 165.300 71.390 165.360 ;
        RECT 69.625 165.160 71.390 165.300 ;
        RECT 69.625 165.115 69.915 165.160 ;
        RECT 71.070 165.100 71.390 165.160 ;
        RECT 86.710 165.300 87.030 165.360 ;
        RECT 92.230 165.300 92.550 165.360 ;
        RECT 86.710 165.160 92.550 165.300 ;
        RECT 86.710 165.100 87.030 165.160 ;
        RECT 92.230 165.100 92.550 165.160 ;
        RECT 101.445 165.115 101.735 165.345 ;
        RECT 103.270 165.300 103.590 165.360 ;
        RECT 117.530 165.300 117.850 165.360 ;
        RECT 103.270 165.160 117.850 165.300 ;
        RECT 28.765 164.960 29.055 165.005 ;
        RECT 37.580 164.960 37.720 165.100 ;
        RECT 28.765 164.820 33.120 164.960 ;
        RECT 37.580 164.820 54.280 164.960 ;
        RECT 28.765 164.775 29.055 164.820 ;
        RECT 32.980 164.680 33.120 164.820 ;
        RECT 29.685 164.620 29.975 164.665 ;
        RECT 31.050 164.620 31.370 164.680 ;
        RECT 29.685 164.480 31.370 164.620 ;
        RECT 29.685 164.435 29.975 164.480 ;
        RECT 31.050 164.420 31.370 164.480 ;
        RECT 32.890 164.620 33.210 164.680 ;
        RECT 35.205 164.620 35.495 164.665 ;
        RECT 32.890 164.480 35.495 164.620 ;
        RECT 32.890 164.420 33.210 164.480 ;
        RECT 35.205 164.435 35.495 164.480 ;
        RECT 43.930 164.620 44.250 164.680 ;
        RECT 44.405 164.620 44.695 164.665 ;
        RECT 43.930 164.480 44.695 164.620 ;
        RECT 43.930 164.420 44.250 164.480 ;
        RECT 44.405 164.435 44.695 164.480 ;
        RECT 45.310 164.420 45.630 164.680 ;
        RECT 48.085 164.620 48.375 164.665 ;
        RECT 51.305 164.620 51.595 164.665 ;
        RECT 53.590 164.620 53.910 164.680 ;
        RECT 48.085 164.480 53.910 164.620 ;
        RECT 54.140 164.620 54.280 164.820 ;
        RECT 67.020 164.820 68.080 164.960 ;
        RECT 67.020 164.680 67.160 164.820 ;
        RECT 54.510 164.620 54.830 164.680 ;
        RECT 54.140 164.480 54.830 164.620 ;
        RECT 48.085 164.435 48.375 164.480 ;
        RECT 51.305 164.435 51.595 164.480 ;
        RECT 53.590 164.420 53.910 164.480 ;
        RECT 54.510 164.420 54.830 164.480 ;
        RECT 62.790 164.665 63.110 164.680 ;
        RECT 62.790 164.620 63.140 164.665 ;
        RECT 62.790 164.480 63.305 164.620 ;
        RECT 62.790 164.435 63.140 164.480 ;
        RECT 66.025 164.435 66.315 164.665 ;
        RECT 66.930 164.620 67.250 164.680 ;
        RECT 66.835 164.480 67.250 164.620 ;
        RECT 62.790 164.420 63.110 164.435 ;
        RECT 35.650 164.280 35.970 164.340 ;
        RECT 36.570 164.280 36.890 164.340 ;
        RECT 35.650 164.140 36.890 164.280 ;
        RECT 35.650 164.080 35.970 164.140 ;
        RECT 36.570 164.080 36.890 164.140 ;
        RECT 46.690 164.080 47.010 164.340 ;
        RECT 50.385 164.280 50.675 164.325 ;
        RECT 50.830 164.280 51.150 164.340 ;
        RECT 58.190 164.280 58.510 164.340 ;
        RECT 50.385 164.140 58.510 164.280 ;
        RECT 50.385 164.095 50.675 164.140 ;
        RECT 50.830 164.080 51.150 164.140 ;
        RECT 58.190 164.080 58.510 164.140 ;
        RECT 59.595 164.280 59.885 164.325 ;
        RECT 62.115 164.280 62.405 164.325 ;
        RECT 63.305 164.280 63.595 164.325 ;
        RECT 59.595 164.140 63.595 164.280 ;
        RECT 59.595 164.095 59.885 164.140 ;
        RECT 62.115 164.095 62.405 164.140 ;
        RECT 63.305 164.095 63.595 164.140 ;
        RECT 64.170 164.080 64.490 164.340 ;
        RECT 66.100 164.280 66.240 164.435 ;
        RECT 66.930 164.420 67.250 164.480 ;
        RECT 67.390 164.420 67.710 164.680 ;
        RECT 67.940 164.620 68.080 164.820 ;
        RECT 70.610 164.760 70.930 165.020 ;
        RECT 81.650 164.960 81.970 165.020 ;
        RECT 89.485 164.960 89.775 165.005 ;
        RECT 90.850 164.960 91.170 165.020 ;
        RECT 96.370 164.960 96.690 165.020 ;
        RECT 98.685 164.960 98.975 165.005 ;
        RECT 81.650 164.820 86.940 164.960 ;
        RECT 81.650 164.760 81.970 164.820 ;
        RECT 67.940 164.480 69.460 164.620 ;
        RECT 66.100 164.140 69.000 164.280 ;
        RECT 47.610 163.940 47.930 164.000 ;
        RECT 68.860 163.985 69.000 164.140 ;
        RECT 60.030 163.940 60.320 163.985 ;
        RECT 61.600 163.940 61.890 163.985 ;
        RECT 63.700 163.940 63.990 163.985 ;
        RECT 47.610 163.800 59.800 163.940 ;
        RECT 47.610 163.740 47.930 163.800 ;
        RECT 26.910 163.600 27.230 163.660 ;
        RECT 27.845 163.600 28.135 163.645 ;
        RECT 26.910 163.460 28.135 163.600 ;
        RECT 26.910 163.400 27.230 163.460 ;
        RECT 27.845 163.415 28.135 163.460 ;
        RECT 35.665 163.600 35.955 163.645 ;
        RECT 47.150 163.600 47.470 163.660 ;
        RECT 35.665 163.460 47.470 163.600 ;
        RECT 35.665 163.415 35.955 163.460 ;
        RECT 47.150 163.400 47.470 163.460 ;
        RECT 51.765 163.600 52.055 163.645 ;
        RECT 52.210 163.600 52.530 163.660 ;
        RECT 51.765 163.460 52.530 163.600 ;
        RECT 59.660 163.600 59.800 163.800 ;
        RECT 60.030 163.800 63.990 163.940 ;
        RECT 60.030 163.755 60.320 163.800 ;
        RECT 61.600 163.755 61.890 163.800 ;
        RECT 63.700 163.755 63.990 163.800 ;
        RECT 68.785 163.755 69.075 163.985 ;
        RECT 69.320 163.940 69.460 164.480 ;
        RECT 71.990 164.420 72.310 164.680 ;
        RECT 72.925 164.620 73.215 164.665 ;
        RECT 74.765 164.620 75.055 164.665 ;
        RECT 72.925 164.480 75.055 164.620 ;
        RECT 72.925 164.435 73.215 164.480 ;
        RECT 74.765 164.435 75.055 164.480 ;
        RECT 76.590 164.620 76.910 164.680 ;
        RECT 78.890 164.620 79.210 164.680 ;
        RECT 76.590 164.480 79.210 164.620 ;
        RECT 76.590 164.420 76.910 164.480 ;
        RECT 78.890 164.420 79.210 164.480 ;
        RECT 81.190 164.620 81.510 164.680 ;
        RECT 82.125 164.620 82.415 164.665 ;
        RECT 81.190 164.480 82.415 164.620 ;
        RECT 81.190 164.420 81.510 164.480 ;
        RECT 82.125 164.435 82.415 164.480 ;
        RECT 83.045 164.435 83.335 164.665 ;
        RECT 70.610 164.280 70.930 164.340 ;
        RECT 71.085 164.280 71.375 164.325 ;
        RECT 70.610 164.140 71.375 164.280 ;
        RECT 70.610 164.080 70.930 164.140 ;
        RECT 71.085 164.095 71.375 164.140 ;
        RECT 81.650 164.280 81.970 164.340 ;
        RECT 83.120 164.280 83.260 164.435 ;
        RECT 86.800 164.340 86.940 164.820 ;
        RECT 89.485 164.820 91.170 164.960 ;
        RECT 89.485 164.775 89.775 164.820 ;
        RECT 90.850 164.760 91.170 164.820 ;
        RECT 96.000 164.820 98.975 164.960 ;
        RECT 101.520 164.960 101.660 165.115 ;
        RECT 103.270 165.100 103.590 165.160 ;
        RECT 117.530 165.100 117.850 165.160 ;
        RECT 130.425 165.300 130.715 165.345 ;
        RECT 132.710 165.300 133.030 165.360 ;
        RECT 130.425 165.160 133.030 165.300 ;
        RECT 130.425 165.115 130.715 165.160 ;
        RECT 132.710 165.100 133.030 165.160 ;
        RECT 134.180 165.160 135.700 165.300 ;
        RECT 105.110 164.960 105.430 165.020 ;
        RECT 108.790 164.960 109.110 165.020 ;
        RECT 101.520 164.820 109.110 164.960 ;
        RECT 89.025 164.620 89.315 164.665 ;
        RECT 95.005 164.620 95.295 164.665 ;
        RECT 96.000 164.620 96.140 164.820 ;
        RECT 96.370 164.760 96.690 164.820 ;
        RECT 98.685 164.775 98.975 164.820 ;
        RECT 105.110 164.760 105.430 164.820 ;
        RECT 108.790 164.760 109.110 164.820 ;
        RECT 128.570 164.960 128.890 165.020 ;
        RECT 129.045 164.960 129.335 165.005 ;
        RECT 129.965 164.960 130.255 165.005 ;
        RECT 132.265 164.960 132.555 165.005 ;
        RECT 133.170 164.960 133.490 165.020 ;
        RECT 128.570 164.820 129.720 164.960 ;
        RECT 128.570 164.760 128.890 164.820 ;
        RECT 129.045 164.775 129.335 164.820 ;
        RECT 89.025 164.480 96.140 164.620 ;
        RECT 89.025 164.435 89.315 164.480 ;
        RECT 95.005 164.435 95.295 164.480 ;
        RECT 97.765 164.435 98.055 164.665 ;
        RECT 99.605 164.620 99.895 164.665 ;
        RECT 100.525 164.620 100.815 164.665 ;
        RECT 99.605 164.480 100.815 164.620 ;
        RECT 99.605 164.435 99.895 164.480 ;
        RECT 100.525 164.435 100.815 164.480 ;
        RECT 103.730 164.620 104.050 164.680 ;
        RECT 105.585 164.620 105.875 164.665 ;
        RECT 109.265 164.620 109.555 164.665 ;
        RECT 103.730 164.480 109.555 164.620 ;
        RECT 81.650 164.140 83.260 164.280 ;
        RECT 86.710 164.280 87.030 164.340 ;
        RECT 93.625 164.280 93.915 164.325 ;
        RECT 95.910 164.280 96.230 164.340 ;
        RECT 86.710 164.140 96.230 164.280 ;
        RECT 81.650 164.080 81.970 164.140 ;
        RECT 86.710 164.080 87.030 164.140 ;
        RECT 93.625 164.095 93.915 164.140 ;
        RECT 95.910 164.080 96.230 164.140 ;
        RECT 96.385 164.280 96.675 164.325 ;
        RECT 97.840 164.280 97.980 164.435 ;
        RECT 103.730 164.420 104.050 164.480 ;
        RECT 105.585 164.435 105.875 164.480 ;
        RECT 109.265 164.435 109.555 164.480 ;
        RECT 113.865 164.620 114.155 164.665 ;
        RECT 114.310 164.620 114.630 164.680 ;
        RECT 113.865 164.480 114.630 164.620 ;
        RECT 113.865 164.435 114.155 164.480 ;
        RECT 114.310 164.420 114.630 164.480 ;
        RECT 115.200 164.620 115.490 164.665 ;
        RECT 120.750 164.620 121.070 164.680 ;
        RECT 115.200 164.480 121.070 164.620 ;
        RECT 115.200 164.435 115.490 164.480 ;
        RECT 120.750 164.420 121.070 164.480 ;
        RECT 96.385 164.140 97.980 164.280 ;
        RECT 114.745 164.280 115.035 164.325 ;
        RECT 115.935 164.280 116.225 164.325 ;
        RECT 118.455 164.280 118.745 164.325 ;
        RECT 121.685 164.280 121.975 164.325 ;
        RECT 127.190 164.280 127.510 164.340 ;
        RECT 114.745 164.140 118.745 164.280 ;
        RECT 96.385 164.095 96.675 164.140 ;
        RECT 114.745 164.095 115.035 164.140 ;
        RECT 115.935 164.095 116.225 164.140 ;
        RECT 118.455 164.095 118.745 164.140 ;
        RECT 120.840 164.140 127.510 164.280 ;
        RECT 129.580 164.280 129.720 164.820 ;
        RECT 129.965 164.820 133.490 164.960 ;
        RECT 129.965 164.775 130.255 164.820 ;
        RECT 132.265 164.775 132.555 164.820 ;
        RECT 133.170 164.760 133.490 164.820 ;
        RECT 133.630 164.760 133.950 165.020 ;
        RECT 134.180 165.005 134.320 165.160 ;
        RECT 135.010 165.005 135.330 165.020 ;
        RECT 134.105 164.775 134.395 165.005 ;
        RECT 135.010 164.775 135.395 165.005 ;
        RECT 135.560 164.960 135.700 165.160 ;
        RECT 135.930 165.100 136.250 165.360 ;
        RECT 136.390 164.960 136.710 165.020 ;
        RECT 135.560 164.820 136.710 164.960 ;
        RECT 135.010 164.760 135.330 164.775 ;
        RECT 136.390 164.760 136.710 164.820 ;
        RECT 130.425 164.620 130.715 164.665 ;
        RECT 131.330 164.620 131.650 164.680 ;
        RECT 131.805 164.620 132.095 164.665 ;
        RECT 130.425 164.480 132.095 164.620 ;
        RECT 130.425 164.435 130.715 164.480 ;
        RECT 131.330 164.420 131.650 164.480 ;
        RECT 131.805 164.435 132.095 164.480 ;
        RECT 132.725 164.620 133.015 164.665 ;
        RECT 133.720 164.620 133.860 164.760 ;
        RECT 132.725 164.480 133.860 164.620 ;
        RECT 139.610 164.620 139.930 164.680 ;
        RECT 141.970 164.620 142.260 164.665 ;
        RECT 139.610 164.480 142.260 164.620 ;
        RECT 132.725 164.435 133.015 164.480 ;
        RECT 131.880 164.280 132.020 164.435 ;
        RECT 139.610 164.420 139.930 164.480 ;
        RECT 141.970 164.435 142.260 164.480 ;
        RECT 134.550 164.280 134.870 164.340 ;
        RECT 138.715 164.280 139.005 164.325 ;
        RECT 141.235 164.280 141.525 164.325 ;
        RECT 142.425 164.280 142.715 164.325 ;
        RECT 129.580 164.140 130.640 164.280 ;
        RECT 131.880 164.140 136.620 164.280 ;
        RECT 87.170 163.940 87.490 164.000 ;
        RECT 96.460 163.940 96.600 164.095 ;
        RECT 69.320 163.800 87.490 163.940 ;
        RECT 87.170 163.740 87.490 163.800 ;
        RECT 88.640 163.800 96.600 163.940 ;
        RECT 98.670 163.940 98.990 164.000 ;
        RECT 100.510 163.940 100.830 164.000 ;
        RECT 106.505 163.940 106.795 163.985 ;
        RECT 98.670 163.800 106.795 163.940 ;
        RECT 88.640 163.660 88.780 163.800 ;
        RECT 98.670 163.740 98.990 163.800 ;
        RECT 100.510 163.740 100.830 163.800 ;
        RECT 106.505 163.755 106.795 163.800 ;
        RECT 108.790 163.740 109.110 164.000 ;
        RECT 120.840 163.985 120.980 164.140 ;
        RECT 121.685 164.095 121.975 164.140 ;
        RECT 127.190 164.080 127.510 164.140 ;
        RECT 130.500 164.000 130.640 164.140 ;
        RECT 134.550 164.080 134.870 164.140 ;
        RECT 114.350 163.940 114.640 163.985 ;
        RECT 116.450 163.940 116.740 163.985 ;
        RECT 118.020 163.940 118.310 163.985 ;
        RECT 114.350 163.800 118.310 163.940 ;
        RECT 114.350 163.755 114.640 163.800 ;
        RECT 116.450 163.755 116.740 163.800 ;
        RECT 118.020 163.755 118.310 163.800 ;
        RECT 120.765 163.755 121.055 163.985 ;
        RECT 130.410 163.740 130.730 164.000 ;
        RECT 130.870 163.740 131.190 164.000 ;
        RECT 132.710 163.940 133.030 164.000 ;
        RECT 136.480 163.985 136.620 164.140 ;
        RECT 138.715 164.140 142.715 164.280 ;
        RECT 138.715 164.095 139.005 164.140 ;
        RECT 141.235 164.095 141.525 164.140 ;
        RECT 142.425 164.095 142.715 164.140 ;
        RECT 143.305 164.280 143.595 164.325 ;
        RECT 147.890 164.280 148.210 164.340 ;
        RECT 143.305 164.140 148.210 164.280 ;
        RECT 143.305 164.095 143.595 164.140 ;
        RECT 147.890 164.080 148.210 164.140 ;
        RECT 132.710 163.800 135.240 163.940 ;
        RECT 132.710 163.740 133.030 163.800 ;
        RECT 66.930 163.600 67.250 163.660 ;
        RECT 59.660 163.460 67.250 163.600 ;
        RECT 51.765 163.415 52.055 163.460 ;
        RECT 52.210 163.400 52.530 163.460 ;
        RECT 66.930 163.400 67.250 163.460 ;
        RECT 69.690 163.600 70.010 163.660 ;
        RECT 71.530 163.600 71.850 163.660 ;
        RECT 69.690 163.460 71.850 163.600 ;
        RECT 69.690 163.400 70.010 163.460 ;
        RECT 71.530 163.400 71.850 163.460 ;
        RECT 75.685 163.600 75.975 163.645 ;
        RECT 76.130 163.600 76.450 163.660 ;
        RECT 75.685 163.460 76.450 163.600 ;
        RECT 75.685 163.415 75.975 163.460 ;
        RECT 76.130 163.400 76.450 163.460 ;
        RECT 80.745 163.600 81.035 163.645 ;
        RECT 81.190 163.600 81.510 163.660 ;
        RECT 86.250 163.600 86.570 163.660 ;
        RECT 80.745 163.460 86.570 163.600 ;
        RECT 80.745 163.415 81.035 163.460 ;
        RECT 81.190 163.400 81.510 163.460 ;
        RECT 86.250 163.400 86.570 163.460 ;
        RECT 88.550 163.400 88.870 163.660 ;
        RECT 96.845 163.600 97.135 163.645 ;
        RECT 102.350 163.600 102.670 163.660 ;
        RECT 106.030 163.600 106.350 163.660 ;
        RECT 96.845 163.460 106.350 163.600 ;
        RECT 96.845 163.415 97.135 163.460 ;
        RECT 102.350 163.400 102.670 163.460 ;
        RECT 106.030 163.400 106.350 163.460 ;
        RECT 123.970 163.600 124.290 163.660 ;
        RECT 124.445 163.600 124.735 163.645 ;
        RECT 123.970 163.460 124.735 163.600 ;
        RECT 123.970 163.400 124.290 163.460 ;
        RECT 124.445 163.415 124.735 163.460 ;
        RECT 133.630 163.400 133.950 163.660 ;
        RECT 135.100 163.645 135.240 163.800 ;
        RECT 136.405 163.755 136.695 163.985 ;
        RECT 139.150 163.940 139.440 163.985 ;
        RECT 140.720 163.940 141.010 163.985 ;
        RECT 142.820 163.940 143.110 163.985 ;
        RECT 139.150 163.800 143.110 163.940 ;
        RECT 139.150 163.755 139.440 163.800 ;
        RECT 140.720 163.755 141.010 163.800 ;
        RECT 142.820 163.755 143.110 163.800 ;
        RECT 135.025 163.415 135.315 163.645 ;
        RECT 22.700 162.780 157.020 163.260 ;
        RECT 27.830 162.580 28.150 162.640 ;
        RECT 29.670 162.580 29.990 162.640 ;
        RECT 33.365 162.580 33.655 162.625 ;
        RECT 27.830 162.440 33.655 162.580 ;
        RECT 27.830 162.380 28.150 162.440 ;
        RECT 29.670 162.380 29.990 162.440 ;
        RECT 33.365 162.395 33.655 162.440 ;
        RECT 41.170 162.580 41.490 162.640 ;
        RECT 44.405 162.580 44.695 162.625 ;
        RECT 41.170 162.440 44.695 162.580 ;
        RECT 41.170 162.380 41.490 162.440 ;
        RECT 44.405 162.395 44.695 162.440 ;
        RECT 49.450 162.380 49.770 162.640 ;
        RECT 55.905 162.580 56.195 162.625 ;
        RECT 57.730 162.580 58.050 162.640 ;
        RECT 55.905 162.440 58.050 162.580 ;
        RECT 55.905 162.395 56.195 162.440 ;
        RECT 57.730 162.380 58.050 162.440 ;
        RECT 62.805 162.580 63.095 162.625 ;
        RECT 63.250 162.580 63.570 162.640 ;
        RECT 65.090 162.580 65.410 162.640 ;
        RECT 62.805 162.440 65.410 162.580 ;
        RECT 62.805 162.395 63.095 162.440 ;
        RECT 63.250 162.380 63.570 162.440 ;
        RECT 65.090 162.380 65.410 162.440 ;
        RECT 70.625 162.580 70.915 162.625 ;
        RECT 76.590 162.580 76.910 162.640 ;
        RECT 70.625 162.440 76.910 162.580 ;
        RECT 70.625 162.395 70.915 162.440 ;
        RECT 76.590 162.380 76.910 162.440 ;
        RECT 88.550 162.580 88.870 162.640 ;
        RECT 120.750 162.580 121.070 162.640 ;
        RECT 121.225 162.580 121.515 162.625 ;
        RECT 131.345 162.580 131.635 162.625 ;
        RECT 131.790 162.580 132.110 162.640 ;
        RECT 88.550 162.440 93.380 162.580 ;
        RECT 88.550 162.380 88.870 162.440 ;
        RECT 24.650 162.240 24.940 162.285 ;
        RECT 26.750 162.240 27.040 162.285 ;
        RECT 28.320 162.240 28.610 162.285 ;
        RECT 24.650 162.100 28.610 162.240 ;
        RECT 24.650 162.055 24.940 162.100 ;
        RECT 26.750 162.055 27.040 162.100 ;
        RECT 28.320 162.055 28.610 162.100 ;
        RECT 30.130 162.240 30.450 162.300 ;
        RECT 31.525 162.240 31.815 162.285 ;
        RECT 30.130 162.100 31.815 162.240 ;
        RECT 30.130 162.040 30.450 162.100 ;
        RECT 31.525 162.055 31.815 162.100 ;
        RECT 36.610 162.240 36.900 162.285 ;
        RECT 38.710 162.240 39.000 162.285 ;
        RECT 40.280 162.240 40.570 162.285 ;
        RECT 47.610 162.240 47.930 162.300 ;
        RECT 36.610 162.100 40.570 162.240 ;
        RECT 36.610 162.055 36.900 162.100 ;
        RECT 38.710 162.055 39.000 162.100 ;
        RECT 40.280 162.055 40.570 162.100 ;
        RECT 47.240 162.100 47.930 162.240 ;
        RECT 25.045 161.900 25.335 161.945 ;
        RECT 26.235 161.900 26.525 161.945 ;
        RECT 28.755 161.900 29.045 161.945 ;
        RECT 36.125 161.900 36.415 161.945 ;
        RECT 25.045 161.760 29.045 161.900 ;
        RECT 25.045 161.715 25.335 161.760 ;
        RECT 26.235 161.715 26.525 161.760 ;
        RECT 28.755 161.715 29.045 161.760 ;
        RECT 29.300 161.760 36.415 161.900 ;
        RECT 24.150 161.560 24.470 161.620 ;
        RECT 29.300 161.560 29.440 161.760 ;
        RECT 36.125 161.715 36.415 161.760 ;
        RECT 37.005 161.900 37.295 161.945 ;
        RECT 38.195 161.900 38.485 161.945 ;
        RECT 40.715 161.900 41.005 161.945 ;
        RECT 37.005 161.760 41.005 161.900 ;
        RECT 37.005 161.715 37.295 161.760 ;
        RECT 38.195 161.715 38.485 161.760 ;
        RECT 40.715 161.715 41.005 161.760 ;
        RECT 24.150 161.420 29.440 161.560 ;
        RECT 24.150 161.360 24.470 161.420 ;
        RECT 24.610 161.220 24.930 161.280 ;
        RECT 25.390 161.220 25.680 161.265 ;
        RECT 24.610 161.080 25.680 161.220 ;
        RECT 24.610 161.020 24.930 161.080 ;
        RECT 25.390 161.035 25.680 161.080 ;
        RECT 34.730 161.220 35.050 161.280 ;
        RECT 37.350 161.220 37.640 161.265 ;
        RECT 34.730 161.080 37.640 161.220 ;
        RECT 34.730 161.020 35.050 161.080 ;
        RECT 37.350 161.035 37.640 161.080 ;
        RECT 40.710 161.220 41.030 161.280 ;
        RECT 45.325 161.220 45.615 161.265 ;
        RECT 40.710 161.080 45.615 161.220 ;
        RECT 47.240 161.220 47.380 162.100 ;
        RECT 47.610 162.040 47.930 162.100 ;
        RECT 53.590 162.240 53.910 162.300 ;
        RECT 64.630 162.240 64.950 162.300 ;
        RECT 53.590 162.100 64.950 162.240 ;
        RECT 53.590 162.040 53.910 162.100 ;
        RECT 64.630 162.040 64.950 162.100 ;
        RECT 73.370 162.240 73.660 162.285 ;
        RECT 74.940 162.240 75.230 162.285 ;
        RECT 77.040 162.240 77.330 162.285 ;
        RECT 73.370 162.100 77.330 162.240 ;
        RECT 73.370 162.055 73.660 162.100 ;
        RECT 74.940 162.055 75.230 162.100 ;
        RECT 77.040 162.055 77.330 162.100 ;
        RECT 77.510 162.240 77.830 162.300 ;
        RECT 92.690 162.240 93.010 162.300 ;
        RECT 77.510 162.100 89.240 162.240 ;
        RECT 77.510 162.040 77.830 162.100 ;
        RECT 54.970 161.900 55.290 161.960 ;
        RECT 59.110 161.900 59.430 161.960 ;
        RECT 72.935 161.900 73.225 161.945 ;
        RECT 75.455 161.900 75.745 161.945 ;
        RECT 76.645 161.900 76.935 161.945 ;
        RECT 47.700 161.760 55.290 161.900 ;
        RECT 47.700 161.605 47.840 161.760 ;
        RECT 54.970 161.700 55.290 161.760 ;
        RECT 55.980 161.760 68.310 161.900 ;
        RECT 47.625 161.375 47.915 161.605 ;
        RECT 49.005 161.375 49.295 161.605 ;
        RECT 48.545 161.220 48.835 161.265 ;
        RECT 47.240 161.080 48.835 161.220 ;
        RECT 40.710 161.020 41.030 161.080 ;
        RECT 45.325 161.035 45.615 161.080 ;
        RECT 48.545 161.035 48.835 161.080 ;
        RECT 31.065 160.880 31.355 160.925 ;
        RECT 32.890 160.880 33.210 160.940 ;
        RECT 31.065 160.740 33.210 160.880 ;
        RECT 31.065 160.695 31.355 160.740 ;
        RECT 32.890 160.680 33.210 160.740 ;
        RECT 33.350 160.680 33.670 160.940 ;
        RECT 34.270 160.680 34.590 160.940 ;
        RECT 36.570 160.880 36.890 160.940 ;
        RECT 43.025 160.880 43.315 160.925 ;
        RECT 36.570 160.740 43.315 160.880 ;
        RECT 36.570 160.680 36.890 160.740 ;
        RECT 43.025 160.695 43.315 160.740 ;
        RECT 43.470 160.680 43.790 160.940 ;
        RECT 44.390 160.925 44.710 160.940 ;
        RECT 44.325 160.695 44.710 160.925 ;
        RECT 46.705 160.880 46.995 160.925 ;
        RECT 47.610 160.880 47.930 160.940 ;
        RECT 46.705 160.740 47.930 160.880 ;
        RECT 49.080 160.880 49.220 161.375 ;
        RECT 50.370 161.360 50.690 161.620 ;
        RECT 51.290 161.360 51.610 161.620 ;
        RECT 52.210 161.360 52.530 161.620 ;
        RECT 53.145 161.560 53.435 161.605 ;
        RECT 53.590 161.560 53.910 161.620 ;
        RECT 55.980 161.560 56.120 161.760 ;
        RECT 59.110 161.700 59.430 161.760 ;
        RECT 53.145 161.420 53.910 161.560 ;
        RECT 53.145 161.375 53.435 161.420 ;
        RECT 53.590 161.360 53.910 161.420 ;
        RECT 54.600 161.420 56.120 161.560 ;
        RECT 50.845 161.220 51.135 161.265 ;
        RECT 54.600 161.220 54.740 161.420 ;
        RECT 56.365 161.375 56.655 161.605 ;
        RECT 68.170 161.560 68.310 161.760 ;
        RECT 72.935 161.760 76.935 161.900 ;
        RECT 72.935 161.715 73.225 161.760 ;
        RECT 75.455 161.715 75.745 161.760 ;
        RECT 76.645 161.715 76.935 161.760 ;
        RECT 78.890 161.900 79.210 161.960 ;
        RECT 80.270 161.900 80.590 161.960 ;
        RECT 85.345 161.900 85.635 161.945 ;
        RECT 88.550 161.900 88.870 161.960 ;
        RECT 78.890 161.760 82.110 161.900 ;
        RECT 78.890 161.700 79.210 161.760 ;
        RECT 80.270 161.700 80.590 161.760 ;
        RECT 76.130 161.605 76.450 161.620 ;
        RECT 76.130 161.560 76.480 161.605 ;
        RECT 77.050 161.560 77.370 161.620 ;
        RECT 77.525 161.560 77.815 161.605 ;
        RECT 68.170 161.420 75.900 161.560 ;
        RECT 50.845 161.080 54.740 161.220 ;
        RECT 54.970 161.220 55.290 161.280 ;
        RECT 56.440 161.220 56.580 161.375 ;
        RECT 54.970 161.080 56.580 161.220 ;
        RECT 59.585 161.220 59.875 161.265 ;
        RECT 63.725 161.220 64.015 161.265 ;
        RECT 59.585 161.080 64.015 161.220 ;
        RECT 50.845 161.035 51.135 161.080 ;
        RECT 54.970 161.020 55.290 161.080 ;
        RECT 59.585 161.035 59.875 161.080 ;
        RECT 63.725 161.035 64.015 161.080 ;
        RECT 64.630 161.220 64.950 161.280 ;
        RECT 75.210 161.220 75.530 161.280 ;
        RECT 64.630 161.080 75.530 161.220 ;
        RECT 64.630 161.020 64.950 161.080 ;
        RECT 75.210 161.020 75.530 161.080 ;
        RECT 57.270 160.880 57.590 160.940 ;
        RECT 49.080 160.740 57.590 160.880 ;
        RECT 46.705 160.695 46.995 160.740 ;
        RECT 44.390 160.680 44.710 160.695 ;
        RECT 47.610 160.680 47.930 160.740 ;
        RECT 57.270 160.680 57.590 160.740 ;
        RECT 61.870 160.680 62.190 160.940 ;
        RECT 62.790 160.925 63.110 160.940 ;
        RECT 62.725 160.695 63.110 160.925 ;
        RECT 75.760 160.880 75.900 161.420 ;
        RECT 76.130 161.420 76.645 161.560 ;
        RECT 77.050 161.420 77.815 161.560 ;
        RECT 76.130 161.375 76.480 161.420 ;
        RECT 76.130 161.360 76.450 161.375 ;
        RECT 77.050 161.360 77.370 161.420 ;
        RECT 77.525 161.375 77.815 161.420 ;
        RECT 80.730 161.360 81.050 161.620 ;
        RECT 81.970 161.560 82.110 161.760 ;
        RECT 85.345 161.760 88.870 161.900 ;
        RECT 85.345 161.715 85.635 161.760 ;
        RECT 88.550 161.700 88.870 161.760 ;
        RECT 82.585 161.560 82.875 161.605 ;
        RECT 81.970 161.420 82.875 161.560 ;
        RECT 82.585 161.375 82.875 161.420 ;
        RECT 86.265 161.375 86.555 161.605 ;
        RECT 79.350 161.220 79.670 161.280 ;
        RECT 81.650 161.220 81.970 161.280 ;
        RECT 86.340 161.220 86.480 161.375 ;
        RECT 79.350 161.080 86.480 161.220 ;
        RECT 79.350 161.020 79.670 161.080 ;
        RECT 81.650 161.020 81.970 161.080 ;
        RECT 82.570 160.880 82.890 160.940 ;
        RECT 75.760 160.740 82.890 160.880 ;
        RECT 62.790 160.680 63.110 160.695 ;
        RECT 82.570 160.680 82.890 160.740 ;
        RECT 85.330 160.880 85.650 160.940 ;
        RECT 87.645 160.880 87.935 160.925 ;
        RECT 85.330 160.740 87.935 160.880 ;
        RECT 89.100 160.880 89.240 162.100 ;
        RECT 89.560 162.100 93.010 162.240 ;
        RECT 89.560 161.605 89.700 162.100 ;
        RECT 92.690 162.040 93.010 162.100 ;
        RECT 90.865 161.900 91.155 161.945 ;
        RECT 91.770 161.900 92.090 161.960 ;
        RECT 90.865 161.760 92.090 161.900 ;
        RECT 90.865 161.715 91.155 161.760 ;
        RECT 91.770 161.700 92.090 161.760 ;
        RECT 89.485 161.375 89.775 161.605 ;
        RECT 89.945 161.560 90.235 161.605 ;
        RECT 92.705 161.560 92.995 161.605 ;
        RECT 89.945 161.420 92.995 161.560 ;
        RECT 93.240 161.560 93.380 162.440 ;
        RECT 120.750 162.440 121.515 162.580 ;
        RECT 120.750 162.380 121.070 162.440 ;
        RECT 121.225 162.395 121.515 162.440 ;
        RECT 130.270 162.440 132.110 162.580 ;
        RECT 93.610 162.240 93.930 162.300 ;
        RECT 104.190 162.240 104.510 162.300 ;
        RECT 93.610 162.100 104.510 162.240 ;
        RECT 93.610 162.040 93.930 162.100 ;
        RECT 104.190 162.040 104.510 162.100 ;
        RECT 106.070 162.240 106.360 162.285 ;
        RECT 108.170 162.240 108.460 162.285 ;
        RECT 109.740 162.240 110.030 162.285 ;
        RECT 106.070 162.100 110.030 162.240 ;
        RECT 106.070 162.055 106.360 162.100 ;
        RECT 108.170 162.055 108.460 162.100 ;
        RECT 109.740 162.055 110.030 162.100 ;
        RECT 112.485 162.240 112.775 162.285 ;
        RECT 129.490 162.240 129.810 162.300 ;
        RECT 130.270 162.240 130.410 162.440 ;
        RECT 131.345 162.395 131.635 162.440 ;
        RECT 131.790 162.380 132.110 162.440 ;
        RECT 132.250 162.580 132.570 162.640 ;
        RECT 135.485 162.580 135.775 162.625 ;
        RECT 132.250 162.440 135.775 162.580 ;
        RECT 132.250 162.380 132.570 162.440 ;
        RECT 135.485 162.395 135.775 162.440 ;
        RECT 136.405 162.580 136.695 162.625 ;
        RECT 137.310 162.580 137.630 162.640 ;
        RECT 147.890 162.580 148.210 162.640 ;
        RECT 136.405 162.440 137.630 162.580 ;
        RECT 136.405 162.395 136.695 162.440 ;
        RECT 137.310 162.380 137.630 162.440 ;
        RECT 146.600 162.440 148.210 162.580 ;
        RECT 112.485 162.100 116.380 162.240 ;
        RECT 112.485 162.055 112.775 162.100 ;
        RECT 95.910 161.900 96.230 161.960 ;
        RECT 116.240 161.945 116.380 162.100 ;
        RECT 129.490 162.100 130.410 162.240 ;
        RECT 130.870 162.240 131.190 162.300 ;
        RECT 130.870 162.100 131.560 162.240 ;
        RECT 129.490 162.040 129.810 162.100 ;
        RECT 130.870 162.040 131.190 162.100 ;
        RECT 105.585 161.900 105.875 161.945 ;
        RECT 95.910 161.760 105.875 161.900 ;
        RECT 95.910 161.700 96.230 161.760 ;
        RECT 105.585 161.715 105.875 161.760 ;
        RECT 106.465 161.900 106.755 161.945 ;
        RECT 107.655 161.900 107.945 161.945 ;
        RECT 110.175 161.900 110.465 161.945 ;
        RECT 106.465 161.760 110.465 161.900 ;
        RECT 106.465 161.715 106.755 161.760 ;
        RECT 107.655 161.715 107.945 161.760 ;
        RECT 110.175 161.715 110.465 161.760 ;
        RECT 116.165 161.900 116.455 161.945 ;
        RECT 121.670 161.900 121.990 161.960 ;
        RECT 131.420 161.900 131.560 162.100 ;
        RECT 133.630 162.040 133.950 162.300 ;
        RECT 139.165 162.055 139.455 162.285 ;
        RECT 141.910 162.240 142.200 162.285 ;
        RECT 143.480 162.240 143.770 162.285 ;
        RECT 145.580 162.240 145.870 162.285 ;
        RECT 141.910 162.100 145.870 162.240 ;
        RECT 141.910 162.055 142.200 162.100 ;
        RECT 143.480 162.055 143.770 162.100 ;
        RECT 145.580 162.055 145.870 162.100 ;
        RECT 139.240 161.900 139.380 162.055 ;
        RECT 146.600 161.945 146.740 162.440 ;
        RECT 147.890 162.380 148.210 162.440 ;
        RECT 147.010 162.240 147.300 162.285 ;
        RECT 149.110 162.240 149.400 162.285 ;
        RECT 150.680 162.240 150.970 162.285 ;
        RECT 147.010 162.100 150.970 162.240 ;
        RECT 147.010 162.055 147.300 162.100 ;
        RECT 149.110 162.055 149.400 162.100 ;
        RECT 150.680 162.055 150.970 162.100 ;
        RECT 116.165 161.760 121.990 161.900 ;
        RECT 116.165 161.715 116.455 161.760 ;
        RECT 121.670 161.700 121.990 161.760 ;
        RECT 130.500 161.760 139.380 161.900 ;
        RECT 141.475 161.900 141.765 161.945 ;
        RECT 143.995 161.900 144.285 161.945 ;
        RECT 145.185 161.900 145.475 161.945 ;
        RECT 141.475 161.760 145.475 161.900 ;
        RECT 93.625 161.560 93.915 161.605 ;
        RECT 96.370 161.560 96.690 161.620 ;
        RECT 93.240 161.420 93.915 161.560 ;
        RECT 89.945 161.375 90.235 161.420 ;
        RECT 92.705 161.375 92.995 161.420 ;
        RECT 93.625 161.375 93.915 161.420 ;
        RECT 94.160 161.420 96.690 161.560 ;
        RECT 92.780 161.220 92.920 161.375 ;
        RECT 94.160 161.220 94.300 161.420 ;
        RECT 96.370 161.360 96.690 161.420 ;
        RECT 100.510 161.360 100.830 161.620 ;
        RECT 100.970 161.560 101.290 161.620 ;
        RECT 100.970 161.420 104.420 161.560 ;
        RECT 100.970 161.360 101.290 161.420 ;
        RECT 92.780 161.080 94.300 161.220 ;
        RECT 95.450 161.220 95.770 161.280 ;
        RECT 102.825 161.220 103.115 161.265 ;
        RECT 95.450 161.080 103.115 161.220 ;
        RECT 95.450 161.020 95.770 161.080 ;
        RECT 102.825 161.035 103.115 161.080 ;
        RECT 98.210 160.880 98.530 160.940 ;
        RECT 89.100 160.740 98.530 160.880 ;
        RECT 85.330 160.680 85.650 160.740 ;
        RECT 87.645 160.695 87.935 160.740 ;
        RECT 98.210 160.680 98.530 160.740 ;
        RECT 99.590 160.880 99.910 160.940 ;
        RECT 101.445 160.880 101.735 160.925 ;
        RECT 101.890 160.880 102.210 160.940 ;
        RECT 104.280 160.925 104.420 161.420 ;
        RECT 120.750 161.360 121.070 161.620 ;
        RECT 122.130 161.360 122.450 161.620 ;
        RECT 123.970 161.360 124.290 161.620 ;
        RECT 125.350 161.360 125.670 161.620 ;
        RECT 126.270 161.605 126.590 161.620 ;
        RECT 126.105 161.375 126.590 161.605 ;
        RECT 127.895 161.560 128.185 161.605 ;
        RECT 129.950 161.560 130.270 161.620 ;
        RECT 127.895 161.420 130.270 161.560 ;
        RECT 130.500 161.560 130.640 161.760 ;
        RECT 141.475 161.715 141.765 161.760 ;
        RECT 143.995 161.715 144.285 161.760 ;
        RECT 145.185 161.715 145.475 161.760 ;
        RECT 146.065 161.900 146.355 161.945 ;
        RECT 146.525 161.900 146.815 161.945 ;
        RECT 146.065 161.760 146.815 161.900 ;
        RECT 146.065 161.715 146.355 161.760 ;
        RECT 146.525 161.715 146.815 161.760 ;
        RECT 147.405 161.900 147.695 161.945 ;
        RECT 148.595 161.900 148.885 161.945 ;
        RECT 151.115 161.900 151.405 161.945 ;
        RECT 147.405 161.760 151.405 161.900 ;
        RECT 147.405 161.715 147.695 161.760 ;
        RECT 148.595 161.715 148.885 161.760 ;
        RECT 151.115 161.715 151.405 161.760 ;
        RECT 130.845 161.560 131.135 161.605 ;
        RECT 130.500 161.420 131.135 161.560 ;
        RECT 127.895 161.375 128.185 161.420 ;
        RECT 126.270 161.360 126.590 161.375 ;
        RECT 129.950 161.360 130.270 161.420 ;
        RECT 130.845 161.375 131.135 161.420 ;
        RECT 106.950 161.265 107.270 161.280 ;
        RECT 106.920 161.035 107.270 161.265 ;
        RECT 106.950 161.020 107.270 161.035 ;
        RECT 109.710 161.220 110.030 161.280 ;
        RECT 113.405 161.220 113.695 161.265 ;
        RECT 122.605 161.220 122.895 161.265 ;
        RECT 109.710 161.080 113.695 161.220 ;
        RECT 109.710 161.020 110.030 161.080 ;
        RECT 113.405 161.035 113.695 161.080 ;
        RECT 113.940 161.080 122.895 161.220 ;
        RECT 99.590 160.740 102.210 160.880 ;
        RECT 99.590 160.680 99.910 160.740 ;
        RECT 101.445 160.695 101.735 160.740 ;
        RECT 101.890 160.680 102.210 160.740 ;
        RECT 104.205 160.880 104.495 160.925 ;
        RECT 112.010 160.880 112.330 160.940 ;
        RECT 113.940 160.880 114.080 161.080 ;
        RECT 122.605 161.035 122.895 161.080 ;
        RECT 123.065 161.035 123.355 161.265 ;
        RECT 124.890 161.220 125.210 161.280 ;
        RECT 126.745 161.220 127.035 161.265 ;
        RECT 124.890 161.080 127.035 161.220 ;
        RECT 104.205 160.740 114.080 160.880 ;
        RECT 114.310 160.880 114.630 160.940 ;
        RECT 117.545 160.880 117.835 160.925 ;
        RECT 114.310 160.740 117.835 160.880 ;
        RECT 104.205 160.695 104.495 160.740 ;
        RECT 112.010 160.680 112.330 160.740 ;
        RECT 114.310 160.680 114.630 160.740 ;
        RECT 117.545 160.695 117.835 160.740 ;
        RECT 118.910 160.880 119.230 160.940 ;
        RECT 123.140 160.880 123.280 161.035 ;
        RECT 124.890 161.020 125.210 161.080 ;
        RECT 126.745 161.035 127.035 161.080 ;
        RECT 127.205 161.220 127.495 161.265 ;
        RECT 129.490 161.220 129.810 161.280 ;
        RECT 127.205 161.080 129.810 161.220 ;
        RECT 127.205 161.035 127.495 161.080 ;
        RECT 129.490 161.020 129.810 161.080 ;
        RECT 133.170 161.220 133.490 161.280 ;
        RECT 144.210 161.220 144.530 161.280 ;
        RECT 147.890 161.265 148.210 161.280 ;
        RECT 144.730 161.220 145.020 161.265 ;
        RECT 133.170 161.080 143.520 161.220 ;
        RECT 133.170 161.020 133.490 161.080 ;
        RECT 118.910 160.740 123.280 160.880 ;
        RECT 128.585 160.880 128.875 160.925 ;
        RECT 131.790 160.880 132.110 160.940 ;
        RECT 128.585 160.740 132.110 160.880 ;
        RECT 118.910 160.680 119.230 160.740 ;
        RECT 128.585 160.695 128.875 160.740 ;
        RECT 131.790 160.680 132.110 160.740 ;
        RECT 135.485 160.880 135.775 160.925 ;
        RECT 136.390 160.880 136.710 160.940 ;
        RECT 135.485 160.740 136.710 160.880 ;
        RECT 143.380 160.880 143.520 161.080 ;
        RECT 144.210 161.080 145.020 161.220 ;
        RECT 144.210 161.020 144.530 161.080 ;
        RECT 144.730 161.035 145.020 161.080 ;
        RECT 147.860 161.035 148.210 161.265 ;
        RECT 147.890 161.020 148.210 161.035 ;
        RECT 153.425 160.880 153.715 160.925 ;
        RECT 154.790 160.880 155.110 160.940 ;
        RECT 143.380 160.740 155.110 160.880 ;
        RECT 135.485 160.695 135.775 160.740 ;
        RECT 136.390 160.680 136.710 160.740 ;
        RECT 153.425 160.695 153.715 160.740 ;
        RECT 154.790 160.680 155.110 160.740 ;
        RECT 22.700 160.060 157.820 160.540 ;
        RECT 24.610 159.660 24.930 159.920 ;
        RECT 26.910 159.905 27.230 159.920 ;
        RECT 26.005 159.675 26.295 159.905 ;
        RECT 26.845 159.675 27.230 159.905 ;
        RECT 36.110 159.860 36.430 159.920 ;
        RECT 68.770 159.860 69.090 159.920 ;
        RECT 25.545 159.180 25.835 159.225 ;
        RECT 26.080 159.180 26.220 159.675 ;
        RECT 26.910 159.660 27.230 159.675 ;
        RECT 33.670 159.720 69.090 159.860 ;
        RECT 27.830 159.320 28.150 159.580 ;
        RECT 32.905 159.520 33.195 159.565 ;
        RECT 33.670 159.520 33.810 159.720 ;
        RECT 36.110 159.660 36.430 159.720 ;
        RECT 32.905 159.380 33.810 159.520 ;
        RECT 32.905 159.335 33.195 159.380 ;
        RECT 43.930 159.320 44.250 159.580 ;
        RECT 45.785 159.520 46.075 159.565 ;
        RECT 44.480 159.380 46.075 159.520 ;
        RECT 25.545 159.040 26.220 159.180 ;
        RECT 33.365 159.180 33.655 159.225 ;
        RECT 34.270 159.180 34.590 159.240 ;
        RECT 33.365 159.040 34.590 159.180 ;
        RECT 25.545 158.995 25.835 159.040 ;
        RECT 33.365 158.995 33.655 159.040 ;
        RECT 34.270 158.980 34.590 159.040 ;
        RECT 36.125 159.180 36.415 159.225 ;
        RECT 36.570 159.180 36.890 159.240 ;
        RECT 38.425 159.180 38.715 159.225 ;
        RECT 44.480 159.180 44.620 159.380 ;
        RECT 45.785 159.335 46.075 159.380 ;
        RECT 46.230 159.520 46.550 159.580 ;
        RECT 53.590 159.520 53.910 159.580 ;
        RECT 54.600 159.565 54.740 159.720 ;
        RECT 68.770 159.660 69.090 159.720 ;
        RECT 93.625 159.860 93.915 159.905 ;
        RECT 96.370 159.860 96.690 159.920 ;
        RECT 93.625 159.720 96.690 159.860 ;
        RECT 93.625 159.675 93.915 159.720 ;
        RECT 96.370 159.660 96.690 159.720 ;
        RECT 98.670 159.860 98.990 159.920 ;
        RECT 98.670 159.720 103.500 159.860 ;
        RECT 98.670 159.660 98.990 159.720 ;
        RECT 46.230 159.380 53.910 159.520 ;
        RECT 46.230 159.320 46.550 159.380 ;
        RECT 53.590 159.320 53.910 159.380 ;
        RECT 54.525 159.335 54.815 159.565 ;
        RECT 62.330 159.320 62.650 159.580 ;
        RECT 67.405 159.520 67.695 159.565 ;
        RECT 69.230 159.520 69.550 159.580 ;
        RECT 79.350 159.520 79.670 159.580 ;
        RECT 80.730 159.520 81.050 159.580 ;
        RECT 63.495 159.350 63.785 159.395 ;
        RECT 67.405 159.380 69.550 159.520 ;
        RECT 63.495 159.240 63.895 159.350 ;
        RECT 67.405 159.335 67.695 159.380 ;
        RECT 69.230 159.320 69.550 159.380 ;
        RECT 77.600 159.380 79.670 159.520 ;
        RECT 36.125 159.040 38.715 159.180 ;
        RECT 36.125 158.995 36.415 159.040 ;
        RECT 36.570 158.980 36.890 159.040 ;
        RECT 38.425 158.995 38.715 159.040 ;
        RECT 38.960 159.040 44.620 159.180 ;
        RECT 24.150 158.840 24.470 158.900 ;
        RECT 28.765 158.840 29.055 158.885 ;
        RECT 24.150 158.700 29.055 158.840 ;
        RECT 24.150 158.640 24.470 158.700 ;
        RECT 28.765 158.655 29.055 158.700 ;
        RECT 33.810 158.840 34.130 158.900 ;
        RECT 35.665 158.840 35.955 158.885 ;
        RECT 38.960 158.840 39.100 159.040 ;
        RECT 45.325 158.995 45.615 159.225 ;
        RECT 33.810 158.700 39.100 158.840 ;
        RECT 33.810 158.640 34.130 158.700 ;
        RECT 35.665 158.655 35.955 158.700 ;
        RECT 40.710 158.640 41.030 158.900 ;
        RECT 41.630 158.640 41.950 158.900 ;
        RECT 42.090 158.640 42.410 158.900 ;
        RECT 42.550 158.640 42.870 158.900 ;
        RECT 43.025 158.840 43.315 158.885 ;
        RECT 43.025 158.700 44.620 158.840 ;
        RECT 43.025 158.655 43.315 158.700 ;
        RECT 44.480 158.560 44.620 158.700 ;
        RECT 34.285 158.500 34.575 158.545 ;
        RECT 34.730 158.500 35.050 158.560 ;
        RECT 34.285 158.360 35.050 158.500 ;
        RECT 34.285 158.315 34.575 158.360 ;
        RECT 34.730 158.300 35.050 158.360 ;
        RECT 44.390 158.300 44.710 158.560 ;
        RECT 45.400 158.500 45.540 158.995 ;
        RECT 47.150 158.980 47.470 159.240 ;
        RECT 50.830 159.180 51.150 159.240 ;
        RECT 54.050 159.180 54.370 159.240 ;
        RECT 50.830 159.040 54.370 159.180 ;
        RECT 50.830 158.980 51.150 159.040 ;
        RECT 54.050 158.980 54.370 159.040 ;
        RECT 60.490 159.225 60.810 159.240 ;
        RECT 60.490 158.995 60.840 159.225 ;
        RECT 62.790 159.180 63.110 159.240 ;
        RECT 63.495 159.180 64.030 159.240 ;
        RECT 66.485 159.180 66.775 159.225 ;
        RECT 62.790 159.040 66.775 159.180 ;
        RECT 60.490 158.980 60.810 158.995 ;
        RECT 62.790 158.980 63.110 159.040 ;
        RECT 63.710 158.980 64.030 159.040 ;
        RECT 66.485 158.995 66.775 159.040 ;
        RECT 68.310 158.980 68.630 159.240 ;
        RECT 71.545 158.995 71.835 159.225 ;
        RECT 72.465 159.180 72.755 159.225 ;
        RECT 73.845 159.180 74.135 159.225 ;
        RECT 72.465 159.040 74.135 159.180 ;
        RECT 72.465 158.995 72.755 159.040 ;
        RECT 73.845 158.995 74.135 159.040 ;
        RECT 48.530 158.840 48.850 158.900 ;
        RECT 50.385 158.840 50.675 158.885 ;
        RECT 48.530 158.700 50.675 158.840 ;
        RECT 48.530 158.640 48.850 158.700 ;
        RECT 50.385 158.655 50.675 158.700 ;
        RECT 57.295 158.840 57.585 158.885 ;
        RECT 59.815 158.840 60.105 158.885 ;
        RECT 61.005 158.840 61.295 158.885 ;
        RECT 57.295 158.700 61.295 158.840 ;
        RECT 57.295 158.655 57.585 158.700 ;
        RECT 59.815 158.655 60.105 158.700 ;
        RECT 61.005 158.655 61.295 158.700 ;
        RECT 61.885 158.840 62.175 158.885 ;
        RECT 64.170 158.840 64.490 158.900 ;
        RECT 67.850 158.840 68.170 158.900 ;
        RECT 61.885 158.700 68.170 158.840 ;
        RECT 61.885 158.655 62.175 158.700 ;
        RECT 64.170 158.640 64.490 158.700 ;
        RECT 67.850 158.640 68.170 158.700 ;
        RECT 70.610 158.640 70.930 158.900 ;
        RECT 71.620 158.840 71.760 158.995 ;
        RECT 77.050 158.980 77.370 159.240 ;
        RECT 76.590 158.840 76.910 158.900 ;
        RECT 77.600 158.885 77.740 159.380 ;
        RECT 79.350 159.320 79.670 159.380 ;
        RECT 80.440 159.320 81.050 159.520 ;
        RECT 80.440 159.210 80.805 159.320 ;
        RECT 80.515 159.165 80.805 159.210 ;
        RECT 81.665 159.180 81.955 159.225 ;
        RECT 81.280 159.040 81.955 159.180 ;
        RECT 77.525 158.840 77.815 158.885 ;
        RECT 71.620 158.700 75.440 158.840 ;
        RECT 54.970 158.500 55.290 158.560 ;
        RECT 45.400 158.360 55.290 158.500 ;
        RECT 26.925 158.160 27.215 158.205 ;
        RECT 31.970 158.160 32.290 158.220 ;
        RECT 26.925 158.020 32.290 158.160 ;
        RECT 26.925 157.975 27.215 158.020 ;
        RECT 31.970 157.960 32.290 158.020 ;
        RECT 39.805 158.160 40.095 158.205 ;
        RECT 45.400 158.160 45.540 158.360 ;
        RECT 54.970 158.300 55.290 158.360 ;
        RECT 57.730 158.500 58.020 158.545 ;
        RECT 59.300 158.500 59.590 158.545 ;
        RECT 61.400 158.500 61.690 158.545 ;
        RECT 68.310 158.500 68.630 158.560 ;
        RECT 57.730 158.360 61.690 158.500 ;
        RECT 57.730 158.315 58.020 158.360 ;
        RECT 59.300 158.315 59.590 158.360 ;
        RECT 61.400 158.315 61.690 158.360 ;
        RECT 62.880 158.360 68.630 158.500 ;
        RECT 70.700 158.500 70.840 158.640 ;
        RECT 75.300 158.545 75.440 158.700 ;
        RECT 76.590 158.700 77.815 158.840 ;
        RECT 76.590 158.640 76.910 158.700 ;
        RECT 77.525 158.655 77.815 158.700 ;
        RECT 78.430 158.640 78.750 158.900 ;
        RECT 81.280 158.545 81.420 159.040 ;
        RECT 81.665 158.995 81.955 159.040 ;
        RECT 84.870 158.980 85.190 159.240 ;
        RECT 85.330 158.980 85.650 159.240 ;
        RECT 86.710 158.980 87.030 159.240 ;
        RECT 88.090 159.225 88.410 159.240 ;
        RECT 88.060 158.995 88.410 159.225 ;
        RECT 95.925 159.180 96.215 159.225 ;
        RECT 96.370 159.180 96.690 159.240 ;
        RECT 95.925 159.040 96.690 159.180 ;
        RECT 95.925 158.995 96.215 159.040 ;
        RECT 88.090 158.980 88.410 158.995 ;
        RECT 96.370 158.980 96.690 159.040 ;
        RECT 96.830 158.980 97.150 159.240 ;
        RECT 97.290 158.980 97.610 159.240 ;
        RECT 100.970 158.980 101.290 159.240 ;
        RECT 101.905 158.995 102.195 159.225 ;
        RECT 103.360 159.180 103.500 159.720 ;
        RECT 106.950 159.660 107.270 159.920 ;
        RECT 114.785 159.675 115.075 159.905 ;
        RECT 120.750 159.860 121.070 159.920 ;
        RECT 122.145 159.860 122.435 159.905 ;
        RECT 120.750 159.720 122.435 159.860 ;
        RECT 114.310 159.520 114.630 159.580 ;
        RECT 112.100 159.380 114.630 159.520 ;
        RECT 114.860 159.520 115.000 159.675 ;
        RECT 120.750 159.660 121.070 159.720 ;
        RECT 122.145 159.675 122.435 159.720 ;
        RECT 116.470 159.520 116.760 159.565 ;
        RECT 114.860 159.380 116.760 159.520 ;
        RECT 122.220 159.520 122.360 159.675 ;
        RECT 124.890 159.660 125.210 159.920 ;
        RECT 125.350 159.860 125.670 159.920 ;
        RECT 126.285 159.860 126.575 159.905 ;
        RECT 125.350 159.720 126.575 159.860 ;
        RECT 125.350 159.660 125.670 159.720 ;
        RECT 126.285 159.675 126.575 159.720 ;
        RECT 126.730 159.860 127.050 159.920 ;
        RECT 129.045 159.860 129.335 159.905 ;
        RECT 126.730 159.720 129.335 159.860 ;
        RECT 126.730 159.660 127.050 159.720 ;
        RECT 129.045 159.675 129.335 159.720 ;
        RECT 147.890 159.660 148.210 159.920 ;
        RECT 129.950 159.520 130.270 159.580 ;
        RECT 122.220 159.380 130.270 159.520 ;
        RECT 104.665 159.180 104.955 159.225 ;
        RECT 103.360 159.040 104.955 159.180 ;
        RECT 104.665 158.995 104.955 159.040 ;
        RECT 105.110 159.180 105.430 159.240 ;
        RECT 105.585 159.180 105.875 159.225 ;
        RECT 105.110 159.040 105.875 159.180 ;
        RECT 84.960 158.840 85.100 158.980 ;
        RECT 81.640 158.700 85.100 158.840 ;
        RECT 87.605 158.840 87.895 158.885 ;
        RECT 88.795 158.840 89.085 158.885 ;
        RECT 91.315 158.840 91.605 158.885 ;
        RECT 87.605 158.700 91.605 158.840 ;
        RECT 70.700 158.360 74.980 158.500 ;
        RECT 39.805 158.020 45.540 158.160 ;
        RECT 46.690 158.160 47.010 158.220 ;
        RECT 62.880 158.160 63.020 158.360 ;
        RECT 68.310 158.300 68.630 158.360 ;
        RECT 46.690 158.020 63.020 158.160 ;
        RECT 39.805 157.975 40.095 158.020 ;
        RECT 46.690 157.960 47.010 158.020 ;
        RECT 63.250 157.960 63.570 158.220 ;
        RECT 64.170 157.960 64.490 158.220 ;
        RECT 71.070 158.160 71.390 158.220 ;
        RECT 72.925 158.160 73.215 158.205 ;
        RECT 71.070 158.020 73.215 158.160 ;
        RECT 74.840 158.160 74.980 158.360 ;
        RECT 75.225 158.315 75.515 158.545 ;
        RECT 79.900 158.360 80.960 158.500 ;
        RECT 79.900 158.160 80.040 158.360 ;
        RECT 74.840 158.020 80.040 158.160 ;
        RECT 71.070 157.960 71.390 158.020 ;
        RECT 72.925 157.975 73.215 158.020 ;
        RECT 80.270 157.960 80.590 158.220 ;
        RECT 80.820 158.160 80.960 158.360 ;
        RECT 81.205 158.315 81.495 158.545 ;
        RECT 81.640 158.160 81.780 158.700 ;
        RECT 87.605 158.655 87.895 158.700 ;
        RECT 88.795 158.655 89.085 158.700 ;
        RECT 91.315 158.655 91.605 158.700 ;
        RECT 94.990 158.640 95.310 158.900 ;
        RECT 98.210 158.840 98.530 158.900 ;
        RECT 101.980 158.840 102.120 158.995 ;
        RECT 105.110 158.980 105.430 159.040 ;
        RECT 105.585 158.995 105.875 159.040 ;
        RECT 107.885 158.995 108.175 159.225 ;
        RECT 98.210 158.700 102.120 158.840 ;
        RECT 106.505 158.840 106.795 158.885 ;
        RECT 107.960 158.840 108.100 158.995 ;
        RECT 108.330 158.980 108.650 159.240 ;
        RECT 108.790 158.980 109.110 159.240 ;
        RECT 109.710 158.980 110.030 159.240 ;
        RECT 112.100 159.225 112.240 159.380 ;
        RECT 114.310 159.320 114.630 159.380 ;
        RECT 116.470 159.335 116.760 159.380 ;
        RECT 129.950 159.320 130.270 159.380 ;
        RECT 131.330 159.320 131.650 159.580 ;
        RECT 136.390 159.320 136.710 159.580 ;
        RECT 137.310 159.565 137.630 159.580 ;
        RECT 137.310 159.335 137.695 159.565 ;
        RECT 152.045 159.520 152.335 159.565 ;
        RECT 144.300 159.380 152.335 159.520 ;
        RECT 137.310 159.320 137.630 159.335 ;
        RECT 112.025 158.995 112.315 159.225 ;
        RECT 112.945 158.995 113.235 159.225 ;
        RECT 109.250 158.840 109.570 158.900 ;
        RECT 106.505 158.700 109.570 158.840 ;
        RECT 98.210 158.640 98.530 158.700 ;
        RECT 106.505 158.655 106.795 158.700 ;
        RECT 109.250 158.640 109.570 158.700 ;
        RECT 87.210 158.500 87.500 158.545 ;
        RECT 89.310 158.500 89.600 158.545 ;
        RECT 90.880 158.500 91.170 158.545 ;
        RECT 87.210 158.360 91.170 158.500 ;
        RECT 87.210 158.315 87.500 158.360 ;
        RECT 89.310 158.315 89.600 158.360 ;
        RECT 90.880 158.315 91.170 158.360 ;
        RECT 108.790 158.500 109.110 158.560 ;
        RECT 113.020 158.500 113.160 158.995 ;
        RECT 113.390 158.980 113.710 159.240 ;
        RECT 113.865 159.180 114.155 159.225 ;
        RECT 122.130 159.180 122.450 159.240 ;
        RECT 113.865 159.040 122.450 159.180 ;
        RECT 113.865 158.995 114.155 159.040 ;
        RECT 122.130 158.980 122.450 159.040 ;
        RECT 122.605 159.180 122.895 159.225 ;
        RECT 128.585 159.180 128.875 159.225 ;
        RECT 131.420 159.180 131.560 159.320 ;
        RECT 122.605 159.040 131.560 159.180 ;
        RECT 132.725 159.180 133.015 159.225 ;
        RECT 135.930 159.180 136.250 159.240 ;
        RECT 144.300 159.225 144.440 159.380 ;
        RECT 152.045 159.335 152.335 159.380 ;
        RECT 132.725 159.040 136.250 159.180 ;
        RECT 122.605 158.995 122.895 159.040 ;
        RECT 128.585 158.995 128.875 159.040 ;
        RECT 132.725 158.995 133.015 159.040 ;
        RECT 135.930 158.980 136.250 159.040 ;
        RECT 144.225 158.995 144.515 159.225 ;
        RECT 146.985 159.180 147.275 159.225 ;
        RECT 147.905 159.180 148.195 159.225 ;
        RECT 146.140 159.040 147.275 159.180 ;
        RECT 114.770 158.840 115.090 158.900 ;
        RECT 115.245 158.840 115.535 158.885 ;
        RECT 114.770 158.700 115.535 158.840 ;
        RECT 114.770 158.640 115.090 158.700 ;
        RECT 115.245 158.655 115.535 158.700 ;
        RECT 116.125 158.840 116.415 158.885 ;
        RECT 117.315 158.840 117.605 158.885 ;
        RECT 119.835 158.840 120.125 158.885 ;
        RECT 116.125 158.700 120.125 158.840 ;
        RECT 116.125 158.655 116.415 158.700 ;
        RECT 117.315 158.655 117.605 158.700 ;
        RECT 119.835 158.655 120.125 158.700 ;
        RECT 131.345 158.840 131.635 158.885 ;
        RECT 133.170 158.840 133.490 158.900 ;
        RECT 131.345 158.700 133.490 158.840 ;
        RECT 131.345 158.655 131.635 158.700 ;
        RECT 133.170 158.640 133.490 158.700 ;
        RECT 144.685 158.840 144.975 158.885 ;
        RECT 145.130 158.840 145.450 158.900 ;
        RECT 144.685 158.700 145.450 158.840 ;
        RECT 144.685 158.655 144.975 158.700 ;
        RECT 145.130 158.640 145.450 158.700 ;
        RECT 115.730 158.500 116.020 158.545 ;
        RECT 117.830 158.500 118.120 158.545 ;
        RECT 119.400 158.500 119.690 158.545 ;
        RECT 108.790 158.360 113.620 158.500 ;
        RECT 108.790 158.300 109.110 158.360 ;
        RECT 80.820 158.020 81.780 158.160 ;
        RECT 82.110 157.960 82.430 158.220 ;
        RECT 86.265 158.160 86.555 158.205 ;
        RECT 87.630 158.160 87.950 158.220 ;
        RECT 86.265 158.020 87.950 158.160 ;
        RECT 86.265 157.975 86.555 158.020 ;
        RECT 87.630 157.960 87.950 158.020 ;
        RECT 88.550 158.160 88.870 158.220 ;
        RECT 98.670 158.160 98.990 158.220 ;
        RECT 88.550 158.020 98.990 158.160 ;
        RECT 88.550 157.960 88.870 158.020 ;
        RECT 98.670 157.960 98.990 158.020 ;
        RECT 101.430 157.960 101.750 158.220 ;
        RECT 113.480 158.160 113.620 158.360 ;
        RECT 115.730 158.360 119.690 158.500 ;
        RECT 115.730 158.315 116.020 158.360 ;
        RECT 117.830 158.315 118.120 158.360 ;
        RECT 119.400 158.315 119.690 158.360 ;
        RECT 121.670 158.500 121.990 158.560 ;
        RECT 126.745 158.500 127.035 158.545 ;
        RECT 121.670 158.360 127.035 158.500 ;
        RECT 121.670 158.300 121.990 158.360 ;
        RECT 118.910 158.160 119.230 158.220 ;
        RECT 123.140 158.205 123.280 158.360 ;
        RECT 126.745 158.315 127.035 158.360 ;
        RECT 127.190 158.500 127.510 158.560 ;
        RECT 129.505 158.500 129.795 158.545 ;
        RECT 127.190 158.360 129.795 158.500 ;
        RECT 127.190 158.300 127.510 158.360 ;
        RECT 129.505 158.315 129.795 158.360 ;
        RECT 136.390 158.500 136.710 158.560 ;
        RECT 146.140 158.545 146.280 159.040 ;
        RECT 146.985 158.995 147.275 159.040 ;
        RECT 147.520 159.040 148.195 159.180 ;
        RECT 136.390 158.360 145.820 158.500 ;
        RECT 136.390 158.300 136.710 158.360 ;
        RECT 113.480 158.020 119.230 158.160 ;
        RECT 118.910 157.960 119.230 158.020 ;
        RECT 123.065 157.975 123.355 158.205 ;
        RECT 132.250 157.960 132.570 158.220 ;
        RECT 137.325 158.160 137.615 158.205 ;
        RECT 137.770 158.160 138.090 158.220 ;
        RECT 137.325 158.020 138.090 158.160 ;
        RECT 137.325 157.975 137.615 158.020 ;
        RECT 137.770 157.960 138.090 158.020 ;
        RECT 138.245 158.160 138.535 158.205 ;
        RECT 138.690 158.160 139.010 158.220 ;
        RECT 138.245 158.020 139.010 158.160 ;
        RECT 145.680 158.160 145.820 158.360 ;
        RECT 146.065 158.315 146.355 158.545 ;
        RECT 147.520 158.160 147.660 159.040 ;
        RECT 147.905 158.995 148.195 159.040 ;
        RECT 154.790 158.980 155.110 159.240 ;
        RECT 145.680 158.020 147.660 158.160 ;
        RECT 138.245 157.975 138.535 158.020 ;
        RECT 138.690 157.960 139.010 158.020 ;
        RECT 22.700 157.340 157.020 157.820 ;
        RECT 29.225 157.140 29.515 157.185 ;
        RECT 31.510 157.140 31.830 157.200 ;
        RECT 29.225 157.000 31.830 157.140 ;
        RECT 29.225 156.955 29.515 157.000 ;
        RECT 31.510 156.940 31.830 157.000 ;
        RECT 32.445 157.140 32.735 157.185 ;
        RECT 33.350 157.140 33.670 157.200 ;
        RECT 32.445 157.000 33.670 157.140 ;
        RECT 32.445 156.955 32.735 157.000 ;
        RECT 33.350 156.940 33.670 157.000 ;
        RECT 39.345 157.140 39.635 157.185 ;
        RECT 42.105 157.140 42.395 157.185 ;
        RECT 42.550 157.140 42.870 157.200 ;
        RECT 39.345 157.000 40.020 157.140 ;
        RECT 39.345 156.955 39.635 157.000 ;
        RECT 30.130 156.460 30.450 156.520 ;
        RECT 33.825 156.460 34.115 156.505 ;
        RECT 30.130 156.320 31.740 156.460 ;
        RECT 30.130 156.260 30.450 156.320 ;
        RECT 30.605 156.120 30.895 156.165 ;
        RECT 31.050 156.120 31.370 156.180 ;
        RECT 31.600 156.165 31.740 156.320 ;
        RECT 32.060 156.320 34.115 156.460 ;
        RECT 32.060 156.180 32.200 156.320 ;
        RECT 33.825 156.275 34.115 156.320 ;
        RECT 30.605 155.980 31.370 156.120 ;
        RECT 30.605 155.935 30.895 155.980 ;
        RECT 31.050 155.920 31.370 155.980 ;
        RECT 31.525 155.935 31.815 156.165 ;
        RECT 31.970 155.920 32.290 156.180 ;
        RECT 32.905 155.935 33.195 156.165 ;
        RECT 27.830 155.780 28.150 155.840 ;
        RECT 30.145 155.780 30.435 155.825 ;
        RECT 27.830 155.640 30.435 155.780 ;
        RECT 32.980 155.780 33.120 155.935 ;
        RECT 33.350 155.920 33.670 156.180 ;
        RECT 34.285 155.935 34.575 156.165 ;
        RECT 36.570 156.120 36.890 156.180 ;
        RECT 37.965 156.120 38.255 156.165 ;
        RECT 36.570 155.980 38.255 156.120 ;
        RECT 33.810 155.780 34.130 155.840 ;
        RECT 32.980 155.640 34.130 155.780 ;
        RECT 27.830 155.580 28.150 155.640 ;
        RECT 30.145 155.595 30.435 155.640 ;
        RECT 33.810 155.580 34.130 155.640 ;
        RECT 25.990 155.440 26.310 155.500 ;
        RECT 29.210 155.485 29.530 155.500 ;
        RECT 28.305 155.440 28.595 155.485 ;
        RECT 25.990 155.300 28.595 155.440 ;
        RECT 25.990 155.240 26.310 155.300 ;
        RECT 28.305 155.255 28.595 155.300 ;
        RECT 29.145 155.440 29.530 155.485 ;
        RECT 30.605 155.440 30.895 155.485 ;
        RECT 29.145 155.300 30.895 155.440 ;
        RECT 29.145 155.255 29.530 155.300 ;
        RECT 30.605 155.255 30.895 155.300 ;
        RECT 32.430 155.440 32.750 155.500 ;
        RECT 34.360 155.440 34.500 155.935 ;
        RECT 36.570 155.920 36.890 155.980 ;
        RECT 37.965 155.935 38.255 155.980 ;
        RECT 32.430 155.300 34.500 155.440 ;
        RECT 38.870 155.440 39.190 155.500 ;
        RECT 39.880 155.440 40.020 157.000 ;
        RECT 42.105 157.000 42.870 157.140 ;
        RECT 42.105 156.955 42.395 157.000 ;
        RECT 42.550 156.940 42.870 157.000 ;
        RECT 45.325 157.140 45.615 157.185 ;
        RECT 46.230 157.140 46.550 157.200 ;
        RECT 45.325 157.000 46.550 157.140 ;
        RECT 45.325 156.955 45.615 157.000 ;
        RECT 46.230 156.940 46.550 157.000 ;
        RECT 53.590 157.140 53.910 157.200 ;
        RECT 54.985 157.140 55.275 157.185 ;
        RECT 53.590 157.000 55.275 157.140 ;
        RECT 53.590 156.940 53.910 157.000 ;
        RECT 54.985 156.955 55.275 157.000 ;
        RECT 59.585 157.140 59.875 157.185 ;
        RECT 60.490 157.140 60.810 157.200 ;
        RECT 59.585 157.000 60.810 157.140 ;
        RECT 59.585 156.955 59.875 157.000 ;
        RECT 60.490 156.940 60.810 157.000 ;
        RECT 61.885 157.140 62.175 157.185 ;
        RECT 62.330 157.140 62.650 157.200 ;
        RECT 61.885 157.000 62.650 157.140 ;
        RECT 61.885 156.955 62.175 157.000 ;
        RECT 62.330 156.940 62.650 157.000 ;
        RECT 76.590 156.940 76.910 157.200 ;
        RECT 88.090 157.140 88.410 157.200 ;
        RECT 88.565 157.140 88.855 157.185 ;
        RECT 88.090 157.000 88.855 157.140 ;
        RECT 88.090 156.940 88.410 157.000 ;
        RECT 88.565 156.955 88.855 157.000 ;
        RECT 96.830 157.140 97.150 157.200 ;
        RECT 98.670 157.140 98.990 157.200 ;
        RECT 99.605 157.140 99.895 157.185 ;
        RECT 119.370 157.140 119.690 157.200 ;
        RECT 130.410 157.140 130.730 157.200 ;
        RECT 96.830 157.000 99.895 157.140 ;
        RECT 96.830 156.940 97.150 157.000 ;
        RECT 98.670 156.940 98.990 157.000 ;
        RECT 99.605 156.955 99.895 157.000 ;
        RECT 101.980 157.000 119.690 157.140 ;
        RECT 41.630 156.800 41.950 156.860 ;
        RECT 43.485 156.800 43.775 156.845 ;
        RECT 41.630 156.660 43.775 156.800 ;
        RECT 41.630 156.600 41.950 156.660 ;
        RECT 43.485 156.615 43.775 156.660 ;
        RECT 48.570 156.800 48.860 156.845 ;
        RECT 50.670 156.800 50.960 156.845 ;
        RECT 52.240 156.800 52.530 156.845 ;
        RECT 48.570 156.660 52.530 156.800 ;
        RECT 48.570 156.615 48.860 156.660 ;
        RECT 50.670 156.615 50.960 156.660 ;
        RECT 52.240 156.615 52.530 156.660 ;
        RECT 64.630 156.800 64.920 156.845 ;
        RECT 66.200 156.800 66.490 156.845 ;
        RECT 68.300 156.800 68.590 156.845 ;
        RECT 64.630 156.660 68.590 156.800 ;
        RECT 64.630 156.615 64.920 156.660 ;
        RECT 66.200 156.615 66.490 156.660 ;
        RECT 68.300 156.615 68.590 156.660 ;
        RECT 70.190 156.800 70.480 156.845 ;
        RECT 72.290 156.800 72.580 156.845 ;
        RECT 73.860 156.800 74.150 156.845 ;
        RECT 70.190 156.660 74.150 156.800 ;
        RECT 70.190 156.615 70.480 156.660 ;
        RECT 72.290 156.615 72.580 156.660 ;
        RECT 73.860 156.615 74.150 156.660 ;
        RECT 91.810 156.800 92.100 156.845 ;
        RECT 93.910 156.800 94.200 156.845 ;
        RECT 95.480 156.800 95.770 156.845 ;
        RECT 91.810 156.660 95.770 156.800 ;
        RECT 91.810 156.615 92.100 156.660 ;
        RECT 93.910 156.615 94.200 156.660 ;
        RECT 95.480 156.615 95.770 156.660 ;
        RECT 99.130 156.800 99.450 156.860 ;
        RECT 101.980 156.800 102.120 157.000 ;
        RECT 119.370 156.940 119.690 157.000 ;
        RECT 119.920 157.000 130.730 157.140 ;
        RECT 99.130 156.660 102.120 156.800 ;
        RECT 102.350 156.800 102.640 156.845 ;
        RECT 103.920 156.800 104.210 156.845 ;
        RECT 106.020 156.800 106.310 156.845 ;
        RECT 102.350 156.660 106.310 156.800 ;
        RECT 99.130 156.600 99.450 156.660 ;
        RECT 102.350 156.615 102.640 156.660 ;
        RECT 103.920 156.615 104.210 156.660 ;
        RECT 106.020 156.615 106.310 156.660 ;
        RECT 108.790 156.800 109.110 156.860 ;
        RECT 109.265 156.800 109.555 156.845 ;
        RECT 108.790 156.660 109.555 156.800 ;
        RECT 108.790 156.600 109.110 156.660 ;
        RECT 109.265 156.615 109.555 156.660 ;
        RECT 40.265 156.275 40.555 156.505 ;
        RECT 40.710 156.460 41.030 156.520 ;
        RECT 45.785 156.460 46.075 156.505 ;
        RECT 47.150 156.460 47.470 156.520 ;
        RECT 40.710 156.320 42.780 156.460 ;
        RECT 40.340 156.120 40.480 156.275 ;
        RECT 40.710 156.260 41.030 156.320 ;
        RECT 41.170 156.120 41.490 156.180 ;
        RECT 42.640 156.165 42.780 156.320 ;
        RECT 45.785 156.320 47.470 156.460 ;
        RECT 45.785 156.275 46.075 156.320 ;
        RECT 47.150 156.260 47.470 156.320 ;
        RECT 48.965 156.460 49.255 156.505 ;
        RECT 50.155 156.460 50.445 156.505 ;
        RECT 52.675 156.460 52.965 156.505 ;
        RECT 48.965 156.320 52.965 156.460 ;
        RECT 48.965 156.275 49.255 156.320 ;
        RECT 50.155 156.275 50.445 156.320 ;
        RECT 52.675 156.275 52.965 156.320 ;
        RECT 64.195 156.460 64.485 156.505 ;
        RECT 66.715 156.460 67.005 156.505 ;
        RECT 67.905 156.460 68.195 156.505 ;
        RECT 64.195 156.320 68.195 156.460 ;
        RECT 64.195 156.275 64.485 156.320 ;
        RECT 66.715 156.275 67.005 156.320 ;
        RECT 67.905 156.275 68.195 156.320 ;
        RECT 70.585 156.460 70.875 156.505 ;
        RECT 71.775 156.460 72.065 156.505 ;
        RECT 74.295 156.460 74.585 156.505 ;
        RECT 70.585 156.320 74.585 156.460 ;
        RECT 70.585 156.275 70.875 156.320 ;
        RECT 71.775 156.275 72.065 156.320 ;
        RECT 74.295 156.275 74.585 156.320 ;
        RECT 86.710 156.460 87.030 156.520 ;
        RECT 91.325 156.460 91.615 156.505 ;
        RECT 86.710 156.320 91.615 156.460 ;
        RECT 86.710 156.260 87.030 156.320 ;
        RECT 91.325 156.275 91.615 156.320 ;
        RECT 92.205 156.460 92.495 156.505 ;
        RECT 93.395 156.460 93.685 156.505 ;
        RECT 95.915 156.460 96.205 156.505 ;
        RECT 92.205 156.320 96.205 156.460 ;
        RECT 92.205 156.275 92.495 156.320 ;
        RECT 93.395 156.275 93.685 156.320 ;
        RECT 95.915 156.275 96.205 156.320 ;
        RECT 101.915 156.460 102.205 156.505 ;
        RECT 104.435 156.460 104.725 156.505 ;
        RECT 105.625 156.460 105.915 156.505 ;
        RECT 101.915 156.320 105.915 156.460 ;
        RECT 101.915 156.275 102.205 156.320 ;
        RECT 104.435 156.275 104.725 156.320 ;
        RECT 105.625 156.275 105.915 156.320 ;
        RECT 106.505 156.460 106.795 156.505 ;
        RECT 109.710 156.460 110.030 156.520 ;
        RECT 106.505 156.320 110.030 156.460 ;
        RECT 106.505 156.275 106.795 156.320 ;
        RECT 109.710 156.260 110.030 156.320 ;
        RECT 113.390 156.460 113.710 156.520 ;
        RECT 116.625 156.460 116.915 156.505 ;
        RECT 119.920 156.460 120.060 157.000 ;
        RECT 130.410 156.940 130.730 157.000 ;
        RECT 136.865 157.140 137.155 157.185 ;
        RECT 137.310 157.140 137.630 157.200 ;
        RECT 136.865 157.000 137.630 157.140 ;
        RECT 136.865 156.955 137.155 157.000 ;
        RECT 137.310 156.940 137.630 157.000 ;
        RECT 141.005 156.800 141.295 156.845 ;
        RECT 121.760 156.660 128.800 156.800 ;
        RECT 113.390 156.320 120.060 156.460 ;
        RECT 120.290 156.460 120.610 156.520 ;
        RECT 121.760 156.505 121.900 156.660 ;
        RECT 128.660 156.520 128.800 156.660 ;
        RECT 138.320 156.660 141.295 156.800 ;
        RECT 120.290 156.320 121.440 156.460 ;
        RECT 113.390 156.260 113.710 156.320 ;
        RECT 116.625 156.275 116.915 156.320 ;
        RECT 120.290 156.260 120.610 156.320 ;
        RECT 41.645 156.120 41.935 156.165 ;
        RECT 40.340 155.980 41.935 156.120 ;
        RECT 41.170 155.920 41.490 155.980 ;
        RECT 41.645 155.935 41.935 155.980 ;
        RECT 42.565 155.935 42.855 156.165 ;
        RECT 44.390 155.920 44.710 156.180 ;
        RECT 48.085 156.120 48.375 156.165 ;
        RECT 48.530 156.120 48.850 156.180 ;
        RECT 48.085 155.980 48.850 156.120 ;
        RECT 48.085 155.935 48.375 155.980 ;
        RECT 48.530 155.920 48.850 155.980 ;
        RECT 57.270 155.920 57.590 156.180 ;
        RECT 58.665 156.120 58.955 156.165 ;
        RECT 61.870 156.120 62.190 156.180 ;
        RECT 58.665 155.980 62.190 156.120 ;
        RECT 58.665 155.935 58.955 155.980 ;
        RECT 61.870 155.920 62.190 155.980 ;
        RECT 68.310 156.120 68.630 156.180 ;
        RECT 71.070 156.165 71.390 156.180 ;
        RECT 68.785 156.120 69.075 156.165 ;
        RECT 69.705 156.120 69.995 156.165 ;
        RECT 71.040 156.120 71.390 156.165 ;
        RECT 68.310 155.980 69.995 156.120 ;
        RECT 70.875 155.980 71.390 156.120 ;
        RECT 68.310 155.920 68.630 155.980 ;
        RECT 68.785 155.935 69.075 155.980 ;
        RECT 69.705 155.935 69.995 155.980 ;
        RECT 71.040 155.935 71.390 155.980 ;
        RECT 71.070 155.920 71.390 155.935 ;
        RECT 87.630 155.920 87.950 156.180 ;
        RECT 89.945 156.120 90.235 156.165 ;
        RECT 94.070 156.120 94.390 156.180 ;
        RECT 89.945 155.980 94.390 156.120 ;
        RECT 89.945 155.935 90.235 155.980 ;
        RECT 94.070 155.920 94.390 155.980 ;
        RECT 101.430 156.120 101.750 156.180 ;
        RECT 105.170 156.120 105.460 156.165 ;
        RECT 101.430 155.980 105.460 156.120 ;
        RECT 101.430 155.920 101.750 155.980 ;
        RECT 105.170 155.935 105.460 155.980 ;
        RECT 108.345 155.935 108.635 156.165 ;
        RECT 109.250 156.120 109.570 156.180 ;
        RECT 118.005 156.120 118.295 156.165 ;
        RECT 109.250 155.980 118.295 156.120 ;
        RECT 47.610 155.780 47.930 155.840 ;
        RECT 49.310 155.780 49.600 155.825 ;
        RECT 62.330 155.780 62.650 155.840 ;
        RECT 47.610 155.640 49.600 155.780 ;
        RECT 47.610 155.580 47.930 155.640 ;
        RECT 49.310 155.595 49.600 155.640 ;
        RECT 50.000 155.640 62.650 155.780 ;
        RECT 50.000 155.440 50.140 155.640 ;
        RECT 62.330 155.580 62.650 155.640 ;
        RECT 65.090 155.780 65.410 155.840 ;
        RECT 67.450 155.780 67.740 155.825 ;
        RECT 92.550 155.780 92.840 155.825 ;
        RECT 65.090 155.640 67.740 155.780 ;
        RECT 65.090 155.580 65.410 155.640 ;
        RECT 67.450 155.595 67.740 155.640 ;
        RECT 90.940 155.640 92.840 155.780 ;
        RECT 108.420 155.780 108.560 155.935 ;
        RECT 109.250 155.920 109.570 155.980 ;
        RECT 118.005 155.935 118.295 155.980 ;
        RECT 111.550 155.780 111.870 155.840 ;
        RECT 116.150 155.780 116.470 155.840 ;
        RECT 108.420 155.640 116.470 155.780 ;
        RECT 118.080 155.780 118.220 155.935 ;
        RECT 118.450 155.920 118.770 156.180 ;
        RECT 119.845 156.120 120.135 156.165 ;
        RECT 120.750 156.120 121.070 156.180 ;
        RECT 119.845 155.980 121.070 156.120 ;
        RECT 121.300 156.120 121.440 156.320 ;
        RECT 121.685 156.275 121.975 156.505 ;
        RECT 124.445 156.460 124.735 156.505 ;
        RECT 124.445 156.320 127.880 156.460 ;
        RECT 124.445 156.275 124.735 156.320 ;
        RECT 125.350 156.120 125.670 156.180 ;
        RECT 121.300 155.980 125.670 156.120 ;
        RECT 119.845 155.935 120.135 155.980 ;
        RECT 120.750 155.920 121.070 155.980 ;
        RECT 125.350 155.920 125.670 155.980 ;
        RECT 125.825 156.120 126.115 156.165 ;
        RECT 127.190 156.120 127.510 156.180 ;
        RECT 127.740 156.165 127.880 156.320 ;
        RECT 128.570 156.260 128.890 156.520 ;
        RECT 132.250 156.460 132.570 156.520 ;
        RECT 129.120 156.320 132.570 156.460 ;
        RECT 125.825 155.980 127.510 156.120 ;
        RECT 125.825 155.935 126.115 155.980 ;
        RECT 118.080 155.640 118.680 155.780 ;
        RECT 38.870 155.300 50.140 155.440 ;
        RECT 57.745 155.440 58.035 155.485 ;
        RECT 59.570 155.440 59.890 155.500 ;
        RECT 83.030 155.440 83.350 155.500 ;
        RECT 90.940 155.485 91.080 155.640 ;
        RECT 92.550 155.595 92.840 155.640 ;
        RECT 111.550 155.580 111.870 155.640 ;
        RECT 116.150 155.580 116.470 155.640 ;
        RECT 57.745 155.300 83.350 155.440 ;
        RECT 29.210 155.240 29.530 155.255 ;
        RECT 32.430 155.240 32.750 155.300 ;
        RECT 38.870 155.240 39.190 155.300 ;
        RECT 57.745 155.255 58.035 155.300 ;
        RECT 59.570 155.240 59.890 155.300 ;
        RECT 83.030 155.240 83.350 155.300 ;
        RECT 90.865 155.255 91.155 155.485 ;
        RECT 96.370 155.440 96.690 155.500 ;
        RECT 98.225 155.440 98.515 155.485 ;
        RECT 96.370 155.300 98.515 155.440 ;
        RECT 96.370 155.240 96.690 155.300 ;
        RECT 98.225 155.255 98.515 155.300 ;
        RECT 110.170 155.440 110.490 155.500 ;
        RECT 113.405 155.440 113.695 155.485 ;
        RECT 110.170 155.300 113.695 155.440 ;
        RECT 110.170 155.240 110.490 155.300 ;
        RECT 113.405 155.255 113.695 155.300 ;
        RECT 117.070 155.240 117.390 155.500 ;
        RECT 118.540 155.440 118.680 155.640 ;
        RECT 118.910 155.580 119.230 155.840 ;
        RECT 122.130 155.780 122.450 155.840 ;
        RECT 125.900 155.780 126.040 155.935 ;
        RECT 127.190 155.920 127.510 155.980 ;
        RECT 127.665 155.935 127.955 156.165 ;
        RECT 128.110 156.120 128.430 156.180 ;
        RECT 129.120 156.120 129.260 156.320 ;
        RECT 132.250 156.260 132.570 156.320 ;
        RECT 128.110 155.980 129.260 156.120 ;
        RECT 128.110 155.920 128.430 155.980 ;
        RECT 129.490 155.920 129.810 156.180 ;
        RECT 129.950 155.920 130.270 156.180 ;
        RECT 130.885 156.120 131.175 156.165 ;
        RECT 131.345 156.120 131.635 156.165 ;
        RECT 130.885 155.980 131.635 156.120 ;
        RECT 130.885 155.935 131.175 155.980 ;
        RECT 131.345 155.935 131.635 155.980 ;
        RECT 131.790 155.920 132.110 156.180 ;
        RECT 132.710 155.920 133.030 156.180 ;
        RECT 133.630 156.120 133.950 156.180 ;
        RECT 138.320 156.165 138.460 156.660 ;
        RECT 141.005 156.615 141.295 156.660 ;
        RECT 143.750 156.800 144.040 156.845 ;
        RECT 145.320 156.800 145.610 156.845 ;
        RECT 147.420 156.800 147.710 156.845 ;
        RECT 143.750 156.660 147.710 156.800 ;
        RECT 143.750 156.615 144.040 156.660 ;
        RECT 145.320 156.615 145.610 156.660 ;
        RECT 147.420 156.615 147.710 156.660 ;
        RECT 143.315 156.460 143.605 156.505 ;
        RECT 145.835 156.460 146.125 156.505 ;
        RECT 147.025 156.460 147.315 156.505 ;
        RECT 143.315 156.320 147.315 156.460 ;
        RECT 143.315 156.275 143.605 156.320 ;
        RECT 145.835 156.275 146.125 156.320 ;
        RECT 147.025 156.275 147.315 156.320 ;
        RECT 135.025 156.120 135.315 156.165 ;
        RECT 137.325 156.120 137.615 156.165 ;
        RECT 133.630 155.980 137.615 156.120 ;
        RECT 133.630 155.920 133.950 155.980 ;
        RECT 135.025 155.935 135.315 155.980 ;
        RECT 137.325 155.935 137.615 155.980 ;
        RECT 138.245 155.935 138.535 156.165 ;
        RECT 138.690 156.120 139.010 156.180 ;
        RECT 139.625 156.120 139.915 156.165 ;
        RECT 138.690 155.980 139.915 156.120 ;
        RECT 119.460 155.640 126.040 155.780 ;
        RECT 119.460 155.440 119.600 155.640 ;
        RECT 122.130 155.580 122.450 155.640 ;
        RECT 126.270 155.580 126.590 155.840 ;
        RECT 126.745 155.780 127.035 155.825 ;
        RECT 134.090 155.780 134.410 155.840 ;
        RECT 135.930 155.780 136.250 155.840 ;
        RECT 138.320 155.780 138.460 155.935 ;
        RECT 138.690 155.920 139.010 155.980 ;
        RECT 139.625 155.935 139.915 155.980 ;
        RECT 147.905 155.935 148.195 156.165 ;
        RECT 149.270 156.120 149.590 156.180 ;
        RECT 149.745 156.120 150.035 156.165 ;
        RECT 149.270 155.980 150.035 156.120 ;
        RECT 146.570 155.780 146.860 155.825 ;
        RECT 126.745 155.640 127.880 155.780 ;
        RECT 126.745 155.595 127.035 155.640 ;
        RECT 127.740 155.500 127.880 155.640 ;
        RECT 134.090 155.640 138.460 155.780 ;
        RECT 140.620 155.640 146.860 155.780 ;
        RECT 147.980 155.780 148.120 155.935 ;
        RECT 149.270 155.920 149.590 155.980 ;
        RECT 149.745 155.935 150.035 155.980 ;
        RECT 153.885 155.780 154.175 155.825 ;
        RECT 155.250 155.780 155.570 155.840 ;
        RECT 147.980 155.640 155.570 155.780 ;
        RECT 134.090 155.580 134.410 155.640 ;
        RECT 135.930 155.580 136.250 155.640 ;
        RECT 118.540 155.300 119.600 155.440 ;
        RECT 124.890 155.240 125.210 155.500 ;
        RECT 125.350 155.440 125.670 155.500 ;
        RECT 127.650 155.440 127.970 155.500 ;
        RECT 125.350 155.300 127.970 155.440 ;
        RECT 125.350 155.240 125.670 155.300 ;
        RECT 127.650 155.240 127.970 155.300 ;
        RECT 133.630 155.240 133.950 155.500 ;
        RECT 137.770 155.240 138.090 155.500 ;
        RECT 140.620 155.485 140.760 155.640 ;
        RECT 146.570 155.595 146.860 155.640 ;
        RECT 153.885 155.595 154.175 155.640 ;
        RECT 155.250 155.580 155.570 155.640 ;
        RECT 140.545 155.255 140.835 155.485 ;
        RECT 22.700 154.620 157.820 155.100 ;
        RECT 31.050 154.220 31.370 154.480 ;
        RECT 31.510 154.220 31.830 154.480 ;
        RECT 40.725 154.420 41.015 154.465 ;
        RECT 42.090 154.420 42.410 154.480 ;
        RECT 40.725 154.280 42.410 154.420 ;
        RECT 40.725 154.235 41.015 154.280 ;
        RECT 42.090 154.220 42.410 154.280 ;
        RECT 65.090 154.220 65.410 154.480 ;
        RECT 74.750 154.420 75.070 154.480 ;
        RECT 82.570 154.420 82.890 154.480 ;
        RECT 68.940 154.280 82.890 154.420 ;
        RECT 31.140 154.080 31.280 154.220 ;
        RECT 32.445 154.080 32.735 154.125 ;
        RECT 38.410 154.080 38.730 154.140 ;
        RECT 39.345 154.080 39.635 154.125 ;
        RECT 31.140 153.940 36.800 154.080 ;
        RECT 32.445 153.895 32.735 153.940 ;
        RECT 36.660 153.800 36.800 153.940 ;
        RECT 38.410 153.940 39.635 154.080 ;
        RECT 38.410 153.880 38.730 153.940 ;
        RECT 39.345 153.895 39.635 153.940 ;
        RECT 25.530 153.785 25.850 153.800 ;
        RECT 25.500 153.555 25.850 153.785 ;
        RECT 25.530 153.540 25.850 153.555 ;
        RECT 30.130 153.740 30.450 153.800 ;
        RECT 33.350 153.740 33.670 153.800 ;
        RECT 30.130 153.600 33.670 153.740 ;
        RECT 30.130 153.540 30.450 153.600 ;
        RECT 33.350 153.540 33.670 153.600 ;
        RECT 33.810 153.540 34.130 153.800 ;
        RECT 36.570 153.540 36.890 153.800 ;
        RECT 37.045 153.740 37.335 153.785 ;
        RECT 37.965 153.740 38.255 153.785 ;
        RECT 37.045 153.600 38.255 153.740 ;
        RECT 37.045 153.555 37.335 153.600 ;
        RECT 37.965 153.555 38.255 153.600 ;
        RECT 38.870 153.540 39.190 153.800 ;
        RECT 39.805 153.740 40.095 153.785 ;
        RECT 42.180 153.740 42.320 154.220 ;
        RECT 63.265 154.080 63.555 154.125 ;
        RECT 68.940 154.080 69.080 154.280 ;
        RECT 74.750 154.220 75.070 154.280 ;
        RECT 82.570 154.220 82.890 154.280 ;
        RECT 94.070 154.220 94.390 154.480 ;
        RECT 95.005 154.420 95.295 154.465 ;
        RECT 96.830 154.420 97.150 154.480 ;
        RECT 98.210 154.420 98.530 154.480 ;
        RECT 98.765 154.420 99.055 154.465 ;
        RECT 95.005 154.280 98.530 154.420 ;
        RECT 95.005 154.235 95.295 154.280 ;
        RECT 96.830 154.220 97.150 154.280 ;
        RECT 98.210 154.220 98.530 154.280 ;
        RECT 98.760 154.235 99.055 154.420 ;
        RECT 82.110 154.080 82.430 154.140 ;
        RECT 63.265 153.940 69.080 154.080 ;
        RECT 69.320 153.940 82.430 154.080 ;
        RECT 63.265 153.895 63.555 153.940 ;
        RECT 69.320 153.800 69.460 153.940 ;
        RECT 43.025 153.740 43.315 153.785 ;
        RECT 39.805 153.600 41.860 153.740 ;
        RECT 42.180 153.600 43.315 153.740 ;
        RECT 39.805 153.555 40.095 153.600 ;
        RECT 24.150 153.200 24.470 153.460 ;
        RECT 25.045 153.400 25.335 153.445 ;
        RECT 26.235 153.400 26.525 153.445 ;
        RECT 28.755 153.400 29.045 153.445 ;
        RECT 25.045 153.260 29.045 153.400 ;
        RECT 25.045 153.215 25.335 153.260 ;
        RECT 26.235 153.215 26.525 153.260 ;
        RECT 28.755 153.215 29.045 153.260 ;
        RECT 24.650 153.060 24.940 153.105 ;
        RECT 26.750 153.060 27.040 153.105 ;
        RECT 28.320 153.060 28.610 153.105 ;
        RECT 24.650 152.920 28.610 153.060 ;
        RECT 24.650 152.875 24.940 152.920 ;
        RECT 26.750 152.875 27.040 152.920 ;
        RECT 28.320 152.875 28.610 152.920 ;
        RECT 41.170 153.060 41.490 153.120 ;
        RECT 41.720 153.060 41.860 153.600 ;
        RECT 43.025 153.555 43.315 153.600 ;
        RECT 43.470 153.540 43.790 153.800 ;
        RECT 44.865 153.740 45.155 153.785 ;
        RECT 45.310 153.740 45.630 153.800 ;
        RECT 44.865 153.600 45.630 153.740 ;
        RECT 44.865 153.555 45.155 153.600 ;
        RECT 45.310 153.540 45.630 153.600 ;
        RECT 50.800 153.740 51.090 153.785 ;
        RECT 53.590 153.740 53.910 153.800 ;
        RECT 50.800 153.600 53.910 153.740 ;
        RECT 50.800 153.555 51.090 153.600 ;
        RECT 53.590 153.540 53.910 153.600 ;
        RECT 57.270 153.740 57.590 153.800 ;
        RECT 62.805 153.740 63.095 153.785 ;
        RECT 57.270 153.600 63.095 153.740 ;
        RECT 57.270 153.540 57.590 153.600 ;
        RECT 62.805 153.555 63.095 153.600 ;
        RECT 42.090 153.400 42.410 153.460 ;
        RECT 44.390 153.400 44.710 153.460 ;
        RECT 42.090 153.260 44.710 153.400 ;
        RECT 42.090 153.200 42.410 153.260 ;
        RECT 44.390 153.200 44.710 153.260 ;
        RECT 48.530 153.400 48.850 153.460 ;
        RECT 49.465 153.400 49.755 153.445 ;
        RECT 48.530 153.260 49.755 153.400 ;
        RECT 48.530 153.200 48.850 153.260 ;
        RECT 49.465 153.215 49.755 153.260 ;
        RECT 50.345 153.400 50.635 153.445 ;
        RECT 51.535 153.400 51.825 153.445 ;
        RECT 54.055 153.400 54.345 153.445 ;
        RECT 58.665 153.400 58.955 153.445 ;
        RECT 50.345 153.260 54.345 153.400 ;
        RECT 50.345 153.215 50.635 153.260 ;
        RECT 51.535 153.215 51.825 153.260 ;
        RECT 54.055 153.215 54.345 153.260 ;
        RECT 56.440 153.260 58.955 153.400 ;
        RECT 62.880 153.400 63.020 153.555 ;
        RECT 64.170 153.540 64.490 153.800 ;
        RECT 67.405 153.555 67.695 153.785 ;
        RECT 68.325 153.740 68.615 153.785 ;
        RECT 69.230 153.740 69.550 153.800 ;
        RECT 68.325 153.600 69.550 153.740 ;
        RECT 68.325 153.555 68.615 153.600 ;
        RECT 66.485 153.400 66.775 153.445 ;
        RECT 62.880 153.260 66.775 153.400 ;
        RECT 67.480 153.400 67.620 153.555 ;
        RECT 69.230 153.540 69.550 153.600 ;
        RECT 76.605 153.740 76.895 153.785 ;
        RECT 77.050 153.740 77.370 153.800 ;
        RECT 78.980 153.785 79.120 153.940 ;
        RECT 82.110 153.880 82.430 153.940 ;
        RECT 83.425 154.080 83.715 154.125 ;
        RECT 83.950 154.080 84.270 154.140 ;
        RECT 83.425 153.940 84.270 154.080 ;
        RECT 83.425 153.895 83.715 153.940 ;
        RECT 83.950 153.880 84.270 153.940 ;
        RECT 84.425 154.080 84.715 154.125 ;
        RECT 84.885 154.080 85.175 154.125 ;
        RECT 84.425 153.940 85.175 154.080 ;
        RECT 84.425 153.895 84.715 153.940 ;
        RECT 84.885 153.895 85.175 153.940 ;
        RECT 96.370 154.080 96.690 154.140 ;
        RECT 97.765 154.080 98.055 154.125 ;
        RECT 98.760 154.080 98.900 154.235 ;
        RECT 113.390 154.220 113.710 154.480 ;
        RECT 118.910 154.420 119.230 154.480 ;
        RECT 125.350 154.420 125.670 154.480 ;
        RECT 128.110 154.420 128.430 154.480 ;
        RECT 118.910 154.280 125.670 154.420 ;
        RECT 118.910 154.220 119.230 154.280 ;
        RECT 125.350 154.220 125.670 154.280 ;
        RECT 126.360 154.280 128.430 154.420 ;
        RECT 109.710 154.080 110.030 154.140 ;
        RECT 117.040 154.080 117.330 154.125 ;
        RECT 124.890 154.080 125.210 154.140 ;
        RECT 96.370 153.940 98.055 154.080 ;
        RECT 96.370 153.880 96.690 153.940 ;
        RECT 97.765 153.895 98.055 153.940 ;
        RECT 98.300 153.940 98.900 154.080 ;
        RECT 106.580 153.940 115.000 154.080 ;
        RECT 98.300 153.800 98.440 153.940 ;
        RECT 76.605 153.600 77.370 153.740 ;
        RECT 76.605 153.555 76.895 153.600 ;
        RECT 77.050 153.540 77.370 153.600 ;
        RECT 78.905 153.555 79.195 153.785 ;
        RECT 80.285 153.740 80.575 153.785 ;
        RECT 81.650 153.740 81.970 153.800 ;
        RECT 89.485 153.740 89.775 153.785 ;
        RECT 80.285 153.600 88.780 153.740 ;
        RECT 80.285 153.555 80.575 153.600 ;
        RECT 81.650 153.540 81.970 153.600 ;
        RECT 70.150 153.400 70.470 153.460 ;
        RECT 74.290 153.400 74.610 153.460 ;
        RECT 67.480 153.260 74.610 153.400 ;
        RECT 56.440 153.105 56.580 153.260 ;
        RECT 58.665 153.215 58.955 153.260 ;
        RECT 66.485 153.215 66.775 153.260 ;
        RECT 70.150 153.200 70.470 153.260 ;
        RECT 74.290 153.200 74.610 153.260 ;
        RECT 75.685 153.215 75.975 153.445 ;
        RECT 76.145 153.400 76.435 153.445 ;
        RECT 83.490 153.400 83.810 153.460 ;
        RECT 76.145 153.260 83.810 153.400 ;
        RECT 76.145 153.215 76.435 153.260 ;
        RECT 49.950 153.060 50.240 153.105 ;
        RECT 52.050 153.060 52.340 153.105 ;
        RECT 53.620 153.060 53.910 153.105 ;
        RECT 41.170 152.920 48.760 153.060 ;
        RECT 41.170 152.860 41.490 152.920 ;
        RECT 34.730 152.520 35.050 152.780 ;
        RECT 45.325 152.720 45.615 152.765 ;
        RECT 48.070 152.720 48.390 152.780 ;
        RECT 45.325 152.580 48.390 152.720 ;
        RECT 48.620 152.720 48.760 152.920 ;
        RECT 49.950 152.920 53.910 153.060 ;
        RECT 49.950 152.875 50.240 152.920 ;
        RECT 52.050 152.875 52.340 152.920 ;
        RECT 53.620 152.875 53.910 152.920 ;
        RECT 56.365 152.875 56.655 153.105 ;
        RECT 75.760 153.060 75.900 153.215 ;
        RECT 83.490 153.200 83.810 153.260 ;
        RECT 84.410 153.400 84.730 153.460 ;
        RECT 87.645 153.400 87.935 153.445 ;
        RECT 88.090 153.400 88.410 153.460 ;
        RECT 84.410 153.260 88.410 153.400 ;
        RECT 84.410 153.200 84.730 153.260 ;
        RECT 87.645 153.215 87.935 153.260 ;
        RECT 88.090 153.200 88.410 153.260 ;
        RECT 80.270 153.060 80.590 153.120 ;
        RECT 75.760 152.920 80.590 153.060 ;
        RECT 88.640 153.060 88.780 153.600 ;
        RECT 89.485 153.600 93.380 153.740 ;
        RECT 89.485 153.555 89.775 153.600 ;
        RECT 93.240 153.460 93.380 153.600 ;
        RECT 98.210 153.540 98.530 153.800 ;
        RECT 98.670 153.740 98.990 153.800 ;
        RECT 106.580 153.785 106.720 153.940 ;
        RECT 109.710 153.880 110.030 153.940 ;
        RECT 107.870 153.785 108.190 153.800 ;
        RECT 100.985 153.740 101.275 153.785 ;
        RECT 98.670 153.600 101.275 153.740 ;
        RECT 98.670 153.540 98.990 153.600 ;
        RECT 100.985 153.555 101.275 153.600 ;
        RECT 106.505 153.555 106.795 153.785 ;
        RECT 107.840 153.555 108.190 153.785 ;
        RECT 107.870 153.540 108.190 153.555 ;
        RECT 114.860 153.460 115.000 153.940 ;
        RECT 117.040 153.940 125.210 154.080 ;
        RECT 117.040 153.895 117.330 153.940 ;
        RECT 124.890 153.880 125.210 153.940 ;
        RECT 126.360 153.785 126.500 154.280 ;
        RECT 128.110 154.220 128.430 154.280 ;
        RECT 129.045 154.420 129.335 154.465 ;
        RECT 132.710 154.420 133.030 154.480 ;
        RECT 135.930 154.420 136.250 154.480 ;
        RECT 129.045 154.280 133.030 154.420 ;
        RECT 129.045 154.235 129.335 154.280 ;
        RECT 132.710 154.220 133.030 154.280 ;
        RECT 134.180 154.280 136.250 154.420 ;
        RECT 127.205 154.080 127.495 154.125 ;
        RECT 128.570 154.080 128.890 154.140 ;
        RECT 131.790 154.080 132.110 154.140 ;
        RECT 133.170 154.125 133.490 154.140 ;
        RECT 127.205 153.940 128.890 154.080 ;
        RECT 127.205 153.895 127.495 153.940 ;
        RECT 126.285 153.555 126.575 153.785 ;
        RECT 93.150 153.200 93.470 153.460 ;
        RECT 102.350 153.400 102.670 153.460 ;
        RECT 93.700 153.260 102.670 153.400 ;
        RECT 93.700 153.060 93.840 153.260 ;
        RECT 102.350 153.200 102.670 153.260 ;
        RECT 107.385 153.400 107.675 153.445 ;
        RECT 108.575 153.400 108.865 153.445 ;
        RECT 111.095 153.400 111.385 153.445 ;
        RECT 107.385 153.260 111.385 153.400 ;
        RECT 107.385 153.215 107.675 153.260 ;
        RECT 108.575 153.215 108.865 153.260 ;
        RECT 111.095 153.215 111.385 153.260 ;
        RECT 114.770 153.400 115.090 153.460 ;
        RECT 115.705 153.400 115.995 153.445 ;
        RECT 114.770 153.260 115.995 153.400 ;
        RECT 114.770 153.200 115.090 153.260 ;
        RECT 115.705 153.215 115.995 153.260 ;
        RECT 116.585 153.400 116.875 153.445 ;
        RECT 117.775 153.400 118.065 153.445 ;
        RECT 120.295 153.400 120.585 153.445 ;
        RECT 116.585 153.260 120.585 153.400 ;
        RECT 116.585 153.215 116.875 153.260 ;
        RECT 117.775 153.215 118.065 153.260 ;
        RECT 120.295 153.215 120.585 153.260 ;
        RECT 88.640 152.920 93.840 153.060 ;
        RECT 96.845 153.060 97.135 153.105 ;
        RECT 106.990 153.060 107.280 153.105 ;
        RECT 109.090 153.060 109.380 153.105 ;
        RECT 110.660 153.060 110.950 153.105 ;
        RECT 96.845 152.920 99.360 153.060 ;
        RECT 56.440 152.720 56.580 152.875 ;
        RECT 80.270 152.860 80.590 152.920 ;
        RECT 96.845 152.875 97.135 152.920 ;
        RECT 99.220 152.780 99.360 152.920 ;
        RECT 106.990 152.920 110.950 153.060 ;
        RECT 106.990 152.875 107.280 152.920 ;
        RECT 109.090 152.875 109.380 152.920 ;
        RECT 110.660 152.875 110.950 152.920 ;
        RECT 116.190 153.060 116.480 153.105 ;
        RECT 118.290 153.060 118.580 153.105 ;
        RECT 119.860 153.060 120.150 153.105 ;
        RECT 116.190 152.920 120.150 153.060 ;
        RECT 116.190 152.875 116.480 152.920 ;
        RECT 118.290 152.875 118.580 152.920 ;
        RECT 119.860 152.875 120.150 152.920 ;
        RECT 122.605 153.060 122.895 153.105 ;
        RECT 127.280 153.060 127.420 153.895 ;
        RECT 128.570 153.880 128.890 153.940 ;
        RECT 131.420 153.940 132.940 154.080 ;
        RECT 127.665 153.555 127.955 153.785 ;
        RECT 128.125 153.740 128.415 153.785 ;
        RECT 130.410 153.740 130.730 153.800 ;
        RECT 131.420 153.785 131.560 153.940 ;
        RECT 131.790 153.880 132.110 153.940 ;
        RECT 128.125 153.600 130.730 153.740 ;
        RECT 128.125 153.555 128.415 153.600 ;
        RECT 127.740 153.400 127.880 153.555 ;
        RECT 130.410 153.540 130.730 153.600 ;
        RECT 131.345 153.555 131.635 153.785 ;
        RECT 132.265 153.555 132.555 153.785 ;
        RECT 132.800 153.740 132.940 153.940 ;
        RECT 133.170 153.895 133.775 154.125 ;
        RECT 133.170 153.880 133.490 153.895 ;
        RECT 134.180 153.740 134.320 154.280 ;
        RECT 135.930 154.220 136.250 154.280 ;
        RECT 137.785 154.235 138.075 154.465 ;
        RECT 140.545 154.235 140.835 154.465 ;
        RECT 134.565 153.895 134.855 154.125 ;
        RECT 132.800 153.600 134.320 153.740 ;
        RECT 134.640 153.740 134.780 153.895 ;
        RECT 136.850 153.880 137.170 154.140 ;
        RECT 137.860 154.080 138.000 154.235 ;
        RECT 140.620 154.080 140.760 154.235 ;
        RECT 146.570 154.080 146.860 154.125 ;
        RECT 137.860 153.940 139.840 154.080 ;
        RECT 140.620 153.940 146.860 154.080 ;
        RECT 139.700 153.785 139.840 153.940 ;
        RECT 146.570 153.895 146.860 153.940 ;
        RECT 139.165 153.740 139.455 153.785 ;
        RECT 134.640 153.600 139.455 153.740 ;
        RECT 139.165 153.555 139.455 153.600 ;
        RECT 139.625 153.555 139.915 153.785 ;
        RECT 131.420 153.400 131.560 153.555 ;
        RECT 127.740 153.260 131.560 153.400 ;
        RECT 132.340 153.400 132.480 153.555 ;
        RECT 137.770 153.400 138.090 153.460 ;
        RECT 132.340 153.260 138.090 153.400 ;
        RECT 137.770 153.200 138.090 153.260 ;
        RECT 122.605 152.920 127.420 153.060 ;
        RECT 131.805 153.060 132.095 153.105 ;
        RECT 131.805 152.920 134.780 153.060 ;
        RECT 122.605 152.875 122.895 152.920 ;
        RECT 131.805 152.875 132.095 152.920 ;
        RECT 48.620 152.580 56.580 152.720 ;
        RECT 45.325 152.535 45.615 152.580 ;
        RECT 48.070 152.520 48.390 152.580 ;
        RECT 61.870 152.520 62.190 152.780 ;
        RECT 78.430 152.520 78.750 152.780 ;
        RECT 82.110 152.720 82.430 152.780 ;
        RECT 82.585 152.720 82.875 152.765 ;
        RECT 82.110 152.580 82.875 152.720 ;
        RECT 82.110 152.520 82.430 152.580 ;
        RECT 82.585 152.535 82.875 152.580 ;
        RECT 83.505 152.720 83.795 152.765 ;
        RECT 85.790 152.720 86.110 152.780 ;
        RECT 83.505 152.580 86.110 152.720 ;
        RECT 83.505 152.535 83.795 152.580 ;
        RECT 85.790 152.520 86.110 152.580 ;
        RECT 89.010 152.520 89.330 152.780 ;
        RECT 89.945 152.720 90.235 152.765 ;
        RECT 90.390 152.720 90.710 152.780 ;
        RECT 89.945 152.580 90.710 152.720 ;
        RECT 89.945 152.535 90.235 152.580 ;
        RECT 90.390 152.520 90.710 152.580 ;
        RECT 94.990 152.520 95.310 152.780 ;
        RECT 98.670 152.520 98.990 152.780 ;
        RECT 99.130 152.720 99.450 152.780 ;
        RECT 99.605 152.720 99.895 152.765 ;
        RECT 99.130 152.580 99.895 152.720 ;
        RECT 99.130 152.520 99.450 152.580 ;
        RECT 99.605 152.535 99.895 152.580 ;
        RECT 104.190 152.520 104.510 152.780 ;
        RECT 132.725 152.720 133.015 152.765 ;
        RECT 133.170 152.720 133.490 152.780 ;
        RECT 132.725 152.580 133.490 152.720 ;
        RECT 132.725 152.535 133.015 152.580 ;
        RECT 133.170 152.520 133.490 152.580 ;
        RECT 133.645 152.720 133.935 152.765 ;
        RECT 134.090 152.720 134.410 152.780 ;
        RECT 133.645 152.580 134.410 152.720 ;
        RECT 134.640 152.720 134.780 152.920 ;
        RECT 135.010 152.860 135.330 153.120 ;
        RECT 135.930 153.060 136.250 153.120 ;
        RECT 138.705 153.060 138.995 153.105 ;
        RECT 135.930 152.920 138.995 153.060 ;
        RECT 139.240 153.060 139.380 153.555 ;
        RECT 143.315 153.400 143.605 153.445 ;
        RECT 145.835 153.400 146.125 153.445 ;
        RECT 147.025 153.400 147.315 153.445 ;
        RECT 143.315 153.260 147.315 153.400 ;
        RECT 143.315 153.215 143.605 153.260 ;
        RECT 145.835 153.215 146.125 153.260 ;
        RECT 147.025 153.215 147.315 153.260 ;
        RECT 147.905 153.400 148.195 153.445 ;
        RECT 155.250 153.400 155.570 153.460 ;
        RECT 147.905 153.260 155.570 153.400 ;
        RECT 147.905 153.215 148.195 153.260 ;
        RECT 155.250 153.200 155.570 153.260 ;
        RECT 141.005 153.060 141.295 153.105 ;
        RECT 139.240 152.920 141.295 153.060 ;
        RECT 135.930 152.860 136.250 152.920 ;
        RECT 138.705 152.875 138.995 152.920 ;
        RECT 141.005 152.875 141.295 152.920 ;
        RECT 143.750 153.060 144.040 153.105 ;
        RECT 145.320 153.060 145.610 153.105 ;
        RECT 147.420 153.060 147.710 153.105 ;
        RECT 143.750 152.920 147.710 153.060 ;
        RECT 143.750 152.875 144.040 152.920 ;
        RECT 145.320 152.875 145.610 152.920 ;
        RECT 147.420 152.875 147.710 152.920 ;
        RECT 136.865 152.720 137.155 152.765 ;
        RECT 134.640 152.580 137.155 152.720 ;
        RECT 133.645 152.535 133.935 152.580 ;
        RECT 134.090 152.520 134.410 152.580 ;
        RECT 136.865 152.535 137.155 152.580 ;
        RECT 22.700 151.900 157.020 152.380 ;
        RECT 25.085 151.700 25.375 151.745 ;
        RECT 25.530 151.700 25.850 151.760 ;
        RECT 25.085 151.560 25.850 151.700 ;
        RECT 25.085 151.515 25.375 151.560 ;
        RECT 25.530 151.500 25.850 151.560 ;
        RECT 27.370 151.700 27.690 151.760 ;
        RECT 31.985 151.700 32.275 151.745 ;
        RECT 27.370 151.560 32.275 151.700 ;
        RECT 27.370 151.500 27.690 151.560 ;
        RECT 31.985 151.515 32.275 151.560 ;
        RECT 32.905 151.700 33.195 151.745 ;
        RECT 33.810 151.700 34.130 151.760 ;
        RECT 32.905 151.560 34.130 151.700 ;
        RECT 32.905 151.515 33.195 151.560 ;
        RECT 33.810 151.500 34.130 151.560 ;
        RECT 34.285 151.700 34.575 151.745 ;
        RECT 36.570 151.700 36.890 151.760 ;
        RECT 34.285 151.560 36.890 151.700 ;
        RECT 34.285 151.515 34.575 151.560 ;
        RECT 36.570 151.500 36.890 151.560 ;
        RECT 41.170 151.500 41.490 151.760 ;
        RECT 42.090 151.500 42.410 151.760 ;
        RECT 53.590 151.500 53.910 151.760 ;
        RECT 57.285 151.700 57.575 151.745 ;
        RECT 59.585 151.700 59.875 151.745 ;
        RECT 60.490 151.700 60.810 151.760 ;
        RECT 63.725 151.700 64.015 151.745 ;
        RECT 57.285 151.560 64.015 151.700 ;
        RECT 57.285 151.515 57.575 151.560 ;
        RECT 59.585 151.515 59.875 151.560 ;
        RECT 60.490 151.500 60.810 151.560 ;
        RECT 63.725 151.515 64.015 151.560 ;
        RECT 84.410 151.500 84.730 151.760 ;
        RECT 85.790 151.500 86.110 151.760 ;
        RECT 89.010 151.700 89.330 151.760 ;
        RECT 97.305 151.700 97.595 151.745 ;
        RECT 89.010 151.560 97.595 151.700 ;
        RECT 89.010 151.500 89.330 151.560 ;
        RECT 97.305 151.515 97.595 151.560 ;
        RECT 100.970 151.500 101.290 151.760 ;
        RECT 104.665 151.700 104.955 151.745 ;
        RECT 107.870 151.700 108.190 151.760 ;
        RECT 104.665 151.560 108.190 151.700 ;
        RECT 104.665 151.515 104.955 151.560 ;
        RECT 107.870 151.500 108.190 151.560 ;
        RECT 120.750 151.700 121.070 151.760 ;
        RECT 123.065 151.700 123.355 151.745 ;
        RECT 120.750 151.560 123.355 151.700 ;
        RECT 120.750 151.500 121.070 151.560 ;
        RECT 123.065 151.515 123.355 151.560 ;
        RECT 133.170 151.700 133.490 151.760 ;
        RECT 135.010 151.700 135.330 151.760 ;
        RECT 133.170 151.560 135.330 151.700 ;
        RECT 133.170 151.500 133.490 151.560 ;
        RECT 135.010 151.500 135.330 151.560 ;
        RECT 30.130 151.360 30.450 151.420 ;
        RECT 33.365 151.360 33.655 151.405 ;
        RECT 48.990 151.360 49.310 151.420 ;
        RECT 58.665 151.360 58.955 151.405 ;
        RECT 30.130 151.220 33.655 151.360 ;
        RECT 30.130 151.160 30.450 151.220 ;
        RECT 33.365 151.175 33.655 151.220 ;
        RECT 48.620 151.220 49.310 151.360 ;
        RECT 36.585 151.020 36.875 151.065 ;
        RECT 37.950 151.020 38.270 151.080 ;
        RECT 33.670 150.880 38.270 151.020 ;
        RECT 25.990 150.480 26.310 150.740 ;
        RECT 28.765 150.680 29.055 150.725 ;
        RECT 29.210 150.680 29.530 150.740 ;
        RECT 28.765 150.540 29.530 150.680 ;
        RECT 28.765 150.495 29.055 150.540 ;
        RECT 29.210 150.480 29.530 150.540 ;
        RECT 29.685 150.495 29.975 150.725 ;
        RECT 33.670 150.680 33.810 150.880 ;
        RECT 36.585 150.835 36.875 150.880 ;
        RECT 37.950 150.820 38.270 150.880 ;
        RECT 48.070 150.820 48.390 151.080 ;
        RECT 37.045 150.680 37.335 150.725 ;
        RECT 39.805 150.680 40.095 150.725 ;
        RECT 31.600 150.540 33.810 150.680 ;
        RECT 35.280 150.540 40.095 150.680 ;
        RECT 29.760 150.340 29.900 150.495 ;
        RECT 31.600 150.340 31.740 150.540 ;
        RECT 29.760 150.200 31.740 150.340 ;
        RECT 32.430 150.340 32.750 150.400 ;
        RECT 35.280 150.385 35.420 150.540 ;
        RECT 37.045 150.495 37.335 150.540 ;
        RECT 39.805 150.495 40.095 150.540 ;
        RECT 43.010 150.680 43.330 150.740 ;
        RECT 44.405 150.680 44.695 150.725 ;
        RECT 43.010 150.540 44.695 150.680 ;
        RECT 43.010 150.480 43.330 150.540 ;
        RECT 44.405 150.495 44.695 150.540 ;
        RECT 44.865 150.680 45.155 150.725 ;
        RECT 47.625 150.680 47.915 150.725 ;
        RECT 48.620 150.680 48.760 151.220 ;
        RECT 48.990 151.160 49.310 151.220 ;
        RECT 55.060 151.220 58.955 151.360 ;
        RECT 44.865 150.540 47.380 150.680 ;
        RECT 44.865 150.495 45.155 150.540 ;
        RECT 47.240 150.385 47.380 150.540 ;
        RECT 47.625 150.540 48.760 150.680 ;
        RECT 47.625 150.495 47.915 150.540 ;
        RECT 48.990 150.480 49.310 150.740 ;
        RECT 49.465 150.495 49.755 150.725 ;
        RECT 54.525 150.680 54.815 150.725 ;
        RECT 55.060 150.680 55.200 151.220 ;
        RECT 58.665 151.175 58.955 151.220 ;
        RECT 78.010 151.360 78.300 151.405 ;
        RECT 80.110 151.360 80.400 151.405 ;
        RECT 81.680 151.360 81.970 151.405 ;
        RECT 78.010 151.220 81.970 151.360 ;
        RECT 78.010 151.175 78.300 151.220 ;
        RECT 80.110 151.175 80.400 151.220 ;
        RECT 81.680 151.175 81.970 151.220 ;
        RECT 88.130 151.360 88.420 151.405 ;
        RECT 90.230 151.360 90.520 151.405 ;
        RECT 91.800 151.360 92.090 151.405 ;
        RECT 88.130 151.220 92.090 151.360 ;
        RECT 88.130 151.175 88.420 151.220 ;
        RECT 90.230 151.175 90.520 151.220 ;
        RECT 91.800 151.175 92.090 151.220 ;
        RECT 93.150 151.360 93.470 151.420 ;
        RECT 94.545 151.360 94.835 151.405 ;
        RECT 93.150 151.220 94.835 151.360 ;
        RECT 93.150 151.160 93.470 151.220 ;
        RECT 94.545 151.175 94.835 151.220 ;
        RECT 106.490 151.360 106.810 151.420 ;
        RECT 108.790 151.360 109.110 151.420 ;
        RECT 106.490 151.220 109.110 151.360 ;
        RECT 106.490 151.160 106.810 151.220 ;
        RECT 108.790 151.160 109.110 151.220 ;
        RECT 116.190 151.360 116.480 151.405 ;
        RECT 118.290 151.360 118.580 151.405 ;
        RECT 119.860 151.360 120.150 151.405 ;
        RECT 116.190 151.220 120.150 151.360 ;
        RECT 116.190 151.175 116.480 151.220 ;
        RECT 118.290 151.175 118.580 151.220 ;
        RECT 119.860 151.175 120.150 151.220 ;
        RECT 130.410 151.360 130.730 151.420 ;
        RECT 150.650 151.360 150.940 151.405 ;
        RECT 152.220 151.360 152.510 151.405 ;
        RECT 154.320 151.360 154.610 151.405 ;
        RECT 130.410 151.220 132.480 151.360 ;
        RECT 130.410 151.160 130.730 151.220 ;
        RECT 78.405 151.020 78.695 151.065 ;
        RECT 79.595 151.020 79.885 151.065 ;
        RECT 82.115 151.020 82.405 151.065 ;
        RECT 55.520 150.880 56.580 151.020 ;
        RECT 55.520 150.725 55.660 150.880 ;
        RECT 54.525 150.540 55.200 150.680 ;
        RECT 54.525 150.495 54.815 150.540 ;
        RECT 55.445 150.495 55.735 150.725 ;
        RECT 35.205 150.340 35.495 150.385 ;
        RECT 32.430 150.200 35.495 150.340 ;
        RECT 32.430 150.140 32.750 150.200 ;
        RECT 35.205 150.155 35.495 150.200 ;
        RECT 47.165 150.155 47.455 150.385 ;
        RECT 48.070 150.340 48.390 150.400 ;
        RECT 49.540 150.340 49.680 150.495 ;
        RECT 55.890 150.480 56.210 150.740 ;
        RECT 56.440 150.680 56.580 150.880 ;
        RECT 78.405 150.880 82.405 151.020 ;
        RECT 78.405 150.835 78.695 150.880 ;
        RECT 79.595 150.835 79.885 150.880 ;
        RECT 82.115 150.835 82.405 150.880 ;
        RECT 88.525 151.020 88.815 151.065 ;
        RECT 89.715 151.020 90.005 151.065 ;
        RECT 92.235 151.020 92.525 151.065 ;
        RECT 88.525 150.880 92.525 151.020 ;
        RECT 88.525 150.835 88.815 150.880 ;
        RECT 89.715 150.835 90.005 150.880 ;
        RECT 92.235 150.835 92.525 150.880 ;
        RECT 101.905 150.835 102.195 151.065 ;
        RECT 109.250 151.020 109.570 151.080 ;
        RECT 105.660 150.880 109.570 151.020 ;
        RECT 58.650 150.680 58.970 150.740 ;
        RECT 56.440 150.540 58.970 150.680 ;
        RECT 58.650 150.480 58.970 150.540 ;
        RECT 77.510 150.480 77.830 150.740 ;
        RECT 86.710 150.680 87.030 150.740 ;
        RECT 87.645 150.680 87.935 150.725 ;
        RECT 90.390 150.680 90.710 150.740 ;
        RECT 86.710 150.540 87.935 150.680 ;
        RECT 86.710 150.480 87.030 150.540 ;
        RECT 87.645 150.495 87.935 150.540 ;
        RECT 88.180 150.540 90.710 150.680 ;
        RECT 56.365 150.340 56.655 150.385 ;
        RECT 59.425 150.340 59.715 150.385 ;
        RECT 60.505 150.340 60.795 150.385 ;
        RECT 61.870 150.340 62.190 150.400 ;
        RECT 48.070 150.200 49.680 150.340 ;
        RECT 55.520 150.200 56.655 150.340 ;
        RECT 48.070 150.140 48.390 150.200 ;
        RECT 29.685 150.000 29.975 150.045 ;
        RECT 31.985 150.000 32.275 150.045 ;
        RECT 29.685 149.860 32.275 150.000 ;
        RECT 29.685 149.815 29.975 149.860 ;
        RECT 31.985 149.815 32.275 149.860 ;
        RECT 33.350 150.000 33.670 150.060 ;
        RECT 34.155 150.000 34.445 150.045 ;
        RECT 33.350 149.860 34.445 150.000 ;
        RECT 33.350 149.800 33.670 149.860 ;
        RECT 34.155 149.815 34.445 149.860 ;
        RECT 43.010 150.000 43.330 150.060 ;
        RECT 43.485 150.000 43.775 150.045 ;
        RECT 43.010 149.860 43.775 150.000 ;
        RECT 43.010 149.800 43.330 149.860 ;
        RECT 43.485 149.815 43.775 149.860 ;
        RECT 46.705 150.000 46.995 150.045 ;
        RECT 49.450 150.000 49.770 150.060 ;
        RECT 46.705 149.860 49.770 150.000 ;
        RECT 46.705 149.815 46.995 149.860 ;
        RECT 49.450 149.800 49.770 149.860 ;
        RECT 52.210 150.000 52.530 150.060 ;
        RECT 55.520 150.000 55.660 150.200 ;
        RECT 56.365 150.155 56.655 150.200 ;
        RECT 57.440 150.200 59.720 150.340 ;
        RECT 57.440 150.060 57.580 150.200 ;
        RECT 59.425 150.155 59.720 150.200 ;
        RECT 60.505 150.200 62.190 150.340 ;
        RECT 60.505 150.155 60.795 150.200 ;
        RECT 52.210 149.860 55.660 150.000 ;
        RECT 57.270 150.045 57.590 150.060 ;
        RECT 52.210 149.800 52.530 149.860 ;
        RECT 57.270 149.815 57.655 150.045 ;
        RECT 57.270 149.800 57.590 149.815 ;
        RECT 58.190 149.800 58.510 150.060 ;
        RECT 59.580 150.000 59.720 150.155 ;
        RECT 61.870 150.140 62.190 150.200 ;
        RECT 62.790 150.140 63.110 150.400 ;
        RECT 67.390 150.340 67.710 150.400 ;
        RECT 68.770 150.340 69.090 150.400 ;
        RECT 67.390 150.200 69.090 150.340 ;
        RECT 67.390 150.140 67.710 150.200 ;
        RECT 68.770 150.140 69.090 150.200 ;
        RECT 75.210 150.140 75.530 150.400 ;
        RECT 78.860 150.340 79.150 150.385 ;
        RECT 81.190 150.340 81.510 150.400 ;
        RECT 78.860 150.200 81.510 150.340 ;
        RECT 78.860 150.155 79.150 150.200 ;
        RECT 81.190 150.140 81.510 150.200 ;
        RECT 84.885 150.340 85.175 150.385 ;
        RECT 88.180 150.340 88.320 150.540 ;
        RECT 90.390 150.480 90.710 150.540 ;
        RECT 95.910 150.480 96.230 150.740 ;
        RECT 96.370 150.480 96.690 150.740 ;
        RECT 97.765 150.680 98.055 150.725 ;
        RECT 98.670 150.680 98.990 150.740 ;
        RECT 97.765 150.540 98.990 150.680 ;
        RECT 97.765 150.495 98.055 150.540 ;
        RECT 98.670 150.480 98.990 150.540 ;
        RECT 99.130 150.480 99.450 150.740 ;
        RECT 100.065 150.680 100.355 150.725 ;
        RECT 100.510 150.680 100.830 150.740 ;
        RECT 100.065 150.540 100.830 150.680 ;
        RECT 100.065 150.495 100.355 150.540 ;
        RECT 100.510 150.480 100.830 150.540 ;
        RECT 84.885 150.200 88.320 150.340 ;
        RECT 88.870 150.340 89.160 150.385 ;
        RECT 97.290 150.340 97.610 150.400 ;
        RECT 101.980 150.340 102.120 150.835 ;
        RECT 102.365 150.680 102.655 150.725 ;
        RECT 104.190 150.680 104.510 150.740 ;
        RECT 105.660 150.725 105.800 150.880 ;
        RECT 109.250 150.820 109.570 150.880 ;
        RECT 116.585 151.020 116.875 151.065 ;
        RECT 117.775 151.020 118.065 151.065 ;
        RECT 120.295 151.020 120.585 151.065 ;
        RECT 130.885 151.020 131.175 151.065 ;
        RECT 131.330 151.020 131.650 151.080 ;
        RECT 116.585 150.880 120.585 151.020 ;
        RECT 116.585 150.835 116.875 150.880 ;
        RECT 117.775 150.835 118.065 150.880 ;
        RECT 120.295 150.835 120.585 150.880 ;
        RECT 130.040 150.880 131.650 151.020 ;
        RECT 102.365 150.540 104.510 150.680 ;
        RECT 102.365 150.495 102.655 150.540 ;
        RECT 104.190 150.480 104.510 150.540 ;
        RECT 105.585 150.495 105.875 150.725 ;
        RECT 106.490 150.480 106.810 150.740 ;
        RECT 107.425 150.680 107.715 150.725 ;
        RECT 110.170 150.680 110.490 150.740 ;
        RECT 107.425 150.540 110.490 150.680 ;
        RECT 107.425 150.495 107.715 150.540 ;
        RECT 110.170 150.480 110.490 150.540 ;
        RECT 112.025 150.680 112.315 150.725 ;
        RECT 114.770 150.680 115.090 150.740 ;
        RECT 115.705 150.680 115.995 150.725 ;
        RECT 112.025 150.540 115.995 150.680 ;
        RECT 112.025 150.495 112.315 150.540 ;
        RECT 114.770 150.480 115.090 150.540 ;
        RECT 115.705 150.495 115.995 150.540 ;
        RECT 125.810 150.480 126.130 150.740 ;
        RECT 126.745 150.680 127.035 150.725 ;
        RECT 130.040 150.680 130.180 150.880 ;
        RECT 130.885 150.835 131.175 150.880 ;
        RECT 131.330 150.820 131.650 150.880 ;
        RECT 126.745 150.540 130.180 150.680 ;
        RECT 126.745 150.495 127.035 150.540 ;
        RECT 130.425 150.495 130.715 150.725 ;
        RECT 84.885 150.155 85.175 150.200 ;
        RECT 88.870 150.155 89.240 150.340 ;
        RECT 63.710 150.045 64.030 150.060 ;
        RECT 63.710 150.000 64.095 150.045 ;
        RECT 59.580 149.860 64.095 150.000 ;
        RECT 63.710 149.815 64.095 149.860 ;
        RECT 63.710 149.800 64.030 149.815 ;
        RECT 64.630 149.800 64.950 150.060 ;
        RECT 83.950 150.000 84.270 150.060 ;
        RECT 85.885 150.000 86.175 150.045 ;
        RECT 83.950 149.860 86.175 150.000 ;
        RECT 83.950 149.800 84.270 149.860 ;
        RECT 85.885 149.815 86.175 149.860 ;
        RECT 86.710 149.800 87.030 150.060 ;
        RECT 87.630 150.000 87.950 150.060 ;
        RECT 89.100 150.000 89.240 150.155 ;
        RECT 97.290 150.200 102.120 150.340 ;
        RECT 97.290 150.140 97.610 150.200 ;
        RECT 106.030 150.140 106.350 150.400 ;
        RECT 107.870 150.140 108.190 150.400 ;
        RECT 112.470 150.340 112.790 150.400 ;
        RECT 115.230 150.340 115.550 150.400 ;
        RECT 112.470 150.200 115.550 150.340 ;
        RECT 112.470 150.140 112.790 150.200 ;
        RECT 115.230 150.140 115.550 150.200 ;
        RECT 117.040 150.340 117.330 150.385 ;
        RECT 125.350 150.340 125.670 150.400 ;
        RECT 117.040 150.200 125.670 150.340 ;
        RECT 117.040 150.155 117.330 150.200 ;
        RECT 125.350 150.140 125.670 150.200 ;
        RECT 87.630 149.860 89.240 150.000 ;
        RECT 87.630 149.800 87.950 149.860 ;
        RECT 94.990 149.800 95.310 150.060 ;
        RECT 98.225 150.000 98.515 150.045 ;
        RECT 98.670 150.000 98.990 150.060 ;
        RECT 98.225 149.860 98.990 150.000 ;
        RECT 107.960 150.000 108.100 150.140 ;
        RECT 122.130 150.000 122.450 150.060 ;
        RECT 107.960 149.860 122.450 150.000 ;
        RECT 98.225 149.815 98.515 149.860 ;
        RECT 98.670 149.800 98.990 149.860 ;
        RECT 122.130 149.800 122.450 149.860 ;
        RECT 122.605 150.000 122.895 150.045 ;
        RECT 126.820 150.000 126.960 150.495 ;
        RECT 122.605 149.860 126.960 150.000 ;
        RECT 129.030 150.000 129.350 150.060 ;
        RECT 129.965 150.000 130.255 150.045 ;
        RECT 129.030 149.860 130.255 150.000 ;
        RECT 130.500 150.000 130.640 150.495 ;
        RECT 131.790 150.480 132.110 150.740 ;
        RECT 132.340 150.725 132.480 151.220 ;
        RECT 150.650 151.220 154.610 151.360 ;
        RECT 150.650 151.175 150.940 151.220 ;
        RECT 152.220 151.175 152.510 151.220 ;
        RECT 154.320 151.175 154.610 151.220 ;
        RECT 134.090 151.020 134.410 151.080 ;
        RECT 150.215 151.020 150.505 151.065 ;
        RECT 152.735 151.020 153.025 151.065 ;
        RECT 153.925 151.020 154.215 151.065 ;
        RECT 134.090 150.880 135.700 151.020 ;
        RECT 134.090 150.820 134.410 150.880 ;
        RECT 132.265 150.495 132.555 150.725 ;
        RECT 133.630 150.480 133.950 150.740 ;
        RECT 135.010 150.480 135.330 150.740 ;
        RECT 135.560 150.680 135.700 150.880 ;
        RECT 150.215 150.880 154.215 151.020 ;
        RECT 150.215 150.835 150.505 150.880 ;
        RECT 152.735 150.835 153.025 150.880 ;
        RECT 153.925 150.835 154.215 150.880 ;
        RECT 136.390 150.680 136.710 150.740 ;
        RECT 137.785 150.680 138.075 150.725 ;
        RECT 145.590 150.680 145.910 150.740 ;
        RECT 135.560 150.540 145.910 150.680 ;
        RECT 136.390 150.480 136.710 150.540 ;
        RECT 137.785 150.495 138.075 150.540 ;
        RECT 145.590 150.480 145.910 150.540 ;
        RECT 154.805 150.680 155.095 150.725 ;
        RECT 155.250 150.680 155.570 150.740 ;
        RECT 154.805 150.540 155.570 150.680 ;
        RECT 154.805 150.495 155.095 150.540 ;
        RECT 155.250 150.480 155.570 150.540 ;
        RECT 134.550 150.340 134.870 150.400 ;
        RECT 136.850 150.340 137.170 150.400 ;
        RECT 134.550 150.200 137.170 150.340 ;
        RECT 134.550 150.140 134.870 150.200 ;
        RECT 136.850 150.140 137.170 150.200 ;
        RECT 148.810 150.340 149.130 150.400 ;
        RECT 153.470 150.340 153.760 150.385 ;
        RECT 148.810 150.200 153.760 150.340 ;
        RECT 148.810 150.140 149.130 150.200 ;
        RECT 153.470 150.155 153.760 150.200 ;
        RECT 132.250 150.000 132.570 150.060 ;
        RECT 130.500 149.860 132.570 150.000 ;
        RECT 122.605 149.815 122.895 149.860 ;
        RECT 129.030 149.800 129.350 149.860 ;
        RECT 129.965 149.815 130.255 149.860 ;
        RECT 132.250 149.800 132.570 149.860 ;
        RECT 133.185 150.000 133.475 150.045 ;
        RECT 134.105 150.000 134.395 150.045 ;
        RECT 133.185 149.860 134.395 150.000 ;
        RECT 133.185 149.815 133.475 149.860 ;
        RECT 134.105 149.815 134.395 149.860 ;
        RECT 135.945 150.000 136.235 150.045 ;
        RECT 136.390 150.000 136.710 150.060 ;
        RECT 135.945 149.860 136.710 150.000 ;
        RECT 135.945 149.815 136.235 149.860 ;
        RECT 136.390 149.800 136.710 149.860 ;
        RECT 143.750 150.000 144.070 150.060 ;
        RECT 147.905 150.000 148.195 150.045 ;
        RECT 143.750 149.860 148.195 150.000 ;
        RECT 143.750 149.800 144.070 149.860 ;
        RECT 147.905 149.815 148.195 149.860 ;
        RECT 22.700 149.180 157.820 149.660 ;
        RECT 32.430 148.780 32.750 149.040 ;
        RECT 48.990 148.980 49.310 149.040 ;
        RECT 50.385 148.980 50.675 149.025 ;
        RECT 48.990 148.840 50.675 148.980 ;
        RECT 48.990 148.780 49.310 148.840 ;
        RECT 50.385 148.795 50.675 148.840 ;
        RECT 51.750 148.980 52.070 149.040 ;
        RECT 59.585 148.980 59.875 149.025 ;
        RECT 62.790 148.980 63.110 149.040 ;
        RECT 51.750 148.840 63.110 148.980 ;
        RECT 51.750 148.780 52.070 148.840 ;
        RECT 59.585 148.795 59.875 148.840 ;
        RECT 62.790 148.780 63.110 148.840 ;
        RECT 75.210 148.980 75.530 149.040 ;
        RECT 91.785 148.980 92.075 149.025 ;
        RECT 122.130 148.980 122.450 149.040 ;
        RECT 122.605 148.980 122.895 149.025 ;
        RECT 126.270 148.980 126.590 149.040 ;
        RECT 75.210 148.840 116.380 148.980 ;
        RECT 75.210 148.780 75.530 148.840 ;
        RECT 91.785 148.795 92.075 148.840 ;
        RECT 34.730 148.640 35.050 148.700 ;
        RECT 38.010 148.640 38.300 148.685 ;
        RECT 52.670 148.640 52.990 148.700 ;
        RECT 77.510 148.640 77.830 148.700 ;
        RECT 34.730 148.500 38.300 148.640 ;
        RECT 34.730 148.440 35.050 148.500 ;
        RECT 38.010 148.455 38.300 148.500 ;
        RECT 49.080 148.500 52.990 148.640 ;
        RECT 39.345 148.300 39.635 148.345 ;
        RECT 48.530 148.300 48.850 148.360 ;
        RECT 49.080 148.345 49.220 148.500 ;
        RECT 52.670 148.440 52.990 148.500 ;
        RECT 59.200 148.500 77.830 148.640 ;
        RECT 39.345 148.160 48.850 148.300 ;
        RECT 39.345 148.115 39.635 148.160 ;
        RECT 48.530 148.100 48.850 148.160 ;
        RECT 49.005 148.115 49.295 148.345 ;
        RECT 49.910 148.100 50.230 148.360 ;
        RECT 50.370 148.100 50.690 148.360 ;
        RECT 51.305 148.115 51.595 148.345 ;
        RECT 56.350 148.300 56.670 148.360 ;
        RECT 59.200 148.345 59.340 148.500 ;
        RECT 57.790 148.300 58.080 148.345 ;
        RECT 56.350 148.160 58.080 148.300 ;
        RECT 34.755 147.960 35.045 148.005 ;
        RECT 37.275 147.960 37.565 148.005 ;
        RECT 38.465 147.960 38.755 148.005 ;
        RECT 51.380 147.960 51.520 148.115 ;
        RECT 56.350 148.100 56.670 148.160 ;
        RECT 57.790 148.115 58.080 148.160 ;
        RECT 59.125 148.115 59.415 148.345 ;
        RECT 62.790 148.300 63.110 148.360 ;
        RECT 65.150 148.300 65.440 148.345 ;
        RECT 62.790 148.160 65.440 148.300 ;
        RECT 62.790 148.100 63.110 148.160 ;
        RECT 65.150 148.115 65.440 148.160 ;
        RECT 66.560 148.005 66.700 148.500 ;
        RECT 73.920 148.345 74.060 148.500 ;
        RECT 77.510 148.440 77.830 148.500 ;
        RECT 81.190 148.440 81.510 148.700 ;
        RECT 85.805 148.640 86.095 148.685 ;
        RECT 87.170 148.640 87.490 148.700 ;
        RECT 85.805 148.500 87.490 148.640 ;
        RECT 85.805 148.455 86.095 148.500 ;
        RECT 87.170 148.440 87.490 148.500 ;
        RECT 87.630 148.440 87.950 148.700 ;
        RECT 88.565 148.640 88.855 148.685 ;
        RECT 95.910 148.640 96.230 148.700 ;
        RECT 116.240 148.685 116.380 148.840 ;
        RECT 122.130 148.840 126.590 148.980 ;
        RECT 122.130 148.780 122.450 148.840 ;
        RECT 122.605 148.795 122.895 148.840 ;
        RECT 126.270 148.780 126.590 148.840 ;
        RECT 126.730 148.980 127.050 149.040 ;
        RECT 129.505 148.980 129.795 149.025 ;
        RECT 135.010 148.980 135.330 149.040 ;
        RECT 126.730 148.840 127.880 148.980 ;
        RECT 126.730 148.780 127.050 148.840 ;
        RECT 127.740 148.685 127.880 148.840 ;
        RECT 129.505 148.840 135.330 148.980 ;
        RECT 129.505 148.795 129.795 148.840 ;
        RECT 135.010 148.780 135.330 148.840 ;
        RECT 148.810 148.780 149.130 149.040 ;
        RECT 88.565 148.500 96.230 148.640 ;
        RECT 88.565 148.455 88.855 148.500 ;
        RECT 91.860 148.360 92.000 148.500 ;
        RECT 95.910 148.440 96.230 148.500 ;
        RECT 98.225 148.640 98.515 148.685 ;
        RECT 98.225 148.500 114.540 148.640 ;
        RECT 98.225 148.455 98.515 148.500 ;
        RECT 72.565 148.300 72.855 148.345 ;
        RECT 72.565 148.160 73.600 148.300 ;
        RECT 72.565 148.115 72.855 148.160 ;
        RECT 34.755 147.820 38.755 147.960 ;
        RECT 34.755 147.775 35.045 147.820 ;
        RECT 37.275 147.775 37.565 147.820 ;
        RECT 38.465 147.775 38.755 147.820 ;
        RECT 49.540 147.820 51.520 147.960 ;
        RECT 54.535 147.960 54.825 148.005 ;
        RECT 57.055 147.960 57.345 148.005 ;
        RECT 58.245 147.960 58.535 148.005 ;
        RECT 54.535 147.820 58.535 147.960 ;
        RECT 35.190 147.620 35.480 147.665 ;
        RECT 36.760 147.620 37.050 147.665 ;
        RECT 38.860 147.620 39.150 147.665 ;
        RECT 35.190 147.480 39.150 147.620 ;
        RECT 35.190 147.435 35.480 147.480 ;
        RECT 36.760 147.435 37.050 147.480 ;
        RECT 38.860 147.435 39.150 147.480 ;
        RECT 44.850 147.280 45.170 147.340 ;
        RECT 49.540 147.325 49.680 147.820 ;
        RECT 54.535 147.775 54.825 147.820 ;
        RECT 57.055 147.775 57.345 147.820 ;
        RECT 58.245 147.775 58.535 147.820 ;
        RECT 61.895 147.960 62.185 148.005 ;
        RECT 64.415 147.960 64.705 148.005 ;
        RECT 65.605 147.960 65.895 148.005 ;
        RECT 61.895 147.820 65.895 147.960 ;
        RECT 61.895 147.775 62.185 147.820 ;
        RECT 64.415 147.775 64.705 147.820 ;
        RECT 65.605 147.775 65.895 147.820 ;
        RECT 66.485 147.960 66.775 148.005 ;
        RECT 67.850 147.960 68.170 148.020 ;
        RECT 66.485 147.820 68.170 147.960 ;
        RECT 66.485 147.775 66.775 147.820 ;
        RECT 67.850 147.760 68.170 147.820 ;
        RECT 69.255 147.960 69.545 148.005 ;
        RECT 71.775 147.960 72.065 148.005 ;
        RECT 72.965 147.960 73.255 148.005 ;
        RECT 69.255 147.820 73.255 147.960 ;
        RECT 73.460 147.960 73.600 148.160 ;
        RECT 73.845 148.115 74.135 148.345 ;
        RECT 76.145 148.115 76.435 148.345 ;
        RECT 73.460 147.820 74.060 147.960 ;
        RECT 69.255 147.775 69.545 147.820 ;
        RECT 71.775 147.775 72.065 147.820 ;
        RECT 72.965 147.775 73.255 147.820 ;
        RECT 52.210 147.420 52.530 147.680 ;
        RECT 54.970 147.620 55.260 147.665 ;
        RECT 56.540 147.620 56.830 147.665 ;
        RECT 58.640 147.620 58.930 147.665 ;
        RECT 54.970 147.480 58.930 147.620 ;
        RECT 54.970 147.435 55.260 147.480 ;
        RECT 56.540 147.435 56.830 147.480 ;
        RECT 58.640 147.435 58.930 147.480 ;
        RECT 62.330 147.620 62.620 147.665 ;
        RECT 63.900 147.620 64.190 147.665 ;
        RECT 66.000 147.620 66.290 147.665 ;
        RECT 62.330 147.480 66.290 147.620 ;
        RECT 62.330 147.435 62.620 147.480 ;
        RECT 63.900 147.435 64.190 147.480 ;
        RECT 66.000 147.435 66.290 147.480 ;
        RECT 69.690 147.620 69.980 147.665 ;
        RECT 71.260 147.620 71.550 147.665 ;
        RECT 73.360 147.620 73.650 147.665 ;
        RECT 69.690 147.480 73.650 147.620 ;
        RECT 73.920 147.620 74.060 147.820 ;
        RECT 75.210 147.760 75.530 148.020 ;
        RECT 76.220 147.960 76.360 148.115 ;
        RECT 77.050 148.100 77.370 148.360 ;
        RECT 78.430 148.100 78.750 148.360 ;
        RECT 82.110 148.100 82.430 148.360 ;
        RECT 83.030 148.100 83.350 148.360 ;
        RECT 83.505 148.300 83.795 148.345 ;
        RECT 85.330 148.300 85.650 148.360 ;
        RECT 83.505 148.160 85.650 148.300 ;
        RECT 83.505 148.115 83.795 148.160 ;
        RECT 85.330 148.100 85.650 148.160 ;
        RECT 86.710 148.100 87.030 148.360 ;
        RECT 88.090 148.100 88.410 148.360 ;
        RECT 91.770 148.100 92.090 148.360 ;
        RECT 103.270 148.300 103.590 148.360 ;
        RECT 106.090 148.300 106.380 148.345 ;
        RECT 103.270 148.160 106.380 148.300 ;
        RECT 103.270 148.100 103.590 148.160 ;
        RECT 106.090 148.115 106.380 148.160 ;
        RECT 108.330 148.300 108.650 148.360 ;
        RECT 109.165 148.300 109.455 148.345 ;
        RECT 108.330 148.160 109.455 148.300 ;
        RECT 108.330 148.100 108.650 148.160 ;
        RECT 109.165 148.115 109.455 148.160 ;
        RECT 83.120 147.960 83.260 148.100 ;
        RECT 102.835 147.960 103.125 148.005 ;
        RECT 105.355 147.960 105.645 148.005 ;
        RECT 106.545 147.960 106.835 148.005 ;
        RECT 76.220 147.820 78.200 147.960 ;
        RECT 83.120 147.820 100.280 147.960 ;
        RECT 78.060 147.680 78.200 147.820 ;
        RECT 77.525 147.620 77.815 147.665 ;
        RECT 73.920 147.480 77.815 147.620 ;
        RECT 69.690 147.435 69.980 147.480 ;
        RECT 71.260 147.435 71.550 147.480 ;
        RECT 73.360 147.435 73.650 147.480 ;
        RECT 77.525 147.435 77.815 147.480 ;
        RECT 77.970 147.620 78.290 147.680 ;
        RECT 99.590 147.620 99.910 147.680 ;
        RECT 77.970 147.480 99.910 147.620 ;
        RECT 77.970 147.420 78.290 147.480 ;
        RECT 99.590 147.420 99.910 147.480 ;
        RECT 49.465 147.280 49.755 147.325 ;
        RECT 44.850 147.140 49.755 147.280 ;
        RECT 44.850 147.080 45.170 147.140 ;
        RECT 49.465 147.095 49.755 147.140 ;
        RECT 61.870 147.280 62.190 147.340 ;
        RECT 66.945 147.280 67.235 147.325 ;
        RECT 75.210 147.280 75.530 147.340 ;
        RECT 61.870 147.140 75.530 147.280 ;
        RECT 100.140 147.280 100.280 147.820 ;
        RECT 102.835 147.820 106.835 147.960 ;
        RECT 102.835 147.775 103.125 147.820 ;
        RECT 105.355 147.775 105.645 147.820 ;
        RECT 106.545 147.775 106.835 147.820 ;
        RECT 107.425 147.960 107.715 148.005 ;
        RECT 107.885 147.960 108.175 148.005 ;
        RECT 107.425 147.820 108.175 147.960 ;
        RECT 107.425 147.775 107.715 147.820 ;
        RECT 107.885 147.775 108.175 147.820 ;
        RECT 108.765 147.960 109.055 148.005 ;
        RECT 109.955 147.960 110.245 148.005 ;
        RECT 112.475 147.960 112.765 148.005 ;
        RECT 108.765 147.820 112.765 147.960 ;
        RECT 108.765 147.775 109.055 147.820 ;
        RECT 109.955 147.775 110.245 147.820 ;
        RECT 112.475 147.775 112.765 147.820 ;
        RECT 100.510 147.420 100.830 147.680 ;
        RECT 103.270 147.620 103.560 147.665 ;
        RECT 104.840 147.620 105.130 147.665 ;
        RECT 106.940 147.620 107.230 147.665 ;
        RECT 103.270 147.480 107.230 147.620 ;
        RECT 103.270 147.435 103.560 147.480 ;
        RECT 104.840 147.435 105.130 147.480 ;
        RECT 106.940 147.435 107.230 147.480 ;
        RECT 107.410 147.280 107.730 147.340 ;
        RECT 100.140 147.140 107.730 147.280 ;
        RECT 107.960 147.280 108.100 147.775 ;
        RECT 108.370 147.620 108.660 147.665 ;
        RECT 110.470 147.620 110.760 147.665 ;
        RECT 112.040 147.620 112.330 147.665 ;
        RECT 108.370 147.480 112.330 147.620 ;
        RECT 114.400 147.620 114.540 148.500 ;
        RECT 116.165 148.455 116.455 148.685 ;
        RECT 127.665 148.455 127.955 148.685 ;
        RECT 128.570 148.640 128.890 148.700 ;
        RECT 128.570 148.500 131.100 148.640 ;
        RECT 128.570 148.440 128.890 148.500 ;
        RECT 115.230 148.300 115.550 148.360 ;
        RECT 126.730 148.300 127.050 148.360 ;
        RECT 115.230 148.160 127.050 148.300 ;
        RECT 115.230 148.100 115.550 148.160 ;
        RECT 126.730 148.100 127.050 148.160 ;
        RECT 127.190 148.100 127.510 148.360 ;
        RECT 128.110 148.100 128.430 148.360 ;
        RECT 129.030 148.100 129.350 148.360 ;
        RECT 130.960 148.345 131.100 148.500 ;
        RECT 131.330 148.440 131.650 148.700 ;
        RECT 131.880 148.500 134.320 148.640 ;
        RECT 130.425 148.115 130.715 148.345 ;
        RECT 130.885 148.300 131.175 148.345 ;
        RECT 131.880 148.300 132.020 148.500 ;
        RECT 130.885 148.160 132.020 148.300 ;
        RECT 132.250 148.300 132.570 148.360 ;
        RECT 132.250 148.160 133.400 148.300 ;
        RECT 130.885 148.115 131.175 148.160 ;
        RECT 124.430 147.960 124.750 148.020 ;
        RECT 130.500 147.960 130.640 148.115 ;
        RECT 132.250 148.100 132.570 148.160 ;
        RECT 124.430 147.820 130.640 147.960 ;
        RECT 124.430 147.760 124.750 147.820 ;
        RECT 132.710 147.760 133.030 148.020 ;
        RECT 133.260 147.960 133.400 148.160 ;
        RECT 133.630 148.100 133.950 148.360 ;
        RECT 134.180 148.300 134.320 148.500 ;
        RECT 134.550 148.440 134.870 148.700 ;
        RECT 136.850 148.640 137.170 148.700 ;
        RECT 135.100 148.500 137.170 148.640 ;
        RECT 135.100 148.300 135.240 148.500 ;
        RECT 136.850 148.440 137.170 148.500 ;
        RECT 134.180 148.160 135.240 148.300 ;
        RECT 135.930 148.100 136.250 148.360 ;
        RECT 147.430 148.300 147.750 148.360 ;
        RECT 147.905 148.300 148.195 148.345 ;
        RECT 147.430 148.160 148.195 148.300 ;
        RECT 147.430 148.100 147.750 148.160 ;
        RECT 147.905 148.115 148.195 148.160 ;
        RECT 135.485 147.960 135.775 148.005 ;
        RECT 133.260 147.820 135.775 147.960 ;
        RECT 135.485 147.775 135.775 147.820 ;
        RECT 144.670 147.620 144.990 147.680 ;
        RECT 114.400 147.480 144.990 147.620 ;
        RECT 108.370 147.435 108.660 147.480 ;
        RECT 110.470 147.435 110.760 147.480 ;
        RECT 112.040 147.435 112.330 147.480 ;
        RECT 144.670 147.420 144.990 147.480 ;
        RECT 114.310 147.280 114.630 147.340 ;
        RECT 107.960 147.140 114.630 147.280 ;
        RECT 61.870 147.080 62.190 147.140 ;
        RECT 66.945 147.095 67.235 147.140 ;
        RECT 75.210 147.080 75.530 147.140 ;
        RECT 107.410 147.080 107.730 147.140 ;
        RECT 114.310 147.080 114.630 147.140 ;
        RECT 114.785 147.280 115.075 147.325 ;
        RECT 115.690 147.280 116.010 147.340 ;
        RECT 124.430 147.280 124.750 147.340 ;
        RECT 114.785 147.140 124.750 147.280 ;
        RECT 114.785 147.095 115.075 147.140 ;
        RECT 115.690 147.080 116.010 147.140 ;
        RECT 124.430 147.080 124.750 147.140 ;
        RECT 125.350 147.280 125.670 147.340 ;
        RECT 126.285 147.280 126.575 147.325 ;
        RECT 125.350 147.140 126.575 147.280 ;
        RECT 125.350 147.080 125.670 147.140 ;
        RECT 126.285 147.095 126.575 147.140 ;
        RECT 132.250 147.280 132.570 147.340 ;
        RECT 134.090 147.280 134.410 147.340 ;
        RECT 132.250 147.140 134.410 147.280 ;
        RECT 132.250 147.080 132.570 147.140 ;
        RECT 134.090 147.080 134.410 147.140 ;
        RECT 22.700 146.460 157.020 146.940 ;
        RECT 45.310 146.260 45.630 146.320 ;
        RECT 46.245 146.260 46.535 146.305 ;
        RECT 45.310 146.120 46.535 146.260 ;
        RECT 45.310 146.060 45.630 146.120 ;
        RECT 46.245 146.075 46.535 146.120 ;
        RECT 50.370 146.060 50.690 146.320 ;
        RECT 56.350 146.060 56.670 146.320 ;
        RECT 62.790 146.060 63.110 146.320 ;
        RECT 85.790 146.260 86.110 146.320 ;
        RECT 89.025 146.260 89.315 146.305 ;
        RECT 85.790 146.120 89.315 146.260 ;
        RECT 85.790 146.060 86.110 146.120 ;
        RECT 89.025 146.075 89.315 146.120 ;
        RECT 98.685 146.260 98.975 146.305 ;
        RECT 101.905 146.260 102.195 146.305 ;
        RECT 98.685 146.120 102.195 146.260 ;
        RECT 98.685 146.075 98.975 146.120 ;
        RECT 101.905 146.075 102.195 146.120 ;
        RECT 103.270 146.060 103.590 146.320 ;
        RECT 106.965 146.260 107.255 146.305 ;
        RECT 108.330 146.260 108.650 146.320 ;
        RECT 106.965 146.120 108.650 146.260 ;
        RECT 106.965 146.075 107.255 146.120 ;
        RECT 108.330 146.060 108.650 146.120 ;
        RECT 112.025 146.260 112.315 146.305 ;
        RECT 112.930 146.260 113.250 146.320 ;
        RECT 112.025 146.120 113.250 146.260 ;
        RECT 112.025 146.075 112.315 146.120 ;
        RECT 112.930 146.060 113.250 146.120 ;
        RECT 121.685 146.260 121.975 146.305 ;
        RECT 125.810 146.260 126.130 146.320 ;
        RECT 127.650 146.260 127.970 146.320 ;
        RECT 132.250 146.260 132.570 146.320 ;
        RECT 133.645 146.260 133.935 146.305 ;
        RECT 136.390 146.260 136.710 146.320 ;
        RECT 121.685 146.120 127.970 146.260 ;
        RECT 121.685 146.075 121.975 146.120 ;
        RECT 125.810 146.060 126.130 146.120 ;
        RECT 127.650 146.060 127.970 146.120 ;
        RECT 128.200 146.120 130.410 146.260 ;
        RECT 52.210 145.720 52.530 145.980 ;
        RECT 71.570 145.920 71.860 145.965 ;
        RECT 73.670 145.920 73.960 145.965 ;
        RECT 75.240 145.920 75.530 145.965 ;
        RECT 99.605 145.920 99.895 145.965 ;
        RECT 101.430 145.920 101.750 145.980 ;
        RECT 71.570 145.780 75.530 145.920 ;
        RECT 71.570 145.735 71.860 145.780 ;
        RECT 73.670 145.735 73.960 145.780 ;
        RECT 75.240 145.735 75.530 145.780 ;
        RECT 80.820 145.780 99.360 145.920 ;
        RECT 43.025 145.580 43.315 145.625 ;
        RECT 46.230 145.580 46.550 145.640 ;
        RECT 43.025 145.440 46.550 145.580 ;
        RECT 43.025 145.395 43.315 145.440 ;
        RECT 46.230 145.380 46.550 145.440 ;
        RECT 48.070 145.580 48.390 145.640 ;
        RECT 52.300 145.580 52.440 145.720 ;
        RECT 48.070 145.440 52.440 145.580 ;
        RECT 48.070 145.380 48.390 145.440 ;
        RECT 26.450 145.040 26.770 145.300 ;
        RECT 30.130 145.040 30.450 145.300 ;
        RECT 31.050 145.240 31.370 145.300 ;
        RECT 32.445 145.240 32.735 145.285 ;
        RECT 31.050 145.100 32.735 145.240 ;
        RECT 31.050 145.040 31.370 145.100 ;
        RECT 32.445 145.055 32.735 145.100 ;
        RECT 42.550 145.040 42.870 145.300 ;
        RECT 44.850 145.040 45.170 145.300 ;
        RECT 47.165 145.055 47.455 145.285 ;
        RECT 47.610 145.240 47.930 145.300 ;
        RECT 48.620 145.285 48.760 145.440 ;
        RECT 52.670 145.380 52.990 145.640 ;
        RECT 57.730 145.580 58.050 145.640 ;
        RECT 80.820 145.625 80.960 145.780 ;
        RECT 71.965 145.580 72.255 145.625 ;
        RECT 73.155 145.580 73.445 145.625 ;
        RECT 75.675 145.580 75.965 145.625 ;
        RECT 57.730 145.440 65.320 145.580 ;
        RECT 57.730 145.380 58.050 145.440 ;
        RECT 47.610 145.100 48.125 145.240 ;
        RECT 30.220 144.900 30.360 145.040 ;
        RECT 33.350 144.900 33.670 144.960 ;
        RECT 30.220 144.760 33.670 144.900 ;
        RECT 33.350 144.700 33.670 144.760 ;
        RECT 43.930 144.900 44.250 144.960 ;
        RECT 47.240 144.900 47.380 145.055 ;
        RECT 47.610 145.040 47.930 145.100 ;
        RECT 48.545 145.055 48.835 145.285 ;
        RECT 49.695 145.240 49.985 145.285 ;
        RECT 51.750 145.240 52.070 145.300 ;
        RECT 49.695 145.100 52.070 145.240 ;
        RECT 49.695 145.055 49.985 145.100 ;
        RECT 51.750 145.040 52.070 145.100 ;
        RECT 52.225 145.240 52.515 145.285 ;
        RECT 52.760 145.240 52.900 145.380 ;
        RECT 52.225 145.100 52.900 145.240 ;
        RECT 57.285 145.240 57.575 145.285 ;
        RECT 58.190 145.240 58.510 145.300 ;
        RECT 58.740 145.285 58.880 145.440 ;
        RECT 57.285 145.100 58.510 145.240 ;
        RECT 52.225 145.055 52.515 145.100 ;
        RECT 57.285 145.055 57.575 145.100 ;
        RECT 58.190 145.040 58.510 145.100 ;
        RECT 58.665 145.055 58.955 145.285 ;
        RECT 63.725 145.240 64.015 145.285 ;
        RECT 64.630 145.240 64.950 145.300 ;
        RECT 65.180 145.285 65.320 145.440 ;
        RECT 71.965 145.440 75.965 145.580 ;
        RECT 71.965 145.395 72.255 145.440 ;
        RECT 73.155 145.395 73.445 145.440 ;
        RECT 75.675 145.395 75.965 145.440 ;
        RECT 80.745 145.395 81.035 145.625 ;
        RECT 81.205 145.395 81.495 145.625 ;
        RECT 86.265 145.580 86.555 145.625 ;
        RECT 96.845 145.580 97.135 145.625 ;
        RECT 98.670 145.580 98.990 145.640 ;
        RECT 86.265 145.440 92.920 145.580 ;
        RECT 86.265 145.395 86.555 145.440 ;
        RECT 63.725 145.100 64.950 145.240 ;
        RECT 63.725 145.055 64.015 145.100 ;
        RECT 64.630 145.040 64.950 145.100 ;
        RECT 65.105 145.055 65.395 145.285 ;
        RECT 71.085 145.240 71.375 145.285 ;
        RECT 69.780 145.100 71.375 145.240 ;
        RECT 43.930 144.760 47.380 144.900 ;
        RECT 49.005 144.900 49.295 144.945 ;
        RECT 52.685 144.900 52.975 144.945 ;
        RECT 49.005 144.760 52.975 144.900 ;
        RECT 43.930 144.700 44.250 144.760 ;
        RECT 49.005 144.715 49.295 144.760 ;
        RECT 52.685 144.715 52.975 144.760 ;
        RECT 66.025 144.900 66.315 144.945 ;
        RECT 67.390 144.900 67.710 144.960 ;
        RECT 66.025 144.760 67.710 144.900 ;
        RECT 66.025 144.715 66.315 144.760 ;
        RECT 67.390 144.700 67.710 144.760 ;
        RECT 67.850 144.900 68.170 144.960 ;
        RECT 69.780 144.945 69.920 145.100 ;
        RECT 71.085 145.055 71.375 145.100 ;
        RECT 76.130 145.240 76.450 145.300 ;
        RECT 80.270 145.240 80.590 145.300 ;
        RECT 81.280 145.240 81.420 145.395 ;
        RECT 76.130 145.100 81.420 145.240 ;
        RECT 76.130 145.040 76.450 145.100 ;
        RECT 80.270 145.040 80.590 145.100 ;
        RECT 86.710 145.040 87.030 145.300 ;
        RECT 91.770 145.285 92.090 145.300 ;
        RECT 92.780 145.285 92.920 145.440 ;
        RECT 93.695 145.440 95.680 145.580 ;
        RECT 93.695 145.285 93.835 145.440 ;
        RECT 95.540 145.300 95.680 145.440 ;
        RECT 96.845 145.440 98.990 145.580 ;
        RECT 99.220 145.580 99.360 145.780 ;
        RECT 99.605 145.780 101.750 145.920 ;
        RECT 99.605 145.735 99.895 145.780 ;
        RECT 101.430 145.720 101.750 145.780 ;
        RECT 115.270 145.920 115.560 145.965 ;
        RECT 117.370 145.920 117.660 145.965 ;
        RECT 118.940 145.920 119.230 145.965 ;
        RECT 115.270 145.780 119.230 145.920 ;
        RECT 115.270 145.735 115.560 145.780 ;
        RECT 117.370 145.735 117.660 145.780 ;
        RECT 118.940 145.735 119.230 145.780 ;
        RECT 126.745 145.920 127.035 145.965 ;
        RECT 127.190 145.920 127.510 145.980 ;
        RECT 126.745 145.780 127.510 145.920 ;
        RECT 126.745 145.735 127.035 145.780 ;
        RECT 127.190 145.720 127.510 145.780 ;
        RECT 102.810 145.580 103.130 145.640 ;
        RECT 109.250 145.580 109.570 145.640 ;
        RECT 99.220 145.440 106.260 145.580 ;
        RECT 96.845 145.395 97.135 145.440 ;
        RECT 98.670 145.380 98.990 145.440 ;
        RECT 102.810 145.380 103.130 145.440 ;
        RECT 91.760 145.240 92.090 145.285 ;
        RECT 91.575 145.100 92.090 145.240 ;
        RECT 91.760 145.055 92.090 145.100 ;
        RECT 92.705 145.055 92.995 145.285 ;
        RECT 93.620 145.055 93.910 145.285 ;
        RECT 94.085 145.240 94.375 145.285 ;
        RECT 94.990 145.240 95.310 145.300 ;
        RECT 94.085 145.100 95.310 145.240 ;
        RECT 94.085 145.055 94.375 145.100 ;
        RECT 91.770 145.040 92.090 145.055 ;
        RECT 69.705 144.900 69.995 144.945 ;
        RECT 67.850 144.760 69.995 144.900 ;
        RECT 67.850 144.700 68.170 144.760 ;
        RECT 69.705 144.715 69.995 144.760 ;
        RECT 72.420 144.900 72.710 144.945 ;
        RECT 74.750 144.900 75.070 144.960 ;
        RECT 72.420 144.760 75.070 144.900 ;
        RECT 72.420 144.715 72.710 144.760 ;
        RECT 74.750 144.700 75.070 144.760 ;
        RECT 75.670 144.900 75.990 144.960 ;
        RECT 83.950 144.900 84.270 144.960 ;
        RECT 88.865 144.900 89.155 144.945 ;
        RECT 75.670 144.760 78.660 144.900 ;
        RECT 75.670 144.700 75.990 144.760 ;
        RECT 25.530 144.360 25.850 144.620 ;
        RECT 29.210 144.360 29.530 144.620 ;
        RECT 29.670 144.560 29.990 144.620 ;
        RECT 31.525 144.560 31.815 144.605 ;
        RECT 29.670 144.420 31.815 144.560 ;
        RECT 29.670 144.360 29.990 144.420 ;
        RECT 31.525 144.375 31.815 144.420 ;
        RECT 44.405 144.560 44.695 144.605 ;
        RECT 47.150 144.560 47.470 144.620 ;
        RECT 44.405 144.420 47.470 144.560 ;
        RECT 44.405 144.375 44.695 144.420 ;
        RECT 47.150 144.360 47.470 144.420 ;
        RECT 49.910 144.560 50.230 144.620 ;
        RECT 51.290 144.560 51.610 144.620 ;
        RECT 49.910 144.420 51.610 144.560 ;
        RECT 49.910 144.360 50.230 144.420 ;
        RECT 51.290 144.360 51.610 144.420 ;
        RECT 58.205 144.560 58.495 144.605 ;
        RECT 59.110 144.560 59.430 144.620 ;
        RECT 58.205 144.420 59.430 144.560 ;
        RECT 58.205 144.375 58.495 144.420 ;
        RECT 59.110 144.360 59.430 144.420 ;
        RECT 61.410 144.560 61.730 144.620 ;
        RECT 64.645 144.560 64.935 144.605 ;
        RECT 61.410 144.420 64.935 144.560 ;
        RECT 61.410 144.360 61.730 144.420 ;
        RECT 64.645 144.375 64.935 144.420 ;
        RECT 77.050 144.560 77.370 144.620 ;
        RECT 78.520 144.605 78.660 144.760 ;
        RECT 83.950 144.760 89.155 144.900 ;
        RECT 83.950 144.700 84.270 144.760 ;
        RECT 88.865 144.715 89.155 144.760 ;
        RECT 89.945 144.900 90.235 144.945 ;
        RECT 89.945 144.760 91.540 144.900 ;
        RECT 89.945 144.715 90.235 144.760 ;
        RECT 91.400 144.620 91.540 144.760 ;
        RECT 92.245 144.715 92.535 144.945 ;
        RECT 92.780 144.900 92.920 145.055 ;
        RECT 94.990 145.040 95.310 145.100 ;
        RECT 95.450 145.040 95.770 145.300 ;
        RECT 101.430 145.240 101.750 145.300 ;
        RECT 106.120 145.285 106.260 145.440 ;
        RECT 107.960 145.440 109.570 145.580 ;
        RECT 107.960 145.285 108.100 145.440 ;
        RECT 109.250 145.380 109.570 145.440 ;
        RECT 115.665 145.580 115.955 145.625 ;
        RECT 116.855 145.580 117.145 145.625 ;
        RECT 119.375 145.580 119.665 145.625 ;
        RECT 115.665 145.440 119.665 145.580 ;
        RECT 115.665 145.395 115.955 145.440 ;
        RECT 116.855 145.395 117.145 145.440 ;
        RECT 119.375 145.395 119.665 145.440 ;
        RECT 102.365 145.240 102.655 145.285 ;
        RECT 101.430 145.100 102.655 145.240 ;
        RECT 101.430 145.040 101.750 145.100 ;
        RECT 102.365 145.055 102.655 145.100 ;
        RECT 106.045 145.055 106.335 145.285 ;
        RECT 107.885 145.055 108.175 145.285 ;
        RECT 108.330 145.040 108.650 145.300 ;
        RECT 108.790 145.040 109.110 145.300 ;
        RECT 109.710 145.040 110.030 145.300 ;
        RECT 110.630 145.040 110.950 145.300 ;
        RECT 114.770 145.040 115.090 145.300 ;
        RECT 124.430 145.040 124.750 145.300 ;
        RECT 125.810 145.285 126.130 145.300 ;
        RECT 124.905 145.055 125.195 145.285 ;
        RECT 125.810 145.055 126.345 145.285 ;
        RECT 94.545 144.900 94.835 144.945 ;
        RECT 92.780 144.760 94.835 144.900 ;
        RECT 94.545 144.715 94.835 144.760 ;
        RECT 99.130 144.900 99.450 144.960 ;
        RECT 100.065 144.900 100.355 144.945 ;
        RECT 99.130 144.760 100.355 144.900 ;
        RECT 77.985 144.560 78.275 144.605 ;
        RECT 77.050 144.420 78.275 144.560 ;
        RECT 77.050 144.360 77.370 144.420 ;
        RECT 77.985 144.375 78.275 144.420 ;
        RECT 78.445 144.375 78.735 144.605 ;
        RECT 80.270 144.360 80.590 144.620 ;
        RECT 88.090 144.360 88.410 144.620 ;
        RECT 90.850 144.360 91.170 144.620 ;
        RECT 91.310 144.360 91.630 144.620 ;
        RECT 92.320 144.560 92.460 144.715 ;
        RECT 99.130 144.700 99.450 144.760 ;
        RECT 100.065 144.715 100.355 144.760 ;
        RECT 100.510 144.900 100.830 144.960 ;
        RECT 100.985 144.900 101.275 144.945 ;
        RECT 100.510 144.760 101.275 144.900 ;
        RECT 100.510 144.700 100.830 144.760 ;
        RECT 100.985 144.715 101.275 144.760 ;
        RECT 116.120 144.900 116.410 144.945 ;
        RECT 117.070 144.900 117.390 144.960 ;
        RECT 116.120 144.760 117.390 144.900 ;
        RECT 124.980 144.900 125.120 145.055 ;
        RECT 125.810 145.040 126.130 145.055 ;
        RECT 126.730 145.040 127.050 145.300 ;
        RECT 128.200 145.285 128.340 146.120 ;
        RECT 130.270 145.920 130.410 146.120 ;
        RECT 132.250 146.120 133.935 146.260 ;
        RECT 132.250 146.060 132.570 146.120 ;
        RECT 133.645 146.075 133.935 146.120 ;
        RECT 134.180 146.120 136.710 146.260 ;
        RECT 134.180 145.920 134.320 146.120 ;
        RECT 136.390 146.060 136.710 146.120 ;
        RECT 136.850 146.260 137.170 146.320 ;
        RECT 141.005 146.260 141.295 146.305 ;
        RECT 136.850 146.120 141.295 146.260 ;
        RECT 136.850 146.060 137.170 146.120 ;
        RECT 141.005 146.075 141.295 146.120 ;
        RECT 145.145 146.260 145.435 146.305 ;
        RECT 146.525 146.260 146.815 146.305 ;
        RECT 145.145 146.120 146.815 146.260 ;
        RECT 145.145 146.075 145.435 146.120 ;
        RECT 146.525 146.075 146.815 146.120 ;
        RECT 147.430 146.060 147.750 146.320 ;
        RECT 130.270 145.780 134.320 145.920 ;
        RECT 135.485 145.920 135.775 145.965 ;
        RECT 137.785 145.920 138.075 145.965 ;
        RECT 141.910 145.920 142.230 145.980 ;
        RECT 135.485 145.780 142.230 145.920 ;
        RECT 135.485 145.735 135.775 145.780 ;
        RECT 137.785 145.735 138.075 145.780 ;
        RECT 141.910 145.720 142.230 145.780 ;
        RECT 144.210 145.920 144.530 145.980 ;
        RECT 148.365 145.920 148.655 145.965 ;
        RECT 144.210 145.780 148.655 145.920 ;
        RECT 144.210 145.720 144.530 145.780 ;
        RECT 148.365 145.735 148.655 145.780 ;
        RECT 151.110 145.920 151.400 145.965 ;
        RECT 152.680 145.920 152.970 145.965 ;
        RECT 154.780 145.920 155.070 145.965 ;
        RECT 151.110 145.780 155.070 145.920 ;
        RECT 151.110 145.735 151.400 145.780 ;
        RECT 152.680 145.735 152.970 145.780 ;
        RECT 154.780 145.735 155.070 145.780 ;
        RECT 129.030 145.580 129.350 145.640 ;
        RECT 132.710 145.580 133.030 145.640 ;
        RECT 135.930 145.580 136.250 145.640 ;
        RECT 150.675 145.580 150.965 145.625 ;
        RECT 153.195 145.580 153.485 145.625 ;
        RECT 154.385 145.580 154.675 145.625 ;
        RECT 129.030 145.440 133.030 145.580 ;
        RECT 129.030 145.380 129.350 145.440 ;
        RECT 132.710 145.380 133.030 145.440 ;
        RECT 134.180 145.440 136.250 145.580 ;
        RECT 128.125 145.055 128.415 145.285 ;
        RECT 129.965 145.055 130.255 145.285 ;
        RECT 131.345 145.240 131.635 145.285 ;
        RECT 134.180 145.240 134.320 145.440 ;
        RECT 135.930 145.380 136.250 145.440 ;
        RECT 141.540 145.440 143.060 145.580 ;
        RECT 141.540 145.285 141.680 145.440 ;
        RECT 131.345 145.100 134.320 145.240 ;
        RECT 131.345 145.055 131.635 145.100 ;
        RECT 136.865 145.055 137.155 145.285 ;
        RECT 139.165 145.240 139.455 145.285 ;
        RECT 137.400 145.100 139.455 145.240 ;
        RECT 128.570 144.900 128.890 144.960 ;
        RECT 124.980 144.760 128.890 144.900 ;
        RECT 130.040 144.900 130.180 145.055 ;
        RECT 131.790 144.900 132.110 144.960 ;
        RECT 130.040 144.760 132.110 144.900 ;
        RECT 116.120 144.715 116.410 144.760 ;
        RECT 117.070 144.700 117.390 144.760 ;
        RECT 128.570 144.700 128.890 144.760 ;
        RECT 131.790 144.700 132.110 144.760 ;
        RECT 132.265 144.900 132.555 144.945 ;
        RECT 133.645 144.900 133.935 144.945 ;
        RECT 132.265 144.760 133.935 144.900 ;
        RECT 132.265 144.715 132.555 144.760 ;
        RECT 133.645 144.715 133.935 144.760 ;
        RECT 134.090 144.900 134.410 144.960 ;
        RECT 136.940 144.900 137.080 145.055 ;
        RECT 134.090 144.760 137.080 144.900 ;
        RECT 134.090 144.700 134.410 144.760 ;
        RECT 95.910 144.560 96.230 144.620 ;
        RECT 92.320 144.420 96.230 144.560 ;
        RECT 95.910 144.360 96.230 144.420 ;
        RECT 96.370 144.360 96.690 144.620 ;
        RECT 96.830 144.560 97.150 144.620 ;
        RECT 98.685 144.560 98.975 144.605 ;
        RECT 96.830 144.420 98.975 144.560 ;
        RECT 96.830 144.360 97.150 144.420 ;
        RECT 98.685 144.375 98.975 144.420 ;
        RECT 105.585 144.560 105.875 144.605 ;
        RECT 107.870 144.560 108.190 144.620 ;
        RECT 108.790 144.560 109.110 144.620 ;
        RECT 105.585 144.420 109.110 144.560 ;
        RECT 105.585 144.375 105.875 144.420 ;
        RECT 107.870 144.360 108.190 144.420 ;
        RECT 108.790 144.360 109.110 144.420 ;
        RECT 123.525 144.560 123.815 144.605 ;
        RECT 127.665 144.560 127.955 144.605 ;
        RECT 123.525 144.420 127.955 144.560 ;
        RECT 123.525 144.375 123.815 144.420 ;
        RECT 127.665 144.375 127.955 144.420 ;
        RECT 130.410 144.360 130.730 144.620 ;
        RECT 132.725 144.560 133.015 144.605 ;
        RECT 137.400 144.560 137.540 145.100 ;
        RECT 139.165 145.055 139.455 145.100 ;
        RECT 141.465 145.055 141.755 145.285 ;
        RECT 141.910 145.240 142.230 145.300 ;
        RECT 142.920 145.285 143.060 145.440 ;
        RECT 150.675 145.440 154.675 145.580 ;
        RECT 150.675 145.395 150.965 145.440 ;
        RECT 153.195 145.395 153.485 145.440 ;
        RECT 154.385 145.395 154.675 145.440 ;
        RECT 142.845 145.240 143.135 145.285 ;
        RECT 143.750 145.240 144.070 145.300 ;
        RECT 144.225 145.240 144.515 145.285 ;
        RECT 141.910 145.100 142.600 145.240 ;
        RECT 141.910 145.040 142.230 145.100 ;
        RECT 142.460 144.900 142.600 145.100 ;
        RECT 142.845 145.100 144.515 145.240 ;
        RECT 142.845 145.055 143.135 145.100 ;
        RECT 143.750 145.040 144.070 145.100 ;
        RECT 144.225 145.055 144.515 145.100 ;
        RECT 155.250 145.040 155.570 145.300 ;
        RECT 143.305 144.900 143.595 144.945 ;
        RECT 142.460 144.760 143.595 144.900 ;
        RECT 143.305 144.715 143.595 144.760 ;
        RECT 145.590 144.900 145.910 144.960 ;
        RECT 147.430 144.900 147.750 144.960 ;
        RECT 145.590 144.760 147.750 144.900 ;
        RECT 145.590 144.700 145.910 144.760 ;
        RECT 147.430 144.700 147.750 144.760 ;
        RECT 152.950 144.900 153.270 144.960 ;
        RECT 153.930 144.900 154.220 144.945 ;
        RECT 152.950 144.760 154.220 144.900 ;
        RECT 152.950 144.700 153.270 144.760 ;
        RECT 153.930 144.715 154.220 144.760 ;
        RECT 132.725 144.420 137.540 144.560 ;
        RECT 139.610 144.560 139.930 144.620 ;
        RECT 140.085 144.560 140.375 144.605 ;
        RECT 139.610 144.420 140.375 144.560 ;
        RECT 132.725 144.375 133.015 144.420 ;
        RECT 139.610 144.360 139.930 144.420 ;
        RECT 140.085 144.375 140.375 144.420 ;
        RECT 142.845 144.560 143.135 144.605 ;
        RECT 146.605 144.560 146.895 144.605 ;
        RECT 148.810 144.560 149.130 144.620 ;
        RECT 150.650 144.560 150.970 144.620 ;
        RECT 142.845 144.420 150.970 144.560 ;
        RECT 142.845 144.375 143.135 144.420 ;
        RECT 146.605 144.375 146.895 144.420 ;
        RECT 148.810 144.360 149.130 144.420 ;
        RECT 150.650 144.360 150.970 144.420 ;
        RECT 22.700 143.740 157.820 144.220 ;
        RECT 31.050 143.340 31.370 143.600 ;
        RECT 42.105 143.540 42.395 143.585 ;
        RECT 42.550 143.540 42.870 143.600 ;
        RECT 42.105 143.400 42.870 143.540 ;
        RECT 42.105 143.355 42.395 143.400 ;
        RECT 42.550 143.340 42.870 143.400 ;
        RECT 43.930 143.540 44.250 143.600 ;
        RECT 44.405 143.540 44.695 143.585 ;
        RECT 43.930 143.400 44.695 143.540 ;
        RECT 43.930 143.340 44.250 143.400 ;
        RECT 44.405 143.355 44.695 143.400 ;
        RECT 53.065 143.540 53.355 143.585 ;
        RECT 56.350 143.540 56.670 143.600 ;
        RECT 60.505 143.540 60.795 143.585 ;
        RECT 53.065 143.400 55.245 143.540 ;
        RECT 53.065 143.355 53.355 143.400 ;
        RECT 25.530 143.245 25.850 143.260 ;
        RECT 25.500 143.200 25.850 143.245 ;
        RECT 25.335 143.060 25.850 143.200 ;
        RECT 25.500 143.015 25.850 143.060 ;
        RECT 25.530 143.000 25.850 143.015 ;
        RECT 24.150 142.660 24.470 142.920 ;
        RECT 31.140 142.860 31.280 143.340 ;
        RECT 43.485 143.200 43.775 143.245 ;
        RECT 47.610 143.200 47.930 143.260 ;
        RECT 54.065 143.200 54.355 143.245 ;
        RECT 33.670 143.060 41.860 143.200 ;
        RECT 32.905 142.860 33.195 142.905 ;
        RECT 33.670 142.860 33.810 143.060 ;
        RECT 31.140 142.720 33.810 142.860 ;
        RECT 35.190 142.860 35.510 142.920 ;
        RECT 41.720 142.905 41.860 143.060 ;
        RECT 43.485 143.060 47.930 143.200 ;
        RECT 43.485 143.015 43.775 143.060 ;
        RECT 40.265 142.860 40.555 142.905 ;
        RECT 35.190 142.720 40.555 142.860 ;
        RECT 32.905 142.675 33.195 142.720 ;
        RECT 35.190 142.660 35.510 142.720 ;
        RECT 40.265 142.675 40.555 142.720 ;
        RECT 41.645 142.860 41.935 142.905 ;
        RECT 42.550 142.860 42.870 142.920 ;
        RECT 41.645 142.720 42.870 142.860 ;
        RECT 41.645 142.675 41.935 142.720 ;
        RECT 42.550 142.660 42.870 142.720 ;
        RECT 43.025 142.675 43.315 142.905 ;
        RECT 45.325 142.675 45.615 142.905 ;
        RECT 25.045 142.520 25.335 142.565 ;
        RECT 26.235 142.520 26.525 142.565 ;
        RECT 28.755 142.520 29.045 142.565 ;
        RECT 25.045 142.380 29.045 142.520 ;
        RECT 25.045 142.335 25.335 142.380 ;
        RECT 26.235 142.335 26.525 142.380 ;
        RECT 28.755 142.335 29.045 142.380 ;
        RECT 31.985 142.335 32.275 142.565 ;
        RECT 24.650 142.180 24.940 142.225 ;
        RECT 26.750 142.180 27.040 142.225 ;
        RECT 28.320 142.180 28.610 142.225 ;
        RECT 24.650 142.040 28.610 142.180 ;
        RECT 32.060 142.180 32.200 142.335 ;
        RECT 32.430 142.320 32.750 142.580 ;
        RECT 33.350 142.320 33.670 142.580 ;
        RECT 39.805 142.520 40.095 142.565 ;
        RECT 40.710 142.520 41.030 142.580 ;
        RECT 39.805 142.380 41.030 142.520 ;
        RECT 39.805 142.335 40.095 142.380 ;
        RECT 40.710 142.320 41.030 142.380 ;
        RECT 36.110 142.180 36.430 142.240 ;
        RECT 43.100 142.180 43.240 142.675 ;
        RECT 45.400 142.520 45.540 142.675 ;
        RECT 45.770 142.660 46.090 142.920 ;
        RECT 47.240 142.905 47.380 143.060 ;
        RECT 47.610 143.000 47.930 143.060 ;
        RECT 53.680 143.060 54.355 143.200 ;
        RECT 47.165 142.675 47.455 142.905 ;
        RECT 51.305 142.860 51.595 142.905 ;
        RECT 52.210 142.860 52.530 142.920 ;
        RECT 51.305 142.720 52.530 142.860 ;
        RECT 53.680 142.860 53.820 143.060 ;
        RECT 54.065 143.015 54.355 143.060 ;
        RECT 54.510 143.000 54.830 143.260 ;
        RECT 55.105 143.200 55.245 143.400 ;
        RECT 56.350 143.400 60.795 143.540 ;
        RECT 56.350 143.340 56.670 143.400 ;
        RECT 60.505 143.355 60.795 143.400 ;
        RECT 70.150 143.340 70.470 143.600 ;
        RECT 74.750 143.340 75.070 143.600 ;
        RECT 78.445 143.540 78.735 143.585 ;
        RECT 80.270 143.540 80.590 143.600 ;
        RECT 78.445 143.400 80.590 143.540 ;
        RECT 78.445 143.355 78.735 143.400 ;
        RECT 80.270 143.340 80.590 143.400 ;
        RECT 86.710 143.540 87.030 143.600 ;
        RECT 87.645 143.540 87.935 143.585 ;
        RECT 86.710 143.400 87.935 143.540 ;
        RECT 86.710 143.340 87.030 143.400 ;
        RECT 87.645 143.355 87.935 143.400 ;
        RECT 91.310 143.540 91.630 143.600 ;
        RECT 92.245 143.540 92.535 143.585 ;
        RECT 91.310 143.400 92.535 143.540 ;
        RECT 55.525 143.200 55.815 143.245 ;
        RECT 57.270 143.200 57.590 143.260 ;
        RECT 55.105 143.060 57.590 143.200 ;
        RECT 55.525 143.015 55.815 143.060 ;
        RECT 57.270 143.000 57.590 143.060 ;
        RECT 56.825 142.860 57.115 142.905 ;
        RECT 53.680 142.720 57.115 142.860 ;
        RECT 51.305 142.675 51.595 142.720 ;
        RECT 52.210 142.660 52.530 142.720 ;
        RECT 56.825 142.675 57.115 142.720 ;
        RECT 66.945 142.860 67.235 142.905 ;
        RECT 69.705 142.860 69.995 142.905 ;
        RECT 71.070 142.860 71.390 142.920 ;
        RECT 66.945 142.720 68.080 142.860 ;
        RECT 66.945 142.675 67.235 142.720 ;
        RECT 57.270 142.520 57.590 142.580 ;
        RECT 59.585 142.520 59.875 142.565 ;
        RECT 45.400 142.380 59.875 142.520 ;
        RECT 57.270 142.320 57.590 142.380 ;
        RECT 59.585 142.335 59.875 142.380 ;
        RECT 63.250 142.320 63.570 142.580 ;
        RECT 56.365 142.180 56.655 142.225 ;
        RECT 59.110 142.180 59.430 142.240 ;
        RECT 67.940 142.225 68.080 142.720 ;
        RECT 69.705 142.720 71.390 142.860 ;
        RECT 69.705 142.675 69.995 142.720 ;
        RECT 71.070 142.660 71.390 142.720 ;
        RECT 75.670 142.660 75.990 142.920 ;
        RECT 77.050 142.660 77.370 142.920 ;
        RECT 77.510 142.660 77.830 142.920 ;
        RECT 82.110 142.905 82.430 142.920 ;
        RECT 82.080 142.675 82.430 142.905 ;
        RECT 87.720 142.860 87.860 143.355 ;
        RECT 91.310 143.340 91.630 143.400 ;
        RECT 92.245 143.355 92.535 143.400 ;
        RECT 97.765 143.540 98.055 143.585 ;
        RECT 98.210 143.540 98.530 143.600 ;
        RECT 97.765 143.400 98.530 143.540 ;
        RECT 97.765 143.355 98.055 143.400 ;
        RECT 98.210 143.340 98.530 143.400 ;
        RECT 109.710 143.540 110.030 143.600 ;
        RECT 112.485 143.540 112.775 143.585 ;
        RECT 109.710 143.400 112.775 143.540 ;
        RECT 109.710 143.340 110.030 143.400 ;
        RECT 112.485 143.355 112.775 143.400 ;
        RECT 126.285 143.540 126.575 143.585 ;
        RECT 126.730 143.540 127.050 143.600 ;
        RECT 126.285 143.400 127.050 143.540 ;
        RECT 126.285 143.355 126.575 143.400 ;
        RECT 126.730 143.340 127.050 143.400 ;
        RECT 134.105 143.540 134.395 143.585 ;
        RECT 135.930 143.540 136.250 143.600 ;
        RECT 134.105 143.400 136.250 143.540 ;
        RECT 134.105 143.355 134.395 143.400 ;
        RECT 135.930 143.340 136.250 143.400 ;
        RECT 141.910 143.540 142.230 143.600 ;
        RECT 142.385 143.540 142.675 143.585 ;
        RECT 141.910 143.400 142.675 143.540 ;
        RECT 141.910 143.340 142.230 143.400 ;
        RECT 142.385 143.355 142.675 143.400 ;
        RECT 143.305 143.540 143.595 143.585 ;
        RECT 144.210 143.540 144.530 143.600 ;
        RECT 143.305 143.400 144.530 143.540 ;
        RECT 143.305 143.355 143.595 143.400 ;
        RECT 144.210 143.340 144.530 143.400 ;
        RECT 147.445 143.540 147.735 143.585 ;
        RECT 150.205 143.540 150.495 143.585 ;
        RECT 147.445 143.400 150.495 143.540 ;
        RECT 147.445 143.355 147.735 143.400 ;
        RECT 150.205 143.355 150.495 143.400 ;
        RECT 152.950 143.340 153.270 143.600 ;
        RECT 93.625 143.200 93.915 143.245 ;
        RECT 96.370 143.200 96.690 143.260 ;
        RECT 109.250 143.200 109.570 143.260 ;
        RECT 118.925 143.200 119.215 143.245 ;
        RECT 93.625 143.060 96.690 143.200 ;
        RECT 93.625 143.015 93.915 143.060 ;
        RECT 96.370 143.000 96.690 143.060 ;
        RECT 97.840 143.060 104.420 143.200 ;
        RECT 89.025 142.860 89.315 142.905 ;
        RECT 87.720 142.720 89.315 142.860 ;
        RECT 89.025 142.675 89.315 142.720 ;
        RECT 90.850 142.860 91.170 142.920 ;
        RECT 92.705 142.860 92.995 142.905 ;
        RECT 90.850 142.720 92.995 142.860 ;
        RECT 82.110 142.660 82.430 142.675 ;
        RECT 90.850 142.660 91.170 142.720 ;
        RECT 92.705 142.675 92.995 142.720 ;
        RECT 94.085 142.675 94.375 142.905 ;
        RECT 94.545 142.860 94.835 142.905 ;
        RECT 95.450 142.860 95.770 142.920 ;
        RECT 94.545 142.720 95.770 142.860 ;
        RECT 94.545 142.675 94.835 142.720 ;
        RECT 70.625 142.520 70.915 142.565 ;
        RECT 79.350 142.520 79.670 142.580 ;
        RECT 80.745 142.520 81.035 142.565 ;
        RECT 70.625 142.380 75.900 142.520 ;
        RECT 70.625 142.335 70.915 142.380 ;
        RECT 75.760 142.240 75.900 142.380 ;
        RECT 79.350 142.380 81.035 142.520 ;
        RECT 79.350 142.320 79.670 142.380 ;
        RECT 80.745 142.335 81.035 142.380 ;
        RECT 81.625 142.520 81.915 142.565 ;
        RECT 82.815 142.520 83.105 142.565 ;
        RECT 85.335 142.520 85.625 142.565 ;
        RECT 81.625 142.380 85.625 142.520 ;
        RECT 81.625 142.335 81.915 142.380 ;
        RECT 82.815 142.335 83.105 142.380 ;
        RECT 85.335 142.335 85.625 142.380 ;
        RECT 32.060 142.040 50.140 142.180 ;
        RECT 24.650 141.995 24.940 142.040 ;
        RECT 26.750 141.995 27.040 142.040 ;
        RECT 28.320 141.995 28.610 142.040 ;
        RECT 36.110 141.980 36.430 142.040 ;
        RECT 34.270 141.640 34.590 141.900 ;
        RECT 36.570 141.640 36.890 141.900 ;
        RECT 41.185 141.840 41.475 141.885 ;
        RECT 41.630 141.840 41.950 141.900 ;
        RECT 41.185 141.700 41.950 141.840 ;
        RECT 41.185 141.655 41.475 141.700 ;
        RECT 41.630 141.640 41.950 141.700 ;
        RECT 46.705 141.840 46.995 141.885 ;
        RECT 47.610 141.840 47.930 141.900 ;
        RECT 46.705 141.700 47.930 141.840 ;
        RECT 46.705 141.655 46.995 141.700 ;
        RECT 47.610 141.640 47.930 141.700 ;
        RECT 48.070 141.840 48.390 141.900 ;
        RECT 50.000 141.885 50.140 142.040 ;
        RECT 56.365 142.040 59.430 142.180 ;
        RECT 56.365 141.995 56.655 142.040 ;
        RECT 59.110 141.980 59.430 142.040 ;
        RECT 67.865 141.995 68.155 142.225 ;
        RECT 75.670 141.980 75.990 142.240 ;
        RECT 81.230 142.180 81.520 142.225 ;
        RECT 83.330 142.180 83.620 142.225 ;
        RECT 84.900 142.180 85.190 142.225 ;
        RECT 81.230 142.040 85.190 142.180 ;
        RECT 94.160 142.180 94.300 142.675 ;
        RECT 95.450 142.660 95.770 142.720 ;
        RECT 95.925 142.520 96.215 142.565 ;
        RECT 96.830 142.520 97.150 142.580 ;
        RECT 95.925 142.380 97.150 142.520 ;
        RECT 95.925 142.335 96.215 142.380 ;
        RECT 96.830 142.320 97.150 142.380 ;
        RECT 96.370 142.180 96.690 142.240 ;
        RECT 97.840 142.180 97.980 143.060 ;
        RECT 98.225 142.675 98.515 142.905 ;
        RECT 98.685 142.860 98.975 142.905 ;
        RECT 99.130 142.860 99.450 142.920 ;
        RECT 104.280 142.905 104.420 143.060 ;
        RECT 109.250 143.060 119.215 143.200 ;
        RECT 109.250 143.000 109.570 143.060 ;
        RECT 118.925 143.015 119.215 143.060 ;
        RECT 125.810 143.200 126.130 143.260 ;
        RECT 142.845 143.200 143.135 143.245 ;
        RECT 143.750 143.200 144.070 143.260 ;
        RECT 155.250 143.200 155.570 143.260 ;
        RECT 125.810 143.060 142.140 143.200 ;
        RECT 125.810 143.000 126.130 143.060 ;
        RECT 98.685 142.720 99.450 142.860 ;
        RECT 98.685 142.675 98.975 142.720 ;
        RECT 98.300 142.520 98.440 142.675 ;
        RECT 99.130 142.660 99.450 142.720 ;
        RECT 99.605 142.860 99.895 142.905 ;
        RECT 101.445 142.860 101.735 142.905 ;
        RECT 99.605 142.720 101.735 142.860 ;
        RECT 99.605 142.675 99.895 142.720 ;
        RECT 101.445 142.675 101.735 142.720 ;
        RECT 104.205 142.675 104.495 142.905 ;
        RECT 104.650 142.860 104.970 142.920 ;
        RECT 105.125 142.860 105.415 142.905 ;
        RECT 104.650 142.720 105.415 142.860 ;
        RECT 104.650 142.660 104.970 142.720 ;
        RECT 105.125 142.675 105.415 142.720 ;
        RECT 108.805 142.675 109.095 142.905 ;
        RECT 109.725 142.860 110.015 142.905 ;
        RECT 111.090 142.860 111.410 142.920 ;
        RECT 109.725 142.720 111.410 142.860 ;
        RECT 109.725 142.675 110.015 142.720 ;
        RECT 108.880 142.520 109.020 142.675 ;
        RECT 111.090 142.660 111.410 142.720 ;
        RECT 115.690 142.660 116.010 142.920 ;
        RECT 118.005 142.675 118.295 142.905 ;
        RECT 118.450 142.860 118.770 142.920 ;
        RECT 119.370 142.860 119.690 142.920 ;
        RECT 118.450 142.720 119.690 142.860 ;
        RECT 111.550 142.520 111.870 142.580 ;
        RECT 118.080 142.520 118.220 142.675 ;
        RECT 118.450 142.660 118.770 142.720 ;
        RECT 119.370 142.660 119.690 142.720 ;
        RECT 119.845 142.860 120.135 142.905 ;
        RECT 121.670 142.860 121.990 142.920 ;
        RECT 119.845 142.720 121.990 142.860 ;
        RECT 119.845 142.675 120.135 142.720 ;
        RECT 121.670 142.660 121.990 142.720 ;
        RECT 124.890 142.860 125.210 142.920 ;
        RECT 126.975 142.860 127.265 142.905 ;
        RECT 124.890 142.720 127.265 142.860 ;
        RECT 124.890 142.660 125.210 142.720 ;
        RECT 126.975 142.675 127.265 142.720 ;
        RECT 127.650 142.660 127.970 142.920 ;
        RECT 128.110 142.660 128.430 142.920 ;
        RECT 128.815 142.905 128.955 143.060 ;
        RECT 128.765 142.675 129.055 142.905 ;
        RECT 129.490 142.660 129.810 142.920 ;
        RECT 130.870 142.905 131.190 142.920 ;
        RECT 129.965 142.675 130.255 142.905 ;
        RECT 130.735 142.675 131.190 142.905 ;
        RECT 98.300 142.380 99.360 142.520 ;
        RECT 108.880 142.380 118.220 142.520 ;
        RECT 130.040 142.520 130.180 142.675 ;
        RECT 130.870 142.660 131.190 142.675 ;
        RECT 139.610 142.905 139.930 142.920 ;
        RECT 139.610 142.860 139.960 142.905 ;
        RECT 142.000 142.860 142.140 143.060 ;
        RECT 142.845 143.060 144.070 143.200 ;
        RECT 142.845 143.015 143.135 143.060 ;
        RECT 143.750 143.000 144.070 143.060 ;
        RECT 149.360 143.060 155.570 143.200 ;
        RECT 143.290 142.860 143.610 142.920 ;
        RECT 148.350 142.860 148.670 142.920 ;
        RECT 139.610 142.720 140.125 142.860 ;
        RECT 142.000 142.720 148.670 142.860 ;
        RECT 139.610 142.675 139.960 142.720 ;
        RECT 139.610 142.660 139.930 142.675 ;
        RECT 143.290 142.660 143.610 142.720 ;
        RECT 148.350 142.660 148.670 142.720 ;
        RECT 148.810 142.660 149.130 142.920 ;
        RECT 136.415 142.520 136.705 142.565 ;
        RECT 138.935 142.520 139.225 142.565 ;
        RECT 140.125 142.520 140.415 142.565 ;
        RECT 130.040 142.380 130.410 142.520 ;
        RECT 94.160 142.040 97.980 142.180 ;
        RECT 81.230 141.995 81.520 142.040 ;
        RECT 83.330 141.995 83.620 142.040 ;
        RECT 84.900 141.995 85.190 142.040 ;
        RECT 96.370 141.980 96.690 142.040 ;
        RECT 49.005 141.840 49.295 141.885 ;
        RECT 48.070 141.700 49.295 141.840 ;
        RECT 48.070 141.640 48.390 141.700 ;
        RECT 49.005 141.655 49.295 141.700 ;
        RECT 49.925 141.655 50.215 141.885 ;
        RECT 52.210 141.640 52.530 141.900 ;
        RECT 53.145 141.840 53.435 141.885 ;
        RECT 55.445 141.840 55.735 141.885 ;
        RECT 60.490 141.840 60.810 141.900 ;
        RECT 53.145 141.700 60.810 141.840 ;
        RECT 53.145 141.655 53.435 141.700 ;
        RECT 55.445 141.655 55.735 141.700 ;
        RECT 60.490 141.640 60.810 141.700 ;
        RECT 65.090 141.840 65.410 141.900 ;
        RECT 66.025 141.840 66.315 141.885 ;
        RECT 65.090 141.700 66.315 141.840 ;
        RECT 65.090 141.640 65.410 141.700 ;
        RECT 66.025 141.655 66.315 141.700 ;
        RECT 93.610 141.840 93.930 141.900 ;
        RECT 95.465 141.840 95.755 141.885 ;
        RECT 93.610 141.700 95.755 141.840 ;
        RECT 93.610 141.640 93.930 141.700 ;
        RECT 95.465 141.655 95.755 141.700 ;
        RECT 96.845 141.840 97.135 141.885 ;
        RECT 98.670 141.840 98.990 141.900 ;
        RECT 99.220 141.885 99.360 142.380 ;
        RECT 111.550 142.320 111.870 142.380 ;
        RECT 130.270 142.240 130.410 142.380 ;
        RECT 136.415 142.380 140.415 142.520 ;
        RECT 136.415 142.335 136.705 142.380 ;
        RECT 138.935 142.335 139.225 142.380 ;
        RECT 140.125 142.335 140.415 142.380 ;
        RECT 141.005 142.520 141.295 142.565 ;
        RECT 149.360 142.520 149.500 143.060 ;
        RECT 155.250 143.000 155.570 143.060 ;
        RECT 149.730 142.860 150.050 142.920 ;
        RECT 150.205 142.860 150.495 142.905 ;
        RECT 149.730 142.720 150.495 142.860 ;
        RECT 149.730 142.660 150.050 142.720 ;
        RECT 150.205 142.675 150.495 142.720 ;
        RECT 150.650 142.860 150.970 142.920 ;
        RECT 151.125 142.860 151.415 142.905 ;
        RECT 150.650 142.720 151.415 142.860 ;
        RECT 150.650 142.660 150.970 142.720 ;
        RECT 151.125 142.675 151.415 142.720 ;
        RECT 152.030 142.660 152.350 142.920 ;
        RECT 141.005 142.380 149.500 142.520 ;
        RECT 141.005 142.335 141.295 142.380 ;
        RECT 104.190 142.180 104.510 142.240 ;
        RECT 116.610 142.180 116.930 142.240 ;
        RECT 104.190 142.040 116.930 142.180 ;
        RECT 130.270 142.040 130.730 142.240 ;
        RECT 104.190 141.980 104.510 142.040 ;
        RECT 116.610 141.980 116.930 142.040 ;
        RECT 130.410 141.980 130.730 142.040 ;
        RECT 131.805 142.180 132.095 142.225 ;
        RECT 132.250 142.180 132.570 142.240 ;
        RECT 134.550 142.180 134.870 142.240 ;
        RECT 131.805 142.040 134.870 142.180 ;
        RECT 131.805 141.995 132.095 142.040 ;
        RECT 132.250 141.980 132.570 142.040 ;
        RECT 134.550 141.980 134.870 142.040 ;
        RECT 136.850 142.180 137.140 142.225 ;
        RECT 138.420 142.180 138.710 142.225 ;
        RECT 140.520 142.180 140.810 142.225 ;
        RECT 136.850 142.040 140.810 142.180 ;
        RECT 136.850 141.995 137.140 142.040 ;
        RECT 138.420 141.995 138.710 142.040 ;
        RECT 140.520 141.995 140.810 142.040 ;
        RECT 144.225 142.180 144.515 142.225 ;
        RECT 144.670 142.180 144.990 142.240 ;
        RECT 144.225 142.040 144.990 142.180 ;
        RECT 144.225 141.995 144.515 142.040 ;
        RECT 144.670 141.980 144.990 142.040 ;
        RECT 145.130 142.180 145.450 142.240 ;
        RECT 145.605 142.180 145.895 142.225 ;
        RECT 148.825 142.180 149.115 142.225 ;
        RECT 145.130 142.040 149.115 142.180 ;
        RECT 145.130 141.980 145.450 142.040 ;
        RECT 145.605 141.995 145.895 142.040 ;
        RECT 148.825 141.995 149.115 142.040 ;
        RECT 96.845 141.700 98.990 141.840 ;
        RECT 96.845 141.655 97.135 141.700 ;
        RECT 98.670 141.640 98.990 141.700 ;
        RECT 99.145 141.840 99.435 141.885 ;
        RECT 103.730 141.840 104.050 141.900 ;
        RECT 99.145 141.700 104.050 141.840 ;
        RECT 99.145 141.655 99.435 141.700 ;
        RECT 103.730 141.640 104.050 141.700 ;
        RECT 106.045 141.840 106.335 141.885 ;
        RECT 107.870 141.840 108.190 141.900 ;
        RECT 106.045 141.700 108.190 141.840 ;
        RECT 106.045 141.655 106.335 141.700 ;
        RECT 107.870 141.640 108.190 141.700 ;
        RECT 117.085 141.840 117.375 141.885 ;
        RECT 117.530 141.840 117.850 141.900 ;
        RECT 117.085 141.700 117.850 141.840 ;
        RECT 117.085 141.655 117.375 141.700 ;
        RECT 117.530 141.640 117.850 141.700 ;
        RECT 141.450 141.640 141.770 141.900 ;
        RECT 147.430 141.640 147.750 141.900 ;
        RECT 148.365 141.840 148.655 141.885 ;
        RECT 152.030 141.840 152.350 141.900 ;
        RECT 148.365 141.700 152.350 141.840 ;
        RECT 148.365 141.655 148.655 141.700 ;
        RECT 152.030 141.640 152.350 141.700 ;
        RECT 22.700 141.020 157.020 141.500 ;
        RECT 26.450 140.620 26.770 140.880 ;
        RECT 27.370 140.620 27.690 140.880 ;
        RECT 31.050 140.620 31.370 140.880 ;
        RECT 34.285 140.820 34.575 140.865 ;
        RECT 33.670 140.680 34.575 140.820 ;
        RECT 27.460 140.140 27.600 140.620 ;
        RECT 29.210 140.280 29.530 140.540 ;
        RECT 31.985 140.480 32.275 140.525 ;
        RECT 32.430 140.480 32.750 140.540 ;
        RECT 31.985 140.340 32.750 140.480 ;
        RECT 31.985 140.295 32.275 140.340 ;
        RECT 32.430 140.280 32.750 140.340 ;
        RECT 33.670 140.200 33.810 140.680 ;
        RECT 34.285 140.635 34.575 140.680 ;
        RECT 35.190 140.620 35.510 140.880 ;
        RECT 36.110 140.620 36.430 140.880 ;
        RECT 44.865 140.820 45.155 140.865 ;
        RECT 45.770 140.820 46.090 140.880 ;
        RECT 44.865 140.680 46.090 140.820 ;
        RECT 44.865 140.635 45.155 140.680 ;
        RECT 45.770 140.620 46.090 140.680 ;
        RECT 46.230 140.820 46.550 140.880 ;
        RECT 49.005 140.820 49.295 140.865 ;
        RECT 51.290 140.820 51.610 140.880 ;
        RECT 46.230 140.680 47.840 140.820 ;
        RECT 46.230 140.620 46.550 140.680 ;
        RECT 33.350 140.140 33.810 140.200 ;
        RECT 27.460 140.000 33.810 140.140 ;
        RECT 33.350 139.940 33.670 140.000 ;
        RECT 36.200 139.800 36.340 140.620 ;
        RECT 38.870 140.480 39.160 140.525 ;
        RECT 40.440 140.480 40.730 140.525 ;
        RECT 42.540 140.480 42.830 140.525 ;
        RECT 47.150 140.480 47.470 140.540 ;
        RECT 38.870 140.340 42.830 140.480 ;
        RECT 38.870 140.295 39.160 140.340 ;
        RECT 40.440 140.295 40.730 140.340 ;
        RECT 42.540 140.295 42.830 140.340 ;
        RECT 45.860 140.340 47.470 140.480 ;
        RECT 47.700 140.480 47.840 140.680 ;
        RECT 49.005 140.680 51.610 140.820 ;
        RECT 49.005 140.635 49.295 140.680 ;
        RECT 51.290 140.620 51.610 140.680 ;
        RECT 54.065 140.820 54.355 140.865 ;
        RECT 63.250 140.820 63.570 140.880 ;
        RECT 54.065 140.680 63.570 140.820 ;
        RECT 54.065 140.635 54.355 140.680 ;
        RECT 54.140 140.480 54.280 140.635 ;
        RECT 63.250 140.620 63.570 140.680 ;
        RECT 82.110 140.820 82.430 140.880 ;
        RECT 83.045 140.820 83.335 140.865 ;
        RECT 82.110 140.680 83.335 140.820 ;
        RECT 82.110 140.620 82.430 140.680 ;
        RECT 83.045 140.635 83.335 140.680 ;
        RECT 96.830 140.820 97.150 140.880 ;
        RECT 103.270 140.820 103.590 140.880 ;
        RECT 96.830 140.680 103.590 140.820 ;
        RECT 96.830 140.620 97.150 140.680 ;
        RECT 103.270 140.620 103.590 140.680 ;
        RECT 110.170 140.820 110.490 140.880 ;
        RECT 121.685 140.820 121.975 140.865 ;
        RECT 110.170 140.680 121.975 140.820 ;
        RECT 110.170 140.620 110.490 140.680 ;
        RECT 121.685 140.635 121.975 140.680 ;
        RECT 128.585 140.820 128.875 140.865 ;
        RECT 130.410 140.820 130.730 140.880 ;
        RECT 128.585 140.680 130.730 140.820 ;
        RECT 128.585 140.635 128.875 140.680 ;
        RECT 130.410 140.620 130.730 140.680 ;
        RECT 47.700 140.340 54.280 140.480 ;
        RECT 56.810 140.480 57.100 140.525 ;
        RECT 58.380 140.480 58.670 140.525 ;
        RECT 60.480 140.480 60.770 140.525 ;
        RECT 56.810 140.340 60.770 140.480 ;
        RECT 45.860 140.185 46.000 140.340 ;
        RECT 47.150 140.280 47.470 140.340 ;
        RECT 56.810 140.295 57.100 140.340 ;
        RECT 58.380 140.295 58.670 140.340 ;
        RECT 60.480 140.295 60.770 140.340 ;
        RECT 64.210 140.480 64.500 140.525 ;
        RECT 66.310 140.480 66.600 140.525 ;
        RECT 67.880 140.480 68.170 140.525 ;
        RECT 64.210 140.340 68.170 140.480 ;
        RECT 64.210 140.295 64.500 140.340 ;
        RECT 66.310 140.295 66.600 140.340 ;
        RECT 67.880 140.295 68.170 140.340 ;
        RECT 89.050 140.480 89.340 140.525 ;
        RECT 91.150 140.480 91.440 140.525 ;
        RECT 92.720 140.480 93.010 140.525 ;
        RECT 89.050 140.340 93.010 140.480 ;
        RECT 89.050 140.295 89.340 140.340 ;
        RECT 91.150 140.295 91.440 140.340 ;
        RECT 92.720 140.295 93.010 140.340 ;
        RECT 95.465 140.480 95.755 140.525 ;
        RECT 95.910 140.480 96.230 140.540 ;
        RECT 95.465 140.340 96.230 140.480 ;
        RECT 95.465 140.295 95.755 140.340 ;
        RECT 95.910 140.280 96.230 140.340 ;
        RECT 96.370 140.480 96.690 140.540 ;
        RECT 101.445 140.480 101.735 140.525 ;
        RECT 96.370 140.340 101.735 140.480 ;
        RECT 96.370 140.280 96.690 140.340 ;
        RECT 101.445 140.295 101.735 140.340 ;
        RECT 104.190 140.480 104.480 140.525 ;
        RECT 105.760 140.480 106.050 140.525 ;
        RECT 107.860 140.480 108.150 140.525 ;
        RECT 109.710 140.480 110.030 140.540 ;
        RECT 114.810 140.480 115.100 140.525 ;
        RECT 116.910 140.480 117.200 140.525 ;
        RECT 118.480 140.480 118.770 140.525 ;
        RECT 104.190 140.340 108.150 140.480 ;
        RECT 104.190 140.295 104.480 140.340 ;
        RECT 105.760 140.295 106.050 140.340 ;
        RECT 107.860 140.295 108.150 140.340 ;
        RECT 108.420 140.340 114.540 140.480 ;
        RECT 38.435 140.140 38.725 140.185 ;
        RECT 40.955 140.140 41.245 140.185 ;
        RECT 42.145 140.140 42.435 140.185 ;
        RECT 38.435 140.000 42.435 140.140 ;
        RECT 38.435 139.955 38.725 140.000 ;
        RECT 40.955 139.955 41.245 140.000 ;
        RECT 42.145 139.955 42.435 140.000 ;
        RECT 45.785 139.955 46.075 140.185 ;
        RECT 46.690 140.140 47.010 140.200 ;
        RECT 49.465 140.140 49.755 140.185 ;
        RECT 52.670 140.140 52.990 140.200 ;
        RECT 46.690 140.000 52.990 140.140 ;
        RECT 46.690 139.940 47.010 140.000 ;
        RECT 49.465 139.955 49.755 140.000 ;
        RECT 52.670 139.940 52.990 140.000 ;
        RECT 56.375 140.140 56.665 140.185 ;
        RECT 58.895 140.140 59.185 140.185 ;
        RECT 60.085 140.140 60.375 140.185 ;
        RECT 56.375 140.000 60.375 140.140 ;
        RECT 56.375 139.955 56.665 140.000 ;
        RECT 58.895 139.955 59.185 140.000 ;
        RECT 60.085 139.955 60.375 140.000 ;
        RECT 64.605 140.140 64.895 140.185 ;
        RECT 65.795 140.140 66.085 140.185 ;
        RECT 68.315 140.140 68.605 140.185 ;
        RECT 64.605 140.000 68.605 140.140 ;
        RECT 64.605 139.955 64.895 140.000 ;
        RECT 65.795 139.955 66.085 140.000 ;
        RECT 68.315 139.955 68.605 140.000 ;
        RECT 75.685 140.140 75.975 140.185 ;
        RECT 77.050 140.140 77.370 140.200 ;
        RECT 88.090 140.140 88.410 140.200 ;
        RECT 75.685 140.000 77.370 140.140 ;
        RECT 75.685 139.955 75.975 140.000 ;
        RECT 77.050 139.940 77.370 140.000 ;
        RECT 84.040 140.000 88.410 140.140 ;
        RECT 33.670 139.660 36.340 139.800 ;
        RECT 41.630 139.845 41.950 139.860 ;
        RECT 41.630 139.800 41.980 139.845 ;
        RECT 41.630 139.660 42.145 139.800 ;
        RECT 27.385 139.460 27.675 139.505 ;
        RECT 29.670 139.460 29.990 139.520 ;
        RECT 27.385 139.320 29.990 139.460 ;
        RECT 27.385 139.275 27.675 139.320 ;
        RECT 29.670 139.260 29.990 139.320 ;
        RECT 30.145 139.460 30.435 139.505 ;
        RECT 33.670 139.460 33.810 139.660 ;
        RECT 41.630 139.615 41.980 139.660 ;
        RECT 43.025 139.615 43.315 139.845 ;
        RECT 41.630 139.600 41.950 139.615 ;
        RECT 30.145 139.320 33.810 139.460 ;
        RECT 30.145 139.275 30.435 139.320 ;
        RECT 34.270 139.260 34.590 139.520 ;
        RECT 43.100 139.460 43.240 139.615 ;
        RECT 44.390 139.600 44.710 139.860 ;
        RECT 44.850 139.800 45.170 139.860 ;
        RECT 47.165 139.800 47.455 139.845 ;
        RECT 44.850 139.660 47.455 139.800 ;
        RECT 44.850 139.600 45.170 139.660 ;
        RECT 47.165 139.615 47.455 139.660 ;
        RECT 48.070 139.600 48.390 139.860 ;
        RECT 52.210 139.600 52.530 139.860 ;
        RECT 53.130 139.600 53.450 139.860 ;
        RECT 53.605 139.800 53.895 139.845 ;
        RECT 57.730 139.800 58.050 139.860 ;
        RECT 53.605 139.660 58.050 139.800 ;
        RECT 53.605 139.615 53.895 139.660 ;
        RECT 57.730 139.600 58.050 139.660 ;
        RECT 60.965 139.800 61.255 139.845 ;
        RECT 61.870 139.800 62.190 139.860 ;
        RECT 65.090 139.845 65.410 139.860 ;
        RECT 63.725 139.800 64.015 139.845 ;
        RECT 65.060 139.800 65.410 139.845 ;
        RECT 71.085 139.800 71.375 139.845 ;
        RECT 60.965 139.660 64.015 139.800 ;
        RECT 64.895 139.660 65.410 139.800 ;
        RECT 60.965 139.615 61.255 139.660 ;
        RECT 61.870 139.600 62.190 139.660 ;
        RECT 63.725 139.615 64.015 139.660 ;
        RECT 65.060 139.615 65.410 139.660 ;
        RECT 65.090 139.600 65.410 139.615 ;
        RECT 70.700 139.660 71.375 139.800 ;
        RECT 50.370 139.460 50.690 139.520 ;
        RECT 43.100 139.320 50.690 139.460 ;
        RECT 50.370 139.260 50.690 139.320 ;
        RECT 58.190 139.460 58.510 139.520 ;
        RECT 59.630 139.460 59.920 139.505 ;
        RECT 58.190 139.320 59.920 139.460 ;
        RECT 58.190 139.260 58.510 139.320 ;
        RECT 59.630 139.275 59.920 139.320 ;
        RECT 70.700 139.180 70.840 139.660 ;
        RECT 71.085 139.615 71.375 139.660 ;
        RECT 75.210 139.600 75.530 139.860 ;
        RECT 84.040 139.845 84.180 140.000 ;
        RECT 88.090 139.940 88.410 140.000 ;
        RECT 89.445 140.140 89.735 140.185 ;
        RECT 90.635 140.140 90.925 140.185 ;
        RECT 93.155 140.140 93.445 140.185 ;
        RECT 89.445 140.000 93.445 140.140 ;
        RECT 89.445 139.955 89.735 140.000 ;
        RECT 90.635 139.955 90.925 140.000 ;
        RECT 93.155 139.955 93.445 140.000 ;
        RECT 98.670 139.940 98.990 140.200 ;
        RECT 108.420 140.185 108.560 140.340 ;
        RECT 109.710 140.280 110.030 140.340 ;
        RECT 103.755 140.140 104.045 140.185 ;
        RECT 106.275 140.140 106.565 140.185 ;
        RECT 107.465 140.140 107.755 140.185 ;
        RECT 103.755 140.000 107.755 140.140 ;
        RECT 103.755 139.955 104.045 140.000 ;
        RECT 106.275 139.955 106.565 140.000 ;
        RECT 107.465 139.955 107.755 140.000 ;
        RECT 108.345 139.955 108.635 140.185 ;
        RECT 83.965 139.615 84.255 139.845 ;
        RECT 85.330 139.600 85.650 139.860 ;
        RECT 87.630 139.800 87.950 139.860 ;
        RECT 88.565 139.800 88.855 139.845 ;
        RECT 104.190 139.800 104.510 139.860 ;
        RECT 87.630 139.660 88.855 139.800 ;
        RECT 87.630 139.600 87.950 139.660 ;
        RECT 88.565 139.615 88.855 139.660 ;
        RECT 89.100 139.660 104.510 139.800 ;
        RECT 83.490 139.460 83.810 139.520 ;
        RECT 89.100 139.460 89.240 139.660 ;
        RECT 104.190 139.600 104.510 139.660 ;
        RECT 107.065 139.800 107.355 139.845 ;
        RECT 107.870 139.800 108.190 139.860 ;
        RECT 107.065 139.660 108.190 139.800 ;
        RECT 107.065 139.615 107.355 139.660 ;
        RECT 107.870 139.600 108.190 139.660 ;
        RECT 109.725 139.800 110.015 139.845 ;
        RECT 110.170 139.800 110.490 139.860 ;
        RECT 109.725 139.660 110.490 139.800 ;
        RECT 109.725 139.615 110.015 139.660 ;
        RECT 110.170 139.600 110.490 139.660 ;
        RECT 111.550 139.600 111.870 139.860 ;
        RECT 114.400 139.845 114.540 140.340 ;
        RECT 114.810 140.340 118.770 140.480 ;
        RECT 114.810 140.295 115.100 140.340 ;
        RECT 116.910 140.295 117.200 140.340 ;
        RECT 118.480 140.295 118.770 140.340 ;
        RECT 148.850 140.480 149.140 140.525 ;
        RECT 150.950 140.480 151.240 140.525 ;
        RECT 152.520 140.480 152.810 140.525 ;
        RECT 148.850 140.340 152.810 140.480 ;
        RECT 148.850 140.295 149.140 140.340 ;
        RECT 150.950 140.295 151.240 140.340 ;
        RECT 152.520 140.295 152.810 140.340 ;
        RECT 115.205 140.140 115.495 140.185 ;
        RECT 116.395 140.140 116.685 140.185 ;
        RECT 118.915 140.140 119.205 140.185 ;
        RECT 115.205 140.000 119.205 140.140 ;
        RECT 115.205 139.955 115.495 140.000 ;
        RECT 116.395 139.955 116.685 140.000 ;
        RECT 118.915 139.955 119.205 140.000 ;
        RECT 127.650 140.140 127.970 140.200 ;
        RECT 139.625 140.140 139.915 140.185 ;
        RECT 127.650 140.000 139.915 140.140 ;
        RECT 127.650 139.940 127.970 140.000 ;
        RECT 139.625 139.955 139.915 140.000 ;
        RECT 149.245 140.140 149.535 140.185 ;
        RECT 150.435 140.140 150.725 140.185 ;
        RECT 152.955 140.140 153.245 140.185 ;
        RECT 149.245 140.000 153.245 140.140 ;
        RECT 149.245 139.955 149.535 140.000 ;
        RECT 150.435 139.955 150.725 140.000 ;
        RECT 152.955 139.955 153.245 140.000 ;
        RECT 114.325 139.800 114.615 139.845 ;
        RECT 114.770 139.800 115.090 139.860 ;
        RECT 114.325 139.660 116.380 139.800 ;
        RECT 114.325 139.615 114.615 139.660 ;
        RECT 114.770 139.600 115.090 139.660 ;
        RECT 116.240 139.520 116.380 139.660 ;
        RECT 124.890 139.600 125.210 139.860 ;
        RECT 127.190 139.600 127.510 139.860 ;
        RECT 131.330 139.800 131.650 139.860 ;
        RECT 133.645 139.800 133.935 139.845 ;
        RECT 131.330 139.660 133.935 139.800 ;
        RECT 131.330 139.600 131.650 139.660 ;
        RECT 133.645 139.615 133.935 139.660 ;
        RECT 134.550 139.800 134.870 139.860 ;
        RECT 135.485 139.800 135.775 139.845 ;
        RECT 134.550 139.660 135.775 139.800 ;
        RECT 134.550 139.600 134.870 139.660 ;
        RECT 135.485 139.615 135.775 139.660 ;
        RECT 135.930 139.600 136.250 139.860 ;
        RECT 140.085 139.615 140.375 139.845 ;
        RECT 140.530 139.800 140.850 139.860 ;
        RECT 141.005 139.800 141.295 139.845 ;
        RECT 140.530 139.660 141.295 139.800 ;
        RECT 83.490 139.320 89.240 139.460 ;
        RECT 89.900 139.460 90.190 139.505 ;
        RECT 95.925 139.460 96.215 139.505 ;
        RECT 89.900 139.320 96.215 139.460 ;
        RECT 83.490 139.260 83.810 139.320 ;
        RECT 89.900 139.275 90.190 139.320 ;
        RECT 95.925 139.275 96.215 139.320 ;
        RECT 109.250 139.460 109.570 139.520 ;
        RECT 110.645 139.460 110.935 139.505 ;
        RECT 109.250 139.320 110.935 139.460 ;
        RECT 109.250 139.260 109.570 139.320 ;
        RECT 110.645 139.275 110.935 139.320 ;
        RECT 111.090 139.460 111.410 139.520 ;
        RECT 112.010 139.460 112.330 139.520 ;
        RECT 115.550 139.460 115.840 139.505 ;
        RECT 111.090 139.320 112.330 139.460 ;
        RECT 111.090 139.260 111.410 139.320 ;
        RECT 112.010 139.260 112.330 139.320 ;
        RECT 112.560 139.320 115.840 139.460 ;
        RECT 29.210 139.120 29.530 139.180 ;
        RECT 31.145 139.120 31.435 139.165 ;
        RECT 29.210 138.980 31.435 139.120 ;
        RECT 29.210 138.920 29.530 138.980 ;
        RECT 31.145 138.935 31.435 138.980 ;
        RECT 40.710 139.120 41.030 139.180 ;
        RECT 46.690 139.120 47.010 139.180 ;
        RECT 40.710 138.980 47.010 139.120 ;
        RECT 40.710 138.920 41.030 138.980 ;
        RECT 46.690 138.920 47.010 138.980 ;
        RECT 47.150 139.120 47.470 139.180 ;
        RECT 47.625 139.120 47.915 139.165 ;
        RECT 47.150 138.980 47.915 139.120 ;
        RECT 47.150 138.920 47.470 138.980 ;
        RECT 47.625 138.935 47.915 138.980 ;
        RECT 51.305 139.120 51.595 139.165 ;
        RECT 51.750 139.120 52.070 139.180 ;
        RECT 51.305 138.980 52.070 139.120 ;
        RECT 51.305 138.935 51.595 138.980 ;
        RECT 51.750 138.920 52.070 138.980 ;
        RECT 70.610 138.920 70.930 139.180 ;
        RECT 71.530 138.920 71.850 139.180 ;
        RECT 73.370 138.920 73.690 139.180 ;
        RECT 82.570 139.120 82.890 139.180 ;
        RECT 84.885 139.120 85.175 139.165 ;
        RECT 87.170 139.120 87.490 139.180 ;
        RECT 82.570 138.980 87.490 139.120 ;
        RECT 82.570 138.920 82.890 138.980 ;
        RECT 84.885 138.935 85.175 138.980 ;
        RECT 87.170 138.920 87.490 138.980 ;
        RECT 89.010 139.120 89.330 139.180 ;
        RECT 104.190 139.120 104.510 139.180 ;
        RECT 106.030 139.120 106.350 139.180 ;
        RECT 112.560 139.165 112.700 139.320 ;
        RECT 115.550 139.275 115.840 139.320 ;
        RECT 116.150 139.260 116.470 139.520 ;
        RECT 128.585 139.460 128.875 139.505 ;
        RECT 129.950 139.460 130.270 139.520 ;
        RECT 137.770 139.460 138.090 139.520 ;
        RECT 128.585 139.320 130.270 139.460 ;
        RECT 128.585 139.275 128.875 139.320 ;
        RECT 129.950 139.260 130.270 139.320 ;
        RECT 135.100 139.320 138.090 139.460 ;
        RECT 140.160 139.460 140.300 139.615 ;
        RECT 140.530 139.600 140.850 139.660 ;
        RECT 141.005 139.615 141.295 139.660 ;
        RECT 145.130 139.600 145.450 139.860 ;
        RECT 148.350 139.600 148.670 139.860 ;
        RECT 144.670 139.460 144.990 139.520 ;
        RECT 146.065 139.460 146.355 139.505 ;
        RECT 149.700 139.460 149.990 139.505 ;
        RECT 150.190 139.460 150.510 139.520 ;
        RECT 140.160 139.320 147.660 139.460 ;
        RECT 89.010 138.980 106.350 139.120 ;
        RECT 89.010 138.920 89.330 138.980 ;
        RECT 104.190 138.920 104.510 138.980 ;
        RECT 106.030 138.920 106.350 138.980 ;
        RECT 112.485 138.935 112.775 139.165 ;
        RECT 121.225 139.120 121.515 139.165 ;
        RECT 124.890 139.120 125.210 139.180 ;
        RECT 121.225 138.980 125.210 139.120 ;
        RECT 121.225 138.935 121.515 138.980 ;
        RECT 124.890 138.920 125.210 138.980 ;
        RECT 127.665 139.120 127.955 139.165 ;
        RECT 131.790 139.120 132.110 139.180 ;
        RECT 135.100 139.165 135.240 139.320 ;
        RECT 137.770 139.260 138.090 139.320 ;
        RECT 144.670 139.260 144.990 139.320 ;
        RECT 146.065 139.275 146.355 139.320 ;
        RECT 127.665 138.980 132.110 139.120 ;
        RECT 127.665 138.935 127.955 138.980 ;
        RECT 131.790 138.920 132.110 138.980 ;
        RECT 135.025 138.935 135.315 139.165 ;
        RECT 141.910 139.120 142.230 139.180 ;
        RECT 144.225 139.120 144.515 139.165 ;
        RECT 141.910 138.980 144.515 139.120 ;
        RECT 141.910 138.920 142.230 138.980 ;
        RECT 144.225 138.935 144.515 138.980 ;
        RECT 146.510 139.120 146.830 139.180 ;
        RECT 146.985 139.120 147.275 139.165 ;
        RECT 146.510 138.980 147.275 139.120 ;
        RECT 147.520 139.120 147.660 139.320 ;
        RECT 149.700 139.320 150.510 139.460 ;
        RECT 149.700 139.275 149.990 139.320 ;
        RECT 150.190 139.260 150.510 139.320 ;
        RECT 155.265 139.120 155.555 139.165 ;
        RECT 147.520 138.980 155.555 139.120 ;
        RECT 146.510 138.920 146.830 138.980 ;
        RECT 146.985 138.935 147.275 138.980 ;
        RECT 155.265 138.935 155.555 138.980 ;
        RECT 22.700 138.300 157.820 138.780 ;
        RECT 27.830 138.100 28.150 138.160 ;
        RECT 31.970 138.100 32.290 138.160 ;
        RECT 27.830 137.960 32.290 138.100 ;
        RECT 27.830 137.900 28.150 137.960 ;
        RECT 31.600 137.465 31.740 137.960 ;
        RECT 31.970 137.900 32.290 137.960 ;
        RECT 33.350 138.100 33.670 138.160 ;
        RECT 41.630 138.100 41.950 138.160 ;
        RECT 33.350 137.960 41.950 138.100 ;
        RECT 33.350 137.900 33.670 137.960 ;
        RECT 41.630 137.900 41.950 137.960 ;
        RECT 44.405 138.100 44.695 138.145 ;
        RECT 44.850 138.100 45.170 138.160 ;
        RECT 44.405 137.960 45.170 138.100 ;
        RECT 44.405 137.915 44.695 137.960 ;
        RECT 44.850 137.900 45.170 137.960 ;
        RECT 47.150 137.900 47.470 138.160 ;
        RECT 57.270 137.900 57.590 138.160 ;
        RECT 58.190 137.900 58.510 138.160 ;
        RECT 60.030 137.900 60.350 138.160 ;
        RECT 68.325 138.100 68.615 138.145 ;
        RECT 70.610 138.100 70.930 138.160 ;
        RECT 68.325 137.960 70.930 138.100 ;
        RECT 68.325 137.915 68.615 137.960 ;
        RECT 70.610 137.900 70.930 137.960 ;
        RECT 71.070 137.900 71.390 138.160 ;
        RECT 76.590 138.100 76.910 138.160 ;
        RECT 77.525 138.100 77.815 138.145 ;
        RECT 76.590 137.960 77.815 138.100 ;
        RECT 76.590 137.900 76.910 137.960 ;
        RECT 77.525 137.915 77.815 137.960 ;
        RECT 83.950 138.100 84.270 138.160 ;
        RECT 84.755 138.100 85.045 138.145 ;
        RECT 88.550 138.100 88.870 138.160 ;
        RECT 89.945 138.100 90.235 138.145 ;
        RECT 92.230 138.100 92.550 138.160 ;
        RECT 83.950 137.960 90.235 138.100 ;
        RECT 83.950 137.900 84.270 137.960 ;
        RECT 84.755 137.915 85.045 137.960 ;
        RECT 88.550 137.900 88.870 137.960 ;
        RECT 89.945 137.915 90.235 137.960 ;
        RECT 90.940 137.960 92.550 138.100 ;
        RECT 34.590 137.760 34.880 137.805 ;
        RECT 57.360 137.760 57.500 137.900 ;
        RECT 90.940 137.820 91.080 137.960 ;
        RECT 92.230 137.900 92.550 137.960 ;
        RECT 96.370 138.100 96.690 138.160 ;
        RECT 102.365 138.100 102.655 138.145 ;
        RECT 103.825 138.100 104.115 138.145 ;
        RECT 96.370 137.960 101.660 138.100 ;
        RECT 96.370 137.900 96.690 137.960 ;
        RECT 32.060 137.620 34.880 137.760 ;
        RECT 31.525 137.235 31.815 137.465 ;
        RECT 30.605 137.080 30.895 137.125 ;
        RECT 32.060 137.080 32.200 137.620 ;
        RECT 34.590 137.575 34.880 137.620 ;
        RECT 44.940 137.620 57.500 137.760 ;
        RECT 57.730 137.760 58.050 137.820 ;
        RECT 68.785 137.760 69.075 137.805 ;
        RECT 73.370 137.760 73.690 137.820 ;
        RECT 83.490 137.760 83.810 137.820 ;
        RECT 57.730 137.620 60.720 137.760 ;
        RECT 32.430 137.220 32.750 137.480 ;
        RECT 32.905 137.420 33.195 137.465 ;
        RECT 36.570 137.420 36.890 137.480 ;
        RECT 44.940 137.465 45.080 137.620 ;
        RECT 57.730 137.560 58.050 137.620 ;
        RECT 32.905 137.280 36.890 137.420 ;
        RECT 32.905 137.235 33.195 137.280 ;
        RECT 36.570 137.220 36.890 137.280 ;
        RECT 42.105 137.420 42.395 137.465 ;
        RECT 42.105 137.280 44.620 137.420 ;
        RECT 42.105 137.235 42.395 137.280 ;
        RECT 30.605 136.940 32.200 137.080 ;
        RECT 30.605 136.895 30.895 136.940 ;
        RECT 33.365 136.895 33.655 137.125 ;
        RECT 34.245 137.080 34.535 137.125 ;
        RECT 35.435 137.080 35.725 137.125 ;
        RECT 37.955 137.080 38.245 137.125 ;
        RECT 34.245 136.940 38.245 137.080 ;
        RECT 44.480 137.080 44.620 137.280 ;
        RECT 44.865 137.235 45.155 137.465 ;
        RECT 46.230 137.420 46.550 137.480 ;
        RECT 45.400 137.280 46.550 137.420 ;
        RECT 45.400 137.080 45.540 137.280 ;
        RECT 46.230 137.220 46.550 137.280 ;
        RECT 50.370 137.220 50.690 137.480 ;
        RECT 51.750 137.465 52.070 137.480 ;
        RECT 51.720 137.420 52.070 137.465 ;
        RECT 51.555 137.280 52.070 137.420 ;
        RECT 51.720 137.235 52.070 137.280 ;
        RECT 51.750 137.220 52.070 137.235 ;
        RECT 53.130 137.420 53.450 137.480 ;
        RECT 54.050 137.420 54.370 137.480 ;
        RECT 53.130 137.280 58.880 137.420 ;
        RECT 53.130 137.220 53.450 137.280 ;
        RECT 54.050 137.220 54.370 137.280 ;
        RECT 44.480 136.940 45.540 137.080 ;
        RECT 51.265 137.080 51.555 137.125 ;
        RECT 52.455 137.080 52.745 137.125 ;
        RECT 54.975 137.080 55.265 137.125 ;
        RECT 51.265 136.940 55.265 137.080 ;
        RECT 58.740 137.080 58.880 137.280 ;
        RECT 59.110 137.220 59.430 137.480 ;
        RECT 60.580 137.465 60.720 137.620 ;
        RECT 68.785 137.620 73.690 137.760 ;
        RECT 68.785 137.575 69.075 137.620 ;
        RECT 73.370 137.560 73.690 137.620 ;
        RECT 73.920 137.620 83.810 137.760 ;
        RECT 60.505 137.235 60.795 137.465 ;
        RECT 70.625 137.420 70.915 137.465 ;
        RECT 61.040 137.280 71.300 137.420 ;
        RECT 61.040 137.080 61.180 137.280 ;
        RECT 70.625 137.235 70.915 137.280 ;
        RECT 58.740 136.940 61.180 137.080 ;
        RECT 65.550 137.080 65.870 137.140 ;
        RECT 69.245 137.080 69.535 137.125 ;
        RECT 65.550 136.940 69.535 137.080 ;
        RECT 71.160 137.080 71.300 137.280 ;
        RECT 71.530 137.220 71.850 137.480 ;
        RECT 73.920 137.420 74.060 137.620 ;
        RECT 83.490 137.560 83.810 137.620 ;
        RECT 85.805 137.760 86.095 137.805 ;
        RECT 86.265 137.760 86.555 137.805 ;
        RECT 85.805 137.620 86.555 137.760 ;
        RECT 85.805 137.575 86.095 137.620 ;
        RECT 86.265 137.575 86.555 137.620 ;
        RECT 90.850 137.560 91.170 137.820 ;
        RECT 92.705 137.760 92.995 137.805 ;
        RECT 99.130 137.760 99.450 137.820 ;
        RECT 101.520 137.805 101.660 137.960 ;
        RECT 102.365 137.960 104.115 138.100 ;
        RECT 102.365 137.915 102.655 137.960 ;
        RECT 103.825 137.915 104.115 137.960 ;
        RECT 104.650 137.900 104.970 138.160 ;
        RECT 105.585 138.100 105.875 138.145 ;
        RECT 108.330 138.100 108.650 138.160 ;
        RECT 111.550 138.100 111.870 138.160 ;
        RECT 105.585 137.960 111.870 138.100 ;
        RECT 105.585 137.915 105.875 137.960 ;
        RECT 108.330 137.900 108.650 137.960 ;
        RECT 111.550 137.900 111.870 137.960 ;
        RECT 113.405 138.100 113.695 138.145 ;
        RECT 113.405 137.960 117.300 138.100 ;
        RECT 113.405 137.915 113.695 137.960 ;
        RECT 100.525 137.760 100.815 137.805 ;
        RECT 92.705 137.620 94.760 137.760 ;
        RECT 92.705 137.575 92.995 137.620 ;
        RECT 72.080 137.280 74.060 137.420 ;
        RECT 72.080 137.080 72.220 137.280 ;
        RECT 77.050 137.220 77.370 137.480 ;
        RECT 88.090 137.420 88.410 137.480 ;
        RECT 91.785 137.420 92.075 137.465 ;
        RECT 88.090 137.280 92.075 137.420 ;
        RECT 88.090 137.220 88.410 137.280 ;
        RECT 91.785 137.235 92.075 137.280 ;
        RECT 92.230 137.220 92.550 137.480 ;
        RECT 93.610 137.220 93.930 137.480 ;
        RECT 94.620 137.465 94.760 137.620 ;
        RECT 99.130 137.620 100.815 137.760 ;
        RECT 99.130 137.560 99.450 137.620 ;
        RECT 100.525 137.575 100.815 137.620 ;
        RECT 101.445 137.575 101.735 137.805 ;
        RECT 102.825 137.760 103.115 137.805 ;
        RECT 103.270 137.760 103.590 137.820 ;
        RECT 109.710 137.760 110.030 137.820 ;
        RECT 102.825 137.620 103.590 137.760 ;
        RECT 102.825 137.575 103.115 137.620 ;
        RECT 103.270 137.560 103.590 137.620 ;
        RECT 106.580 137.620 110.030 137.760 ;
        RECT 94.545 137.235 94.835 137.465 ;
        RECT 95.005 137.420 95.295 137.465 ;
        RECT 95.910 137.420 96.230 137.480 ;
        RECT 95.005 137.280 96.230 137.420 ;
        RECT 95.005 137.235 95.295 137.280 ;
        RECT 95.910 137.220 96.230 137.280 ;
        RECT 96.370 137.220 96.690 137.480 ;
        RECT 97.750 137.220 98.070 137.480 ;
        RECT 99.590 137.420 99.910 137.480 ;
        RECT 99.220 137.280 99.910 137.420 ;
        RECT 71.160 136.940 72.220 137.080 ;
        RECT 75.670 137.080 75.990 137.140 ;
        RECT 77.985 137.080 78.275 137.125 ;
        RECT 75.670 136.940 78.275 137.080 ;
        RECT 34.245 136.895 34.535 136.940 ;
        RECT 35.435 136.895 35.725 136.940 ;
        RECT 37.955 136.895 38.245 136.940 ;
        RECT 51.265 136.895 51.555 136.940 ;
        RECT 52.455 136.895 52.745 136.940 ;
        RECT 54.975 136.895 55.265 136.940 ;
        RECT 32.890 136.740 33.210 136.800 ;
        RECT 33.440 136.740 33.580 136.895 ;
        RECT 65.550 136.880 65.870 136.940 ;
        RECT 69.245 136.895 69.535 136.940 ;
        RECT 75.670 136.880 75.990 136.940 ;
        RECT 77.985 136.895 78.275 136.940 ;
        RECT 89.010 136.880 89.330 137.140 ;
        RECT 95.450 136.880 95.770 137.140 ;
        RECT 99.220 137.125 99.360 137.280 ;
        RECT 99.590 137.220 99.910 137.280 ;
        RECT 102.350 137.420 102.670 137.480 ;
        RECT 105.125 137.420 105.415 137.465 ;
        RECT 102.350 137.280 105.415 137.420 ;
        RECT 102.350 137.220 102.670 137.280 ;
        RECT 105.125 137.235 105.415 137.280 ;
        RECT 106.030 137.220 106.350 137.480 ;
        RECT 106.580 137.465 106.720 137.620 ;
        RECT 109.710 137.560 110.030 137.620 ;
        RECT 107.870 137.465 108.190 137.480 ;
        RECT 117.160 137.465 117.300 137.960 ;
        RECT 121.670 137.900 121.990 138.160 ;
        RECT 129.490 137.900 129.810 138.160 ;
        RECT 129.950 137.900 130.270 138.160 ;
        RECT 140.530 137.900 140.850 138.160 ;
        RECT 143.290 138.100 143.610 138.160 ;
        RECT 143.765 138.100 144.055 138.145 ;
        RECT 143.290 137.960 144.055 138.100 ;
        RECT 143.290 137.900 143.610 137.960 ;
        RECT 143.765 137.915 144.055 137.960 ;
        RECT 146.510 137.900 146.830 138.160 ;
        RECT 147.445 137.915 147.735 138.145 ;
        RECT 124.890 137.760 125.210 137.820 ;
        RECT 129.580 137.760 129.720 137.900 ;
        RECT 134.550 137.760 134.870 137.820 ;
        RECT 141.450 137.760 141.770 137.820 ;
        RECT 142.830 137.760 143.150 137.820 ;
        RECT 124.890 137.620 128.800 137.760 ;
        RECT 129.580 137.620 132.940 137.760 ;
        RECT 124.890 137.560 125.210 137.620 ;
        RECT 106.505 137.235 106.795 137.465 ;
        RECT 107.840 137.235 108.190 137.465 ;
        RECT 117.085 137.420 117.375 137.465 ;
        RECT 118.910 137.420 119.230 137.480 ;
        RECT 117.085 137.280 119.230 137.420 ;
        RECT 117.085 137.235 117.375 137.280 ;
        RECT 107.870 137.220 108.190 137.235 ;
        RECT 118.910 137.220 119.230 137.280 ;
        RECT 127.650 137.420 127.970 137.480 ;
        RECT 128.660 137.465 128.800 137.620 ;
        RECT 128.125 137.420 128.415 137.465 ;
        RECT 127.650 137.280 128.415 137.420 ;
        RECT 127.650 137.220 127.970 137.280 ;
        RECT 128.125 137.235 128.415 137.280 ;
        RECT 128.585 137.235 128.875 137.465 ;
        RECT 130.885 137.235 131.175 137.465 ;
        RECT 99.145 136.895 99.435 137.125 ;
        RECT 107.385 137.080 107.675 137.125 ;
        RECT 108.575 137.080 108.865 137.125 ;
        RECT 111.095 137.080 111.385 137.125 ;
        RECT 107.385 136.940 111.385 137.080 ;
        RECT 107.385 136.895 107.675 136.940 ;
        RECT 108.575 136.895 108.865 136.940 ;
        RECT 111.095 136.895 111.385 136.940 ;
        RECT 121.210 136.880 121.530 137.140 ;
        RECT 124.905 137.080 125.195 137.125 ;
        RECT 125.350 137.080 125.670 137.140 ;
        RECT 124.905 136.940 125.670 137.080 ;
        RECT 124.905 136.895 125.195 136.940 ;
        RECT 125.350 136.880 125.670 136.940 ;
        RECT 126.285 136.895 126.575 137.125 ;
        RECT 126.745 137.080 127.035 137.125 ;
        RECT 127.190 137.080 127.510 137.140 ;
        RECT 126.745 136.940 127.510 137.080 ;
        RECT 130.960 137.080 131.100 137.235 ;
        RECT 131.330 137.220 131.650 137.480 ;
        RECT 131.790 137.220 132.110 137.480 ;
        RECT 132.800 137.465 132.940 137.620 ;
        RECT 134.550 137.620 136.160 137.760 ;
        RECT 134.550 137.560 134.870 137.620 ;
        RECT 132.725 137.235 133.015 137.465 ;
        RECT 133.645 137.420 133.935 137.465 ;
        RECT 134.090 137.420 134.410 137.480 ;
        RECT 135.010 137.465 135.330 137.480 ;
        RECT 133.645 137.280 134.410 137.420 ;
        RECT 133.645 137.235 133.935 137.280 ;
        RECT 134.090 137.220 134.410 137.280 ;
        RECT 134.980 137.235 135.330 137.465 ;
        RECT 136.020 137.420 136.160 137.620 ;
        RECT 141.450 137.620 144.900 137.760 ;
        RECT 141.450 137.560 141.770 137.620 ;
        RECT 142.830 137.560 143.150 137.620 ;
        RECT 136.020 137.280 141.680 137.420 ;
        RECT 135.010 137.220 135.330 137.235 ;
        RECT 133.170 137.080 133.490 137.140 ;
        RECT 141.540 137.125 141.680 137.280 ;
        RECT 141.910 137.220 142.230 137.480 ;
        RECT 144.210 137.220 144.530 137.480 ;
        RECT 144.760 137.465 144.900 137.620 ;
        RECT 144.685 137.235 144.975 137.465 ;
        RECT 147.520 137.420 147.660 137.915 ;
        RECT 150.190 137.900 150.510 138.160 ;
        RECT 149.285 137.420 149.575 137.465 ;
        RECT 147.520 137.280 149.575 137.420 ;
        RECT 149.285 137.235 149.575 137.280 ;
        RECT 130.960 136.940 133.490 137.080 ;
        RECT 126.745 136.895 127.035 136.940 ;
        RECT 32.890 136.600 33.580 136.740 ;
        RECT 33.850 136.740 34.140 136.785 ;
        RECT 35.950 136.740 36.240 136.785 ;
        RECT 37.520 136.740 37.810 136.785 ;
        RECT 44.390 136.740 44.710 136.800 ;
        RECT 50.870 136.740 51.160 136.785 ;
        RECT 52.970 136.740 53.260 136.785 ;
        RECT 54.540 136.740 54.830 136.785 ;
        RECT 33.850 136.600 37.810 136.740 ;
        RECT 32.890 136.540 33.210 136.600 ;
        RECT 33.850 136.555 34.140 136.600 ;
        RECT 35.950 136.555 36.240 136.600 ;
        RECT 37.520 136.555 37.810 136.600 ;
        RECT 39.880 136.600 45.540 136.740 ;
        RECT 32.430 136.400 32.750 136.460 ;
        RECT 39.880 136.400 40.020 136.600 ;
        RECT 44.390 136.540 44.710 136.600 ;
        RECT 32.430 136.260 40.020 136.400 ;
        RECT 40.265 136.400 40.555 136.445 ;
        RECT 40.710 136.400 41.030 136.460 ;
        RECT 40.265 136.260 41.030 136.400 ;
        RECT 32.430 136.200 32.750 136.260 ;
        RECT 40.265 136.215 40.555 136.260 ;
        RECT 40.710 136.200 41.030 136.260 ;
        RECT 42.550 136.200 42.870 136.460 ;
        RECT 45.400 136.445 45.540 136.600 ;
        RECT 50.870 136.600 54.830 136.740 ;
        RECT 50.870 136.555 51.160 136.600 ;
        RECT 52.970 136.555 53.260 136.600 ;
        RECT 54.540 136.555 54.830 136.600 ;
        RECT 106.990 136.740 107.280 136.785 ;
        RECT 109.090 136.740 109.380 136.785 ;
        RECT 110.660 136.740 110.950 136.785 ;
        RECT 106.990 136.600 110.950 136.740 ;
        RECT 126.360 136.740 126.500 136.895 ;
        RECT 127.190 136.880 127.510 136.940 ;
        RECT 133.170 136.880 133.490 136.940 ;
        RECT 134.525 137.080 134.815 137.125 ;
        RECT 135.715 137.080 136.005 137.125 ;
        RECT 138.235 137.080 138.525 137.125 ;
        RECT 134.525 136.940 138.525 137.080 ;
        RECT 134.525 136.895 134.815 136.940 ;
        RECT 135.715 136.895 136.005 136.940 ;
        RECT 138.235 136.895 138.525 136.940 ;
        RECT 141.465 136.895 141.755 137.125 ;
        RECT 128.110 136.740 128.430 136.800 ;
        RECT 126.360 136.600 128.430 136.740 ;
        RECT 106.990 136.555 107.280 136.600 ;
        RECT 109.090 136.555 109.380 136.600 ;
        RECT 110.660 136.555 110.950 136.600 ;
        RECT 128.110 136.540 128.430 136.600 ;
        RECT 134.130 136.740 134.420 136.785 ;
        RECT 136.230 136.740 136.520 136.785 ;
        RECT 137.800 136.740 138.090 136.785 ;
        RECT 134.130 136.600 138.090 136.740 ;
        RECT 134.130 136.555 134.420 136.600 ;
        RECT 136.230 136.555 136.520 136.600 ;
        RECT 137.800 136.555 138.090 136.600 ;
        RECT 45.325 136.215 45.615 136.445 ;
        RECT 66.470 136.200 66.790 136.460 ;
        RECT 75.210 136.200 75.530 136.460 ;
        RECT 83.030 136.400 83.350 136.460 ;
        RECT 83.965 136.400 84.255 136.445 ;
        RECT 83.030 136.260 84.255 136.400 ;
        RECT 83.030 136.200 83.350 136.260 ;
        RECT 83.965 136.215 84.255 136.260 ;
        RECT 84.885 136.400 85.175 136.445 ;
        RECT 85.790 136.400 86.110 136.460 ;
        RECT 84.885 136.260 86.110 136.400 ;
        RECT 84.885 136.215 85.175 136.260 ;
        RECT 85.790 136.200 86.110 136.260 ;
        RECT 97.305 136.400 97.595 136.445 ;
        RECT 98.225 136.400 98.515 136.445 ;
        RECT 97.305 136.260 98.515 136.400 ;
        RECT 97.305 136.215 97.595 136.260 ;
        RECT 98.225 136.215 98.515 136.260 ;
        RECT 98.670 136.200 98.990 136.460 ;
        RECT 103.730 136.200 104.050 136.460 ;
        RECT 113.850 136.200 114.170 136.460 ;
        RECT 116.610 136.400 116.930 136.460 ;
        RECT 118.005 136.400 118.295 136.445 ;
        RECT 116.610 136.260 118.295 136.400 ;
        RECT 116.610 136.200 116.930 136.260 ;
        RECT 118.005 136.215 118.295 136.260 ;
        RECT 144.210 136.400 144.530 136.460 ;
        RECT 146.525 136.400 146.815 136.445 ;
        RECT 147.430 136.400 147.750 136.460 ;
        RECT 144.210 136.260 147.750 136.400 ;
        RECT 144.210 136.200 144.530 136.260 ;
        RECT 146.525 136.215 146.815 136.260 ;
        RECT 147.430 136.200 147.750 136.260 ;
        RECT 22.700 135.580 157.020 136.060 ;
        RECT 26.925 135.380 27.215 135.425 ;
        RECT 30.145 135.380 30.435 135.425 ;
        RECT 26.925 135.240 30.435 135.380 ;
        RECT 26.925 135.195 27.215 135.240 ;
        RECT 30.145 135.195 30.435 135.240 ;
        RECT 41.630 135.180 41.950 135.440 ;
        RECT 75.210 135.380 75.530 135.440 ;
        RECT 71.620 135.240 75.530 135.380 ;
        RECT 31.050 135.040 31.370 135.100 ;
        RECT 32.430 135.040 32.750 135.100 ;
        RECT 27.920 134.900 32.750 135.040 ;
        RECT 27.920 134.405 28.060 134.900 ;
        RECT 31.050 134.840 31.370 134.900 ;
        RECT 32.430 134.840 32.750 134.900 ;
        RECT 29.210 134.700 29.530 134.760 ;
        RECT 36.125 134.700 36.415 134.745 ;
        RECT 29.210 134.560 36.415 134.700 ;
        RECT 29.210 134.500 29.530 134.560 ;
        RECT 36.125 134.515 36.415 134.560 ;
        RECT 43.485 134.700 43.775 134.745 ;
        RECT 48.990 134.700 49.310 134.760 ;
        RECT 43.485 134.560 49.310 134.700 ;
        RECT 43.485 134.515 43.775 134.560 ;
        RECT 48.990 134.500 49.310 134.560 ;
        RECT 27.845 134.175 28.135 134.405 ;
        RECT 28.765 134.360 29.055 134.405 ;
        RECT 29.670 134.360 29.990 134.420 ;
        RECT 31.525 134.360 31.815 134.405 ;
        RECT 28.765 134.220 31.815 134.360 ;
        RECT 28.765 134.175 29.055 134.220 ;
        RECT 29.670 134.160 29.990 134.220 ;
        RECT 31.525 134.175 31.815 134.220 ;
        RECT 31.970 134.160 32.290 134.420 ;
        RECT 32.430 134.160 32.750 134.420 ;
        RECT 36.570 134.360 36.890 134.420 ;
        RECT 38.885 134.360 39.175 134.405 ;
        RECT 36.570 134.220 39.175 134.360 ;
        RECT 36.570 134.160 36.890 134.220 ;
        RECT 38.885 134.175 39.175 134.220 ;
        RECT 42.565 134.360 42.855 134.405 ;
        RECT 43.010 134.360 43.330 134.420 ;
        RECT 42.565 134.220 43.330 134.360 ;
        RECT 42.565 134.175 42.855 134.220 ;
        RECT 43.010 134.160 43.330 134.220 ;
        RECT 43.930 134.360 44.250 134.420 ;
        RECT 46.705 134.360 46.995 134.405 ;
        RECT 43.930 134.220 46.995 134.360 ;
        RECT 43.930 134.160 44.250 134.220 ;
        RECT 46.705 134.175 46.995 134.220 ;
        RECT 52.210 134.360 52.530 134.420 ;
        RECT 55.445 134.360 55.735 134.405 ;
        RECT 52.210 134.220 55.735 134.360 ;
        RECT 52.210 134.160 52.530 134.220 ;
        RECT 55.445 134.175 55.735 134.220 ;
        RECT 70.625 134.360 70.915 134.405 ;
        RECT 71.620 134.360 71.760 135.240 ;
        RECT 75.210 135.180 75.530 135.240 ;
        RECT 85.790 135.380 86.110 135.440 ;
        RECT 88.565 135.380 88.855 135.425 ;
        RECT 85.790 135.240 88.855 135.380 ;
        RECT 85.790 135.180 86.110 135.240 ;
        RECT 88.565 135.195 88.855 135.240 ;
        RECT 90.865 135.380 91.155 135.425 ;
        RECT 95.450 135.380 95.770 135.440 ;
        RECT 90.865 135.240 95.770 135.380 ;
        RECT 90.865 135.195 91.155 135.240 ;
        RECT 95.450 135.180 95.770 135.240 ;
        RECT 97.305 135.380 97.595 135.425 ;
        RECT 97.750 135.380 98.070 135.440 ;
        RECT 97.305 135.240 98.070 135.380 ;
        RECT 97.305 135.195 97.595 135.240 ;
        RECT 97.750 135.180 98.070 135.240 ;
        RECT 107.425 135.380 107.715 135.425 ;
        RECT 107.870 135.380 108.190 135.440 ;
        RECT 107.425 135.240 108.190 135.380 ;
        RECT 107.425 135.195 107.715 135.240 ;
        RECT 107.870 135.180 108.190 135.240 ;
        RECT 130.885 135.380 131.175 135.425 ;
        RECT 131.790 135.380 132.110 135.440 ;
        RECT 130.885 135.240 132.110 135.380 ;
        RECT 130.885 135.195 131.175 135.240 ;
        RECT 131.790 135.180 132.110 135.240 ;
        RECT 135.010 135.180 135.330 135.440 ;
        RECT 72.490 135.040 72.780 135.085 ;
        RECT 74.590 135.040 74.880 135.085 ;
        RECT 76.160 135.040 76.450 135.085 ;
        RECT 72.490 134.900 76.450 135.040 ;
        RECT 72.490 134.855 72.780 134.900 ;
        RECT 74.590 134.855 74.880 134.900 ;
        RECT 76.160 134.855 76.450 134.900 ;
        RECT 79.850 135.040 80.140 135.085 ;
        RECT 81.950 135.040 82.240 135.085 ;
        RECT 83.520 135.040 83.810 135.085 ;
        RECT 79.850 134.900 83.810 135.040 ;
        RECT 79.850 134.855 80.140 134.900 ;
        RECT 81.950 134.855 82.240 134.900 ;
        RECT 83.520 134.855 83.810 134.900 ;
        RECT 116.650 135.040 116.940 135.085 ;
        RECT 118.750 135.040 119.040 135.085 ;
        RECT 120.320 135.040 120.610 135.085 ;
        RECT 116.650 134.900 120.610 135.040 ;
        RECT 116.650 134.855 116.940 134.900 ;
        RECT 118.750 134.855 119.040 134.900 ;
        RECT 120.320 134.855 120.610 134.900 ;
        RECT 130.425 135.040 130.715 135.085 ;
        RECT 131.345 135.040 131.635 135.085 ;
        RECT 130.425 134.900 131.635 135.040 ;
        RECT 130.425 134.855 130.715 134.900 ;
        RECT 131.345 134.855 131.635 134.900 ;
        RECT 145.630 135.040 145.920 135.085 ;
        RECT 147.730 135.040 148.020 135.085 ;
        RECT 149.300 135.040 149.590 135.085 ;
        RECT 145.630 134.900 149.590 135.040 ;
        RECT 145.630 134.855 145.920 134.900 ;
        RECT 147.730 134.855 148.020 134.900 ;
        RECT 149.300 134.855 149.590 134.900 ;
        RECT 72.885 134.700 73.175 134.745 ;
        RECT 74.075 134.700 74.365 134.745 ;
        RECT 76.595 134.700 76.885 134.745 ;
        RECT 72.885 134.560 76.885 134.700 ;
        RECT 72.885 134.515 73.175 134.560 ;
        RECT 74.075 134.515 74.365 134.560 ;
        RECT 76.595 134.515 76.885 134.560 ;
        RECT 80.245 134.700 80.535 134.745 ;
        RECT 81.435 134.700 81.725 134.745 ;
        RECT 83.955 134.700 84.245 134.745 ;
        RECT 80.245 134.560 84.245 134.700 ;
        RECT 80.245 134.515 80.535 134.560 ;
        RECT 81.435 134.515 81.725 134.560 ;
        RECT 83.955 134.515 84.245 134.560 ;
        RECT 96.385 134.700 96.675 134.745 ;
        RECT 117.045 134.700 117.335 134.745 ;
        RECT 118.235 134.700 118.525 134.745 ;
        RECT 120.755 134.700 121.045 134.745 ;
        RECT 96.385 134.560 98.440 134.700 ;
        RECT 96.385 134.515 96.675 134.560 ;
        RECT 98.300 134.420 98.440 134.560 ;
        RECT 117.045 134.560 121.045 134.700 ;
        RECT 117.045 134.515 117.335 134.560 ;
        RECT 118.235 134.515 118.525 134.560 ;
        RECT 120.755 134.515 121.045 134.560 ;
        RECT 123.985 134.700 124.275 134.745 ;
        RECT 127.190 134.700 127.510 134.760 ;
        RECT 128.110 134.700 128.430 134.760 ;
        RECT 123.985 134.560 127.880 134.700 ;
        RECT 123.985 134.515 124.275 134.560 ;
        RECT 127.190 134.500 127.510 134.560 ;
        RECT 70.625 134.220 71.760 134.360 ;
        RECT 72.005 134.360 72.295 134.405 ;
        RECT 79.350 134.360 79.670 134.420 ;
        RECT 89.010 134.360 89.330 134.420 ;
        RECT 90.405 134.360 90.695 134.405 ;
        RECT 72.005 134.220 79.670 134.360 ;
        RECT 70.625 134.175 70.915 134.220 ;
        RECT 72.005 134.175 72.295 134.220 ;
        RECT 31.065 134.020 31.355 134.065 ;
        RECT 32.060 134.020 32.200 134.160 ;
        RECT 40.710 134.020 41.030 134.080 ;
        RECT 31.065 133.880 41.030 134.020 ;
        RECT 31.065 133.835 31.355 133.880 ;
        RECT 40.710 133.820 41.030 133.880 ;
        RECT 68.310 134.020 68.630 134.080 ;
        RECT 72.080 134.020 72.220 134.175 ;
        RECT 79.350 134.160 79.670 134.220 ;
        RECT 86.340 134.220 90.695 134.360 ;
        RECT 73.230 134.020 73.520 134.065 ;
        RECT 68.310 133.880 72.220 134.020 ;
        RECT 72.540 133.880 73.520 134.020 ;
        RECT 68.310 133.820 68.630 133.880 ;
        RECT 27.370 133.680 27.690 133.740 ;
        RECT 29.225 133.680 29.515 133.725 ;
        RECT 27.370 133.540 29.515 133.680 ;
        RECT 27.370 133.480 27.690 133.540 ;
        RECT 29.225 133.495 29.515 133.540 ;
        RECT 30.065 133.680 30.355 133.725 ;
        RECT 31.985 133.680 32.275 133.725 ;
        RECT 30.065 133.540 32.275 133.680 ;
        RECT 30.065 133.495 30.355 133.540 ;
        RECT 31.985 133.495 32.275 133.540 ;
        RECT 43.010 133.680 43.330 133.740 ;
        RECT 43.945 133.680 44.235 133.725 ;
        RECT 43.010 133.540 44.235 133.680 ;
        RECT 43.010 133.480 43.330 133.540 ;
        RECT 43.945 133.495 44.235 133.540 ;
        RECT 52.670 133.480 52.990 133.740 ;
        RECT 71.545 133.680 71.835 133.725 ;
        RECT 72.540 133.680 72.680 133.880 ;
        RECT 73.230 133.835 73.520 133.880 ;
        RECT 80.700 134.020 80.990 134.065 ;
        RECT 82.110 134.020 82.430 134.080 ;
        RECT 80.700 133.880 82.430 134.020 ;
        RECT 80.700 133.835 80.990 133.880 ;
        RECT 82.110 133.820 82.430 133.880 ;
        RECT 71.545 133.540 72.680 133.680 ;
        RECT 76.130 133.680 76.450 133.740 ;
        RECT 86.340 133.725 86.480 134.220 ;
        RECT 89.010 134.160 89.330 134.220 ;
        RECT 90.405 134.175 90.695 134.220 ;
        RECT 95.910 134.160 96.230 134.420 ;
        RECT 97.305 134.175 97.595 134.405 ;
        RECT 88.550 134.065 88.870 134.080 ;
        RECT 88.485 133.835 88.870 134.065 ;
        RECT 89.485 134.020 89.775 134.065 ;
        RECT 92.230 134.020 92.550 134.080 ;
        RECT 97.380 134.020 97.520 134.175 ;
        RECT 98.210 134.160 98.530 134.420 ;
        RECT 108.330 134.160 108.650 134.420 ;
        RECT 109.250 134.160 109.570 134.420 ;
        RECT 110.185 134.360 110.475 134.405 ;
        RECT 113.850 134.360 114.170 134.420 ;
        RECT 110.185 134.220 114.170 134.360 ;
        RECT 110.185 134.175 110.475 134.220 ;
        RECT 113.850 134.160 114.170 134.220 ;
        RECT 116.150 134.160 116.470 134.420 ;
        RECT 117.530 134.405 117.850 134.420 ;
        RECT 117.500 134.360 117.850 134.405 ;
        RECT 117.335 134.220 117.850 134.360 ;
        RECT 117.500 134.175 117.850 134.220 ;
        RECT 117.530 134.160 117.850 134.175 ;
        RECT 118.910 134.360 119.230 134.420 ;
        RECT 123.525 134.360 123.815 134.405 ;
        RECT 118.910 134.220 123.815 134.360 ;
        RECT 118.910 134.160 119.230 134.220 ;
        RECT 123.525 134.175 123.815 134.220 ;
        RECT 125.350 134.160 125.670 134.420 ;
        RECT 125.810 134.360 126.130 134.420 ;
        RECT 127.740 134.405 127.880 134.560 ;
        RECT 128.110 134.560 130.410 134.700 ;
        RECT 128.110 134.500 128.430 134.560 ;
        RECT 126.285 134.360 126.575 134.405 ;
        RECT 125.810 134.220 126.575 134.360 ;
        RECT 125.810 134.160 126.130 134.220 ;
        RECT 126.285 134.175 126.575 134.220 ;
        RECT 126.745 134.175 127.035 134.405 ;
        RECT 127.665 134.175 127.955 134.405 ;
        RECT 89.485 133.880 97.520 134.020 ;
        RECT 89.485 133.835 89.775 133.880 ;
        RECT 88.550 133.820 88.870 133.835 ;
        RECT 92.230 133.820 92.550 133.880 ;
        RECT 108.790 133.820 109.110 134.080 ;
        RECT 78.905 133.680 79.195 133.725 ;
        RECT 76.130 133.540 79.195 133.680 ;
        RECT 71.545 133.495 71.835 133.540 ;
        RECT 76.130 133.480 76.450 133.540 ;
        RECT 78.905 133.495 79.195 133.540 ;
        RECT 86.265 133.495 86.555 133.725 ;
        RECT 86.710 133.680 87.030 133.740 ;
        RECT 87.645 133.680 87.935 133.725 ;
        RECT 86.710 133.540 87.935 133.680 ;
        RECT 86.710 133.480 87.030 133.540 ;
        RECT 87.645 133.495 87.935 133.540 ;
        RECT 123.065 133.680 123.355 133.725 ;
        RECT 125.350 133.680 125.670 133.740 ;
        RECT 123.065 133.540 125.670 133.680 ;
        RECT 123.065 133.495 123.355 133.540 ;
        RECT 125.350 133.480 125.670 133.540 ;
        RECT 126.285 133.680 126.575 133.725 ;
        RECT 126.820 133.680 126.960 134.175 ;
        RECT 128.570 134.160 128.890 134.420 ;
        RECT 129.030 134.360 129.350 134.420 ;
        RECT 129.505 134.360 129.795 134.405 ;
        RECT 129.030 134.220 129.795 134.360 ;
        RECT 130.270 134.360 130.410 134.560 ;
        RECT 137.770 134.500 138.090 134.760 ;
        RECT 144.210 134.700 144.530 134.760 ;
        RECT 141.540 134.560 144.530 134.700 ;
        RECT 139.165 134.360 139.455 134.405 ;
        RECT 130.270 134.220 139.455 134.360 ;
        RECT 129.030 134.160 129.350 134.220 ;
        RECT 129.505 134.175 129.795 134.220 ;
        RECT 139.165 134.175 139.455 134.220 ;
        RECT 140.085 134.360 140.375 134.405 ;
        RECT 140.990 134.360 141.310 134.420 ;
        RECT 141.540 134.405 141.680 134.560 ;
        RECT 144.210 134.500 144.530 134.560 ;
        RECT 146.025 134.700 146.315 134.745 ;
        RECT 147.215 134.700 147.505 134.745 ;
        RECT 149.735 134.700 150.025 134.745 ;
        RECT 146.025 134.560 150.025 134.700 ;
        RECT 146.025 134.515 146.315 134.560 ;
        RECT 147.215 134.515 147.505 134.560 ;
        RECT 149.735 134.515 150.025 134.560 ;
        RECT 140.085 134.220 141.310 134.360 ;
        RECT 140.085 134.175 140.375 134.220 ;
        RECT 131.330 134.020 131.650 134.080 ;
        RECT 130.270 133.880 131.650 134.020 ;
        RECT 130.270 133.680 130.410 133.880 ;
        RECT 131.330 133.820 131.650 133.880 ;
        RECT 133.170 133.820 133.490 134.080 ;
        RECT 139.240 134.020 139.380 134.175 ;
        RECT 140.990 134.160 141.310 134.220 ;
        RECT 141.465 134.175 141.755 134.405 ;
        RECT 142.370 134.160 142.690 134.420 ;
        RECT 142.830 134.160 143.150 134.420 ;
        RECT 143.290 134.160 143.610 134.420 ;
        RECT 145.145 134.360 145.435 134.405 ;
        RECT 148.350 134.360 148.670 134.420 ;
        RECT 145.145 134.220 148.670 134.360 ;
        RECT 145.145 134.175 145.435 134.220 ;
        RECT 148.350 134.160 148.670 134.220 ;
        RECT 144.685 134.020 144.975 134.065 ;
        RECT 146.370 134.020 146.660 134.065 ;
        RECT 139.240 133.880 143.060 134.020 ;
        RECT 126.285 133.540 130.410 133.680 ;
        RECT 141.005 133.680 141.295 133.725 ;
        RECT 141.910 133.680 142.230 133.740 ;
        RECT 141.005 133.540 142.230 133.680 ;
        RECT 142.920 133.680 143.060 133.880 ;
        RECT 144.685 133.880 146.660 134.020 ;
        RECT 144.685 133.835 144.975 133.880 ;
        RECT 146.370 133.835 146.660 133.880 ;
        RECT 151.110 133.680 151.430 133.740 ;
        RECT 152.045 133.680 152.335 133.725 ;
        RECT 142.920 133.540 152.335 133.680 ;
        RECT 126.285 133.495 126.575 133.540 ;
        RECT 141.005 133.495 141.295 133.540 ;
        RECT 141.910 133.480 142.230 133.540 ;
        RECT 151.110 133.480 151.430 133.540 ;
        RECT 152.045 133.495 152.335 133.540 ;
        RECT 22.700 132.860 157.820 133.340 ;
        RECT 28.765 132.660 29.055 132.705 ;
        RECT 28.765 132.520 30.360 132.660 ;
        RECT 28.765 132.475 29.055 132.520 ;
        RECT 26.925 131.980 27.215 132.025 ;
        RECT 27.370 131.980 27.690 132.040 ;
        RECT 26.925 131.840 27.690 131.980 ;
        RECT 26.925 131.795 27.215 131.840 ;
        RECT 27.370 131.780 27.690 131.840 ;
        RECT 28.290 131.780 28.610 132.040 ;
        RECT 29.210 131.780 29.530 132.040 ;
        RECT 30.220 131.980 30.360 132.520 ;
        RECT 36.570 132.460 36.890 132.720 ;
        RECT 52.210 132.460 52.530 132.720 ;
        RECT 52.685 132.660 52.975 132.705 ;
        RECT 54.970 132.660 55.290 132.720 ;
        RECT 65.105 132.660 65.395 132.705 ;
        RECT 52.685 132.520 57.500 132.660 ;
        RECT 52.685 132.475 52.975 132.520 ;
        RECT 54.970 132.460 55.290 132.520 ;
        RECT 37.950 132.320 38.270 132.380 ;
        RECT 39.190 132.320 39.480 132.365 ;
        RECT 37.950 132.180 39.480 132.320 ;
        RECT 37.950 132.120 38.270 132.180 ;
        RECT 39.190 132.135 39.480 132.180 ;
        RECT 50.830 132.320 51.150 132.380 ;
        RECT 57.360 132.320 57.500 132.520 ;
        RECT 64.260 132.520 65.395 132.660 ;
        RECT 63.725 132.320 64.015 132.365 ;
        RECT 50.830 132.180 53.360 132.320 ;
        RECT 57.360 132.180 64.015 132.320 ;
        RECT 50.830 132.120 51.150 132.180 ;
        RECT 30.965 131.980 31.255 132.025 ;
        RECT 30.220 131.840 31.255 131.980 ;
        RECT 30.965 131.795 31.255 131.840 ;
        RECT 32.890 131.980 33.210 132.040 ;
        RECT 45.310 131.980 45.630 132.040 ;
        RECT 53.220 132.025 53.360 132.180 ;
        RECT 63.725 132.135 64.015 132.180 ;
        RECT 46.245 131.980 46.535 132.025 ;
        RECT 32.890 131.840 38.180 131.980 ;
        RECT 32.890 131.780 33.210 131.840 ;
        RECT 38.040 131.685 38.180 131.840 ;
        RECT 45.310 131.840 46.535 131.980 ;
        RECT 45.310 131.780 45.630 131.840 ;
        RECT 46.245 131.795 46.535 131.840 ;
        RECT 53.145 131.795 53.435 132.025 ;
        RECT 54.525 131.795 54.815 132.025 ;
        RECT 56.365 131.980 56.655 132.025 ;
        RECT 60.950 131.980 61.270 132.040 ;
        RECT 56.365 131.840 61.270 131.980 ;
        RECT 56.365 131.795 56.655 131.840 ;
        RECT 29.685 131.640 29.975 131.685 ;
        RECT 27.000 131.500 29.975 131.640 ;
        RECT 27.000 131.360 27.140 131.500 ;
        RECT 29.685 131.455 29.975 131.500 ;
        RECT 30.565 131.640 30.855 131.685 ;
        RECT 31.755 131.640 32.045 131.685 ;
        RECT 34.275 131.640 34.565 131.685 ;
        RECT 30.565 131.500 34.565 131.640 ;
        RECT 30.565 131.455 30.855 131.500 ;
        RECT 31.755 131.455 32.045 131.500 ;
        RECT 34.275 131.455 34.565 131.500 ;
        RECT 37.965 131.455 38.255 131.685 ;
        RECT 38.845 131.640 39.135 131.685 ;
        RECT 40.035 131.640 40.325 131.685 ;
        RECT 42.555 131.640 42.845 131.685 ;
        RECT 38.845 131.500 42.845 131.640 ;
        RECT 38.845 131.455 39.135 131.500 ;
        RECT 40.035 131.455 40.325 131.500 ;
        RECT 42.555 131.455 42.845 131.500 ;
        RECT 50.845 131.640 51.135 131.685 ;
        RECT 51.290 131.640 51.610 131.700 ;
        RECT 50.845 131.500 51.610 131.640 ;
        RECT 50.845 131.455 51.135 131.500 ;
        RECT 26.910 131.100 27.230 131.360 ;
        RECT 25.990 130.760 26.310 131.020 ;
        RECT 29.760 130.960 29.900 131.455 ;
        RECT 30.170 131.300 30.460 131.345 ;
        RECT 32.270 131.300 32.560 131.345 ;
        RECT 33.840 131.300 34.130 131.345 ;
        RECT 30.170 131.160 34.130 131.300 ;
        RECT 30.170 131.115 30.460 131.160 ;
        RECT 32.270 131.115 32.560 131.160 ;
        RECT 33.840 131.115 34.130 131.160 ;
        RECT 32.890 130.960 33.210 131.020 ;
        RECT 29.760 130.820 33.210 130.960 ;
        RECT 38.040 130.960 38.180 131.455 ;
        RECT 51.290 131.440 51.610 131.500 ;
        RECT 54.065 131.455 54.355 131.685 ;
        RECT 54.600 131.640 54.740 131.795 ;
        RECT 60.950 131.780 61.270 131.840 ;
        RECT 61.425 131.980 61.715 132.025 ;
        RECT 64.260 131.980 64.400 132.520 ;
        RECT 65.105 132.475 65.395 132.520 ;
        RECT 66.945 132.660 67.235 132.705 ;
        RECT 71.530 132.660 71.850 132.720 ;
        RECT 66.945 132.520 71.850 132.660 ;
        RECT 66.945 132.475 67.235 132.520 ;
        RECT 71.530 132.460 71.850 132.520 ;
        RECT 77.050 132.660 77.370 132.720 ;
        RECT 77.985 132.660 78.275 132.705 ;
        RECT 77.050 132.520 78.275 132.660 ;
        RECT 77.050 132.460 77.370 132.520 ;
        RECT 77.985 132.475 78.275 132.520 ;
        RECT 82.110 132.460 82.430 132.720 ;
        RECT 85.345 132.660 85.635 132.705 ;
        RECT 92.230 132.660 92.550 132.720 ;
        RECT 94.545 132.660 94.835 132.705 ;
        RECT 85.345 132.520 92.000 132.660 ;
        RECT 85.345 132.475 85.635 132.520 ;
        RECT 64.645 132.320 64.935 132.365 ;
        RECT 66.470 132.320 66.790 132.380 ;
        RECT 83.965 132.320 84.255 132.365 ;
        RECT 64.645 132.180 66.790 132.320 ;
        RECT 64.645 132.135 64.935 132.180 ;
        RECT 66.470 132.120 66.790 132.180 ;
        RECT 82.200 132.180 84.255 132.320 ;
        RECT 82.200 132.040 82.340 132.180 ;
        RECT 83.965 132.135 84.255 132.180 ;
        RECT 87.185 132.320 87.475 132.365 ;
        RECT 88.870 132.320 89.160 132.365 ;
        RECT 87.185 132.180 89.160 132.320 ;
        RECT 91.860 132.320 92.000 132.520 ;
        RECT 92.230 132.520 94.835 132.660 ;
        RECT 92.230 132.460 92.550 132.520 ;
        RECT 94.545 132.475 94.835 132.520 ;
        RECT 108.330 132.660 108.650 132.720 ;
        RECT 108.330 132.520 114.540 132.660 ;
        RECT 108.330 132.460 108.650 132.520 ;
        RECT 102.810 132.320 103.130 132.380 ;
        RECT 107.425 132.320 107.715 132.365 ;
        RECT 91.860 132.180 103.130 132.320 ;
        RECT 87.185 132.135 87.475 132.180 ;
        RECT 88.870 132.135 89.160 132.180 ;
        RECT 102.810 132.120 103.130 132.180 ;
        RECT 104.280 132.180 107.715 132.320 ;
        RECT 104.280 132.040 104.420 132.180 ;
        RECT 107.425 132.135 107.715 132.180 ;
        RECT 109.250 132.320 109.570 132.380 ;
        RECT 113.865 132.320 114.155 132.365 ;
        RECT 109.250 132.180 114.155 132.320 ;
        RECT 114.400 132.320 114.540 132.520 ;
        RECT 115.705 132.475 115.995 132.705 ;
        RECT 121.210 132.660 121.530 132.720 ;
        RECT 123.065 132.660 123.355 132.705 ;
        RECT 121.210 132.520 123.355 132.660 ;
        RECT 115.780 132.320 115.920 132.475 ;
        RECT 121.210 132.460 121.530 132.520 ;
        RECT 123.065 132.475 123.355 132.520 ;
        RECT 129.950 132.660 130.270 132.720 ;
        RECT 133.170 132.660 133.490 132.720 ;
        RECT 129.950 132.520 133.490 132.660 ;
        RECT 117.390 132.320 117.680 132.365 ;
        RECT 114.400 132.180 115.000 132.320 ;
        RECT 115.780 132.180 117.680 132.320 ;
        RECT 123.140 132.320 123.280 132.475 ;
        RECT 129.950 132.460 130.270 132.520 ;
        RECT 133.170 132.460 133.490 132.520 ;
        RECT 135.025 132.660 135.315 132.705 ;
        RECT 135.930 132.660 136.250 132.720 ;
        RECT 141.005 132.660 141.295 132.705 ;
        RECT 135.025 132.520 141.295 132.660 ;
        RECT 135.025 132.475 135.315 132.520 ;
        RECT 135.930 132.460 136.250 132.520 ;
        RECT 141.005 132.475 141.295 132.520 ;
        RECT 142.370 132.660 142.690 132.720 ;
        RECT 143.305 132.660 143.595 132.705 ;
        RECT 142.370 132.520 143.595 132.660 ;
        RECT 142.370 132.460 142.690 132.520 ;
        RECT 143.305 132.475 143.595 132.520 ;
        RECT 123.140 132.180 128.340 132.320 ;
        RECT 109.250 132.120 109.570 132.180 ;
        RECT 113.865 132.135 114.155 132.180 ;
        RECT 76.130 131.980 76.450 132.040 ;
        RECT 61.425 131.840 64.400 131.980 ;
        RECT 65.640 131.840 76.450 131.980 ;
        RECT 61.425 131.795 61.715 131.840 ;
        RECT 65.640 131.700 65.780 131.840 ;
        RECT 76.130 131.780 76.450 131.840 ;
        RECT 77.065 131.795 77.355 132.025 ;
        RECT 65.550 131.640 65.870 131.700 ;
        RECT 54.600 131.500 65.870 131.640 ;
        RECT 38.450 131.300 38.740 131.345 ;
        RECT 40.550 131.300 40.840 131.345 ;
        RECT 42.120 131.300 42.410 131.345 ;
        RECT 54.140 131.300 54.280 131.455 ;
        RECT 65.550 131.440 65.870 131.500 ;
        RECT 66.010 131.640 66.330 131.700 ;
        RECT 67.405 131.640 67.695 131.685 ;
        RECT 66.010 131.500 67.695 131.640 ;
        RECT 66.010 131.440 66.330 131.500 ;
        RECT 67.405 131.455 67.695 131.500 ;
        RECT 67.865 131.640 68.155 131.685 ;
        RECT 76.590 131.640 76.910 131.700 ;
        RECT 67.865 131.500 76.910 131.640 ;
        RECT 77.140 131.640 77.280 131.795 ;
        RECT 82.110 131.780 82.430 132.040 ;
        RECT 83.030 131.780 83.350 132.040 ;
        RECT 84.425 131.980 84.715 132.025 ;
        RECT 84.870 131.980 85.190 132.040 ;
        RECT 84.425 131.840 85.190 131.980 ;
        RECT 84.425 131.795 84.715 131.840 ;
        RECT 84.870 131.780 85.190 131.840 ;
        RECT 86.265 131.980 86.555 132.025 ;
        RECT 86.710 131.980 87.030 132.040 ;
        RECT 86.265 131.840 87.030 131.980 ;
        RECT 86.265 131.795 86.555 131.840 ;
        RECT 86.710 131.780 87.030 131.840 ;
        RECT 87.630 131.780 87.950 132.040 ;
        RECT 88.180 131.840 97.520 131.980 ;
        RECT 77.510 131.640 77.830 131.700 ;
        RECT 88.180 131.640 88.320 131.840 ;
        RECT 77.140 131.500 88.320 131.640 ;
        RECT 88.525 131.640 88.815 131.685 ;
        RECT 89.715 131.640 90.005 131.685 ;
        RECT 92.235 131.640 92.525 131.685 ;
        RECT 88.525 131.500 92.525 131.640 ;
        RECT 67.865 131.455 68.155 131.500 ;
        RECT 67.940 131.300 68.080 131.455 ;
        RECT 76.590 131.440 76.910 131.500 ;
        RECT 77.510 131.440 77.830 131.500 ;
        RECT 88.525 131.455 88.815 131.500 ;
        RECT 89.715 131.455 90.005 131.500 ;
        RECT 92.235 131.455 92.525 131.500 ;
        RECT 95.910 131.640 96.230 131.700 ;
        RECT 96.845 131.640 97.135 131.685 ;
        RECT 95.910 131.500 97.135 131.640 ;
        RECT 97.380 131.640 97.520 131.840 ;
        RECT 97.750 131.780 98.070 132.040 ;
        RECT 104.190 131.780 104.510 132.040 ;
        RECT 105.110 131.980 105.430 132.040 ;
        RECT 105.585 131.980 105.875 132.025 ;
        RECT 106.505 131.980 106.795 132.025 ;
        RECT 105.110 131.840 106.795 131.980 ;
        RECT 105.110 131.780 105.430 131.840 ;
        RECT 105.585 131.795 105.875 131.840 ;
        RECT 106.505 131.795 106.795 131.840 ;
        RECT 112.945 131.795 113.235 132.025 ;
        RECT 113.390 131.980 113.710 132.040 ;
        RECT 114.860 132.025 115.000 132.180 ;
        RECT 117.390 132.135 117.680 132.180 ;
        RECT 114.325 131.980 114.615 132.025 ;
        RECT 113.390 131.840 114.615 131.980 ;
        RECT 109.710 131.640 110.030 131.700 ;
        RECT 97.380 131.500 110.030 131.640 ;
        RECT 113.020 131.640 113.160 131.795 ;
        RECT 113.390 131.780 113.710 131.840 ;
        RECT 114.325 131.795 114.615 131.840 ;
        RECT 114.785 131.795 115.075 132.025 ;
        RECT 116.150 131.780 116.470 132.040 ;
        RECT 116.610 131.780 116.930 132.040 ;
        RECT 125.350 131.980 125.670 132.040 ;
        RECT 127.665 131.980 127.955 132.025 ;
        RECT 125.350 131.840 127.955 131.980 ;
        RECT 128.200 131.980 128.340 132.180 ;
        RECT 129.030 132.120 129.350 132.380 ;
        RECT 130.410 132.120 130.730 132.380 ;
        RECT 133.630 132.320 133.950 132.380 ;
        RECT 134.565 132.320 134.855 132.365 ;
        RECT 133.630 132.180 134.855 132.320 ;
        RECT 133.630 132.120 133.950 132.180 ;
        RECT 134.565 132.135 134.855 132.180 ;
        RECT 129.965 131.985 130.255 132.025 ;
        RECT 129.580 131.980 130.255 131.985 ;
        RECT 128.200 131.845 130.255 131.980 ;
        RECT 128.200 131.840 129.720 131.845 ;
        RECT 125.350 131.780 125.670 131.840 ;
        RECT 127.665 131.795 127.955 131.840 ;
        RECT 129.965 131.795 130.255 131.845 ;
        RECT 132.250 131.980 132.570 132.040 ;
        RECT 134.105 131.980 134.395 132.025 ;
        RECT 132.250 131.840 134.395 131.980 ;
        RECT 132.250 131.780 132.570 131.840 ;
        RECT 134.105 131.795 134.395 131.840 ;
        RECT 136.405 131.980 136.695 132.025 ;
        RECT 140.545 131.980 140.835 132.025 ;
        RECT 141.005 131.980 141.295 132.025 ;
        RECT 136.405 131.840 141.295 131.980 ;
        RECT 136.405 131.795 136.695 131.840 ;
        RECT 140.545 131.795 140.835 131.840 ;
        RECT 141.005 131.795 141.295 131.840 ;
        RECT 141.910 131.780 142.230 132.040 ;
        RECT 142.830 131.780 143.150 132.040 ;
        RECT 143.290 131.980 143.610 132.040 ;
        RECT 143.765 131.980 144.055 132.025 ;
        RECT 143.290 131.840 144.055 131.980 ;
        RECT 143.290 131.780 143.610 131.840 ;
        RECT 143.765 131.795 144.055 131.840 ;
        RECT 144.670 131.980 144.990 132.040 ;
        RECT 145.605 131.980 145.895 132.025 ;
        RECT 144.670 131.840 145.895 131.980 ;
        RECT 116.700 131.640 116.840 131.780 ;
        RECT 113.020 131.500 116.840 131.640 ;
        RECT 117.045 131.640 117.335 131.685 ;
        RECT 118.235 131.640 118.525 131.685 ;
        RECT 120.755 131.640 121.045 131.685 ;
        RECT 117.045 131.500 121.045 131.640 ;
        RECT 95.910 131.440 96.230 131.500 ;
        RECT 96.845 131.455 97.135 131.500 ;
        RECT 109.710 131.440 110.030 131.500 ;
        RECT 117.045 131.455 117.335 131.500 ;
        RECT 118.235 131.455 118.525 131.500 ;
        RECT 120.755 131.455 121.045 131.500 ;
        RECT 125.810 131.640 126.130 131.700 ;
        RECT 127.205 131.640 127.495 131.685 ;
        RECT 125.810 131.500 127.495 131.640 ;
        RECT 125.810 131.440 126.130 131.500 ;
        RECT 127.205 131.455 127.495 131.500 ;
        RECT 128.570 131.640 128.890 131.700 ;
        RECT 129.505 131.640 129.795 131.685 ;
        RECT 128.570 131.500 129.795 131.640 ;
        RECT 38.450 131.160 42.410 131.300 ;
        RECT 38.450 131.115 38.740 131.160 ;
        RECT 40.550 131.115 40.840 131.160 ;
        RECT 42.120 131.115 42.410 131.160 ;
        RECT 44.940 131.160 54.280 131.300 ;
        RECT 54.600 131.160 68.080 131.300 ;
        RECT 88.130 131.300 88.420 131.345 ;
        RECT 90.230 131.300 90.520 131.345 ;
        RECT 91.800 131.300 92.090 131.345 ;
        RECT 88.130 131.160 92.090 131.300 ;
        RECT 42.550 130.960 42.870 131.020 ;
        RECT 38.040 130.820 42.870 130.960 ;
        RECT 32.890 130.760 33.210 130.820 ;
        RECT 42.550 130.760 42.870 130.820 ;
        RECT 43.930 130.960 44.250 131.020 ;
        RECT 44.940 131.005 45.080 131.160 ;
        RECT 44.865 130.960 45.155 131.005 ;
        RECT 43.930 130.820 45.155 130.960 ;
        RECT 43.930 130.760 44.250 130.820 ;
        RECT 44.865 130.775 45.155 130.820 ;
        RECT 45.325 130.960 45.615 131.005 ;
        RECT 45.770 130.960 46.090 131.020 ;
        RECT 45.325 130.820 46.090 130.960 ;
        RECT 45.325 130.775 45.615 130.820 ;
        RECT 45.770 130.760 46.090 130.820 ;
        RECT 48.990 130.960 49.310 131.020 ;
        RECT 51.290 130.960 51.610 131.020 ;
        RECT 54.600 130.960 54.740 131.160 ;
        RECT 88.130 131.115 88.420 131.160 ;
        RECT 90.230 131.115 90.520 131.160 ;
        RECT 91.800 131.115 92.090 131.160 ;
        RECT 105.585 131.300 105.875 131.345 ;
        RECT 107.870 131.300 108.190 131.360 ;
        RECT 105.585 131.160 108.190 131.300 ;
        RECT 105.585 131.115 105.875 131.160 ;
        RECT 107.870 131.100 108.190 131.160 ;
        RECT 116.650 131.300 116.940 131.345 ;
        RECT 118.750 131.300 119.040 131.345 ;
        RECT 120.320 131.300 120.610 131.345 ;
        RECT 116.650 131.160 120.610 131.300 ;
        RECT 127.280 131.300 127.420 131.455 ;
        RECT 128.570 131.440 128.890 131.500 ;
        RECT 129.505 131.455 129.795 131.500 ;
        RECT 137.785 131.640 138.075 131.685 ;
        RECT 138.230 131.640 138.550 131.700 ;
        RECT 137.785 131.500 138.550 131.640 ;
        RECT 137.785 131.455 138.075 131.500 ;
        RECT 138.230 131.440 138.550 131.500 ;
        RECT 134.550 131.300 134.870 131.360 ;
        RECT 127.280 131.160 134.870 131.300 ;
        RECT 116.650 131.115 116.940 131.160 ;
        RECT 118.750 131.115 119.040 131.160 ;
        RECT 120.320 131.115 120.610 131.160 ;
        RECT 134.550 131.100 134.870 131.160 ;
        RECT 135.945 131.300 136.235 131.345 ;
        RECT 142.000 131.300 142.140 131.780 ;
        RECT 143.840 131.640 143.980 131.795 ;
        RECT 144.670 131.780 144.990 131.840 ;
        RECT 145.605 131.795 145.895 131.840 ;
        RECT 146.525 131.980 146.815 132.025 ;
        RECT 152.950 131.980 153.270 132.040 ;
        RECT 146.525 131.840 153.270 131.980 ;
        RECT 146.525 131.795 146.815 131.840 ;
        RECT 152.950 131.780 153.270 131.840 ;
        RECT 147.905 131.640 148.195 131.685 ;
        RECT 143.840 131.500 148.195 131.640 ;
        RECT 147.905 131.455 148.195 131.500 ;
        RECT 151.110 131.440 151.430 131.700 ;
        RECT 154.790 131.440 155.110 131.700 ;
        RECT 135.945 131.160 142.140 131.300 ;
        RECT 147.445 131.300 147.735 131.345 ;
        RECT 153.870 131.300 154.190 131.360 ;
        RECT 147.445 131.160 154.190 131.300 ;
        RECT 135.945 131.115 136.235 131.160 ;
        RECT 147.445 131.115 147.735 131.160 ;
        RECT 153.870 131.100 154.190 131.160 ;
        RECT 48.990 130.820 54.740 130.960 ;
        RECT 48.990 130.760 49.310 130.820 ;
        RECT 51.290 130.760 51.610 130.820 ;
        RECT 55.890 130.760 56.210 131.020 ;
        RECT 57.285 130.960 57.575 131.005 ;
        RECT 58.650 130.960 58.970 131.020 ;
        RECT 57.285 130.820 58.970 130.960 ;
        RECT 57.285 130.775 57.575 130.820 ;
        RECT 58.650 130.760 58.970 130.820 ;
        RECT 62.330 130.760 62.650 131.020 ;
        RECT 62.805 130.960 63.095 131.005 ;
        RECT 63.710 130.960 64.030 131.020 ;
        RECT 62.805 130.820 64.030 130.960 ;
        RECT 62.805 130.775 63.095 130.820 ;
        RECT 63.710 130.760 64.030 130.820 ;
        RECT 98.685 130.960 98.975 131.005 ;
        RECT 103.270 130.960 103.590 131.020 ;
        RECT 105.110 130.960 105.430 131.020 ;
        RECT 98.685 130.820 105.430 130.960 ;
        RECT 98.685 130.775 98.975 130.820 ;
        RECT 103.270 130.760 103.590 130.820 ;
        RECT 105.110 130.760 105.430 130.820 ;
        RECT 108.345 130.960 108.635 131.005 ;
        RECT 114.310 130.960 114.630 131.020 ;
        RECT 108.345 130.820 114.630 130.960 ;
        RECT 108.345 130.775 108.635 130.820 ;
        RECT 114.310 130.760 114.630 130.820 ;
        RECT 126.285 130.960 126.575 131.005 ;
        RECT 129.950 130.960 130.270 131.020 ;
        RECT 126.285 130.820 130.270 130.960 ;
        RECT 126.285 130.775 126.575 130.820 ;
        RECT 129.950 130.760 130.270 130.820 ;
        RECT 132.710 130.760 133.030 131.020 ;
        RECT 152.045 130.960 152.335 131.005 ;
        RECT 153.410 130.960 153.730 131.020 ;
        RECT 152.045 130.820 153.730 130.960 ;
        RECT 152.045 130.775 152.335 130.820 ;
        RECT 153.410 130.760 153.730 130.820 ;
        RECT 22.700 130.140 157.020 130.620 ;
        RECT 31.065 129.940 31.355 129.985 ;
        RECT 32.430 129.940 32.750 130.000 ;
        RECT 31.065 129.800 32.750 129.940 ;
        RECT 31.065 129.755 31.355 129.800 ;
        RECT 32.430 129.740 32.750 129.800 ;
        RECT 37.950 129.940 38.270 130.000 ;
        RECT 40.265 129.940 40.555 129.985 ;
        RECT 37.950 129.800 40.555 129.940 ;
        RECT 37.950 129.740 38.270 129.800 ;
        RECT 40.265 129.755 40.555 129.800 ;
        RECT 50.845 129.940 51.135 129.985 ;
        RECT 54.510 129.940 54.830 130.000 ;
        RECT 55.890 129.940 56.210 130.000 ;
        RECT 50.845 129.800 56.210 129.940 ;
        RECT 50.845 129.755 51.135 129.800 ;
        RECT 54.510 129.740 54.830 129.800 ;
        RECT 55.890 129.740 56.210 129.800 ;
        RECT 60.490 129.940 60.810 130.000 ;
        RECT 84.425 129.940 84.715 129.985 ;
        RECT 84.870 129.940 85.190 130.000 ;
        RECT 60.490 129.800 82.110 129.940 ;
        RECT 60.490 129.740 60.810 129.800 ;
        RECT 24.650 129.600 24.940 129.645 ;
        RECT 26.750 129.600 27.040 129.645 ;
        RECT 28.320 129.600 28.610 129.645 ;
        RECT 24.650 129.460 28.610 129.600 ;
        RECT 24.650 129.415 24.940 129.460 ;
        RECT 26.750 129.415 27.040 129.460 ;
        RECT 28.320 129.415 28.610 129.460 ;
        RECT 44.430 129.600 44.720 129.645 ;
        RECT 46.530 129.600 46.820 129.645 ;
        RECT 48.100 129.600 48.390 129.645 ;
        RECT 44.430 129.460 48.390 129.600 ;
        RECT 44.430 129.415 44.720 129.460 ;
        RECT 46.530 129.415 46.820 129.460 ;
        RECT 48.100 129.415 48.390 129.460 ;
        RECT 51.790 129.600 52.080 129.645 ;
        RECT 53.890 129.600 54.180 129.645 ;
        RECT 55.460 129.600 55.750 129.645 ;
        RECT 51.790 129.460 55.750 129.600 ;
        RECT 51.790 129.415 52.080 129.460 ;
        RECT 53.890 129.415 54.180 129.460 ;
        RECT 55.460 129.415 55.750 129.460 ;
        RECT 62.370 129.600 62.660 129.645 ;
        RECT 64.470 129.600 64.760 129.645 ;
        RECT 66.040 129.600 66.330 129.645 ;
        RECT 62.370 129.460 66.330 129.600 ;
        RECT 62.370 129.415 62.660 129.460 ;
        RECT 64.470 129.415 64.760 129.460 ;
        RECT 66.040 129.415 66.330 129.460 ;
        RECT 69.730 129.600 70.020 129.645 ;
        RECT 71.830 129.600 72.120 129.645 ;
        RECT 73.400 129.600 73.690 129.645 ;
        RECT 69.730 129.460 73.690 129.600 ;
        RECT 69.730 129.415 70.020 129.460 ;
        RECT 71.830 129.415 72.120 129.460 ;
        RECT 73.400 129.415 73.690 129.460 ;
        RECT 76.145 129.600 76.435 129.645 ;
        RECT 81.970 129.600 82.110 129.800 ;
        RECT 84.425 129.800 85.190 129.940 ;
        RECT 84.425 129.755 84.715 129.800 ;
        RECT 84.870 129.740 85.190 129.800 ;
        RECT 129.030 129.940 129.350 130.000 ;
        RECT 138.230 129.940 138.550 130.000 ;
        RECT 129.030 129.800 138.550 129.940 ;
        RECT 129.030 129.740 129.350 129.800 ;
        RECT 138.230 129.740 138.550 129.800 ;
        RECT 151.570 129.940 151.890 130.000 ;
        RECT 154.790 129.940 155.110 130.000 ;
        RECT 155.265 129.940 155.555 129.985 ;
        RECT 151.570 129.800 155.555 129.940 ;
        RECT 151.570 129.740 151.890 129.800 ;
        RECT 154.790 129.740 155.110 129.800 ;
        RECT 155.265 129.755 155.555 129.800 ;
        RECT 94.070 129.600 94.390 129.660 ;
        RECT 76.145 129.460 76.820 129.600 ;
        RECT 81.970 129.460 94.390 129.600 ;
        RECT 76.145 129.415 76.435 129.460 ;
        RECT 25.045 129.260 25.335 129.305 ;
        RECT 26.235 129.260 26.525 129.305 ;
        RECT 28.755 129.260 29.045 129.305 ;
        RECT 25.045 129.120 29.045 129.260 ;
        RECT 25.045 129.075 25.335 129.120 ;
        RECT 26.235 129.075 26.525 129.120 ;
        RECT 28.755 129.075 29.045 129.120 ;
        RECT 40.710 129.260 41.030 129.320 ;
        RECT 40.710 129.120 41.860 129.260 ;
        RECT 40.710 129.060 41.030 129.120 ;
        RECT 24.165 128.920 24.455 128.965 ;
        RECT 26.910 128.920 27.230 128.980 ;
        RECT 41.720 128.965 41.860 129.120 ;
        RECT 43.010 129.060 43.330 129.320 ;
        RECT 43.470 129.060 43.790 129.320 ;
        RECT 76.680 129.305 76.820 129.460 ;
        RECT 94.070 129.400 94.390 129.460 ;
        RECT 98.710 129.600 99.000 129.645 ;
        RECT 100.810 129.600 101.100 129.645 ;
        RECT 102.380 129.600 102.670 129.645 ;
        RECT 98.710 129.460 102.670 129.600 ;
        RECT 98.710 129.415 99.000 129.460 ;
        RECT 100.810 129.415 101.100 129.460 ;
        RECT 102.380 129.415 102.670 129.460 ;
        RECT 131.830 129.600 132.120 129.645 ;
        RECT 133.930 129.600 134.220 129.645 ;
        RECT 135.500 129.600 135.790 129.645 ;
        RECT 131.830 129.460 135.790 129.600 ;
        RECT 131.830 129.415 132.120 129.460 ;
        RECT 133.930 129.415 134.220 129.460 ;
        RECT 135.500 129.415 135.790 129.460 ;
        RECT 148.850 129.600 149.140 129.645 ;
        RECT 150.950 129.600 151.240 129.645 ;
        RECT 152.520 129.600 152.810 129.645 ;
        RECT 148.850 129.460 152.810 129.600 ;
        RECT 148.850 129.415 149.140 129.460 ;
        RECT 150.950 129.415 151.240 129.460 ;
        RECT 152.520 129.415 152.810 129.460 ;
        RECT 44.825 129.260 45.115 129.305 ;
        RECT 46.015 129.260 46.305 129.305 ;
        RECT 48.535 129.260 48.825 129.305 ;
        RECT 44.825 129.120 48.825 129.260 ;
        RECT 44.825 129.075 45.115 129.120 ;
        RECT 46.015 129.075 46.305 129.120 ;
        RECT 48.535 129.075 48.825 129.120 ;
        RECT 52.185 129.260 52.475 129.305 ;
        RECT 53.375 129.260 53.665 129.305 ;
        RECT 55.895 129.260 56.185 129.305 ;
        RECT 52.185 129.120 56.185 129.260 ;
        RECT 52.185 129.075 52.475 129.120 ;
        RECT 53.375 129.075 53.665 129.120 ;
        RECT 55.895 129.075 56.185 129.120 ;
        RECT 62.765 129.260 63.055 129.305 ;
        RECT 63.955 129.260 64.245 129.305 ;
        RECT 66.475 129.260 66.765 129.305 ;
        RECT 62.765 129.120 66.765 129.260 ;
        RECT 62.765 129.075 63.055 129.120 ;
        RECT 63.955 129.075 64.245 129.120 ;
        RECT 66.475 129.075 66.765 129.120 ;
        RECT 70.125 129.260 70.415 129.305 ;
        RECT 71.315 129.260 71.605 129.305 ;
        RECT 73.835 129.260 74.125 129.305 ;
        RECT 70.125 129.120 74.125 129.260 ;
        RECT 70.125 129.075 70.415 129.120 ;
        RECT 71.315 129.075 71.605 129.120 ;
        RECT 73.835 129.075 74.125 129.120 ;
        RECT 76.605 129.075 76.895 129.305 ;
        RECT 81.650 129.260 81.970 129.320 ;
        RECT 88.090 129.260 88.410 129.320 ;
        RECT 81.280 129.120 83.720 129.260 ;
        RECT 24.165 128.780 27.230 128.920 ;
        RECT 24.165 128.735 24.455 128.780 ;
        RECT 26.910 128.720 27.230 128.780 ;
        RECT 41.185 128.735 41.475 128.965 ;
        RECT 41.645 128.735 41.935 128.965 ;
        RECT 42.550 128.920 42.870 128.980 ;
        RECT 43.945 128.920 44.235 128.965 ;
        RECT 50.370 128.920 50.690 128.980 ;
        RECT 52.670 128.965 52.990 128.980 ;
        RECT 51.305 128.920 51.595 128.965 ;
        RECT 52.640 128.920 52.990 128.965 ;
        RECT 42.550 128.780 51.595 128.920 ;
        RECT 52.475 128.780 52.990 128.920 ;
        RECT 25.500 128.580 25.790 128.625 ;
        RECT 25.990 128.580 26.310 128.640 ;
        RECT 25.500 128.440 26.310 128.580 ;
        RECT 25.500 128.395 25.790 128.440 ;
        RECT 25.990 128.380 26.310 128.440 ;
        RECT 41.260 128.240 41.400 128.735 ;
        RECT 42.550 128.720 42.870 128.780 ;
        RECT 43.945 128.735 44.235 128.780 ;
        RECT 50.370 128.720 50.690 128.780 ;
        RECT 51.305 128.735 51.595 128.780 ;
        RECT 52.640 128.735 52.990 128.780 ;
        RECT 52.670 128.720 52.990 128.735 ;
        RECT 58.650 128.720 58.970 128.980 ;
        RECT 59.570 128.720 59.890 128.980 ;
        RECT 61.870 128.920 62.190 128.980 ;
        RECT 67.850 128.920 68.170 128.980 ;
        RECT 69.245 128.920 69.535 128.965 ;
        RECT 61.870 128.780 69.535 128.920 ;
        RECT 61.870 128.720 62.190 128.780 ;
        RECT 67.850 128.720 68.170 128.780 ;
        RECT 69.245 128.735 69.535 128.780 ;
        RECT 70.580 128.920 70.870 128.965 ;
        RECT 75.670 128.920 75.990 128.980 ;
        RECT 81.280 128.965 81.420 129.120 ;
        RECT 81.650 129.060 81.970 129.120 ;
        RECT 70.580 128.780 75.990 128.920 ;
        RECT 70.580 128.735 70.870 128.780 ;
        RECT 75.670 128.720 75.990 128.780 ;
        RECT 81.205 128.735 81.495 128.965 ;
        RECT 82.585 128.735 82.875 128.965 ;
        RECT 45.280 128.580 45.570 128.625 ;
        RECT 45.770 128.580 46.090 128.640 ;
        RECT 44.020 128.440 46.090 128.580 ;
        RECT 44.020 128.240 44.160 128.440 ;
        RECT 45.280 128.395 45.570 128.440 ;
        RECT 45.770 128.380 46.090 128.440 ;
        RECT 50.830 128.580 51.150 128.640 ;
        RECT 59.125 128.580 59.415 128.625 ;
        RECT 50.830 128.440 59.415 128.580 ;
        RECT 50.830 128.380 51.150 128.440 ;
        RECT 59.125 128.395 59.415 128.440 ;
        RECT 62.330 128.580 62.650 128.640 ;
        RECT 63.110 128.580 63.400 128.625 ;
        RECT 62.330 128.440 63.400 128.580 ;
        RECT 62.330 128.380 62.650 128.440 ;
        RECT 63.110 128.395 63.400 128.440 ;
        RECT 80.730 128.580 81.050 128.640 ;
        RECT 82.125 128.580 82.415 128.625 ;
        RECT 82.660 128.580 82.800 128.735 ;
        RECT 83.030 128.720 83.350 128.980 ;
        RECT 83.580 128.965 83.720 129.120 ;
        RECT 84.500 129.120 88.410 129.260 ;
        RECT 84.500 128.965 84.640 129.120 ;
        RECT 88.090 129.060 88.410 129.120 ;
        RECT 99.105 129.260 99.395 129.305 ;
        RECT 100.295 129.260 100.585 129.305 ;
        RECT 102.815 129.260 103.105 129.305 ;
        RECT 129.490 129.260 129.810 129.320 ;
        RECT 99.105 129.120 103.105 129.260 ;
        RECT 99.105 129.075 99.395 129.120 ;
        RECT 100.295 129.075 100.585 129.120 ;
        RECT 102.815 129.075 103.105 129.120 ;
        RECT 105.660 129.120 129.810 129.260 ;
        RECT 83.505 128.735 83.795 128.965 ;
        RECT 84.425 128.735 84.715 128.965 ;
        RECT 85.345 128.920 85.635 128.965 ;
        RECT 90.850 128.920 91.170 128.980 ;
        RECT 85.345 128.780 91.170 128.920 ;
        RECT 85.345 128.735 85.635 128.780 ;
        RECT 90.850 128.720 91.170 128.780 ;
        RECT 91.310 128.920 91.630 128.980 ;
        RECT 98.225 128.920 98.515 128.965 ;
        RECT 100.970 128.920 101.290 128.980 ;
        RECT 105.660 128.920 105.800 129.120 ;
        RECT 129.490 129.060 129.810 129.120 ;
        RECT 132.225 129.260 132.515 129.305 ;
        RECT 133.415 129.260 133.705 129.305 ;
        RECT 135.935 129.260 136.225 129.305 ;
        RECT 132.225 129.120 136.225 129.260 ;
        RECT 132.225 129.075 132.515 129.120 ;
        RECT 133.415 129.075 133.705 129.120 ;
        RECT 135.935 129.075 136.225 129.120 ;
        RECT 144.225 129.260 144.515 129.305 ;
        RECT 145.130 129.260 145.450 129.320 ;
        RECT 144.225 129.120 145.450 129.260 ;
        RECT 144.225 129.075 144.515 129.120 ;
        RECT 145.130 129.060 145.450 129.120 ;
        RECT 148.350 129.060 148.670 129.320 ;
        RECT 149.245 129.260 149.535 129.305 ;
        RECT 150.435 129.260 150.725 129.305 ;
        RECT 152.955 129.260 153.245 129.305 ;
        RECT 149.245 129.120 153.245 129.260 ;
        RECT 149.245 129.075 149.535 129.120 ;
        RECT 150.435 129.075 150.725 129.120 ;
        RECT 152.955 129.075 153.245 129.120 ;
        RECT 91.310 128.780 98.515 128.920 ;
        RECT 91.310 128.720 91.630 128.780 ;
        RECT 98.225 128.735 98.515 128.780 ;
        RECT 99.220 128.780 105.800 128.920 ;
        RECT 106.045 128.920 106.335 128.965 ;
        RECT 109.265 128.920 109.555 128.965 ;
        RECT 106.045 128.780 109.555 128.920 ;
        RECT 87.630 128.580 87.950 128.640 ;
        RECT 91.400 128.580 91.540 128.720 ;
        RECT 80.730 128.440 82.800 128.580 ;
        RECT 83.120 128.440 84.640 128.580 ;
        RECT 80.730 128.380 81.050 128.440 ;
        RECT 82.125 128.395 82.415 128.440 ;
        RECT 41.260 128.100 44.160 128.240 ;
        RECT 58.205 128.240 58.495 128.285 ;
        RECT 58.650 128.240 58.970 128.300 ;
        RECT 58.205 128.100 58.970 128.240 ;
        RECT 58.205 128.055 58.495 128.100 ;
        RECT 58.650 128.040 58.970 128.100 ;
        RECT 67.850 128.240 68.170 128.300 ;
        RECT 68.785 128.240 69.075 128.285 ;
        RECT 67.850 128.100 69.075 128.240 ;
        RECT 67.850 128.040 68.170 128.100 ;
        RECT 68.785 128.055 69.075 128.100 ;
        RECT 78.430 128.240 78.750 128.300 ;
        RECT 79.825 128.240 80.115 128.285 ;
        RECT 78.430 128.100 80.115 128.240 ;
        RECT 78.430 128.040 78.750 128.100 ;
        RECT 79.825 128.055 80.115 128.100 ;
        RECT 80.285 128.240 80.575 128.285 ;
        RECT 83.120 128.240 83.260 128.440 ;
        RECT 84.500 128.300 84.640 128.440 ;
        RECT 87.630 128.440 91.540 128.580 ;
        RECT 94.070 128.580 94.390 128.640 ;
        RECT 95.465 128.580 95.755 128.625 ;
        RECT 95.910 128.580 96.230 128.640 ;
        RECT 94.070 128.440 96.230 128.580 ;
        RECT 87.630 128.380 87.950 128.440 ;
        RECT 94.070 128.380 94.390 128.440 ;
        RECT 95.465 128.395 95.755 128.440 ;
        RECT 95.910 128.380 96.230 128.440 ;
        RECT 96.385 128.580 96.675 128.625 ;
        RECT 99.220 128.580 99.360 128.780 ;
        RECT 100.970 128.720 101.290 128.780 ;
        RECT 106.045 128.735 106.335 128.780 ;
        RECT 109.265 128.735 109.555 128.780 ;
        RECT 109.710 128.920 110.030 128.980 ;
        RECT 110.185 128.920 110.475 128.965 ;
        RECT 109.710 128.780 110.475 128.920 ;
        RECT 96.385 128.440 99.360 128.580 ;
        RECT 99.560 128.580 99.850 128.625 ;
        RECT 104.190 128.580 104.510 128.640 ;
        RECT 99.560 128.440 104.510 128.580 ;
        RECT 96.385 128.395 96.675 128.440 ;
        RECT 99.560 128.395 99.850 128.440 ;
        RECT 104.190 128.380 104.510 128.440 ;
        RECT 80.285 128.100 83.260 128.240 ;
        RECT 80.285 128.055 80.575 128.100 ;
        RECT 84.410 128.040 84.730 128.300 ;
        RECT 105.125 128.240 105.415 128.285 ;
        RECT 106.120 128.240 106.260 128.735 ;
        RECT 109.340 128.580 109.480 128.735 ;
        RECT 109.710 128.720 110.030 128.780 ;
        RECT 110.185 128.735 110.475 128.780 ;
        RECT 111.105 128.920 111.395 128.965 ;
        RECT 111.565 128.920 111.855 128.965 ;
        RECT 111.105 128.780 111.855 128.920 ;
        RECT 111.105 128.735 111.395 128.780 ;
        RECT 111.565 128.735 111.855 128.780 ;
        RECT 130.410 128.920 130.730 128.980 ;
        RECT 131.345 128.920 131.635 128.965 ;
        RECT 134.090 128.920 134.410 128.980 ;
        RECT 145.605 128.920 145.895 128.965 ;
        RECT 130.410 128.780 134.410 128.920 ;
        RECT 130.410 128.720 130.730 128.780 ;
        RECT 131.345 128.735 131.635 128.780 ;
        RECT 134.090 128.720 134.410 128.780 ;
        RECT 144.300 128.780 145.895 128.920 ;
        RECT 125.350 128.580 125.670 128.640 ;
        RECT 132.710 128.625 133.030 128.640 ;
        RECT 132.680 128.580 133.030 128.625 ;
        RECT 109.340 128.440 125.670 128.580 ;
        RECT 132.515 128.440 133.030 128.580 ;
        RECT 125.350 128.380 125.670 128.440 ;
        RECT 132.680 128.395 133.030 128.440 ;
        RECT 132.710 128.380 133.030 128.395 ;
        RECT 136.390 128.580 136.710 128.640 ;
        RECT 141.005 128.580 141.295 128.625 ;
        RECT 144.300 128.580 144.440 128.780 ;
        RECT 145.605 128.735 145.895 128.780 ;
        RECT 136.390 128.440 144.440 128.580 ;
        RECT 136.390 128.380 136.710 128.440 ;
        RECT 141.005 128.395 141.295 128.440 ;
        RECT 144.670 128.380 144.990 128.640 ;
        RECT 149.700 128.580 149.990 128.625 ;
        RECT 152.030 128.580 152.350 128.640 ;
        RECT 149.700 128.440 152.350 128.580 ;
        RECT 149.700 128.395 149.990 128.440 ;
        RECT 152.030 128.380 152.350 128.440 ;
        RECT 105.125 128.100 106.260 128.240 ;
        RECT 107.410 128.240 107.730 128.300 ;
        RECT 108.805 128.240 109.095 128.285 ;
        RECT 107.410 128.100 109.095 128.240 ;
        RECT 105.125 128.055 105.415 128.100 ;
        RECT 107.410 128.040 107.730 128.100 ;
        RECT 108.805 128.055 109.095 128.100 ;
        RECT 109.710 128.240 110.030 128.300 ;
        RECT 112.485 128.240 112.775 128.285 ;
        RECT 109.710 128.100 112.775 128.240 ;
        RECT 109.710 128.040 110.030 128.100 ;
        RECT 112.485 128.055 112.775 128.100 ;
        RECT 136.850 128.240 137.170 128.300 ;
        RECT 144.760 128.240 144.900 128.380 ;
        RECT 136.850 128.100 144.900 128.240 ;
        RECT 146.525 128.240 146.815 128.285 ;
        RECT 154.330 128.240 154.650 128.300 ;
        RECT 146.525 128.100 154.650 128.240 ;
        RECT 136.850 128.040 137.170 128.100 ;
        RECT 146.525 128.055 146.815 128.100 ;
        RECT 154.330 128.040 154.650 128.100 ;
        RECT 22.700 127.420 157.820 127.900 ;
        RECT 30.130 127.220 30.450 127.280 ;
        RECT 36.570 127.220 36.890 127.280 ;
        RECT 67.390 127.220 67.710 127.280 ;
        RECT 28.380 127.080 30.450 127.220 ;
        RECT 28.380 126.940 28.520 127.080 ;
        RECT 30.130 127.020 30.450 127.080 ;
        RECT 33.440 127.080 36.890 127.220 ;
        RECT 28.290 126.680 28.610 126.940 ;
        RECT 33.440 126.925 33.580 127.080 ;
        RECT 36.570 127.020 36.890 127.080 ;
        RECT 38.500 127.080 67.710 127.220 ;
        RECT 38.500 126.925 38.640 127.080 ;
        RECT 67.390 127.020 67.710 127.080 ;
        RECT 104.190 127.020 104.510 127.280 ;
        RECT 132.265 127.035 132.555 127.265 ;
        RECT 137.785 127.035 138.075 127.265 ;
        RECT 138.690 127.220 139.010 127.280 ;
        RECT 138.690 127.080 139.380 127.220 ;
        RECT 29.225 126.880 29.515 126.925 ;
        RECT 33.365 126.880 33.655 126.925 ;
        RECT 29.225 126.740 33.655 126.880 ;
        RECT 29.225 126.695 29.515 126.740 ;
        RECT 33.365 126.695 33.655 126.740 ;
        RECT 34.445 126.880 34.735 126.925 ;
        RECT 34.445 126.740 35.880 126.880 ;
        RECT 34.445 126.695 34.735 126.740 ;
        RECT 35.740 126.600 35.880 126.740 ;
        RECT 38.425 126.695 38.715 126.925 ;
        RECT 45.310 126.680 45.630 126.940 ;
        RECT 50.845 126.880 51.135 126.925 ;
        RECT 52.225 126.880 52.515 126.925 ;
        RECT 48.620 126.740 52.515 126.880 ;
        RECT 29.685 126.355 29.975 126.585 ;
        RECT 27.830 125.520 28.150 125.580 ;
        RECT 28.305 125.520 28.595 125.565 ;
        RECT 27.830 125.380 28.595 125.520 ;
        RECT 29.760 125.520 29.900 126.355 ;
        RECT 35.650 126.340 35.970 126.600 ;
        RECT 36.570 126.340 36.890 126.600 ;
        RECT 43.930 126.340 44.250 126.600 ;
        RECT 44.405 126.540 44.695 126.585 ;
        RECT 47.150 126.540 47.470 126.600 ;
        RECT 44.405 126.400 47.470 126.540 ;
        RECT 44.405 126.355 44.695 126.400 ;
        RECT 47.150 126.340 47.470 126.400 ;
        RECT 42.550 126.000 42.870 126.260 ;
        RECT 44.020 126.200 44.160 126.340 ;
        RECT 48.620 126.200 48.760 126.740 ;
        RECT 50.845 126.695 51.135 126.740 ;
        RECT 52.225 126.695 52.515 126.740 ;
        RECT 59.570 126.880 59.890 126.940 ;
        RECT 61.885 126.880 62.175 126.925 ;
        RECT 59.570 126.740 62.175 126.880 ;
        RECT 59.570 126.680 59.890 126.740 ;
        RECT 61.885 126.695 62.175 126.740 ;
        RECT 76.590 126.680 76.910 126.940 ;
        RECT 97.750 126.880 98.070 126.940 ;
        RECT 106.965 126.880 107.255 126.925 ;
        RECT 97.750 126.740 107.255 126.880 ;
        RECT 97.750 126.680 98.070 126.740 ;
        RECT 106.965 126.695 107.255 126.740 ;
        RECT 107.410 126.680 107.730 126.940 ;
        RECT 130.410 126.880 130.730 126.940 ;
        RECT 109.800 126.740 114.080 126.880 ;
        RECT 109.800 126.600 109.940 126.740 ;
        RECT 54.525 126.540 54.815 126.585 ;
        RECT 58.190 126.540 58.510 126.600 ;
        RECT 54.525 126.400 58.510 126.540 ;
        RECT 54.525 126.355 54.815 126.400 ;
        RECT 58.190 126.340 58.510 126.400 ;
        RECT 58.650 126.340 58.970 126.600 ;
        RECT 60.950 126.540 61.270 126.600 ;
        RECT 64.185 126.540 64.475 126.585 ;
        RECT 60.950 126.400 64.475 126.540 ;
        RECT 60.950 126.340 61.270 126.400 ;
        RECT 64.185 126.355 64.475 126.400 ;
        RECT 44.020 126.060 48.760 126.200 ;
        RECT 54.065 126.200 54.355 126.245 ;
        RECT 57.270 126.200 57.590 126.260 ;
        RECT 54.065 126.060 57.590 126.200 ;
        RECT 54.065 126.015 54.355 126.060 ;
        RECT 57.270 126.000 57.590 126.060 ;
        RECT 63.710 126.000 64.030 126.260 ;
        RECT 64.260 126.200 64.400 126.355 ;
        RECT 67.850 126.340 68.170 126.600 ;
        RECT 76.130 126.540 76.450 126.600 ;
        RECT 77.065 126.540 77.355 126.585 ;
        RECT 76.130 126.400 77.355 126.540 ;
        RECT 76.130 126.340 76.450 126.400 ;
        RECT 77.065 126.355 77.355 126.400 ;
        RECT 78.430 126.340 78.750 126.600 ;
        RECT 78.905 126.540 79.195 126.585 ;
        RECT 79.350 126.540 79.670 126.600 ;
        RECT 80.270 126.585 80.590 126.600 ;
        RECT 92.690 126.585 93.010 126.600 ;
        RECT 78.905 126.400 79.670 126.540 ;
        RECT 78.905 126.355 79.195 126.400 ;
        RECT 79.350 126.340 79.670 126.400 ;
        RECT 80.240 126.355 80.590 126.585 ;
        RECT 92.660 126.355 93.010 126.585 ;
        RECT 80.270 126.340 80.590 126.355 ;
        RECT 92.690 126.340 93.010 126.355 ;
        RECT 105.110 126.340 105.430 126.600 ;
        RECT 105.585 126.540 105.875 126.585 ;
        RECT 109.710 126.540 110.030 126.600 ;
        RECT 105.585 126.400 110.030 126.540 ;
        RECT 105.585 126.355 105.875 126.400 ;
        RECT 109.710 126.340 110.030 126.400 ;
        RECT 110.630 126.540 110.950 126.600 ;
        RECT 113.450 126.540 113.740 126.585 ;
        RECT 110.630 126.400 113.740 126.540 ;
        RECT 113.940 126.540 114.080 126.740 ;
        RECT 115.320 126.740 130.730 126.880 ;
        RECT 132.340 126.880 132.480 127.035 ;
        RECT 135.010 126.880 135.330 126.940 ;
        RECT 132.340 126.740 136.160 126.880 ;
        RECT 115.320 126.585 115.460 126.740 ;
        RECT 130.410 126.680 130.730 126.740 ;
        RECT 135.010 126.680 135.330 126.740 ;
        RECT 114.785 126.540 115.075 126.585 ;
        RECT 115.245 126.540 115.535 126.585 ;
        RECT 116.525 126.540 116.815 126.585 ;
        RECT 113.940 126.400 114.540 126.540 ;
        RECT 110.630 126.340 110.950 126.400 ;
        RECT 113.450 126.355 113.740 126.400 ;
        RECT 79.785 126.200 80.075 126.245 ;
        RECT 80.975 126.200 81.265 126.245 ;
        RECT 83.495 126.200 83.785 126.245 ;
        RECT 89.025 126.200 89.315 126.245 ;
        RECT 64.260 126.060 67.160 126.200 ;
        RECT 49.005 125.860 49.295 125.905 ;
        RECT 54.970 125.860 55.290 125.920 ;
        RECT 55.445 125.860 55.735 125.905 ;
        RECT 34.360 125.720 35.880 125.860 ;
        RECT 31.050 125.520 31.370 125.580 ;
        RECT 34.360 125.565 34.500 125.720 ;
        RECT 34.285 125.520 34.575 125.565 ;
        RECT 29.760 125.380 34.575 125.520 ;
        RECT 27.830 125.320 28.150 125.380 ;
        RECT 28.305 125.335 28.595 125.380 ;
        RECT 31.050 125.320 31.370 125.380 ;
        RECT 34.285 125.335 34.575 125.380 ;
        RECT 34.730 125.520 35.050 125.580 ;
        RECT 35.740 125.565 35.880 125.720 ;
        RECT 49.005 125.720 54.280 125.860 ;
        RECT 49.005 125.675 49.295 125.720 ;
        RECT 35.205 125.520 35.495 125.565 ;
        RECT 34.730 125.380 35.495 125.520 ;
        RECT 34.730 125.320 35.050 125.380 ;
        RECT 35.205 125.335 35.495 125.380 ;
        RECT 35.665 125.335 35.955 125.565 ;
        RECT 37.505 125.520 37.795 125.565 ;
        RECT 49.450 125.520 49.770 125.580 ;
        RECT 37.505 125.380 49.770 125.520 ;
        RECT 37.505 125.335 37.795 125.380 ;
        RECT 49.450 125.320 49.770 125.380 ;
        RECT 50.830 125.320 51.150 125.580 ;
        RECT 51.290 125.520 51.610 125.580 ;
        RECT 54.140 125.565 54.280 125.720 ;
        RECT 54.970 125.720 55.735 125.860 ;
        RECT 54.970 125.660 55.290 125.720 ;
        RECT 55.445 125.675 55.735 125.720 ;
        RECT 66.010 125.660 66.330 125.920 ;
        RECT 67.020 125.905 67.160 126.060 ;
        RECT 79.785 126.060 83.785 126.200 ;
        RECT 79.785 126.015 80.075 126.060 ;
        RECT 80.975 126.015 81.265 126.060 ;
        RECT 83.495 126.015 83.785 126.060 ;
        RECT 85.880 126.060 89.315 126.200 ;
        RECT 66.945 125.675 67.235 125.905 ;
        RECT 79.390 125.860 79.680 125.905 ;
        RECT 81.490 125.860 81.780 125.905 ;
        RECT 83.060 125.860 83.350 125.905 ;
        RECT 79.390 125.720 83.350 125.860 ;
        RECT 79.390 125.675 79.680 125.720 ;
        RECT 81.490 125.675 81.780 125.720 ;
        RECT 83.060 125.675 83.350 125.720 ;
        RECT 85.880 125.580 86.020 126.060 ;
        RECT 89.025 126.015 89.315 126.060 ;
        RECT 91.310 126.000 91.630 126.260 ;
        RECT 92.205 126.200 92.495 126.245 ;
        RECT 93.395 126.200 93.685 126.245 ;
        RECT 95.915 126.200 96.205 126.245 ;
        RECT 92.205 126.060 96.205 126.200 ;
        RECT 92.205 126.015 92.495 126.060 ;
        RECT 93.395 126.015 93.685 126.060 ;
        RECT 95.915 126.015 96.205 126.060 ;
        RECT 101.430 126.200 101.750 126.260 ;
        RECT 103.285 126.200 103.575 126.245 ;
        RECT 101.430 126.060 103.575 126.200 ;
        RECT 101.430 126.000 101.750 126.060 ;
        RECT 103.285 126.015 103.575 126.060 ;
        RECT 110.195 126.200 110.485 126.245 ;
        RECT 112.715 126.200 113.005 126.245 ;
        RECT 113.905 126.200 114.195 126.245 ;
        RECT 110.195 126.060 114.195 126.200 ;
        RECT 114.400 126.200 114.540 126.400 ;
        RECT 114.785 126.400 115.535 126.540 ;
        RECT 114.785 126.355 115.075 126.400 ;
        RECT 115.245 126.355 115.535 126.400 ;
        RECT 115.780 126.400 116.815 126.540 ;
        RECT 115.780 126.200 115.920 126.400 ;
        RECT 116.525 126.355 116.815 126.400 ;
        RECT 123.065 126.540 123.355 126.585 ;
        RECT 125.350 126.540 125.670 126.600 ;
        RECT 123.065 126.400 125.670 126.540 ;
        RECT 123.065 126.355 123.355 126.400 ;
        RECT 125.350 126.340 125.670 126.400 ;
        RECT 126.270 126.340 126.590 126.600 ;
        RECT 131.345 126.540 131.635 126.585 ;
        RECT 130.270 126.400 131.635 126.540 ;
        RECT 114.400 126.060 115.920 126.200 ;
        RECT 116.125 126.200 116.415 126.245 ;
        RECT 117.315 126.200 117.605 126.245 ;
        RECT 119.835 126.200 120.125 126.245 ;
        RECT 116.125 126.060 120.125 126.200 ;
        RECT 110.195 126.015 110.485 126.060 ;
        RECT 112.715 126.015 113.005 126.060 ;
        RECT 113.905 126.015 114.195 126.060 ;
        RECT 116.125 126.015 116.415 126.060 ;
        RECT 117.315 126.015 117.605 126.060 ;
        RECT 119.835 126.015 120.125 126.060 ;
        RECT 91.810 125.860 92.100 125.905 ;
        RECT 93.910 125.860 94.200 125.905 ;
        RECT 95.480 125.860 95.770 125.905 ;
        RECT 91.810 125.720 95.770 125.860 ;
        RECT 91.810 125.675 92.100 125.720 ;
        RECT 93.910 125.675 94.200 125.720 ;
        RECT 95.480 125.675 95.770 125.720 ;
        RECT 98.225 125.860 98.515 125.905 ;
        RECT 101.520 125.860 101.660 126.000 ;
        RECT 98.225 125.720 101.660 125.860 ;
        RECT 110.630 125.860 110.920 125.905 ;
        RECT 112.200 125.860 112.490 125.905 ;
        RECT 114.300 125.860 114.590 125.905 ;
        RECT 110.630 125.720 114.590 125.860 ;
        RECT 98.225 125.675 98.515 125.720 ;
        RECT 110.630 125.675 110.920 125.720 ;
        RECT 112.200 125.675 112.490 125.720 ;
        RECT 114.300 125.675 114.590 125.720 ;
        RECT 115.730 125.860 116.020 125.905 ;
        RECT 117.830 125.860 118.120 125.905 ;
        RECT 119.400 125.860 119.690 125.905 ;
        RECT 115.730 125.720 119.690 125.860 ;
        RECT 126.360 125.860 126.500 126.340 ;
        RECT 128.570 126.200 128.890 126.260 ;
        RECT 130.270 126.200 130.410 126.400 ;
        RECT 131.345 126.355 131.635 126.400 ;
        RECT 133.170 126.540 133.490 126.600 ;
        RECT 136.020 126.585 136.160 126.740 ;
        RECT 134.565 126.540 134.855 126.585 ;
        RECT 133.170 126.400 134.855 126.540 ;
        RECT 133.170 126.340 133.490 126.400 ;
        RECT 134.565 126.355 134.855 126.400 ;
        RECT 135.485 126.355 135.775 126.585 ;
        RECT 135.945 126.355 136.235 126.585 ;
        RECT 128.570 126.060 130.410 126.200 ;
        RECT 135.560 126.200 135.700 126.355 ;
        RECT 136.390 126.340 136.710 126.600 ;
        RECT 137.860 126.540 138.000 127.035 ;
        RECT 138.690 127.020 139.010 127.080 ;
        RECT 139.240 126.880 139.380 127.080 ;
        RECT 145.130 127.020 145.450 127.280 ;
        RECT 146.525 126.880 146.815 126.925 ;
        RECT 139.240 126.740 146.815 126.880 ;
        RECT 146.525 126.695 146.815 126.740 ;
        RECT 148.350 126.880 148.670 126.940 ;
        RECT 150.205 126.880 150.495 126.925 ;
        RECT 148.350 126.740 150.495 126.880 ;
        RECT 148.350 126.680 148.670 126.740 ;
        RECT 150.205 126.695 150.495 126.740 ;
        RECT 139.525 126.540 139.815 126.585 ;
        RECT 137.860 126.400 139.815 126.540 ;
        RECT 139.525 126.355 139.815 126.400 ;
        RECT 152.950 126.540 153.270 126.600 ;
        RECT 153.425 126.540 153.715 126.585 ;
        RECT 152.950 126.400 153.715 126.540 ;
        RECT 152.950 126.340 153.270 126.400 ;
        RECT 153.425 126.355 153.715 126.400 ;
        RECT 153.885 126.355 154.175 126.585 ;
        RECT 137.310 126.200 137.630 126.260 ;
        RECT 135.560 126.060 137.630 126.200 ;
        RECT 128.570 126.000 128.890 126.060 ;
        RECT 137.310 126.000 137.630 126.060 ;
        RECT 138.245 126.015 138.535 126.245 ;
        RECT 139.125 126.200 139.415 126.245 ;
        RECT 140.315 126.200 140.605 126.245 ;
        RECT 142.835 126.200 143.125 126.245 ;
        RECT 139.125 126.060 143.125 126.200 ;
        RECT 139.125 126.015 139.415 126.060 ;
        RECT 140.315 126.015 140.605 126.060 ;
        RECT 142.835 126.015 143.125 126.060 ;
        RECT 144.670 126.200 144.990 126.260 ;
        RECT 153.960 126.200 154.100 126.355 ;
        RECT 154.330 126.340 154.650 126.600 ;
        RECT 154.790 126.540 155.110 126.600 ;
        RECT 155.265 126.540 155.555 126.585 ;
        RECT 154.790 126.400 155.555 126.540 ;
        RECT 154.790 126.340 155.110 126.400 ;
        RECT 155.265 126.355 155.555 126.400 ;
        RECT 144.670 126.060 154.100 126.200 ;
        RECT 129.950 125.860 130.270 125.920 ;
        RECT 137.770 125.860 138.090 125.920 ;
        RECT 126.360 125.720 138.090 125.860 ;
        RECT 115.730 125.675 116.020 125.720 ;
        RECT 117.830 125.675 118.120 125.720 ;
        RECT 119.400 125.675 119.690 125.720 ;
        RECT 129.950 125.660 130.270 125.720 ;
        RECT 137.770 125.660 138.090 125.720 ;
        RECT 51.765 125.520 52.055 125.565 ;
        RECT 51.290 125.380 52.055 125.520 ;
        RECT 51.290 125.320 51.610 125.380 ;
        RECT 51.765 125.335 52.055 125.380 ;
        RECT 54.065 125.520 54.355 125.565 ;
        RECT 54.510 125.520 54.830 125.580 ;
        RECT 54.065 125.380 54.830 125.520 ;
        RECT 54.065 125.335 54.355 125.380 ;
        RECT 54.510 125.320 54.830 125.380 ;
        RECT 85.790 125.320 86.110 125.580 ;
        RECT 86.250 125.320 86.570 125.580 ;
        RECT 87.170 125.520 87.490 125.580 ;
        RECT 94.990 125.520 95.310 125.580 ;
        RECT 87.170 125.380 95.310 125.520 ;
        RECT 87.170 125.320 87.490 125.380 ;
        RECT 94.990 125.320 95.310 125.380 ;
        RECT 100.510 125.320 100.830 125.580 ;
        RECT 107.885 125.520 108.175 125.565 ;
        RECT 113.390 125.520 113.710 125.580 ;
        RECT 107.885 125.380 113.710 125.520 ;
        RECT 107.885 125.335 108.175 125.380 ;
        RECT 113.390 125.320 113.710 125.380 ;
        RECT 122.145 125.520 122.435 125.565 ;
        RECT 123.510 125.520 123.830 125.580 ;
        RECT 122.145 125.380 123.830 125.520 ;
        RECT 122.145 125.335 122.435 125.380 ;
        RECT 123.510 125.320 123.830 125.380 ;
        RECT 125.365 125.520 125.655 125.565 ;
        RECT 136.850 125.520 137.170 125.580 ;
        RECT 125.365 125.380 137.170 125.520 ;
        RECT 138.320 125.520 138.460 126.015 ;
        RECT 144.670 126.000 144.990 126.060 ;
        RECT 138.730 125.860 139.020 125.905 ;
        RECT 140.830 125.860 141.120 125.905 ;
        RECT 142.400 125.860 142.690 125.905 ;
        RECT 148.350 125.860 148.670 125.920 ;
        RECT 138.730 125.720 142.690 125.860 ;
        RECT 138.730 125.675 139.020 125.720 ;
        RECT 140.830 125.675 141.120 125.720 ;
        RECT 142.400 125.675 142.690 125.720 ;
        RECT 142.920 125.720 148.670 125.860 ;
        RECT 142.920 125.520 143.060 125.720 ;
        RECT 148.350 125.660 148.670 125.720 ;
        RECT 138.320 125.380 143.060 125.520 ;
        RECT 148.810 125.520 149.130 125.580 ;
        RECT 152.045 125.520 152.335 125.565 ;
        RECT 148.810 125.380 152.335 125.520 ;
        RECT 125.365 125.335 125.655 125.380 ;
        RECT 136.850 125.320 137.170 125.380 ;
        RECT 148.810 125.320 149.130 125.380 ;
        RECT 152.045 125.335 152.335 125.380 ;
        RECT 22.700 124.700 157.020 125.180 ;
        RECT 31.050 124.500 31.370 124.560 ;
        RECT 35.650 124.500 35.970 124.560 ;
        RECT 36.125 124.500 36.415 124.545 ;
        RECT 31.050 124.360 33.810 124.500 ;
        RECT 31.050 124.300 31.370 124.360 ;
        RECT 24.650 124.160 24.940 124.205 ;
        RECT 26.750 124.160 27.040 124.205 ;
        RECT 28.320 124.160 28.610 124.205 ;
        RECT 24.650 124.020 28.610 124.160 ;
        RECT 24.650 123.975 24.940 124.020 ;
        RECT 26.750 123.975 27.040 124.020 ;
        RECT 28.320 123.975 28.610 124.020 ;
        RECT 25.045 123.820 25.335 123.865 ;
        RECT 26.235 123.820 26.525 123.865 ;
        RECT 28.755 123.820 29.045 123.865 ;
        RECT 25.045 123.680 29.045 123.820 ;
        RECT 25.045 123.635 25.335 123.680 ;
        RECT 26.235 123.635 26.525 123.680 ;
        RECT 28.755 123.635 29.045 123.680 ;
        RECT 24.165 123.480 24.455 123.525 ;
        RECT 26.910 123.480 27.230 123.540 ;
        RECT 24.165 123.340 27.230 123.480 ;
        RECT 33.670 123.480 33.810 124.360 ;
        RECT 35.650 124.360 36.415 124.500 ;
        RECT 35.650 124.300 35.970 124.360 ;
        RECT 36.125 124.315 36.415 124.360 ;
        RECT 74.290 124.500 74.610 124.560 ;
        RECT 80.270 124.500 80.590 124.560 ;
        RECT 80.745 124.500 81.035 124.545 ;
        RECT 74.290 124.360 76.820 124.500 ;
        RECT 74.290 124.300 74.610 124.360 ;
        RECT 38.870 124.160 39.160 124.205 ;
        RECT 40.440 124.160 40.730 124.205 ;
        RECT 42.540 124.160 42.830 124.205 ;
        RECT 38.870 124.020 42.830 124.160 ;
        RECT 38.870 123.975 39.160 124.020 ;
        RECT 40.440 123.975 40.730 124.020 ;
        RECT 42.540 123.975 42.830 124.020 ;
        RECT 62.330 124.160 62.650 124.220 ;
        RECT 62.805 124.160 63.095 124.205 ;
        RECT 70.150 124.160 70.470 124.220 ;
        RECT 62.330 124.020 70.470 124.160 ;
        RECT 62.330 123.960 62.650 124.020 ;
        RECT 62.805 123.975 63.095 124.020 ;
        RECT 70.150 123.960 70.470 124.020 ;
        RECT 71.070 124.160 71.360 124.205 ;
        RECT 72.640 124.160 72.930 124.205 ;
        RECT 74.740 124.160 75.030 124.205 ;
        RECT 71.070 124.020 75.030 124.160 ;
        RECT 71.070 123.975 71.360 124.020 ;
        RECT 72.640 123.975 72.930 124.020 ;
        RECT 74.740 123.975 75.030 124.020 ;
        RECT 38.435 123.820 38.725 123.865 ;
        RECT 40.955 123.820 41.245 123.865 ;
        RECT 42.145 123.820 42.435 123.865 ;
        RECT 38.435 123.680 42.435 123.820 ;
        RECT 38.435 123.635 38.725 123.680 ;
        RECT 40.955 123.635 41.245 123.680 ;
        RECT 42.145 123.635 42.435 123.680 ;
        RECT 70.635 123.820 70.925 123.865 ;
        RECT 73.155 123.820 73.445 123.865 ;
        RECT 74.345 123.820 74.635 123.865 ;
        RECT 75.685 123.820 75.975 123.865 ;
        RECT 70.635 123.680 74.635 123.820 ;
        RECT 70.635 123.635 70.925 123.680 ;
        RECT 73.155 123.635 73.445 123.680 ;
        RECT 74.345 123.635 74.635 123.680 ;
        RECT 74.840 123.680 75.975 123.820 ;
        RECT 74.840 123.540 74.980 123.680 ;
        RECT 75.685 123.635 75.975 123.680 ;
        RECT 34.745 123.480 35.035 123.525 ;
        RECT 37.030 123.480 37.350 123.540 ;
        RECT 33.670 123.340 37.350 123.480 ;
        RECT 24.165 123.295 24.455 123.340 ;
        RECT 26.910 123.280 27.230 123.340 ;
        RECT 34.745 123.295 35.035 123.340 ;
        RECT 37.030 123.280 37.350 123.340 ;
        RECT 42.550 123.480 42.870 123.540 ;
        RECT 43.025 123.480 43.315 123.525 ;
        RECT 42.550 123.340 43.315 123.480 ;
        RECT 42.550 123.280 42.870 123.340 ;
        RECT 43.025 123.295 43.315 123.340 ;
        RECT 45.325 123.480 45.615 123.525 ;
        RECT 45.770 123.480 46.090 123.540 ;
        RECT 45.325 123.340 46.090 123.480 ;
        RECT 45.325 123.295 45.615 123.340 ;
        RECT 45.770 123.280 46.090 123.340 ;
        RECT 46.245 123.480 46.535 123.525 ;
        RECT 47.150 123.480 47.470 123.540 ;
        RECT 46.245 123.340 47.470 123.480 ;
        RECT 46.245 123.295 46.535 123.340 ;
        RECT 47.150 123.280 47.470 123.340 ;
        RECT 52.670 123.280 52.990 123.540 ;
        RECT 53.130 123.280 53.450 123.540 ;
        RECT 53.605 123.480 53.895 123.525 ;
        RECT 54.050 123.480 54.370 123.540 ;
        RECT 53.605 123.340 54.370 123.480 ;
        RECT 53.605 123.295 53.895 123.340 ;
        RECT 54.050 123.280 54.370 123.340 ;
        RECT 60.490 123.480 60.810 123.540 ;
        RECT 60.965 123.480 61.255 123.525 ;
        RECT 61.885 123.480 62.175 123.525 ;
        RECT 63.725 123.480 64.015 123.525 ;
        RECT 60.490 123.340 64.015 123.480 ;
        RECT 60.490 123.280 60.810 123.340 ;
        RECT 60.965 123.295 61.255 123.340 ;
        RECT 61.885 123.295 62.175 123.340 ;
        RECT 63.725 123.295 64.015 123.340 ;
        RECT 74.750 123.280 75.070 123.540 ;
        RECT 76.680 123.525 76.820 124.360 ;
        RECT 80.270 124.360 81.035 124.500 ;
        RECT 80.270 124.300 80.590 124.360 ;
        RECT 80.745 124.315 81.035 124.360 ;
        RECT 84.425 124.500 84.715 124.545 ;
        RECT 86.250 124.500 86.570 124.560 ;
        RECT 84.425 124.360 86.570 124.500 ;
        RECT 84.425 124.315 84.715 124.360 ;
        RECT 86.250 124.300 86.570 124.360 ;
        RECT 92.230 124.300 92.550 124.560 ;
        RECT 92.690 124.500 93.010 124.560 ;
        RECT 93.625 124.500 93.915 124.545 ;
        RECT 92.690 124.360 93.915 124.500 ;
        RECT 92.690 124.300 93.010 124.360 ;
        RECT 93.625 124.315 93.915 124.360 ;
        RECT 94.990 124.500 95.310 124.560 ;
        RECT 97.305 124.500 97.595 124.545 ;
        RECT 100.510 124.500 100.830 124.560 ;
        RECT 94.990 124.360 97.060 124.500 ;
        RECT 94.990 124.300 95.310 124.360 ;
        RECT 83.505 124.160 83.795 124.205 ;
        RECT 81.970 124.020 83.795 124.160 ;
        RECT 81.970 123.820 82.110 124.020 ;
        RECT 83.505 123.975 83.795 124.020 ;
        RECT 86.725 124.160 87.015 124.205 ;
        RECT 92.320 124.160 92.460 124.300 ;
        RECT 95.450 124.160 95.770 124.220 ;
        RECT 86.725 124.020 95.770 124.160 ;
        RECT 86.725 123.975 87.015 124.020 ;
        RECT 95.450 123.960 95.770 124.020 ;
        RECT 96.385 123.975 96.675 124.205 ;
        RECT 96.920 124.160 97.060 124.360 ;
        RECT 97.305 124.360 100.830 124.500 ;
        RECT 97.305 124.315 97.595 124.360 ;
        RECT 100.510 124.300 100.830 124.360 ;
        RECT 110.185 124.500 110.475 124.545 ;
        RECT 110.630 124.500 110.950 124.560 ;
        RECT 110.185 124.360 110.950 124.500 ;
        RECT 110.185 124.315 110.475 124.360 ;
        RECT 110.630 124.300 110.950 124.360 ;
        RECT 116.625 124.500 116.915 124.545 ;
        RECT 118.005 124.500 118.295 124.545 ;
        RECT 116.625 124.360 118.295 124.500 ;
        RECT 116.625 124.315 116.915 124.360 ;
        RECT 118.005 124.315 118.295 124.360 ;
        RECT 120.305 124.315 120.595 124.545 ;
        RECT 123.525 124.500 123.815 124.545 ;
        RECT 126.730 124.500 127.050 124.560 ;
        RECT 123.525 124.360 127.050 124.500 ;
        RECT 123.525 124.315 123.815 124.360 ;
        RECT 112.930 124.160 113.250 124.220 ;
        RECT 96.920 124.020 113.250 124.160 ;
        RECT 90.850 123.820 91.170 123.880 ;
        RECT 81.740 123.680 82.110 123.820 ;
        RECT 84.500 123.680 86.940 123.820 ;
        RECT 81.740 123.525 81.880 123.680 ;
        RECT 75.225 123.295 75.515 123.525 ;
        RECT 76.605 123.295 76.895 123.525 ;
        RECT 81.665 123.295 81.955 123.525 ;
        RECT 25.500 123.140 25.790 123.185 ;
        RECT 26.450 123.140 26.770 123.200 ;
        RECT 25.500 123.000 26.770 123.140 ;
        RECT 25.500 122.955 25.790 123.000 ;
        RECT 26.450 122.940 26.770 123.000 ;
        RECT 40.710 123.140 41.030 123.200 ;
        RECT 41.690 123.140 41.980 123.185 ;
        RECT 40.710 123.000 41.980 123.140 ;
        RECT 40.710 122.940 41.030 123.000 ;
        RECT 41.690 122.955 41.980 123.000 ;
        RECT 43.470 123.140 43.790 123.200 ;
        RECT 53.220 123.140 53.360 123.280 ;
        RECT 43.470 123.000 53.360 123.140 ;
        RECT 71.530 123.140 71.850 123.200 ;
        RECT 73.890 123.140 74.180 123.185 ;
        RECT 71.530 123.000 74.180 123.140 ;
        RECT 43.470 122.940 43.790 123.000 ;
        RECT 71.530 122.940 71.850 123.000 ;
        RECT 73.890 122.955 74.180 123.000 ;
        RECT 28.750 122.800 29.070 122.860 ;
        RECT 31.525 122.800 31.815 122.845 ;
        RECT 28.750 122.660 31.815 122.800 ;
        RECT 28.750 122.600 29.070 122.660 ;
        RECT 31.525 122.615 31.815 122.660 ;
        RECT 39.330 122.800 39.650 122.860 ;
        RECT 43.010 122.800 43.330 122.860 ;
        RECT 44.405 122.800 44.695 122.845 ;
        RECT 39.330 122.660 44.695 122.800 ;
        RECT 39.330 122.600 39.650 122.660 ;
        RECT 43.010 122.600 43.330 122.660 ;
        RECT 44.405 122.615 44.695 122.660 ;
        RECT 53.145 122.800 53.435 122.845 ;
        RECT 53.590 122.800 53.910 122.860 ;
        RECT 53.145 122.660 53.910 122.800 ;
        RECT 53.145 122.615 53.435 122.660 ;
        RECT 53.590 122.600 53.910 122.660 ;
        RECT 59.570 122.800 59.890 122.860 ;
        RECT 60.045 122.800 60.335 122.845 ;
        RECT 59.570 122.660 60.335 122.800 ;
        RECT 59.570 122.600 59.890 122.660 ;
        RECT 60.045 122.615 60.335 122.660 ;
        RECT 64.630 122.600 64.950 122.860 ;
        RECT 68.325 122.800 68.615 122.845 ;
        RECT 69.690 122.800 70.010 122.860 ;
        RECT 68.325 122.660 70.010 122.800 ;
        RECT 75.300 122.800 75.440 123.295 ;
        RECT 83.030 123.280 83.350 123.540 ;
        RECT 77.510 123.140 77.830 123.200 ;
        RECT 80.730 123.140 81.050 123.200 ;
        RECT 84.500 123.140 84.640 123.680 ;
        RECT 86.800 123.540 86.940 123.680 ;
        RECT 87.260 123.680 91.170 123.820 ;
        RECT 85.805 123.480 86.095 123.525 ;
        RECT 85.805 123.340 86.480 123.480 ;
        RECT 85.805 123.295 86.095 123.340 ;
        RECT 77.510 123.000 84.640 123.140 ;
        RECT 84.870 123.140 85.190 123.200 ;
        RECT 85.345 123.140 85.635 123.185 ;
        RECT 84.870 123.000 85.635 123.140 ;
        RECT 86.340 123.140 86.480 123.340 ;
        RECT 86.710 123.280 87.030 123.540 ;
        RECT 87.260 123.140 87.400 123.680 ;
        RECT 90.850 123.620 91.170 123.680 ;
        RECT 91.310 123.820 91.630 123.880 ;
        RECT 92.705 123.820 92.995 123.865 ;
        RECT 93.150 123.820 93.470 123.880 ;
        RECT 96.460 123.820 96.600 123.975 ;
        RECT 91.310 123.680 93.470 123.820 ;
        RECT 91.310 123.620 91.630 123.680 ;
        RECT 92.705 123.635 92.995 123.680 ;
        RECT 93.150 123.620 93.470 123.680 ;
        RECT 94.620 123.680 96.600 123.820 ;
        RECT 88.550 123.280 88.870 123.540 ;
        RECT 94.620 123.525 94.760 123.680 ;
        RECT 94.545 123.295 94.835 123.525 ;
        RECT 95.450 123.480 95.770 123.540 ;
        RECT 95.925 123.480 96.215 123.525 ;
        RECT 95.450 123.340 96.215 123.480 ;
        RECT 95.450 123.280 95.770 123.340 ;
        RECT 95.925 123.295 96.215 123.340 ;
        RECT 103.730 123.280 104.050 123.540 ;
        RECT 106.580 123.525 106.720 124.020 ;
        RECT 112.930 123.960 113.250 124.020 ;
        RECT 117.085 123.975 117.375 124.205 ;
        RECT 117.530 124.160 117.850 124.220 ;
        RECT 120.380 124.160 120.520 124.315 ;
        RECT 126.730 124.300 127.050 124.360 ;
        RECT 128.570 124.300 128.890 124.560 ;
        RECT 130.410 124.500 130.730 124.560 ;
        RECT 129.120 124.360 130.730 124.500 ;
        RECT 117.530 124.020 120.520 124.160 ;
        RECT 122.605 124.160 122.895 124.205 ;
        RECT 124.890 124.160 125.210 124.220 ;
        RECT 122.605 124.020 125.210 124.160 ;
        RECT 117.160 123.820 117.300 123.975 ;
        RECT 117.530 123.960 117.850 124.020 ;
        RECT 122.605 123.975 122.895 124.020 ;
        RECT 124.890 123.960 125.210 124.020 ;
        RECT 125.350 124.160 125.670 124.220 ;
        RECT 127.665 124.160 127.955 124.205 ;
        RECT 125.350 124.020 127.955 124.160 ;
        RECT 125.350 123.960 125.670 124.020 ;
        RECT 127.665 123.975 127.955 124.020 ;
        RECT 123.510 123.820 123.830 123.880 ;
        RECT 129.120 123.865 129.260 124.360 ;
        RECT 130.410 124.300 130.730 124.360 ;
        RECT 143.765 124.315 144.055 124.545 ;
        RECT 129.530 124.160 129.820 124.205 ;
        RECT 131.630 124.160 131.920 124.205 ;
        RECT 133.200 124.160 133.490 124.205 ;
        RECT 129.530 124.020 133.490 124.160 ;
        RECT 129.530 123.975 129.820 124.020 ;
        RECT 131.630 123.975 131.920 124.020 ;
        RECT 133.200 123.975 133.490 124.020 ;
        RECT 135.930 124.160 136.250 124.220 ;
        RECT 143.840 124.160 143.980 124.315 ;
        RECT 135.930 124.020 143.980 124.160 ;
        RECT 147.930 124.160 148.220 124.205 ;
        RECT 150.030 124.160 150.320 124.205 ;
        RECT 151.600 124.160 151.890 124.205 ;
        RECT 147.930 124.020 151.890 124.160 ;
        RECT 135.930 123.960 136.250 124.020 ;
        RECT 142.000 123.865 142.140 124.020 ;
        RECT 147.930 123.975 148.220 124.020 ;
        RECT 150.030 123.975 150.320 124.020 ;
        RECT 151.600 123.975 151.890 124.020 ;
        RECT 126.285 123.820 126.575 123.865 ;
        RECT 111.180 123.680 117.300 123.820 ;
        RECT 119.920 123.680 123.280 123.820 ;
        RECT 105.585 123.480 105.875 123.525 ;
        RECT 105.585 123.340 106.260 123.480 ;
        RECT 105.585 123.295 105.875 123.340 ;
        RECT 86.340 123.000 87.400 123.140 ;
        RECT 92.690 123.140 93.010 123.200 ;
        RECT 98.225 123.140 98.515 123.185 ;
        RECT 92.690 123.000 98.515 123.140 ;
        RECT 106.120 123.140 106.260 123.340 ;
        RECT 106.505 123.295 106.795 123.525 ;
        RECT 106.965 123.480 107.255 123.525 ;
        RECT 107.870 123.480 108.190 123.540 ;
        RECT 111.180 123.525 111.320 123.680 ;
        RECT 106.965 123.340 110.860 123.480 ;
        RECT 106.965 123.295 107.255 123.340 ;
        RECT 107.870 123.280 108.190 123.340 ;
        RECT 110.170 123.140 110.490 123.200 ;
        RECT 106.120 123.000 110.490 123.140 ;
        RECT 110.720 123.140 110.860 123.340 ;
        RECT 111.105 123.295 111.395 123.525 ;
        RECT 112.470 123.480 112.790 123.540 ;
        RECT 111.640 123.340 112.790 123.480 ;
        RECT 111.640 123.140 111.780 123.340 ;
        RECT 112.470 123.280 112.790 123.340 ;
        RECT 113.390 123.280 113.710 123.540 ;
        RECT 114.770 123.480 115.090 123.540 ;
        RECT 119.920 123.525 120.060 123.680 ;
        RECT 113.940 123.340 115.090 123.480 ;
        RECT 110.720 123.000 111.780 123.140 ;
        RECT 112.025 123.140 112.315 123.185 ;
        RECT 113.940 123.140 114.080 123.340 ;
        RECT 114.770 123.280 115.090 123.340 ;
        RECT 119.845 123.295 120.135 123.525 ;
        RECT 121.670 123.280 121.990 123.540 ;
        RECT 123.140 123.480 123.280 123.680 ;
        RECT 123.510 123.680 126.575 123.820 ;
        RECT 123.510 123.620 123.830 123.680 ;
        RECT 126.285 123.635 126.575 123.680 ;
        RECT 129.045 123.635 129.335 123.865 ;
        RECT 129.925 123.820 130.215 123.865 ;
        RECT 131.115 123.820 131.405 123.865 ;
        RECT 133.635 123.820 133.925 123.865 ;
        RECT 129.925 123.680 133.925 123.820 ;
        RECT 129.925 123.635 130.215 123.680 ;
        RECT 131.115 123.635 131.405 123.680 ;
        RECT 133.635 123.635 133.925 123.680 ;
        RECT 141.925 123.635 142.215 123.865 ;
        RECT 148.325 123.820 148.615 123.865 ;
        RECT 149.515 123.820 149.805 123.865 ;
        RECT 152.035 123.820 152.325 123.865 ;
        RECT 148.325 123.680 152.325 123.820 ;
        RECT 148.325 123.635 148.615 123.680 ;
        RECT 149.515 123.635 149.805 123.680 ;
        RECT 152.035 123.635 152.325 123.680 ;
        RECT 124.445 123.480 124.735 123.525 ;
        RECT 129.490 123.480 129.810 123.540 ;
        RECT 123.140 123.340 124.200 123.480 ;
        RECT 112.025 123.000 114.080 123.140 ;
        RECT 115.230 123.140 115.550 123.200 ;
        RECT 118.925 123.140 119.215 123.185 ;
        RECT 115.230 123.000 119.215 123.140 ;
        RECT 124.060 123.140 124.200 123.340 ;
        RECT 124.445 123.340 129.810 123.480 ;
        RECT 124.445 123.295 124.735 123.340 ;
        RECT 129.490 123.280 129.810 123.340 ;
        RECT 136.850 123.280 137.170 123.540 ;
        RECT 137.325 123.480 137.615 123.525 ;
        RECT 138.690 123.480 139.010 123.540 ;
        RECT 143.765 123.480 144.055 123.525 ;
        RECT 137.325 123.340 144.055 123.480 ;
        RECT 137.325 123.295 137.615 123.340 ;
        RECT 138.690 123.280 139.010 123.340 ;
        RECT 143.765 123.295 144.055 123.340 ;
        RECT 144.210 123.280 144.530 123.540 ;
        RECT 145.130 123.280 145.450 123.540 ;
        RECT 147.445 123.480 147.735 123.525 ;
        RECT 147.890 123.480 148.210 123.540 ;
        RECT 148.810 123.525 149.130 123.540 ;
        RECT 148.780 123.480 149.130 123.525 ;
        RECT 147.445 123.340 148.210 123.480 ;
        RECT 148.615 123.340 149.130 123.480 ;
        RECT 147.445 123.295 147.735 123.340 ;
        RECT 147.890 123.280 148.210 123.340 ;
        RECT 148.780 123.295 149.130 123.340 ;
        RECT 148.810 123.280 149.130 123.295 ;
        RECT 126.270 123.140 126.590 123.200 ;
        RECT 124.060 123.000 126.590 123.140 ;
        RECT 77.510 122.940 77.830 123.000 ;
        RECT 80.730 122.940 81.050 123.000 ;
        RECT 84.870 122.940 85.190 123.000 ;
        RECT 85.345 122.955 85.635 123.000 ;
        RECT 92.690 122.940 93.010 123.000 ;
        RECT 98.225 122.955 98.515 123.000 ;
        RECT 110.170 122.940 110.490 123.000 ;
        RECT 112.025 122.955 112.315 123.000 ;
        RECT 115.230 122.940 115.550 123.000 ;
        RECT 118.925 122.955 119.215 123.000 ;
        RECT 126.270 122.940 126.590 123.000 ;
        RECT 130.380 123.140 130.670 123.185 ;
        RECT 130.870 123.140 131.190 123.200 ;
        RECT 130.380 123.000 131.190 123.140 ;
        RECT 136.940 123.140 137.080 123.280 ;
        RECT 138.245 123.140 138.535 123.185 ;
        RECT 141.910 123.140 142.230 123.200 ;
        RECT 136.940 123.000 142.230 123.140 ;
        RECT 130.380 122.955 130.670 123.000 ;
        RECT 130.870 122.940 131.190 123.000 ;
        RECT 138.245 122.955 138.535 123.000 ;
        RECT 141.910 122.940 142.230 123.000 ;
        RECT 79.350 122.800 79.670 122.860 ;
        RECT 75.300 122.660 79.670 122.800 ;
        RECT 68.325 122.615 68.615 122.660 ;
        RECT 69.690 122.600 70.010 122.660 ;
        RECT 79.350 122.600 79.670 122.660 ;
        RECT 82.110 122.800 82.430 122.860 ;
        RECT 84.410 122.845 84.730 122.860 ;
        RECT 82.585 122.800 82.875 122.845 ;
        RECT 82.110 122.660 82.875 122.800 ;
        RECT 82.110 122.600 82.430 122.660 ;
        RECT 82.585 122.615 82.875 122.660 ;
        RECT 84.345 122.615 84.730 122.845 ;
        RECT 84.410 122.600 84.730 122.615 ;
        RECT 94.990 122.800 95.310 122.860 ;
        RECT 95.465 122.800 95.755 122.845 ;
        RECT 94.990 122.660 95.755 122.800 ;
        RECT 94.990 122.600 95.310 122.660 ;
        RECT 95.465 122.615 95.755 122.660 ;
        RECT 95.910 122.800 96.230 122.860 ;
        RECT 97.175 122.800 97.465 122.845 ;
        RECT 95.910 122.660 97.465 122.800 ;
        RECT 95.910 122.600 96.230 122.660 ;
        RECT 97.175 122.615 97.465 122.660 ;
        RECT 100.970 122.600 101.290 122.860 ;
        RECT 104.650 122.600 104.970 122.860 ;
        RECT 114.310 122.800 114.630 122.860 ;
        RECT 117.875 122.800 118.165 122.845 ;
        RECT 114.310 122.660 118.165 122.800 ;
        RECT 114.310 122.600 114.630 122.660 ;
        RECT 117.875 122.615 118.165 122.660 ;
        RECT 136.390 122.600 136.710 122.860 ;
        RECT 137.770 122.800 138.090 122.860 ;
        RECT 139.165 122.800 139.455 122.845 ;
        RECT 137.770 122.660 139.455 122.800 ;
        RECT 137.770 122.600 138.090 122.660 ;
        RECT 139.165 122.615 139.455 122.660 ;
        RECT 142.830 122.600 143.150 122.860 ;
        RECT 154.330 122.600 154.650 122.860 ;
        RECT 22.700 121.980 157.820 122.460 ;
        RECT 26.450 121.580 26.770 121.840 ;
        RECT 36.570 121.580 36.890 121.840 ;
        RECT 38.425 121.780 38.715 121.825 ;
        RECT 40.710 121.780 41.030 121.840 ;
        RECT 38.425 121.640 41.030 121.780 ;
        RECT 38.425 121.595 38.715 121.640 ;
        RECT 40.710 121.580 41.030 121.640 ;
        RECT 50.385 121.780 50.675 121.825 ;
        RECT 52.670 121.780 52.990 121.840 ;
        RECT 50.385 121.640 52.990 121.780 ;
        RECT 50.385 121.595 50.675 121.640 ;
        RECT 52.670 121.580 52.990 121.640 ;
        RECT 59.125 121.595 59.415 121.825 ;
        RECT 82.110 121.780 82.430 121.840 ;
        RECT 87.170 121.780 87.490 121.840 ;
        RECT 91.770 121.825 92.090 121.840 ;
        RECT 81.970 121.640 87.490 121.780 ;
        RECT 33.365 121.440 33.655 121.485 ;
        RECT 34.745 121.440 35.035 121.485 ;
        RECT 33.365 121.300 35.035 121.440 ;
        RECT 33.365 121.255 33.655 121.300 ;
        RECT 34.745 121.255 35.035 121.300 ;
        RECT 39.805 121.440 40.095 121.485 ;
        RECT 41.950 121.440 42.240 121.485 ;
        RECT 54.510 121.440 54.830 121.500 ;
        RECT 59.200 121.440 59.340 121.595 ;
        RECT 81.970 121.580 82.430 121.640 ;
        RECT 87.170 121.580 87.490 121.640 ;
        RECT 90.405 121.780 90.695 121.825 ;
        RECT 91.705 121.780 92.090 121.825 ;
        RECT 95.450 121.780 95.770 121.840 ;
        RECT 90.405 121.640 95.770 121.780 ;
        RECT 90.405 121.595 90.695 121.640 ;
        RECT 91.705 121.595 92.090 121.640 ;
        RECT 91.770 121.580 92.090 121.595 ;
        RECT 95.450 121.580 95.770 121.640 ;
        RECT 110.170 121.780 110.490 121.840 ;
        RECT 114.310 121.825 114.630 121.840 ;
        RECT 113.405 121.780 113.695 121.825 ;
        RECT 110.170 121.640 113.695 121.780 ;
        RECT 110.170 121.580 110.490 121.640 ;
        RECT 113.405 121.595 113.695 121.640 ;
        RECT 114.245 121.595 114.630 121.825 ;
        RECT 123.985 121.595 124.275 121.825 ;
        RECT 114.310 121.580 114.630 121.595 ;
        RECT 61.870 121.440 62.190 121.500 ;
        RECT 39.805 121.300 42.240 121.440 ;
        RECT 39.805 121.255 40.095 121.300 ;
        RECT 41.950 121.255 42.240 121.300 ;
        RECT 51.840 121.300 59.340 121.440 ;
        RECT 59.660 121.300 62.190 121.440 ;
        RECT 51.840 121.160 51.980 121.300 ;
        RECT 54.510 121.240 54.830 121.300 ;
        RECT 35.650 120.900 35.970 121.160 ;
        RECT 37.030 120.900 37.350 121.160 ;
        RECT 37.505 120.915 37.795 121.145 ;
        RECT 29.210 120.560 29.530 120.820 ;
        RECT 37.580 120.760 37.720 120.915 ;
        RECT 39.330 120.900 39.650 121.160 ;
        RECT 40.265 121.100 40.555 121.145 ;
        RECT 50.830 121.100 51.150 121.160 ;
        RECT 40.265 120.960 51.150 121.100 ;
        RECT 40.265 120.915 40.555 120.960 ;
        RECT 50.830 120.900 51.150 120.960 ;
        RECT 51.290 120.900 51.610 121.160 ;
        RECT 51.750 120.900 52.070 121.160 ;
        RECT 53.590 121.145 53.910 121.160 ;
        RECT 59.660 121.145 59.800 121.300 ;
        RECT 61.870 121.240 62.190 121.300 ;
        RECT 68.785 121.440 69.075 121.485 ;
        RECT 81.970 121.440 82.110 121.580 ;
        RECT 68.785 121.300 82.110 121.440 ;
        RECT 86.710 121.440 87.030 121.500 ;
        RECT 88.565 121.440 88.855 121.485 ;
        RECT 86.710 121.300 88.855 121.440 ;
        RECT 68.785 121.255 69.075 121.300 ;
        RECT 86.710 121.240 87.030 121.300 ;
        RECT 88.565 121.255 88.855 121.300 ;
        RECT 89.485 121.440 89.775 121.485 ;
        RECT 90.850 121.440 91.170 121.500 ;
        RECT 89.485 121.300 91.170 121.440 ;
        RECT 89.485 121.255 89.775 121.300 ;
        RECT 90.850 121.240 91.170 121.300 ;
        RECT 92.690 121.240 93.010 121.500 ;
        RECT 99.145 121.440 99.435 121.485 ;
        RECT 100.970 121.440 101.290 121.500 ;
        RECT 99.145 121.300 101.290 121.440 ;
        RECT 99.145 121.255 99.435 121.300 ;
        RECT 100.970 121.240 101.290 121.300 ;
        RECT 103.240 121.440 103.530 121.485 ;
        RECT 104.650 121.440 104.970 121.500 ;
        RECT 103.240 121.300 104.970 121.440 ;
        RECT 103.240 121.255 103.530 121.300 ;
        RECT 104.650 121.240 104.970 121.300 ;
        RECT 115.230 121.240 115.550 121.500 ;
        RECT 122.300 121.440 122.590 121.485 ;
        RECT 124.060 121.440 124.200 121.595 ;
        RECT 126.270 121.580 126.590 121.840 ;
        RECT 129.965 121.780 130.255 121.825 ;
        RECT 130.870 121.780 131.190 121.840 ;
        RECT 146.970 121.780 147.290 121.840 ;
        RECT 129.965 121.640 131.190 121.780 ;
        RECT 129.965 121.595 130.255 121.640 ;
        RECT 130.870 121.580 131.190 121.640 ;
        RECT 134.640 121.640 147.290 121.780 ;
        RECT 128.585 121.440 128.875 121.485 ;
        RECT 133.630 121.440 133.950 121.500 ;
        RECT 122.300 121.300 124.200 121.440 ;
        RECT 124.520 121.300 126.500 121.440 ;
        RECT 122.300 121.255 122.590 121.300 ;
        RECT 53.560 121.100 53.910 121.145 ;
        RECT 53.395 120.960 53.910 121.100 ;
        RECT 53.560 120.915 53.910 120.960 ;
        RECT 59.585 120.915 59.875 121.145 ;
        RECT 60.920 121.100 61.210 121.145 ;
        RECT 66.945 121.100 67.235 121.145 ;
        RECT 60.920 120.960 67.235 121.100 ;
        RECT 60.920 120.915 61.210 120.960 ;
        RECT 66.945 120.915 67.235 120.960 ;
        RECT 53.590 120.900 53.910 120.915 ;
        RECT 67.850 120.900 68.170 121.160 ;
        RECT 69.230 120.900 69.550 121.160 ;
        RECT 69.690 120.900 70.010 121.160 ;
        RECT 74.290 121.100 74.610 121.160 ;
        RECT 74.765 121.100 75.055 121.145 ;
        RECT 74.290 120.960 75.055 121.100 ;
        RECT 74.290 120.900 74.610 120.960 ;
        RECT 74.765 120.915 75.055 120.960 ;
        RECT 75.685 121.100 75.975 121.145 ;
        RECT 77.510 121.100 77.830 121.160 ;
        RECT 75.685 120.960 77.830 121.100 ;
        RECT 75.685 120.915 75.975 120.960 ;
        RECT 77.510 120.900 77.830 120.960 ;
        RECT 98.210 120.900 98.530 121.160 ;
        RECT 99.605 121.100 99.895 121.145 ;
        RECT 100.050 121.100 100.370 121.160 ;
        RECT 124.520 121.100 124.660 121.300 ;
        RECT 99.605 120.960 100.370 121.100 ;
        RECT 99.605 120.915 99.895 120.960 ;
        RECT 100.050 120.900 100.370 120.960 ;
        RECT 116.700 120.960 124.660 121.100 ;
        RECT 34.360 120.620 37.720 120.760 ;
        RECT 31.510 120.220 31.830 120.480 ;
        RECT 34.360 120.465 34.500 120.620 ;
        RECT 40.725 120.575 41.015 120.805 ;
        RECT 41.605 120.760 41.895 120.805 ;
        RECT 42.795 120.760 43.085 120.805 ;
        RECT 45.315 120.760 45.605 120.805 ;
        RECT 41.605 120.620 45.605 120.760 ;
        RECT 41.605 120.575 41.895 120.620 ;
        RECT 42.795 120.575 43.085 120.620 ;
        RECT 45.315 120.575 45.605 120.620 ;
        RECT 48.990 120.760 49.310 120.820 ;
        RECT 50.370 120.760 50.690 120.820 ;
        RECT 48.990 120.620 50.690 120.760 ;
        RECT 34.285 120.235 34.575 120.465 ;
        RECT 33.350 119.880 33.670 120.140 ;
        RECT 40.800 120.080 40.940 120.575 ;
        RECT 48.990 120.560 49.310 120.620 ;
        RECT 50.370 120.560 50.690 120.620 ;
        RECT 52.225 120.575 52.515 120.805 ;
        RECT 53.105 120.760 53.395 120.805 ;
        RECT 54.295 120.760 54.585 120.805 ;
        RECT 56.815 120.760 57.105 120.805 ;
        RECT 53.105 120.620 57.105 120.760 ;
        RECT 53.105 120.575 53.395 120.620 ;
        RECT 54.295 120.575 54.585 120.620 ;
        RECT 56.815 120.575 57.105 120.620 ;
        RECT 60.465 120.760 60.755 120.805 ;
        RECT 61.655 120.760 61.945 120.805 ;
        RECT 64.175 120.760 64.465 120.805 ;
        RECT 60.465 120.620 64.465 120.760 ;
        RECT 60.465 120.575 60.755 120.620 ;
        RECT 61.655 120.575 61.945 120.620 ;
        RECT 64.175 120.575 64.465 120.620 ;
        RECT 85.330 120.760 85.650 120.820 ;
        RECT 86.265 120.760 86.555 120.805 ;
        RECT 85.330 120.620 86.555 120.760 ;
        RECT 41.210 120.420 41.500 120.465 ;
        RECT 43.310 120.420 43.600 120.465 ;
        RECT 44.880 120.420 45.170 120.465 ;
        RECT 41.210 120.280 45.170 120.420 ;
        RECT 41.210 120.235 41.500 120.280 ;
        RECT 43.310 120.235 43.600 120.280 ;
        RECT 44.880 120.235 45.170 120.280 ;
        RECT 46.690 120.420 47.010 120.480 ;
        RECT 52.300 120.420 52.440 120.575 ;
        RECT 85.330 120.560 85.650 120.620 ;
        RECT 86.265 120.575 86.555 120.620 ;
        RECT 96.830 120.560 97.150 120.820 ;
        RECT 101.890 120.560 102.210 120.820 ;
        RECT 102.785 120.760 103.075 120.805 ;
        RECT 103.975 120.760 104.265 120.805 ;
        RECT 106.495 120.760 106.785 120.805 ;
        RECT 109.725 120.760 110.015 120.805 ;
        RECT 116.700 120.760 116.840 120.960 ;
        RECT 124.890 120.900 125.210 121.160 ;
        RECT 126.360 121.145 126.500 121.300 ;
        RECT 127.280 121.300 128.340 121.440 ;
        RECT 127.280 121.160 127.420 121.300 ;
        RECT 126.285 120.915 126.575 121.145 ;
        RECT 127.190 120.900 127.510 121.160 ;
        RECT 127.650 120.900 127.970 121.160 ;
        RECT 128.200 121.100 128.340 121.300 ;
        RECT 128.585 121.300 133.950 121.440 ;
        RECT 128.585 121.255 128.875 121.300 ;
        RECT 133.630 121.240 133.950 121.300 ;
        RECT 132.250 121.100 132.570 121.160 ;
        RECT 128.200 120.960 132.570 121.100 ;
        RECT 132.250 120.900 132.570 120.960 ;
        RECT 102.785 120.620 106.785 120.760 ;
        RECT 102.785 120.575 103.075 120.620 ;
        RECT 103.975 120.575 104.265 120.620 ;
        RECT 106.495 120.575 106.785 120.620 ;
        RECT 108.880 120.620 110.015 120.760 ;
        RECT 46.690 120.280 52.440 120.420 ;
        RECT 52.710 120.420 53.000 120.465 ;
        RECT 54.810 120.420 55.100 120.465 ;
        RECT 56.380 120.420 56.670 120.465 ;
        RECT 52.710 120.280 56.670 120.420 ;
        RECT 46.690 120.220 47.010 120.280 ;
        RECT 52.710 120.235 53.000 120.280 ;
        RECT 54.810 120.235 55.100 120.280 ;
        RECT 56.380 120.235 56.670 120.280 ;
        RECT 60.070 120.420 60.360 120.465 ;
        RECT 62.170 120.420 62.460 120.465 ;
        RECT 63.740 120.420 64.030 120.465 ;
        RECT 60.070 120.280 64.030 120.420 ;
        RECT 60.070 120.235 60.360 120.280 ;
        RECT 62.170 120.235 62.460 120.280 ;
        RECT 63.740 120.235 64.030 120.280 ;
        RECT 64.630 120.420 64.950 120.480 ;
        RECT 97.750 120.420 98.070 120.480 ;
        RECT 64.630 120.280 98.070 120.420 ;
        RECT 64.630 120.220 64.950 120.280 ;
        RECT 97.750 120.220 98.070 120.280 ;
        RECT 102.390 120.420 102.680 120.465 ;
        RECT 104.490 120.420 104.780 120.465 ;
        RECT 106.060 120.420 106.350 120.465 ;
        RECT 102.390 120.280 106.350 120.420 ;
        RECT 102.390 120.235 102.680 120.280 ;
        RECT 104.490 120.235 104.780 120.280 ;
        RECT 106.060 120.235 106.350 120.280 ;
        RECT 108.330 120.420 108.650 120.480 ;
        RECT 108.880 120.465 109.020 120.620 ;
        RECT 109.725 120.575 110.015 120.620 ;
        RECT 112.560 120.620 116.840 120.760 ;
        RECT 108.805 120.420 109.095 120.465 ;
        RECT 108.330 120.280 109.095 120.420 ;
        RECT 108.330 120.220 108.650 120.280 ;
        RECT 108.805 120.235 109.095 120.280 ;
        RECT 42.550 120.080 42.870 120.140 ;
        RECT 46.780 120.080 46.920 120.220 ;
        RECT 40.800 119.940 46.920 120.080 ;
        RECT 47.150 120.080 47.470 120.140 ;
        RECT 47.625 120.080 47.915 120.125 ;
        RECT 47.150 119.940 47.915 120.080 ;
        RECT 42.550 119.880 42.870 119.940 ;
        RECT 47.150 119.880 47.470 119.940 ;
        RECT 47.625 119.895 47.915 119.940 ;
        RECT 66.470 119.880 66.790 120.140 ;
        RECT 72.925 120.080 73.215 120.125 ;
        RECT 74.290 120.080 74.610 120.140 ;
        RECT 72.925 119.940 74.610 120.080 ;
        RECT 72.925 119.895 73.215 119.940 ;
        RECT 74.290 119.880 74.610 119.940 ;
        RECT 75.685 120.080 75.975 120.125 ;
        RECT 76.590 120.080 76.910 120.140 ;
        RECT 75.685 119.940 76.910 120.080 ;
        RECT 75.685 119.895 75.975 119.940 ;
        RECT 76.590 119.880 76.910 119.940 ;
        RECT 83.505 120.080 83.795 120.125 ;
        RECT 83.950 120.080 84.270 120.140 ;
        RECT 83.505 119.940 84.270 120.080 ;
        RECT 83.505 119.895 83.795 119.940 ;
        RECT 83.950 119.880 84.270 119.940 ;
        RECT 90.865 120.080 91.155 120.125 ;
        RECT 91.310 120.080 91.630 120.140 ;
        RECT 90.865 119.940 91.630 120.080 ;
        RECT 90.865 119.895 91.155 119.940 ;
        RECT 91.310 119.880 91.630 119.940 ;
        RECT 91.785 120.080 92.075 120.125 ;
        RECT 93.625 120.080 93.915 120.125 ;
        RECT 91.785 119.940 93.915 120.080 ;
        RECT 91.785 119.895 92.075 119.940 ;
        RECT 93.625 119.895 93.915 119.940 ;
        RECT 97.290 119.880 97.610 120.140 ;
        RECT 107.870 120.080 108.190 120.140 ;
        RECT 112.560 120.080 112.700 120.620 ;
        RECT 116.700 120.480 116.840 120.620 ;
        RECT 118.935 120.760 119.225 120.805 ;
        RECT 121.455 120.760 121.745 120.805 ;
        RECT 122.645 120.760 122.935 120.805 ;
        RECT 118.935 120.620 122.935 120.760 ;
        RECT 118.935 120.575 119.225 120.620 ;
        RECT 121.455 120.575 121.745 120.620 ;
        RECT 122.645 120.575 122.935 120.620 ;
        RECT 123.510 120.760 123.830 120.820 ;
        RECT 130.410 120.760 130.730 120.820 ;
        RECT 123.510 120.620 130.730 120.760 ;
        RECT 123.510 120.560 123.830 120.620 ;
        RECT 130.410 120.560 130.730 120.620 ;
        RECT 133.185 120.760 133.475 120.805 ;
        RECT 133.645 120.760 133.935 120.805 ;
        RECT 133.185 120.620 133.935 120.760 ;
        RECT 133.185 120.575 133.475 120.620 ;
        RECT 133.645 120.575 133.935 120.620 ;
        RECT 112.945 120.420 113.235 120.465 ;
        RECT 112.945 120.280 114.540 120.420 ;
        RECT 112.945 120.235 113.235 120.280 ;
        RECT 114.400 120.125 114.540 120.280 ;
        RECT 116.610 120.220 116.930 120.480 ;
        RECT 119.370 120.420 119.660 120.465 ;
        RECT 120.940 120.420 121.230 120.465 ;
        RECT 123.040 120.420 123.330 120.465 ;
        RECT 119.370 120.280 123.330 120.420 ;
        RECT 119.370 120.235 119.660 120.280 ;
        RECT 120.940 120.235 121.230 120.280 ;
        RECT 123.040 120.235 123.330 120.280 ;
        RECT 129.505 120.420 129.795 120.465 ;
        RECT 134.640 120.420 134.780 121.640 ;
        RECT 146.970 121.580 147.290 121.640 ;
        RECT 152.045 121.780 152.335 121.825 ;
        RECT 152.950 121.780 153.270 121.840 ;
        RECT 152.045 121.640 153.270 121.780 ;
        RECT 152.045 121.595 152.335 121.640 ;
        RECT 152.950 121.580 153.270 121.640 ;
        RECT 137.770 121.440 138.090 121.500 ;
        RECT 144.670 121.440 144.990 121.500 ;
        RECT 148.350 121.440 148.670 121.500 ;
        RECT 135.100 121.300 138.090 121.440 ;
        RECT 135.100 121.145 135.240 121.300 ;
        RECT 137.770 121.240 138.090 121.300 ;
        RECT 138.780 121.300 148.670 121.440 ;
        RECT 135.025 120.915 135.315 121.145 ;
        RECT 135.485 120.915 135.775 121.145 ;
        RECT 135.945 121.100 136.235 121.145 ;
        RECT 136.390 121.100 136.710 121.160 ;
        RECT 138.780 121.145 138.920 121.300 ;
        RECT 144.670 121.240 144.990 121.300 ;
        RECT 148.350 121.240 148.670 121.300 ;
        RECT 149.360 121.300 154.560 121.440 ;
        RECT 149.360 121.145 149.500 121.300 ;
        RECT 154.420 121.160 154.560 121.300 ;
        RECT 135.945 120.960 136.710 121.100 ;
        RECT 135.945 120.915 136.235 120.960 ;
        RECT 129.505 120.280 134.780 120.420 ;
        RECT 135.010 120.420 135.330 120.480 ;
        RECT 135.560 120.420 135.700 120.915 ;
        RECT 136.390 120.900 136.710 120.960 ;
        RECT 136.865 121.100 137.155 121.145 ;
        RECT 137.325 121.100 137.615 121.145 ;
        RECT 136.865 120.960 137.615 121.100 ;
        RECT 136.865 120.915 137.155 120.960 ;
        RECT 137.325 120.915 137.615 120.960 ;
        RECT 138.245 120.915 138.535 121.145 ;
        RECT 138.705 120.915 138.995 121.145 ;
        RECT 139.165 121.100 139.455 121.145 ;
        RECT 139.165 120.960 140.300 121.100 ;
        RECT 139.165 120.915 139.455 120.960 ;
        RECT 136.940 120.760 137.080 120.915 ;
        RECT 136.480 120.620 137.080 120.760 ;
        RECT 136.480 120.480 136.620 120.620 ;
        RECT 135.010 120.280 135.700 120.420 ;
        RECT 129.505 120.235 129.795 120.280 ;
        RECT 135.010 120.220 135.330 120.280 ;
        RECT 107.870 119.940 112.700 120.080 ;
        RECT 107.870 119.880 108.190 119.940 ;
        RECT 114.325 119.895 114.615 120.125 ;
        RECT 135.560 120.080 135.700 120.280 ;
        RECT 136.390 120.220 136.710 120.480 ;
        RECT 136.850 120.420 137.170 120.480 ;
        RECT 138.320 120.420 138.460 120.915 ;
        RECT 136.850 120.280 138.460 120.420 ;
        RECT 136.850 120.220 137.170 120.280 ;
        RECT 138.780 120.080 138.920 120.915 ;
        RECT 135.560 119.940 138.920 120.080 ;
        RECT 140.160 120.080 140.300 120.960 ;
        RECT 149.285 120.915 149.575 121.145 ;
        RECT 150.665 121.100 150.955 121.145 ;
        RECT 152.950 121.100 153.270 121.160 ;
        RECT 150.665 120.960 153.270 121.100 ;
        RECT 150.665 120.915 150.955 120.960 ;
        RECT 152.950 120.900 153.270 120.960 ;
        RECT 154.330 121.100 154.650 121.160 ;
        RECT 154.805 121.100 155.095 121.145 ;
        RECT 154.330 120.960 155.095 121.100 ;
        RECT 154.330 120.900 154.650 120.960 ;
        RECT 154.805 120.915 155.095 120.960 ;
        RECT 144.210 120.560 144.530 120.820 ;
        RECT 147.445 120.575 147.735 120.805 ;
        RECT 150.205 120.760 150.495 120.805 ;
        RECT 155.250 120.760 155.570 120.820 ;
        RECT 150.205 120.620 155.570 120.760 ;
        RECT 150.205 120.575 150.495 120.620 ;
        RECT 140.545 120.420 140.835 120.465 ;
        RECT 147.520 120.420 147.660 120.575 ;
        RECT 155.250 120.560 155.570 120.620 ;
        RECT 140.545 120.280 147.660 120.420 ;
        RECT 140.545 120.235 140.835 120.280 ;
        RECT 141.005 120.080 141.295 120.125 ;
        RECT 141.450 120.080 141.770 120.140 ;
        RECT 140.160 119.940 141.770 120.080 ;
        RECT 141.005 119.895 141.295 119.940 ;
        RECT 141.450 119.880 141.770 119.940 ;
        RECT 144.670 119.880 144.990 120.140 ;
        RECT 145.130 120.080 145.450 120.140 ;
        RECT 148.365 120.080 148.655 120.125 ;
        RECT 145.130 119.940 148.655 120.080 ;
        RECT 145.130 119.880 145.450 119.940 ;
        RECT 148.365 119.895 148.655 119.940 ;
        RECT 150.665 120.080 150.955 120.125 ;
        RECT 151.110 120.080 151.430 120.140 ;
        RECT 150.665 119.940 151.430 120.080 ;
        RECT 150.665 119.895 150.955 119.940 ;
        RECT 151.110 119.880 151.430 119.940 ;
        RECT 22.700 119.260 157.020 119.740 ;
        RECT 26.925 119.060 27.215 119.105 ;
        RECT 29.210 119.060 29.530 119.120 ;
        RECT 26.925 118.920 29.530 119.060 ;
        RECT 26.925 118.875 27.215 118.920 ;
        RECT 29.210 118.860 29.530 118.920 ;
        RECT 42.550 119.060 42.870 119.120 ;
        RECT 43.945 119.060 44.235 119.105 ;
        RECT 42.550 118.920 44.235 119.060 ;
        RECT 42.550 118.860 42.870 118.920 ;
        RECT 43.945 118.875 44.235 118.920 ;
        RECT 45.770 119.060 46.090 119.120 ;
        RECT 53.605 119.060 53.895 119.105 ;
        RECT 54.050 119.060 54.370 119.120 ;
        RECT 45.770 118.920 48.760 119.060 ;
        RECT 28.290 118.720 28.610 118.780 ;
        RECT 29.685 118.720 29.975 118.765 ;
        RECT 28.290 118.580 29.975 118.720 ;
        RECT 28.290 118.520 28.610 118.580 ;
        RECT 29.685 118.535 29.975 118.580 ;
        RECT 30.130 118.720 30.450 118.780 ;
        RECT 34.730 118.720 35.050 118.780 ;
        RECT 38.410 118.720 38.730 118.780 ;
        RECT 44.020 118.720 44.160 118.875 ;
        RECT 45.770 118.860 46.090 118.920 ;
        RECT 47.150 118.720 47.470 118.780 ;
        RECT 48.620 118.720 48.760 118.920 ;
        RECT 53.605 118.920 54.370 119.060 ;
        RECT 53.605 118.875 53.895 118.920 ;
        RECT 54.050 118.860 54.370 118.920 ;
        RECT 64.645 119.060 64.935 119.105 ;
        RECT 66.025 119.060 66.315 119.105 ;
        RECT 64.645 118.920 66.315 119.060 ;
        RECT 64.645 118.875 64.935 118.920 ;
        RECT 66.025 118.875 66.315 118.920 ;
        RECT 71.530 119.060 71.850 119.120 ;
        RECT 72.005 119.060 72.295 119.105 ;
        RECT 71.530 118.920 72.295 119.060 ;
        RECT 71.530 118.860 71.850 118.920 ;
        RECT 72.005 118.875 72.295 118.920 ;
        RECT 73.385 119.060 73.675 119.105 ;
        RECT 74.290 119.060 74.610 119.120 ;
        RECT 73.385 118.920 74.610 119.060 ;
        RECT 73.385 118.875 73.675 118.920 ;
        RECT 74.290 118.860 74.610 118.920 ;
        RECT 80.730 119.060 81.050 119.120 ;
        RECT 83.030 119.060 83.350 119.120 ;
        RECT 80.730 118.920 83.350 119.060 ;
        RECT 80.730 118.860 81.050 118.920 ;
        RECT 83.030 118.860 83.350 118.920 ;
        RECT 83.950 118.860 84.270 119.120 ;
        RECT 97.750 119.060 98.070 119.120 ;
        RECT 102.825 119.060 103.115 119.105 ;
        RECT 103.730 119.060 104.050 119.120 ;
        RECT 105.110 119.060 105.430 119.120 ;
        RECT 97.750 118.920 100.740 119.060 ;
        RECT 97.750 118.860 98.070 118.920 ;
        RECT 54.525 118.720 54.815 118.765 ;
        RECT 30.130 118.580 35.050 118.720 ;
        RECT 30.130 118.520 30.450 118.580 ;
        RECT 34.730 118.520 35.050 118.580 ;
        RECT 37.120 118.580 43.240 118.720 ;
        RECT 44.020 118.580 47.840 118.720 ;
        RECT 48.620 118.580 54.815 118.720 ;
        RECT 28.750 118.180 29.070 118.440 ;
        RECT 29.210 118.180 29.530 118.440 ;
        RECT 27.830 117.840 28.150 118.100 ;
        RECT 29.685 118.040 29.975 118.085 ;
        RECT 30.220 118.040 30.360 118.520 ;
        RECT 29.685 117.900 30.360 118.040 ;
        RECT 31.065 118.040 31.355 118.085 ;
        RECT 31.510 118.040 31.830 118.100 ;
        RECT 31.065 117.900 31.830 118.040 ;
        RECT 29.685 117.855 29.975 117.900 ;
        RECT 31.065 117.855 31.355 117.900 ;
        RECT 31.510 117.840 31.830 117.900 ;
        RECT 33.810 117.840 34.130 118.100 ;
        RECT 37.120 118.085 37.260 118.580 ;
        RECT 38.410 118.520 38.730 118.580 ;
        RECT 42.550 118.180 42.870 118.440 ;
        RECT 43.100 118.380 43.240 118.580 ;
        RECT 47.150 118.520 47.470 118.580 ;
        RECT 47.700 118.425 47.840 118.580 ;
        RECT 54.525 118.535 54.815 118.580 ;
        RECT 65.565 118.720 65.855 118.765 ;
        RECT 67.850 118.720 68.170 118.780 ;
        RECT 65.565 118.580 68.170 118.720 ;
        RECT 65.565 118.535 65.855 118.580 ;
        RECT 67.850 118.520 68.170 118.580 ;
        RECT 68.310 118.720 68.630 118.780 ;
        RECT 70.150 118.720 70.470 118.780 ;
        RECT 73.830 118.720 74.150 118.780 ;
        RECT 68.310 118.580 74.150 118.720 ;
        RECT 68.310 118.520 68.630 118.580 ;
        RECT 70.150 118.520 70.470 118.580 ;
        RECT 73.830 118.520 74.150 118.580 ;
        RECT 76.170 118.720 76.460 118.765 ;
        RECT 78.270 118.720 78.560 118.765 ;
        RECT 79.840 118.720 80.130 118.765 ;
        RECT 76.170 118.580 80.130 118.720 ;
        RECT 76.170 118.535 76.460 118.580 ;
        RECT 78.270 118.535 78.560 118.580 ;
        RECT 79.840 118.535 80.130 118.580 ;
        RECT 82.585 118.720 82.875 118.765 ;
        RECT 85.330 118.720 85.650 118.780 ;
        RECT 82.585 118.580 85.650 118.720 ;
        RECT 82.585 118.535 82.875 118.580 ;
        RECT 85.330 118.520 85.650 118.580 ;
        RECT 88.130 118.720 88.420 118.765 ;
        RECT 90.230 118.720 90.520 118.765 ;
        RECT 91.800 118.720 92.090 118.765 ;
        RECT 88.130 118.580 92.090 118.720 ;
        RECT 88.130 118.535 88.420 118.580 ;
        RECT 90.230 118.535 90.520 118.580 ;
        RECT 91.800 118.535 92.090 118.580 ;
        RECT 96.410 118.720 96.700 118.765 ;
        RECT 98.510 118.720 98.800 118.765 ;
        RECT 100.080 118.720 100.370 118.765 ;
        RECT 96.410 118.580 100.370 118.720 ;
        RECT 100.600 118.720 100.740 118.920 ;
        RECT 102.825 118.920 105.430 119.060 ;
        RECT 102.825 118.875 103.115 118.920 ;
        RECT 103.730 118.860 104.050 118.920 ;
        RECT 105.110 118.860 105.430 118.920 ;
        RECT 105.660 118.920 118.220 119.060 ;
        RECT 105.660 118.720 105.800 118.920 ;
        RECT 100.600 118.580 105.800 118.720 ;
        RECT 113.890 118.720 114.180 118.765 ;
        RECT 115.990 118.720 116.280 118.765 ;
        RECT 117.560 118.720 117.850 118.765 ;
        RECT 113.890 118.580 117.850 118.720 ;
        RECT 118.080 118.720 118.220 118.920 ;
        RECT 121.670 118.860 121.990 119.120 ;
        RECT 134.090 119.060 134.410 119.120 ;
        RECT 135.010 119.060 135.330 119.120 ;
        RECT 122.220 118.920 128.800 119.060 ;
        RECT 122.220 118.720 122.360 118.920 ;
        RECT 118.080 118.580 122.360 118.720 ;
        RECT 124.010 118.720 124.300 118.765 ;
        RECT 126.110 118.720 126.400 118.765 ;
        RECT 127.680 118.720 127.970 118.765 ;
        RECT 124.010 118.580 127.970 118.720 ;
        RECT 96.410 118.535 96.700 118.580 ;
        RECT 98.510 118.535 98.800 118.580 ;
        RECT 100.080 118.535 100.370 118.580 ;
        RECT 113.890 118.535 114.180 118.580 ;
        RECT 115.990 118.535 116.280 118.580 ;
        RECT 117.560 118.535 117.850 118.580 ;
        RECT 124.010 118.535 124.300 118.580 ;
        RECT 126.110 118.535 126.400 118.580 ;
        RECT 127.680 118.535 127.970 118.580 ;
        RECT 44.405 118.380 44.695 118.425 ;
        RECT 43.100 118.240 44.695 118.380 ;
        RECT 44.405 118.195 44.695 118.240 ;
        RECT 47.625 118.195 47.915 118.425 ;
        RECT 50.845 118.380 51.135 118.425 ;
        RECT 55.445 118.380 55.735 118.425 ;
        RECT 64.630 118.380 64.950 118.440 ;
        RECT 50.845 118.240 54.280 118.380 ;
        RECT 50.845 118.195 51.135 118.240 ;
        RECT 37.045 117.855 37.335 118.085 ;
        RECT 38.425 118.040 38.715 118.085 ;
        RECT 37.580 117.900 38.715 118.040 ;
        RECT 31.600 117.700 31.740 117.840 ;
        RECT 34.270 117.700 34.590 117.760 ;
        RECT 37.580 117.700 37.720 117.900 ;
        RECT 38.425 117.855 38.715 117.900 ;
        RECT 41.630 117.840 41.950 118.100 ;
        RECT 42.105 117.855 42.395 118.085 ;
        RECT 43.025 118.040 43.315 118.085 ;
        RECT 43.470 118.040 43.790 118.100 ;
        RECT 43.025 117.900 43.790 118.040 ;
        RECT 43.025 117.855 43.315 117.900 ;
        RECT 31.600 117.560 37.720 117.700 ;
        RECT 37.950 117.700 38.270 117.760 ;
        RECT 42.180 117.700 42.320 117.855 ;
        RECT 43.470 117.840 43.790 117.900 ;
        RECT 45.325 117.855 45.615 118.085 ;
        RECT 43.930 117.700 44.250 117.760 ;
        RECT 37.950 117.560 41.860 117.700 ;
        RECT 42.180 117.560 44.250 117.700 ;
        RECT 34.270 117.500 34.590 117.560 ;
        RECT 37.950 117.500 38.270 117.560 ;
        RECT 30.605 117.360 30.895 117.405 ;
        RECT 31.050 117.360 31.370 117.420 ;
        RECT 30.605 117.220 31.370 117.360 ;
        RECT 30.605 117.175 30.895 117.220 ;
        RECT 31.050 117.160 31.370 117.220 ;
        RECT 32.890 117.160 33.210 117.420 ;
        RECT 36.110 117.160 36.430 117.420 ;
        RECT 40.725 117.360 41.015 117.405 ;
        RECT 41.170 117.360 41.490 117.420 ;
        RECT 40.725 117.220 41.490 117.360 ;
        RECT 41.720 117.360 41.860 117.560 ;
        RECT 43.930 117.500 44.250 117.560 ;
        RECT 45.400 117.360 45.540 117.855 ;
        RECT 51.750 117.840 52.070 118.100 ;
        RECT 52.670 117.840 52.990 118.100 ;
        RECT 54.140 118.085 54.280 118.240 ;
        RECT 55.445 118.240 64.950 118.380 ;
        RECT 55.445 118.195 55.735 118.240 ;
        RECT 64.630 118.180 64.950 118.240 ;
        RECT 66.470 118.380 66.790 118.440 ;
        RECT 67.390 118.380 67.710 118.440 ;
        RECT 68.785 118.380 69.075 118.425 ;
        RECT 66.470 118.240 69.075 118.380 ;
        RECT 66.470 118.180 66.790 118.240 ;
        RECT 67.390 118.180 67.710 118.240 ;
        RECT 68.785 118.195 69.075 118.240 ;
        RECT 69.230 118.380 69.550 118.440 ;
        RECT 76.565 118.380 76.855 118.425 ;
        RECT 77.755 118.380 78.045 118.425 ;
        RECT 80.275 118.380 80.565 118.425 ;
        RECT 88.525 118.380 88.815 118.425 ;
        RECT 89.715 118.380 90.005 118.425 ;
        RECT 92.235 118.380 92.525 118.425 ;
        RECT 69.230 118.240 74.980 118.380 ;
        RECT 69.230 118.180 69.550 118.240 ;
        RECT 69.780 118.085 69.920 118.240 ;
        RECT 54.065 117.855 54.355 118.085 ;
        RECT 69.705 118.040 69.995 118.085 ;
        RECT 71.085 118.040 71.375 118.085 ;
        RECT 69.705 117.900 70.105 118.040 ;
        RECT 71.085 117.900 72.680 118.040 ;
        RECT 69.705 117.855 69.995 117.900 ;
        RECT 71.085 117.855 71.375 117.900 ;
        RECT 63.725 117.700 64.015 117.745 ;
        RECT 64.170 117.700 64.490 117.760 ;
        RECT 68.310 117.700 68.630 117.760 ;
        RECT 63.725 117.560 68.630 117.700 ;
        RECT 63.725 117.515 64.015 117.560 ;
        RECT 64.170 117.500 64.490 117.560 ;
        RECT 68.310 117.500 68.630 117.560 ;
        RECT 41.720 117.220 45.540 117.360 ;
        RECT 46.245 117.360 46.535 117.405 ;
        RECT 49.910 117.360 50.230 117.420 ;
        RECT 46.245 117.220 50.230 117.360 ;
        RECT 40.725 117.175 41.015 117.220 ;
        RECT 41.170 117.160 41.490 117.220 ;
        RECT 46.245 117.175 46.535 117.220 ;
        RECT 49.910 117.160 50.230 117.220 ;
        RECT 50.830 117.360 51.150 117.420 ;
        RECT 55.445 117.360 55.735 117.405 ;
        RECT 50.830 117.220 55.735 117.360 ;
        RECT 50.830 117.160 51.150 117.220 ;
        RECT 55.445 117.175 55.735 117.220 ;
        RECT 64.775 117.360 65.065 117.405 ;
        RECT 68.770 117.360 69.090 117.420 ;
        RECT 64.775 117.220 69.090 117.360 ;
        RECT 64.775 117.175 65.065 117.220 ;
        RECT 68.770 117.160 69.090 117.220 ;
        RECT 70.165 117.360 70.455 117.405 ;
        RECT 71.530 117.360 71.850 117.420 ;
        RECT 72.540 117.405 72.680 117.900 ;
        RECT 73.830 117.700 74.150 117.760 ;
        RECT 74.305 117.700 74.595 117.745 ;
        RECT 73.830 117.560 74.595 117.700 ;
        RECT 74.840 117.700 74.980 118.240 ;
        RECT 76.565 118.240 80.565 118.380 ;
        RECT 76.565 118.195 76.855 118.240 ;
        RECT 77.755 118.195 78.045 118.240 ;
        RECT 80.275 118.195 80.565 118.240 ;
        RECT 80.775 118.240 87.860 118.380 ;
        RECT 75.685 118.040 75.975 118.085 ;
        RECT 79.350 118.040 79.670 118.100 ;
        RECT 80.775 118.040 80.915 118.240 ;
        RECT 75.685 117.900 80.915 118.040 ;
        RECT 75.685 117.855 75.975 117.900 ;
        RECT 79.350 117.840 79.670 117.900 ;
        RECT 85.330 117.840 85.650 118.100 ;
        RECT 86.265 118.040 86.555 118.085 ;
        RECT 87.170 118.040 87.490 118.100 ;
        RECT 87.720 118.085 87.860 118.240 ;
        RECT 88.525 118.240 92.525 118.380 ;
        RECT 88.525 118.195 88.815 118.240 ;
        RECT 89.715 118.195 90.005 118.240 ;
        RECT 92.235 118.195 92.525 118.240 ;
        RECT 96.805 118.380 97.095 118.425 ;
        RECT 97.995 118.380 98.285 118.425 ;
        RECT 100.515 118.380 100.805 118.425 ;
        RECT 96.805 118.240 100.805 118.380 ;
        RECT 96.805 118.195 97.095 118.240 ;
        RECT 97.995 118.195 98.285 118.240 ;
        RECT 100.515 118.195 100.805 118.240 ;
        RECT 101.890 118.380 102.210 118.440 ;
        RECT 113.405 118.380 113.695 118.425 ;
        RECT 101.890 118.240 113.695 118.380 ;
        RECT 101.890 118.180 102.210 118.240 ;
        RECT 113.405 118.195 113.695 118.240 ;
        RECT 114.285 118.380 114.575 118.425 ;
        RECT 115.475 118.380 115.765 118.425 ;
        RECT 117.995 118.380 118.285 118.425 ;
        RECT 114.285 118.240 118.285 118.380 ;
        RECT 114.285 118.195 114.575 118.240 ;
        RECT 115.475 118.195 115.765 118.240 ;
        RECT 117.995 118.195 118.285 118.240 ;
        RECT 123.510 118.180 123.830 118.440 ;
        RECT 124.405 118.380 124.695 118.425 ;
        RECT 125.595 118.380 125.885 118.425 ;
        RECT 128.115 118.380 128.405 118.425 ;
        RECT 124.405 118.240 128.405 118.380 ;
        RECT 128.660 118.380 128.800 118.920 ;
        RECT 134.090 118.920 135.330 119.060 ;
        RECT 134.090 118.860 134.410 118.920 ;
        RECT 135.010 118.860 135.330 118.920 ;
        RECT 139.165 119.060 139.455 119.105 ;
        RECT 144.210 119.060 144.530 119.120 ;
        RECT 139.165 118.920 144.530 119.060 ;
        RECT 139.165 118.875 139.455 118.920 ;
        RECT 144.210 118.860 144.530 118.920 ;
        RECT 155.250 118.860 155.570 119.120 ;
        RECT 130.425 118.720 130.715 118.765 ;
        RECT 138.690 118.720 139.010 118.780 ;
        RECT 130.425 118.580 139.010 118.720 ;
        RECT 130.425 118.535 130.715 118.580 ;
        RECT 133.170 118.380 133.490 118.440 ;
        RECT 136.390 118.380 136.710 118.440 ;
        RECT 137.860 118.425 138.000 118.580 ;
        RECT 138.690 118.520 139.010 118.580 ;
        RECT 141.910 118.720 142.200 118.765 ;
        RECT 143.480 118.720 143.770 118.765 ;
        RECT 145.580 118.720 145.870 118.765 ;
        RECT 141.910 118.580 145.870 118.720 ;
        RECT 141.910 118.535 142.200 118.580 ;
        RECT 143.480 118.535 143.770 118.580 ;
        RECT 145.580 118.535 145.870 118.580 ;
        RECT 148.850 118.720 149.140 118.765 ;
        RECT 150.950 118.720 151.240 118.765 ;
        RECT 152.520 118.720 152.810 118.765 ;
        RECT 148.850 118.580 152.810 118.720 ;
        RECT 148.850 118.535 149.140 118.580 ;
        RECT 150.950 118.535 151.240 118.580 ;
        RECT 152.520 118.535 152.810 118.580 ;
        RECT 128.660 118.240 136.710 118.380 ;
        RECT 124.405 118.195 124.695 118.240 ;
        RECT 125.595 118.195 125.885 118.240 ;
        RECT 128.115 118.195 128.405 118.240 ;
        RECT 86.265 117.900 87.490 118.040 ;
        RECT 86.265 117.855 86.555 117.900 ;
        RECT 87.170 117.840 87.490 117.900 ;
        RECT 87.645 118.040 87.935 118.085 ;
        RECT 93.150 118.040 93.470 118.100 ;
        RECT 95.925 118.040 96.215 118.085 ;
        RECT 101.980 118.040 102.120 118.180 ;
        RECT 87.645 117.900 102.120 118.040 ;
        RECT 87.645 117.855 87.935 117.900 ;
        RECT 93.150 117.840 93.470 117.900 ;
        RECT 95.925 117.855 96.215 117.900 ;
        RECT 107.870 117.840 108.190 118.100 ;
        RECT 108.330 117.840 108.650 118.100 ;
        RECT 112.485 118.040 112.775 118.085 ;
        RECT 112.930 118.040 113.250 118.100 ;
        RECT 112.485 117.900 113.250 118.040 ;
        RECT 112.485 117.855 112.775 117.900 ;
        RECT 112.930 117.840 113.250 117.900 ;
        RECT 116.610 118.040 116.930 118.100 ;
        RECT 120.765 118.040 121.055 118.085 ;
        RECT 116.610 117.900 121.055 118.040 ;
        RECT 116.610 117.840 116.930 117.900 ;
        RECT 120.765 117.855 121.055 117.900 ;
        RECT 121.685 118.040 121.975 118.085 ;
        RECT 127.190 118.040 127.510 118.100 ;
        RECT 121.685 117.900 127.510 118.040 ;
        RECT 121.685 117.855 121.975 117.900 ;
        RECT 127.190 117.840 127.510 117.900 ;
        RECT 129.030 118.040 129.350 118.100 ;
        RECT 132.340 118.085 132.480 118.240 ;
        RECT 133.170 118.180 133.490 118.240 ;
        RECT 136.390 118.180 136.710 118.240 ;
        RECT 137.785 118.195 138.075 118.425 ;
        RECT 141.475 118.380 141.765 118.425 ;
        RECT 143.995 118.380 144.285 118.425 ;
        RECT 145.185 118.380 145.475 118.425 ;
        RECT 141.475 118.240 145.475 118.380 ;
        RECT 141.475 118.195 141.765 118.240 ;
        RECT 143.995 118.195 144.285 118.240 ;
        RECT 145.185 118.195 145.475 118.240 ;
        RECT 146.065 118.380 146.355 118.425 ;
        RECT 147.890 118.380 148.210 118.440 ;
        RECT 148.365 118.380 148.655 118.425 ;
        RECT 146.065 118.240 148.655 118.380 ;
        RECT 146.065 118.195 146.355 118.240 ;
        RECT 147.890 118.180 148.210 118.240 ;
        RECT 148.365 118.195 148.655 118.240 ;
        RECT 149.245 118.380 149.535 118.425 ;
        RECT 150.435 118.380 150.725 118.425 ;
        RECT 152.955 118.380 153.245 118.425 ;
        RECT 149.245 118.240 153.245 118.380 ;
        RECT 149.245 118.195 149.535 118.240 ;
        RECT 150.435 118.195 150.725 118.240 ;
        RECT 152.955 118.195 153.245 118.240 ;
        RECT 144.670 118.085 144.990 118.100 ;
        RECT 129.030 117.900 131.560 118.040 ;
        RECT 129.030 117.840 129.350 117.900 ;
        RECT 77.020 117.700 77.310 117.745 ;
        RECT 77.510 117.700 77.830 117.760 ;
        RECT 74.840 117.560 76.820 117.700 ;
        RECT 73.830 117.500 74.150 117.560 ;
        RECT 74.305 117.515 74.595 117.560 ;
        RECT 76.680 117.420 76.820 117.560 ;
        RECT 77.020 117.560 77.830 117.700 ;
        RECT 77.020 117.515 77.310 117.560 ;
        RECT 77.510 117.500 77.830 117.560 ;
        RECT 82.110 117.700 82.430 117.760 ;
        RECT 83.805 117.700 84.095 117.745 ;
        RECT 84.410 117.700 84.730 117.760 ;
        RECT 82.110 117.560 84.730 117.700 ;
        RECT 82.110 117.500 82.430 117.560 ;
        RECT 83.805 117.515 84.095 117.560 ;
        RECT 84.410 117.500 84.730 117.560 ;
        RECT 84.870 117.500 85.190 117.760 ;
        RECT 88.980 117.700 89.270 117.745 ;
        RECT 90.850 117.700 91.170 117.760 ;
        RECT 97.290 117.745 97.610 117.760 ;
        RECT 97.260 117.700 97.610 117.745 ;
        RECT 100.510 117.700 100.830 117.760 ;
        RECT 88.980 117.560 91.170 117.700 ;
        RECT 97.095 117.560 97.610 117.700 ;
        RECT 88.980 117.515 89.270 117.560 ;
        RECT 90.850 117.500 91.170 117.560 ;
        RECT 97.260 117.515 97.610 117.560 ;
        RECT 97.290 117.500 97.610 117.515 ;
        RECT 97.840 117.560 100.830 117.700 ;
        RECT 70.165 117.220 71.850 117.360 ;
        RECT 70.165 117.175 70.455 117.220 ;
        RECT 71.530 117.160 71.850 117.220 ;
        RECT 72.465 117.175 72.755 117.405 ;
        RECT 73.305 117.360 73.595 117.405 ;
        RECT 74.750 117.360 75.070 117.420 ;
        RECT 73.305 117.220 75.070 117.360 ;
        RECT 73.305 117.175 73.595 117.220 ;
        RECT 74.750 117.160 75.070 117.220 ;
        RECT 76.590 117.160 76.910 117.420 ;
        RECT 78.430 117.360 78.750 117.420 ;
        RECT 83.045 117.360 83.335 117.405 ;
        RECT 78.430 117.220 83.335 117.360 ;
        RECT 78.430 117.160 78.750 117.220 ;
        RECT 83.045 117.175 83.335 117.220 ;
        RECT 85.330 117.360 85.650 117.420 ;
        RECT 85.805 117.360 86.095 117.405 ;
        RECT 85.330 117.220 86.095 117.360 ;
        RECT 85.330 117.160 85.650 117.220 ;
        RECT 85.805 117.175 86.095 117.220 ;
        RECT 94.545 117.360 94.835 117.405 ;
        RECT 96.830 117.360 97.150 117.420 ;
        RECT 97.840 117.360 97.980 117.560 ;
        RECT 100.510 117.500 100.830 117.560 ;
        RECT 109.710 117.500 110.030 117.760 ;
        RECT 110.185 117.700 110.475 117.745 ;
        RECT 112.025 117.700 112.315 117.745 ;
        RECT 110.185 117.560 112.315 117.700 ;
        RECT 110.185 117.515 110.475 117.560 ;
        RECT 112.025 117.515 112.315 117.560 ;
        RECT 114.740 117.700 115.030 117.745 ;
        RECT 116.150 117.700 116.470 117.760 ;
        RECT 114.740 117.560 116.470 117.700 ;
        RECT 114.740 117.515 115.030 117.560 ;
        RECT 116.150 117.500 116.470 117.560 ;
        RECT 124.860 117.700 125.150 117.745 ;
        RECT 130.885 117.700 131.175 117.745 ;
        RECT 124.860 117.560 131.175 117.700 ;
        RECT 131.420 117.700 131.560 117.900 ;
        RECT 132.265 117.855 132.555 118.085 ;
        RECT 134.565 118.040 134.855 118.085 ;
        RECT 135.025 118.040 135.315 118.085 ;
        RECT 134.565 117.900 135.315 118.040 ;
        RECT 134.565 117.855 134.855 117.900 ;
        RECT 135.025 117.855 135.315 117.900 ;
        RECT 144.670 118.040 145.020 118.085 ;
        RECT 151.110 118.040 151.430 118.100 ;
        RECT 144.670 117.900 145.185 118.040 ;
        RECT 145.680 117.900 151.430 118.040 ;
        RECT 144.670 117.855 145.020 117.900 ;
        RECT 144.670 117.840 144.990 117.855 ;
        RECT 132.725 117.700 133.015 117.745 ;
        RECT 131.420 117.560 133.015 117.700 ;
        RECT 124.860 117.515 125.150 117.560 ;
        RECT 130.885 117.515 131.175 117.560 ;
        RECT 132.725 117.515 133.015 117.560 ;
        RECT 133.630 117.700 133.950 117.760 ;
        RECT 145.680 117.700 145.820 117.900 ;
        RECT 151.110 117.840 151.430 117.900 ;
        RECT 133.630 117.560 145.820 117.700 ;
        RECT 146.050 117.700 146.370 117.760 ;
        RECT 149.590 117.700 149.880 117.745 ;
        RECT 146.050 117.560 149.880 117.700 ;
        RECT 133.630 117.500 133.950 117.560 ;
        RECT 146.050 117.500 146.370 117.560 ;
        RECT 149.590 117.515 149.880 117.560 ;
        RECT 94.545 117.220 97.980 117.360 ;
        RECT 99.130 117.360 99.450 117.420 ;
        RECT 106.965 117.360 107.255 117.405 ;
        RECT 99.130 117.220 107.255 117.360 ;
        RECT 94.545 117.175 94.835 117.220 ;
        RECT 96.830 117.160 97.150 117.220 ;
        RECT 99.130 117.160 99.450 117.220 ;
        RECT 106.965 117.175 107.255 117.220 ;
        RECT 120.290 117.160 120.610 117.420 ;
        RECT 133.170 117.160 133.490 117.420 ;
        RECT 136.390 117.360 136.710 117.420 ;
        RECT 150.190 117.360 150.510 117.420 ;
        RECT 136.390 117.220 150.510 117.360 ;
        RECT 136.390 117.160 136.710 117.220 ;
        RECT 150.190 117.160 150.510 117.220 ;
        RECT 22.700 116.540 157.820 117.020 ;
        RECT 30.590 116.340 30.910 116.400 ;
        RECT 30.590 116.200 33.580 116.340 ;
        RECT 30.590 116.140 30.910 116.200 ;
        RECT 26.910 116.000 27.230 116.060 ;
        RECT 32.890 116.045 33.210 116.060 ;
        RECT 32.860 116.000 33.210 116.045 ;
        RECT 24.240 115.860 31.740 116.000 ;
        RECT 32.695 115.860 33.210 116.000 ;
        RECT 33.440 116.000 33.580 116.200 ;
        RECT 38.410 116.140 38.730 116.400 ;
        RECT 41.630 116.340 41.950 116.400 ;
        RECT 45.770 116.340 46.090 116.400 ;
        RECT 74.765 116.340 75.055 116.385 ;
        RECT 41.630 116.200 46.090 116.340 ;
        RECT 41.630 116.140 41.950 116.200 ;
        RECT 45.770 116.140 46.090 116.200 ;
        RECT 67.480 116.200 75.055 116.340 ;
        RECT 58.650 116.000 58.970 116.060 ;
        RECT 33.440 115.860 58.970 116.000 ;
        RECT 24.240 115.705 24.380 115.860 ;
        RECT 26.910 115.800 27.230 115.860 ;
        RECT 25.530 115.705 25.850 115.720 ;
        RECT 31.600 115.705 31.740 115.860 ;
        RECT 32.860 115.815 33.210 115.860 ;
        RECT 32.890 115.800 33.210 115.815 ;
        RECT 58.650 115.800 58.970 115.860 ;
        RECT 66.180 116.000 66.470 116.045 ;
        RECT 67.480 116.000 67.620 116.200 ;
        RECT 74.765 116.155 75.055 116.200 ;
        RECT 77.510 116.140 77.830 116.400 ;
        RECT 79.365 116.340 79.655 116.385 ;
        RECT 81.190 116.340 81.510 116.400 ;
        RECT 79.365 116.200 81.510 116.340 ;
        RECT 79.365 116.155 79.655 116.200 ;
        RECT 81.190 116.140 81.510 116.200 ;
        RECT 87.170 116.140 87.490 116.400 ;
        RECT 89.025 116.340 89.315 116.385 ;
        RECT 90.850 116.340 91.170 116.400 ;
        RECT 89.025 116.200 91.170 116.340 ;
        RECT 89.025 116.155 89.315 116.200 ;
        RECT 90.850 116.140 91.170 116.200 ;
        RECT 91.310 116.140 91.630 116.400 ;
        RECT 98.210 116.140 98.530 116.400 ;
        RECT 116.150 116.140 116.470 116.400 ;
        RECT 127.205 116.340 127.495 116.385 ;
        RECT 132.265 116.340 132.555 116.385 ;
        RECT 133.170 116.340 133.490 116.400 ;
        RECT 127.205 116.200 129.720 116.340 ;
        RECT 127.205 116.155 127.495 116.200 ;
        RECT 66.180 115.860 67.620 116.000 ;
        RECT 66.180 115.815 66.470 115.860 ;
        RECT 67.850 115.800 68.170 116.060 ;
        RECT 68.770 116.045 69.090 116.060 ;
        RECT 68.770 115.815 69.155 116.045 ;
        RECT 69.690 116.000 70.010 116.060 ;
        RECT 91.400 116.000 91.540 116.140 ;
        RECT 69.690 115.860 75.900 116.000 ;
        RECT 68.770 115.800 69.090 115.815 ;
        RECT 69.690 115.800 70.010 115.860 ;
        RECT 24.165 115.475 24.455 115.705 ;
        RECT 25.500 115.475 25.850 115.705 ;
        RECT 31.525 115.475 31.815 115.705 ;
        RECT 37.030 115.660 37.350 115.720 ;
        RECT 37.950 115.660 38.270 115.720 ;
        RECT 37.030 115.520 38.270 115.660 ;
        RECT 25.530 115.460 25.850 115.475 ;
        RECT 37.030 115.460 37.350 115.520 ;
        RECT 37.950 115.460 38.270 115.520 ;
        RECT 41.170 115.460 41.490 115.720 ;
        RECT 42.565 115.660 42.855 115.705 ;
        RECT 43.010 115.660 43.330 115.720 ;
        RECT 42.565 115.520 43.330 115.660 ;
        RECT 42.565 115.475 42.855 115.520 ;
        RECT 43.010 115.460 43.330 115.520 ;
        RECT 43.485 115.660 43.775 115.705 ;
        RECT 44.405 115.660 44.695 115.705 ;
        RECT 43.485 115.520 44.695 115.660 ;
        RECT 43.485 115.475 43.775 115.520 ;
        RECT 44.405 115.475 44.695 115.520 ;
        RECT 46.690 115.660 47.010 115.720 ;
        RECT 49.005 115.660 49.295 115.705 ;
        RECT 46.690 115.520 49.295 115.660 ;
        RECT 46.690 115.460 47.010 115.520 ;
        RECT 49.005 115.475 49.295 115.520 ;
        RECT 49.450 115.660 49.770 115.720 ;
        RECT 75.760 115.705 75.900 115.860 ;
        RECT 90.020 115.860 91.540 116.000 ;
        RECT 50.285 115.660 50.575 115.705 ;
        RECT 49.450 115.520 50.575 115.660 ;
        RECT 49.450 115.460 49.770 115.520 ;
        RECT 50.285 115.475 50.575 115.520 ;
        RECT 67.405 115.660 67.695 115.705 ;
        RECT 67.405 115.520 75.440 115.660 ;
        RECT 67.405 115.475 67.695 115.520 ;
        RECT 25.045 115.320 25.335 115.365 ;
        RECT 26.235 115.320 26.525 115.365 ;
        RECT 28.755 115.320 29.045 115.365 ;
        RECT 25.045 115.180 29.045 115.320 ;
        RECT 25.045 115.135 25.335 115.180 ;
        RECT 26.235 115.135 26.525 115.180 ;
        RECT 28.755 115.135 29.045 115.180 ;
        RECT 32.405 115.320 32.695 115.365 ;
        RECT 33.595 115.320 33.885 115.365 ;
        RECT 36.115 115.320 36.405 115.365 ;
        RECT 32.405 115.180 36.405 115.320 ;
        RECT 32.405 115.135 32.695 115.180 ;
        RECT 33.595 115.135 33.885 115.180 ;
        RECT 36.115 115.135 36.405 115.180 ;
        RECT 43.930 115.320 44.250 115.380 ;
        RECT 47.165 115.320 47.455 115.365 ;
        RECT 43.930 115.180 47.455 115.320 ;
        RECT 43.930 115.120 44.250 115.180 ;
        RECT 47.165 115.135 47.455 115.180 ;
        RECT 49.885 115.320 50.175 115.365 ;
        RECT 51.075 115.320 51.365 115.365 ;
        RECT 53.595 115.320 53.885 115.365 ;
        RECT 49.885 115.180 53.885 115.320 ;
        RECT 49.885 115.135 50.175 115.180 ;
        RECT 51.075 115.135 51.365 115.180 ;
        RECT 53.595 115.135 53.885 115.180 ;
        RECT 59.125 115.135 59.415 115.365 ;
        RECT 62.815 115.320 63.105 115.365 ;
        RECT 65.335 115.320 65.625 115.365 ;
        RECT 66.525 115.320 66.815 115.365 ;
        RECT 62.815 115.180 66.815 115.320 ;
        RECT 62.815 115.135 63.105 115.180 ;
        RECT 65.335 115.135 65.625 115.180 ;
        RECT 66.525 115.135 66.815 115.180 ;
        RECT 67.850 115.320 68.170 115.380 ;
        RECT 72.925 115.320 73.215 115.365 ;
        RECT 67.850 115.180 73.215 115.320 ;
        RECT 75.300 115.320 75.440 115.520 ;
        RECT 75.685 115.475 75.975 115.705 ;
        RECT 76.590 115.460 76.910 115.720 ;
        RECT 77.050 115.460 77.370 115.720 ;
        RECT 78.430 115.460 78.750 115.720 ;
        RECT 79.825 115.660 80.115 115.705 ;
        RECT 80.730 115.660 81.050 115.720 ;
        RECT 79.825 115.520 81.050 115.660 ;
        RECT 79.825 115.475 80.115 115.520 ;
        RECT 80.730 115.460 81.050 115.520 ;
        RECT 81.620 115.660 81.910 115.705 ;
        RECT 83.490 115.660 83.810 115.720 ;
        RECT 90.020 115.705 90.160 115.860 ;
        RECT 94.070 115.800 94.390 116.060 ;
        RECT 114.325 116.000 114.615 116.045 ;
        RECT 118.450 116.000 118.770 116.060 ;
        RECT 97.380 115.860 118.770 116.000 ;
        RECT 81.620 115.520 83.810 115.660 ;
        RECT 81.620 115.475 81.910 115.520 ;
        RECT 83.490 115.460 83.810 115.520 ;
        RECT 89.945 115.475 90.235 115.705 ;
        RECT 90.865 115.475 91.155 115.705 ;
        RECT 91.310 115.660 91.630 115.720 ;
        RECT 92.230 115.660 92.550 115.720 ;
        RECT 91.310 115.520 92.550 115.660 ;
        RECT 79.350 115.320 79.670 115.380 ;
        RECT 75.300 115.280 80.040 115.320 ;
        RECT 80.285 115.280 80.575 115.365 ;
        RECT 75.300 115.180 80.575 115.280 ;
        RECT 24.650 114.980 24.940 115.025 ;
        RECT 26.750 114.980 27.040 115.025 ;
        RECT 28.320 114.980 28.610 115.025 ;
        RECT 24.650 114.840 28.610 114.980 ;
        RECT 24.650 114.795 24.940 114.840 ;
        RECT 26.750 114.795 27.040 114.840 ;
        RECT 28.320 114.795 28.610 114.840 ;
        RECT 32.010 114.980 32.300 115.025 ;
        RECT 34.110 114.980 34.400 115.025 ;
        RECT 35.680 114.980 35.970 115.025 ;
        RECT 32.010 114.840 35.970 114.980 ;
        RECT 32.010 114.795 32.300 114.840 ;
        RECT 34.110 114.795 34.400 114.840 ;
        RECT 35.680 114.795 35.970 114.840 ;
        RECT 49.490 114.980 49.780 115.025 ;
        RECT 51.590 114.980 51.880 115.025 ;
        RECT 53.160 114.980 53.450 115.025 ;
        RECT 49.490 114.840 53.450 114.980 ;
        RECT 49.490 114.795 49.780 114.840 ;
        RECT 51.590 114.795 51.880 114.840 ;
        RECT 53.160 114.795 53.450 114.840 ;
        RECT 54.970 114.980 55.290 115.040 ;
        RECT 56.365 114.980 56.655 115.025 ;
        RECT 54.970 114.840 56.655 114.980 ;
        RECT 54.970 114.780 55.290 114.840 ;
        RECT 56.365 114.795 56.655 114.840 ;
        RECT 31.050 114.440 31.370 114.700 ;
        RECT 40.265 114.640 40.555 114.685 ;
        RECT 40.710 114.640 41.030 114.700 ;
        RECT 40.265 114.500 41.030 114.640 ;
        RECT 40.265 114.455 40.555 114.500 ;
        RECT 40.710 114.440 41.030 114.500 ;
        RECT 55.905 114.640 56.195 114.685 ;
        RECT 57.730 114.640 58.050 114.700 ;
        RECT 59.200 114.640 59.340 115.135 ;
        RECT 67.850 115.120 68.170 115.180 ;
        RECT 72.925 115.135 73.215 115.180 ;
        RECT 79.350 115.120 79.670 115.180 ;
        RECT 79.900 115.140 80.575 115.180 ;
        RECT 80.285 115.135 80.575 115.140 ;
        RECT 81.165 115.320 81.455 115.365 ;
        RECT 82.355 115.320 82.645 115.365 ;
        RECT 84.875 115.320 85.165 115.365 ;
        RECT 90.940 115.320 91.080 115.475 ;
        RECT 91.310 115.460 91.630 115.520 ;
        RECT 92.230 115.460 92.550 115.520 ;
        RECT 97.380 115.320 97.520 115.860 ;
        RECT 114.325 115.815 114.615 115.860 ;
        RECT 118.450 115.800 118.770 115.860 ;
        RECT 99.605 115.660 99.895 115.705 ;
        RECT 100.970 115.660 101.290 115.720 ;
        RECT 99.605 115.520 101.290 115.660 ;
        RECT 99.605 115.475 99.895 115.520 ;
        RECT 100.970 115.460 101.290 115.520 ;
        RECT 112.470 115.660 112.790 115.720 ;
        RECT 113.865 115.660 114.155 115.705 ;
        RECT 112.470 115.520 114.155 115.660 ;
        RECT 112.470 115.460 112.790 115.520 ;
        RECT 113.865 115.475 114.155 115.520 ;
        RECT 114.770 115.660 115.090 115.720 ;
        RECT 115.245 115.660 115.535 115.705 ;
        RECT 114.770 115.520 115.535 115.660 ;
        RECT 114.770 115.460 115.090 115.520 ;
        RECT 115.245 115.475 115.535 115.520 ;
        RECT 128.110 115.650 128.430 115.720 ;
        RECT 129.580 115.705 129.720 116.200 ;
        RECT 132.265 116.200 133.490 116.340 ;
        RECT 132.265 116.155 132.555 116.200 ;
        RECT 133.170 116.140 133.490 116.200 ;
        RECT 135.560 116.200 136.620 116.340 ;
        RECT 135.560 116.000 135.700 116.200 ;
        RECT 130.040 115.860 135.700 116.000 ;
        RECT 129.045 115.650 129.335 115.705 ;
        RECT 128.110 115.510 129.335 115.650 ;
        RECT 128.110 115.460 128.430 115.510 ;
        RECT 129.045 115.475 129.335 115.510 ;
        RECT 129.505 115.475 129.795 115.705 ;
        RECT 81.165 115.180 85.165 115.320 ;
        RECT 81.165 115.135 81.455 115.180 ;
        RECT 82.355 115.135 82.645 115.180 ;
        RECT 84.875 115.135 85.165 115.180 ;
        RECT 86.800 115.180 97.520 115.320 ;
        RECT 97.750 115.320 98.070 115.380 ;
        RECT 98.225 115.320 98.515 115.365 ;
        RECT 97.750 115.180 98.515 115.320 ;
        RECT 63.250 114.980 63.540 115.025 ;
        RECT 64.820 114.980 65.110 115.025 ;
        RECT 66.920 114.980 67.210 115.025 ;
        RECT 70.165 114.980 70.455 115.025 ;
        RECT 63.250 114.840 67.210 114.980 ;
        RECT 63.250 114.795 63.540 114.840 ;
        RECT 64.820 114.795 65.110 114.840 ;
        RECT 66.920 114.795 67.210 114.840 ;
        RECT 68.860 114.840 70.455 114.980 ;
        RECT 55.905 114.500 59.340 114.640 ;
        RECT 60.505 114.640 60.795 114.685 ;
        RECT 65.550 114.640 65.870 114.700 ;
        RECT 68.860 114.685 69.000 114.840 ;
        RECT 70.165 114.795 70.455 114.840 ;
        RECT 80.770 114.980 81.060 115.025 ;
        RECT 82.870 114.980 83.160 115.025 ;
        RECT 84.440 114.980 84.730 115.025 ;
        RECT 80.770 114.840 84.730 114.980 ;
        RECT 80.770 114.795 81.060 114.840 ;
        RECT 82.870 114.795 83.160 114.840 ;
        RECT 84.440 114.795 84.730 114.840 ;
        RECT 60.505 114.500 65.870 114.640 ;
        RECT 55.905 114.455 56.195 114.500 ;
        RECT 57.730 114.440 58.050 114.500 ;
        RECT 60.505 114.455 60.795 114.500 ;
        RECT 65.550 114.440 65.870 114.500 ;
        RECT 68.785 114.455 69.075 114.685 ;
        RECT 69.705 114.640 69.995 114.685 ;
        RECT 71.070 114.640 71.390 114.700 ;
        RECT 69.705 114.500 71.390 114.640 ;
        RECT 69.705 114.455 69.995 114.500 ;
        RECT 71.070 114.440 71.390 114.500 ;
        RECT 71.530 114.640 71.850 114.700 ;
        RECT 81.190 114.640 81.510 114.700 ;
        RECT 86.800 114.640 86.940 115.180 ;
        RECT 97.750 115.120 98.070 115.180 ;
        RECT 98.225 115.135 98.515 115.180 ;
        RECT 99.145 115.320 99.435 115.365 ;
        RECT 100.050 115.320 100.370 115.380 ;
        RECT 99.145 115.180 100.370 115.320 ;
        RECT 99.145 115.135 99.435 115.180 ;
        RECT 100.050 115.120 100.370 115.180 ;
        RECT 109.250 115.320 109.570 115.380 ;
        RECT 110.185 115.320 110.475 115.365 ;
        RECT 109.250 115.180 110.475 115.320 ;
        RECT 109.250 115.120 109.570 115.180 ;
        RECT 110.185 115.135 110.475 115.180 ;
        RECT 118.450 115.320 118.770 115.380 ;
        RECT 120.290 115.320 120.610 115.380 ;
        RECT 121.225 115.320 121.515 115.365 ;
        RECT 118.450 115.180 121.515 115.320 ;
        RECT 118.450 115.120 118.770 115.180 ;
        RECT 120.290 115.120 120.610 115.180 ;
        RECT 121.225 115.135 121.515 115.180 ;
        RECT 128.585 115.320 128.875 115.365 ;
        RECT 130.040 115.320 130.180 115.860 ;
        RECT 135.930 115.800 136.250 116.060 ;
        RECT 136.480 116.000 136.620 116.200 ;
        RECT 136.850 116.140 137.170 116.400 ;
        RECT 137.310 116.340 137.630 116.400 ;
        RECT 139.165 116.340 139.455 116.385 ;
        RECT 145.130 116.340 145.450 116.400 ;
        RECT 137.310 116.200 139.455 116.340 ;
        RECT 137.310 116.140 137.630 116.200 ;
        RECT 139.165 116.155 139.455 116.200 ;
        RECT 139.700 116.200 145.450 116.340 ;
        RECT 139.700 116.000 139.840 116.200 ;
        RECT 145.130 116.140 145.450 116.200 ;
        RECT 146.050 116.140 146.370 116.400 ;
        RECT 152.030 116.140 152.350 116.400 ;
        RECT 136.480 115.860 139.840 116.000 ;
        RECT 140.085 116.000 140.375 116.045 ;
        RECT 141.450 116.000 141.770 116.060 ;
        RECT 140.085 115.860 141.770 116.000 ;
        RECT 140.085 115.815 140.375 115.860 ;
        RECT 141.450 115.800 141.770 115.860 ;
        RECT 146.970 116.000 147.290 116.060 ;
        RECT 154.790 116.000 155.110 116.060 ;
        RECT 146.970 115.860 149.040 116.000 ;
        RECT 146.970 115.800 147.290 115.860 ;
        RECT 132.250 115.660 132.570 115.720 ;
        RECT 133.645 115.660 133.935 115.705 ;
        RECT 132.250 115.520 133.935 115.660 ;
        RECT 132.250 115.460 132.570 115.520 ;
        RECT 133.645 115.475 133.935 115.520 ;
        RECT 134.565 115.660 134.855 115.705 ;
        RECT 135.025 115.660 135.315 115.705 ;
        RECT 137.785 115.660 138.075 115.705 ;
        RECT 141.005 115.660 141.295 115.705 ;
        RECT 141.910 115.660 142.230 115.720 ;
        RECT 134.565 115.520 142.230 115.660 ;
        RECT 134.565 115.475 134.855 115.520 ;
        RECT 135.025 115.475 135.315 115.520 ;
        RECT 137.785 115.475 138.075 115.520 ;
        RECT 141.005 115.475 141.295 115.520 ;
        RECT 141.910 115.460 142.230 115.520 ;
        RECT 147.905 115.475 148.195 115.705 ;
        RECT 128.585 115.180 130.180 115.320 ;
        RECT 130.410 115.320 130.730 115.380 ;
        RECT 130.885 115.320 131.175 115.365 ;
        RECT 130.410 115.180 131.175 115.320 ;
        RECT 128.585 115.135 128.875 115.180 ;
        RECT 130.410 115.120 130.730 115.180 ;
        RECT 130.885 115.135 131.175 115.180 ;
        RECT 143.305 115.320 143.595 115.365 ;
        RECT 146.525 115.320 146.815 115.365 ;
        RECT 143.305 115.180 146.815 115.320 ;
        RECT 147.980 115.320 148.120 115.475 ;
        RECT 148.350 115.460 148.670 115.720 ;
        RECT 148.900 115.705 149.040 115.860 ;
        RECT 150.280 115.860 155.110 116.000 ;
        RECT 150.280 115.720 150.420 115.860 ;
        RECT 154.790 115.800 155.110 115.860 ;
        RECT 148.825 115.475 149.115 115.705 ;
        RECT 149.745 115.660 150.035 115.705 ;
        RECT 150.190 115.660 150.510 115.720 ;
        RECT 149.745 115.520 150.510 115.660 ;
        RECT 149.745 115.475 150.035 115.520 ;
        RECT 150.190 115.460 150.510 115.520 ;
        RECT 153.410 115.460 153.730 115.720 ;
        RECT 153.885 115.475 154.175 115.705 ;
        RECT 150.650 115.320 150.970 115.380 ;
        RECT 147.980 115.180 150.970 115.320 ;
        RECT 143.305 115.135 143.595 115.180 ;
        RECT 146.525 115.135 146.815 115.180 ;
        RECT 150.650 115.120 150.970 115.180 ;
        RECT 88.090 114.980 88.410 115.040 ;
        RECT 93.165 114.980 93.455 115.025 ;
        RECT 142.830 114.980 143.150 115.040 ;
        RECT 88.090 114.840 93.455 114.980 ;
        RECT 88.090 114.780 88.410 114.840 ;
        RECT 93.165 114.795 93.455 114.840 ;
        RECT 129.120 114.840 143.150 114.980 ;
        RECT 71.530 114.500 86.940 114.640 ;
        RECT 110.630 114.640 110.950 114.700 ;
        RECT 113.405 114.640 113.695 114.685 ;
        RECT 110.630 114.500 113.695 114.640 ;
        RECT 71.530 114.440 71.850 114.500 ;
        RECT 81.190 114.440 81.510 114.500 ;
        RECT 110.630 114.440 110.950 114.500 ;
        RECT 113.405 114.455 113.695 114.500 ;
        RECT 115.690 114.640 116.010 114.700 ;
        RECT 129.120 114.685 129.260 114.840 ;
        RECT 142.830 114.780 143.150 114.840 ;
        RECT 148.350 114.980 148.670 115.040 ;
        RECT 153.960 114.980 154.100 115.475 ;
        RECT 154.330 115.460 154.650 115.720 ;
        RECT 154.880 115.660 155.020 115.800 ;
        RECT 155.265 115.660 155.555 115.705 ;
        RECT 154.880 115.520 155.555 115.660 ;
        RECT 155.265 115.475 155.555 115.520 ;
        RECT 148.350 114.840 154.100 114.980 ;
        RECT 148.350 114.780 148.670 114.840 ;
        RECT 118.465 114.640 118.755 114.685 ;
        RECT 115.690 114.500 118.755 114.640 ;
        RECT 115.690 114.440 116.010 114.500 ;
        RECT 118.465 114.455 118.755 114.500 ;
        RECT 129.045 114.455 129.335 114.685 ;
        RECT 131.345 114.640 131.635 114.685 ;
        RECT 132.710 114.640 133.030 114.700 ;
        RECT 131.345 114.500 133.030 114.640 ;
        RECT 131.345 114.455 131.635 114.500 ;
        RECT 132.710 114.440 133.030 114.500 ;
        RECT 135.930 114.640 136.250 114.700 ;
        RECT 138.245 114.640 138.535 114.685 ;
        RECT 135.930 114.500 138.535 114.640 ;
        RECT 135.930 114.440 136.250 114.500 ;
        RECT 138.245 114.455 138.535 114.500 ;
        RECT 22.700 113.820 157.020 114.300 ;
        RECT 25.530 113.620 25.850 113.680 ;
        RECT 26.465 113.620 26.755 113.665 ;
        RECT 25.530 113.480 26.755 113.620 ;
        RECT 25.530 113.420 25.850 113.480 ;
        RECT 26.465 113.435 26.755 113.480 ;
        RECT 37.045 113.620 37.335 113.665 ;
        RECT 37.950 113.620 38.270 113.680 ;
        RECT 41.630 113.620 41.950 113.680 ;
        RECT 37.045 113.480 38.270 113.620 ;
        RECT 37.045 113.435 37.335 113.480 ;
        RECT 37.950 113.420 38.270 113.480 ;
        RECT 38.500 113.480 41.950 113.620 ;
        RECT 36.125 113.280 36.415 113.325 ;
        RECT 38.500 113.280 38.640 113.480 ;
        RECT 41.630 113.420 41.950 113.480 ;
        RECT 43.930 113.620 44.250 113.680 ;
        RECT 45.325 113.620 45.615 113.665 ;
        RECT 43.930 113.480 45.615 113.620 ;
        RECT 43.930 113.420 44.250 113.480 ;
        RECT 45.325 113.435 45.615 113.480 ;
        RECT 48.085 113.620 48.375 113.665 ;
        RECT 49.450 113.620 49.770 113.680 ;
        RECT 48.085 113.480 49.770 113.620 ;
        RECT 48.085 113.435 48.375 113.480 ;
        RECT 49.450 113.420 49.770 113.480 ;
        RECT 54.510 113.620 54.830 113.680 ;
        RECT 55.905 113.620 56.195 113.665 ;
        RECT 54.510 113.480 56.195 113.620 ;
        RECT 54.510 113.420 54.830 113.480 ;
        RECT 55.905 113.435 56.195 113.480 ;
        RECT 36.125 113.140 38.640 113.280 ;
        RECT 38.910 113.280 39.200 113.325 ;
        RECT 41.010 113.280 41.300 113.325 ;
        RECT 42.580 113.280 42.870 113.325 ;
        RECT 38.910 113.140 42.870 113.280 ;
        RECT 36.125 113.095 36.415 113.140 ;
        RECT 38.910 113.095 39.200 113.140 ;
        RECT 41.010 113.095 41.300 113.140 ;
        RECT 42.580 113.095 42.870 113.140 ;
        RECT 31.050 112.940 31.370 113.000 ;
        RECT 32.905 112.940 33.195 112.985 ;
        RECT 39.305 112.940 39.595 112.985 ;
        RECT 40.495 112.940 40.785 112.985 ;
        RECT 43.015 112.940 43.305 112.985 ;
        RECT 31.050 112.800 33.810 112.940 ;
        RECT 31.050 112.740 31.370 112.800 ;
        RECT 32.905 112.755 33.195 112.800 ;
        RECT 26.910 112.600 27.230 112.660 ;
        RECT 29.225 112.600 29.515 112.645 ;
        RECT 26.910 112.460 29.515 112.600 ;
        RECT 33.670 112.600 33.810 112.800 ;
        RECT 39.305 112.800 43.305 112.940 ;
        RECT 39.305 112.755 39.595 112.800 ;
        RECT 40.495 112.755 40.785 112.800 ;
        RECT 43.015 112.755 43.305 112.800 ;
        RECT 53.130 112.940 53.450 113.000 ;
        RECT 55.980 112.940 56.120 113.435 ;
        RECT 57.270 113.420 57.590 113.680 ;
        RECT 64.205 113.620 64.495 113.665 ;
        RECT 65.125 113.620 65.415 113.665 ;
        RECT 64.205 113.480 65.415 113.620 ;
        RECT 64.205 113.435 64.495 113.480 ;
        RECT 65.125 113.435 65.415 113.480 ;
        RECT 67.850 113.420 68.170 113.680 ;
        RECT 80.745 113.620 81.035 113.665 ;
        RECT 83.490 113.620 83.810 113.680 ;
        RECT 80.745 113.480 83.810 113.620 ;
        RECT 80.745 113.435 81.035 113.480 ;
        RECT 83.490 113.420 83.810 113.480 ;
        RECT 84.425 113.620 84.715 113.665 ;
        RECT 86.250 113.620 86.570 113.680 ;
        RECT 87.170 113.620 87.490 113.680 ;
        RECT 84.425 113.480 87.490 113.620 ;
        RECT 84.425 113.435 84.715 113.480 ;
        RECT 86.250 113.420 86.570 113.480 ;
        RECT 87.170 113.420 87.490 113.480 ;
        RECT 92.245 113.620 92.535 113.665 ;
        RECT 98.210 113.620 98.530 113.680 ;
        RECT 100.525 113.620 100.815 113.665 ;
        RECT 100.970 113.620 101.290 113.680 ;
        RECT 92.245 113.480 101.290 113.620 ;
        RECT 92.245 113.435 92.535 113.480 ;
        RECT 98.210 113.420 98.530 113.480 ;
        RECT 100.525 113.435 100.815 113.480 ;
        RECT 100.970 113.420 101.290 113.480 ;
        RECT 109.250 113.420 109.570 113.680 ;
        RECT 110.630 113.420 110.950 113.680 ;
        RECT 114.770 113.420 115.090 113.680 ;
        RECT 115.690 113.420 116.010 113.680 ;
        RECT 129.030 113.420 129.350 113.680 ;
        RECT 131.345 113.620 131.635 113.665 ;
        RECT 143.750 113.620 144.070 113.680 ;
        RECT 148.350 113.620 148.670 113.680 ;
        RECT 131.345 113.480 144.070 113.620 ;
        RECT 131.345 113.435 131.635 113.480 ;
        RECT 143.750 113.420 144.070 113.480 ;
        RECT 144.300 113.480 148.670 113.620 ;
        RECT 70.610 113.280 70.900 113.325 ;
        RECT 72.180 113.280 72.470 113.325 ;
        RECT 74.280 113.280 74.570 113.325 ;
        RECT 70.610 113.140 74.570 113.280 ;
        RECT 70.610 113.095 70.900 113.140 ;
        RECT 72.180 113.095 72.470 113.140 ;
        RECT 74.280 113.095 74.570 113.140 ;
        RECT 94.110 113.280 94.400 113.325 ;
        RECT 96.210 113.280 96.500 113.325 ;
        RECT 97.780 113.280 98.070 113.325 ;
        RECT 94.110 113.140 98.070 113.280 ;
        RECT 94.110 113.095 94.400 113.140 ;
        RECT 96.210 113.095 96.500 113.140 ;
        RECT 97.780 113.095 98.070 113.140 ;
        RECT 102.850 113.280 103.140 113.325 ;
        RECT 104.950 113.280 105.240 113.325 ;
        RECT 106.520 113.280 106.810 113.325 ;
        RECT 102.850 113.140 106.810 113.280 ;
        RECT 102.850 113.095 103.140 113.140 ;
        RECT 104.950 113.095 105.240 113.140 ;
        RECT 106.520 113.095 106.810 113.140 ;
        RECT 124.445 113.280 124.735 113.325 ;
        RECT 124.890 113.280 125.210 113.340 ;
        RECT 135.470 113.280 135.790 113.340 ;
        RECT 124.445 113.140 135.790 113.280 ;
        RECT 124.445 113.095 124.735 113.140 ;
        RECT 124.890 113.080 125.210 113.140 ;
        RECT 135.470 113.080 135.790 113.140 ;
        RECT 70.175 112.940 70.465 112.985 ;
        RECT 72.695 112.940 72.985 112.985 ;
        RECT 73.885 112.940 74.175 112.985 ;
        RECT 53.130 112.800 54.740 112.940 ;
        RECT 55.980 112.800 63.480 112.940 ;
        RECT 53.130 112.740 53.450 112.800 ;
        RECT 37.030 112.600 37.350 112.660 ;
        RECT 33.670 112.460 37.350 112.600 ;
        RECT 26.910 112.400 27.230 112.460 ;
        RECT 29.225 112.415 29.515 112.460 ;
        RECT 37.030 112.400 37.350 112.460 ;
        RECT 38.425 112.600 38.715 112.645 ;
        RECT 46.690 112.600 47.010 112.660 ;
        RECT 38.425 112.460 47.010 112.600 ;
        RECT 38.425 112.415 38.715 112.460 ;
        RECT 46.690 112.400 47.010 112.460 ;
        RECT 47.165 112.415 47.455 112.645 ;
        RECT 48.085 112.600 48.375 112.645 ;
        RECT 51.305 112.600 51.595 112.645 ;
        RECT 48.085 112.460 51.595 112.600 ;
        RECT 48.085 112.415 48.375 112.460 ;
        RECT 51.305 112.415 51.595 112.460 ;
        RECT 53.590 112.600 53.910 112.660 ;
        RECT 54.065 112.600 54.355 112.645 ;
        RECT 53.590 112.460 54.355 112.600 ;
        RECT 54.600 112.600 54.740 112.800 ;
        RECT 57.285 112.600 57.575 112.645 ;
        RECT 54.600 112.460 57.575 112.600 ;
        RECT 37.120 112.260 37.260 112.400 ;
        RECT 37.965 112.260 38.255 112.305 ;
        RECT 37.120 112.120 38.255 112.260 ;
        RECT 37.965 112.075 38.255 112.120 ;
        RECT 39.760 112.260 40.050 112.305 ;
        RECT 40.250 112.260 40.570 112.320 ;
        RECT 39.760 112.120 40.570 112.260 ;
        RECT 39.760 112.075 40.050 112.120 ;
        RECT 40.250 112.060 40.570 112.120 ;
        RECT 29.210 111.920 29.530 111.980 ;
        RECT 37.030 111.965 37.350 111.980 ;
        RECT 30.145 111.920 30.435 111.965 ;
        RECT 29.210 111.780 30.435 111.920 ;
        RECT 29.210 111.720 29.530 111.780 ;
        RECT 30.145 111.735 30.435 111.780 ;
        RECT 36.965 111.735 37.350 111.965 ;
        RECT 47.240 111.920 47.380 112.415 ;
        RECT 53.590 112.400 53.910 112.460 ;
        RECT 54.065 112.415 54.355 112.460 ;
        RECT 57.285 112.415 57.575 112.460 ;
        RECT 57.730 112.400 58.050 112.660 ;
        RECT 58.740 112.645 58.880 112.800 ;
        RECT 58.665 112.415 58.955 112.645 ;
        RECT 60.950 112.600 61.270 112.660 ;
        RECT 63.340 112.645 63.480 112.800 ;
        RECT 70.175 112.800 74.175 112.940 ;
        RECT 70.175 112.755 70.465 112.800 ;
        RECT 72.695 112.755 72.985 112.800 ;
        RECT 73.885 112.755 74.175 112.800 ;
        RECT 74.765 112.940 75.055 112.985 ;
        RECT 79.350 112.940 79.670 113.000 ;
        RECT 74.765 112.800 79.670 112.940 ;
        RECT 74.765 112.755 75.055 112.800 ;
        RECT 79.350 112.740 79.670 112.800 ;
        RECT 93.625 112.755 93.915 112.985 ;
        RECT 94.505 112.940 94.795 112.985 ;
        RECT 95.695 112.940 95.985 112.985 ;
        RECT 98.215 112.940 98.505 112.985 ;
        RECT 94.505 112.800 98.505 112.940 ;
        RECT 94.505 112.755 94.795 112.800 ;
        RECT 95.695 112.755 95.985 112.800 ;
        RECT 98.215 112.755 98.505 112.800 ;
        RECT 101.890 112.940 102.210 113.000 ;
        RECT 102.365 112.940 102.655 112.985 ;
        RECT 101.890 112.800 102.655 112.940 ;
        RECT 62.345 112.600 62.635 112.645 ;
        RECT 60.950 112.460 62.635 112.600 ;
        RECT 60.950 112.400 61.270 112.460 ;
        RECT 62.345 112.415 62.635 112.460 ;
        RECT 63.265 112.415 63.555 112.645 ;
        RECT 81.665 112.415 81.955 112.645 ;
        RECT 82.570 112.600 82.890 112.660 ;
        RECT 83.045 112.600 83.335 112.645 ;
        RECT 82.570 112.460 83.335 112.600 ;
        RECT 52.670 112.260 52.990 112.320 ;
        RECT 55.745 112.260 56.035 112.305 ;
        RECT 52.670 112.120 56.035 112.260 ;
        RECT 52.670 112.060 52.990 112.120 ;
        RECT 55.745 112.075 56.035 112.120 ;
        RECT 56.825 112.260 57.115 112.305 ;
        RECT 57.820 112.260 57.960 112.400 ;
        RECT 56.825 112.120 57.960 112.260 ;
        RECT 71.990 112.260 72.310 112.320 ;
        RECT 73.430 112.260 73.720 112.305 ;
        RECT 71.990 112.120 73.720 112.260 ;
        RECT 81.740 112.260 81.880 112.415 ;
        RECT 82.570 112.400 82.890 112.460 ;
        RECT 83.045 112.415 83.335 112.460 ;
        RECT 92.690 112.400 93.010 112.660 ;
        RECT 93.700 112.600 93.840 112.755 ;
        RECT 101.890 112.740 102.210 112.800 ;
        RECT 102.365 112.755 102.655 112.800 ;
        RECT 103.245 112.940 103.535 112.985 ;
        RECT 104.435 112.940 104.725 112.985 ;
        RECT 106.955 112.940 107.245 112.985 ;
        RECT 103.245 112.800 107.245 112.940 ;
        RECT 103.245 112.755 103.535 112.800 ;
        RECT 104.435 112.755 104.725 112.800 ;
        RECT 106.955 112.755 107.245 112.800 ;
        RECT 123.525 112.940 123.815 112.985 ;
        RECT 125.350 112.940 125.670 113.000 ;
        RECT 130.410 112.940 130.730 113.000 ;
        RECT 123.525 112.800 125.670 112.940 ;
        RECT 123.525 112.755 123.815 112.800 ;
        RECT 125.350 112.740 125.670 112.800 ;
        RECT 128.660 112.800 130.730 112.940 ;
        RECT 101.980 112.600 102.120 112.740 ;
        RECT 128.660 112.660 128.800 112.800 ;
        RECT 130.410 112.740 130.730 112.800 ;
        RECT 132.340 112.800 143.060 112.940 ;
        RECT 93.700 112.460 102.120 112.600 ;
        RECT 115.230 112.400 115.550 112.660 ;
        RECT 118.450 112.400 118.770 112.660 ;
        RECT 119.830 112.400 120.150 112.660 ;
        RECT 124.905 112.600 125.195 112.645 ;
        RECT 123.140 112.460 125.195 112.600 ;
        RECT 84.410 112.305 84.730 112.320 ;
        RECT 81.740 112.120 83.720 112.260 ;
        RECT 56.825 112.075 57.115 112.120 ;
        RECT 71.990 112.060 72.310 112.120 ;
        RECT 73.430 112.075 73.720 112.120 ;
        RECT 54.510 111.920 54.830 111.980 ;
        RECT 54.985 111.920 55.275 111.965 ;
        RECT 47.240 111.780 55.275 111.920 ;
        RECT 37.030 111.720 37.350 111.735 ;
        RECT 54.510 111.720 54.830 111.780 ;
        RECT 54.985 111.735 55.275 111.780 ;
        RECT 66.930 111.920 67.250 111.980 ;
        RECT 67.405 111.920 67.695 111.965 ;
        RECT 66.930 111.780 67.695 111.920 ;
        RECT 66.930 111.720 67.250 111.780 ;
        RECT 67.405 111.735 67.695 111.780 ;
        RECT 76.590 111.920 76.910 111.980 ;
        RECT 82.570 111.920 82.890 111.980 ;
        RECT 83.580 111.965 83.720 112.120 ;
        RECT 84.345 112.075 84.730 112.305 ;
        RECT 84.410 112.060 84.730 112.075 ;
        RECT 84.870 112.260 85.190 112.320 ;
        RECT 85.345 112.260 85.635 112.305 ;
        RECT 88.090 112.260 88.410 112.320 ;
        RECT 84.870 112.120 88.410 112.260 ;
        RECT 84.870 112.060 85.190 112.120 ;
        RECT 85.345 112.075 85.635 112.120 ;
        RECT 88.090 112.060 88.410 112.120 ;
        RECT 91.325 112.260 91.615 112.305 ;
        RECT 92.780 112.260 92.920 112.400 ;
        RECT 93.610 112.260 93.930 112.320 ;
        RECT 91.325 112.120 93.930 112.260 ;
        RECT 91.325 112.075 91.615 112.120 ;
        RECT 93.610 112.060 93.930 112.120 ;
        RECT 94.960 112.260 95.250 112.305 ;
        RECT 96.830 112.260 97.150 112.320 ;
        RECT 94.960 112.120 97.150 112.260 ;
        RECT 94.960 112.075 95.250 112.120 ;
        RECT 96.830 112.060 97.150 112.120 ;
        RECT 103.700 112.260 103.990 112.305 ;
        RECT 104.650 112.260 104.970 112.320 ;
        RECT 103.700 112.120 104.970 112.260 ;
        RECT 103.700 112.075 103.990 112.120 ;
        RECT 104.650 112.060 104.970 112.120 ;
        RECT 111.550 112.260 111.870 112.320 ;
        RECT 115.320 112.260 115.460 112.400 ;
        RECT 116.625 112.260 116.915 112.305 ;
        RECT 111.550 112.120 116.915 112.260 ;
        RECT 111.550 112.060 111.870 112.120 ;
        RECT 116.625 112.075 116.915 112.120 ;
        RECT 76.590 111.780 82.890 111.920 ;
        RECT 76.590 111.720 76.910 111.780 ;
        RECT 82.570 111.720 82.890 111.780 ;
        RECT 83.505 111.735 83.795 111.965 ;
        RECT 91.770 111.920 92.090 111.980 ;
        RECT 92.325 111.920 92.615 111.965 ;
        RECT 91.770 111.780 92.615 111.920 ;
        RECT 91.770 111.720 92.090 111.780 ;
        RECT 92.325 111.735 92.615 111.780 ;
        RECT 93.165 111.920 93.455 111.965 ;
        RECT 97.750 111.920 98.070 111.980 ;
        RECT 93.165 111.780 98.070 111.920 ;
        RECT 93.165 111.735 93.455 111.780 ;
        RECT 97.750 111.720 98.070 111.780 ;
        RECT 105.570 111.920 105.890 111.980 ;
        RECT 109.725 111.920 110.015 111.965 ;
        RECT 105.570 111.780 110.015 111.920 ;
        RECT 105.570 111.720 105.890 111.780 ;
        RECT 109.725 111.735 110.015 111.780 ;
        RECT 110.565 111.920 110.855 111.965 ;
        RECT 114.310 111.920 114.630 111.980 ;
        RECT 115.575 111.920 115.865 111.965 ;
        RECT 110.565 111.780 115.865 111.920 ;
        RECT 110.565 111.735 110.855 111.780 ;
        RECT 114.310 111.720 114.630 111.780 ;
        RECT 115.575 111.735 115.865 111.780 ;
        RECT 117.990 111.720 118.310 111.980 ;
        RECT 121.670 111.920 121.990 111.980 ;
        RECT 123.140 111.965 123.280 112.460 ;
        RECT 124.905 112.415 125.195 112.460 ;
        RECT 128.570 112.400 128.890 112.660 ;
        RECT 129.045 112.600 129.335 112.645 ;
        RECT 129.045 112.585 130.640 112.600 ;
        RECT 131.330 112.585 131.650 112.660 ;
        RECT 129.045 112.460 131.650 112.585 ;
        RECT 129.045 112.415 129.335 112.460 ;
        RECT 130.500 112.445 131.650 112.460 ;
        RECT 131.330 112.400 131.650 112.445 ;
        RECT 131.790 112.400 132.110 112.660 ;
        RECT 127.665 112.260 127.955 112.305 ;
        RECT 129.505 112.260 129.795 112.305 ;
        RECT 129.950 112.260 130.270 112.320 ;
        RECT 127.665 112.120 128.800 112.260 ;
        RECT 127.665 112.075 127.955 112.120 ;
        RECT 123.065 111.920 123.355 111.965 ;
        RECT 121.670 111.780 123.355 111.920 ;
        RECT 121.670 111.720 121.990 111.780 ;
        RECT 123.065 111.735 123.355 111.780 ;
        RECT 123.525 111.920 123.815 111.965 ;
        RECT 124.430 111.920 124.750 111.980 ;
        RECT 123.525 111.780 124.750 111.920 ;
        RECT 128.660 111.920 128.800 112.120 ;
        RECT 129.505 112.120 130.270 112.260 ;
        RECT 129.505 112.075 129.795 112.120 ;
        RECT 129.950 112.060 130.270 112.120 ;
        RECT 130.425 112.260 130.715 112.305 ;
        RECT 132.340 112.260 132.480 112.800 ;
        RECT 132.710 112.400 133.030 112.660 ;
        RECT 133.185 112.415 133.475 112.645 ;
        RECT 133.645 112.600 133.935 112.645 ;
        RECT 139.165 112.600 139.455 112.645 ;
        RECT 133.645 112.460 139.455 112.600 ;
        RECT 133.645 112.415 133.935 112.460 ;
        RECT 139.165 112.415 139.455 112.460 ;
        RECT 141.925 112.415 142.215 112.645 ;
        RECT 130.425 112.120 132.480 112.260 ;
        RECT 133.260 112.260 133.400 112.415 ;
        RECT 133.260 112.120 135.700 112.260 ;
        RECT 130.425 112.075 130.715 112.120 ;
        RECT 134.090 111.920 134.410 111.980 ;
        RECT 128.660 111.780 134.410 111.920 ;
        RECT 123.525 111.735 123.815 111.780 ;
        RECT 124.430 111.720 124.750 111.780 ;
        RECT 134.090 111.720 134.410 111.780 ;
        RECT 135.010 111.720 135.330 111.980 ;
        RECT 135.560 111.920 135.700 112.120 ;
        RECT 135.930 112.060 136.250 112.320 ;
        RECT 136.865 112.260 137.155 112.305 ;
        RECT 138.230 112.260 138.550 112.320 ;
        RECT 142.000 112.260 142.140 112.415 ;
        RECT 136.865 112.120 142.140 112.260 ;
        RECT 142.920 112.260 143.060 112.800 ;
        RECT 144.300 112.645 144.440 113.480 ;
        RECT 148.350 113.420 148.670 113.480 ;
        RECT 152.950 113.620 153.270 113.680 ;
        RECT 154.790 113.620 155.110 113.680 ;
        RECT 155.265 113.620 155.555 113.665 ;
        RECT 152.950 113.480 155.555 113.620 ;
        RECT 152.950 113.420 153.270 113.480 ;
        RECT 154.790 113.420 155.110 113.480 ;
        RECT 155.265 113.435 155.555 113.480 ;
        RECT 148.850 113.280 149.140 113.325 ;
        RECT 150.950 113.280 151.240 113.325 ;
        RECT 152.520 113.280 152.810 113.325 ;
        RECT 148.850 113.140 152.810 113.280 ;
        RECT 148.850 113.095 149.140 113.140 ;
        RECT 150.950 113.095 151.240 113.140 ;
        RECT 152.520 113.095 152.810 113.140 ;
        RECT 147.890 112.940 148.210 113.000 ;
        RECT 148.365 112.940 148.655 112.985 ;
        RECT 145.220 112.800 146.740 112.940 ;
        RECT 144.225 112.415 144.515 112.645 ;
        RECT 144.670 112.400 144.990 112.660 ;
        RECT 145.220 112.260 145.360 112.800 ;
        RECT 145.590 112.400 145.910 112.660 ;
        RECT 146.600 112.645 146.740 112.800 ;
        RECT 147.890 112.800 148.655 112.940 ;
        RECT 147.890 112.740 148.210 112.800 ;
        RECT 148.365 112.755 148.655 112.800 ;
        RECT 149.245 112.940 149.535 112.985 ;
        RECT 150.435 112.940 150.725 112.985 ;
        RECT 152.955 112.940 153.245 112.985 ;
        RECT 149.245 112.800 153.245 112.940 ;
        RECT 149.245 112.755 149.535 112.800 ;
        RECT 150.435 112.755 150.725 112.800 ;
        RECT 152.955 112.755 153.245 112.800 ;
        RECT 146.065 112.415 146.355 112.645 ;
        RECT 146.525 112.600 146.815 112.645 ;
        RECT 152.030 112.600 152.350 112.660 ;
        RECT 146.525 112.460 152.350 112.600 ;
        RECT 146.525 112.415 146.815 112.460 ;
        RECT 142.920 112.120 145.360 112.260 ;
        RECT 136.865 112.075 137.155 112.120 ;
        RECT 138.230 112.060 138.550 112.120 ;
        RECT 137.310 111.920 137.630 111.980 ;
        RECT 135.560 111.780 137.630 111.920 ;
        RECT 137.310 111.720 137.630 111.780 ;
        RECT 137.785 111.920 138.075 111.965 ;
        RECT 142.370 111.920 142.690 111.980 ;
        RECT 137.785 111.780 142.690 111.920 ;
        RECT 137.785 111.735 138.075 111.780 ;
        RECT 142.370 111.720 142.690 111.780 ;
        RECT 142.830 111.920 143.150 111.980 ;
        RECT 143.305 111.920 143.595 111.965 ;
        RECT 146.140 111.920 146.280 112.415 ;
        RECT 152.030 112.400 152.350 112.460 ;
        RECT 147.905 112.260 148.195 112.305 ;
        RECT 149.590 112.260 149.880 112.305 ;
        RECT 147.905 112.120 149.880 112.260 ;
        RECT 147.905 112.075 148.195 112.120 ;
        RECT 149.590 112.075 149.880 112.120 ;
        RECT 142.830 111.780 146.280 111.920 ;
        RECT 142.830 111.720 143.150 111.780 ;
        RECT 143.305 111.735 143.595 111.780 ;
        RECT 22.700 111.100 157.820 111.580 ;
        RECT 26.910 110.700 27.230 110.960 ;
        RECT 32.905 110.900 33.195 110.945 ;
        RECT 36.110 110.900 36.430 110.960 ;
        RECT 32.905 110.760 36.430 110.900 ;
        RECT 32.905 110.715 33.195 110.760 ;
        RECT 36.110 110.700 36.430 110.760 ;
        RECT 53.590 110.700 53.910 110.960 ;
        RECT 54.510 110.700 54.830 110.960 ;
        RECT 65.550 110.900 65.870 110.960 ;
        RECT 66.945 110.900 67.235 110.945 ;
        RECT 69.690 110.900 70.010 110.960 ;
        RECT 65.550 110.760 66.700 110.900 ;
        RECT 65.550 110.700 65.870 110.760 ;
        RECT 52.685 110.560 52.975 110.605 ;
        RECT 54.600 110.560 54.740 110.700 ;
        RECT 52.685 110.420 54.740 110.560 ;
        RECT 64.170 110.560 64.490 110.620 ;
        RECT 65.105 110.560 65.395 110.605 ;
        RECT 66.105 110.560 66.395 110.605 ;
        RECT 64.170 110.420 65.395 110.560 ;
        RECT 52.685 110.375 52.975 110.420 ;
        RECT 64.170 110.360 64.490 110.420 ;
        RECT 65.105 110.375 65.395 110.420 ;
        RECT 65.640 110.420 66.395 110.560 ;
        RECT 27.845 110.220 28.135 110.265 ;
        RECT 28.290 110.220 28.610 110.280 ;
        RECT 27.845 110.080 28.610 110.220 ;
        RECT 27.845 110.035 28.135 110.080 ;
        RECT 28.290 110.020 28.610 110.080 ;
        RECT 29.210 110.020 29.530 110.280 ;
        RECT 34.745 110.220 35.035 110.265 ;
        RECT 41.630 110.220 41.950 110.280 ;
        RECT 34.745 110.080 41.950 110.220 ;
        RECT 34.745 110.035 35.035 110.080 ;
        RECT 41.630 110.020 41.950 110.080 ;
        RECT 51.765 110.220 52.055 110.265 ;
        RECT 53.130 110.220 53.450 110.280 ;
        RECT 51.765 110.080 53.450 110.220 ;
        RECT 51.765 110.035 52.055 110.080 ;
        RECT 53.130 110.020 53.450 110.080 ;
        RECT 54.050 110.220 54.370 110.280 ;
        RECT 54.525 110.220 54.815 110.265 ;
        RECT 54.050 110.080 54.815 110.220 ;
        RECT 54.050 110.020 54.370 110.080 ;
        RECT 54.525 110.035 54.815 110.080 ;
        RECT 54.970 110.020 55.290 110.280 ;
        RECT 56.365 110.220 56.655 110.265 ;
        RECT 57.730 110.220 58.050 110.280 ;
        RECT 56.365 110.080 58.050 110.220 ;
        RECT 56.365 110.035 56.655 110.080 ;
        RECT 57.730 110.020 58.050 110.080 ;
        RECT 28.765 109.880 29.055 109.925 ;
        RECT 31.510 109.880 31.830 109.940 ;
        RECT 37.030 109.880 37.350 109.940 ;
        RECT 28.765 109.740 37.350 109.880 ;
        RECT 28.765 109.695 29.055 109.740 ;
        RECT 31.510 109.680 31.830 109.740 ;
        RECT 37.030 109.680 37.350 109.740 ;
        RECT 50.370 109.880 50.690 109.940 ;
        RECT 53.605 109.880 53.895 109.925 ;
        RECT 50.370 109.740 53.895 109.880 ;
        RECT 50.370 109.680 50.690 109.740 ;
        RECT 53.605 109.695 53.895 109.740 ;
        RECT 55.905 109.880 56.195 109.925 ;
        RECT 60.950 109.880 61.270 109.940 ;
        RECT 55.905 109.740 61.270 109.880 ;
        RECT 55.905 109.695 56.195 109.740 ;
        RECT 31.985 109.540 32.275 109.585 ;
        RECT 33.810 109.540 34.130 109.600 ;
        RECT 31.985 109.400 34.130 109.540 ;
        RECT 31.985 109.355 32.275 109.400 ;
        RECT 33.810 109.340 34.130 109.400 ;
        RECT 54.970 109.540 55.290 109.600 ;
        RECT 55.980 109.540 56.120 109.695 ;
        RECT 60.950 109.680 61.270 109.740 ;
        RECT 54.970 109.400 56.120 109.540 ;
        RECT 58.205 109.540 58.495 109.585 ;
        RECT 64.630 109.540 64.950 109.600 ;
        RECT 58.205 109.400 64.950 109.540 ;
        RECT 65.640 109.540 65.780 110.420 ;
        RECT 66.105 110.375 66.395 110.420 ;
        RECT 66.560 110.220 66.700 110.760 ;
        RECT 66.945 110.760 70.010 110.900 ;
        RECT 66.945 110.715 67.235 110.760 ;
        RECT 69.690 110.700 70.010 110.760 ;
        RECT 71.990 110.700 72.310 110.960 ;
        RECT 79.350 110.900 79.670 110.960 ;
        RECT 74.840 110.760 79.670 110.900 ;
        RECT 67.850 110.360 68.170 110.620 ;
        RECT 70.165 110.560 70.455 110.605 ;
        RECT 74.840 110.560 74.980 110.760 ;
        RECT 79.350 110.700 79.670 110.760 ;
        RECT 82.570 110.900 82.890 110.960 ;
        RECT 92.705 110.900 92.995 110.945 ;
        RECT 96.370 110.900 96.690 110.960 ;
        RECT 82.570 110.760 88.780 110.900 ;
        RECT 82.570 110.700 82.890 110.760 ;
        RECT 88.090 110.560 88.410 110.620 ;
        RECT 70.165 110.420 74.980 110.560 ;
        RECT 75.300 110.420 88.410 110.560 ;
        RECT 70.165 110.375 70.455 110.420 ;
        RECT 67.405 110.220 67.695 110.265 ;
        RECT 66.560 110.080 67.695 110.220 ;
        RECT 67.940 110.220 68.080 110.360 ;
        RECT 68.325 110.220 68.615 110.265 ;
        RECT 67.940 110.080 68.615 110.220 ;
        RECT 67.405 110.035 67.695 110.080 ;
        RECT 68.325 110.035 68.615 110.080 ;
        RECT 69.230 110.220 69.550 110.280 ;
        RECT 69.705 110.220 69.995 110.265 ;
        RECT 69.230 110.080 69.995 110.220 ;
        RECT 69.230 110.020 69.550 110.080 ;
        RECT 69.705 110.035 69.995 110.080 ;
        RECT 71.070 110.020 71.390 110.280 ;
        RECT 75.300 110.265 75.440 110.420 ;
        RECT 75.225 110.035 75.515 110.265 ;
        RECT 76.560 110.220 76.850 110.265 ;
        RECT 77.970 110.220 78.290 110.280 ;
        RECT 85.880 110.265 86.020 110.420 ;
        RECT 88.090 110.360 88.410 110.420 ;
        RECT 87.170 110.265 87.490 110.280 ;
        RECT 76.560 110.080 78.290 110.220 ;
        RECT 76.560 110.035 76.850 110.080 ;
        RECT 77.970 110.020 78.290 110.080 ;
        RECT 85.805 110.035 86.095 110.265 ;
        RECT 87.140 110.035 87.490 110.265 ;
        RECT 88.640 110.220 88.780 110.760 ;
        RECT 92.705 110.760 96.690 110.900 ;
        RECT 92.705 110.715 92.995 110.760 ;
        RECT 96.370 110.700 96.690 110.760 ;
        RECT 96.830 110.700 97.150 110.960 ;
        RECT 98.685 110.900 98.975 110.945 ;
        RECT 98.685 110.760 103.040 110.900 ;
        RECT 98.685 110.715 98.975 110.760 ;
        RECT 91.310 110.560 91.630 110.620 ;
        RECT 91.310 110.420 99.360 110.560 ;
        RECT 91.310 110.360 91.630 110.420 ;
        RECT 88.640 110.080 97.060 110.220 ;
        RECT 87.170 110.020 87.490 110.035 ;
        RECT 66.010 109.880 66.330 109.940 ;
        RECT 67.865 109.880 68.155 109.925 ;
        RECT 66.010 109.740 68.155 109.880 ;
        RECT 66.010 109.680 66.330 109.740 ;
        RECT 67.865 109.695 68.155 109.740 ;
        RECT 76.105 109.880 76.395 109.925 ;
        RECT 77.295 109.880 77.585 109.925 ;
        RECT 79.815 109.880 80.105 109.925 ;
        RECT 76.105 109.740 80.105 109.880 ;
        RECT 76.105 109.695 76.395 109.740 ;
        RECT 77.295 109.695 77.585 109.740 ;
        RECT 79.815 109.695 80.105 109.740 ;
        RECT 86.685 109.880 86.975 109.925 ;
        RECT 87.875 109.880 88.165 109.925 ;
        RECT 90.395 109.880 90.685 109.925 ;
        RECT 86.685 109.740 90.685 109.880 ;
        RECT 86.685 109.695 86.975 109.740 ;
        RECT 87.875 109.695 88.165 109.740 ;
        RECT 90.395 109.695 90.685 109.740 ;
        RECT 96.370 109.680 96.690 109.940 ;
        RECT 96.920 109.880 97.060 110.080 ;
        RECT 97.750 110.020 98.070 110.280 ;
        RECT 99.220 110.265 99.360 110.420 ;
        RECT 99.145 110.035 99.435 110.265 ;
        RECT 99.680 109.880 99.820 110.760 ;
        RECT 102.900 110.620 103.040 110.760 ;
        RECT 104.650 110.700 104.970 110.960 ;
        RECT 118.465 110.900 118.755 110.945 ;
        RECT 119.830 110.900 120.150 110.960 ;
        RECT 115.780 110.760 120.150 110.900 ;
        RECT 102.810 110.560 103.130 110.620 ;
        RECT 106.505 110.560 106.795 110.605 ;
        RECT 102.810 110.420 106.795 110.560 ;
        RECT 102.810 110.360 103.130 110.420 ;
        RECT 106.505 110.375 106.795 110.420 ;
        RECT 100.510 110.020 100.830 110.280 ;
        RECT 100.970 110.220 101.290 110.280 ;
        RECT 101.445 110.220 101.735 110.265 ;
        RECT 100.970 110.080 101.735 110.220 ;
        RECT 100.970 110.020 101.290 110.080 ;
        RECT 101.445 110.035 101.735 110.080 ;
        RECT 105.570 110.020 105.890 110.280 ;
        RECT 106.965 110.035 107.255 110.265 ;
        RECT 108.345 110.220 108.635 110.265 ;
        RECT 109.250 110.220 109.570 110.280 ;
        RECT 115.780 110.265 115.920 110.760 ;
        RECT 118.465 110.715 118.755 110.760 ;
        RECT 119.830 110.700 120.150 110.760 ;
        RECT 122.130 110.900 122.450 110.960 ;
        RECT 128.570 110.900 128.890 110.960 ;
        RECT 122.130 110.760 128.890 110.900 ;
        RECT 122.130 110.700 122.450 110.760 ;
        RECT 128.570 110.700 128.890 110.760 ;
        RECT 129.950 110.700 130.270 110.960 ;
        RECT 132.250 110.700 132.570 110.960 ;
        RECT 135.930 110.900 136.250 110.960 ;
        RECT 137.310 110.900 137.630 110.960 ;
        RECT 133.720 110.760 137.630 110.900 ;
        RECT 117.990 110.360 118.310 110.620 ;
        RECT 123.970 110.605 124.290 110.620 ;
        RECT 123.970 110.560 124.320 110.605 ;
        RECT 123.820 110.420 124.320 110.560 ;
        RECT 123.970 110.375 124.320 110.420 ;
        RECT 127.650 110.560 127.970 110.620 ;
        RECT 130.040 110.560 130.180 110.700 ;
        RECT 133.720 110.560 133.860 110.760 ;
        RECT 135.930 110.700 136.250 110.760 ;
        RECT 137.310 110.700 137.630 110.760 ;
        RECT 137.770 110.900 138.090 110.960 ;
        RECT 142.830 110.900 143.150 110.960 ;
        RECT 137.770 110.760 143.150 110.900 ;
        RECT 137.770 110.700 138.090 110.760 ;
        RECT 142.830 110.700 143.150 110.760 ;
        RECT 150.650 110.900 150.970 110.960 ;
        RECT 152.045 110.900 152.335 110.945 ;
        RECT 150.650 110.760 152.335 110.900 ;
        RECT 150.650 110.700 150.970 110.760 ;
        RECT 152.045 110.715 152.335 110.760 ;
        RECT 127.650 110.420 133.860 110.560 ;
        RECT 134.060 110.560 134.350 110.605 ;
        RECT 135.010 110.560 135.330 110.620 ;
        RECT 134.060 110.420 135.330 110.560 ;
        RECT 123.970 110.360 124.290 110.375 ;
        RECT 127.650 110.360 127.970 110.420 ;
        RECT 134.060 110.375 134.350 110.420 ;
        RECT 135.010 110.360 135.330 110.420 ;
        RECT 145.760 110.560 146.050 110.605 ;
        RECT 147.445 110.560 147.735 110.605 ;
        RECT 145.760 110.420 147.735 110.560 ;
        RECT 145.760 110.375 146.050 110.420 ;
        RECT 147.445 110.375 147.735 110.420 ;
        RECT 108.345 110.080 109.570 110.220 ;
        RECT 108.345 110.035 108.635 110.080 ;
        RECT 96.920 109.740 99.820 109.880 ;
        RECT 107.040 109.880 107.180 110.035 ;
        RECT 109.250 110.020 109.570 110.080 ;
        RECT 115.605 110.080 115.920 110.265 ;
        RECT 116.165 110.220 116.455 110.265 ;
        RECT 120.290 110.220 120.610 110.280 ;
        RECT 116.165 110.080 120.610 110.220 ;
        RECT 115.605 110.035 115.895 110.080 ;
        RECT 116.165 110.035 116.455 110.080 ;
        RECT 120.290 110.020 120.610 110.080 ;
        RECT 125.365 110.220 125.655 110.265 ;
        RECT 129.950 110.220 130.270 110.280 ;
        RECT 132.725 110.220 133.015 110.265 ;
        RECT 125.365 110.080 133.015 110.220 ;
        RECT 125.365 110.035 125.655 110.080 ;
        RECT 129.950 110.020 130.270 110.080 ;
        RECT 132.725 110.035 133.015 110.080 ;
        RECT 155.250 110.020 155.570 110.280 ;
        RECT 112.010 109.880 112.330 109.940 ;
        RECT 117.545 109.880 117.835 109.925 ;
        RECT 107.040 109.740 112.330 109.880 ;
        RECT 112.010 109.680 112.330 109.740 ;
        RECT 117.160 109.740 117.835 109.880 ;
        RECT 68.770 109.540 69.090 109.600 ;
        RECT 71.530 109.540 71.850 109.600 ;
        RECT 74.750 109.540 75.070 109.600 ;
        RECT 65.640 109.400 75.070 109.540 ;
        RECT 54.970 109.340 55.290 109.400 ;
        RECT 58.205 109.355 58.495 109.400 ;
        RECT 64.630 109.340 64.950 109.400 ;
        RECT 68.770 109.340 69.090 109.400 ;
        RECT 71.530 109.340 71.850 109.400 ;
        RECT 74.750 109.340 75.070 109.400 ;
        RECT 75.710 109.540 76.000 109.585 ;
        RECT 77.810 109.540 78.100 109.585 ;
        RECT 79.380 109.540 79.670 109.585 ;
        RECT 86.290 109.540 86.580 109.585 ;
        RECT 88.390 109.540 88.680 109.585 ;
        RECT 89.960 109.540 90.250 109.585 ;
        RECT 114.785 109.540 115.075 109.585 ;
        RECT 75.710 109.400 79.670 109.540 ;
        RECT 75.710 109.355 76.000 109.400 ;
        RECT 77.810 109.355 78.100 109.400 ;
        RECT 79.380 109.355 79.670 109.400 ;
        RECT 81.740 109.400 85.100 109.540 ;
        RECT 32.430 109.200 32.750 109.260 ;
        RECT 32.905 109.200 33.195 109.245 ;
        RECT 33.350 109.200 33.670 109.260 ;
        RECT 32.430 109.060 33.670 109.200 ;
        RECT 32.430 109.000 32.750 109.060 ;
        RECT 32.905 109.015 33.195 109.060 ;
        RECT 33.350 109.000 33.670 109.060 ;
        RECT 50.830 109.000 51.150 109.260 ;
        RECT 65.550 109.200 65.870 109.260 ;
        RECT 66.025 109.200 66.315 109.245 ;
        RECT 65.550 109.060 66.315 109.200 ;
        RECT 65.550 109.000 65.870 109.060 ;
        RECT 66.025 109.015 66.315 109.060 ;
        RECT 66.470 109.200 66.790 109.260 ;
        RECT 81.740 109.200 81.880 109.400 ;
        RECT 66.470 109.060 81.880 109.200 ;
        RECT 82.125 109.200 82.415 109.245 ;
        RECT 84.410 109.200 84.730 109.260 ;
        RECT 82.125 109.060 84.730 109.200 ;
        RECT 84.960 109.200 85.100 109.400 ;
        RECT 86.290 109.400 90.250 109.540 ;
        RECT 86.290 109.355 86.580 109.400 ;
        RECT 88.390 109.355 88.680 109.400 ;
        RECT 89.960 109.355 90.250 109.400 ;
        RECT 92.320 109.400 93.840 109.540 ;
        RECT 92.320 109.200 92.460 109.400 ;
        RECT 84.960 109.060 92.460 109.200 ;
        RECT 66.470 109.000 66.790 109.060 ;
        RECT 82.125 109.015 82.415 109.060 ;
        RECT 84.410 109.000 84.730 109.060 ;
        RECT 93.150 109.000 93.470 109.260 ;
        RECT 93.700 109.200 93.840 109.400 ;
        RECT 100.140 109.400 101.200 109.540 ;
        RECT 100.140 109.200 100.280 109.400 ;
        RECT 93.700 109.060 100.280 109.200 ;
        RECT 100.510 109.000 100.830 109.260 ;
        RECT 101.060 109.200 101.200 109.400 ;
        RECT 107.500 109.400 115.075 109.540 ;
        RECT 107.500 109.200 107.640 109.400 ;
        RECT 114.785 109.355 115.075 109.400 ;
        RECT 101.060 109.060 107.640 109.200 ;
        RECT 107.885 109.200 108.175 109.245 ;
        RECT 109.250 109.200 109.570 109.260 ;
        RECT 107.885 109.060 109.570 109.200 ;
        RECT 107.885 109.015 108.175 109.060 ;
        RECT 109.250 109.000 109.570 109.060 ;
        RECT 109.710 109.200 110.030 109.260 ;
        RECT 117.160 109.200 117.300 109.740 ;
        RECT 117.545 109.695 117.835 109.740 ;
        RECT 120.775 109.880 121.065 109.925 ;
        RECT 123.295 109.880 123.585 109.925 ;
        RECT 124.485 109.880 124.775 109.925 ;
        RECT 120.775 109.740 124.775 109.880 ;
        RECT 120.775 109.695 121.065 109.740 ;
        RECT 123.295 109.695 123.585 109.740 ;
        RECT 124.485 109.695 124.775 109.740 ;
        RECT 129.505 109.880 129.795 109.925 ;
        RECT 131.790 109.880 132.110 109.940 ;
        RECT 129.505 109.740 132.110 109.880 ;
        RECT 129.505 109.695 129.795 109.740 ;
        RECT 131.790 109.680 132.110 109.740 ;
        RECT 133.605 109.880 133.895 109.925 ;
        RECT 134.795 109.880 135.085 109.925 ;
        RECT 137.315 109.880 137.605 109.925 ;
        RECT 133.605 109.740 137.605 109.880 ;
        RECT 133.605 109.695 133.895 109.740 ;
        RECT 134.795 109.695 135.085 109.740 ;
        RECT 137.315 109.695 137.605 109.740 ;
        RECT 142.395 109.880 142.685 109.925 ;
        RECT 144.915 109.880 145.205 109.925 ;
        RECT 146.105 109.880 146.395 109.925 ;
        RECT 142.395 109.740 146.395 109.880 ;
        RECT 142.395 109.695 142.685 109.740 ;
        RECT 144.915 109.695 145.205 109.740 ;
        RECT 146.105 109.695 146.395 109.740 ;
        RECT 146.985 109.880 147.275 109.925 ;
        RECT 147.890 109.880 148.210 109.940 ;
        RECT 146.985 109.740 148.210 109.880 ;
        RECT 146.985 109.695 147.275 109.740 ;
        RECT 147.890 109.680 148.210 109.740 ;
        RECT 150.190 109.680 150.510 109.940 ;
        RECT 121.210 109.540 121.500 109.585 ;
        RECT 122.780 109.540 123.070 109.585 ;
        RECT 124.880 109.540 125.170 109.585 ;
        RECT 121.210 109.400 125.170 109.540 ;
        RECT 121.210 109.355 121.500 109.400 ;
        RECT 122.780 109.355 123.070 109.400 ;
        RECT 124.880 109.355 125.170 109.400 ;
        RECT 133.210 109.540 133.500 109.585 ;
        RECT 135.310 109.540 135.600 109.585 ;
        RECT 136.880 109.540 137.170 109.585 ;
        RECT 133.210 109.400 137.170 109.540 ;
        RECT 133.210 109.355 133.500 109.400 ;
        RECT 135.310 109.355 135.600 109.400 ;
        RECT 136.880 109.355 137.170 109.400 ;
        RECT 137.770 109.540 138.090 109.600 ;
        RECT 140.085 109.540 140.375 109.585 ;
        RECT 137.770 109.400 140.375 109.540 ;
        RECT 137.770 109.340 138.090 109.400 ;
        RECT 140.085 109.355 140.375 109.400 ;
        RECT 142.830 109.540 143.120 109.585 ;
        RECT 144.400 109.540 144.690 109.585 ;
        RECT 146.500 109.540 146.790 109.585 ;
        RECT 142.830 109.400 146.790 109.540 ;
        RECT 142.830 109.355 143.120 109.400 ;
        RECT 144.400 109.355 144.690 109.400 ;
        RECT 146.500 109.355 146.790 109.400 ;
        RECT 122.130 109.200 122.450 109.260 ;
        RECT 109.710 109.060 122.450 109.200 ;
        RECT 109.710 109.000 110.030 109.060 ;
        RECT 122.130 109.000 122.450 109.060 ;
        RECT 128.110 109.200 128.430 109.260 ;
        RECT 130.870 109.200 131.190 109.260 ;
        RECT 128.110 109.060 131.190 109.200 ;
        RECT 128.110 109.000 128.430 109.060 ;
        RECT 130.870 109.000 131.190 109.060 ;
        RECT 138.230 109.200 138.550 109.260 ;
        RECT 139.625 109.200 139.915 109.245 ;
        RECT 138.230 109.060 139.915 109.200 ;
        RECT 138.230 109.000 138.550 109.060 ;
        RECT 139.625 109.015 139.915 109.060 ;
        RECT 146.970 109.200 147.290 109.260 ;
        RECT 155.250 109.200 155.570 109.260 ;
        RECT 146.970 109.060 155.570 109.200 ;
        RECT 146.970 109.000 147.290 109.060 ;
        RECT 155.250 109.000 155.570 109.060 ;
        RECT 22.700 108.380 157.020 108.860 ;
        RECT 37.490 107.980 37.810 108.240 ;
        RECT 46.705 108.180 46.995 108.225 ;
        RECT 50.830 108.180 51.150 108.240 ;
        RECT 46.705 108.040 51.150 108.180 ;
        RECT 46.705 107.995 46.995 108.040 ;
        RECT 50.830 107.980 51.150 108.040 ;
        RECT 76.590 108.180 76.910 108.240 ;
        RECT 84.870 108.180 85.190 108.240 ;
        RECT 76.590 108.040 85.190 108.180 ;
        RECT 76.590 107.980 76.910 108.040 ;
        RECT 84.870 107.980 85.190 108.040 ;
        RECT 87.170 108.180 87.490 108.240 ;
        RECT 88.105 108.180 88.395 108.225 ;
        RECT 87.170 108.040 88.395 108.180 ;
        RECT 87.170 107.980 87.490 108.040 ;
        RECT 88.105 107.995 88.395 108.040 ;
        RECT 91.785 108.180 92.075 108.225 ;
        RECT 93.150 108.180 93.470 108.240 ;
        RECT 91.785 108.040 93.470 108.180 ;
        RECT 91.785 107.995 92.075 108.040 ;
        RECT 93.150 107.980 93.470 108.040 ;
        RECT 100.985 108.180 101.275 108.225 ;
        RECT 102.365 108.180 102.655 108.225 ;
        RECT 114.310 108.180 114.630 108.240 ;
        RECT 100.985 108.040 102.655 108.180 ;
        RECT 100.985 107.995 101.275 108.040 ;
        RECT 102.365 107.995 102.655 108.040 ;
        RECT 104.740 108.040 114.630 108.180 ;
        RECT 49.925 107.840 50.215 107.885 ;
        RECT 68.770 107.840 69.090 107.900 ;
        RECT 76.130 107.840 76.450 107.900 ;
        RECT 81.190 107.840 81.510 107.900 ;
        RECT 104.740 107.840 104.880 108.040 ;
        RECT 114.310 107.980 114.630 108.040 ;
        RECT 120.290 107.980 120.610 108.240 ;
        RECT 120.765 108.180 121.055 108.225 ;
        RECT 125.350 108.180 125.670 108.240 ;
        RECT 120.765 108.040 125.670 108.180 ;
        RECT 120.765 107.995 121.055 108.040 ;
        RECT 125.350 107.980 125.670 108.040 ;
        RECT 146.970 107.980 147.290 108.240 ;
        RECT 154.330 108.180 154.650 108.240 ;
        RECT 147.520 108.040 154.650 108.180 ;
        RECT 47.240 107.700 53.360 107.840 ;
        RECT 34.730 107.500 35.050 107.560 ;
        RECT 34.730 107.360 36.800 107.500 ;
        RECT 34.730 107.300 35.050 107.360 ;
        RECT 32.445 107.160 32.735 107.205 ;
        RECT 32.890 107.160 33.210 107.220 ;
        RECT 32.445 107.020 33.210 107.160 ;
        RECT 32.445 106.975 32.735 107.020 ;
        RECT 32.890 106.960 33.210 107.020 ;
        RECT 33.810 106.960 34.130 107.220 ;
        RECT 36.125 107.160 36.415 107.205 ;
        RECT 34.820 107.020 36.415 107.160 ;
        RECT 34.820 106.540 34.960 107.020 ;
        RECT 36.125 106.975 36.415 107.020 ;
        RECT 36.660 106.820 36.800 107.360 ;
        RECT 37.030 107.160 37.350 107.220 ;
        RECT 39.805 107.160 40.095 107.205 ;
        RECT 37.030 107.020 40.095 107.160 ;
        RECT 37.030 106.960 37.350 107.020 ;
        RECT 39.805 106.975 40.095 107.020 ;
        RECT 40.725 107.160 41.015 107.205 ;
        RECT 41.185 107.160 41.475 107.205 ;
        RECT 40.725 107.020 41.475 107.160 ;
        RECT 40.725 106.975 41.015 107.020 ;
        RECT 41.185 106.975 41.475 107.020 ;
        RECT 43.930 106.960 44.250 107.220 ;
        RECT 37.490 106.820 37.810 106.880 ;
        RECT 36.660 106.680 37.810 106.820 ;
        RECT 37.490 106.620 37.810 106.680 ;
        RECT 46.625 106.820 46.915 106.865 ;
        RECT 47.240 106.820 47.380 107.700 ;
        RECT 49.925 107.655 50.215 107.700 ;
        RECT 48.085 107.500 48.375 107.545 ;
        RECT 50.845 107.500 51.135 107.545 ;
        RECT 48.085 107.360 51.135 107.500 ;
        RECT 48.085 107.315 48.375 107.360 ;
        RECT 50.845 107.315 51.135 107.360 ;
        RECT 53.220 107.220 53.360 107.700 ;
        RECT 68.770 107.700 76.450 107.840 ;
        RECT 68.770 107.640 69.090 107.700 ;
        RECT 76.130 107.640 76.450 107.700 ;
        RECT 79.900 107.700 80.960 107.840 ;
        RECT 54.970 107.300 55.290 107.560 ;
        RECT 69.230 107.500 69.550 107.560 ;
        RECT 65.640 107.360 67.160 107.500 ;
        RECT 65.640 107.220 65.780 107.360 ;
        RECT 49.005 107.160 49.295 107.205 ;
        RECT 49.910 107.160 50.230 107.220 ;
        RECT 47.700 107.020 50.230 107.160 ;
        RECT 47.700 106.865 47.840 107.020 ;
        RECT 49.005 106.975 49.295 107.020 ;
        RECT 49.910 106.960 50.230 107.020 ;
        RECT 50.385 107.160 50.675 107.205 ;
        RECT 50.385 107.020 52.900 107.160 ;
        RECT 50.385 106.975 50.675 107.020 ;
        RECT 52.760 106.865 52.900 107.020 ;
        RECT 53.130 106.960 53.450 107.220 ;
        RECT 54.050 107.160 54.370 107.220 ;
        RECT 55.445 107.160 55.735 107.205 ;
        RECT 54.050 107.020 55.735 107.160 ;
        RECT 54.050 106.960 54.370 107.020 ;
        RECT 55.445 106.975 55.735 107.020 ;
        RECT 64.630 106.960 64.950 107.220 ;
        RECT 65.105 107.160 65.395 107.205 ;
        RECT 65.550 107.160 65.870 107.220 ;
        RECT 65.105 107.020 65.870 107.160 ;
        RECT 65.105 106.975 65.395 107.020 ;
        RECT 65.550 106.960 65.870 107.020 ;
        RECT 66.010 106.960 66.330 107.220 ;
        RECT 66.470 106.960 66.790 107.220 ;
        RECT 67.020 107.205 67.160 107.360 ;
        RECT 69.230 107.360 73.140 107.500 ;
        RECT 69.230 107.300 69.550 107.360 ;
        RECT 66.945 106.975 67.235 107.205 ;
        RECT 67.390 107.160 67.710 107.220 ;
        RECT 67.865 107.160 68.155 107.205 ;
        RECT 67.390 107.020 68.155 107.160 ;
        RECT 67.390 106.960 67.710 107.020 ;
        RECT 67.865 106.975 68.155 107.020 ;
        RECT 71.530 106.960 71.850 107.220 ;
        RECT 73.000 107.205 73.140 107.360 ;
        RECT 72.925 106.975 73.215 107.205 ;
        RECT 74.290 106.960 74.610 107.220 ;
        RECT 76.130 107.160 76.450 107.220 ;
        RECT 79.900 107.205 80.040 107.700 ;
        RECT 80.820 107.500 80.960 107.700 ;
        RECT 81.190 107.700 97.980 107.840 ;
        RECT 81.190 107.640 81.510 107.700 ;
        RECT 83.950 107.500 84.270 107.560 ;
        RECT 80.820 107.360 84.270 107.500 ;
        RECT 83.950 107.300 84.270 107.360 ;
        RECT 84.410 107.300 84.730 107.560 ;
        RECT 84.870 107.500 85.190 107.560 ;
        RECT 84.870 107.360 97.520 107.500 ;
        RECT 84.870 107.300 85.190 107.360 ;
        RECT 78.445 107.160 78.735 107.205 ;
        RECT 76.130 107.020 78.735 107.160 ;
        RECT 76.130 106.960 76.450 107.020 ;
        RECT 78.445 106.975 78.735 107.020 ;
        RECT 79.365 106.975 79.655 107.205 ;
        RECT 79.825 106.975 80.115 107.205 ;
        RECT 46.625 106.680 47.380 106.820 ;
        RECT 46.625 106.635 46.915 106.680 ;
        RECT 47.625 106.635 47.915 106.865 ;
        RECT 52.685 106.820 52.975 106.865 ;
        RECT 58.190 106.820 58.510 106.880 ;
        RECT 52.685 106.680 58.510 106.820 ;
        RECT 64.720 106.820 64.860 106.960 ;
        RECT 79.440 106.820 79.580 106.975 ;
        RECT 80.730 106.960 81.050 107.220 ;
        RECT 81.265 107.160 81.555 107.205 ;
        RECT 84.500 107.160 84.640 107.300 ;
        RECT 85.345 107.160 85.635 107.205 ;
        RECT 81.265 107.020 83.720 107.160 ;
        RECT 84.500 107.020 85.635 107.160 ;
        RECT 81.265 106.975 81.555 107.020 ;
        RECT 80.270 106.820 80.590 106.880 ;
        RECT 64.720 106.680 80.590 106.820 ;
        RECT 83.580 106.820 83.720 107.020 ;
        RECT 85.345 106.975 85.635 107.020 ;
        RECT 86.250 106.960 86.570 107.220 ;
        RECT 89.025 106.975 89.315 107.205 ;
        RECT 85.805 106.820 86.095 106.865 ;
        RECT 83.580 106.680 86.095 106.820 ;
        RECT 89.100 106.820 89.240 106.975 ;
        RECT 89.930 106.960 90.250 107.220 ;
        RECT 90.405 107.160 90.695 107.205 ;
        RECT 91.310 107.160 91.630 107.220 ;
        RECT 93.610 107.160 93.930 107.220 ;
        RECT 96.830 107.160 97.150 107.220 ;
        RECT 90.405 107.020 91.630 107.160 ;
        RECT 90.405 106.975 90.695 107.020 ;
        RECT 91.310 106.960 91.630 107.020 ;
        RECT 92.780 107.020 97.150 107.160 ;
        RECT 92.780 106.880 92.920 107.020 ;
        RECT 93.610 106.960 93.930 107.020 ;
        RECT 96.830 106.960 97.150 107.020 ;
        RECT 89.100 106.680 91.080 106.820 ;
        RECT 52.685 106.635 52.975 106.680 ;
        RECT 58.190 106.620 58.510 106.680 ;
        RECT 80.270 106.620 80.590 106.680 ;
        RECT 85.805 106.635 86.095 106.680 ;
        RECT 31.510 106.480 31.830 106.540 ;
        RECT 32.905 106.480 33.195 106.525 ;
        RECT 31.510 106.340 33.195 106.480 ;
        RECT 31.510 106.280 31.830 106.340 ;
        RECT 32.905 106.295 33.195 106.340 ;
        RECT 34.730 106.280 35.050 106.540 ;
        RECT 36.585 106.480 36.875 106.525 ;
        RECT 37.950 106.480 38.270 106.540 ;
        RECT 39.805 106.480 40.095 106.525 ;
        RECT 36.585 106.340 40.095 106.480 ;
        RECT 36.585 106.295 36.875 106.340 ;
        RECT 37.950 106.280 38.270 106.340 ;
        RECT 39.805 106.295 40.095 106.340 ;
        RECT 45.310 106.480 45.630 106.540 ;
        RECT 45.785 106.480 46.075 106.525 ;
        RECT 45.310 106.340 46.075 106.480 ;
        RECT 45.310 106.280 45.630 106.340 ;
        RECT 45.785 106.295 46.075 106.340 ;
        RECT 51.290 106.480 51.610 106.540 ;
        RECT 52.225 106.480 52.515 106.525 ;
        RECT 51.290 106.340 52.515 106.480 ;
        RECT 51.290 106.280 51.610 106.340 ;
        RECT 52.225 106.295 52.515 106.340 ;
        RECT 57.270 106.280 57.590 106.540 ;
        RECT 63.725 106.480 64.015 106.525 ;
        RECT 64.170 106.480 64.490 106.540 ;
        RECT 63.725 106.340 64.490 106.480 ;
        RECT 63.725 106.295 64.015 106.340 ;
        RECT 64.170 106.280 64.490 106.340 ;
        RECT 64.630 106.480 64.950 106.540 ;
        RECT 67.405 106.480 67.695 106.525 ;
        RECT 64.630 106.340 67.695 106.480 ;
        RECT 64.630 106.280 64.950 106.340 ;
        RECT 67.405 106.295 67.695 106.340 ;
        RECT 70.610 106.280 70.930 106.540 ;
        RECT 72.465 106.480 72.755 106.525 ;
        RECT 75.210 106.480 75.530 106.540 ;
        RECT 72.465 106.340 75.530 106.480 ;
        RECT 72.465 106.295 72.755 106.340 ;
        RECT 75.210 106.280 75.530 106.340 ;
        RECT 75.670 106.480 75.990 106.540 ;
        RECT 77.525 106.480 77.815 106.525 ;
        RECT 75.670 106.340 77.815 106.480 ;
        RECT 75.670 106.280 75.990 106.340 ;
        RECT 77.525 106.295 77.815 106.340 ;
        RECT 81.190 106.480 81.510 106.540 ;
        RECT 90.940 106.525 91.080 106.680 ;
        RECT 92.690 106.620 93.010 106.880 ;
        RECT 97.380 106.820 97.520 107.360 ;
        RECT 97.840 107.205 97.980 107.700 ;
        RECT 101.520 107.700 104.880 107.840 ;
        RECT 97.765 106.975 98.055 107.205 ;
        RECT 98.210 106.960 98.530 107.220 ;
        RECT 99.130 106.960 99.450 107.220 ;
        RECT 99.605 107.160 99.895 107.205 ;
        RECT 100.970 107.160 101.290 107.220 ;
        RECT 99.605 107.020 101.290 107.160 ;
        RECT 99.605 106.975 99.895 107.020 ;
        RECT 100.970 106.960 101.290 107.020 ;
        RECT 100.050 106.820 100.370 106.880 ;
        RECT 101.520 106.820 101.660 107.700 ;
        RECT 105.110 107.640 105.430 107.900 ;
        RECT 109.710 107.840 110.030 107.900 ;
        RECT 108.420 107.700 110.030 107.840 ;
        RECT 105.200 107.500 105.340 107.640 ;
        RECT 106.965 107.500 107.255 107.545 ;
        RECT 105.200 107.360 107.255 107.500 ;
        RECT 106.965 107.315 107.255 107.360 ;
        RECT 105.110 107.160 105.430 107.220 ;
        RECT 107.425 107.160 107.715 107.205 ;
        RECT 105.110 107.020 107.715 107.160 ;
        RECT 108.420 107.160 108.560 107.700 ;
        RECT 109.710 107.640 110.030 107.700 ;
        RECT 113.890 107.840 114.180 107.885 ;
        RECT 115.990 107.840 116.280 107.885 ;
        RECT 117.560 107.840 117.850 107.885 ;
        RECT 113.890 107.700 117.850 107.840 ;
        RECT 113.890 107.655 114.180 107.700 ;
        RECT 115.990 107.655 116.280 107.700 ;
        RECT 117.560 107.655 117.850 107.700 ;
        RECT 122.130 107.840 122.450 107.900 ;
        RECT 123.065 107.840 123.355 107.885 ;
        RECT 122.130 107.700 123.355 107.840 ;
        RECT 122.130 107.640 122.450 107.700 ;
        RECT 123.065 107.655 123.355 107.700 ;
        RECT 125.810 107.840 126.100 107.885 ;
        RECT 127.380 107.840 127.670 107.885 ;
        RECT 129.480 107.840 129.770 107.885 ;
        RECT 147.520 107.840 147.660 108.040 ;
        RECT 154.330 107.980 154.650 108.040 ;
        RECT 125.810 107.700 129.770 107.840 ;
        RECT 125.810 107.655 126.100 107.700 ;
        RECT 127.380 107.655 127.670 107.700 ;
        RECT 129.480 107.655 129.770 107.700 ;
        RECT 145.680 107.700 147.660 107.840 ;
        RECT 147.930 107.840 148.220 107.885 ;
        RECT 150.030 107.840 150.320 107.885 ;
        RECT 151.600 107.840 151.890 107.885 ;
        RECT 147.930 107.700 151.890 107.840 ;
        RECT 108.790 107.500 109.110 107.560 ;
        RECT 113.405 107.500 113.695 107.545 ;
        RECT 108.790 107.360 113.695 107.500 ;
        RECT 108.790 107.300 109.110 107.360 ;
        RECT 113.405 107.315 113.695 107.360 ;
        RECT 114.285 107.500 114.575 107.545 ;
        RECT 115.475 107.500 115.765 107.545 ;
        RECT 117.995 107.500 118.285 107.545 ;
        RECT 114.285 107.360 118.285 107.500 ;
        RECT 114.285 107.315 114.575 107.360 ;
        RECT 115.475 107.315 115.765 107.360 ;
        RECT 117.995 107.315 118.285 107.360 ;
        RECT 125.375 107.500 125.665 107.545 ;
        RECT 127.895 107.500 128.185 107.545 ;
        RECT 129.085 107.500 129.375 107.545 ;
        RECT 125.375 107.360 129.375 107.500 ;
        RECT 125.375 107.315 125.665 107.360 ;
        RECT 127.895 107.315 128.185 107.360 ;
        RECT 129.085 107.315 129.375 107.360 ;
        RECT 130.410 107.300 130.730 107.560 ;
        RECT 132.250 107.500 132.570 107.560 ;
        RECT 134.090 107.500 134.410 107.560 ;
        RECT 141.450 107.500 141.770 107.560 ;
        RECT 143.750 107.500 144.070 107.560 ;
        RECT 132.250 107.360 144.070 107.500 ;
        RECT 132.250 107.300 132.570 107.360 ;
        RECT 134.090 107.300 134.410 107.360 ;
        RECT 108.420 107.020 109.020 107.160 ;
        RECT 105.110 106.960 105.430 107.020 ;
        RECT 107.425 106.975 107.715 107.020 ;
        RECT 108.880 106.865 109.020 107.020 ;
        RECT 109.250 106.960 109.570 107.220 ;
        RECT 110.645 106.975 110.935 107.205 ;
        RECT 111.090 107.160 111.410 107.220 ;
        RECT 111.565 107.160 111.855 107.205 ;
        RECT 111.090 107.020 111.855 107.160 ;
        RECT 97.380 106.680 100.370 106.820 ;
        RECT 100.050 106.620 100.370 106.680 ;
        RECT 101.060 106.680 101.660 106.820 ;
        RECT 101.980 106.680 108.560 106.820 ;
        RECT 91.770 106.525 92.090 106.540 ;
        RECT 81.665 106.480 81.955 106.525 ;
        RECT 81.190 106.340 81.955 106.480 ;
        RECT 81.190 106.280 81.510 106.340 ;
        RECT 81.665 106.295 81.955 106.340 ;
        RECT 90.865 106.295 91.155 106.525 ;
        RECT 91.705 106.295 92.090 106.525 ;
        RECT 91.770 106.280 92.090 106.295 ;
        RECT 96.830 106.280 97.150 106.540 ;
        RECT 101.060 106.525 101.200 106.680 ;
        RECT 101.980 106.525 102.120 106.680 ;
        RECT 101.060 106.340 101.355 106.525 ;
        RECT 101.065 106.295 101.355 106.340 ;
        RECT 101.905 106.295 102.195 106.525 ;
        RECT 106.030 106.280 106.350 106.540 ;
        RECT 108.420 106.480 108.560 106.680 ;
        RECT 108.805 106.635 109.095 106.865 ;
        RECT 110.720 106.820 110.860 106.975 ;
        RECT 111.090 106.960 111.410 107.020 ;
        RECT 111.565 106.975 111.855 107.020 ;
        RECT 112.010 106.960 112.330 107.220 ;
        RECT 121.670 106.960 121.990 107.220 ;
        RECT 122.145 107.160 122.435 107.205 ;
        RECT 124.890 107.160 125.210 107.220 ;
        RECT 122.145 107.020 125.210 107.160 ;
        RECT 122.145 106.975 122.435 107.020 ;
        RECT 124.890 106.960 125.210 107.020 ;
        RECT 129.950 106.960 130.270 107.220 ;
        RECT 133.645 107.160 133.935 107.205 ;
        RECT 135.485 107.160 135.775 107.205 ;
        RECT 133.645 107.020 135.775 107.160 ;
        RECT 133.645 106.975 133.935 107.020 ;
        RECT 135.485 106.975 135.775 107.020 ;
        RECT 135.945 106.975 136.235 107.205 ;
        RECT 109.340 106.680 110.860 106.820 ;
        RECT 112.470 106.820 112.790 106.880 ;
        RECT 114.630 106.820 114.920 106.865 ;
        RECT 112.470 106.680 114.920 106.820 ;
        RECT 109.340 106.480 109.480 106.680 ;
        RECT 112.470 106.620 112.790 106.680 ;
        RECT 114.630 106.635 114.920 106.680 ;
        RECT 119.370 106.820 119.690 106.880 ;
        RECT 120.765 106.820 121.055 106.865 ;
        RECT 119.370 106.680 121.055 106.820 ;
        RECT 119.370 106.620 119.690 106.680 ;
        RECT 120.765 106.635 121.055 106.680 ;
        RECT 128.740 106.820 129.030 106.865 ;
        RECT 134.105 106.820 134.395 106.865 ;
        RECT 128.740 106.680 134.395 106.820 ;
        RECT 136.020 106.820 136.160 106.975 ;
        RECT 136.390 106.960 136.710 107.220 ;
        RECT 137.400 107.205 137.540 107.360 ;
        RECT 141.450 107.300 141.770 107.360 ;
        RECT 143.750 107.300 144.070 107.360 ;
        RECT 137.325 106.975 137.615 107.205 ;
        RECT 137.770 107.160 138.090 107.220 ;
        RECT 145.680 107.205 145.820 107.700 ;
        RECT 147.930 107.655 148.220 107.700 ;
        RECT 150.030 107.655 150.320 107.700 ;
        RECT 151.600 107.655 151.890 107.700 ;
        RECT 148.325 107.500 148.615 107.545 ;
        RECT 149.515 107.500 149.805 107.545 ;
        RECT 152.035 107.500 152.325 107.545 ;
        RECT 148.325 107.360 152.325 107.500 ;
        RECT 148.325 107.315 148.615 107.360 ;
        RECT 149.515 107.315 149.805 107.360 ;
        RECT 152.035 107.315 152.325 107.360 ;
        RECT 141.005 107.160 141.295 107.205 ;
        RECT 137.770 107.020 141.295 107.160 ;
        RECT 137.770 106.960 138.090 107.020 ;
        RECT 141.005 106.975 141.295 107.020 ;
        RECT 145.605 106.975 145.895 107.205 ;
        RECT 146.065 107.160 146.355 107.205 ;
        RECT 146.510 107.160 146.830 107.220 ;
        RECT 146.065 107.020 146.830 107.160 ;
        RECT 146.065 106.975 146.355 107.020 ;
        RECT 146.510 106.960 146.830 107.020 ;
        RECT 147.445 107.160 147.735 107.205 ;
        RECT 147.890 107.160 148.210 107.220 ;
        RECT 147.445 107.020 148.210 107.160 ;
        RECT 147.445 106.975 147.735 107.020 ;
        RECT 147.890 106.960 148.210 107.020 ;
        RECT 139.150 106.820 139.470 106.880 ;
        RECT 136.020 106.680 139.470 106.820 ;
        RECT 128.740 106.635 129.030 106.680 ;
        RECT 134.105 106.635 134.395 106.680 ;
        RECT 139.150 106.620 139.470 106.680 ;
        RECT 143.750 106.820 144.070 106.880 ;
        RECT 146.985 106.820 147.275 106.865 ;
        RECT 148.670 106.820 148.960 106.865 ;
        RECT 143.750 106.680 147.275 106.820 ;
        RECT 143.750 106.620 144.070 106.680 ;
        RECT 146.985 106.635 147.275 106.680 ;
        RECT 147.520 106.680 148.960 106.820 ;
        RECT 147.520 106.540 147.660 106.680 ;
        RECT 148.670 106.635 148.960 106.680 ;
        RECT 108.420 106.340 109.480 106.480 ;
        RECT 109.710 106.280 110.030 106.540 ;
        RECT 144.210 106.280 144.530 106.540 ;
        RECT 144.670 106.280 144.990 106.540 ;
        RECT 147.430 106.280 147.750 106.540 ;
        RECT 22.700 105.660 157.820 106.140 ;
        RECT 36.570 105.460 36.890 105.520 ;
        RECT 36.200 105.320 36.890 105.460 ;
        RECT 34.270 105.120 34.590 105.180 ;
        RECT 33.900 104.980 34.590 105.120 ;
        RECT 31.985 104.780 32.275 104.825 ;
        RECT 32.890 104.780 33.210 104.840 ;
        RECT 33.900 104.825 34.040 104.980 ;
        RECT 34.270 104.920 34.590 104.980 ;
        RECT 35.160 105.120 35.450 105.165 ;
        RECT 36.200 105.120 36.340 105.320 ;
        RECT 36.570 105.260 36.890 105.320 ;
        RECT 40.725 105.460 41.015 105.505 ;
        RECT 43.930 105.460 44.250 105.520 ;
        RECT 40.725 105.320 44.250 105.460 ;
        RECT 40.725 105.275 41.015 105.320 ;
        RECT 43.930 105.260 44.250 105.320 ;
        RECT 53.130 105.460 53.450 105.520 ;
        RECT 54.985 105.460 55.275 105.505 ;
        RECT 53.130 105.320 55.275 105.460 ;
        RECT 53.130 105.260 53.450 105.320 ;
        RECT 54.985 105.275 55.275 105.320 ;
        RECT 57.270 105.460 57.590 105.520 ;
        RECT 71.530 105.460 71.850 105.520 ;
        RECT 74.765 105.460 75.055 105.505 ;
        RECT 57.270 105.320 71.300 105.460 ;
        RECT 57.270 105.260 57.590 105.320 ;
        RECT 56.365 105.120 56.655 105.165 ;
        RECT 58.190 105.120 58.510 105.180 ;
        RECT 35.160 104.980 36.340 105.120 ;
        RECT 42.180 104.980 56.120 105.120 ;
        RECT 35.160 104.935 35.450 104.980 ;
        RECT 31.985 104.640 33.210 104.780 ;
        RECT 31.985 104.595 32.275 104.640 ;
        RECT 32.890 104.580 33.210 104.640 ;
        RECT 33.825 104.595 34.115 104.825 ;
        RECT 42.180 104.780 42.320 104.980 ;
        RECT 34.360 104.640 42.320 104.780 ;
        RECT 42.520 104.780 42.810 104.825 ;
        RECT 44.390 104.780 44.710 104.840 ;
        RECT 42.520 104.640 44.710 104.780 ;
        RECT 31.065 104.255 31.355 104.485 ;
        RECT 31.140 104.100 31.280 104.255 ;
        RECT 31.510 104.240 31.830 104.500 ;
        RECT 32.445 104.440 32.735 104.485 ;
        RECT 33.350 104.440 33.670 104.500 ;
        RECT 34.360 104.440 34.500 104.640 ;
        RECT 42.520 104.595 42.810 104.640 ;
        RECT 44.390 104.580 44.710 104.640 ;
        RECT 51.290 104.580 51.610 104.840 ;
        RECT 54.510 104.580 54.830 104.840 ;
        RECT 55.445 104.595 55.735 104.825 ;
        RECT 32.445 104.300 33.670 104.440 ;
        RECT 32.445 104.255 32.735 104.300 ;
        RECT 33.350 104.240 33.670 104.300 ;
        RECT 33.900 104.300 34.500 104.440 ;
        RECT 34.705 104.440 34.995 104.485 ;
        RECT 35.895 104.440 36.185 104.485 ;
        RECT 38.415 104.440 38.705 104.485 ;
        RECT 34.705 104.300 38.705 104.440 ;
        RECT 33.900 104.100 34.040 104.300 ;
        RECT 34.705 104.255 34.995 104.300 ;
        RECT 35.895 104.255 36.185 104.300 ;
        RECT 38.415 104.255 38.705 104.300 ;
        RECT 41.170 104.240 41.490 104.500 ;
        RECT 42.065 104.440 42.355 104.485 ;
        RECT 43.255 104.440 43.545 104.485 ;
        RECT 45.775 104.440 46.065 104.485 ;
        RECT 54.050 104.440 54.370 104.500 ;
        RECT 55.520 104.440 55.660 104.595 ;
        RECT 42.065 104.300 46.065 104.440 ;
        RECT 42.065 104.255 42.355 104.300 ;
        RECT 43.255 104.255 43.545 104.300 ;
        RECT 45.775 104.255 46.065 104.300 ;
        RECT 48.160 104.300 55.660 104.440 ;
        RECT 55.980 104.440 56.120 104.980 ;
        RECT 56.365 104.980 58.510 105.120 ;
        RECT 56.365 104.935 56.655 104.980 ;
        RECT 58.190 104.920 58.510 104.980 ;
        RECT 62.880 104.825 63.020 105.320 ;
        RECT 68.280 105.120 68.570 105.165 ;
        RECT 70.610 105.120 70.930 105.180 ;
        RECT 63.340 104.980 65.780 105.120 ;
        RECT 63.340 104.840 63.480 104.980 ;
        RECT 65.640 104.840 65.780 104.980 ;
        RECT 68.280 104.980 70.930 105.120 ;
        RECT 68.280 104.935 68.570 104.980 ;
        RECT 70.610 104.920 70.930 104.980 ;
        RECT 56.825 104.780 57.115 104.825 ;
        RECT 57.285 104.780 57.575 104.825 ;
        RECT 56.825 104.640 57.575 104.780 ;
        RECT 56.825 104.595 57.115 104.640 ;
        RECT 57.285 104.595 57.575 104.640 ;
        RECT 59.660 104.640 62.560 104.780 ;
        RECT 59.660 104.440 59.800 104.640 ;
        RECT 55.980 104.300 59.800 104.440 ;
        RECT 48.160 104.145 48.300 104.300 ;
        RECT 54.050 104.240 54.370 104.300 ;
        RECT 60.030 104.240 60.350 104.500 ;
        RECT 62.420 104.440 62.560 104.640 ;
        RECT 62.805 104.595 63.095 104.825 ;
        RECT 63.250 104.580 63.570 104.840 ;
        RECT 64.185 104.595 64.475 104.825 ;
        RECT 63.710 104.440 64.030 104.500 ;
        RECT 64.260 104.440 64.400 104.595 ;
        RECT 64.630 104.580 64.950 104.840 ;
        RECT 65.550 104.580 65.870 104.840 ;
        RECT 66.485 104.780 66.775 104.825 ;
        RECT 70.150 104.780 70.470 104.840 ;
        RECT 66.485 104.640 70.470 104.780 ;
        RECT 71.160 104.780 71.300 105.320 ;
        RECT 71.530 105.320 75.055 105.460 ;
        RECT 71.530 105.260 71.850 105.320 ;
        RECT 74.765 105.275 75.055 105.320 ;
        RECT 77.525 105.460 77.815 105.505 ;
        RECT 77.970 105.460 78.290 105.520 ;
        RECT 77.525 105.320 78.290 105.460 ;
        RECT 77.525 105.275 77.815 105.320 ;
        RECT 77.970 105.260 78.290 105.320 ;
        RECT 79.350 105.460 79.670 105.520 ;
        RECT 90.850 105.460 91.170 105.520 ;
        RECT 99.130 105.460 99.450 105.520 ;
        RECT 79.350 105.320 91.170 105.460 ;
        RECT 79.350 105.260 79.670 105.320 ;
        RECT 90.850 105.260 91.170 105.320 ;
        RECT 94.620 105.320 99.450 105.460 ;
        RECT 71.990 105.120 72.310 105.180 ;
        RECT 75.525 105.120 75.815 105.165 ;
        RECT 71.990 104.980 75.815 105.120 ;
        RECT 71.990 104.920 72.310 104.980 ;
        RECT 75.525 104.935 75.815 104.980 ;
        RECT 76.590 104.920 76.910 105.180 ;
        RECT 81.125 105.120 81.415 105.165 ;
        RECT 81.650 105.120 81.970 105.180 ;
        RECT 79.440 104.980 81.970 105.120 ;
        RECT 79.440 104.840 79.580 104.980 ;
        RECT 81.125 104.935 81.415 104.980 ;
        RECT 81.650 104.920 81.970 104.980 ;
        RECT 82.125 104.935 82.415 105.165 ;
        RECT 83.950 105.120 84.270 105.180 ;
        RECT 86.250 105.120 86.570 105.180 ;
        RECT 83.950 104.980 86.570 105.120 ;
        RECT 71.160 104.640 76.360 104.780 ;
        RECT 66.485 104.595 66.775 104.640 ;
        RECT 70.150 104.580 70.470 104.640 ;
        RECT 66.010 104.440 66.330 104.500 ;
        RECT 62.420 104.300 63.480 104.440 ;
        RECT 31.140 103.960 34.040 104.100 ;
        RECT 34.310 104.100 34.600 104.145 ;
        RECT 36.410 104.100 36.700 104.145 ;
        RECT 37.980 104.100 38.270 104.145 ;
        RECT 34.310 103.960 38.270 104.100 ;
        RECT 34.310 103.915 34.600 103.960 ;
        RECT 36.410 103.915 36.700 103.960 ;
        RECT 37.980 103.915 38.270 103.960 ;
        RECT 41.670 104.100 41.960 104.145 ;
        RECT 43.770 104.100 44.060 104.145 ;
        RECT 45.340 104.100 45.630 104.145 ;
        RECT 41.670 103.960 45.630 104.100 ;
        RECT 41.670 103.915 41.960 103.960 ;
        RECT 43.770 103.915 44.060 103.960 ;
        RECT 45.340 103.915 45.630 103.960 ;
        RECT 48.085 103.915 48.375 104.145 ;
        RECT 62.330 104.100 62.650 104.160 ;
        RECT 48.620 103.960 62.650 104.100 ;
        RECT 63.340 104.100 63.480 104.300 ;
        RECT 63.710 104.300 66.330 104.440 ;
        RECT 63.710 104.240 64.030 104.300 ;
        RECT 66.010 104.240 66.330 104.300 ;
        RECT 66.930 104.240 67.250 104.500 ;
        RECT 67.825 104.440 68.115 104.485 ;
        RECT 69.015 104.440 69.305 104.485 ;
        RECT 71.535 104.440 71.825 104.485 ;
        RECT 67.825 104.300 71.825 104.440 ;
        RECT 67.825 104.255 68.115 104.300 ;
        RECT 69.015 104.255 69.305 104.300 ;
        RECT 71.535 104.255 71.825 104.300 ;
        RECT 67.430 104.100 67.720 104.145 ;
        RECT 69.530 104.100 69.820 104.145 ;
        RECT 71.100 104.100 71.390 104.145 ;
        RECT 63.340 103.960 67.160 104.100 ;
        RECT 33.350 103.560 33.670 103.820 ;
        RECT 37.490 103.760 37.810 103.820 ;
        RECT 48.620 103.760 48.760 103.960 ;
        RECT 62.330 103.900 62.650 103.960 ;
        RECT 37.490 103.620 48.760 103.760 ;
        RECT 54.065 103.760 54.355 103.805 ;
        RECT 54.510 103.760 54.830 103.820 ;
        RECT 54.065 103.620 54.830 103.760 ;
        RECT 37.490 103.560 37.810 103.620 ;
        RECT 54.065 103.575 54.355 103.620 ;
        RECT 54.510 103.560 54.830 103.620 ;
        RECT 61.870 103.560 62.190 103.820 ;
        RECT 65.090 103.760 65.410 103.820 ;
        RECT 66.485 103.760 66.775 103.805 ;
        RECT 65.090 103.620 66.775 103.760 ;
        RECT 67.020 103.760 67.160 103.960 ;
        RECT 67.430 103.960 71.390 104.100 ;
        RECT 67.430 103.915 67.720 103.960 ;
        RECT 69.530 103.915 69.820 103.960 ;
        RECT 71.100 103.915 71.390 103.960 ;
        RECT 68.770 103.760 69.090 103.820 ;
        RECT 67.020 103.620 69.090 103.760 ;
        RECT 65.090 103.560 65.410 103.620 ;
        RECT 66.485 103.575 66.775 103.620 ;
        RECT 68.770 103.560 69.090 103.620 ;
        RECT 71.530 103.760 71.850 103.820 ;
        RECT 73.845 103.760 74.135 103.805 ;
        RECT 74.290 103.760 74.610 103.820 ;
        RECT 71.530 103.620 74.610 103.760 ;
        RECT 71.530 103.560 71.850 103.620 ;
        RECT 73.845 103.575 74.135 103.620 ;
        RECT 74.290 103.560 74.610 103.620 ;
        RECT 75.670 103.560 75.990 103.820 ;
        RECT 76.220 103.760 76.360 104.640 ;
        RECT 78.445 104.595 78.735 104.825 ;
        RECT 78.520 104.440 78.660 104.595 ;
        RECT 79.350 104.580 79.670 104.840 ;
        RECT 79.810 104.580 80.130 104.840 ;
        RECT 82.200 104.440 82.340 104.935 ;
        RECT 83.950 104.920 84.270 104.980 ;
        RECT 84.960 104.840 85.100 104.980 ;
        RECT 86.250 104.920 86.570 104.980 ;
        RECT 84.870 104.580 85.190 104.840 ;
        RECT 85.790 104.580 86.110 104.840 ;
        RECT 93.150 104.580 93.470 104.840 ;
        RECT 94.620 104.825 94.760 105.320 ;
        RECT 99.130 105.260 99.450 105.320 ;
        RECT 100.050 105.460 100.370 105.520 ;
        RECT 101.905 105.460 102.195 105.505 ;
        RECT 105.110 105.460 105.430 105.520 ;
        RECT 111.550 105.460 111.870 105.520 ;
        RECT 113.785 105.460 114.075 105.505 ;
        RECT 114.310 105.460 114.630 105.520 ;
        RECT 100.050 105.320 101.200 105.460 ;
        RECT 100.050 105.260 100.370 105.320 ;
        RECT 96.370 105.120 96.690 105.180 ;
        RECT 101.060 105.120 101.200 105.320 ;
        RECT 101.905 105.320 105.430 105.460 ;
        RECT 101.905 105.275 102.195 105.320 ;
        RECT 105.110 105.260 105.430 105.320 ;
        RECT 107.040 105.320 112.700 105.460 ;
        RECT 107.040 105.120 107.180 105.320 ;
        RECT 111.550 105.260 111.870 105.320 ;
        RECT 96.370 104.980 100.740 105.120 ;
        RECT 101.060 104.980 107.180 105.120 ;
        RECT 107.580 105.120 107.870 105.165 ;
        RECT 109.710 105.120 110.030 105.180 ;
        RECT 112.010 105.120 112.330 105.180 ;
        RECT 107.580 104.980 110.030 105.120 ;
        RECT 96.370 104.920 96.690 104.980 ;
        RECT 93.625 104.595 93.915 104.825 ;
        RECT 94.545 104.595 94.835 104.825 ;
        RECT 95.005 104.780 95.295 104.825 ;
        RECT 100.050 104.780 100.370 104.840 ;
        RECT 100.600 104.825 100.740 104.980 ;
        RECT 107.580 104.935 107.870 104.980 ;
        RECT 109.710 104.920 110.030 104.980 ;
        RECT 110.260 104.980 112.330 105.120 ;
        RECT 112.560 105.120 112.700 105.320 ;
        RECT 113.785 105.320 114.630 105.460 ;
        RECT 113.785 105.275 114.075 105.320 ;
        RECT 114.310 105.260 114.630 105.320 ;
        RECT 129.965 105.460 130.255 105.505 ;
        RECT 136.390 105.460 136.710 105.520 ;
        RECT 129.965 105.320 136.710 105.460 ;
        RECT 129.965 105.275 130.255 105.320 ;
        RECT 136.390 105.260 136.710 105.320 ;
        RECT 137.310 105.460 137.630 105.520 ;
        RECT 150.650 105.460 150.970 105.520 ;
        RECT 137.310 105.320 144.900 105.460 ;
        RECT 137.310 105.260 137.630 105.320 ;
        RECT 114.785 105.120 115.075 105.165 ;
        RECT 112.560 104.980 115.075 105.120 ;
        RECT 95.005 104.640 100.370 104.780 ;
        RECT 95.005 104.595 95.295 104.640 ;
        RECT 82.570 104.440 82.890 104.500 ;
        RECT 92.690 104.440 93.010 104.500 ;
        RECT 78.520 104.300 80.500 104.440 ;
        RECT 82.200 104.300 93.010 104.440 ;
        RECT 93.700 104.440 93.840 104.595 ;
        RECT 100.050 104.580 100.370 104.640 ;
        RECT 100.525 104.595 100.815 104.825 ;
        RECT 100.970 104.580 101.290 104.840 ;
        RECT 110.260 104.825 110.400 104.980 ;
        RECT 112.010 104.920 112.330 104.980 ;
        RECT 114.785 104.935 115.075 104.980 ;
        RECT 127.650 105.120 127.970 105.180 ;
        RECT 128.125 105.120 128.415 105.165 ;
        RECT 127.650 104.980 128.415 105.120 ;
        RECT 127.650 104.920 127.970 104.980 ;
        RECT 128.125 104.935 128.415 104.980 ;
        RECT 129.045 105.120 129.335 105.165 ;
        RECT 144.210 105.120 144.530 105.180 ;
        RECT 129.045 104.980 144.530 105.120 ;
        RECT 129.045 104.935 129.335 104.980 ;
        RECT 101.445 104.595 101.735 104.825 ;
        RECT 110.185 104.595 110.475 104.825 ;
        RECT 97.750 104.440 98.070 104.500 ;
        RECT 93.700 104.300 98.070 104.440 ;
        RECT 80.360 104.145 80.500 104.300 ;
        RECT 82.570 104.240 82.890 104.300 ;
        RECT 92.690 104.240 93.010 104.300 ;
        RECT 97.750 104.240 98.070 104.300 ;
        RECT 98.210 104.240 98.530 104.500 ;
        RECT 80.285 103.915 80.575 104.145 ;
        RECT 97.840 104.100 97.980 104.240 ;
        RECT 101.520 104.100 101.660 104.595 ;
        RECT 110.630 104.580 110.950 104.840 ;
        RECT 111.565 104.780 111.855 104.825 ;
        RECT 111.565 104.640 113.160 104.780 ;
        RECT 111.565 104.595 111.855 104.640 ;
        RECT 104.215 104.440 104.505 104.485 ;
        RECT 106.735 104.440 107.025 104.485 ;
        RECT 107.925 104.440 108.215 104.485 ;
        RECT 104.215 104.300 108.215 104.440 ;
        RECT 104.215 104.255 104.505 104.300 ;
        RECT 106.735 104.255 107.025 104.300 ;
        RECT 107.925 104.255 108.215 104.300 ;
        RECT 108.790 104.240 109.110 104.500 ;
        RECT 112.470 104.240 112.790 104.500 ;
        RECT 101.890 104.100 102.210 104.160 ;
        RECT 80.820 103.960 81.880 104.100 ;
        RECT 97.840 103.960 102.210 104.100 ;
        RECT 80.820 103.760 80.960 103.960 ;
        RECT 76.220 103.620 80.960 103.760 ;
        RECT 81.190 103.560 81.510 103.820 ;
        RECT 81.740 103.760 81.880 103.960 ;
        RECT 101.890 103.900 102.210 103.960 ;
        RECT 104.650 104.100 104.940 104.145 ;
        RECT 106.220 104.100 106.510 104.145 ;
        RECT 108.320 104.100 108.610 104.145 ;
        RECT 104.650 103.960 108.610 104.100 ;
        RECT 104.650 103.915 104.940 103.960 ;
        RECT 106.220 103.915 106.510 103.960 ;
        RECT 108.320 103.915 108.610 103.960 ;
        RECT 84.410 103.760 84.730 103.820 ;
        RECT 81.740 103.620 84.730 103.760 ;
        RECT 84.410 103.560 84.730 103.620 ;
        RECT 84.885 103.760 85.175 103.805 ;
        RECT 86.250 103.760 86.570 103.820 ;
        RECT 84.885 103.620 86.570 103.760 ;
        RECT 84.885 103.575 85.175 103.620 ;
        RECT 86.250 103.560 86.570 103.620 ;
        RECT 92.245 103.760 92.535 103.805 ;
        RECT 94.530 103.760 94.850 103.820 ;
        RECT 92.245 103.620 94.850 103.760 ;
        RECT 92.245 103.575 92.535 103.620 ;
        RECT 94.530 103.560 94.850 103.620 ;
        RECT 95.465 103.760 95.755 103.805 ;
        RECT 95.910 103.760 96.230 103.820 ;
        RECT 95.465 103.620 96.230 103.760 ;
        RECT 95.465 103.575 95.755 103.620 ;
        RECT 95.910 103.560 96.230 103.620 ;
        RECT 105.110 103.760 105.430 103.820 ;
        RECT 108.880 103.760 109.020 104.240 ;
        RECT 113.020 104.145 113.160 104.640 ;
        RECT 120.290 104.580 120.610 104.840 ;
        RECT 131.330 104.780 131.650 104.840 ;
        RECT 131.805 104.780 132.095 104.825 ;
        RECT 131.330 104.640 132.095 104.780 ;
        RECT 131.330 104.580 131.650 104.640 ;
        RECT 131.805 104.595 132.095 104.640 ;
        RECT 132.265 104.595 132.555 104.825 ;
        RECT 132.340 104.440 132.480 104.595 ;
        RECT 132.710 104.580 133.030 104.840 ;
        RECT 133.645 104.780 133.935 104.825 ;
        RECT 134.090 104.780 134.410 104.840 ;
        RECT 133.645 104.640 134.410 104.780 ;
        RECT 133.645 104.595 133.935 104.640 ;
        RECT 134.090 104.580 134.410 104.640 ;
        RECT 135.010 104.580 135.330 104.840 ;
        RECT 135.485 104.595 135.775 104.825 ;
        RECT 135.945 104.780 136.235 104.825 ;
        RECT 136.850 104.780 137.170 104.840 ;
        RECT 135.945 104.640 139.380 104.780 ;
        RECT 135.945 104.595 136.235 104.640 ;
        RECT 135.560 104.440 135.700 104.595 ;
        RECT 136.850 104.580 137.170 104.640 ;
        RECT 132.340 104.300 135.700 104.440 ;
        RECT 112.945 103.915 113.235 104.145 ;
        RECT 135.560 104.100 135.700 104.300 ;
        RECT 137.325 104.440 137.615 104.485 ;
        RECT 137.785 104.440 138.075 104.485 ;
        RECT 137.325 104.300 138.075 104.440 ;
        RECT 139.240 104.440 139.380 104.640 ;
        RECT 141.450 104.580 141.770 104.840 ;
        RECT 142.370 104.580 142.690 104.840 ;
        RECT 142.830 104.580 143.150 104.840 ;
        RECT 143.380 104.825 143.520 104.980 ;
        RECT 144.210 104.920 144.530 104.980 ;
        RECT 143.305 104.595 143.595 104.825 ;
        RECT 144.760 104.780 144.900 105.320 ;
        RECT 149.820 105.320 150.970 105.460 ;
        RECT 145.590 105.120 145.910 105.180 ;
        RECT 149.820 105.165 149.960 105.320 ;
        RECT 150.650 105.260 150.970 105.320 ;
        RECT 152.030 105.260 152.350 105.520 ;
        RECT 148.825 105.120 149.115 105.165 ;
        RECT 145.590 104.980 149.115 105.120 ;
        RECT 145.590 104.920 145.910 104.980 ;
        RECT 148.825 104.935 149.115 104.980 ;
        RECT 149.745 104.935 150.035 105.165 ;
        RECT 150.665 104.780 150.955 104.825 ;
        RECT 144.760 104.640 150.955 104.780 ;
        RECT 150.665 104.595 150.955 104.640 ;
        RECT 154.790 104.580 155.110 104.840 ;
        RECT 145.145 104.440 145.435 104.485 ;
        RECT 139.240 104.300 145.435 104.440 ;
        RECT 137.325 104.255 137.615 104.300 ;
        RECT 137.785 104.255 138.075 104.300 ;
        RECT 145.145 104.255 145.435 104.300 ;
        RECT 145.590 104.440 145.910 104.500 ;
        RECT 147.905 104.440 148.195 104.485 ;
        RECT 145.590 104.300 148.195 104.440 ;
        RECT 145.590 104.240 145.910 104.300 ;
        RECT 147.905 104.255 148.195 104.300 ;
        RECT 139.150 104.100 139.470 104.160 ;
        RECT 142.830 104.100 143.150 104.160 ;
        RECT 135.560 103.960 143.150 104.100 ;
        RECT 139.150 103.900 139.470 103.960 ;
        RECT 142.830 103.900 143.150 103.960 ;
        RECT 144.685 104.100 144.975 104.145 ;
        RECT 150.190 104.100 150.510 104.160 ;
        RECT 144.685 103.960 150.510 104.100 ;
        RECT 144.685 103.915 144.975 103.960 ;
        RECT 150.190 103.900 150.510 103.960 ;
        RECT 105.110 103.620 109.020 103.760 ;
        RECT 113.865 103.760 114.155 103.805 ;
        RECT 117.085 103.760 117.375 103.805 ;
        RECT 113.865 103.620 117.375 103.760 ;
        RECT 105.110 103.560 105.430 103.620 ;
        RECT 113.865 103.575 114.155 103.620 ;
        RECT 117.085 103.575 117.375 103.620 ;
        RECT 130.410 103.560 130.730 103.820 ;
        RECT 138.690 103.760 139.010 103.820 ;
        RECT 141.005 103.760 141.295 103.805 ;
        RECT 138.690 103.620 141.295 103.760 ;
        RECT 138.690 103.560 139.010 103.620 ;
        RECT 141.005 103.575 141.295 103.620 ;
        RECT 22.700 102.940 157.020 103.420 ;
        RECT 36.125 102.740 36.415 102.785 ;
        RECT 36.570 102.740 36.890 102.800 ;
        RECT 36.125 102.600 36.890 102.740 ;
        RECT 36.125 102.555 36.415 102.600 ;
        RECT 36.570 102.540 36.890 102.600 ;
        RECT 44.390 102.540 44.710 102.800 ;
        RECT 57.730 102.740 58.050 102.800 ;
        RECT 58.205 102.740 58.495 102.785 ;
        RECT 57.730 102.600 58.495 102.740 ;
        RECT 57.730 102.540 58.050 102.600 ;
        RECT 58.205 102.555 58.495 102.600 ;
        RECT 82.110 102.740 82.430 102.800 ;
        RECT 85.790 102.740 86.110 102.800 ;
        RECT 93.150 102.740 93.470 102.800 ;
        RECT 82.110 102.600 86.110 102.740 ;
        RECT 82.110 102.540 82.430 102.600 ;
        RECT 85.790 102.540 86.110 102.600 ;
        RECT 87.720 102.600 93.470 102.740 ;
        RECT 34.730 102.200 35.050 102.460 ;
        RECT 52.210 102.400 52.500 102.445 ;
        RECT 53.780 102.400 54.070 102.445 ;
        RECT 55.880 102.400 56.170 102.445 ;
        RECT 52.210 102.260 56.170 102.400 ;
        RECT 52.210 102.215 52.500 102.260 ;
        RECT 53.780 102.215 54.070 102.260 ;
        RECT 55.880 102.215 56.170 102.260 ;
        RECT 58.650 102.400 58.970 102.460 ;
        RECT 80.270 102.400 80.590 102.460 ;
        RECT 58.650 102.260 80.590 102.400 ;
        RECT 58.650 102.200 58.970 102.260 ;
        RECT 80.270 102.200 80.590 102.260 ;
        RECT 80.730 102.400 81.050 102.460 ;
        RECT 87.720 102.400 87.860 102.600 ;
        RECT 93.150 102.540 93.470 102.600 ;
        RECT 95.910 102.540 96.230 102.800 ;
        RECT 96.830 102.740 97.150 102.800 ;
        RECT 111.090 102.740 111.410 102.800 ;
        RECT 96.830 102.600 111.410 102.740 ;
        RECT 96.830 102.540 97.150 102.600 ;
        RECT 111.090 102.540 111.410 102.600 ;
        RECT 131.330 102.740 131.650 102.800 ;
        RECT 132.265 102.740 132.555 102.785 ;
        RECT 131.330 102.600 132.555 102.740 ;
        RECT 131.330 102.540 131.650 102.600 ;
        RECT 132.265 102.555 132.555 102.600 ;
        RECT 138.230 102.540 138.550 102.800 ;
        RECT 145.590 102.740 145.910 102.800 ;
        RECT 143.840 102.600 145.910 102.740 ;
        RECT 80.730 102.260 87.860 102.400 ;
        RECT 88.130 102.400 88.420 102.445 ;
        RECT 90.230 102.400 90.520 102.445 ;
        RECT 91.800 102.400 92.090 102.445 ;
        RECT 88.130 102.260 92.090 102.400 ;
        RECT 80.730 102.200 81.050 102.260 ;
        RECT 88.130 102.215 88.420 102.260 ;
        RECT 90.230 102.215 90.520 102.260 ;
        RECT 91.800 102.215 92.090 102.260 ;
        RECT 94.545 102.400 94.835 102.445 ;
        RECT 98.210 102.400 98.530 102.460 ;
        RECT 118.450 102.400 118.740 102.445 ;
        RECT 120.020 102.400 120.310 102.445 ;
        RECT 122.120 102.400 122.410 102.445 ;
        RECT 94.545 102.260 102.580 102.400 ;
        RECT 94.545 102.215 94.835 102.260 ;
        RECT 98.210 102.200 98.530 102.260 ;
        RECT 32.905 102.060 33.195 102.105 ;
        RECT 33.350 102.060 33.670 102.120 ;
        RECT 32.905 101.920 33.670 102.060 ;
        RECT 32.905 101.875 33.195 101.920 ;
        RECT 33.350 101.860 33.670 101.920 ;
        RECT 35.205 101.875 35.495 102.105 ;
        RECT 51.775 102.060 52.065 102.105 ;
        RECT 54.295 102.060 54.585 102.105 ;
        RECT 55.485 102.060 55.775 102.105 ;
        RECT 51.775 101.920 55.775 102.060 ;
        RECT 51.775 101.875 52.065 101.920 ;
        RECT 54.295 101.875 54.585 101.920 ;
        RECT 55.485 101.875 55.775 101.920 ;
        RECT 56.365 102.060 56.655 102.105 ;
        RECT 66.930 102.060 67.250 102.120 ;
        RECT 75.210 102.060 75.530 102.120 ;
        RECT 81.650 102.060 81.970 102.120 ;
        RECT 85.330 102.060 85.650 102.120 ;
        RECT 56.365 101.920 67.250 102.060 ;
        RECT 56.365 101.875 56.655 101.920 ;
        RECT 30.605 101.720 30.895 101.765 ;
        RECT 31.510 101.720 31.830 101.780 ;
        RECT 30.605 101.580 31.830 101.720 ;
        RECT 30.605 101.535 30.895 101.580 ;
        RECT 31.510 101.520 31.830 101.580 ;
        RECT 32.430 101.720 32.750 101.780 ;
        RECT 34.270 101.720 34.590 101.780 ;
        RECT 32.430 101.580 34.590 101.720 ;
        RECT 35.280 101.720 35.420 101.875 ;
        RECT 66.930 101.860 67.250 101.920 ;
        RECT 67.480 101.920 68.540 102.060 ;
        RECT 37.045 101.720 37.335 101.765 ;
        RECT 35.280 101.580 37.335 101.720 ;
        RECT 32.430 101.520 32.750 101.580 ;
        RECT 34.270 101.520 34.590 101.580 ;
        RECT 37.045 101.535 37.335 101.580 ;
        RECT 37.950 101.720 38.270 101.780 ;
        RECT 39.805 101.720 40.095 101.765 ;
        RECT 37.950 101.580 40.095 101.720 ;
        RECT 37.950 101.520 38.270 101.580 ;
        RECT 39.805 101.535 40.095 101.580 ;
        RECT 40.725 101.720 41.015 101.765 ;
        RECT 41.185 101.720 41.475 101.765 ;
        RECT 40.725 101.580 41.475 101.720 ;
        RECT 40.725 101.535 41.015 101.580 ;
        RECT 41.185 101.535 41.475 101.580 ;
        RECT 43.025 101.720 43.315 101.765 ;
        RECT 43.930 101.720 44.250 101.780 ;
        RECT 43.025 101.580 44.250 101.720 ;
        RECT 43.025 101.535 43.315 101.580 ;
        RECT 43.930 101.520 44.250 101.580 ;
        RECT 45.310 101.520 45.630 101.780 ;
        RECT 59.110 101.520 59.430 101.780 ;
        RECT 59.585 101.720 59.875 101.765 ;
        RECT 59.585 101.580 60.260 101.720 ;
        RECT 59.585 101.535 59.875 101.580 ;
        RECT 29.670 101.180 29.990 101.440 ;
        RECT 33.810 101.380 34.130 101.440 ;
        RECT 40.265 101.380 40.555 101.425 ;
        RECT 33.810 101.240 40.555 101.380 ;
        RECT 33.810 101.180 34.130 101.240 ;
        RECT 40.265 101.195 40.555 101.240 ;
        RECT 42.105 101.195 42.395 101.425 ;
        RECT 54.510 101.380 54.830 101.440 ;
        RECT 55.030 101.380 55.320 101.425 ;
        RECT 54.510 101.240 55.320 101.380 ;
        RECT 31.525 101.040 31.815 101.085 ;
        RECT 34.730 101.040 35.050 101.100 ;
        RECT 31.525 100.900 35.050 101.040 ;
        RECT 31.525 100.855 31.815 100.900 ;
        RECT 34.730 100.840 35.050 100.900 ;
        RECT 37.030 101.040 37.350 101.100 ;
        RECT 42.180 101.040 42.320 101.195 ;
        RECT 54.510 101.180 54.830 101.240 ;
        RECT 55.030 101.195 55.320 101.240 ;
        RECT 37.030 100.900 42.320 101.040 ;
        RECT 49.465 101.040 49.755 101.085 ;
        RECT 57.270 101.040 57.590 101.100 ;
        RECT 49.465 100.900 57.590 101.040 ;
        RECT 60.120 101.040 60.260 101.580 ;
        RECT 60.505 101.535 60.795 101.765 ;
        RECT 60.965 101.720 61.255 101.765 ;
        RECT 63.710 101.720 64.030 101.780 ;
        RECT 60.965 101.580 64.030 101.720 ;
        RECT 60.965 101.535 61.255 101.580 ;
        RECT 60.580 101.380 60.720 101.535 ;
        RECT 63.710 101.520 64.030 101.580 ;
        RECT 65.105 101.535 65.395 101.765 ;
        RECT 65.550 101.720 65.870 101.780 ;
        RECT 66.025 101.720 66.315 101.765 ;
        RECT 67.480 101.720 67.620 101.920 ;
        RECT 65.550 101.580 67.620 101.720 ;
        RECT 65.180 101.380 65.320 101.535 ;
        RECT 65.550 101.520 65.870 101.580 ;
        RECT 66.025 101.535 66.315 101.580 ;
        RECT 67.850 101.520 68.170 101.780 ;
        RECT 68.400 101.765 68.540 101.920 ;
        RECT 75.210 101.920 81.970 102.060 ;
        RECT 75.210 101.860 75.530 101.920 ;
        RECT 68.325 101.535 68.615 101.765 ;
        RECT 69.245 101.720 69.535 101.765 ;
        RECT 71.530 101.720 71.850 101.780 ;
        RECT 69.245 101.580 71.850 101.720 ;
        RECT 69.245 101.535 69.535 101.580 ;
        RECT 71.530 101.520 71.850 101.580 ;
        RECT 68.785 101.380 69.075 101.425 ;
        RECT 60.580 101.240 69.075 101.380 ;
        RECT 68.785 101.195 69.075 101.240 ;
        RECT 63.250 101.040 63.570 101.100 ;
        RECT 60.120 100.900 63.570 101.040 ;
        RECT 37.030 100.840 37.350 100.900 ;
        RECT 49.465 100.855 49.755 100.900 ;
        RECT 57.270 100.840 57.590 100.900 ;
        RECT 63.250 100.840 63.570 100.900 ;
        RECT 64.185 101.040 64.475 101.085 ;
        RECT 64.630 101.040 64.950 101.100 ;
        RECT 64.185 100.900 64.950 101.040 ;
        RECT 64.185 100.855 64.475 100.900 ;
        RECT 64.630 100.840 64.950 100.900 ;
        RECT 76.590 100.840 76.910 101.100 ;
        RECT 77.140 101.040 77.280 101.920 ;
        RECT 81.650 101.860 81.970 101.920 ;
        RECT 82.660 101.920 85.650 102.060 ;
        RECT 77.525 101.720 77.815 101.765 ;
        RECT 78.430 101.720 78.750 101.780 ;
        RECT 77.525 101.580 78.750 101.720 ;
        RECT 77.525 101.535 77.815 101.580 ;
        RECT 78.430 101.520 78.750 101.580 ;
        RECT 78.905 101.720 79.195 101.765 ;
        RECT 79.810 101.720 80.130 101.780 ;
        RECT 78.905 101.580 80.130 101.720 ;
        RECT 78.905 101.535 79.195 101.580 ;
        RECT 79.810 101.520 80.130 101.580 ;
        RECT 80.730 101.520 81.050 101.780 ;
        RECT 81.205 101.535 81.495 101.765 ;
        RECT 81.280 101.380 81.420 101.535 ;
        RECT 82.110 101.520 82.430 101.780 ;
        RECT 82.660 101.765 82.800 101.920 ;
        RECT 85.330 101.860 85.650 101.920 ;
        RECT 88.525 102.060 88.815 102.105 ;
        RECT 89.715 102.060 90.005 102.105 ;
        RECT 92.235 102.060 92.525 102.105 ;
        RECT 88.525 101.920 92.525 102.060 ;
        RECT 88.525 101.875 88.815 101.920 ;
        RECT 89.715 101.875 90.005 101.920 ;
        RECT 92.235 101.875 92.525 101.920 ;
        RECT 97.750 102.060 98.070 102.120 ;
        RECT 97.750 101.920 99.360 102.060 ;
        RECT 97.750 101.860 98.070 101.920 ;
        RECT 82.585 101.535 82.875 101.765 ;
        RECT 84.410 101.520 84.730 101.780 ;
        RECT 84.870 101.520 85.190 101.780 ;
        RECT 85.790 101.520 86.110 101.780 ;
        RECT 86.250 101.520 86.570 101.780 ;
        RECT 87.645 101.720 87.935 101.765 ;
        RECT 88.090 101.720 88.410 101.780 ;
        RECT 99.220 101.765 99.360 101.920 ;
        RECT 101.430 101.860 101.750 102.120 ;
        RECT 98.685 101.720 98.975 101.765 ;
        RECT 87.645 101.580 88.410 101.720 ;
        RECT 87.645 101.535 87.935 101.580 ;
        RECT 88.090 101.520 88.410 101.580 ;
        RECT 88.640 101.580 98.975 101.720 ;
        RECT 84.500 101.380 84.640 101.520 ;
        RECT 88.640 101.380 88.780 101.580 ;
        RECT 98.685 101.535 98.975 101.580 ;
        RECT 99.145 101.535 99.435 101.765 ;
        RECT 99.590 101.720 99.910 101.780 ;
        RECT 100.065 101.720 100.355 101.765 ;
        RECT 99.590 101.580 100.355 101.720 ;
        RECT 99.590 101.520 99.910 101.580 ;
        RECT 100.065 101.535 100.355 101.580 ;
        RECT 100.525 101.535 100.815 101.765 ;
        RECT 100.985 101.720 101.275 101.765 ;
        RECT 101.520 101.720 101.660 101.860 ;
        RECT 100.985 101.580 101.660 101.720 ;
        RECT 100.985 101.535 101.275 101.580 ;
        RECT 81.280 101.240 84.180 101.380 ;
        RECT 84.500 101.240 88.780 101.380 ;
        RECT 84.040 101.100 84.180 101.240 ;
        RECT 88.980 101.195 89.270 101.425 ;
        RECT 91.770 101.380 92.090 101.440 ;
        RECT 95.765 101.380 96.055 101.425 ;
        RECT 91.770 101.240 96.055 101.380 ;
        RECT 78.445 101.040 78.735 101.085 ;
        RECT 77.140 100.900 78.735 101.040 ;
        RECT 78.445 100.855 78.735 100.900 ;
        RECT 79.810 100.840 80.130 101.100 ;
        RECT 83.490 100.840 83.810 101.100 ;
        RECT 83.950 101.040 84.270 101.100 ;
        RECT 84.870 101.040 85.190 101.100 ;
        RECT 83.950 100.900 85.190 101.040 ;
        RECT 83.950 100.840 84.270 100.900 ;
        RECT 84.870 100.840 85.190 100.900 ;
        RECT 87.630 101.040 87.950 101.100 ;
        RECT 89.055 101.040 89.195 101.195 ;
        RECT 91.770 101.180 92.090 101.240 ;
        RECT 95.765 101.195 96.055 101.240 ;
        RECT 96.830 101.180 97.150 101.440 ;
        RECT 100.600 101.380 100.740 101.535 ;
        RECT 101.890 101.520 102.210 101.780 ;
        RECT 102.440 101.765 102.580 102.260 ;
        RECT 118.450 102.260 122.410 102.400 ;
        RECT 118.450 102.215 118.740 102.260 ;
        RECT 120.020 102.215 120.310 102.260 ;
        RECT 122.120 102.215 122.410 102.260 ;
        RECT 125.390 102.400 125.680 102.445 ;
        RECT 127.490 102.400 127.780 102.445 ;
        RECT 129.060 102.400 129.350 102.445 ;
        RECT 125.390 102.260 129.350 102.400 ;
        RECT 125.390 102.215 125.680 102.260 ;
        RECT 127.490 102.215 127.780 102.260 ;
        RECT 129.060 102.215 129.350 102.260 ;
        RECT 131.790 102.400 132.110 102.460 ;
        RECT 143.840 102.400 143.980 102.600 ;
        RECT 145.590 102.540 145.910 102.600 ;
        RECT 147.430 102.540 147.750 102.800 ;
        RECT 131.790 102.260 135.240 102.400 ;
        RECT 131.790 102.200 132.110 102.260 ;
        RECT 135.100 102.105 135.240 102.260 ;
        RECT 136.940 102.260 143.980 102.400 ;
        RECT 148.850 102.400 149.140 102.445 ;
        RECT 150.950 102.400 151.240 102.445 ;
        RECT 152.520 102.400 152.810 102.445 ;
        RECT 148.850 102.260 152.810 102.400 ;
        RECT 118.015 102.060 118.305 102.105 ;
        RECT 120.535 102.060 120.825 102.105 ;
        RECT 121.725 102.060 122.015 102.105 ;
        RECT 118.015 101.920 122.015 102.060 ;
        RECT 118.015 101.875 118.305 101.920 ;
        RECT 120.535 101.875 120.825 101.920 ;
        RECT 121.725 101.875 122.015 101.920 ;
        RECT 125.785 102.060 126.075 102.105 ;
        RECT 126.975 102.060 127.265 102.105 ;
        RECT 129.495 102.060 129.785 102.105 ;
        RECT 125.785 101.920 129.785 102.060 ;
        RECT 125.785 101.875 126.075 101.920 ;
        RECT 126.975 101.875 127.265 101.920 ;
        RECT 129.495 101.875 129.785 101.920 ;
        RECT 135.025 101.875 135.315 102.105 ;
        RECT 102.365 101.535 102.655 101.765 ;
        RECT 103.285 101.535 103.575 101.765 ;
        RECT 101.445 101.380 101.735 101.425 ;
        RECT 100.600 101.240 101.735 101.380 ;
        RECT 101.980 101.380 102.120 101.520 ;
        RECT 103.360 101.380 103.500 101.535 ;
        RECT 113.390 101.520 113.710 101.780 ;
        RECT 114.325 101.720 114.615 101.765 ;
        RECT 117.530 101.720 117.850 101.780 ;
        RECT 114.325 101.580 117.850 101.720 ;
        RECT 114.325 101.535 114.615 101.580 ;
        RECT 117.530 101.520 117.850 101.580 ;
        RECT 122.605 101.720 122.895 101.765 ;
        RECT 124.890 101.720 125.210 101.780 ;
        RECT 122.605 101.580 125.210 101.720 ;
        RECT 122.605 101.535 122.895 101.580 ;
        RECT 124.890 101.520 125.210 101.580 ;
        RECT 126.240 101.720 126.530 101.765 ;
        RECT 130.410 101.720 130.730 101.780 ;
        RECT 126.240 101.580 130.730 101.720 ;
        RECT 126.240 101.535 126.530 101.580 ;
        RECT 130.410 101.520 130.730 101.580 ;
        RECT 133.170 101.720 133.490 101.780 ;
        RECT 136.940 101.765 137.080 102.260 ;
        RECT 148.850 102.215 149.140 102.260 ;
        RECT 150.950 102.215 151.240 102.260 ;
        RECT 152.520 102.215 152.810 102.260 ;
        RECT 155.250 102.200 155.570 102.460 ;
        RECT 137.770 101.860 138.090 102.120 ;
        RECT 140.530 102.060 140.850 102.120 ;
        RECT 141.450 102.060 141.770 102.120 ;
        RECT 149.245 102.060 149.535 102.105 ;
        RECT 150.435 102.060 150.725 102.105 ;
        RECT 152.955 102.060 153.245 102.105 ;
        RECT 140.530 101.920 149.040 102.060 ;
        RECT 140.530 101.860 140.850 101.920 ;
        RECT 141.450 101.860 141.770 101.920 ;
        RECT 136.865 101.720 137.155 101.765 ;
        RECT 139.165 101.720 139.455 101.765 ;
        RECT 133.170 101.580 137.155 101.720 ;
        RECT 133.170 101.520 133.490 101.580 ;
        RECT 136.865 101.535 137.155 101.580 ;
        RECT 137.860 101.580 139.455 101.720 ;
        RECT 101.980 101.240 103.500 101.380 ;
        RECT 104.650 101.380 104.970 101.440 ;
        RECT 119.830 101.380 120.150 101.440 ;
        RECT 121.270 101.380 121.560 101.425 ;
        RECT 104.650 101.240 118.680 101.380 ;
        RECT 101.445 101.195 101.735 101.240 ;
        RECT 104.650 101.180 104.970 101.240 ;
        RECT 87.630 100.900 89.195 101.040 ;
        RECT 87.630 100.840 87.950 100.900 ;
        RECT 94.990 100.840 95.310 101.100 ;
        RECT 97.765 101.040 98.055 101.085 ;
        RECT 98.670 101.040 98.990 101.100 ;
        RECT 97.765 100.900 98.990 101.040 ;
        RECT 97.765 100.855 98.055 100.900 ;
        RECT 98.670 100.840 98.990 100.900 ;
        RECT 99.590 101.040 99.910 101.100 ;
        RECT 102.825 101.040 103.115 101.085 ;
        RECT 99.590 100.900 103.115 101.040 ;
        RECT 99.590 100.840 99.910 100.900 ;
        RECT 102.825 100.855 103.115 100.900 ;
        RECT 113.850 100.840 114.170 101.100 ;
        RECT 115.705 101.040 115.995 101.085 ;
        RECT 117.990 101.040 118.310 101.100 ;
        RECT 115.705 100.900 118.310 101.040 ;
        RECT 118.540 101.040 118.680 101.240 ;
        RECT 119.830 101.240 121.560 101.380 ;
        RECT 119.830 101.180 120.150 101.240 ;
        RECT 121.270 101.195 121.560 101.240 ;
        RECT 129.490 101.380 129.810 101.440 ;
        RECT 137.860 101.380 138.000 101.580 ;
        RECT 139.165 101.535 139.455 101.580 ;
        RECT 142.845 101.720 143.135 101.765 ;
        RECT 143.290 101.720 143.610 101.780 ;
        RECT 144.300 101.765 144.440 101.920 ;
        RECT 142.845 101.580 143.610 101.720 ;
        RECT 142.845 101.535 143.135 101.580 ;
        RECT 143.290 101.520 143.610 101.580 ;
        RECT 144.225 101.535 144.515 101.765 ;
        RECT 145.130 101.520 145.450 101.780 ;
        RECT 145.590 101.520 145.910 101.780 ;
        RECT 146.050 101.520 146.370 101.780 ;
        RECT 147.890 101.720 148.210 101.780 ;
        RECT 148.365 101.720 148.655 101.765 ;
        RECT 147.890 101.580 148.655 101.720 ;
        RECT 148.900 101.720 149.040 101.920 ;
        RECT 149.245 101.920 153.245 102.060 ;
        RECT 149.245 101.875 149.535 101.920 ;
        RECT 150.435 101.875 150.725 101.920 ;
        RECT 152.955 101.875 153.245 101.920 ;
        RECT 151.110 101.720 151.430 101.780 ;
        RECT 148.900 101.580 151.430 101.720 ;
        RECT 147.890 101.520 148.210 101.580 ;
        RECT 148.365 101.535 148.655 101.580 ;
        RECT 151.110 101.520 151.430 101.580 ;
        RECT 129.490 101.240 138.000 101.380 ;
        RECT 138.245 101.380 138.535 101.425 ;
        RECT 144.670 101.380 144.990 101.440 ;
        RECT 147.980 101.380 148.120 101.520 ;
        RECT 138.245 101.240 144.990 101.380 ;
        RECT 129.490 101.180 129.810 101.240 ;
        RECT 138.245 101.195 138.535 101.240 ;
        RECT 144.670 101.180 144.990 101.240 ;
        RECT 145.220 101.240 148.120 101.380 ;
        RECT 148.810 101.380 149.130 101.440 ;
        RECT 149.590 101.380 149.880 101.425 ;
        RECT 148.810 101.240 149.880 101.380 ;
        RECT 126.730 101.040 127.050 101.100 ;
        RECT 118.540 100.900 127.050 101.040 ;
        RECT 115.705 100.855 115.995 100.900 ;
        RECT 117.990 100.840 118.310 100.900 ;
        RECT 126.730 100.840 127.050 100.900 ;
        RECT 130.870 101.040 131.190 101.100 ;
        RECT 135.945 101.040 136.235 101.085 ;
        RECT 130.870 100.900 136.235 101.040 ;
        RECT 130.870 100.840 131.190 100.900 ;
        RECT 135.945 100.855 136.235 100.900 ;
        RECT 143.290 101.040 143.610 101.100 ;
        RECT 145.220 101.040 145.360 101.240 ;
        RECT 148.810 101.180 149.130 101.240 ;
        RECT 149.590 101.195 149.880 101.240 ;
        RECT 143.290 100.900 145.360 101.040 ;
        RECT 145.590 101.040 145.910 101.100 ;
        RECT 150.190 101.040 150.510 101.100 ;
        RECT 145.590 100.900 150.510 101.040 ;
        RECT 143.290 100.840 143.610 100.900 ;
        RECT 145.590 100.840 145.910 100.900 ;
        RECT 150.190 100.840 150.510 100.900 ;
        RECT 22.700 100.220 157.820 100.700 ;
        RECT 26.910 100.020 27.230 100.080 ;
        RECT 40.710 100.020 41.030 100.080 ;
        RECT 24.240 99.880 41.030 100.020 ;
        RECT 24.240 99.385 24.380 99.880 ;
        RECT 26.910 99.820 27.230 99.880 ;
        RECT 40.710 99.820 41.030 99.880 ;
        RECT 58.205 99.835 58.495 100.065 ;
        RECT 80.730 100.020 81.050 100.080 ;
        RECT 63.800 99.880 81.050 100.020 ;
        RECT 33.350 99.725 33.670 99.740 ;
        RECT 33.285 99.495 33.670 99.725 ;
        RECT 33.350 99.480 33.670 99.495 ;
        RECT 34.270 99.480 34.590 99.740 ;
        RECT 37.505 99.680 37.795 99.725 ;
        RECT 36.200 99.540 37.795 99.680 ;
        RECT 58.280 99.680 58.420 99.835 ;
        RECT 63.800 99.680 63.940 99.880 ;
        RECT 80.730 99.820 81.050 99.880 ;
        RECT 87.630 100.020 87.950 100.080 ;
        RECT 89.485 100.020 89.775 100.065 ;
        RECT 87.630 99.880 89.775 100.020 ;
        RECT 87.630 99.820 87.950 99.880 ;
        RECT 89.485 99.835 89.775 99.880 ;
        RECT 90.850 100.020 91.170 100.080 ;
        RECT 117.545 100.020 117.835 100.065 ;
        RECT 90.850 99.880 117.835 100.020 ;
        RECT 90.850 99.820 91.170 99.880 ;
        RECT 117.545 99.835 117.835 99.880 ;
        RECT 119.830 99.820 120.150 100.080 ;
        RECT 133.170 99.820 133.490 100.080 ;
        RECT 142.830 100.020 143.150 100.080 ;
        RECT 145.590 100.020 145.910 100.080 ;
        RECT 142.000 99.880 145.910 100.020 ;
        RECT 74.290 99.680 74.610 99.740 ;
        RECT 58.280 99.540 63.940 99.680 ;
        RECT 25.530 99.385 25.850 99.400 ;
        RECT 24.165 99.155 24.455 99.385 ;
        RECT 25.500 99.155 25.850 99.385 ;
        RECT 25.530 99.140 25.850 99.155 ;
        RECT 31.510 99.340 31.830 99.400 ;
        RECT 35.650 99.340 35.970 99.400 ;
        RECT 36.200 99.340 36.340 99.540 ;
        RECT 37.505 99.495 37.795 99.540 ;
        RECT 31.510 99.200 35.420 99.340 ;
        RECT 31.510 99.140 31.830 99.200 ;
        RECT 25.045 99.000 25.335 99.045 ;
        RECT 26.235 99.000 26.525 99.045 ;
        RECT 28.755 99.000 29.045 99.045 ;
        RECT 25.045 98.860 29.045 99.000 ;
        RECT 25.045 98.815 25.335 98.860 ;
        RECT 26.235 98.815 26.525 98.860 ;
        RECT 28.755 98.815 29.045 98.860 ;
        RECT 29.670 99.000 29.990 99.060 ;
        RECT 29.670 98.860 34.500 99.000 ;
        RECT 29.670 98.800 29.990 98.860 ;
        RECT 24.650 98.660 24.940 98.705 ;
        RECT 26.750 98.660 27.040 98.705 ;
        RECT 28.320 98.660 28.610 98.705 ;
        RECT 24.650 98.520 28.610 98.660 ;
        RECT 24.650 98.475 24.940 98.520 ;
        RECT 26.750 98.475 27.040 98.520 ;
        RECT 28.320 98.475 28.610 98.520 ;
        RECT 30.220 98.320 30.360 98.860 ;
        RECT 30.590 98.660 30.910 98.720 ;
        RECT 33.810 98.660 34.130 98.720 ;
        RECT 30.590 98.520 34.130 98.660 ;
        RECT 34.360 98.660 34.500 98.860 ;
        RECT 34.730 98.800 35.050 99.060 ;
        RECT 35.280 99.000 35.420 99.200 ;
        RECT 35.650 99.200 36.340 99.340 ;
        RECT 35.650 99.140 35.970 99.200 ;
        RECT 37.045 99.155 37.335 99.385 ;
        RECT 37.965 99.155 38.255 99.385 ;
        RECT 56.365 99.340 56.655 99.385 ;
        RECT 57.270 99.340 57.590 99.400 ;
        RECT 60.030 99.340 60.350 99.400 ;
        RECT 63.800 99.385 63.940 99.540 ;
        RECT 71.160 99.540 74.610 99.680 ;
        RECT 56.365 99.200 60.350 99.340 ;
        RECT 56.365 99.155 56.655 99.200 ;
        RECT 37.120 99.000 37.260 99.155 ;
        RECT 35.280 98.860 37.260 99.000 ;
        RECT 38.040 98.660 38.180 99.155 ;
        RECT 57.270 99.140 57.590 99.200 ;
        RECT 60.030 99.140 60.350 99.200 ;
        RECT 63.725 99.155 64.015 99.385 ;
        RECT 64.185 99.155 64.475 99.385 ;
        RECT 54.970 99.000 55.290 99.060 ;
        RECT 55.905 99.000 56.195 99.045 ;
        RECT 54.970 98.860 56.195 99.000 ;
        RECT 54.970 98.800 55.290 98.860 ;
        RECT 55.905 98.815 56.195 98.860 ;
        RECT 63.250 99.000 63.570 99.060 ;
        RECT 64.260 99.000 64.400 99.155 ;
        RECT 65.090 99.140 65.410 99.400 ;
        RECT 65.565 99.340 65.855 99.385 ;
        RECT 66.010 99.340 66.330 99.400 ;
        RECT 71.160 99.385 71.300 99.540 ;
        RECT 74.290 99.480 74.610 99.540 ;
        RECT 76.100 99.680 76.390 99.725 ;
        RECT 76.590 99.680 76.910 99.740 ;
        RECT 94.990 99.680 95.310 99.740 ;
        RECT 76.100 99.540 76.910 99.680 ;
        RECT 76.100 99.495 76.390 99.540 ;
        RECT 76.590 99.480 76.910 99.540 ;
        RECT 90.480 99.540 95.310 99.680 ;
        RECT 65.565 99.200 66.330 99.340 ;
        RECT 65.565 99.155 65.855 99.200 ;
        RECT 66.010 99.140 66.330 99.200 ;
        RECT 71.085 99.155 71.375 99.385 ;
        RECT 71.530 99.340 71.850 99.400 ;
        RECT 72.005 99.340 72.295 99.385 ;
        RECT 71.530 99.200 72.295 99.340 ;
        RECT 71.530 99.140 71.850 99.200 ;
        RECT 72.005 99.155 72.295 99.200 ;
        RECT 83.505 99.155 83.795 99.385 ;
        RECT 63.250 98.860 64.400 99.000 ;
        RECT 66.470 99.000 66.790 99.060 ;
        RECT 74.765 99.000 75.055 99.045 ;
        RECT 66.470 98.860 75.055 99.000 ;
        RECT 63.250 98.800 63.570 98.860 ;
        RECT 66.470 98.800 66.790 98.860 ;
        RECT 74.765 98.815 75.055 98.860 ;
        RECT 75.645 99.000 75.935 99.045 ;
        RECT 76.835 99.000 77.125 99.045 ;
        RECT 79.355 99.000 79.645 99.045 ;
        RECT 75.645 98.860 79.645 99.000 ;
        RECT 75.645 98.815 75.935 98.860 ;
        RECT 76.835 98.815 77.125 98.860 ;
        RECT 79.355 98.815 79.645 98.860 ;
        RECT 34.360 98.520 38.180 98.660 ;
        RECT 59.110 98.660 59.430 98.720 ;
        RECT 67.850 98.660 68.170 98.720 ;
        RECT 75.250 98.660 75.540 98.705 ;
        RECT 77.350 98.660 77.640 98.705 ;
        RECT 78.920 98.660 79.210 98.705 ;
        RECT 83.580 98.660 83.720 99.155 ;
        RECT 83.950 99.140 84.270 99.400 ;
        RECT 84.885 99.155 85.175 99.385 ;
        RECT 84.960 99.000 85.100 99.155 ;
        RECT 85.330 99.140 85.650 99.400 ;
        RECT 90.480 99.385 90.620 99.540 ;
        RECT 94.990 99.480 95.310 99.540 ;
        RECT 96.830 99.680 97.150 99.740 ;
        RECT 101.430 99.680 101.750 99.740 ;
        RECT 96.830 99.540 101.750 99.680 ;
        RECT 96.830 99.480 97.150 99.540 ;
        RECT 101.430 99.480 101.750 99.540 ;
        RECT 113.390 99.680 113.710 99.740 ;
        RECT 117.990 99.680 118.310 99.740 ;
        RECT 124.890 99.680 125.210 99.740 ;
        RECT 126.270 99.680 126.590 99.740 ;
        RECT 129.950 99.680 130.270 99.740 ;
        RECT 113.390 99.540 116.610 99.680 ;
        RECT 113.390 99.480 113.710 99.540 ;
        RECT 90.405 99.155 90.695 99.385 ;
        RECT 90.850 99.340 91.170 99.400 ;
        RECT 91.325 99.340 91.615 99.385 ;
        RECT 90.850 99.200 91.615 99.340 ;
        RECT 90.850 99.140 91.170 99.200 ;
        RECT 91.325 99.155 91.615 99.200 ;
        RECT 91.770 99.140 92.090 99.400 ;
        RECT 97.765 99.155 98.055 99.385 ;
        RECT 85.790 99.000 86.110 99.060 ;
        RECT 97.840 99.000 97.980 99.155 ;
        RECT 98.210 99.140 98.530 99.400 ;
        RECT 99.130 99.140 99.450 99.400 ;
        RECT 99.590 99.140 99.910 99.400 ;
        RECT 106.460 99.340 106.750 99.385 ;
        RECT 107.870 99.340 108.190 99.400 ;
        RECT 106.460 99.200 108.190 99.340 ;
        RECT 116.470 99.340 116.610 99.540 ;
        RECT 117.990 99.540 124.200 99.680 ;
        RECT 117.990 99.480 118.310 99.540 ;
        RECT 117.545 99.340 117.835 99.385 ;
        RECT 116.470 99.200 117.835 99.340 ;
        RECT 106.460 99.155 106.750 99.200 ;
        RECT 107.870 99.140 108.190 99.200 ;
        RECT 117.545 99.155 117.835 99.200 ;
        RECT 120.750 99.140 121.070 99.400 ;
        RECT 122.130 99.140 122.450 99.400 ;
        RECT 124.060 99.385 124.200 99.540 ;
        RECT 124.890 99.540 140.300 99.680 ;
        RECT 124.890 99.480 125.210 99.540 ;
        RECT 126.270 99.480 126.590 99.540 ;
        RECT 129.950 99.480 130.270 99.540 ;
        RECT 123.985 99.155 124.275 99.385 ;
        RECT 126.730 99.340 127.050 99.400 ;
        RECT 128.585 99.340 128.875 99.385 ;
        RECT 129.030 99.340 129.350 99.400 ;
        RECT 126.730 99.200 129.350 99.340 ;
        RECT 126.730 99.140 127.050 99.200 ;
        RECT 128.585 99.155 128.875 99.200 ;
        RECT 129.030 99.140 129.350 99.200 ;
        RECT 138.690 99.385 139.010 99.400 ;
        RECT 138.690 99.340 139.040 99.385 ;
        RECT 138.690 99.200 139.205 99.340 ;
        RECT 138.690 99.155 139.040 99.200 ;
        RECT 138.690 99.140 139.010 99.155 ;
        RECT 84.960 98.860 86.110 99.000 ;
        RECT 85.790 98.800 86.110 98.860 ;
        RECT 92.320 98.860 97.980 99.000 ;
        RECT 98.670 99.000 98.990 99.060 ;
        RECT 103.730 99.000 104.050 99.060 ;
        RECT 98.670 98.860 104.050 99.000 ;
        RECT 59.110 98.520 72.220 98.660 ;
        RECT 30.590 98.460 30.910 98.520 ;
        RECT 33.810 98.460 34.130 98.520 ;
        RECT 59.110 98.460 59.430 98.520 ;
        RECT 67.850 98.460 68.170 98.520 ;
        RECT 31.065 98.320 31.355 98.365 ;
        RECT 30.220 98.180 31.355 98.320 ;
        RECT 31.065 98.135 31.355 98.180 ;
        RECT 32.430 98.120 32.750 98.380 ;
        RECT 32.890 98.320 33.210 98.380 ;
        RECT 33.365 98.320 33.655 98.365 ;
        RECT 32.890 98.180 33.655 98.320 ;
        RECT 32.890 98.120 33.210 98.180 ;
        RECT 33.365 98.135 33.655 98.180 ;
        RECT 35.190 98.320 35.510 98.380 ;
        RECT 36.585 98.320 36.875 98.365 ;
        RECT 35.190 98.180 36.875 98.320 ;
        RECT 35.190 98.120 35.510 98.180 ;
        RECT 36.585 98.135 36.875 98.180 ;
        RECT 61.410 98.320 61.730 98.380 ;
        RECT 62.805 98.320 63.095 98.365 ;
        RECT 61.410 98.180 63.095 98.320 ;
        RECT 61.410 98.120 61.730 98.180 ;
        RECT 62.805 98.135 63.095 98.180 ;
        RECT 71.070 98.320 71.390 98.380 ;
        RECT 71.545 98.320 71.835 98.365 ;
        RECT 71.070 98.180 71.835 98.320 ;
        RECT 72.080 98.320 72.220 98.520 ;
        RECT 75.250 98.520 79.210 98.660 ;
        RECT 75.250 98.475 75.540 98.520 ;
        RECT 77.350 98.475 77.640 98.520 ;
        RECT 78.920 98.475 79.210 98.520 ;
        RECT 79.440 98.520 83.720 98.660 ;
        RECT 79.440 98.320 79.580 98.520 ;
        RECT 72.080 98.180 79.580 98.320 ;
        RECT 71.070 98.120 71.390 98.180 ;
        RECT 71.545 98.135 71.835 98.180 ;
        RECT 81.650 98.120 81.970 98.380 ;
        RECT 82.110 98.320 82.430 98.380 ;
        RECT 82.585 98.320 82.875 98.365 ;
        RECT 82.110 98.180 82.875 98.320 ;
        RECT 83.580 98.320 83.720 98.520 ;
        RECT 92.320 98.320 92.460 98.860 ;
        RECT 98.670 98.800 98.990 98.860 ;
        RECT 103.730 98.800 104.050 98.860 ;
        RECT 105.110 98.800 105.430 99.060 ;
        RECT 106.005 99.000 106.295 99.045 ;
        RECT 107.195 99.000 107.485 99.045 ;
        RECT 109.715 99.000 110.005 99.045 ;
        RECT 115.230 99.000 115.550 99.060 ;
        RECT 115.705 99.000 115.995 99.045 ;
        RECT 106.005 98.860 110.005 99.000 ;
        RECT 106.005 98.815 106.295 98.860 ;
        RECT 107.195 98.815 107.485 98.860 ;
        RECT 109.715 98.815 110.005 98.860 ;
        RECT 112.100 98.860 115.995 99.000 ;
        RECT 112.100 98.705 112.240 98.860 ;
        RECT 115.230 98.800 115.550 98.860 ;
        RECT 115.705 98.815 115.995 98.860 ;
        RECT 116.150 99.000 116.470 99.060 ;
        RECT 116.625 99.000 116.915 99.045 ;
        RECT 116.150 98.860 116.915 99.000 ;
        RECT 116.150 98.800 116.470 98.860 ;
        RECT 116.625 98.815 116.915 98.860 ;
        RECT 117.070 99.000 117.390 99.060 ;
        RECT 119.370 99.000 119.690 99.060 ;
        RECT 117.070 98.860 119.690 99.000 ;
        RECT 117.070 98.800 117.390 98.860 ;
        RECT 119.370 98.800 119.690 98.860 ;
        RECT 120.290 99.000 120.610 99.060 ;
        RECT 140.160 99.045 140.300 99.540 ;
        RECT 140.530 99.140 140.850 99.400 ;
        RECT 141.450 99.140 141.770 99.400 ;
        RECT 142.000 99.385 142.140 99.880 ;
        RECT 142.830 99.820 143.150 99.880 ;
        RECT 145.590 99.820 145.910 99.880 ;
        RECT 147.905 100.020 148.195 100.065 ;
        RECT 148.810 100.020 149.130 100.080 ;
        RECT 147.905 99.880 149.130 100.020 ;
        RECT 147.905 99.835 148.195 99.880 ;
        RECT 148.810 99.820 149.130 99.880 ;
        RECT 149.730 99.820 150.050 100.080 ;
        RECT 144.210 99.680 144.530 99.740 ;
        RECT 142.460 99.540 144.530 99.680 ;
        RECT 142.460 99.385 142.600 99.540 ;
        RECT 144.210 99.480 144.530 99.540 ;
        RECT 146.050 99.680 146.370 99.740 ;
        RECT 149.820 99.680 149.960 99.820 ;
        RECT 152.045 99.680 152.335 99.725 ;
        RECT 146.050 99.540 152.335 99.680 ;
        RECT 146.050 99.480 146.370 99.540 ;
        RECT 152.045 99.495 152.335 99.540 ;
        RECT 141.925 99.155 142.215 99.385 ;
        RECT 142.385 99.155 142.675 99.385 ;
        RECT 149.285 99.155 149.575 99.385 ;
        RECT 149.745 99.155 150.035 99.385 ;
        RECT 150.205 99.340 150.495 99.385 ;
        RECT 150.650 99.340 150.970 99.400 ;
        RECT 150.205 99.200 150.970 99.340 ;
        RECT 150.205 99.155 150.495 99.200 ;
        RECT 121.225 99.000 121.515 99.045 ;
        RECT 123.065 99.000 123.355 99.045 ;
        RECT 120.290 98.860 123.355 99.000 ;
        RECT 120.290 98.800 120.610 98.860 ;
        RECT 121.225 98.815 121.515 98.860 ;
        RECT 123.065 98.815 123.355 98.860 ;
        RECT 124.905 98.815 125.195 99.045 ;
        RECT 135.495 99.000 135.785 99.045 ;
        RECT 138.015 99.000 138.305 99.045 ;
        RECT 139.205 99.000 139.495 99.045 ;
        RECT 135.495 98.860 139.495 99.000 ;
        RECT 135.495 98.815 135.785 98.860 ;
        RECT 138.015 98.815 138.305 98.860 ;
        RECT 139.205 98.815 139.495 98.860 ;
        RECT 140.085 99.000 140.375 99.045 ;
        RECT 143.290 99.000 143.610 99.060 ;
        RECT 140.085 98.860 143.610 99.000 ;
        RECT 140.085 98.815 140.375 98.860 ;
        RECT 105.610 98.660 105.900 98.705 ;
        RECT 107.710 98.660 108.000 98.705 ;
        RECT 109.280 98.660 109.570 98.705 ;
        RECT 105.610 98.520 109.570 98.660 ;
        RECT 105.610 98.475 105.900 98.520 ;
        RECT 107.710 98.475 108.000 98.520 ;
        RECT 109.280 98.475 109.570 98.520 ;
        RECT 112.025 98.475 112.315 98.705 ;
        RECT 121.685 98.660 121.975 98.705 ;
        RECT 123.970 98.660 124.290 98.720 ;
        RECT 121.685 98.520 124.290 98.660 ;
        RECT 121.685 98.475 121.975 98.520 ;
        RECT 123.970 98.460 124.290 98.520 ;
        RECT 83.580 98.180 92.460 98.320 ;
        RECT 96.845 98.320 97.135 98.365 ;
        RECT 104.190 98.320 104.510 98.380 ;
        RECT 96.845 98.180 104.510 98.320 ;
        RECT 82.110 98.120 82.430 98.180 ;
        RECT 82.585 98.135 82.875 98.180 ;
        RECT 96.845 98.135 97.135 98.180 ;
        RECT 104.190 98.120 104.510 98.180 ;
        RECT 112.945 98.320 113.235 98.365 ;
        RECT 114.310 98.320 114.630 98.380 ;
        RECT 112.945 98.180 114.630 98.320 ;
        RECT 112.945 98.135 113.235 98.180 ;
        RECT 114.310 98.120 114.630 98.180 ;
        RECT 119.370 98.320 119.690 98.380 ;
        RECT 124.980 98.320 125.120 98.815 ;
        RECT 143.290 98.800 143.610 98.860 ;
        RECT 143.765 99.000 144.055 99.045 ;
        RECT 144.225 99.000 144.515 99.045 ;
        RECT 149.360 99.000 149.500 99.155 ;
        RECT 143.765 98.860 144.515 99.000 ;
        RECT 143.765 98.815 144.055 98.860 ;
        RECT 144.225 98.815 144.515 98.860 ;
        RECT 148.900 98.860 149.500 99.000 ;
        RECT 149.820 99.000 149.960 99.155 ;
        RECT 150.650 99.140 150.970 99.200 ;
        RECT 151.110 99.140 151.430 99.400 ;
        RECT 154.330 99.340 154.650 99.400 ;
        RECT 154.805 99.340 155.095 99.385 ;
        RECT 154.330 99.200 155.095 99.340 ;
        RECT 154.330 99.140 154.650 99.200 ;
        RECT 154.805 99.155 155.095 99.200 ;
        RECT 149.820 98.860 150.420 99.000 ;
        RECT 135.930 98.660 136.220 98.705 ;
        RECT 137.500 98.660 137.790 98.705 ;
        RECT 139.600 98.660 139.890 98.705 ;
        RECT 135.930 98.520 139.890 98.660 ;
        RECT 135.930 98.475 136.220 98.520 ;
        RECT 137.500 98.475 137.790 98.520 ;
        RECT 139.600 98.475 139.890 98.520 ;
        RECT 119.370 98.180 125.120 98.320 ;
        RECT 129.505 98.320 129.795 98.365 ;
        RECT 140.530 98.320 140.850 98.380 ;
        RECT 129.505 98.180 140.850 98.320 ;
        RECT 119.370 98.120 119.690 98.180 ;
        RECT 129.505 98.135 129.795 98.180 ;
        RECT 140.530 98.120 140.850 98.180 ;
        RECT 144.670 98.320 144.990 98.380 ;
        RECT 147.445 98.320 147.735 98.365 ;
        RECT 144.670 98.180 147.735 98.320 ;
        RECT 148.900 98.320 149.040 98.860 ;
        RECT 150.280 98.720 150.420 98.860 ;
        RECT 150.190 98.460 150.510 98.720 ;
        RECT 152.030 98.320 152.350 98.380 ;
        RECT 148.900 98.180 152.350 98.320 ;
        RECT 144.670 98.120 144.990 98.180 ;
        RECT 147.445 98.135 147.735 98.180 ;
        RECT 152.030 98.120 152.350 98.180 ;
        RECT 22.700 97.500 157.020 97.980 ;
        RECT 25.530 97.100 25.850 97.360 ;
        RECT 30.605 97.300 30.895 97.345 ;
        RECT 32.890 97.300 33.210 97.360 ;
        RECT 30.605 97.160 33.210 97.300 ;
        RECT 30.605 97.115 30.895 97.160 ;
        RECT 32.890 97.100 33.210 97.160 ;
        RECT 33.810 97.100 34.130 97.360 ;
        RECT 36.110 97.300 36.430 97.360 ;
        RECT 43.945 97.300 44.235 97.345 ;
        RECT 45.310 97.300 45.630 97.360 ;
        RECT 75.670 97.300 75.990 97.360 ;
        RECT 36.110 97.160 42.320 97.300 ;
        RECT 36.110 97.100 36.430 97.160 ;
        RECT 31.985 96.960 32.275 97.005 ;
        RECT 35.190 96.960 35.510 97.020 ;
        RECT 31.985 96.820 35.510 96.960 ;
        RECT 31.985 96.775 32.275 96.820 ;
        RECT 35.190 96.760 35.510 96.820 ;
        RECT 37.530 96.960 37.820 97.005 ;
        RECT 39.630 96.960 39.920 97.005 ;
        RECT 41.200 96.960 41.490 97.005 ;
        RECT 37.530 96.820 41.490 96.960 ;
        RECT 37.530 96.775 37.820 96.820 ;
        RECT 39.630 96.775 39.920 96.820 ;
        RECT 41.200 96.775 41.490 96.820 ;
        RECT 32.430 96.620 32.750 96.680 ;
        RECT 26.540 96.480 32.750 96.620 ;
        RECT 26.540 96.325 26.680 96.480 ;
        RECT 32.430 96.420 32.750 96.480 ;
        RECT 37.925 96.620 38.215 96.665 ;
        RECT 39.115 96.620 39.405 96.665 ;
        RECT 41.635 96.620 41.925 96.665 ;
        RECT 37.925 96.480 41.925 96.620 ;
        RECT 42.180 96.620 42.320 97.160 ;
        RECT 43.945 97.160 45.630 97.300 ;
        RECT 43.945 97.115 44.235 97.160 ;
        RECT 45.310 97.100 45.630 97.160 ;
        RECT 72.080 97.160 75.990 97.300 ;
        RECT 44.890 96.960 45.180 97.005 ;
        RECT 46.990 96.960 47.280 97.005 ;
        RECT 48.560 96.960 48.850 97.005 ;
        RECT 44.890 96.820 48.850 96.960 ;
        RECT 44.890 96.775 45.180 96.820 ;
        RECT 46.990 96.775 47.280 96.820 ;
        RECT 48.560 96.775 48.850 96.820 ;
        RECT 51.305 96.960 51.595 97.005 ;
        RECT 52.670 96.960 52.990 97.020 ;
        RECT 51.305 96.820 52.990 96.960 ;
        RECT 51.305 96.775 51.595 96.820 ;
        RECT 52.670 96.760 52.990 96.820 ;
        RECT 62.330 96.960 62.650 97.020 ;
        RECT 72.080 96.960 72.220 97.160 ;
        RECT 75.670 97.100 75.990 97.160 ;
        RECT 78.430 97.100 78.750 97.360 ;
        RECT 79.365 97.300 79.655 97.345 ;
        RECT 80.745 97.300 81.035 97.345 ;
        RECT 79.365 97.160 81.035 97.300 ;
        RECT 79.365 97.115 79.655 97.160 ;
        RECT 80.745 97.115 81.035 97.160 ;
        RECT 84.425 97.300 84.715 97.345 ;
        RECT 85.330 97.300 85.650 97.360 ;
        RECT 84.425 97.160 85.650 97.300 ;
        RECT 84.425 97.115 84.715 97.160 ;
        RECT 85.330 97.100 85.650 97.160 ;
        RECT 90.850 97.100 91.170 97.360 ;
        RECT 107.425 97.300 107.715 97.345 ;
        RECT 107.870 97.300 108.190 97.360 ;
        RECT 95.080 97.160 107.180 97.300 ;
        RECT 62.330 96.820 72.220 96.960 ;
        RECT 72.450 96.960 72.770 97.020 ;
        RECT 88.550 96.960 88.870 97.020 ;
        RECT 95.080 96.960 95.220 97.160 ;
        RECT 72.450 96.820 88.870 96.960 ;
        RECT 62.330 96.760 62.650 96.820 ;
        RECT 65.640 96.665 65.780 96.820 ;
        RECT 72.450 96.760 72.770 96.820 ;
        RECT 88.550 96.760 88.870 96.820 ;
        RECT 89.560 96.820 95.220 96.960 ;
        RECT 95.450 96.960 95.770 97.020 ;
        RECT 97.305 96.960 97.595 97.005 ;
        RECT 95.450 96.820 97.595 96.960 ;
        RECT 45.285 96.620 45.575 96.665 ;
        RECT 46.475 96.620 46.765 96.665 ;
        RECT 48.995 96.620 49.285 96.665 ;
        RECT 42.180 96.480 45.080 96.620 ;
        RECT 37.925 96.435 38.215 96.480 ;
        RECT 39.115 96.435 39.405 96.480 ;
        RECT 41.635 96.435 41.925 96.480 ;
        RECT 26.465 96.095 26.755 96.325 ;
        RECT 29.685 96.095 29.975 96.325 ;
        RECT 29.760 95.940 29.900 96.095 ;
        RECT 30.590 96.080 30.910 96.340 ;
        RECT 32.890 96.280 33.210 96.340 ;
        RECT 33.825 96.280 34.115 96.325 ;
        RECT 31.140 96.140 34.115 96.280 ;
        RECT 31.140 95.940 31.280 96.140 ;
        RECT 32.890 96.080 33.210 96.140 ;
        RECT 33.825 96.095 34.115 96.140 ;
        RECT 35.190 96.080 35.510 96.340 ;
        RECT 37.045 96.280 37.335 96.325 ;
        RECT 40.710 96.280 41.030 96.340 ;
        RECT 44.390 96.280 44.710 96.340 ;
        RECT 37.045 96.140 44.710 96.280 ;
        RECT 44.940 96.280 45.080 96.480 ;
        RECT 45.285 96.480 49.285 96.620 ;
        RECT 45.285 96.435 45.575 96.480 ;
        RECT 46.475 96.435 46.765 96.480 ;
        RECT 48.995 96.435 49.285 96.480 ;
        RECT 65.565 96.435 65.855 96.665 ;
        RECT 66.470 96.620 66.790 96.680 ;
        RECT 76.145 96.620 76.435 96.665 ;
        RECT 88.090 96.620 88.410 96.680 ;
        RECT 66.470 96.480 88.410 96.620 ;
        RECT 66.470 96.420 66.790 96.480 ;
        RECT 76.145 96.435 76.435 96.480 ;
        RECT 88.090 96.420 88.410 96.480 ;
        RECT 54.510 96.280 54.830 96.340 ;
        RECT 55.445 96.280 55.735 96.325 ;
        RECT 44.940 96.140 49.680 96.280 ;
        RECT 37.045 96.095 37.335 96.140 ;
        RECT 40.710 96.080 41.030 96.140 ;
        RECT 44.390 96.080 44.710 96.140 ;
        RECT 33.350 95.940 33.670 96.000 ;
        RECT 29.760 95.800 31.280 95.940 ;
        RECT 32.520 95.800 33.670 95.940 ;
        RECT 32.520 95.645 32.660 95.800 ;
        RECT 33.350 95.740 33.670 95.800 ;
        RECT 38.380 95.940 38.670 95.985 ;
        RECT 41.170 95.940 41.490 96.000 ;
        RECT 38.380 95.800 41.490 95.940 ;
        RECT 38.380 95.755 38.670 95.800 ;
        RECT 41.170 95.740 41.490 95.800 ;
        RECT 45.740 95.940 46.030 95.985 ;
        RECT 48.990 95.940 49.310 96.000 ;
        RECT 45.740 95.800 49.310 95.940 ;
        RECT 49.540 95.940 49.680 96.140 ;
        RECT 54.510 96.140 55.735 96.280 ;
        RECT 54.510 96.080 54.830 96.140 ;
        RECT 55.445 96.095 55.735 96.140 ;
        RECT 67.405 96.095 67.695 96.325 ;
        RECT 67.850 96.280 68.170 96.340 ;
        RECT 68.325 96.280 68.615 96.325 ;
        RECT 67.850 96.140 68.615 96.280 ;
        RECT 66.025 95.940 66.315 95.985 ;
        RECT 49.540 95.800 66.315 95.940 ;
        RECT 67.480 95.940 67.620 96.095 ;
        RECT 67.850 96.080 68.170 96.140 ;
        RECT 68.325 96.095 68.615 96.140 ;
        RECT 69.245 96.280 69.535 96.325 ;
        RECT 72.910 96.280 73.230 96.340 ;
        RECT 81.190 96.280 81.510 96.340 ;
        RECT 69.245 96.140 73.230 96.280 ;
        RECT 69.245 96.095 69.535 96.140 ;
        RECT 72.910 96.080 73.230 96.140 ;
        RECT 75.300 96.140 81.510 96.280 ;
        RECT 71.070 95.940 71.390 96.000 ;
        RECT 67.480 95.800 71.390 95.940 ;
        RECT 45.740 95.755 46.030 95.800 ;
        RECT 48.990 95.740 49.310 95.800 ;
        RECT 66.025 95.755 66.315 95.800 ;
        RECT 71.070 95.740 71.390 95.800 ;
        RECT 71.530 95.940 71.850 96.000 ;
        RECT 72.005 95.940 72.295 95.985 ;
        RECT 71.530 95.800 72.295 95.940 ;
        RECT 71.530 95.740 71.850 95.800 ;
        RECT 72.005 95.755 72.295 95.800 ;
        RECT 72.450 95.740 72.770 96.000 ;
        RECT 32.445 95.415 32.735 95.645 ;
        RECT 54.970 95.600 55.290 95.660 ;
        RECT 56.365 95.600 56.655 95.645 ;
        RECT 54.970 95.460 56.655 95.600 ;
        RECT 54.970 95.400 55.290 95.460 ;
        RECT 56.365 95.415 56.655 95.460 ;
        RECT 60.030 95.600 60.350 95.660 ;
        RECT 75.300 95.600 75.440 96.140 ;
        RECT 75.670 95.940 75.990 96.000 ;
        RECT 79.350 95.985 79.670 96.000 ;
        RECT 80.360 95.985 80.500 96.140 ;
        RECT 81.190 96.080 81.510 96.140 ;
        RECT 81.650 96.280 81.970 96.340 ;
        RECT 83.505 96.280 83.795 96.325 ;
        RECT 84.425 96.280 84.715 96.325 ;
        RECT 81.650 96.140 84.715 96.280 ;
        RECT 81.650 96.080 81.970 96.140 ;
        RECT 83.505 96.095 83.795 96.140 ;
        RECT 84.425 96.095 84.715 96.140 ;
        RECT 84.870 96.280 85.190 96.340 ;
        RECT 85.345 96.280 85.635 96.325 ;
        RECT 84.870 96.140 85.635 96.280 ;
        RECT 84.870 96.080 85.190 96.140 ;
        RECT 85.345 96.095 85.635 96.140 ;
        RECT 75.670 95.800 79.120 95.940 ;
        RECT 75.670 95.740 75.990 95.800 ;
        RECT 60.030 95.460 75.440 95.600 ;
        RECT 78.980 95.600 79.120 95.800 ;
        RECT 79.285 95.755 79.670 95.985 ;
        RECT 80.285 95.755 80.575 95.985 ;
        RECT 89.560 95.940 89.700 96.820 ;
        RECT 95.450 96.760 95.770 96.820 ;
        RECT 97.305 96.775 97.595 96.820 ;
        RECT 93.150 96.620 93.470 96.680 ;
        RECT 104.650 96.620 104.970 96.680 ;
        RECT 90.480 96.480 104.970 96.620 ;
        RECT 80.820 95.800 89.700 95.940 ;
        RECT 89.945 95.940 90.235 95.985 ;
        RECT 90.480 95.940 90.620 96.480 ;
        RECT 93.150 96.420 93.470 96.480 ;
        RECT 104.650 96.420 104.970 96.480 ;
        RECT 94.070 96.280 94.390 96.340 ;
        RECT 94.070 96.140 95.680 96.280 ;
        RECT 94.070 96.080 94.390 96.140 ;
        RECT 91.310 95.985 91.630 96.000 ;
        RECT 95.540 95.985 95.680 96.140 ;
        RECT 96.370 96.080 96.690 96.340 ;
        RECT 96.830 96.290 97.150 96.340 ;
        RECT 96.830 96.150 97.335 96.290 ;
        RECT 96.830 96.080 97.150 96.150 ;
        RECT 97.750 96.080 98.070 96.340 ;
        RECT 102.350 96.080 102.670 96.340 ;
        RECT 89.945 95.800 90.620 95.940 ;
        RECT 79.350 95.740 79.670 95.755 ;
        RECT 80.820 95.600 80.960 95.800 ;
        RECT 89.945 95.755 90.235 95.800 ;
        RECT 91.025 95.755 91.630 95.985 ;
        RECT 94.545 95.755 94.835 95.985 ;
        RECT 95.465 95.755 95.755 95.985 ;
        RECT 107.040 95.940 107.180 97.160 ;
        RECT 107.425 97.160 108.190 97.300 ;
        RECT 107.425 97.115 107.715 97.160 ;
        RECT 107.870 97.100 108.190 97.160 ;
        RECT 113.390 97.300 113.710 97.360 ;
        RECT 113.865 97.300 114.155 97.345 ;
        RECT 113.390 97.160 114.155 97.300 ;
        RECT 113.390 97.100 113.710 97.160 ;
        RECT 113.865 97.115 114.155 97.160 ;
        RECT 117.530 97.100 117.850 97.360 ;
        RECT 122.130 97.300 122.450 97.360 ;
        RECT 122.605 97.300 122.895 97.345 ;
        RECT 122.130 97.160 122.895 97.300 ;
        RECT 122.130 97.100 122.450 97.160 ;
        RECT 122.605 97.115 122.895 97.160 ;
        RECT 132.710 97.300 133.030 97.360 ;
        RECT 135.945 97.300 136.235 97.345 ;
        RECT 132.710 97.160 136.235 97.300 ;
        RECT 132.710 97.100 133.030 97.160 ;
        RECT 135.945 97.115 136.235 97.160 ;
        RECT 109.710 96.960 110.030 97.020 ;
        RECT 110.185 96.960 110.475 97.005 ;
        RECT 116.150 96.960 116.470 97.020 ;
        RECT 109.710 96.820 116.470 96.960 ;
        RECT 109.710 96.760 110.030 96.820 ;
        RECT 110.185 96.775 110.475 96.820 ;
        RECT 116.150 96.760 116.470 96.820 ;
        RECT 141.910 96.960 142.200 97.005 ;
        RECT 143.480 96.960 143.770 97.005 ;
        RECT 145.580 96.960 145.870 97.005 ;
        RECT 141.910 96.820 145.870 96.960 ;
        RECT 141.910 96.775 142.200 96.820 ;
        RECT 143.480 96.775 143.770 96.820 ;
        RECT 145.580 96.775 145.870 96.820 ;
        RECT 148.390 96.960 148.680 97.005 ;
        RECT 150.490 96.960 150.780 97.005 ;
        RECT 152.060 96.960 152.350 97.005 ;
        RECT 148.390 96.820 152.350 96.960 ;
        RECT 148.390 96.775 148.680 96.820 ;
        RECT 150.490 96.775 150.780 96.820 ;
        RECT 152.060 96.775 152.350 96.820 ;
        RECT 109.265 96.435 109.555 96.665 ;
        RECT 117.070 96.620 117.390 96.680 ;
        RECT 111.180 96.480 117.390 96.620 ;
        RECT 108.345 96.280 108.635 96.325 ;
        RECT 109.340 96.280 109.480 96.435 ;
        RECT 108.345 96.140 109.480 96.280 ;
        RECT 108.345 96.095 108.635 96.140 ;
        RECT 111.180 95.940 111.320 96.480 ;
        RECT 117.070 96.420 117.390 96.480 ;
        RECT 118.465 96.620 118.755 96.665 ;
        RECT 120.750 96.620 121.070 96.680 ;
        RECT 140.070 96.620 140.390 96.680 ;
        RECT 118.465 96.480 121.440 96.620 ;
        RECT 118.465 96.435 118.755 96.480 ;
        RECT 120.750 96.420 121.070 96.480 ;
        RECT 113.390 96.080 113.710 96.340 ;
        RECT 114.310 96.080 114.630 96.340 ;
        RECT 115.230 96.280 115.550 96.340 ;
        RECT 115.705 96.280 115.995 96.325 ;
        RECT 115.230 96.140 115.995 96.280 ;
        RECT 115.230 96.080 115.550 96.140 ;
        RECT 115.705 96.095 115.995 96.140 ;
        RECT 107.040 95.800 111.320 95.940 ;
        RECT 91.310 95.740 91.630 95.755 ;
        RECT 78.980 95.460 80.960 95.600 ;
        RECT 60.030 95.400 60.350 95.460 ;
        RECT 91.770 95.400 92.090 95.660 ;
        RECT 93.610 95.600 93.930 95.660 ;
        RECT 94.620 95.600 94.760 95.755 ;
        RECT 111.550 95.740 111.870 96.000 ;
        RECT 113.480 95.940 113.620 96.080 ;
        RECT 116.625 95.940 116.915 95.985 ;
        RECT 113.480 95.800 116.915 95.940 ;
        RECT 117.160 95.940 117.300 96.420 ;
        RECT 117.990 96.080 118.310 96.340 ;
        RECT 118.925 96.280 119.215 96.325 ;
        RECT 119.370 96.280 119.690 96.340 ;
        RECT 118.925 96.140 119.690 96.280 ;
        RECT 118.925 96.095 119.215 96.140 ;
        RECT 119.370 96.080 119.690 96.140 ;
        RECT 120.290 96.080 120.610 96.340 ;
        RECT 121.300 96.325 121.440 96.480 ;
        RECT 127.280 96.480 140.390 96.620 ;
        RECT 121.225 96.095 121.515 96.325 ;
        RECT 122.145 96.280 122.435 96.325 ;
        RECT 123.525 96.280 123.815 96.325 ;
        RECT 122.145 96.140 123.815 96.280 ;
        RECT 122.145 96.095 122.435 96.140 ;
        RECT 123.525 96.095 123.815 96.140 ;
        RECT 123.970 96.080 124.290 96.340 ;
        RECT 127.280 96.325 127.420 96.480 ;
        RECT 140.070 96.420 140.390 96.480 ;
        RECT 141.475 96.620 141.765 96.665 ;
        RECT 143.995 96.620 144.285 96.665 ;
        RECT 145.185 96.620 145.475 96.665 ;
        RECT 141.475 96.480 145.475 96.620 ;
        RECT 141.475 96.435 141.765 96.480 ;
        RECT 143.995 96.435 144.285 96.480 ;
        RECT 145.185 96.435 145.475 96.480 ;
        RECT 148.785 96.620 149.075 96.665 ;
        RECT 149.975 96.620 150.265 96.665 ;
        RECT 152.495 96.620 152.785 96.665 ;
        RECT 148.785 96.480 152.785 96.620 ;
        RECT 148.785 96.435 149.075 96.480 ;
        RECT 149.975 96.435 150.265 96.480 ;
        RECT 152.495 96.435 152.785 96.480 ;
        RECT 127.205 96.095 127.495 96.325 ;
        RECT 127.665 96.280 127.955 96.325 ;
        RECT 128.110 96.280 128.430 96.340 ;
        RECT 127.665 96.140 128.430 96.280 ;
        RECT 127.665 96.095 127.955 96.140 ;
        RECT 128.110 96.080 128.430 96.140 ;
        RECT 128.570 96.080 128.890 96.340 ;
        RECT 136.850 96.080 137.170 96.340 ;
        RECT 141.910 96.280 142.230 96.340 ;
        RECT 137.400 96.140 142.230 96.280 ;
        RECT 122.605 95.940 122.895 95.985 ;
        RECT 117.160 95.800 122.895 95.940 ;
        RECT 116.625 95.755 116.915 95.800 ;
        RECT 122.605 95.755 122.895 95.800 ;
        RECT 129.030 95.940 129.350 96.000 ;
        RECT 137.400 95.940 137.540 96.140 ;
        RECT 141.910 96.080 142.230 96.140 ;
        RECT 144.670 96.325 144.990 96.340 ;
        RECT 144.670 96.280 145.020 96.325 ;
        RECT 146.065 96.280 146.355 96.325 ;
        RECT 147.890 96.280 148.210 96.340 ;
        RECT 144.670 96.140 145.185 96.280 ;
        RECT 146.065 96.140 148.210 96.280 ;
        RECT 144.670 96.095 145.020 96.140 ;
        RECT 146.065 96.095 146.355 96.140 ;
        RECT 144.670 96.080 144.990 96.095 ;
        RECT 129.030 95.800 137.540 95.940 ;
        RECT 137.770 95.940 138.090 96.000 ;
        RECT 140.530 95.940 140.850 96.000 ;
        RECT 137.770 95.800 140.850 95.940 ;
        RECT 129.030 95.740 129.350 95.800 ;
        RECT 137.770 95.740 138.090 95.800 ;
        RECT 140.530 95.740 140.850 95.800 ;
        RECT 145.130 95.940 145.450 96.000 ;
        RECT 146.140 95.940 146.280 96.095 ;
        RECT 147.890 96.080 148.210 96.140 ;
        RECT 145.130 95.800 146.280 95.940 ;
        RECT 148.350 95.940 148.670 96.000 ;
        RECT 149.130 95.940 149.420 95.985 ;
        RECT 148.350 95.800 149.420 95.940 ;
        RECT 145.130 95.740 145.450 95.800 ;
        RECT 148.350 95.740 148.670 95.800 ;
        RECT 149.130 95.755 149.420 95.800 ;
        RECT 93.610 95.460 94.760 95.600 ;
        RECT 101.445 95.600 101.735 95.645 ;
        RECT 101.890 95.600 102.210 95.660 ;
        RECT 101.445 95.460 102.210 95.600 ;
        RECT 93.610 95.400 93.930 95.460 ;
        RECT 101.445 95.415 101.735 95.460 ;
        RECT 101.890 95.400 102.210 95.460 ;
        RECT 126.730 95.400 127.050 95.660 ;
        RECT 127.650 95.600 127.970 95.660 ;
        RECT 128.125 95.600 128.415 95.645 ;
        RECT 127.650 95.460 128.415 95.600 ;
        RECT 127.650 95.400 127.970 95.460 ;
        RECT 128.125 95.415 128.415 95.460 ;
        RECT 137.310 95.600 137.630 95.660 ;
        RECT 139.165 95.600 139.455 95.645 ;
        RECT 143.750 95.600 144.070 95.660 ;
        RECT 137.310 95.460 144.070 95.600 ;
        RECT 137.310 95.400 137.630 95.460 ;
        RECT 139.165 95.415 139.455 95.460 ;
        RECT 143.750 95.400 144.070 95.460 ;
        RECT 146.510 95.600 146.830 95.660 ;
        RECT 154.330 95.600 154.650 95.660 ;
        RECT 154.805 95.600 155.095 95.645 ;
        RECT 146.510 95.460 155.095 95.600 ;
        RECT 146.510 95.400 146.830 95.460 ;
        RECT 154.330 95.400 154.650 95.460 ;
        RECT 154.805 95.415 155.095 95.460 ;
        RECT 22.700 94.780 157.820 95.260 ;
        RECT 72.450 94.580 72.770 94.640 ;
        RECT 40.800 94.440 72.770 94.580 ;
        RECT 40.800 94.285 40.940 94.440 ;
        RECT 72.450 94.380 72.770 94.440 ;
        RECT 72.910 94.580 73.230 94.640 ;
        RECT 111.550 94.580 111.870 94.640 ;
        RECT 112.945 94.580 113.235 94.625 ;
        RECT 72.910 94.440 74.980 94.580 ;
        RECT 72.910 94.380 73.230 94.440 ;
        RECT 40.725 94.055 41.015 94.285 ;
        RECT 44.390 94.240 44.710 94.300 ;
        RECT 41.260 94.100 50.600 94.240 ;
        RECT 32.445 93.715 32.735 93.945 ;
        RECT 33.365 93.900 33.655 93.945 ;
        RECT 35.650 93.900 35.970 93.960 ;
        RECT 33.365 93.760 35.970 93.900 ;
        RECT 33.365 93.715 33.655 93.760 ;
        RECT 32.520 93.560 32.660 93.715 ;
        RECT 35.650 93.700 35.970 93.760 ;
        RECT 37.045 93.900 37.335 93.945 ;
        RECT 41.260 93.900 41.400 94.100 ;
        RECT 44.390 94.040 44.710 94.100 ;
        RECT 37.045 93.760 41.400 93.900 ;
        RECT 37.045 93.715 37.335 93.760 ;
        RECT 42.090 93.700 42.410 93.960 ;
        RECT 49.910 93.700 50.230 93.960 ;
        RECT 50.460 93.900 50.600 94.100 ;
        RECT 53.130 94.040 53.450 94.300 ;
        RECT 54.970 94.240 55.290 94.300 ;
        RECT 74.840 94.285 74.980 94.440 ;
        RECT 83.580 94.440 109.020 94.580 ;
        RECT 55.750 94.240 56.040 94.285 ;
        RECT 67.250 94.240 67.540 94.285 ;
        RECT 54.970 94.100 56.040 94.240 ;
        RECT 54.970 94.040 55.290 94.100 ;
        RECT 55.750 94.055 56.040 94.100 ;
        RECT 65.180 94.100 67.540 94.240 ;
        RECT 54.525 93.900 54.815 93.945 ;
        RECT 50.460 93.760 54.815 93.900 ;
        RECT 54.525 93.715 54.815 93.760 ;
        RECT 61.885 93.900 62.175 93.945 ;
        RECT 61.885 93.760 63.480 93.900 ;
        RECT 61.885 93.715 62.175 93.760 ;
        RECT 36.110 93.560 36.430 93.620 ;
        RECT 63.340 93.605 63.480 93.760 ;
        RECT 32.520 93.420 36.430 93.560 ;
        RECT 36.110 93.360 36.430 93.420 ;
        RECT 55.405 93.560 55.695 93.605 ;
        RECT 56.595 93.560 56.885 93.605 ;
        RECT 59.115 93.560 59.405 93.605 ;
        RECT 55.405 93.420 59.405 93.560 ;
        RECT 55.405 93.375 55.695 93.420 ;
        RECT 56.595 93.375 56.885 93.420 ;
        RECT 59.115 93.375 59.405 93.420 ;
        RECT 63.265 93.375 63.555 93.605 ;
        RECT 41.170 93.020 41.490 93.280 ;
        RECT 48.990 93.020 49.310 93.280 ;
        RECT 51.290 93.020 51.610 93.280 ;
        RECT 54.065 93.220 54.355 93.265 ;
        RECT 54.510 93.220 54.830 93.280 ;
        RECT 54.065 93.080 54.830 93.220 ;
        RECT 54.065 93.035 54.355 93.080 ;
        RECT 54.510 93.020 54.830 93.080 ;
        RECT 55.010 93.220 55.300 93.265 ;
        RECT 57.110 93.220 57.400 93.265 ;
        RECT 58.680 93.220 58.970 93.265 ;
        RECT 55.010 93.080 58.970 93.220 ;
        RECT 55.010 93.035 55.300 93.080 ;
        RECT 57.110 93.035 57.400 93.080 ;
        RECT 58.680 93.035 58.970 93.080 ;
        RECT 64.170 93.020 64.490 93.280 ;
        RECT 25.530 92.880 25.850 92.940 ;
        RECT 32.445 92.880 32.735 92.925 ;
        RECT 25.530 92.740 32.735 92.880 ;
        RECT 25.530 92.680 25.850 92.740 ;
        RECT 32.445 92.695 32.735 92.740 ;
        RECT 34.270 92.880 34.590 92.940 ;
        RECT 53.145 92.880 53.435 92.925 ;
        RECT 60.490 92.880 60.810 92.940 ;
        RECT 34.270 92.740 60.810 92.880 ;
        RECT 34.270 92.680 34.590 92.740 ;
        RECT 53.145 92.695 53.435 92.740 ;
        RECT 60.490 92.680 60.810 92.740 ;
        RECT 60.950 92.880 61.270 92.940 ;
        RECT 61.425 92.880 61.715 92.925 ;
        RECT 60.950 92.740 61.715 92.880 ;
        RECT 60.950 92.680 61.270 92.740 ;
        RECT 61.425 92.695 61.715 92.740 ;
        RECT 62.805 92.880 63.095 92.925 ;
        RECT 65.180 92.880 65.320 94.100 ;
        RECT 67.250 94.055 67.540 94.100 ;
        RECT 74.765 94.055 75.055 94.285 ;
        RECT 83.580 94.240 83.720 94.440 ;
        RECT 76.220 94.100 83.720 94.240 ;
        RECT 66.025 93.900 66.315 93.945 ;
        RECT 66.470 93.900 66.790 93.960 ;
        RECT 66.025 93.760 66.790 93.900 ;
        RECT 66.025 93.715 66.315 93.760 ;
        RECT 66.470 93.700 66.790 93.760 ;
        RECT 68.770 93.900 69.090 93.960 ;
        RECT 74.290 93.900 74.610 93.960 ;
        RECT 75.685 93.900 75.975 93.945 ;
        RECT 68.770 93.760 74.060 93.900 ;
        RECT 68.770 93.700 69.090 93.760 ;
        RECT 65.550 93.360 65.870 93.620 ;
        RECT 66.905 93.560 67.195 93.605 ;
        RECT 68.095 93.560 68.385 93.605 ;
        RECT 70.615 93.560 70.905 93.605 ;
        RECT 66.905 93.420 70.905 93.560 ;
        RECT 73.920 93.560 74.060 93.760 ;
        RECT 74.290 93.760 75.975 93.900 ;
        RECT 74.290 93.700 74.610 93.760 ;
        RECT 75.685 93.715 75.975 93.760 ;
        RECT 76.220 93.560 76.360 94.100 ;
        RECT 80.745 93.900 81.035 93.945 ;
        RECT 80.745 93.760 81.420 93.900 ;
        RECT 80.745 93.715 81.035 93.760 ;
        RECT 73.920 93.420 76.360 93.560 ;
        RECT 66.905 93.375 67.195 93.420 ;
        RECT 68.095 93.375 68.385 93.420 ;
        RECT 70.615 93.375 70.905 93.420 ;
        RECT 81.280 93.280 81.420 93.760 ;
        RECT 83.045 93.715 83.335 93.945 ;
        RECT 81.650 93.360 81.970 93.620 ;
        RECT 66.510 93.220 66.800 93.265 ;
        RECT 68.610 93.220 68.900 93.265 ;
        RECT 70.180 93.220 70.470 93.265 ;
        RECT 66.510 93.080 70.470 93.220 ;
        RECT 66.510 93.035 66.800 93.080 ;
        RECT 68.610 93.035 68.900 93.080 ;
        RECT 70.180 93.035 70.470 93.080 ;
        RECT 81.190 93.220 81.510 93.280 ;
        RECT 82.125 93.220 82.415 93.265 ;
        RECT 81.190 93.080 82.415 93.220 ;
        RECT 83.120 93.220 83.260 93.715 ;
        RECT 83.580 93.560 83.720 94.100 ;
        RECT 83.965 94.240 84.255 94.285 ;
        RECT 85.790 94.240 86.110 94.300 ;
        RECT 91.310 94.240 91.630 94.300 ;
        RECT 95.925 94.240 96.215 94.285 ;
        RECT 105.110 94.240 105.430 94.300 ;
        RECT 83.965 94.100 86.110 94.240 ;
        RECT 83.965 94.055 84.255 94.100 ;
        RECT 85.790 94.040 86.110 94.100 ;
        RECT 86.340 94.100 96.215 94.240 ;
        RECT 86.340 93.945 86.480 94.100 ;
        RECT 91.310 94.040 91.630 94.100 ;
        RECT 95.925 94.055 96.215 94.100 ;
        RECT 100.600 94.100 108.560 94.240 ;
        RECT 84.425 93.900 84.715 93.945 ;
        RECT 86.265 93.900 86.555 93.945 ;
        RECT 84.425 93.760 86.555 93.900 ;
        RECT 84.425 93.715 84.715 93.760 ;
        RECT 86.265 93.715 86.555 93.760 ;
        RECT 88.090 93.700 88.410 93.960 ;
        RECT 89.470 93.945 89.790 93.960 ;
        RECT 89.440 93.715 89.790 93.945 ;
        RECT 89.470 93.700 89.790 93.715 ;
        RECT 95.450 93.700 95.770 93.960 ;
        RECT 96.370 93.700 96.690 93.960 ;
        RECT 97.750 93.700 98.070 93.960 ;
        RECT 98.210 93.900 98.530 93.960 ;
        RECT 100.600 93.945 100.740 94.100 ;
        RECT 105.110 94.040 105.430 94.100 ;
        RECT 101.890 93.945 102.210 93.960 ;
        RECT 99.145 93.900 99.435 93.945 ;
        RECT 98.210 93.760 99.435 93.900 ;
        RECT 98.210 93.700 98.530 93.760 ;
        RECT 99.145 93.715 99.435 93.760 ;
        RECT 100.525 93.715 100.815 93.945 ;
        RECT 101.860 93.900 102.210 93.945 ;
        RECT 101.695 93.760 102.210 93.900 ;
        RECT 101.860 93.715 102.210 93.760 ;
        RECT 101.890 93.700 102.210 93.715 ;
        RECT 108.420 93.620 108.560 94.100 ;
        RECT 108.880 93.900 109.020 94.440 ;
        RECT 111.550 94.440 113.235 94.580 ;
        RECT 111.550 94.380 111.870 94.440 ;
        RECT 112.945 94.395 113.235 94.440 ;
        RECT 124.430 94.580 124.750 94.640 ;
        RECT 124.905 94.580 125.195 94.625 ;
        RECT 124.430 94.440 125.195 94.580 ;
        RECT 124.430 94.380 124.750 94.440 ;
        RECT 124.905 94.395 125.195 94.440 ;
        RECT 133.185 94.580 133.475 94.625 ;
        RECT 135.010 94.580 135.330 94.640 ;
        RECT 136.405 94.580 136.695 94.625 ;
        RECT 133.185 94.440 133.860 94.580 ;
        RECT 133.185 94.395 133.475 94.440 ;
        RECT 112.485 94.240 112.775 94.285 ;
        RECT 129.490 94.240 129.810 94.300 ;
        RECT 112.485 94.100 129.810 94.240 ;
        RECT 112.485 94.055 112.775 94.100 ;
        RECT 129.490 94.040 129.810 94.100 ;
        RECT 115.245 93.900 115.535 93.945 ;
        RECT 108.880 93.760 115.535 93.900 ;
        RECT 115.245 93.715 115.535 93.760 ;
        RECT 117.545 93.715 117.835 93.945 ;
        RECT 85.345 93.560 85.635 93.605 ;
        RECT 83.580 93.420 85.635 93.560 ;
        RECT 85.345 93.375 85.635 93.420 ;
        RECT 85.790 93.360 86.110 93.620 ;
        RECT 86.710 93.360 87.030 93.620 ;
        RECT 88.985 93.560 89.275 93.605 ;
        RECT 90.175 93.560 90.465 93.605 ;
        RECT 92.695 93.560 92.985 93.605 ;
        RECT 88.985 93.420 92.985 93.560 ;
        RECT 88.985 93.375 89.275 93.420 ;
        RECT 90.175 93.375 90.465 93.420 ;
        RECT 92.695 93.375 92.985 93.420 ;
        RECT 101.405 93.560 101.695 93.605 ;
        RECT 102.595 93.560 102.885 93.605 ;
        RECT 105.115 93.560 105.405 93.605 ;
        RECT 101.405 93.420 105.405 93.560 ;
        RECT 101.405 93.375 101.695 93.420 ;
        RECT 102.595 93.375 102.885 93.420 ;
        RECT 105.115 93.375 105.405 93.420 ;
        RECT 108.330 93.360 108.650 93.620 ;
        RECT 113.850 93.360 114.170 93.620 ;
        RECT 114.325 93.375 114.615 93.605 ;
        RECT 114.785 93.560 115.075 93.605 ;
        RECT 117.620 93.560 117.760 93.715 ;
        RECT 117.990 93.700 118.310 93.960 ;
        RECT 118.925 93.715 119.215 93.945 ;
        RECT 119.385 93.900 119.675 93.945 ;
        RECT 120.290 93.900 120.610 93.960 ;
        RECT 119.385 93.760 120.610 93.900 ;
        RECT 119.385 93.715 119.675 93.760 ;
        RECT 118.450 93.560 118.770 93.620 ;
        RECT 114.785 93.420 118.770 93.560 ;
        RECT 119.000 93.560 119.140 93.715 ;
        RECT 120.290 93.700 120.610 93.760 ;
        RECT 121.210 93.900 121.530 93.960 ;
        RECT 121.685 93.900 121.975 93.945 ;
        RECT 121.210 93.760 121.975 93.900 ;
        RECT 121.210 93.700 121.530 93.760 ;
        RECT 121.685 93.715 121.975 93.760 ;
        RECT 123.065 93.900 123.355 93.945 ;
        RECT 123.065 93.760 123.740 93.900 ;
        RECT 123.065 93.715 123.355 93.760 ;
        RECT 119.830 93.560 120.150 93.620 ;
        RECT 120.765 93.560 121.055 93.605 ;
        RECT 119.000 93.420 121.055 93.560 ;
        RECT 114.785 93.375 115.075 93.420 ;
        RECT 86.800 93.220 86.940 93.360 ;
        RECT 83.120 93.080 86.940 93.220 ;
        RECT 88.590 93.220 88.880 93.265 ;
        RECT 90.690 93.220 90.980 93.265 ;
        RECT 92.260 93.220 92.550 93.265 ;
        RECT 88.590 93.080 92.550 93.220 ;
        RECT 81.190 93.020 81.510 93.080 ;
        RECT 82.125 93.035 82.415 93.080 ;
        RECT 88.590 93.035 88.880 93.080 ;
        RECT 90.690 93.035 90.980 93.080 ;
        RECT 92.260 93.035 92.550 93.080 ;
        RECT 93.610 93.220 93.930 93.280 ;
        RECT 95.005 93.220 95.295 93.265 ;
        RECT 97.290 93.220 97.610 93.280 ;
        RECT 93.610 93.080 97.610 93.220 ;
        RECT 93.610 93.020 93.930 93.080 ;
        RECT 95.005 93.035 95.295 93.080 ;
        RECT 97.290 93.020 97.610 93.080 ;
        RECT 101.010 93.220 101.300 93.265 ;
        RECT 103.110 93.220 103.400 93.265 ;
        RECT 104.680 93.220 104.970 93.265 ;
        RECT 110.630 93.220 110.950 93.280 ;
        RECT 114.400 93.220 114.540 93.375 ;
        RECT 118.450 93.360 118.770 93.420 ;
        RECT 119.830 93.360 120.150 93.420 ;
        RECT 120.765 93.375 121.055 93.420 ;
        RECT 117.530 93.220 117.850 93.280 ;
        RECT 101.010 93.080 104.970 93.220 ;
        RECT 101.010 93.035 101.300 93.080 ;
        RECT 103.110 93.035 103.400 93.080 ;
        RECT 104.680 93.035 104.970 93.080 ;
        RECT 105.200 93.080 109.480 93.220 ;
        RECT 62.805 92.740 65.320 92.880 ;
        RECT 62.805 92.695 63.095 92.740 ;
        RECT 76.590 92.680 76.910 92.940 ;
        RECT 79.825 92.880 80.115 92.925 ;
        RECT 80.270 92.880 80.590 92.940 ;
        RECT 79.825 92.740 80.590 92.880 ;
        RECT 79.825 92.695 80.115 92.740 ;
        RECT 80.270 92.680 80.590 92.740 ;
        RECT 87.645 92.880 87.935 92.925 ;
        RECT 89.930 92.880 90.250 92.940 ;
        RECT 87.645 92.740 90.250 92.880 ;
        RECT 87.645 92.695 87.935 92.740 ;
        RECT 89.930 92.680 90.250 92.740 ;
        RECT 92.690 92.880 93.010 92.940 ;
        RECT 105.200 92.880 105.340 93.080 ;
        RECT 92.690 92.740 105.340 92.880 ;
        RECT 107.425 92.880 107.715 92.925 ;
        RECT 108.790 92.880 109.110 92.940 ;
        RECT 107.425 92.740 109.110 92.880 ;
        RECT 109.340 92.880 109.480 93.080 ;
        RECT 110.630 93.080 117.850 93.220 ;
        RECT 123.600 93.220 123.740 93.760 ;
        RECT 123.985 93.715 124.275 93.945 ;
        RECT 124.060 93.560 124.200 93.715 ;
        RECT 124.430 93.700 124.750 93.960 ;
        RECT 125.365 93.900 125.655 93.945 ;
        RECT 126.730 93.900 127.050 93.960 ;
        RECT 127.650 93.945 127.970 93.960 ;
        RECT 133.720 93.945 133.860 94.440 ;
        RECT 135.010 94.440 136.695 94.580 ;
        RECT 135.010 94.380 135.330 94.440 ;
        RECT 136.405 94.395 136.695 94.440 ;
        RECT 140.070 94.380 140.390 94.640 ;
        RECT 141.450 94.580 141.770 94.640 ;
        RECT 143.765 94.580 144.055 94.625 ;
        RECT 141.450 94.440 144.055 94.580 ;
        RECT 141.450 94.380 141.770 94.440 ;
        RECT 143.765 94.395 144.055 94.440 ;
        RECT 144.210 94.380 144.530 94.640 ;
        RECT 147.905 94.580 148.195 94.625 ;
        RECT 148.350 94.580 148.670 94.640 ;
        RECT 150.190 94.580 150.510 94.640 ;
        RECT 147.905 94.440 148.670 94.580 ;
        RECT 147.905 94.395 148.195 94.440 ;
        RECT 148.350 94.380 148.670 94.440 ;
        RECT 149.820 94.440 150.510 94.580 ;
        RECT 135.485 94.240 135.775 94.285 ;
        RECT 140.160 94.240 140.300 94.380 ;
        RECT 135.485 94.100 138.920 94.240 ;
        RECT 135.485 94.055 135.775 94.100 ;
        RECT 127.620 93.900 127.970 93.945 ;
        RECT 125.365 93.760 127.050 93.900 ;
        RECT 127.455 93.760 127.970 93.900 ;
        RECT 125.365 93.715 125.655 93.760 ;
        RECT 125.440 93.560 125.580 93.715 ;
        RECT 126.730 93.700 127.050 93.760 ;
        RECT 127.620 93.715 127.970 93.760 ;
        RECT 133.645 93.715 133.935 93.945 ;
        RECT 134.565 93.900 134.855 93.945 ;
        RECT 136.850 93.900 137.170 93.960 ;
        RECT 134.565 93.760 137.170 93.900 ;
        RECT 134.565 93.715 134.855 93.760 ;
        RECT 127.650 93.700 127.970 93.715 ;
        RECT 124.060 93.420 125.580 93.560 ;
        RECT 126.270 93.360 126.590 93.620 ;
        RECT 127.165 93.560 127.455 93.605 ;
        RECT 128.355 93.560 128.645 93.605 ;
        RECT 130.875 93.560 131.165 93.605 ;
        RECT 127.165 93.420 131.165 93.560 ;
        RECT 133.720 93.560 133.860 93.715 ;
        RECT 136.850 93.700 137.170 93.760 ;
        RECT 137.310 93.700 137.630 93.960 ;
        RECT 137.770 93.900 138.090 93.960 ;
        RECT 138.780 93.945 138.920 94.100 ;
        RECT 139.700 94.100 140.300 94.240 ;
        RECT 140.530 94.240 140.850 94.300 ;
        RECT 141.925 94.240 142.215 94.285 ;
        RECT 142.370 94.240 142.690 94.300 ;
        RECT 140.530 94.100 142.690 94.240 ;
        RECT 139.700 93.945 139.840 94.100 ;
        RECT 140.530 94.040 140.850 94.100 ;
        RECT 141.925 94.055 142.215 94.100 ;
        RECT 142.370 94.040 142.690 94.100 ;
        RECT 142.845 94.240 143.135 94.285 ;
        RECT 146.510 94.240 146.830 94.300 ;
        RECT 142.845 94.100 146.830 94.240 ;
        RECT 142.845 94.055 143.135 94.100 ;
        RECT 146.510 94.040 146.830 94.100 ;
        RECT 138.245 93.900 138.535 93.945 ;
        RECT 137.770 93.760 138.535 93.900 ;
        RECT 137.770 93.700 138.090 93.760 ;
        RECT 138.245 93.715 138.535 93.760 ;
        RECT 138.705 93.715 138.995 93.945 ;
        RECT 139.625 93.715 139.915 93.945 ;
        RECT 140.070 93.700 140.390 93.960 ;
        RECT 141.005 93.715 141.295 93.945 ;
        RECT 143.750 93.900 144.070 93.960 ;
        RECT 146.985 93.900 147.275 93.945 ;
        RECT 143.750 93.760 147.275 93.900 ;
        RECT 141.080 93.560 141.220 93.715 ;
        RECT 143.750 93.700 144.070 93.760 ;
        RECT 146.985 93.715 147.275 93.760 ;
        RECT 149.270 93.700 149.590 93.960 ;
        RECT 149.820 93.945 149.960 94.440 ;
        RECT 150.190 94.380 150.510 94.440 ;
        RECT 152.030 94.380 152.350 94.640 ;
        RECT 149.745 93.715 150.035 93.945 ;
        RECT 150.205 93.715 150.495 93.945 ;
        RECT 133.720 93.420 141.220 93.560 ;
        RECT 150.280 93.560 150.420 93.715 ;
        RECT 151.110 93.700 151.430 93.960 ;
        RECT 155.250 93.700 155.570 93.960 ;
        RECT 153.870 93.560 154.190 93.620 ;
        RECT 150.280 93.420 154.190 93.560 ;
        RECT 127.165 93.375 127.455 93.420 ;
        RECT 128.355 93.375 128.645 93.420 ;
        RECT 130.875 93.375 131.165 93.420 ;
        RECT 153.870 93.360 154.190 93.420 ;
        RECT 124.430 93.220 124.750 93.280 ;
        RECT 123.600 93.080 124.750 93.220 ;
        RECT 110.630 93.020 110.950 93.080 ;
        RECT 117.530 93.020 117.850 93.080 ;
        RECT 124.430 93.020 124.750 93.080 ;
        RECT 126.770 93.220 127.060 93.265 ;
        RECT 128.870 93.220 129.160 93.265 ;
        RECT 130.440 93.220 130.730 93.265 ;
        RECT 139.165 93.220 139.455 93.265 ;
        RECT 126.770 93.080 130.730 93.220 ;
        RECT 126.770 93.035 127.060 93.080 ;
        RECT 128.870 93.035 129.160 93.080 ;
        RECT 130.440 93.035 130.730 93.080 ;
        RECT 132.800 93.080 139.455 93.220 ;
        RECT 112.010 92.880 112.330 92.940 ;
        RECT 109.340 92.740 112.330 92.880 ;
        RECT 92.690 92.680 93.010 92.740 ;
        RECT 107.425 92.695 107.715 92.740 ;
        RECT 108.790 92.680 109.110 92.740 ;
        RECT 112.010 92.680 112.330 92.740 ;
        RECT 114.310 92.880 114.630 92.940 ;
        RECT 116.625 92.880 116.915 92.925 ;
        RECT 114.310 92.740 116.915 92.880 ;
        RECT 114.310 92.680 114.630 92.740 ;
        RECT 116.625 92.695 116.915 92.740 ;
        RECT 129.490 92.880 129.810 92.940 ;
        RECT 132.800 92.880 132.940 93.080 ;
        RECT 139.165 93.035 139.455 93.080 ;
        RECT 129.490 92.740 132.940 92.880 ;
        RECT 129.490 92.680 129.810 92.740 ;
        RECT 22.700 92.060 157.020 92.540 ;
        RECT 30.590 91.860 30.910 91.920 ;
        RECT 32.890 91.860 33.210 91.920 ;
        RECT 30.590 91.720 33.210 91.860 ;
        RECT 30.590 91.660 30.910 91.720 ;
        RECT 32.890 91.660 33.210 91.720 ;
        RECT 36.110 91.660 36.430 91.920 ;
        RECT 41.185 91.675 41.475 91.905 ;
        RECT 24.650 91.520 24.940 91.565 ;
        RECT 26.750 91.520 27.040 91.565 ;
        RECT 28.320 91.520 28.610 91.565 ;
        RECT 24.650 91.380 28.610 91.520 ;
        RECT 41.260 91.520 41.400 91.675 ;
        RECT 42.090 91.660 42.410 91.920 ;
        RECT 49.465 91.675 49.755 91.905 ;
        RECT 49.910 91.860 50.230 91.920 ;
        RECT 50.385 91.860 50.675 91.905 ;
        RECT 49.910 91.720 50.675 91.860 ;
        RECT 42.565 91.520 42.855 91.565 ;
        RECT 41.260 91.380 42.855 91.520 ;
        RECT 49.540 91.520 49.680 91.675 ;
        RECT 49.910 91.660 50.230 91.720 ;
        RECT 50.385 91.675 50.675 91.720 ;
        RECT 53.130 91.860 53.450 91.920 ;
        RECT 56.365 91.860 56.655 91.905 ;
        RECT 53.130 91.720 56.655 91.860 ;
        RECT 53.130 91.660 53.450 91.720 ;
        RECT 56.365 91.675 56.655 91.720 ;
        RECT 65.550 91.860 65.870 91.920 ;
        RECT 66.485 91.860 66.775 91.905 ;
        RECT 65.550 91.720 66.775 91.860 ;
        RECT 65.550 91.660 65.870 91.720 ;
        RECT 66.485 91.675 66.775 91.720 ;
        RECT 67.850 91.860 68.170 91.920 ;
        RECT 69.705 91.860 69.995 91.905 ;
        RECT 67.850 91.720 69.995 91.860 ;
        RECT 67.850 91.660 68.170 91.720 ;
        RECT 69.705 91.675 69.995 91.720 ;
        RECT 71.070 91.860 71.390 91.920 ;
        RECT 85.790 91.860 86.110 91.920 ;
        RECT 89.470 91.860 89.790 91.920 ;
        RECT 90.405 91.860 90.695 91.905 ;
        RECT 71.070 91.720 72.680 91.860 ;
        RECT 71.070 91.660 71.390 91.720 ;
        RECT 60.030 91.520 60.350 91.580 ;
        RECT 49.540 91.380 60.350 91.520 ;
        RECT 24.650 91.335 24.940 91.380 ;
        RECT 26.750 91.335 27.040 91.380 ;
        RECT 28.320 91.335 28.610 91.380 ;
        RECT 42.565 91.335 42.855 91.380 ;
        RECT 60.030 91.320 60.350 91.380 ;
        RECT 64.170 91.520 64.490 91.580 ;
        RECT 67.940 91.520 68.080 91.660 ;
        RECT 64.170 91.380 68.080 91.520 ;
        RECT 64.170 91.320 64.490 91.380 ;
        RECT 25.045 91.180 25.335 91.225 ;
        RECT 26.235 91.180 26.525 91.225 ;
        RECT 28.755 91.180 29.045 91.225 ;
        RECT 25.045 91.040 29.045 91.180 ;
        RECT 25.045 90.995 25.335 91.040 ;
        RECT 26.235 90.995 26.525 91.040 ;
        RECT 28.755 90.995 29.045 91.040 ;
        RECT 34.745 91.180 35.035 91.225 ;
        RECT 36.570 91.180 36.890 91.240 ;
        RECT 37.045 91.180 37.335 91.225 ;
        RECT 34.745 91.040 37.335 91.180 ;
        RECT 34.745 90.995 35.035 91.040 ;
        RECT 36.570 90.980 36.890 91.040 ;
        RECT 37.045 90.995 37.335 91.040 ;
        RECT 44.390 91.180 44.710 91.240 ;
        RECT 47.625 91.180 47.915 91.225 ;
        RECT 50.845 91.180 51.135 91.225 ;
        RECT 44.390 91.040 51.135 91.180 ;
        RECT 44.390 90.980 44.710 91.040 ;
        RECT 24.165 90.840 24.455 90.885 ;
        RECT 26.910 90.840 27.230 90.900 ;
        RECT 28.290 90.840 28.610 90.900 ;
        RECT 24.165 90.700 28.610 90.840 ;
        RECT 24.165 90.655 24.455 90.700 ;
        RECT 26.910 90.640 27.230 90.700 ;
        RECT 28.290 90.640 28.610 90.700 ;
        RECT 32.445 90.840 32.735 90.885 ;
        RECT 32.890 90.840 33.210 90.900 ;
        RECT 32.445 90.700 33.210 90.840 ;
        RECT 32.445 90.655 32.735 90.700 ;
        RECT 32.890 90.640 33.210 90.700 ;
        RECT 37.490 90.640 37.810 90.900 ;
        RECT 37.965 90.655 38.255 90.885 ;
        RECT 38.425 90.840 38.715 90.885 ;
        RECT 43.010 90.840 43.330 90.900 ;
        RECT 43.485 90.840 43.775 90.885 ;
        RECT 38.425 90.700 42.780 90.840 ;
        RECT 38.425 90.655 38.715 90.700 ;
        RECT 25.530 90.545 25.850 90.560 ;
        RECT 25.500 90.500 25.850 90.545 ;
        RECT 25.335 90.360 25.850 90.500 ;
        RECT 25.500 90.315 25.850 90.360 ;
        RECT 25.530 90.300 25.850 90.315 ;
        RECT 36.110 90.500 36.430 90.560 ;
        RECT 38.040 90.500 38.180 90.655 ;
        RECT 36.110 90.360 38.180 90.500 ;
        RECT 36.110 90.300 36.430 90.360 ;
        RECT 40.250 90.300 40.570 90.560 ;
        RECT 31.050 89.960 31.370 90.220 ;
        RECT 41.170 90.205 41.490 90.220 ;
        RECT 41.170 89.975 41.555 90.205 ;
        RECT 42.640 90.160 42.780 90.700 ;
        RECT 43.010 90.700 43.775 90.840 ;
        RECT 43.010 90.640 43.330 90.700 ;
        RECT 43.485 90.655 43.775 90.700 ;
        RECT 43.930 90.640 44.250 90.900 ;
        RECT 44.850 90.840 45.170 90.900 ;
        RECT 45.400 90.885 45.540 91.040 ;
        RECT 47.625 90.995 47.915 91.040 ;
        RECT 50.845 90.995 51.135 91.040 ;
        RECT 51.290 91.180 51.610 91.240 ;
        RECT 54.510 91.180 54.830 91.240 ;
        RECT 51.290 91.040 54.830 91.180 ;
        RECT 51.290 90.980 51.610 91.040 ;
        RECT 44.480 90.700 45.170 90.840 ;
        RECT 44.480 90.500 44.620 90.700 ;
        RECT 44.850 90.640 45.170 90.700 ;
        RECT 45.325 90.655 45.615 90.885 ;
        RECT 47.165 90.840 47.455 90.885 ;
        RECT 49.910 90.840 50.230 90.900 ;
        RECT 52.210 90.840 52.530 90.900 ;
        RECT 52.760 90.885 52.900 91.040 ;
        RECT 54.510 90.980 54.830 91.040 ;
        RECT 57.285 91.180 57.575 91.225 ;
        RECT 58.190 91.180 58.510 91.240 ;
        RECT 60.505 91.180 60.795 91.225 ;
        RECT 57.285 91.040 60.795 91.180 ;
        RECT 57.285 90.995 57.575 91.040 ;
        RECT 47.165 90.700 50.230 90.840 ;
        RECT 52.015 90.700 52.530 90.840 ;
        RECT 47.165 90.655 47.455 90.700 ;
        RECT 49.910 90.640 50.230 90.700 ;
        RECT 52.210 90.640 52.530 90.700 ;
        RECT 52.685 90.655 52.975 90.885 ;
        RECT 53.145 90.840 53.435 90.885 ;
        RECT 53.590 90.840 53.910 90.900 ;
        RECT 53.145 90.700 53.910 90.840 ;
        RECT 53.145 90.655 53.435 90.700 ;
        RECT 53.590 90.640 53.910 90.700 ;
        RECT 54.050 90.640 54.370 90.900 ;
        RECT 55.905 90.840 56.195 90.885 ;
        RECT 57.360 90.840 57.500 90.995 ;
        RECT 58.190 90.980 58.510 91.040 ;
        RECT 60.505 90.995 60.795 91.040 ;
        RECT 66.930 91.180 67.250 91.240 ;
        RECT 67.865 91.180 68.155 91.225 ;
        RECT 66.930 91.040 71.760 91.180 ;
        RECT 66.930 90.980 67.250 91.040 ;
        RECT 67.865 90.995 68.155 91.040 ;
        RECT 55.905 90.700 57.500 90.840 ;
        RECT 55.905 90.655 56.195 90.700 ;
        RECT 57.745 90.655 58.035 90.885 ;
        RECT 60.045 90.840 60.335 90.885 ;
        RECT 60.950 90.840 61.270 90.900 ;
        RECT 61.885 90.840 62.175 90.885 ;
        RECT 60.045 90.700 60.720 90.840 ;
        RECT 60.045 90.655 60.335 90.700 ;
        RECT 46.705 90.500 46.995 90.545 ;
        RECT 52.300 90.500 52.440 90.640 ;
        RECT 55.445 90.500 55.735 90.545 ;
        RECT 44.480 90.360 46.995 90.500 ;
        RECT 46.705 90.315 46.995 90.360 ;
        RECT 47.240 90.360 50.140 90.500 ;
        RECT 52.300 90.360 55.735 90.500 ;
        RECT 57.820 90.500 57.960 90.655 ;
        RECT 58.650 90.500 58.970 90.560 ;
        RECT 60.580 90.500 60.720 90.700 ;
        RECT 60.950 90.700 62.175 90.840 ;
        RECT 60.950 90.640 61.270 90.700 ;
        RECT 61.885 90.655 62.175 90.700 ;
        RECT 67.405 90.655 67.695 90.885 ;
        RECT 62.790 90.500 63.110 90.560 ;
        RECT 57.820 90.360 60.260 90.500 ;
        RECT 60.580 90.360 63.110 90.500 ;
        RECT 67.480 90.500 67.620 90.655 ;
        RECT 68.310 90.640 68.630 90.900 ;
        RECT 68.770 90.640 69.090 90.900 ;
        RECT 70.625 90.825 70.915 90.885 ;
        RECT 71.620 90.840 71.760 91.040 ;
        RECT 72.540 90.885 72.680 91.720 ;
        RECT 85.790 91.720 88.780 91.860 ;
        RECT 85.790 91.660 86.110 91.720 ;
        RECT 81.190 91.520 81.510 91.580 ;
        RECT 88.105 91.520 88.395 91.565 ;
        RECT 81.190 91.380 88.395 91.520 ;
        RECT 88.640 91.520 88.780 91.720 ;
        RECT 89.470 91.720 90.695 91.860 ;
        RECT 89.470 91.660 89.790 91.720 ;
        RECT 90.405 91.675 90.695 91.720 ;
        RECT 90.850 91.860 91.170 91.920 ;
        RECT 94.085 91.860 94.375 91.905 ;
        RECT 90.850 91.720 94.375 91.860 ;
        RECT 90.850 91.660 91.170 91.720 ;
        RECT 94.085 91.675 94.375 91.720 ;
        RECT 98.210 91.660 98.530 91.920 ;
        RECT 100.985 91.860 101.275 91.905 ;
        RECT 101.430 91.860 101.750 91.920 ;
        RECT 100.985 91.720 101.750 91.860 ;
        RECT 100.985 91.675 101.275 91.720 ;
        RECT 101.430 91.660 101.750 91.720 ;
        RECT 101.905 91.860 102.195 91.905 ;
        RECT 102.350 91.860 102.670 91.920 ;
        RECT 111.565 91.860 111.855 91.905 ;
        RECT 101.905 91.720 102.670 91.860 ;
        RECT 101.905 91.675 102.195 91.720 ;
        RECT 102.350 91.660 102.670 91.720 ;
        RECT 106.580 91.720 111.855 91.860 ;
        RECT 98.300 91.520 98.440 91.660 ;
        RECT 88.640 91.380 95.220 91.520 ;
        RECT 81.190 91.320 81.510 91.380 ;
        RECT 83.120 91.225 83.260 91.380 ;
        RECT 88.105 91.335 88.395 91.380 ;
        RECT 81.665 91.180 81.955 91.225 ;
        RECT 78.980 91.040 81.955 91.180 ;
        RECT 72.005 90.840 72.295 90.885 ;
        RECT 70.625 90.685 71.300 90.825 ;
        RECT 71.620 90.700 72.295 90.840 ;
        RECT 70.625 90.655 70.915 90.685 ;
        RECT 71.160 90.500 71.300 90.685 ;
        RECT 72.005 90.655 72.295 90.700 ;
        RECT 72.465 90.655 72.755 90.885 ;
        RECT 73.385 90.840 73.675 90.885 ;
        RECT 76.590 90.840 76.910 90.900 ;
        RECT 78.980 90.885 79.120 91.040 ;
        RECT 81.665 90.995 81.955 91.040 ;
        RECT 83.045 90.995 83.335 91.225 ;
        RECT 89.930 90.980 90.250 91.240 ;
        RECT 92.690 91.180 93.010 91.240 ;
        RECT 90.940 91.040 93.010 91.180 ;
        RECT 73.385 90.700 76.910 90.840 ;
        RECT 73.385 90.655 73.675 90.700 ;
        RECT 76.590 90.640 76.910 90.700 ;
        RECT 78.905 90.655 79.195 90.885 ;
        RECT 80.270 90.640 80.590 90.900 ;
        RECT 81.205 90.840 81.495 90.885 ;
        RECT 82.570 90.840 82.890 90.900 ;
        RECT 81.205 90.700 82.890 90.840 ;
        RECT 81.205 90.655 81.495 90.700 ;
        RECT 82.570 90.640 82.890 90.700 ;
        RECT 83.505 90.655 83.795 90.885 ;
        RECT 83.965 90.840 84.255 90.885 ;
        RECT 90.940 90.840 91.080 91.040 ;
        RECT 92.690 90.980 93.010 91.040 ;
        RECT 95.080 90.900 95.220 91.380 ;
        RECT 96.460 91.380 98.440 91.520 ;
        RECT 99.145 91.520 99.435 91.565 ;
        RECT 103.285 91.520 103.575 91.565 ;
        RECT 99.145 91.380 103.575 91.520 ;
        RECT 83.965 90.700 91.080 90.840 ;
        RECT 91.325 90.840 91.615 90.885 ;
        RECT 91.770 90.840 92.090 90.900 ;
        RECT 91.325 90.700 92.090 90.840 ;
        RECT 83.965 90.655 84.255 90.700 ;
        RECT 91.325 90.655 91.615 90.700 ;
        RECT 72.925 90.500 73.215 90.545 ;
        RECT 67.480 90.360 73.215 90.500 ;
        RECT 43.470 90.160 43.790 90.220 ;
        RECT 47.240 90.160 47.380 90.360 ;
        RECT 42.640 90.020 47.380 90.160 ;
        RECT 41.170 89.960 41.490 89.975 ;
        RECT 43.470 89.960 43.790 90.020 ;
        RECT 49.450 89.960 49.770 90.220 ;
        RECT 50.000 90.160 50.140 90.360 ;
        RECT 55.445 90.315 55.735 90.360 ;
        RECT 58.650 90.300 58.970 90.360 ;
        RECT 54.970 90.160 55.290 90.220 ;
        RECT 50.000 90.020 55.290 90.160 ;
        RECT 54.970 89.960 55.290 90.020 ;
        RECT 59.110 90.160 59.430 90.220 ;
        RECT 59.585 90.160 59.875 90.205 ;
        RECT 59.110 90.020 59.875 90.160 ;
        RECT 60.120 90.160 60.260 90.360 ;
        RECT 62.790 90.300 63.110 90.360 ;
        RECT 72.925 90.315 73.215 90.360 ;
        RECT 81.650 90.500 81.970 90.560 ;
        RECT 83.580 90.500 83.720 90.655 ;
        RECT 81.650 90.360 83.720 90.500 ;
        RECT 81.650 90.300 81.970 90.360 ;
        RECT 63.725 90.160 64.015 90.205 ;
        RECT 60.120 90.020 64.015 90.160 ;
        RECT 59.110 89.960 59.430 90.020 ;
        RECT 59.585 89.975 59.875 90.020 ;
        RECT 63.725 89.975 64.015 90.020 ;
        RECT 68.310 90.160 68.630 90.220 ;
        RECT 71.530 90.160 71.850 90.220 ;
        RECT 68.310 90.020 71.850 90.160 ;
        RECT 68.310 89.960 68.630 90.020 ;
        RECT 71.530 89.960 71.850 90.020 ;
        RECT 76.590 90.160 76.910 90.220 ;
        RECT 77.985 90.160 78.275 90.205 ;
        RECT 76.590 90.020 78.275 90.160 ;
        RECT 76.590 89.960 76.910 90.020 ;
        RECT 77.985 89.975 78.275 90.020 ;
        RECT 78.430 90.160 78.750 90.220 ;
        RECT 84.040 90.160 84.180 90.655 ;
        RECT 91.770 90.640 92.090 90.700 ;
        RECT 94.990 90.640 95.310 90.900 ;
        RECT 95.465 90.840 95.755 90.885 ;
        RECT 95.910 90.840 96.230 90.900 ;
        RECT 96.460 90.885 96.600 91.380 ;
        RECT 99.145 91.335 99.435 91.380 ;
        RECT 103.285 91.335 103.575 91.380 ;
        RECT 99.220 91.180 99.360 91.335 ;
        RECT 98.300 91.040 99.360 91.180 ;
        RECT 95.465 90.700 96.230 90.840 ;
        RECT 95.465 90.655 95.755 90.700 ;
        RECT 95.910 90.640 96.230 90.700 ;
        RECT 96.385 90.655 96.675 90.885 ;
        RECT 96.845 90.840 97.135 90.885 ;
        RECT 97.750 90.840 98.070 90.900 ;
        RECT 98.300 90.840 98.440 91.040 ;
        RECT 96.845 90.700 98.440 90.840 ;
        RECT 98.685 90.840 98.975 90.885 ;
        RECT 98.685 90.700 103.500 90.840 ;
        RECT 96.845 90.655 97.135 90.700 ;
        RECT 97.750 90.640 98.070 90.700 ;
        RECT 98.685 90.655 98.975 90.700 ;
        RECT 103.360 90.560 103.500 90.700 ;
        RECT 104.650 90.640 104.970 90.900 ;
        RECT 105.110 90.640 105.430 90.900 ;
        RECT 105.570 90.640 105.890 90.900 ;
        RECT 106.580 90.885 106.720 91.720 ;
        RECT 111.565 91.675 111.855 91.720 ;
        RECT 112.010 91.860 112.330 91.920 ;
        RECT 112.010 91.720 114.080 91.860 ;
        RECT 112.010 91.660 112.330 91.720 ;
        RECT 108.345 91.520 108.635 91.565 ;
        RECT 109.250 91.520 109.570 91.580 ;
        RECT 108.345 91.380 109.570 91.520 ;
        RECT 108.345 91.335 108.635 91.380 ;
        RECT 109.250 91.320 109.570 91.380 ;
        RECT 109.710 91.520 110.030 91.580 ;
        RECT 113.405 91.520 113.695 91.565 ;
        RECT 109.710 91.380 113.695 91.520 ;
        RECT 113.940 91.520 114.080 91.720 ;
        RECT 114.310 91.660 114.630 91.920 ;
        RECT 117.530 91.660 117.850 91.920 ;
        RECT 124.430 91.860 124.750 91.920 ;
        RECT 128.110 91.860 128.430 91.920 ;
        RECT 124.430 91.720 128.430 91.860 ;
        RECT 124.430 91.660 124.750 91.720 ;
        RECT 128.110 91.660 128.430 91.720 ;
        RECT 128.570 91.660 128.890 91.920 ;
        RECT 149.270 91.860 149.590 91.920 ;
        RECT 151.585 91.860 151.875 91.905 ;
        RECT 149.270 91.720 151.875 91.860 ;
        RECT 149.270 91.660 149.590 91.720 ;
        RECT 151.585 91.675 151.875 91.720 ;
        RECT 117.085 91.520 117.375 91.565 ;
        RECT 117.990 91.520 118.310 91.580 ;
        RECT 143.790 91.520 144.080 91.565 ;
        RECT 145.890 91.520 146.180 91.565 ;
        RECT 147.460 91.520 147.750 91.565 ;
        RECT 113.940 91.380 114.540 91.520 ;
        RECT 109.710 91.320 110.030 91.380 ;
        RECT 113.405 91.335 113.695 91.380 ;
        RECT 113.850 91.180 114.170 91.240 ;
        RECT 109.340 91.040 114.170 91.180 ;
        RECT 114.400 91.180 114.540 91.380 ;
        RECT 117.085 91.380 118.310 91.520 ;
        RECT 117.085 91.335 117.375 91.380 ;
        RECT 117.990 91.320 118.310 91.380 ;
        RECT 118.540 91.380 130.410 91.520 ;
        RECT 118.540 91.180 118.680 91.380 ;
        RECT 114.400 91.040 118.680 91.180 ;
        RECT 126.820 91.040 129.260 91.180 ;
        RECT 109.340 90.885 109.480 91.040 ;
        RECT 113.850 90.980 114.170 91.040 ;
        RECT 106.505 90.655 106.795 90.885 ;
        RECT 109.265 90.655 109.555 90.885 ;
        RECT 103.270 90.500 103.590 90.560 ;
        RECT 106.580 90.500 106.720 90.655 ;
        RECT 110.630 90.640 110.950 90.900 ;
        RECT 111.090 90.640 111.410 90.900 ;
        RECT 112.025 90.655 112.315 90.885 ;
        RECT 118.450 90.840 118.770 90.900 ;
        RECT 114.860 90.700 118.770 90.840 ;
        RECT 103.270 90.360 106.720 90.500 ;
        RECT 108.790 90.500 109.110 90.560 ;
        RECT 112.100 90.500 112.240 90.655 ;
        RECT 114.860 90.500 115.000 90.700 ;
        RECT 118.450 90.640 118.770 90.700 ;
        RECT 119.830 90.640 120.150 90.900 ;
        RECT 120.290 90.840 120.610 90.900 ;
        RECT 126.820 90.885 126.960 91.040 ;
        RECT 120.765 90.840 121.055 90.885 ;
        RECT 120.290 90.700 121.055 90.840 ;
        RECT 120.290 90.640 120.610 90.700 ;
        RECT 120.765 90.655 121.055 90.700 ;
        RECT 126.745 90.655 127.035 90.885 ;
        RECT 127.205 90.840 127.495 90.885 ;
        RECT 129.120 90.840 129.260 91.040 ;
        RECT 129.490 90.980 129.810 91.240 ;
        RECT 130.270 91.180 130.410 91.380 ;
        RECT 143.790 91.380 147.750 91.520 ;
        RECT 143.790 91.335 144.080 91.380 ;
        RECT 145.890 91.335 146.180 91.380 ;
        RECT 147.460 91.335 147.750 91.380 ;
        RECT 130.885 91.180 131.175 91.225 ;
        RECT 130.270 91.040 131.175 91.180 ;
        RECT 130.885 90.995 131.175 91.040 ;
        RECT 144.185 91.180 144.475 91.225 ;
        RECT 145.375 91.180 145.665 91.225 ;
        RECT 147.895 91.180 148.185 91.225 ;
        RECT 144.185 91.040 148.185 91.180 ;
        RECT 144.185 90.995 144.475 91.040 ;
        RECT 145.375 90.995 145.665 91.040 ;
        RECT 147.895 90.995 148.185 91.040 ;
        RECT 154.330 90.980 154.650 91.240 ;
        RECT 129.950 90.840 130.270 90.900 ;
        RECT 127.205 90.700 128.800 90.840 ;
        RECT 129.120 90.700 130.270 90.840 ;
        RECT 127.205 90.655 127.495 90.700 ;
        RECT 108.790 90.360 112.240 90.500 ;
        RECT 113.940 90.360 115.000 90.500 ;
        RECT 115.230 90.500 115.550 90.560 ;
        RECT 125.810 90.500 126.130 90.560 ;
        RECT 115.230 90.360 126.130 90.500 ;
        RECT 103.270 90.300 103.590 90.360 ;
        RECT 108.790 90.300 109.110 90.360 ;
        RECT 78.430 90.020 84.180 90.160 ;
        RECT 85.330 90.160 85.650 90.220 ;
        RECT 87.645 90.160 87.935 90.205 ;
        RECT 85.330 90.020 87.935 90.160 ;
        RECT 78.430 89.960 78.750 90.020 ;
        RECT 85.330 89.960 85.650 90.020 ;
        RECT 87.645 89.975 87.935 90.020 ;
        RECT 100.970 89.960 101.290 90.220 ;
        RECT 110.185 90.160 110.475 90.205 ;
        RECT 113.940 90.160 114.080 90.360 ;
        RECT 115.230 90.300 115.550 90.360 ;
        RECT 125.810 90.300 126.130 90.360 ;
        RECT 128.125 90.315 128.415 90.545 ;
        RECT 128.660 90.500 128.800 90.700 ;
        RECT 129.950 90.640 130.270 90.700 ;
        RECT 130.425 90.840 130.715 90.885 ;
        RECT 135.010 90.840 135.330 90.900 ;
        RECT 135.945 90.840 136.235 90.885 ;
        RECT 130.425 90.700 136.235 90.840 ;
        RECT 130.425 90.655 130.715 90.700 ;
        RECT 130.500 90.500 130.640 90.655 ;
        RECT 135.010 90.640 135.330 90.700 ;
        RECT 135.945 90.655 136.235 90.700 ;
        RECT 136.390 90.640 136.710 90.900 ;
        RECT 137.325 90.655 137.615 90.885 ;
        RECT 128.660 90.360 130.640 90.500 ;
        RECT 137.400 90.500 137.540 90.655 ;
        RECT 137.770 90.640 138.090 90.900 ;
        RECT 141.925 90.840 142.215 90.885 ;
        RECT 142.830 90.840 143.150 90.900 ;
        RECT 141.925 90.700 143.150 90.840 ;
        RECT 141.925 90.655 142.215 90.700 ;
        RECT 142.830 90.640 143.150 90.700 ;
        RECT 143.305 90.840 143.595 90.885 ;
        RECT 143.305 90.700 145.360 90.840 ;
        RECT 143.305 90.655 143.595 90.700 ;
        RECT 145.220 90.560 145.360 90.700 ;
        RECT 138.690 90.500 139.010 90.560 ;
        RECT 144.530 90.500 144.820 90.545 ;
        RECT 137.400 90.360 139.010 90.500 ;
        RECT 110.185 90.020 114.080 90.160 ;
        RECT 114.245 90.160 114.535 90.205 ;
        RECT 117.530 90.160 117.850 90.220 ;
        RECT 114.245 90.020 117.850 90.160 ;
        RECT 128.200 90.160 128.340 90.315 ;
        RECT 138.690 90.300 139.010 90.360 ;
        RECT 142.920 90.360 144.820 90.500 ;
        RECT 129.490 90.160 129.810 90.220 ;
        RECT 128.200 90.020 129.810 90.160 ;
        RECT 110.185 89.975 110.475 90.020 ;
        RECT 114.245 89.975 114.535 90.020 ;
        RECT 117.530 89.960 117.850 90.020 ;
        RECT 129.490 89.960 129.810 90.020 ;
        RECT 132.710 90.160 133.030 90.220 ;
        RECT 142.920 90.205 143.060 90.360 ;
        RECT 144.530 90.315 144.820 90.360 ;
        RECT 145.130 90.300 145.450 90.560 ;
        RECT 135.025 90.160 135.315 90.205 ;
        RECT 132.710 90.020 135.315 90.160 ;
        RECT 132.710 89.960 133.030 90.020 ;
        RECT 135.025 89.975 135.315 90.020 ;
        RECT 142.845 89.975 143.135 90.205 ;
        RECT 150.190 89.960 150.510 90.220 ;
        RECT 22.700 89.340 157.820 89.820 ;
        RECT 30.590 88.940 30.910 89.200 ;
        RECT 49.450 89.140 49.770 89.200 ;
        RECT 49.925 89.140 50.215 89.185 ;
        RECT 54.050 89.140 54.370 89.200 ;
        RECT 49.450 89.000 50.215 89.140 ;
        RECT 49.450 88.940 49.770 89.000 ;
        RECT 49.925 88.955 50.215 89.000 ;
        RECT 50.920 89.000 54.370 89.140 ;
        RECT 31.985 88.800 32.275 88.845 ;
        RECT 32.890 88.800 33.210 88.860 ;
        RECT 31.985 88.660 35.420 88.800 ;
        RECT 31.985 88.615 32.275 88.660 ;
        RECT 32.890 88.600 33.210 88.660 ;
        RECT 30.145 88.460 30.435 88.505 ;
        RECT 30.590 88.460 30.910 88.520 ;
        RECT 30.145 88.320 30.910 88.460 ;
        RECT 30.145 88.275 30.435 88.320 ;
        RECT 30.590 88.260 30.910 88.320 ;
        RECT 31.050 88.460 31.370 88.520 ;
        RECT 31.525 88.460 31.815 88.505 ;
        RECT 31.050 88.320 31.815 88.460 ;
        RECT 31.050 88.260 31.370 88.320 ;
        RECT 31.525 88.275 31.815 88.320 ;
        RECT 32.445 88.275 32.735 88.505 ;
        RECT 34.185 88.460 34.475 88.505 ;
        RECT 34.185 88.275 34.500 88.460 ;
        RECT 30.680 88.120 30.820 88.260 ;
        RECT 32.520 88.120 32.660 88.275 ;
        RECT 30.680 87.980 32.660 88.120 ;
        RECT 32.905 88.120 33.195 88.165 ;
        RECT 33.350 88.120 33.670 88.180 ;
        RECT 32.905 87.980 33.670 88.120 ;
        RECT 34.360 88.120 34.500 88.275 ;
        RECT 34.730 88.260 35.050 88.520 ;
        RECT 35.280 88.505 35.420 88.660 ;
        RECT 36.570 88.600 36.890 88.860 ;
        RECT 42.565 88.615 42.855 88.845 ;
        RECT 35.205 88.275 35.495 88.505 ;
        RECT 36.110 88.460 36.430 88.520 ;
        RECT 37.505 88.460 37.795 88.505 ;
        RECT 36.110 88.320 37.795 88.460 ;
        RECT 36.110 88.260 36.430 88.320 ;
        RECT 37.505 88.275 37.795 88.320 ;
        RECT 37.950 88.260 38.270 88.520 ;
        RECT 41.170 88.460 41.490 88.520 ;
        RECT 42.640 88.460 42.780 88.615 ;
        RECT 41.170 88.320 42.780 88.460 ;
        RECT 41.170 88.260 41.490 88.320 ;
        RECT 44.390 88.260 44.710 88.520 ;
        RECT 44.850 88.260 45.170 88.520 ;
        RECT 45.310 88.260 45.630 88.520 ;
        RECT 46.230 88.260 46.550 88.520 ;
        RECT 49.910 88.460 50.230 88.520 ;
        RECT 50.920 88.505 51.060 89.000 ;
        RECT 54.050 88.940 54.370 89.000 ;
        RECT 54.510 89.140 54.830 89.200 ;
        RECT 57.285 89.140 57.575 89.185 ;
        RECT 54.510 89.000 57.575 89.140 ;
        RECT 54.510 88.940 54.830 89.000 ;
        RECT 57.285 88.955 57.575 89.000 ;
        RECT 58.190 88.940 58.510 89.200 ;
        RECT 78.430 89.140 78.750 89.200 ;
        RECT 58.740 89.000 78.750 89.140 ;
        RECT 54.600 88.800 54.740 88.940 ;
        RECT 52.760 88.660 54.740 88.800 ;
        RECT 54.970 88.800 55.290 88.860 ;
        RECT 58.740 88.800 58.880 89.000 ;
        RECT 78.430 88.940 78.750 89.000 ;
        RECT 82.570 89.140 82.890 89.200 ;
        RECT 83.965 89.140 84.255 89.185 ;
        RECT 82.570 89.000 84.255 89.140 ;
        RECT 82.570 88.940 82.890 89.000 ;
        RECT 83.965 88.955 84.255 89.000 ;
        RECT 86.710 89.140 87.030 89.200 ;
        RECT 88.105 89.140 88.395 89.185 ;
        RECT 86.710 89.000 88.395 89.140 ;
        RECT 86.710 88.940 87.030 89.000 ;
        RECT 88.105 88.955 88.395 89.000 ;
        RECT 100.970 89.140 101.290 89.200 ;
        RECT 102.365 89.140 102.655 89.185 ;
        RECT 115.230 89.140 115.550 89.200 ;
        RECT 100.970 89.000 102.655 89.140 ;
        RECT 100.970 88.940 101.290 89.000 ;
        RECT 102.365 88.955 102.655 89.000 ;
        RECT 104.280 89.000 115.550 89.140 ;
        RECT 54.970 88.660 58.880 88.800 ;
        RECT 63.250 88.800 63.570 88.860 ;
        RECT 76.100 88.800 76.390 88.845 ;
        RECT 76.590 88.800 76.910 88.860 ;
        RECT 104.280 88.800 104.420 89.000 ;
        RECT 115.230 88.940 115.550 89.000 ;
        RECT 117.990 88.940 118.310 89.200 ;
        RECT 118.450 89.140 118.770 89.200 ;
        RECT 120.765 89.140 121.055 89.185 ;
        RECT 118.450 89.000 121.055 89.140 ;
        RECT 118.450 88.940 118.770 89.000 ;
        RECT 120.765 88.955 121.055 89.000 ;
        RECT 142.370 89.140 142.690 89.200 ;
        RECT 152.030 89.140 152.350 89.200 ;
        RECT 142.370 89.000 148.120 89.140 ;
        RECT 142.370 88.940 142.690 89.000 ;
        RECT 106.045 88.800 106.335 88.845 ;
        RECT 63.250 88.660 75.900 88.800 ;
        RECT 50.845 88.460 51.135 88.505 ;
        RECT 49.910 88.320 51.135 88.460 ;
        RECT 49.910 88.260 50.230 88.320 ;
        RECT 50.845 88.275 51.135 88.320 ;
        RECT 51.305 88.275 51.595 88.505 ;
        RECT 42.105 88.120 42.395 88.165 ;
        RECT 43.010 88.120 43.330 88.180 ;
        RECT 34.360 87.980 37.720 88.120 ;
        RECT 32.905 87.935 33.195 87.980 ;
        RECT 33.350 87.920 33.670 87.980 ;
        RECT 35.650 87.780 35.970 87.840 ;
        RECT 36.585 87.780 36.875 87.825 ;
        RECT 35.650 87.640 36.875 87.780 ;
        RECT 35.650 87.580 35.970 87.640 ;
        RECT 36.585 87.595 36.875 87.640 ;
        RECT 37.580 87.500 37.720 87.980 ;
        RECT 42.105 87.980 43.330 88.120 ;
        RECT 42.105 87.935 42.395 87.980 ;
        RECT 43.010 87.920 43.330 87.980 ;
        RECT 43.485 88.120 43.775 88.165 ;
        RECT 43.930 88.120 44.250 88.180 ;
        RECT 47.165 88.120 47.455 88.165 ;
        RECT 43.485 87.980 47.455 88.120 ;
        RECT 51.380 88.120 51.520 88.275 ;
        RECT 52.210 88.260 52.530 88.520 ;
        RECT 52.760 88.505 52.900 88.660 ;
        RECT 54.970 88.600 55.290 88.660 ;
        RECT 63.250 88.600 63.570 88.660 ;
        RECT 52.685 88.275 52.975 88.505 ;
        RECT 53.130 88.260 53.450 88.520 ;
        RECT 54.050 88.260 54.370 88.520 ;
        RECT 66.470 88.460 66.790 88.520 ;
        RECT 74.765 88.460 75.055 88.505 ;
        RECT 66.470 88.320 75.055 88.460 ;
        RECT 75.760 88.460 75.900 88.660 ;
        RECT 76.100 88.660 76.910 88.800 ;
        RECT 76.100 88.615 76.390 88.660 ;
        RECT 76.590 88.600 76.910 88.660 ;
        RECT 77.140 88.660 104.420 88.800 ;
        RECT 104.740 88.660 106.335 88.800 ;
        RECT 77.140 88.460 77.280 88.660 ;
        RECT 104.740 88.520 104.880 88.660 ;
        RECT 106.045 88.615 106.335 88.660 ;
        RECT 108.330 88.800 108.650 88.860 ;
        RECT 125.810 88.800 126.130 88.860 ;
        RECT 126.745 88.800 127.035 88.845 ;
        RECT 127.190 88.800 127.510 88.860 ;
        RECT 108.330 88.660 110.860 88.800 ;
        RECT 108.330 88.600 108.650 88.660 ;
        RECT 75.760 88.320 77.280 88.460 ;
        RECT 77.510 88.460 77.830 88.520 ;
        RECT 82.125 88.460 82.415 88.505 ;
        RECT 77.510 88.320 82.415 88.460 ;
        RECT 66.470 88.260 66.790 88.320 ;
        RECT 74.765 88.275 75.055 88.320 ;
        RECT 77.510 88.260 77.830 88.320 ;
        RECT 82.125 88.275 82.415 88.320 ;
        RECT 82.570 88.460 82.890 88.520 ;
        RECT 83.045 88.460 83.335 88.505 ;
        RECT 82.570 88.320 83.335 88.460 ;
        RECT 82.570 88.260 82.890 88.320 ;
        RECT 83.045 88.275 83.335 88.320 ;
        RECT 85.330 88.260 85.650 88.520 ;
        RECT 87.645 88.275 87.935 88.505 ;
        RECT 88.565 88.460 88.855 88.505 ;
        RECT 90.850 88.460 91.170 88.520 ;
        RECT 88.565 88.320 91.170 88.460 ;
        RECT 88.565 88.275 88.855 88.320 ;
        RECT 53.590 88.120 53.910 88.180 ;
        RECT 54.985 88.120 55.275 88.165 ;
        RECT 51.380 87.980 55.275 88.120 ;
        RECT 43.485 87.935 43.775 87.980 ;
        RECT 43.930 87.920 44.250 87.980 ;
        RECT 47.165 87.935 47.455 87.980 ;
        RECT 53.590 87.920 53.910 87.980 ;
        RECT 54.985 87.935 55.275 87.980 ;
        RECT 75.645 88.120 75.935 88.165 ;
        RECT 76.835 88.120 77.125 88.165 ;
        RECT 79.355 88.120 79.645 88.165 ;
        RECT 75.645 87.980 79.645 88.120 ;
        RECT 75.645 87.935 75.935 87.980 ;
        RECT 76.835 87.935 77.125 87.980 ;
        RECT 79.355 87.935 79.645 87.980 ;
        RECT 80.730 88.120 81.050 88.180 ;
        RECT 81.650 88.120 81.970 88.180 ;
        RECT 87.720 88.120 87.860 88.275 ;
        RECT 90.850 88.260 91.170 88.320 ;
        RECT 103.270 88.260 103.590 88.520 ;
        RECT 103.745 88.275 104.035 88.505 ;
        RECT 80.730 87.980 87.860 88.120 ;
        RECT 103.820 88.120 103.960 88.275 ;
        RECT 104.650 88.260 104.970 88.520 ;
        RECT 105.110 88.260 105.430 88.520 ;
        RECT 106.505 88.460 106.795 88.505 ;
        RECT 107.885 88.460 108.175 88.505 ;
        RECT 106.505 88.320 107.640 88.460 ;
        RECT 106.505 88.275 106.795 88.320 ;
        RECT 105.570 88.120 105.890 88.180 ;
        RECT 106.965 88.120 107.255 88.165 ;
        RECT 103.820 87.980 107.255 88.120 ;
        RECT 107.500 88.120 107.640 88.320 ;
        RECT 107.885 88.320 108.560 88.460 ;
        RECT 107.885 88.275 108.175 88.320 ;
        RECT 108.420 88.180 108.560 88.320 ;
        RECT 108.790 88.260 109.110 88.520 ;
        RECT 109.265 88.460 109.555 88.505 ;
        RECT 109.710 88.460 110.030 88.520 ;
        RECT 109.265 88.320 110.030 88.460 ;
        RECT 109.265 88.275 109.555 88.320 ;
        RECT 109.710 88.260 110.030 88.320 ;
        RECT 110.720 88.180 110.860 88.660 ;
        RECT 119.460 88.660 120.980 88.800 ;
        RECT 112.010 88.505 112.330 88.520 ;
        RECT 111.925 88.275 112.330 88.505 ;
        RECT 118.925 88.460 119.215 88.505 ;
        RECT 119.460 88.460 119.600 88.660 ;
        RECT 118.925 88.320 119.600 88.460 ;
        RECT 119.845 88.460 120.135 88.505 ;
        RECT 120.305 88.460 120.595 88.505 ;
        RECT 119.845 88.320 120.595 88.460 ;
        RECT 120.840 88.460 120.980 88.660 ;
        RECT 125.810 88.660 127.510 88.800 ;
        RECT 125.810 88.600 126.130 88.660 ;
        RECT 126.745 88.615 127.035 88.660 ;
        RECT 127.190 88.600 127.510 88.660 ;
        RECT 127.825 88.800 128.115 88.845 ;
        RECT 129.950 88.800 130.270 88.860 ;
        RECT 146.510 88.800 146.830 88.860 ;
        RECT 127.825 88.660 130.410 88.800 ;
        RECT 127.825 88.615 128.115 88.660 ;
        RECT 129.950 88.600 130.410 88.660 ;
        RECT 121.210 88.460 121.530 88.520 ;
        RECT 120.840 88.320 121.530 88.460 ;
        RECT 130.270 88.460 130.410 88.600 ;
        RECT 142.920 88.660 147.660 88.800 ;
        RECT 135.485 88.460 135.775 88.505 ;
        RECT 130.270 88.320 135.775 88.460 ;
        RECT 118.925 88.275 119.215 88.320 ;
        RECT 119.845 88.275 120.135 88.320 ;
        RECT 120.305 88.275 120.595 88.320 ;
        RECT 112.010 88.260 112.330 88.275 ;
        RECT 108.330 88.120 108.650 88.180 ;
        RECT 110.170 88.120 110.490 88.180 ;
        RECT 107.500 87.980 108.100 88.120 ;
        RECT 80.730 87.920 81.050 87.980 ;
        RECT 81.650 87.920 81.970 87.980 ;
        RECT 105.570 87.920 105.890 87.980 ;
        RECT 106.965 87.935 107.255 87.980 ;
        RECT 107.960 87.840 108.100 87.980 ;
        RECT 108.330 87.980 110.490 88.120 ;
        RECT 108.330 87.920 108.650 87.980 ;
        RECT 110.170 87.920 110.490 87.980 ;
        RECT 110.630 87.920 110.950 88.180 ;
        RECT 111.525 88.120 111.815 88.165 ;
        RECT 112.715 88.120 113.005 88.165 ;
        RECT 115.235 88.120 115.525 88.165 ;
        RECT 119.920 88.120 120.060 88.275 ;
        RECT 121.210 88.260 121.530 88.320 ;
        RECT 135.485 88.275 135.775 88.320 ;
        RECT 136.390 88.260 136.710 88.520 ;
        RECT 137.770 88.260 138.090 88.520 ;
        RECT 138.690 88.460 139.010 88.520 ;
        RECT 140.545 88.460 140.835 88.505 ;
        RECT 138.690 88.320 140.835 88.460 ;
        RECT 138.690 88.260 139.010 88.320 ;
        RECT 140.545 88.275 140.835 88.320 ;
        RECT 141.005 88.460 141.295 88.505 ;
        RECT 142.920 88.460 143.060 88.660 ;
        RECT 141.005 88.320 143.060 88.460 ;
        RECT 141.005 88.275 141.295 88.320 ;
        RECT 143.305 88.275 143.595 88.505 ;
        RECT 111.525 87.980 115.525 88.120 ;
        RECT 111.525 87.935 111.815 87.980 ;
        RECT 112.715 87.935 113.005 87.980 ;
        RECT 115.235 87.935 115.525 87.980 ;
        RECT 117.620 87.980 120.060 88.120 ;
        RECT 137.860 88.120 138.000 88.260 ;
        RECT 141.925 88.120 142.215 88.165 ;
        RECT 137.860 87.980 142.215 88.120 ;
        RECT 143.380 88.120 143.520 88.275 ;
        RECT 143.750 88.260 144.070 88.520 ;
        RECT 144.225 88.275 144.515 88.505 ;
        RECT 144.760 88.460 144.900 88.660 ;
        RECT 146.510 88.600 146.830 88.660 ;
        RECT 145.145 88.460 145.435 88.505 ;
        RECT 144.760 88.320 145.435 88.460 ;
        RECT 145.145 88.275 145.435 88.320 ;
        RECT 144.300 88.120 144.440 88.275 ;
        RECT 145.590 88.260 145.910 88.520 ;
        RECT 146.050 88.260 146.370 88.520 ;
        RECT 146.970 88.260 147.290 88.520 ;
        RECT 147.520 88.505 147.660 88.660 ;
        RECT 147.445 88.275 147.735 88.505 ;
        RECT 147.980 88.460 148.120 89.000 ;
        RECT 152.030 89.000 153.180 89.140 ;
        RECT 152.030 88.940 152.350 89.000 ;
        RECT 153.040 88.845 153.180 89.000 ;
        RECT 152.965 88.615 153.255 88.845 ;
        RECT 148.825 88.460 149.115 88.505 ;
        RECT 147.980 88.320 149.115 88.460 ;
        RECT 148.825 88.275 149.115 88.320 ;
        RECT 147.060 88.120 147.200 88.260 ;
        RECT 143.380 87.980 143.980 88.120 ;
        RECT 144.300 87.980 147.200 88.120 ;
        RECT 148.900 88.120 149.040 88.275 ;
        RECT 149.730 88.260 150.050 88.520 ;
        RECT 150.650 88.260 150.970 88.520 ;
        RECT 152.045 88.275 152.335 88.505 ;
        RECT 152.120 88.120 152.260 88.275 ;
        RECT 153.870 88.260 154.190 88.520 ;
        RECT 148.900 87.980 152.260 88.120 ;
        RECT 59.110 87.780 59.430 87.840 ;
        RECT 60.045 87.780 60.335 87.825 ;
        RECT 59.110 87.640 60.335 87.780 ;
        RECT 59.110 87.580 59.430 87.640 ;
        RECT 60.045 87.595 60.335 87.640 ;
        RECT 75.250 87.780 75.540 87.825 ;
        RECT 77.350 87.780 77.640 87.825 ;
        RECT 78.920 87.780 79.210 87.825 ;
        RECT 93.150 87.780 93.470 87.840 ;
        RECT 75.250 87.640 79.210 87.780 ;
        RECT 75.250 87.595 75.540 87.640 ;
        RECT 77.350 87.595 77.640 87.640 ;
        RECT 78.920 87.595 79.210 87.640 ;
        RECT 81.280 87.640 93.470 87.780 ;
        RECT 37.490 87.440 37.810 87.500 ;
        RECT 40.265 87.440 40.555 87.485 ;
        RECT 37.490 87.300 40.555 87.440 ;
        RECT 37.490 87.240 37.810 87.300 ;
        RECT 40.265 87.255 40.555 87.300 ;
        RECT 58.205 87.440 58.495 87.485 ;
        RECT 58.650 87.440 58.970 87.500 ;
        RECT 58.205 87.300 58.970 87.440 ;
        RECT 58.205 87.255 58.495 87.300 ;
        RECT 58.650 87.240 58.970 87.300 ;
        RECT 65.090 87.440 65.410 87.500 ;
        RECT 81.280 87.440 81.420 87.640 ;
        RECT 93.150 87.580 93.470 87.640 ;
        RECT 107.870 87.580 108.190 87.840 ;
        RECT 117.620 87.825 117.760 87.980 ;
        RECT 141.925 87.935 142.215 87.980 ;
        RECT 111.130 87.780 111.420 87.825 ;
        RECT 113.230 87.780 113.520 87.825 ;
        RECT 114.800 87.780 115.090 87.825 ;
        RECT 111.130 87.640 115.090 87.780 ;
        RECT 111.130 87.595 111.420 87.640 ;
        RECT 113.230 87.595 113.520 87.640 ;
        RECT 114.800 87.595 115.090 87.640 ;
        RECT 117.545 87.595 117.835 87.825 ;
        RECT 132.710 87.780 133.030 87.840 ;
        RECT 127.740 87.640 133.030 87.780 ;
        RECT 65.090 87.300 81.420 87.440 ;
        RECT 65.090 87.240 65.410 87.300 ;
        RECT 81.650 87.240 81.970 87.500 ;
        RECT 86.250 87.240 86.570 87.500 ;
        RECT 110.185 87.440 110.475 87.485 ;
        RECT 112.010 87.440 112.330 87.500 ;
        RECT 127.740 87.485 127.880 87.640 ;
        RECT 132.710 87.580 133.030 87.640 ;
        RECT 135.010 87.580 135.330 87.840 ;
        RECT 143.840 87.780 143.980 87.980 ;
        RECT 146.050 87.780 146.370 87.840 ;
        RECT 143.840 87.640 146.370 87.780 ;
        RECT 146.050 87.580 146.370 87.640 ;
        RECT 110.185 87.300 112.330 87.440 ;
        RECT 110.185 87.255 110.475 87.300 ;
        RECT 112.010 87.240 112.330 87.300 ;
        RECT 127.665 87.255 127.955 87.485 ;
        RECT 128.110 87.440 128.430 87.500 ;
        RECT 128.585 87.440 128.875 87.485 ;
        RECT 128.110 87.300 128.875 87.440 ;
        RECT 128.110 87.240 128.430 87.300 ;
        RECT 128.585 87.255 128.875 87.300 ;
        RECT 143.750 87.440 144.070 87.500 ;
        RECT 145.590 87.440 145.910 87.500 ;
        RECT 143.750 87.300 145.910 87.440 ;
        RECT 143.750 87.240 144.070 87.300 ;
        RECT 145.590 87.240 145.910 87.300 ;
        RECT 148.350 87.240 148.670 87.500 ;
        RECT 22.700 86.620 157.020 87.100 ;
        RECT 34.745 86.420 35.035 86.465 ;
        RECT 39.345 86.420 39.635 86.465 ;
        RECT 34.745 86.280 39.635 86.420 ;
        RECT 34.745 86.235 35.035 86.280 ;
        RECT 39.345 86.235 39.635 86.280 ;
        RECT 43.010 86.420 43.330 86.480 ;
        RECT 43.485 86.420 43.775 86.465 ;
        RECT 43.010 86.280 43.775 86.420 ;
        RECT 43.010 86.220 43.330 86.280 ;
        RECT 43.485 86.235 43.775 86.280 ;
        RECT 49.910 86.220 50.230 86.480 ;
        RECT 57.285 86.420 57.575 86.465 ;
        RECT 58.665 86.420 58.955 86.465 ;
        RECT 57.285 86.280 58.955 86.420 ;
        RECT 57.285 86.235 57.575 86.280 ;
        RECT 58.665 86.235 58.955 86.280 ;
        RECT 65.565 86.420 65.855 86.465 ;
        RECT 66.945 86.420 67.235 86.465 ;
        RECT 65.565 86.280 67.235 86.420 ;
        RECT 65.565 86.235 65.855 86.280 ;
        RECT 66.945 86.235 67.235 86.280 ;
        RECT 69.690 86.420 70.010 86.480 ;
        RECT 77.510 86.420 77.830 86.480 ;
        RECT 69.690 86.280 77.830 86.420 ;
        RECT 69.690 86.220 70.010 86.280 ;
        RECT 77.510 86.220 77.830 86.280 ;
        RECT 80.360 86.280 81.880 86.420 ;
        RECT 37.950 85.880 38.270 86.140 ;
        RECT 46.230 86.080 46.550 86.140 ;
        RECT 43.560 85.940 46.550 86.080 ;
        RECT 34.360 85.600 37.260 85.740 ;
        RECT 34.360 85.445 34.500 85.600 ;
        RECT 37.120 85.445 37.260 85.600 ;
        RECT 43.560 85.460 43.700 85.940 ;
        RECT 46.230 85.880 46.550 85.940 ;
        RECT 66.010 86.080 66.330 86.140 ;
        RECT 66.485 86.080 66.775 86.125 ;
        RECT 71.530 86.080 71.850 86.140 ;
        RECT 79.825 86.080 80.115 86.125 ;
        RECT 66.010 85.940 66.775 86.080 ;
        RECT 66.010 85.880 66.330 85.940 ;
        RECT 66.485 85.895 66.775 85.940 ;
        RECT 67.940 85.940 71.850 86.080 ;
        RECT 45.310 85.740 45.630 85.800 ;
        RECT 54.050 85.740 54.370 85.800 ;
        RECT 44.020 85.600 45.630 85.740 ;
        RECT 34.285 85.215 34.575 85.445 ;
        RECT 35.205 85.400 35.495 85.445 ;
        RECT 36.125 85.400 36.415 85.445 ;
        RECT 34.820 85.260 36.415 85.400 ;
        RECT 34.820 85.120 34.960 85.260 ;
        RECT 35.205 85.215 35.495 85.260 ;
        RECT 36.125 85.215 36.415 85.260 ;
        RECT 37.045 85.400 37.335 85.445 ;
        RECT 37.490 85.400 37.810 85.460 ;
        RECT 37.045 85.260 37.810 85.400 ;
        RECT 37.045 85.215 37.335 85.260 ;
        RECT 37.490 85.200 37.810 85.260 ;
        RECT 41.645 85.400 41.935 85.445 ;
        RECT 42.550 85.400 42.870 85.460 ;
        RECT 41.645 85.260 42.870 85.400 ;
        RECT 41.645 85.215 41.935 85.260 ;
        RECT 42.550 85.200 42.870 85.260 ;
        RECT 43.025 85.400 43.315 85.445 ;
        RECT 43.470 85.400 43.790 85.460 ;
        RECT 44.020 85.445 44.160 85.600 ;
        RECT 45.310 85.540 45.630 85.600 ;
        RECT 49.540 85.600 54.370 85.740 ;
        RECT 43.025 85.260 43.790 85.400 ;
        RECT 43.025 85.215 43.315 85.260 ;
        RECT 43.470 85.200 43.790 85.260 ;
        RECT 43.945 85.215 44.235 85.445 ;
        RECT 44.390 85.200 44.710 85.460 ;
        RECT 48.070 85.400 48.390 85.460 ;
        RECT 49.540 85.445 49.680 85.600 ;
        RECT 54.050 85.540 54.370 85.600 ;
        RECT 49.465 85.400 49.755 85.445 ;
        RECT 48.070 85.260 49.755 85.400 ;
        RECT 48.070 85.200 48.390 85.260 ;
        RECT 49.465 85.215 49.755 85.260 ;
        RECT 50.385 85.215 50.675 85.445 ;
        RECT 50.830 85.400 51.150 85.460 ;
        RECT 51.765 85.400 52.055 85.445 ;
        RECT 50.830 85.260 52.055 85.400 ;
        RECT 34.730 84.860 35.050 85.120 ;
        RECT 37.950 85.060 38.270 85.120 ;
        RECT 39.185 85.060 39.475 85.105 ;
        RECT 37.950 84.920 39.475 85.060 ;
        RECT 37.950 84.860 38.270 84.920 ;
        RECT 39.185 84.875 39.475 84.920 ;
        RECT 40.250 84.860 40.570 85.120 ;
        RECT 50.460 85.060 50.600 85.215 ;
        RECT 50.830 85.200 51.150 85.260 ;
        RECT 51.765 85.215 52.055 85.260 ;
        RECT 55.445 85.400 55.735 85.445 ;
        RECT 57.270 85.400 57.590 85.460 ;
        RECT 55.445 85.260 57.590 85.400 ;
        RECT 55.445 85.215 55.735 85.260 ;
        RECT 57.270 85.200 57.590 85.260 ;
        RECT 60.490 85.400 60.810 85.460 ;
        RECT 65.090 85.400 65.410 85.460 ;
        RECT 67.940 85.445 68.080 85.940 ;
        RECT 71.530 85.880 71.850 85.940 ;
        RECT 73.000 85.940 80.115 86.080 ;
        RECT 68.400 85.600 70.380 85.740 ;
        RECT 68.400 85.445 68.540 85.600 ;
        RECT 70.240 85.460 70.380 85.600 ;
        RECT 60.490 85.260 65.410 85.400 ;
        RECT 60.490 85.200 60.810 85.260 ;
        RECT 52.670 85.060 52.990 85.120 ;
        RECT 50.460 84.920 52.990 85.060 ;
        RECT 52.670 84.860 52.990 84.920 ;
        RECT 54.970 85.060 55.290 85.120 ;
        RECT 56.365 85.060 56.655 85.105 ;
        RECT 54.970 84.920 56.655 85.060 ;
        RECT 54.970 84.860 55.290 84.920 ;
        RECT 56.365 84.875 56.655 84.920 ;
        RECT 57.745 85.060 58.035 85.105 ;
        RECT 63.250 85.060 63.570 85.120 ;
        RECT 64.720 85.105 64.860 85.260 ;
        RECT 65.090 85.200 65.410 85.260 ;
        RECT 67.865 85.215 68.155 85.445 ;
        RECT 68.325 85.215 68.615 85.445 ;
        RECT 69.230 85.200 69.550 85.460 ;
        RECT 69.690 85.200 70.010 85.460 ;
        RECT 70.150 85.200 70.470 85.460 ;
        RECT 71.620 85.445 71.760 85.880 ;
        RECT 71.545 85.400 71.835 85.445 ;
        RECT 72.450 85.400 72.770 85.460 ;
        RECT 73.000 85.445 73.140 85.940 ;
        RECT 79.825 85.895 80.115 85.940 ;
        RECT 80.360 85.740 80.500 86.280 ;
        RECT 81.740 86.140 81.880 86.280 ;
        RECT 82.570 86.220 82.890 86.480 ;
        RECT 100.985 86.420 101.275 86.465 ;
        RECT 101.430 86.420 101.750 86.480 ;
        RECT 100.985 86.280 101.750 86.420 ;
        RECT 100.985 86.235 101.275 86.280 ;
        RECT 101.430 86.220 101.750 86.280 ;
        RECT 136.390 86.420 136.710 86.480 ;
        RECT 137.785 86.420 138.075 86.465 ;
        RECT 136.390 86.280 138.075 86.420 ;
        RECT 136.390 86.220 136.710 86.280 ;
        RECT 137.785 86.235 138.075 86.280 ;
        RECT 141.910 86.220 142.230 86.480 ;
        RECT 142.830 86.220 143.150 86.480 ;
        RECT 146.510 86.220 146.830 86.480 ;
        RECT 146.970 86.420 147.290 86.480 ;
        RECT 148.825 86.420 149.115 86.465 ;
        RECT 146.970 86.280 149.115 86.420 ;
        RECT 146.970 86.220 147.290 86.280 ;
        RECT 148.825 86.235 149.115 86.280 ;
        RECT 81.650 86.080 81.970 86.140 ;
        RECT 82.660 86.080 82.800 86.220 ;
        RECT 90.390 86.080 90.680 86.125 ;
        RECT 91.960 86.080 92.250 86.125 ;
        RECT 94.060 86.080 94.350 86.125 ;
        RECT 81.650 85.880 82.110 86.080 ;
        RECT 82.660 85.940 83.260 86.080 ;
        RECT 78.520 85.600 80.500 85.740 ;
        RECT 81.970 85.740 82.110 85.880 ;
        RECT 81.970 85.600 82.800 85.740 ;
        RECT 71.545 85.260 72.770 85.400 ;
        RECT 71.545 85.215 71.835 85.260 ;
        RECT 72.450 85.200 72.770 85.260 ;
        RECT 72.925 85.215 73.215 85.445 ;
        RECT 74.305 85.400 74.595 85.445 ;
        RECT 77.510 85.400 77.830 85.460 ;
        RECT 78.520 85.445 78.660 85.600 ;
        RECT 74.305 85.260 77.830 85.400 ;
        RECT 74.305 85.215 74.595 85.260 ;
        RECT 57.745 84.920 63.570 85.060 ;
        RECT 57.745 84.875 58.035 84.920 ;
        RECT 38.410 84.520 38.730 84.780 ;
        RECT 40.340 84.720 40.480 84.860 ;
        RECT 57.820 84.720 57.960 84.875 ;
        RECT 63.250 84.860 63.570 84.920 ;
        RECT 64.645 84.875 64.935 85.105 ;
        RECT 65.725 85.060 66.015 85.105 ;
        RECT 66.930 85.060 67.250 85.120 ;
        RECT 70.625 85.060 70.915 85.105 ;
        RECT 65.725 84.920 70.915 85.060 ;
        RECT 65.725 84.875 66.015 84.920 ;
        RECT 66.930 84.860 67.250 84.920 ;
        RECT 70.625 84.875 70.915 84.920 ;
        RECT 40.340 84.580 57.960 84.720 ;
        RECT 58.650 84.765 58.970 84.780 ;
        RECT 58.650 84.535 59.035 84.765 ;
        RECT 58.650 84.520 58.970 84.535 ;
        RECT 59.570 84.520 59.890 84.780 ;
        RECT 69.230 84.720 69.550 84.780 ;
        RECT 73.000 84.720 73.140 85.215 ;
        RECT 77.510 85.200 77.830 85.260 ;
        RECT 78.445 85.215 78.735 85.445 ;
        RECT 78.890 85.200 79.210 85.460 ;
        RECT 81.190 85.200 81.510 85.460 ;
        RECT 81.650 85.200 81.970 85.460 ;
        RECT 82.660 85.445 82.800 85.600 ;
        RECT 82.585 85.215 82.875 85.445 ;
        RECT 79.825 85.060 80.115 85.105 ;
        RECT 83.120 85.060 83.260 85.940 ;
        RECT 90.390 85.940 94.350 86.080 ;
        RECT 90.390 85.895 90.680 85.940 ;
        RECT 91.960 85.895 92.250 85.940 ;
        RECT 94.060 85.895 94.350 85.940 ;
        RECT 98.670 85.880 98.990 86.140 ;
        RECT 129.070 86.080 129.360 86.125 ;
        RECT 131.170 86.080 131.460 86.125 ;
        RECT 132.740 86.080 133.030 86.125 ;
        RECT 129.070 85.940 133.030 86.080 ;
        RECT 129.070 85.895 129.360 85.940 ;
        RECT 131.170 85.895 131.460 85.940 ;
        RECT 132.740 85.895 133.030 85.940 ;
        RECT 86.250 85.740 86.570 85.800 ;
        RECT 89.955 85.740 90.245 85.785 ;
        RECT 92.475 85.740 92.765 85.785 ;
        RECT 93.665 85.740 93.955 85.785 ;
        RECT 86.250 85.600 89.700 85.740 ;
        RECT 86.250 85.540 86.570 85.600 ;
        RECT 85.790 85.200 86.110 85.460 ;
        RECT 86.725 85.400 87.015 85.445 ;
        RECT 89.560 85.400 89.700 85.600 ;
        RECT 89.955 85.600 93.955 85.740 ;
        RECT 89.955 85.555 90.245 85.600 ;
        RECT 92.475 85.555 92.765 85.600 ;
        RECT 93.665 85.555 93.955 85.600 ;
        RECT 94.545 85.740 94.835 85.785 ;
        RECT 98.760 85.740 98.900 85.880 ;
        RECT 94.545 85.600 98.900 85.740 ;
        RECT 126.270 85.740 126.590 85.800 ;
        RECT 128.585 85.740 128.875 85.785 ;
        RECT 126.270 85.600 128.875 85.740 ;
        RECT 94.545 85.555 94.835 85.600 ;
        RECT 126.270 85.540 126.590 85.600 ;
        RECT 128.585 85.555 128.875 85.600 ;
        RECT 129.465 85.740 129.755 85.785 ;
        RECT 130.655 85.740 130.945 85.785 ;
        RECT 133.175 85.740 133.465 85.785 ;
        RECT 129.465 85.600 133.465 85.740 ;
        RECT 129.465 85.555 129.755 85.600 ;
        RECT 130.655 85.555 130.945 85.600 ;
        RECT 133.175 85.555 133.465 85.600 ;
        RECT 137.770 85.740 138.090 85.800 ;
        RECT 140.085 85.740 140.375 85.785 ;
        RECT 149.730 85.740 150.050 85.800 ;
        RECT 137.770 85.600 140.375 85.740 ;
        RECT 137.770 85.540 138.090 85.600 ;
        RECT 140.085 85.555 140.375 85.600 ;
        RECT 146.140 85.600 150.050 85.740 ;
        RECT 93.210 85.400 93.500 85.445 ;
        RECT 97.765 85.400 98.055 85.445 ;
        RECT 86.725 85.260 87.860 85.400 ;
        RECT 89.560 85.260 93.500 85.400 ;
        RECT 86.725 85.215 87.015 85.260 ;
        RECT 79.825 84.920 83.260 85.060 ;
        RECT 79.825 84.875 80.115 84.920 ;
        RECT 87.720 84.780 87.860 85.260 ;
        RECT 93.210 85.215 93.500 85.260 ;
        RECT 96.460 85.260 98.055 85.400 ;
        RECT 96.460 85.120 96.600 85.260 ;
        RECT 97.765 85.215 98.055 85.260 ;
        RECT 98.685 85.215 98.975 85.445 ;
        RECT 102.810 85.400 103.130 85.460 ;
        RECT 105.110 85.400 105.430 85.460 ;
        RECT 102.810 85.260 105.430 85.400 ;
        RECT 96.370 84.860 96.690 85.120 ;
        RECT 97.290 85.060 97.610 85.120 ;
        RECT 98.760 85.060 98.900 85.215 ;
        RECT 102.810 85.200 103.130 85.260 ;
        RECT 105.110 85.200 105.430 85.260 ;
        RECT 105.570 85.400 105.890 85.460 ;
        RECT 106.045 85.400 106.335 85.445 ;
        RECT 105.570 85.260 106.335 85.400 ;
        RECT 105.570 85.200 105.890 85.260 ;
        RECT 106.045 85.215 106.335 85.260 ;
        RECT 106.965 85.400 107.255 85.445 ;
        RECT 109.250 85.400 109.570 85.460 ;
        RECT 106.965 85.260 109.570 85.400 ;
        RECT 106.965 85.215 107.255 85.260 ;
        RECT 97.290 84.920 98.900 85.060 ;
        RECT 106.120 85.060 106.260 85.215 ;
        RECT 109.250 85.200 109.570 85.260 ;
        RECT 127.205 85.400 127.495 85.445 ;
        RECT 128.110 85.400 128.430 85.460 ;
        RECT 127.205 85.260 128.430 85.400 ;
        RECT 127.205 85.215 127.495 85.260 ;
        RECT 128.110 85.200 128.430 85.260 ;
        RECT 134.550 85.400 134.870 85.460 ;
        RECT 136.865 85.400 137.155 85.445 ;
        RECT 134.550 85.260 137.155 85.400 ;
        RECT 134.550 85.200 134.870 85.260 ;
        RECT 136.865 85.215 137.155 85.260 ;
        RECT 145.590 85.400 145.910 85.460 ;
        RECT 146.140 85.445 146.280 85.600 ;
        RECT 149.730 85.540 150.050 85.600 ;
        RECT 146.065 85.400 146.355 85.445 ;
        RECT 145.590 85.260 146.355 85.400 ;
        RECT 145.590 85.200 145.910 85.260 ;
        RECT 146.065 85.215 146.355 85.260 ;
        RECT 146.985 85.400 147.275 85.445 ;
        RECT 150.190 85.400 150.510 85.460 ;
        RECT 150.665 85.400 150.955 85.445 ;
        RECT 146.985 85.260 150.955 85.400 ;
        RECT 146.985 85.215 147.275 85.260 ;
        RECT 150.190 85.200 150.510 85.260 ;
        RECT 150.665 85.215 150.955 85.260 ;
        RECT 108.790 85.060 109.110 85.120 ;
        RECT 129.810 85.060 130.100 85.105 ;
        RECT 106.120 84.920 109.110 85.060 ;
        RECT 97.290 84.860 97.610 84.920 ;
        RECT 108.790 84.860 109.110 84.920 ;
        RECT 128.200 84.920 130.100 85.060 ;
        RECT 69.230 84.580 73.140 84.720 ;
        RECT 80.730 84.720 81.050 84.780 ;
        RECT 85.805 84.720 86.095 84.765 ;
        RECT 80.730 84.580 86.095 84.720 ;
        RECT 69.230 84.520 69.550 84.580 ;
        RECT 80.730 84.520 81.050 84.580 ;
        RECT 85.805 84.535 86.095 84.580 ;
        RECT 87.630 84.520 87.950 84.780 ;
        RECT 95.465 84.720 95.755 84.765 ;
        RECT 95.910 84.720 96.230 84.780 ;
        RECT 95.465 84.580 96.230 84.720 ;
        RECT 95.465 84.535 95.755 84.580 ;
        RECT 95.910 84.520 96.230 84.580 ;
        RECT 97.750 84.520 98.070 84.780 ;
        RECT 100.050 84.520 100.370 84.780 ;
        RECT 100.985 84.720 101.275 84.765 ;
        RECT 102.350 84.720 102.670 84.780 ;
        RECT 100.985 84.580 102.670 84.720 ;
        RECT 100.985 84.535 101.275 84.580 ;
        RECT 102.350 84.520 102.670 84.580 ;
        RECT 106.030 84.720 106.350 84.780 ;
        RECT 107.870 84.720 108.190 84.780 ;
        RECT 128.200 84.765 128.340 84.920 ;
        RECT 129.810 84.875 130.100 84.920 ;
        RECT 135.945 84.875 136.235 85.105 ;
        RECT 141.925 85.060 142.215 85.105 ;
        RECT 148.350 85.060 148.670 85.120 ;
        RECT 141.925 84.920 148.670 85.060 ;
        RECT 141.925 84.875 142.215 84.920 ;
        RECT 106.030 84.580 108.190 84.720 ;
        RECT 106.030 84.520 106.350 84.580 ;
        RECT 107.870 84.520 108.190 84.580 ;
        RECT 128.125 84.535 128.415 84.765 ;
        RECT 135.470 84.720 135.790 84.780 ;
        RECT 136.020 84.720 136.160 84.875 ;
        RECT 148.350 84.860 148.670 84.920 ;
        RECT 149.730 84.860 150.050 85.120 ;
        RECT 135.470 84.580 136.160 84.720 ;
        RECT 135.470 84.520 135.790 84.580 ;
        RECT 22.700 83.900 157.820 84.380 ;
        RECT 37.030 83.700 37.350 83.760 ;
        RECT 37.505 83.700 37.795 83.745 ;
        RECT 37.030 83.560 37.795 83.700 ;
        RECT 37.030 83.500 37.350 83.560 ;
        RECT 37.505 83.515 37.795 83.560 ;
        RECT 44.390 83.500 44.710 83.760 ;
        RECT 48.070 83.500 48.390 83.760 ;
        RECT 69.705 83.515 69.995 83.745 ;
        RECT 38.410 83.360 38.730 83.420 ;
        RECT 44.480 83.360 44.620 83.500 ;
        RECT 66.470 83.360 66.790 83.420 ;
        RECT 32.980 83.220 38.730 83.360 ;
        RECT 32.980 83.065 33.120 83.220 ;
        RECT 38.410 83.160 38.730 83.220 ;
        RECT 43.100 83.220 44.620 83.360 ;
        RECT 62.880 83.220 66.790 83.360 ;
        RECT 69.780 83.360 69.920 83.515 ;
        RECT 70.150 83.500 70.470 83.760 ;
        RECT 72.450 83.500 72.770 83.760 ;
        RECT 78.890 83.700 79.210 83.760 ;
        RECT 81.650 83.700 81.970 83.760 ;
        RECT 78.890 83.560 81.970 83.700 ;
        RECT 78.890 83.500 79.210 83.560 ;
        RECT 81.650 83.500 81.970 83.560 ;
        RECT 85.790 83.700 86.110 83.760 ;
        RECT 85.790 83.560 90.160 83.700 ;
        RECT 85.790 83.500 86.110 83.560 ;
        RECT 72.005 83.360 72.295 83.405 ;
        RECT 87.630 83.360 87.950 83.420 ;
        RECT 90.020 83.405 90.160 83.560 ;
        RECT 90.850 83.500 91.170 83.760 ;
        RECT 91.785 83.700 92.075 83.745 ;
        RECT 97.290 83.700 97.610 83.760 ;
        RECT 91.785 83.560 97.610 83.700 ;
        RECT 91.785 83.515 92.075 83.560 ;
        RECT 97.290 83.500 97.610 83.560 ;
        RECT 102.350 83.500 102.670 83.760 ;
        RECT 105.585 83.700 105.875 83.745 ;
        RECT 102.900 83.560 107.640 83.700 ;
        RECT 89.025 83.360 89.315 83.405 ;
        RECT 69.780 83.220 73.600 83.360 ;
        RECT 32.905 82.835 33.195 83.065 ;
        RECT 35.190 82.820 35.510 83.080 ;
        RECT 36.125 83.020 36.415 83.065 ;
        RECT 40.710 83.020 41.030 83.080 ;
        RECT 36.125 82.880 41.030 83.020 ;
        RECT 36.125 82.835 36.415 82.880 ;
        RECT 40.710 82.820 41.030 82.880 ;
        RECT 41.170 82.820 41.490 83.080 ;
        RECT 42.550 82.820 42.870 83.080 ;
        RECT 43.100 83.065 43.240 83.220 ;
        RECT 43.025 82.835 43.315 83.065 ;
        RECT 44.390 82.820 44.710 83.080 ;
        RECT 49.925 83.020 50.215 83.065 ;
        RECT 50.830 83.020 51.150 83.080 ;
        RECT 49.925 82.880 51.150 83.020 ;
        RECT 49.925 82.835 50.215 82.880 ;
        RECT 50.830 82.820 51.150 82.880 ;
        RECT 51.290 82.820 51.610 83.080 ;
        RECT 60.950 83.065 61.270 83.080 ;
        RECT 62.880 83.065 63.020 83.220 ;
        RECT 66.470 83.160 66.790 83.220 ;
        RECT 72.005 83.175 72.295 83.220 ;
        RECT 64.170 83.065 64.490 83.080 ;
        RECT 60.950 82.835 61.300 83.065 ;
        RECT 62.345 83.020 62.635 83.065 ;
        RECT 62.805 83.020 63.095 83.065 ;
        RECT 62.345 82.880 63.095 83.020 ;
        RECT 62.345 82.835 62.635 82.880 ;
        RECT 62.805 82.835 63.095 82.880 ;
        RECT 64.140 82.835 64.490 83.065 ;
        RECT 60.950 82.820 61.270 82.835 ;
        RECT 64.170 82.820 64.490 82.835 ;
        RECT 70.610 83.020 70.930 83.080 ;
        RECT 73.460 83.065 73.600 83.220 ;
        RECT 87.630 83.220 89.315 83.360 ;
        RECT 87.630 83.160 87.950 83.220 ;
        RECT 89.025 83.175 89.315 83.220 ;
        RECT 89.945 83.360 90.235 83.405 ;
        RECT 92.690 83.360 93.010 83.420 ;
        RECT 89.945 83.220 93.010 83.360 ;
        RECT 89.945 83.175 90.235 83.220 ;
        RECT 92.690 83.160 93.010 83.220 ;
        RECT 97.750 83.360 98.070 83.420 ;
        RECT 102.900 83.360 103.040 83.560 ;
        RECT 105.585 83.515 105.875 83.560 ;
        RECT 106.030 83.360 106.350 83.420 ;
        RECT 106.965 83.360 107.255 83.405 ;
        RECT 97.750 83.220 103.040 83.360 ;
        RECT 103.360 83.220 107.255 83.360 ;
        RECT 97.750 83.160 98.070 83.220 ;
        RECT 97.290 83.065 97.610 83.080 ;
        RECT 71.085 83.020 71.375 83.065 ;
        RECT 72.465 83.020 72.755 83.065 ;
        RECT 70.610 82.880 72.755 83.020 ;
        RECT 70.610 82.820 70.930 82.880 ;
        RECT 71.085 82.835 71.375 82.880 ;
        RECT 72.465 82.835 72.755 82.880 ;
        RECT 73.385 82.835 73.675 83.065 ;
        RECT 97.290 82.835 97.640 83.065 ;
        RECT 100.050 83.020 100.370 83.080 ;
        RECT 103.360 83.065 103.500 83.220 ;
        RECT 106.030 83.160 106.350 83.220 ;
        RECT 106.965 83.175 107.255 83.220 ;
        RECT 100.985 83.020 101.275 83.065 ;
        RECT 100.050 82.880 101.275 83.020 ;
        RECT 97.290 82.820 97.610 82.835 ;
        RECT 100.050 82.820 100.370 82.880 ;
        RECT 100.985 82.835 101.275 82.880 ;
        RECT 103.285 82.835 103.575 83.065 ;
        RECT 39.760 82.680 40.050 82.725 ;
        RECT 42.100 82.680 42.390 82.725 ;
        RECT 39.760 82.540 42.390 82.680 ;
        RECT 39.760 82.495 40.050 82.540 ;
        RECT 42.100 82.495 42.390 82.540 ;
        RECT 43.490 82.680 43.780 82.725 ;
        RECT 45.830 82.680 46.120 82.725 ;
        RECT 43.490 82.540 46.120 82.680 ;
        RECT 43.490 82.495 43.780 82.540 ;
        RECT 45.830 82.495 46.120 82.540 ;
        RECT 50.390 82.680 50.680 82.725 ;
        RECT 52.730 82.680 53.020 82.725 ;
        RECT 50.390 82.540 53.020 82.680 ;
        RECT 50.390 82.495 50.680 82.540 ;
        RECT 52.730 82.495 53.020 82.540 ;
        RECT 57.755 82.680 58.045 82.725 ;
        RECT 60.275 82.680 60.565 82.725 ;
        RECT 61.465 82.680 61.755 82.725 ;
        RECT 57.755 82.540 61.755 82.680 ;
        RECT 57.755 82.495 58.045 82.540 ;
        RECT 60.275 82.495 60.565 82.540 ;
        RECT 61.465 82.495 61.755 82.540 ;
        RECT 63.685 82.680 63.975 82.725 ;
        RECT 64.875 82.680 65.165 82.725 ;
        RECT 67.395 82.680 67.685 82.725 ;
        RECT 63.685 82.540 67.685 82.680 ;
        RECT 63.685 82.495 63.975 82.540 ;
        RECT 64.875 82.495 65.165 82.540 ;
        RECT 67.395 82.495 67.685 82.540 ;
        RECT 94.095 82.680 94.385 82.725 ;
        RECT 96.615 82.680 96.905 82.725 ;
        RECT 97.805 82.680 98.095 82.725 ;
        RECT 94.095 82.540 98.095 82.680 ;
        RECT 94.095 82.495 94.385 82.540 ;
        RECT 96.615 82.495 96.905 82.540 ;
        RECT 97.805 82.495 98.095 82.540 ;
        RECT 98.670 82.480 98.990 82.740 ;
        RECT 103.745 82.495 104.035 82.725 ;
        RECT 107.500 82.680 107.640 83.560 ;
        RECT 126.285 83.515 126.575 83.745 ;
        RECT 127.125 83.700 127.415 83.745 ;
        RECT 129.030 83.700 129.350 83.760 ;
        RECT 127.125 83.560 129.350 83.700 ;
        RECT 127.125 83.515 127.415 83.560 ;
        RECT 108.790 83.160 109.110 83.420 ;
        RECT 109.250 83.160 109.570 83.420 ;
        RECT 108.880 83.020 109.020 83.160 ;
        RECT 110.185 83.020 110.475 83.065 ;
        RECT 108.880 82.880 110.475 83.020 ;
        RECT 110.185 82.835 110.475 82.880 ;
        RECT 119.830 82.820 120.150 83.080 ;
        RECT 125.365 83.020 125.655 83.065 ;
        RECT 126.360 83.020 126.500 83.515 ;
        RECT 129.030 83.500 129.350 83.560 ;
        RECT 135.010 83.500 135.330 83.760 ;
        RECT 145.145 83.700 145.435 83.745 ;
        RECT 146.050 83.700 146.370 83.760 ;
        RECT 145.145 83.560 146.370 83.700 ;
        RECT 145.145 83.515 145.435 83.560 ;
        RECT 146.050 83.500 146.370 83.560 ;
        RECT 127.650 83.360 127.970 83.420 ;
        RECT 128.125 83.360 128.415 83.405 ;
        RECT 129.490 83.360 129.810 83.420 ;
        RECT 127.650 83.220 128.415 83.360 ;
        RECT 127.650 83.160 127.970 83.220 ;
        RECT 128.125 83.175 128.415 83.220 ;
        RECT 129.120 83.220 129.810 83.360 ;
        RECT 125.365 82.880 126.500 83.020 ;
        RECT 125.365 82.835 125.655 82.880 ;
        RECT 128.570 82.820 128.890 83.080 ;
        RECT 108.805 82.680 109.095 82.725 ;
        RECT 107.500 82.540 109.095 82.680 ;
        RECT 108.805 82.495 109.095 82.540 ;
        RECT 40.265 82.340 40.555 82.385 ;
        RECT 41.640 82.340 41.930 82.385 ;
        RECT 40.265 82.200 41.930 82.340 ;
        RECT 40.265 82.155 40.555 82.200 ;
        RECT 41.640 82.155 41.930 82.200 ;
        RECT 43.950 82.340 44.240 82.385 ;
        RECT 45.325 82.340 45.615 82.385 ;
        RECT 43.950 82.200 45.615 82.340 ;
        RECT 43.950 82.155 44.240 82.200 ;
        RECT 45.325 82.155 45.615 82.200 ;
        RECT 50.850 82.340 51.140 82.385 ;
        RECT 52.225 82.340 52.515 82.385 ;
        RECT 50.850 82.200 52.515 82.340 ;
        RECT 50.850 82.155 51.140 82.200 ;
        RECT 52.225 82.155 52.515 82.200 ;
        RECT 54.970 82.340 55.290 82.400 ;
        RECT 55.890 82.340 56.210 82.400 ;
        RECT 54.970 82.200 56.210 82.340 ;
        RECT 54.970 82.140 55.290 82.200 ;
        RECT 55.890 82.140 56.210 82.200 ;
        RECT 58.190 82.340 58.480 82.385 ;
        RECT 59.760 82.340 60.050 82.385 ;
        RECT 61.860 82.340 62.150 82.385 ;
        RECT 58.190 82.200 62.150 82.340 ;
        RECT 58.190 82.155 58.480 82.200 ;
        RECT 59.760 82.155 60.050 82.200 ;
        RECT 61.860 82.155 62.150 82.200 ;
        RECT 63.290 82.340 63.580 82.385 ;
        RECT 65.390 82.340 65.680 82.385 ;
        RECT 66.960 82.340 67.250 82.385 ;
        RECT 63.290 82.200 67.250 82.340 ;
        RECT 63.290 82.155 63.580 82.200 ;
        RECT 65.390 82.155 65.680 82.200 ;
        RECT 66.960 82.155 67.250 82.200 ;
        RECT 94.530 82.340 94.820 82.385 ;
        RECT 96.100 82.340 96.390 82.385 ;
        RECT 98.200 82.340 98.490 82.385 ;
        RECT 94.530 82.200 98.490 82.340 ;
        RECT 103.820 82.340 103.960 82.495 ;
        RECT 118.450 82.480 118.770 82.740 ;
        RECT 118.930 82.680 119.220 82.725 ;
        RECT 121.270 82.680 121.560 82.725 ;
        RECT 129.120 82.680 129.260 83.220 ;
        RECT 129.490 83.160 129.810 83.220 ;
        RECT 143.290 83.360 143.610 83.420 ;
        RECT 143.290 83.220 145.820 83.360 ;
        RECT 143.290 83.160 143.610 83.220 ;
        RECT 134.550 82.820 134.870 83.080 ;
        RECT 135.470 82.820 135.790 83.080 ;
        RECT 145.680 83.065 145.820 83.220 ;
        RECT 145.605 82.835 145.895 83.065 ;
        RECT 118.930 82.540 121.560 82.680 ;
        RECT 118.930 82.495 119.220 82.540 ;
        RECT 121.270 82.495 121.560 82.540 ;
        RECT 123.600 82.540 129.260 82.680 ;
        RECT 145.680 82.680 145.820 82.835 ;
        RECT 146.050 82.820 146.370 83.080 ;
        RECT 146.970 83.020 147.290 83.080 ;
        RECT 147.445 83.020 147.735 83.065 ;
        RECT 146.970 82.880 147.735 83.020 ;
        RECT 146.970 82.820 147.290 82.880 ;
        RECT 147.445 82.835 147.735 82.880 ;
        RECT 148.350 82.820 148.670 83.080 ;
        RECT 147.905 82.680 148.195 82.725 ;
        RECT 145.680 82.540 148.195 82.680 ;
        RECT 109.710 82.340 110.030 82.400 ;
        RECT 123.600 82.385 123.740 82.540 ;
        RECT 147.905 82.495 148.195 82.540 ;
        RECT 111.565 82.340 111.855 82.385 ;
        RECT 103.820 82.200 107.180 82.340 ;
        RECT 94.530 82.155 94.820 82.200 ;
        RECT 96.100 82.155 96.390 82.200 ;
        RECT 98.200 82.155 98.490 82.200 ;
        RECT 25.530 82.000 25.850 82.060 ;
        RECT 26.005 82.000 26.295 82.045 ;
        RECT 25.530 81.860 26.295 82.000 ;
        RECT 25.530 81.800 25.850 81.860 ;
        RECT 26.005 81.815 26.295 81.860 ;
        RECT 31.970 81.800 32.290 82.060 ;
        RECT 35.650 81.800 35.970 82.060 ;
        RECT 55.445 82.000 55.735 82.045 ;
        RECT 57.270 82.000 57.590 82.060 ;
        RECT 55.445 81.860 57.590 82.000 ;
        RECT 55.445 81.815 55.735 81.860 ;
        RECT 57.270 81.800 57.590 81.860 ;
        RECT 82.125 82.000 82.415 82.045 ;
        RECT 82.570 82.000 82.890 82.060 ;
        RECT 82.125 81.860 82.890 82.000 ;
        RECT 82.125 81.815 82.415 81.860 ;
        RECT 82.570 81.800 82.890 81.860 ;
        RECT 101.430 82.000 101.750 82.060 ;
        RECT 101.905 82.000 102.195 82.045 ;
        RECT 101.430 81.860 102.195 82.000 ;
        RECT 101.430 81.800 101.750 81.860 ;
        RECT 101.905 81.815 102.195 81.860 ;
        RECT 102.810 82.000 103.130 82.060 ;
        RECT 107.040 82.045 107.180 82.200 ;
        RECT 109.710 82.200 111.855 82.340 ;
        RECT 109.710 82.140 110.030 82.200 ;
        RECT 111.565 82.155 111.855 82.200 ;
        RECT 119.390 82.340 119.680 82.385 ;
        RECT 120.765 82.340 121.055 82.385 ;
        RECT 119.390 82.200 121.055 82.340 ;
        RECT 119.390 82.155 119.680 82.200 ;
        RECT 120.765 82.155 121.055 82.200 ;
        RECT 123.525 82.155 123.815 82.385 ;
        RECT 141.450 82.140 141.770 82.400 ;
        RECT 106.045 82.000 106.335 82.045 ;
        RECT 102.810 81.860 106.335 82.000 ;
        RECT 102.810 81.800 103.130 81.860 ;
        RECT 106.045 81.815 106.335 81.860 ;
        RECT 106.965 82.000 107.255 82.045 ;
        RECT 111.105 82.000 111.395 82.045 ;
        RECT 106.965 81.860 111.395 82.000 ;
        RECT 106.965 81.815 107.255 81.860 ;
        RECT 111.105 81.815 111.395 81.860 ;
        RECT 114.310 82.000 114.630 82.060 ;
        RECT 114.785 82.000 115.075 82.045 ;
        RECT 114.310 81.860 115.075 82.000 ;
        RECT 114.310 81.800 114.630 81.860 ;
        RECT 114.785 81.815 115.075 81.860 ;
        RECT 116.610 81.800 116.930 82.060 ;
        RECT 124.430 81.800 124.750 82.060 ;
        RECT 127.205 82.000 127.495 82.045 ;
        RECT 130.425 82.000 130.715 82.045 ;
        RECT 127.205 81.860 130.715 82.000 ;
        RECT 127.205 81.815 127.495 81.860 ;
        RECT 130.425 81.815 130.715 81.860 ;
        RECT 132.710 81.800 133.030 82.060 ;
        RECT 142.830 82.000 143.150 82.060 ;
        RECT 143.305 82.000 143.595 82.045 ;
        RECT 142.830 81.860 143.595 82.000 ;
        RECT 142.830 81.800 143.150 81.860 ;
        RECT 143.305 81.815 143.595 81.860 ;
        RECT 143.750 82.000 144.070 82.060 ;
        RECT 144.225 82.000 144.515 82.045 ;
        RECT 143.750 81.860 144.515 82.000 ;
        RECT 143.750 81.800 144.070 81.860 ;
        RECT 144.225 81.815 144.515 81.860 ;
        RECT 146.510 82.000 146.830 82.060 ;
        RECT 146.985 82.000 147.275 82.045 ;
        RECT 146.510 81.860 147.275 82.000 ;
        RECT 146.510 81.800 146.830 81.860 ;
        RECT 146.985 81.815 147.275 81.860 ;
        RECT 22.700 81.180 157.020 81.660 ;
        RECT 35.190 80.780 35.510 81.040 ;
        RECT 41.170 80.980 41.490 81.040 ;
        RECT 47.165 80.980 47.455 81.025 ;
        RECT 41.170 80.840 47.455 80.980 ;
        RECT 41.170 80.780 41.490 80.840 ;
        RECT 47.165 80.795 47.455 80.840 ;
        RECT 51.290 80.780 51.610 81.040 ;
        RECT 52.210 80.980 52.530 81.040 ;
        RECT 57.745 80.980 58.035 81.025 ;
        RECT 58.650 80.980 58.970 81.040 ;
        RECT 52.210 80.840 55.660 80.980 ;
        RECT 52.210 80.780 52.530 80.840 ;
        RECT 28.790 80.640 29.080 80.685 ;
        RECT 30.890 80.640 31.180 80.685 ;
        RECT 32.460 80.640 32.750 80.685 ;
        RECT 28.790 80.500 32.750 80.640 ;
        RECT 28.790 80.455 29.080 80.500 ;
        RECT 30.890 80.455 31.180 80.500 ;
        RECT 32.460 80.455 32.750 80.500 ;
        RECT 41.650 80.640 41.940 80.685 ;
        RECT 43.025 80.640 43.315 80.685 ;
        RECT 41.650 80.500 43.315 80.640 ;
        RECT 41.650 80.455 41.940 80.500 ;
        RECT 43.025 80.455 43.315 80.500 ;
        RECT 43.930 80.640 44.250 80.700 ;
        RECT 45.785 80.640 46.075 80.685 ;
        RECT 54.510 80.640 54.830 80.700 ;
        RECT 43.930 80.500 46.075 80.640 ;
        RECT 43.930 80.440 44.250 80.500 ;
        RECT 45.785 80.455 46.075 80.500 ;
        RECT 46.320 80.500 54.830 80.640 ;
        RECT 28.290 80.100 28.610 80.360 ;
        RECT 29.185 80.300 29.475 80.345 ;
        RECT 30.375 80.300 30.665 80.345 ;
        RECT 32.895 80.300 33.185 80.345 ;
        RECT 29.185 80.160 33.185 80.300 ;
        RECT 29.185 80.115 29.475 80.160 ;
        RECT 30.375 80.115 30.665 80.160 ;
        RECT 32.895 80.115 33.185 80.160 ;
        RECT 41.190 80.300 41.480 80.345 ;
        RECT 43.530 80.300 43.820 80.345 ;
        RECT 41.190 80.160 43.820 80.300 ;
        RECT 41.190 80.115 41.480 80.160 ;
        RECT 43.530 80.115 43.820 80.160 ;
        RECT 46.320 80.020 46.460 80.500 ;
        RECT 50.370 80.300 50.690 80.360 ;
        RECT 53.220 80.345 53.360 80.500 ;
        RECT 54.510 80.440 54.830 80.500 ;
        RECT 55.520 80.640 55.660 80.840 ;
        RECT 57.745 80.840 58.970 80.980 ;
        RECT 57.745 80.795 58.035 80.840 ;
        RECT 58.650 80.780 58.970 80.840 ;
        RECT 60.045 80.980 60.335 81.025 ;
        RECT 60.950 80.980 61.270 81.040 ;
        RECT 60.045 80.840 61.270 80.980 ;
        RECT 60.045 80.795 60.335 80.840 ;
        RECT 60.950 80.780 61.270 80.840 ;
        RECT 64.170 80.980 64.490 81.040 ;
        RECT 65.105 80.980 65.395 81.025 ;
        RECT 64.170 80.840 65.395 80.980 ;
        RECT 64.170 80.780 64.490 80.840 ;
        RECT 65.105 80.795 65.395 80.840 ;
        RECT 77.985 80.980 78.275 81.025 ;
        RECT 78.890 80.980 79.210 81.040 ;
        RECT 77.985 80.840 79.210 80.980 ;
        RECT 77.985 80.795 78.275 80.840 ;
        RECT 78.890 80.780 79.210 80.840 ;
        RECT 92.690 80.780 93.010 81.040 ;
        RECT 95.910 80.980 96.230 81.040 ;
        RECT 96.385 80.980 96.675 81.025 ;
        RECT 95.910 80.840 96.675 80.980 ;
        RECT 95.910 80.780 96.230 80.840 ;
        RECT 96.385 80.795 96.675 80.840 ;
        RECT 97.290 80.980 97.610 81.040 ;
        RECT 97.765 80.980 98.055 81.025 ;
        RECT 97.290 80.840 98.055 80.980 ;
        RECT 97.290 80.780 97.610 80.840 ;
        RECT 97.765 80.795 98.055 80.840 ;
        RECT 98.670 80.980 98.990 81.040 ;
        RECT 110.630 80.980 110.950 81.040 ;
        RECT 128.125 80.980 128.415 81.025 ;
        RECT 128.570 80.980 128.890 81.040 ;
        RECT 98.670 80.840 121.440 80.980 ;
        RECT 98.670 80.780 98.990 80.840 ;
        RECT 59.110 80.640 59.430 80.700 ;
        RECT 61.410 80.640 61.730 80.700 ;
        RECT 55.520 80.500 61.730 80.640 ;
        RECT 52.225 80.300 52.515 80.345 ;
        RECT 50.370 80.160 52.515 80.300 ;
        RECT 50.370 80.100 50.690 80.160 ;
        RECT 52.225 80.115 52.515 80.160 ;
        RECT 53.145 80.115 53.435 80.345 ;
        RECT 53.605 80.300 53.895 80.345 ;
        RECT 54.985 80.300 55.275 80.345 ;
        RECT 53.605 80.160 55.275 80.300 ;
        RECT 53.605 80.115 53.895 80.160 ;
        RECT 54.985 80.115 55.275 80.160 ;
        RECT 27.845 79.775 28.135 80.005 ;
        RECT 29.640 79.960 29.930 80.005 ;
        RECT 31.970 79.960 32.290 80.020 ;
        RECT 29.640 79.820 32.290 79.960 ;
        RECT 29.640 79.775 29.930 79.820 ;
        RECT 27.920 79.620 28.060 79.775 ;
        RECT 31.970 79.760 32.290 79.820 ;
        RECT 35.190 79.960 35.510 80.020 ;
        RECT 36.125 79.960 36.415 80.005 ;
        RECT 35.190 79.820 36.415 79.960 ;
        RECT 35.190 79.760 35.510 79.820 ;
        RECT 36.125 79.775 36.415 79.820 ;
        RECT 40.265 79.960 40.555 80.005 ;
        RECT 40.725 79.960 41.015 80.005 ;
        RECT 40.265 79.820 41.015 79.960 ;
        RECT 40.265 79.775 40.555 79.820 ;
        RECT 40.725 79.775 41.015 79.820 ;
        RECT 42.105 79.960 42.395 80.005 ;
        RECT 44.850 79.960 45.170 80.020 ;
        RECT 42.105 79.820 45.170 79.960 ;
        RECT 42.105 79.775 42.395 79.820 ;
        RECT 44.850 79.760 45.170 79.820 ;
        RECT 46.230 79.760 46.550 80.020 ;
        RECT 47.165 79.775 47.455 80.005 ;
        RECT 49.450 79.970 49.770 80.020 ;
        RECT 49.925 79.970 50.215 80.015 ;
        RECT 49.450 79.830 50.215 79.970 ;
        RECT 36.570 79.620 36.890 79.680 ;
        RECT 27.920 79.480 36.890 79.620 ;
        RECT 36.570 79.420 36.890 79.480 ;
        RECT 37.045 79.620 37.335 79.665 ;
        RECT 41.170 79.620 41.490 79.680 ;
        RECT 37.045 79.480 41.490 79.620 ;
        RECT 37.045 79.435 37.335 79.480 ;
        RECT 41.170 79.420 41.490 79.480 ;
        RECT 26.910 79.080 27.230 79.340 ;
        RECT 37.950 79.080 38.270 79.340 ;
        RECT 47.240 79.280 47.380 79.775 ;
        RECT 49.450 79.760 49.770 79.830 ;
        RECT 49.925 79.785 50.215 79.830 ;
        RECT 50.830 79.760 51.150 80.020 ;
        RECT 55.520 80.005 55.660 80.500 ;
        RECT 59.110 80.440 59.430 80.500 ;
        RECT 61.410 80.440 61.730 80.500 ;
        RECT 73.850 80.640 74.140 80.685 ;
        RECT 75.225 80.640 75.515 80.685 ;
        RECT 73.850 80.500 75.515 80.640 ;
        RECT 73.850 80.455 74.140 80.500 ;
        RECT 75.225 80.455 75.515 80.500 ;
        RECT 79.350 80.640 79.670 80.700 ;
        RECT 81.650 80.640 81.970 80.700 ;
        RECT 79.350 80.500 81.970 80.640 ;
        RECT 79.350 80.440 79.670 80.500 ;
        RECT 81.650 80.440 81.970 80.500 ;
        RECT 82.590 80.640 82.880 80.685 ;
        RECT 83.965 80.640 84.255 80.685 ;
        RECT 82.590 80.500 84.255 80.640 ;
        RECT 82.590 80.455 82.880 80.500 ;
        RECT 83.965 80.455 84.255 80.500 ;
        RECT 88.570 80.640 88.860 80.685 ;
        RECT 89.945 80.640 90.235 80.685 ;
        RECT 88.570 80.500 90.235 80.640 ;
        RECT 88.570 80.455 88.860 80.500 ;
        RECT 89.945 80.455 90.235 80.500 ;
        RECT 55.890 80.300 56.210 80.360 ;
        RECT 73.390 80.300 73.680 80.345 ;
        RECT 75.730 80.300 76.020 80.345 ;
        RECT 55.890 80.160 58.420 80.300 ;
        RECT 55.890 80.100 56.210 80.160 ;
        RECT 52.685 79.775 52.975 80.005 ;
        RECT 54.525 79.775 54.815 80.005 ;
        RECT 55.445 79.775 55.735 80.005 ;
        RECT 52.760 79.620 52.900 79.775 ;
        RECT 54.600 79.620 54.740 79.775 ;
        RECT 57.270 79.760 57.590 80.020 ;
        RECT 58.280 80.005 58.420 80.160 ;
        RECT 73.390 80.160 76.020 80.300 ;
        RECT 73.390 80.115 73.680 80.160 ;
        RECT 75.730 80.115 76.020 80.160 ;
        RECT 82.130 80.300 82.420 80.345 ;
        RECT 84.470 80.300 84.760 80.345 ;
        RECT 82.130 80.160 84.760 80.300 ;
        RECT 82.130 80.115 82.420 80.160 ;
        RECT 84.470 80.115 84.760 80.160 ;
        RECT 88.110 80.300 88.400 80.345 ;
        RECT 90.450 80.300 90.740 80.345 ;
        RECT 97.750 80.300 98.070 80.360 ;
        RECT 101.060 80.345 101.200 80.840 ;
        RECT 110.630 80.780 110.950 80.840 ;
        RECT 101.470 80.640 101.760 80.685 ;
        RECT 103.570 80.640 103.860 80.685 ;
        RECT 105.140 80.640 105.430 80.685 ;
        RECT 101.470 80.500 105.430 80.640 ;
        RECT 101.470 80.455 101.760 80.500 ;
        RECT 103.570 80.455 103.860 80.500 ;
        RECT 105.140 80.455 105.430 80.500 ;
        RECT 107.885 80.640 108.175 80.685 ;
        RECT 109.250 80.640 109.570 80.700 ;
        RECT 107.885 80.500 109.570 80.640 ;
        RECT 107.885 80.455 108.175 80.500 ;
        RECT 109.250 80.440 109.570 80.500 ;
        RECT 115.250 80.640 115.540 80.685 ;
        RECT 116.625 80.640 116.915 80.685 ;
        RECT 115.250 80.500 116.915 80.640 ;
        RECT 115.250 80.455 115.540 80.500 ;
        RECT 116.625 80.455 116.915 80.500 ;
        RECT 118.450 80.640 118.770 80.700 ;
        RECT 119.845 80.640 120.135 80.685 ;
        RECT 118.450 80.500 120.135 80.640 ;
        RECT 118.450 80.440 118.770 80.500 ;
        RECT 119.845 80.455 120.135 80.500 ;
        RECT 88.110 80.160 90.740 80.300 ;
        RECT 88.110 80.115 88.400 80.160 ;
        RECT 90.450 80.115 90.740 80.160 ;
        RECT 96.690 80.160 98.070 80.300 ;
        RECT 58.205 79.775 58.495 80.005 ;
        RECT 59.125 79.960 59.415 80.005 ;
        RECT 59.570 79.960 59.890 80.020 ;
        RECT 59.125 79.820 59.890 79.960 ;
        RECT 59.125 79.775 59.415 79.820 ;
        RECT 59.570 79.760 59.890 79.820 ;
        RECT 66.010 79.760 66.330 80.020 ;
        RECT 72.465 79.960 72.755 80.005 ;
        RECT 72.925 79.960 73.215 80.005 ;
        RECT 72.465 79.820 73.215 79.960 ;
        RECT 72.465 79.775 72.755 79.820 ;
        RECT 72.925 79.775 73.215 79.820 ;
        RECT 73.830 79.960 74.150 80.020 ;
        RECT 74.305 79.960 74.595 80.005 ;
        RECT 73.830 79.820 74.595 79.960 ;
        RECT 73.830 79.760 74.150 79.820 ;
        RECT 74.305 79.775 74.595 79.820 ;
        RECT 79.365 79.960 79.655 80.005 ;
        RECT 79.810 79.960 80.130 80.020 ;
        RECT 79.365 79.820 80.130 79.960 ;
        RECT 79.365 79.775 79.655 79.820 ;
        RECT 79.810 79.760 80.130 79.820 ;
        RECT 81.665 79.960 81.955 80.005 ;
        RECT 82.570 79.960 82.890 80.020 ;
        RECT 81.665 79.820 82.890 79.960 ;
        RECT 81.665 79.775 81.955 79.820 ;
        RECT 82.570 79.760 82.890 79.820 ;
        RECT 83.030 79.760 83.350 80.020 ;
        RECT 83.490 79.760 83.810 80.020 ;
        RECT 87.170 79.960 87.490 80.020 ;
        RECT 87.645 79.960 87.935 80.005 ;
        RECT 87.170 79.820 87.935 79.960 ;
        RECT 87.170 79.760 87.490 79.820 ;
        RECT 87.645 79.775 87.935 79.820 ;
        RECT 88.550 79.960 88.870 80.020 ;
        RECT 89.025 79.960 89.315 80.005 ;
        RECT 88.550 79.820 89.315 79.960 ;
        RECT 88.550 79.760 88.870 79.820 ;
        RECT 89.025 79.775 89.315 79.820 ;
        RECT 54.970 79.620 55.290 79.680 ;
        RECT 57.730 79.620 58.050 79.680 ;
        RECT 52.760 79.480 58.050 79.620 ;
        RECT 54.970 79.420 55.290 79.480 ;
        RECT 57.730 79.420 58.050 79.480 ;
        RECT 76.590 79.620 76.910 79.680 ;
        RECT 80.285 79.620 80.575 79.665 ;
        RECT 83.580 79.620 83.720 79.760 ;
        RECT 76.590 79.480 83.720 79.620 ;
        RECT 93.150 79.620 93.470 79.680 ;
        RECT 96.690 79.665 96.830 80.160 ;
        RECT 97.750 80.100 98.070 80.160 ;
        RECT 100.985 80.115 101.275 80.345 ;
        RECT 101.865 80.300 102.155 80.345 ;
        RECT 103.055 80.300 103.345 80.345 ;
        RECT 105.575 80.300 105.865 80.345 ;
        RECT 111.550 80.300 111.870 80.360 ;
        RECT 101.865 80.160 105.865 80.300 ;
        RECT 101.865 80.115 102.155 80.160 ;
        RECT 103.055 80.115 103.345 80.160 ;
        RECT 105.575 80.115 105.865 80.160 ;
        RECT 109.800 80.160 111.870 80.300 ;
        RECT 98.685 79.960 98.975 80.005 ;
        RECT 97.380 79.820 98.975 79.960 ;
        RECT 95.465 79.620 95.755 79.665 ;
        RECT 93.150 79.480 95.755 79.620 ;
        RECT 76.590 79.420 76.910 79.480 ;
        RECT 80.285 79.435 80.575 79.480 ;
        RECT 93.150 79.420 93.470 79.480 ;
        RECT 95.465 79.435 95.755 79.480 ;
        RECT 96.545 79.435 96.835 79.665 ;
        RECT 50.830 79.280 51.150 79.340 ;
        RECT 47.240 79.140 51.150 79.280 ;
        RECT 50.830 79.080 51.150 79.140 ;
        RECT 81.205 79.280 81.495 79.325 ;
        RECT 83.490 79.280 83.810 79.340 ;
        RECT 81.205 79.140 83.810 79.280 ;
        RECT 81.205 79.095 81.495 79.140 ;
        RECT 83.490 79.080 83.810 79.140 ;
        RECT 86.725 79.280 87.015 79.325 ;
        RECT 95.910 79.280 96.230 79.340 ;
        RECT 97.380 79.325 97.520 79.820 ;
        RECT 98.685 79.775 98.975 79.820 ;
        RECT 101.430 79.960 101.750 80.020 ;
        RECT 109.800 80.005 109.940 80.160 ;
        RECT 111.550 80.100 111.870 80.160 ;
        RECT 114.310 80.100 114.630 80.360 ;
        RECT 121.300 80.345 121.440 80.840 ;
        RECT 128.125 80.840 128.890 80.980 ;
        RECT 128.125 80.795 128.415 80.840 ;
        RECT 128.570 80.780 128.890 80.840 ;
        RECT 129.030 80.980 129.350 81.040 ;
        RECT 141.450 80.980 141.770 81.040 ;
        RECT 129.030 80.840 141.770 80.980 ;
        RECT 129.030 80.780 129.350 80.840 ;
        RECT 121.710 80.640 122.000 80.685 ;
        RECT 123.810 80.640 124.100 80.685 ;
        RECT 125.380 80.640 125.670 80.685 ;
        RECT 121.710 80.500 125.670 80.640 ;
        RECT 121.710 80.455 122.000 80.500 ;
        RECT 123.810 80.455 124.100 80.500 ;
        RECT 125.380 80.455 125.670 80.500 ;
        RECT 133.650 80.640 133.940 80.685 ;
        RECT 135.025 80.640 135.315 80.685 ;
        RECT 133.650 80.500 135.315 80.640 ;
        RECT 133.650 80.455 133.940 80.500 ;
        RECT 135.025 80.455 135.315 80.500 ;
        RECT 137.785 80.640 138.075 80.685 ;
        RECT 138.230 80.640 138.550 80.700 ;
        RECT 137.785 80.500 138.550 80.640 ;
        RECT 137.785 80.455 138.075 80.500 ;
        RECT 138.230 80.440 138.550 80.500 ;
        RECT 114.790 80.300 115.080 80.345 ;
        RECT 117.130 80.300 117.420 80.345 ;
        RECT 114.790 80.160 117.420 80.300 ;
        RECT 114.790 80.115 115.080 80.160 ;
        RECT 117.130 80.115 117.420 80.160 ;
        RECT 121.225 80.115 121.515 80.345 ;
        RECT 122.105 80.300 122.395 80.345 ;
        RECT 123.295 80.300 123.585 80.345 ;
        RECT 125.815 80.300 126.105 80.345 ;
        RECT 122.105 80.160 126.105 80.300 ;
        RECT 122.105 80.115 122.395 80.160 ;
        RECT 123.295 80.115 123.585 80.160 ;
        RECT 125.815 80.115 126.105 80.160 ;
        RECT 132.710 80.100 133.030 80.360 ;
        RECT 141.080 80.345 141.220 80.840 ;
        RECT 141.450 80.780 141.770 80.840 ;
        RECT 145.630 80.640 145.920 80.685 ;
        RECT 147.730 80.640 148.020 80.685 ;
        RECT 149.300 80.640 149.590 80.685 ;
        RECT 145.630 80.500 149.590 80.640 ;
        RECT 145.630 80.455 145.920 80.500 ;
        RECT 147.730 80.455 148.020 80.500 ;
        RECT 149.300 80.455 149.590 80.500 ;
        RECT 133.190 80.300 133.480 80.345 ;
        RECT 135.530 80.300 135.820 80.345 ;
        RECT 133.190 80.160 135.820 80.300 ;
        RECT 133.190 80.115 133.480 80.160 ;
        RECT 135.530 80.115 135.820 80.160 ;
        RECT 141.005 80.115 141.295 80.345 ;
        RECT 143.290 80.100 143.610 80.360 ;
        RECT 145.130 80.100 145.450 80.360 ;
        RECT 146.025 80.300 146.315 80.345 ;
        RECT 147.215 80.300 147.505 80.345 ;
        RECT 149.735 80.300 150.025 80.345 ;
        RECT 146.025 80.160 150.025 80.300 ;
        RECT 146.025 80.115 146.315 80.160 ;
        RECT 147.215 80.115 147.505 80.160 ;
        RECT 149.735 80.115 150.025 80.160 ;
        RECT 102.265 79.960 102.555 80.005 ;
        RECT 101.430 79.820 102.555 79.960 ;
        RECT 101.430 79.760 101.750 79.820 ;
        RECT 102.265 79.775 102.555 79.820 ;
        RECT 109.725 79.775 110.015 80.005 ;
        RECT 110.630 79.760 110.950 80.020 ;
        RECT 115.690 79.760 116.010 80.020 ;
        RECT 122.560 79.960 122.850 80.005 ;
        RECT 124.430 79.960 124.750 80.020 ;
        RECT 122.560 79.820 124.750 79.960 ;
        RECT 122.560 79.775 122.850 79.820 ;
        RECT 124.430 79.760 124.750 79.820 ;
        RECT 128.570 79.760 128.890 80.020 ;
        RECT 129.490 79.760 129.810 80.020 ;
        RECT 130.410 79.960 130.730 80.020 ;
        RECT 130.885 79.960 131.175 80.005 ;
        RECT 130.410 79.820 131.175 79.960 ;
        RECT 130.410 79.760 130.730 79.820 ;
        RECT 130.885 79.775 131.175 79.820 ;
        RECT 134.105 79.960 134.395 80.005 ;
        RECT 135.930 79.960 136.250 80.020 ;
        RECT 134.105 79.820 136.250 79.960 ;
        RECT 134.105 79.775 134.395 79.820 ;
        RECT 135.930 79.760 136.250 79.820 ;
        RECT 142.830 79.760 143.150 80.020 ;
        RECT 146.510 80.005 146.830 80.020 ;
        RECT 146.480 79.960 146.830 80.005 ;
        RECT 146.315 79.820 146.830 79.960 ;
        RECT 146.480 79.775 146.830 79.820 ;
        RECT 146.510 79.760 146.830 79.775 ;
        RECT 86.725 79.140 96.230 79.280 ;
        RECT 86.725 79.095 87.015 79.140 ;
        RECT 95.910 79.080 96.230 79.140 ;
        RECT 97.305 79.095 97.595 79.325 ;
        RECT 110.170 79.080 110.490 79.340 ;
        RECT 119.370 79.080 119.690 79.340 ;
        RECT 141.910 79.280 142.230 79.340 ;
        RECT 144.225 79.280 144.515 79.325 ;
        RECT 141.910 79.140 144.515 79.280 ;
        RECT 141.910 79.080 142.230 79.140 ;
        RECT 144.225 79.095 144.515 79.140 ;
        RECT 148.350 79.280 148.670 79.340 ;
        RECT 152.045 79.280 152.335 79.325 ;
        RECT 148.350 79.140 152.335 79.280 ;
        RECT 148.350 79.080 148.670 79.140 ;
        RECT 152.045 79.095 152.335 79.140 ;
        RECT 22.700 78.460 157.820 78.940 ;
        RECT 30.590 78.060 30.910 78.320 ;
        RECT 34.730 78.060 35.050 78.320 ;
        RECT 36.570 78.260 36.890 78.320 ;
        RECT 36.570 78.120 41.400 78.260 ;
        RECT 36.570 78.060 36.890 78.120 ;
        RECT 37.950 77.920 38.270 77.980 ;
        RECT 34.820 77.780 38.270 77.920 ;
        RECT 41.260 77.920 41.400 78.120 ;
        RECT 44.390 78.060 44.710 78.320 ;
        RECT 44.850 78.060 45.170 78.320 ;
        RECT 49.005 78.075 49.295 78.305 ;
        RECT 49.450 78.260 49.770 78.320 ;
        RECT 58.650 78.260 58.970 78.320 ;
        RECT 61.410 78.260 61.730 78.320 ;
        RECT 49.450 78.120 61.730 78.260 ;
        RECT 49.080 77.920 49.220 78.075 ;
        RECT 49.450 78.060 49.770 78.120 ;
        RECT 41.260 77.780 49.220 77.920 ;
        RECT 25.530 77.380 25.850 77.640 ;
        RECT 26.910 77.380 27.230 77.640 ;
        RECT 34.820 77.625 34.960 77.780 ;
        RECT 37.950 77.720 38.270 77.780 ;
        RECT 49.910 77.720 50.230 77.980 ;
        RECT 52.210 77.920 52.530 77.980 ;
        RECT 53.220 77.965 53.360 78.120 ;
        RECT 58.650 78.060 58.970 78.120 ;
        RECT 61.410 78.060 61.730 78.120 ;
        RECT 61.885 78.260 62.175 78.305 ;
        RECT 62.790 78.260 63.110 78.320 ;
        RECT 61.885 78.120 63.110 78.260 ;
        RECT 61.885 78.075 62.175 78.120 ;
        RECT 62.790 78.060 63.110 78.120 ;
        RECT 73.830 78.060 74.150 78.320 ;
        RECT 80.745 78.260 81.035 78.305 ;
        RECT 83.030 78.260 83.350 78.320 ;
        RECT 80.745 78.120 83.350 78.260 ;
        RECT 80.745 78.075 81.035 78.120 ;
        RECT 83.030 78.060 83.350 78.120 ;
        RECT 86.725 78.260 87.015 78.305 ;
        RECT 88.550 78.260 88.870 78.320 ;
        RECT 86.725 78.120 88.870 78.260 ;
        RECT 86.725 78.075 87.015 78.120 ;
        RECT 88.550 78.060 88.870 78.120 ;
        RECT 94.070 78.260 94.390 78.320 ;
        RECT 95.925 78.260 96.215 78.305 ;
        RECT 94.070 78.120 96.215 78.260 ;
        RECT 94.070 78.060 94.390 78.120 ;
        RECT 95.925 78.075 96.215 78.120 ;
        RECT 113.390 78.260 113.710 78.320 ;
        RECT 113.865 78.260 114.155 78.305 ;
        RECT 113.390 78.120 114.155 78.260 ;
        RECT 113.390 78.060 113.710 78.120 ;
        RECT 113.865 78.075 114.155 78.120 ;
        RECT 115.690 78.060 116.010 78.320 ;
        RECT 121.210 78.060 121.530 78.320 ;
        RECT 129.965 78.075 130.255 78.305 ;
        RECT 134.550 78.260 134.870 78.320 ;
        RECT 135.485 78.260 135.775 78.305 ;
        RECT 134.550 78.120 135.775 78.260 ;
        RECT 51.840 77.780 52.530 77.920 ;
        RECT 34.745 77.395 35.035 77.625 ;
        RECT 35.650 77.380 35.970 77.640 ;
        RECT 43.470 77.380 43.790 77.640 ;
        RECT 45.770 77.380 46.090 77.640 ;
        RECT 51.840 77.625 51.980 77.780 ;
        RECT 52.210 77.720 52.530 77.780 ;
        RECT 53.145 77.735 53.435 77.965 ;
        RECT 79.350 77.920 79.670 77.980 ;
        RECT 56.900 77.780 62.560 77.920 ;
        RECT 56.900 77.625 57.040 77.780 ;
        RECT 51.765 77.395 52.055 77.625 ;
        RECT 54.065 77.580 54.355 77.625 ;
        RECT 55.445 77.580 55.735 77.625 ;
        RECT 54.065 77.440 55.735 77.580 ;
        RECT 54.065 77.395 54.355 77.440 ;
        RECT 55.445 77.395 55.735 77.440 ;
        RECT 56.825 77.395 57.115 77.625 ;
        RECT 57.730 77.580 58.050 77.640 ;
        RECT 62.420 77.625 62.560 77.780 ;
        RECT 76.680 77.780 79.670 77.920 ;
        RECT 58.205 77.580 58.495 77.625 ;
        RECT 57.730 77.440 58.495 77.580 ;
        RECT 57.730 77.380 58.050 77.440 ;
        RECT 58.205 77.395 58.495 77.440 ;
        RECT 62.345 77.395 62.635 77.625 ;
        RECT 72.925 77.395 73.215 77.625 ;
        RECT 75.225 77.580 75.515 77.625 ;
        RECT 75.670 77.580 75.990 77.640 ;
        RECT 75.225 77.440 75.990 77.580 ;
        RECT 75.225 77.395 75.515 77.440 ;
        RECT 26.010 77.240 26.300 77.285 ;
        RECT 28.350 77.240 28.640 77.285 ;
        RECT 26.010 77.100 28.640 77.240 ;
        RECT 26.010 77.055 26.300 77.100 ;
        RECT 28.350 77.055 28.640 77.100 ;
        RECT 57.290 77.240 57.580 77.285 ;
        RECT 59.630 77.240 59.920 77.285 ;
        RECT 57.290 77.100 59.920 77.240 ;
        RECT 57.290 77.055 57.580 77.100 ;
        RECT 59.630 77.055 59.920 77.100 ;
        RECT 26.470 76.900 26.760 76.945 ;
        RECT 27.845 76.900 28.135 76.945 ;
        RECT 26.470 76.760 28.135 76.900 ;
        RECT 26.470 76.715 26.760 76.760 ;
        RECT 27.845 76.715 28.135 76.760 ;
        RECT 54.510 76.900 54.830 76.960 ;
        RECT 55.430 76.900 55.750 76.960 ;
        RECT 54.510 76.760 55.750 76.900 ;
        RECT 54.510 76.700 54.830 76.760 ;
        RECT 55.430 76.700 55.750 76.760 ;
        RECT 57.750 76.900 58.040 76.945 ;
        RECT 59.125 76.900 59.415 76.945 ;
        RECT 57.750 76.760 59.415 76.900 ;
        RECT 73.000 76.900 73.140 77.395 ;
        RECT 75.670 77.380 75.990 77.440 ;
        RECT 76.130 77.380 76.450 77.640 ;
        RECT 76.680 77.625 76.820 77.780 ;
        RECT 79.350 77.720 79.670 77.780 ;
        RECT 79.810 77.920 80.130 77.980 ;
        RECT 81.665 77.920 81.955 77.965 ;
        RECT 79.810 77.780 81.955 77.920 ;
        RECT 79.810 77.720 80.130 77.780 ;
        RECT 81.665 77.735 81.955 77.780 ;
        RECT 83.490 77.720 83.810 77.980 ;
        RECT 116.610 77.720 116.930 77.980 ;
        RECT 130.040 77.920 130.180 78.075 ;
        RECT 134.550 78.060 134.870 78.120 ;
        RECT 135.485 78.075 135.775 78.120 ;
        RECT 135.930 78.060 136.250 78.320 ;
        RECT 141.910 78.060 142.230 78.320 ;
        RECT 142.830 78.260 143.150 78.320 ;
        RECT 145.605 78.260 145.895 78.305 ;
        RECT 142.830 78.120 145.895 78.260 ;
        RECT 142.830 78.060 143.150 78.120 ;
        RECT 145.605 78.075 145.895 78.120 ;
        RECT 146.525 77.920 146.815 77.965 ;
        RECT 146.970 77.920 147.290 77.980 ;
        RECT 130.040 77.780 130.410 77.920 ;
        RECT 76.605 77.395 76.895 77.625 ;
        RECT 77.510 77.580 77.830 77.640 ;
        RECT 82.585 77.580 82.875 77.625 ;
        RECT 77.510 77.440 82.875 77.580 ;
        RECT 77.510 77.380 77.830 77.440 ;
        RECT 82.585 77.395 82.875 77.440 ;
        RECT 85.790 77.380 86.110 77.640 ;
        RECT 87.170 77.380 87.490 77.640 ;
        RECT 92.230 77.380 92.550 77.640 ;
        RECT 108.805 77.580 109.095 77.625 ;
        RECT 109.710 77.580 110.030 77.640 ;
        RECT 108.805 77.440 110.030 77.580 ;
        RECT 108.805 77.395 109.095 77.440 ;
        RECT 109.710 77.380 110.030 77.440 ;
        RECT 110.170 77.380 110.490 77.640 ;
        RECT 114.770 77.380 115.090 77.640 ;
        RECT 116.165 77.580 116.455 77.625 ;
        RECT 116.700 77.580 116.840 77.720 ;
        RECT 116.165 77.440 116.840 77.580 ;
        RECT 117.545 77.580 117.835 77.625 ;
        RECT 123.510 77.580 123.830 77.640 ;
        RECT 117.545 77.440 123.830 77.580 ;
        RECT 116.165 77.395 116.455 77.440 ;
        RECT 117.545 77.395 117.835 77.440 ;
        RECT 123.510 77.380 123.830 77.440 ;
        RECT 129.030 77.380 129.350 77.640 ;
        RECT 130.270 77.580 130.410 77.780 ;
        RECT 146.525 77.780 147.290 77.920 ;
        RECT 146.525 77.735 146.815 77.780 ;
        RECT 146.970 77.720 147.290 77.780 ;
        RECT 147.445 77.920 147.735 77.965 ;
        RECT 148.350 77.920 148.670 77.980 ;
        RECT 147.445 77.780 148.670 77.920 ;
        RECT 147.445 77.735 147.735 77.780 ;
        RECT 148.350 77.720 148.670 77.780 ;
        RECT 131.805 77.580 132.095 77.625 ;
        RECT 130.270 77.440 132.095 77.580 ;
        RECT 131.805 77.395 132.095 77.440 ;
        RECT 136.850 77.380 137.170 77.640 ;
        RECT 140.085 77.580 140.375 77.625 ;
        RECT 143.750 77.580 144.070 77.640 ;
        RECT 140.085 77.440 144.070 77.580 ;
        RECT 140.085 77.395 140.375 77.440 ;
        RECT 143.750 77.380 144.070 77.440 ;
        RECT 77.065 77.240 77.355 77.285 ;
        RECT 78.445 77.240 78.735 77.285 ;
        RECT 77.065 77.100 78.735 77.240 ;
        RECT 77.065 77.055 77.355 77.100 ;
        RECT 78.445 77.055 78.735 77.100 ;
        RECT 78.890 77.040 79.210 77.300 ;
        RECT 79.350 77.040 79.670 77.300 ;
        RECT 79.825 77.055 80.115 77.285 ;
        RECT 90.405 77.240 90.695 77.285 ;
        RECT 90.865 77.240 91.155 77.285 ;
        RECT 90.405 77.100 91.155 77.240 ;
        RECT 90.405 77.055 90.695 77.100 ;
        RECT 90.865 77.055 91.155 77.100 ;
        RECT 91.330 77.240 91.620 77.285 ;
        RECT 93.670 77.240 93.960 77.285 ;
        RECT 91.330 77.100 93.960 77.240 ;
        RECT 91.330 77.055 91.620 77.100 ;
        RECT 93.670 77.055 93.960 77.100 ;
        RECT 109.270 77.240 109.560 77.285 ;
        RECT 111.610 77.240 111.900 77.285 ;
        RECT 109.270 77.100 111.900 77.240 ;
        RECT 109.270 77.055 109.560 77.100 ;
        RECT 111.610 77.055 111.900 77.100 ;
        RECT 116.630 77.240 116.920 77.285 ;
        RECT 118.970 77.240 119.260 77.285 ;
        RECT 116.630 77.100 119.260 77.240 ;
        RECT 116.630 77.055 116.920 77.100 ;
        RECT 118.970 77.055 119.260 77.100 ;
        RECT 75.210 76.900 75.530 76.960 ;
        RECT 73.000 76.760 75.530 76.900 ;
        RECT 57.750 76.715 58.040 76.760 ;
        RECT 59.125 76.715 59.415 76.760 ;
        RECT 75.210 76.700 75.530 76.760 ;
        RECT 75.685 76.900 75.975 76.945 ;
        RECT 76.130 76.900 76.450 76.960 ;
        RECT 79.900 76.900 80.040 77.055 ;
        RECT 130.410 77.040 130.730 77.300 ;
        RECT 130.890 77.240 131.180 77.285 ;
        RECT 133.230 77.240 133.520 77.285 ;
        RECT 130.890 77.100 133.520 77.240 ;
        RECT 130.890 77.055 131.180 77.100 ;
        RECT 133.230 77.055 133.520 77.100 ;
        RECT 75.685 76.760 80.040 76.900 ;
        RECT 81.650 76.900 81.970 76.960 ;
        RECT 84.425 76.900 84.715 76.945 ;
        RECT 81.650 76.760 84.715 76.900 ;
        RECT 75.685 76.715 75.975 76.760 ;
        RECT 76.130 76.700 76.450 76.760 ;
        RECT 81.650 76.700 81.970 76.760 ;
        RECT 84.425 76.715 84.715 76.760 ;
        RECT 91.790 76.900 92.080 76.945 ;
        RECT 93.165 76.900 93.455 76.945 ;
        RECT 91.790 76.760 93.455 76.900 ;
        RECT 91.790 76.715 92.080 76.760 ;
        RECT 93.165 76.715 93.455 76.760 ;
        RECT 109.730 76.900 110.020 76.945 ;
        RECT 111.105 76.900 111.395 76.945 ;
        RECT 109.730 76.760 111.395 76.900 ;
        RECT 109.730 76.715 110.020 76.760 ;
        RECT 111.105 76.715 111.395 76.760 ;
        RECT 117.090 76.900 117.380 76.945 ;
        RECT 118.465 76.900 118.755 76.945 ;
        RECT 117.090 76.760 118.755 76.900 ;
        RECT 117.090 76.715 117.380 76.760 ;
        RECT 118.465 76.715 118.755 76.760 ;
        RECT 131.350 76.900 131.640 76.945 ;
        RECT 132.725 76.900 133.015 76.945 ;
        RECT 131.350 76.760 133.015 76.900 ;
        RECT 131.350 76.715 131.640 76.760 ;
        RECT 132.725 76.715 133.015 76.760 ;
        RECT 142.845 76.900 143.135 76.945 ;
        RECT 146.050 76.900 146.370 76.960 ;
        RECT 142.845 76.760 146.370 76.900 ;
        RECT 142.845 76.715 143.135 76.760 ;
        RECT 146.050 76.700 146.370 76.760 ;
        RECT 33.365 76.560 33.655 76.605 ;
        RECT 34.730 76.560 35.050 76.620 ;
        RECT 33.365 76.420 35.050 76.560 ;
        RECT 33.365 76.375 33.655 76.420 ;
        RECT 34.730 76.360 35.050 76.420 ;
        RECT 49.925 76.560 50.215 76.605 ;
        RECT 50.370 76.560 50.690 76.620 ;
        RECT 49.925 76.420 50.690 76.560 ;
        RECT 49.925 76.375 50.215 76.420 ;
        RECT 50.370 76.360 50.690 76.420 ;
        RECT 66.930 76.360 67.250 76.620 ;
        RECT 68.310 76.360 68.630 76.620 ;
        RECT 101.430 76.560 101.750 76.620 ;
        RECT 101.905 76.560 102.195 76.605 ;
        RECT 101.430 76.420 102.195 76.560 ;
        RECT 101.430 76.360 101.750 76.420 ;
        RECT 101.905 76.375 102.195 76.420 ;
        RECT 141.925 76.560 142.215 76.605 ;
        RECT 142.370 76.560 142.690 76.620 ;
        RECT 141.925 76.420 142.690 76.560 ;
        RECT 141.925 76.375 142.215 76.420 ;
        RECT 142.370 76.360 142.690 76.420 ;
        RECT 22.700 75.740 157.020 76.220 ;
        RECT 41.170 75.340 41.490 75.600 ;
        RECT 57.730 75.340 58.050 75.600 ;
        RECT 75.210 75.340 75.530 75.600 ;
        RECT 76.130 75.340 76.450 75.600 ;
        RECT 85.790 75.540 86.110 75.600 ;
        RECT 88.105 75.540 88.395 75.585 ;
        RECT 85.790 75.400 88.395 75.540 ;
        RECT 85.790 75.340 86.110 75.400 ;
        RECT 88.105 75.355 88.395 75.400 ;
        RECT 89.945 75.355 90.235 75.585 ;
        RECT 91.325 75.540 91.615 75.585 ;
        RECT 92.230 75.540 92.550 75.600 ;
        RECT 91.325 75.400 92.550 75.540 ;
        RECT 91.325 75.355 91.615 75.400 ;
        RECT 28.770 75.200 29.060 75.245 ;
        RECT 30.145 75.200 30.435 75.245 ;
        RECT 28.770 75.060 30.435 75.200 ;
        RECT 28.770 75.015 29.060 75.060 ;
        RECT 30.145 75.015 30.435 75.060 ;
        RECT 37.050 75.200 37.340 75.245 ;
        RECT 38.425 75.200 38.715 75.245 ;
        RECT 44.390 75.200 44.710 75.260 ;
        RECT 46.230 75.200 46.550 75.260 ;
        RECT 37.050 75.060 38.715 75.200 ;
        RECT 37.050 75.015 37.340 75.060 ;
        RECT 38.425 75.015 38.715 75.060 ;
        RECT 42.180 75.060 46.550 75.200 ;
        RECT 28.310 74.860 28.600 74.905 ;
        RECT 30.650 74.860 30.940 74.905 ;
        RECT 28.310 74.720 30.940 74.860 ;
        RECT 28.310 74.675 28.600 74.720 ;
        RECT 30.650 74.675 30.940 74.720 ;
        RECT 34.730 74.860 35.050 74.920 ;
        RECT 36.125 74.860 36.415 74.905 ;
        RECT 34.730 74.720 36.415 74.860 ;
        RECT 34.730 74.660 35.050 74.720 ;
        RECT 36.125 74.675 36.415 74.720 ;
        RECT 36.590 74.860 36.880 74.905 ;
        RECT 38.930 74.860 39.220 74.905 ;
        RECT 36.590 74.720 39.220 74.860 ;
        RECT 36.590 74.675 36.880 74.720 ;
        RECT 38.930 74.675 39.220 74.720 ;
        RECT 27.385 74.520 27.675 74.565 ;
        RECT 27.845 74.520 28.135 74.565 ;
        RECT 27.385 74.380 28.135 74.520 ;
        RECT 27.385 74.335 27.675 74.380 ;
        RECT 27.845 74.335 28.135 74.380 ;
        RECT 29.225 74.335 29.515 74.565 ;
        RECT 29.300 74.180 29.440 74.335 ;
        RECT 34.270 74.320 34.590 74.580 ;
        RECT 37.030 74.520 37.350 74.580 ;
        RECT 37.505 74.520 37.795 74.565 ;
        RECT 37.030 74.380 37.795 74.520 ;
        RECT 37.030 74.320 37.350 74.380 ;
        RECT 37.505 74.335 37.795 74.380 ;
        RECT 41.645 74.520 41.935 74.565 ;
        RECT 42.180 74.520 42.320 75.060 ;
        RECT 44.390 75.000 44.710 75.060 ;
        RECT 46.230 75.000 46.550 75.060 ;
        RECT 67.870 75.200 68.160 75.245 ;
        RECT 69.245 75.200 69.535 75.245 ;
        RECT 67.870 75.060 69.535 75.200 ;
        RECT 67.870 75.015 68.160 75.060 ;
        RECT 69.245 75.015 69.535 75.060 ;
        RECT 77.510 75.200 77.830 75.260 ;
        RECT 77.985 75.200 78.275 75.245 ;
        RECT 80.270 75.200 80.590 75.260 ;
        RECT 77.510 75.060 80.590 75.200 ;
        RECT 90.020 75.200 90.160 75.355 ;
        RECT 92.230 75.340 92.550 75.400 ;
        RECT 99.145 75.355 99.435 75.585 ;
        RECT 111.565 75.355 111.855 75.585 ;
        RECT 112.485 75.540 112.775 75.585 ;
        RECT 114.770 75.540 115.090 75.600 ;
        RECT 112.485 75.400 115.090 75.540 ;
        RECT 112.485 75.355 112.775 75.400 ;
        RECT 95.925 75.200 96.215 75.245 ;
        RECT 99.220 75.200 99.360 75.355 ;
        RECT 90.020 75.060 99.360 75.200 ;
        RECT 102.370 75.200 102.660 75.245 ;
        RECT 103.745 75.200 104.035 75.245 ;
        RECT 102.370 75.060 104.035 75.200 ;
        RECT 111.640 75.200 111.780 75.355 ;
        RECT 114.770 75.340 115.090 75.400 ;
        RECT 131.790 75.340 132.110 75.600 ;
        RECT 132.725 75.540 133.015 75.585 ;
        RECT 136.850 75.540 137.170 75.600 ;
        RECT 132.725 75.400 137.170 75.540 ;
        RECT 132.725 75.355 133.015 75.400 ;
        RECT 136.850 75.340 137.170 75.400 ;
        RECT 146.525 75.540 146.815 75.585 ;
        RECT 146.970 75.540 147.290 75.600 ;
        RECT 146.525 75.400 147.290 75.540 ;
        RECT 146.525 75.355 146.815 75.400 ;
        RECT 146.970 75.340 147.290 75.400 ;
        RECT 113.865 75.200 114.155 75.245 ;
        RECT 116.150 75.200 116.470 75.260 ;
        RECT 142.390 75.200 142.680 75.245 ;
        RECT 143.765 75.200 144.055 75.245 ;
        RECT 111.640 75.060 115.920 75.200 ;
        RECT 77.510 75.000 77.830 75.060 ;
        RECT 77.985 75.015 78.275 75.060 ;
        RECT 80.270 75.000 80.590 75.060 ;
        RECT 95.925 75.015 96.215 75.060 ;
        RECT 102.370 75.015 102.660 75.060 ;
        RECT 103.745 75.015 104.035 75.060 ;
        RECT 113.865 75.015 114.155 75.060 ;
        RECT 64.645 74.860 64.935 74.905 ;
        RECT 42.640 74.720 64.935 74.860 ;
        RECT 42.640 74.565 42.780 74.720 ;
        RECT 41.645 74.380 42.320 74.520 ;
        RECT 41.645 74.335 41.935 74.380 ;
        RECT 42.565 74.335 42.855 74.565 ;
        RECT 50.385 74.520 50.675 74.565 ;
        RECT 50.830 74.520 51.150 74.580 ;
        RECT 50.385 74.380 51.150 74.520 ;
        RECT 50.385 74.335 50.675 74.380 ;
        RECT 40.710 74.180 41.030 74.240 ;
        RECT 42.105 74.180 42.395 74.225 ;
        RECT 29.300 74.040 42.395 74.180 ;
        RECT 50.460 74.180 50.600 74.335 ;
        RECT 50.830 74.320 51.150 74.380 ;
        RECT 51.305 74.520 51.595 74.565 ;
        RECT 54.970 74.520 55.290 74.580 ;
        RECT 56.365 74.520 56.655 74.565 ;
        RECT 51.305 74.380 56.655 74.520 ;
        RECT 51.305 74.335 51.595 74.380 ;
        RECT 54.970 74.320 55.290 74.380 ;
        RECT 56.365 74.335 56.655 74.380 ;
        RECT 58.190 74.520 58.510 74.580 ;
        RECT 58.740 74.565 58.880 74.720 ;
        RECT 64.645 74.675 64.935 74.720 ;
        RECT 66.930 74.660 67.250 74.920 ;
        RECT 67.410 74.860 67.700 74.905 ;
        RECT 69.750 74.860 70.040 74.905 ;
        RECT 75.670 74.860 75.990 74.920 ;
        RECT 96.385 74.860 96.675 74.905 ;
        RECT 67.410 74.720 70.040 74.860 ;
        RECT 67.410 74.675 67.700 74.720 ;
        RECT 69.750 74.675 70.040 74.720 ;
        RECT 72.540 74.720 75.990 74.860 ;
        RECT 58.665 74.520 58.955 74.565 ;
        RECT 58.190 74.380 58.955 74.520 ;
        RECT 58.190 74.320 58.510 74.380 ;
        RECT 58.665 74.335 58.955 74.380 ;
        RECT 59.110 74.320 59.430 74.580 ;
        RECT 60.030 74.320 60.350 74.580 ;
        RECT 60.490 74.320 60.810 74.580 ;
        RECT 63.710 74.520 64.030 74.580 ;
        RECT 64.185 74.520 64.475 74.565 ;
        RECT 61.040 74.380 64.475 74.520 ;
        RECT 54.510 74.180 54.830 74.240 ;
        RECT 55.445 74.180 55.735 74.225 ;
        RECT 50.460 74.040 51.520 74.180 ;
        RECT 40.710 73.980 41.030 74.040 ;
        RECT 42.105 73.995 42.395 74.040 ;
        RECT 31.510 73.840 31.830 73.900 ;
        RECT 32.905 73.840 33.195 73.885 ;
        RECT 31.510 73.700 33.195 73.840 ;
        RECT 31.510 73.640 31.830 73.700 ;
        RECT 32.905 73.655 33.195 73.700 ;
        RECT 35.205 73.840 35.495 73.885 ;
        RECT 36.110 73.840 36.430 73.900 ;
        RECT 35.205 73.700 36.430 73.840 ;
        RECT 35.205 73.655 35.495 73.700 ;
        RECT 36.110 73.640 36.430 73.700 ;
        RECT 49.910 73.840 50.230 73.900 ;
        RECT 50.845 73.840 51.135 73.885 ;
        RECT 49.910 73.700 51.135 73.840 ;
        RECT 51.380 73.840 51.520 74.040 ;
        RECT 54.510 74.040 55.735 74.180 ;
        RECT 54.510 73.980 54.830 74.040 ;
        RECT 55.445 73.995 55.735 74.040 ;
        RECT 57.285 74.180 57.575 74.225 ;
        RECT 61.040 74.180 61.180 74.380 ;
        RECT 63.710 74.320 64.030 74.380 ;
        RECT 64.185 74.335 64.475 74.380 ;
        RECT 65.090 74.320 65.410 74.580 ;
        RECT 72.540 74.565 72.680 74.720 ;
        RECT 75.670 74.660 75.990 74.720 ;
        RECT 83.120 74.720 86.020 74.860 ;
        RECT 68.325 74.335 68.615 74.565 ;
        RECT 72.465 74.335 72.755 74.565 ;
        RECT 73.385 74.520 73.675 74.565 ;
        RECT 76.130 74.520 76.450 74.580 ;
        RECT 78.890 74.520 79.210 74.580 ;
        RECT 81.650 74.520 81.970 74.580 ;
        RECT 83.120 74.565 83.260 74.720 ;
        RECT 83.045 74.520 83.335 74.565 ;
        RECT 73.385 74.380 83.335 74.520 ;
        RECT 73.385 74.335 73.675 74.380 ;
        RECT 57.285 74.040 61.180 74.180 ;
        RECT 62.790 74.180 63.110 74.240 ;
        RECT 65.180 74.180 65.320 74.320 ;
        RECT 62.790 74.040 65.320 74.180 ;
        RECT 68.400 74.180 68.540 74.335 ;
        RECT 76.130 74.320 76.450 74.380 ;
        RECT 78.890 74.320 79.210 74.380 ;
        RECT 81.650 74.320 81.970 74.380 ;
        RECT 83.045 74.335 83.335 74.380 ;
        RECT 83.950 74.320 84.270 74.580 ;
        RECT 85.880 74.565 86.020 74.720 ;
        RECT 95.080 74.720 96.675 74.860 ;
        RECT 85.805 74.335 86.095 74.565 ;
        RECT 86.265 74.520 86.555 74.565 ;
        RECT 89.025 74.520 89.315 74.565 ;
        RECT 86.265 74.380 89.315 74.520 ;
        RECT 86.265 74.335 86.555 74.380 ;
        RECT 89.025 74.335 89.315 74.380 ;
        RECT 89.945 74.335 90.235 74.565 ;
        RECT 90.405 74.520 90.695 74.565 ;
        RECT 90.850 74.520 91.170 74.580 ;
        RECT 90.405 74.380 91.170 74.520 ;
        RECT 90.405 74.335 90.695 74.380 ;
        RECT 72.925 74.180 73.215 74.225 ;
        RECT 68.400 74.040 73.215 74.180 ;
        RECT 57.285 73.995 57.575 74.040 ;
        RECT 57.360 73.840 57.500 73.995 ;
        RECT 62.790 73.980 63.110 74.040 ;
        RECT 72.925 73.995 73.215 74.040 ;
        RECT 88.550 74.180 88.870 74.240 ;
        RECT 90.020 74.180 90.160 74.335 ;
        RECT 90.850 74.320 91.170 74.380 ;
        RECT 93.610 74.520 93.930 74.580 ;
        RECT 95.080 74.565 95.220 74.720 ;
        RECT 96.385 74.675 96.675 74.720 ;
        RECT 101.430 74.660 101.750 74.920 ;
        RECT 101.910 74.860 102.200 74.905 ;
        RECT 104.250 74.860 104.540 74.905 ;
        RECT 101.910 74.720 104.540 74.860 ;
        RECT 101.910 74.675 102.200 74.720 ;
        RECT 104.250 74.675 104.540 74.720 ;
        RECT 111.550 74.860 111.870 74.920 ;
        RECT 115.780 74.905 115.920 75.060 ;
        RECT 116.150 75.060 127.835 75.200 ;
        RECT 116.150 75.000 116.610 75.060 ;
        RECT 116.470 74.905 116.610 75.000 ;
        RECT 111.550 74.720 114.540 74.860 ;
        RECT 111.550 74.660 111.870 74.720 ;
        RECT 95.005 74.520 95.295 74.565 ;
        RECT 95.925 74.520 96.215 74.565 ;
        RECT 97.290 74.520 97.610 74.580 ;
        RECT 93.610 74.380 95.295 74.520 ;
        RECT 93.610 74.320 93.930 74.380 ;
        RECT 95.005 74.335 95.295 74.380 ;
        RECT 95.540 74.380 97.610 74.520 ;
        RECT 88.550 74.040 90.160 74.180 ;
        RECT 88.550 73.980 88.870 74.040 ;
        RECT 51.380 73.700 57.500 73.840 ;
        RECT 57.730 73.840 58.050 73.900 ;
        RECT 61.885 73.840 62.175 73.885 ;
        RECT 57.730 73.700 62.175 73.840 ;
        RECT 49.910 73.640 50.230 73.700 ;
        RECT 50.845 73.655 51.135 73.700 ;
        RECT 57.730 73.640 58.050 73.700 ;
        RECT 61.885 73.655 62.175 73.700 ;
        RECT 72.005 73.840 72.295 73.885 ;
        RECT 74.290 73.840 74.610 73.900 ;
        RECT 72.005 73.700 74.610 73.840 ;
        RECT 72.005 73.655 72.295 73.700 ;
        RECT 74.290 73.640 74.610 73.700 ;
        RECT 75.670 73.840 75.990 73.900 ;
        RECT 76.145 73.840 76.435 73.885 ;
        RECT 75.670 73.700 76.435 73.840 ;
        RECT 75.670 73.640 75.990 73.700 ;
        RECT 76.145 73.655 76.435 73.700 ;
        RECT 83.490 73.640 83.810 73.900 ;
        RECT 83.950 73.840 84.270 73.900 ;
        RECT 95.540 73.840 95.680 74.380 ;
        RECT 95.925 74.335 96.215 74.380 ;
        RECT 97.290 74.320 97.610 74.380 ;
        RECT 98.225 74.520 98.515 74.565 ;
        RECT 99.145 74.520 99.435 74.565 ;
        RECT 98.225 74.380 99.435 74.520 ;
        RECT 98.225 74.335 98.515 74.380 ;
        RECT 99.145 74.335 99.435 74.380 ;
        RECT 99.590 74.320 99.910 74.580 ;
        RECT 102.350 74.520 102.670 74.580 ;
        RECT 102.825 74.520 103.115 74.565 ;
        RECT 102.350 74.380 103.115 74.520 ;
        RECT 102.350 74.320 102.670 74.380 ;
        RECT 102.825 74.335 103.115 74.380 ;
        RECT 103.730 74.520 104.050 74.580 ;
        RECT 107.885 74.520 108.175 74.565 ;
        RECT 103.730 74.380 108.175 74.520 ;
        RECT 103.730 74.320 104.050 74.380 ;
        RECT 107.885 74.335 108.175 74.380 ;
        RECT 109.725 74.520 110.015 74.565 ;
        RECT 111.090 74.520 111.410 74.580 ;
        RECT 113.390 74.520 113.710 74.580 ;
        RECT 109.725 74.380 111.410 74.520 ;
        RECT 112.100 74.500 113.710 74.520 ;
        RECT 109.725 74.335 110.015 74.380 ;
        RECT 106.950 74.180 107.270 74.240 ;
        RECT 100.600 74.040 107.270 74.180 ;
        RECT 107.960 74.180 108.100 74.335 ;
        RECT 111.090 74.320 111.410 74.380 ;
        RECT 111.640 74.380 113.710 74.500 ;
        RECT 111.640 74.360 112.240 74.380 ;
        RECT 111.640 74.180 111.780 74.360 ;
        RECT 113.390 74.320 113.710 74.380 ;
        RECT 113.850 74.520 114.170 74.580 ;
        RECT 114.400 74.565 114.540 74.720 ;
        RECT 115.705 74.675 115.995 74.905 ;
        RECT 116.470 74.720 116.870 74.905 ;
        RECT 116.580 74.675 116.870 74.720 ;
        RECT 117.050 74.860 117.340 74.905 ;
        RECT 118.465 74.860 118.755 74.905 ;
        RECT 117.050 74.720 118.755 74.860 ;
        RECT 117.050 74.675 117.340 74.720 ;
        RECT 118.465 74.675 118.755 74.720 ;
        RECT 114.325 74.520 114.615 74.565 ;
        RECT 113.850 74.380 114.615 74.520 ;
        RECT 113.850 74.320 114.170 74.380 ;
        RECT 114.325 74.335 114.615 74.380 ;
        RECT 114.770 74.520 115.090 74.580 ;
        RECT 123.140 74.565 123.280 75.060 ;
        RECT 123.510 74.860 123.830 74.920 ;
        RECT 126.730 74.860 127.050 74.920 ;
        RECT 123.510 74.720 127.050 74.860 ;
        RECT 123.510 74.660 123.830 74.720 ;
        RECT 126.730 74.660 127.050 74.720 ;
        RECT 127.695 74.565 127.835 75.060 ;
        RECT 142.390 75.060 144.055 75.200 ;
        RECT 142.390 75.015 142.680 75.060 ;
        RECT 143.765 75.015 144.055 75.060 ;
        RECT 128.125 74.860 128.415 74.905 ;
        RECT 131.345 74.860 131.635 74.905 ;
        RECT 128.125 74.720 131.635 74.860 ;
        RECT 128.125 74.675 128.415 74.720 ;
        RECT 131.345 74.675 131.635 74.720 ;
        RECT 141.930 74.860 142.220 74.905 ;
        RECT 144.270 74.860 144.560 74.905 ;
        RECT 141.930 74.720 144.560 74.860 ;
        RECT 141.930 74.675 142.220 74.720 ;
        RECT 144.270 74.675 144.560 74.720 ;
        RECT 116.165 74.520 116.455 74.565 ;
        RECT 118.005 74.520 118.295 74.565 ;
        RECT 114.770 74.380 118.295 74.520 ;
        RECT 114.770 74.320 115.090 74.380 ;
        RECT 116.165 74.335 116.455 74.380 ;
        RECT 118.005 74.335 118.295 74.380 ;
        RECT 118.925 74.335 119.215 74.565 ;
        RECT 123.065 74.335 123.355 74.565 ;
        RECT 123.985 74.335 124.275 74.565 ;
        RECT 127.665 74.335 127.955 74.565 ;
        RECT 107.960 74.040 111.780 74.180 ;
        RECT 112.470 74.180 112.790 74.240 ;
        RECT 119.000 74.180 119.140 74.335 ;
        RECT 120.750 74.180 121.070 74.240 ;
        RECT 112.470 74.040 121.070 74.180 ;
        RECT 83.950 73.700 95.680 73.840 ;
        RECT 95.910 73.840 96.230 73.900 ;
        RECT 100.600 73.840 100.740 74.040 ;
        RECT 106.950 73.980 107.270 74.040 ;
        RECT 112.470 73.980 112.790 74.040 ;
        RECT 120.750 73.980 121.070 74.040 ;
        RECT 122.130 74.180 122.450 74.240 ;
        RECT 124.060 74.180 124.200 74.335 ;
        RECT 130.870 74.320 131.190 74.580 ;
        RECT 134.550 74.520 134.870 74.580 ;
        RECT 135.025 74.520 135.315 74.565 ;
        RECT 135.930 74.520 136.250 74.580 ;
        RECT 134.550 74.380 135.315 74.520 ;
        RECT 134.550 74.320 134.870 74.380 ;
        RECT 135.025 74.335 135.315 74.380 ;
        RECT 135.560 74.380 136.250 74.520 ;
        RECT 135.560 74.180 135.700 74.380 ;
        RECT 135.930 74.320 136.250 74.380 ;
        RECT 137.325 74.520 137.615 74.565 ;
        RECT 138.690 74.520 139.010 74.580 ;
        RECT 137.325 74.380 139.010 74.520 ;
        RECT 137.325 74.335 137.615 74.380 ;
        RECT 138.690 74.320 139.010 74.380 ;
        RECT 141.005 74.520 141.295 74.565 ;
        RECT 141.465 74.520 141.755 74.565 ;
        RECT 141.005 74.380 141.755 74.520 ;
        RECT 141.005 74.335 141.295 74.380 ;
        RECT 141.465 74.335 141.755 74.380 ;
        RECT 142.845 74.335 143.135 74.565 ;
        RECT 142.920 74.180 143.060 74.335 ;
        RECT 122.130 74.040 124.200 74.180 ;
        RECT 122.130 73.980 122.450 74.040 ;
        RECT 95.910 73.700 100.740 73.840 ;
        RECT 100.985 73.840 101.275 73.885 ;
        RECT 101.430 73.840 101.750 73.900 ;
        RECT 100.985 73.700 101.750 73.840 ;
        RECT 83.950 73.640 84.270 73.700 ;
        RECT 95.910 73.640 96.230 73.700 ;
        RECT 100.985 73.655 101.275 73.700 ;
        RECT 101.430 73.640 101.750 73.700 ;
        RECT 105.110 73.840 105.430 73.900 ;
        RECT 106.505 73.840 106.795 73.885 ;
        RECT 105.110 73.700 106.795 73.840 ;
        RECT 105.110 73.640 105.430 73.700 ;
        RECT 106.505 73.655 106.795 73.700 ;
        RECT 108.805 73.840 109.095 73.885 ;
        RECT 109.250 73.840 109.570 73.900 ;
        RECT 108.805 73.700 109.570 73.840 ;
        RECT 108.805 73.655 109.095 73.700 ;
        RECT 109.250 73.640 109.570 73.700 ;
        RECT 111.550 73.640 111.870 73.900 ;
        RECT 114.785 73.840 115.075 73.885 ;
        RECT 119.830 73.840 120.150 73.900 ;
        RECT 114.785 73.700 120.150 73.840 ;
        RECT 124.060 73.840 124.200 74.040 ;
        RECT 131.420 74.040 135.700 74.180 ;
        RECT 138.320 74.040 143.060 74.180 ;
        RECT 131.420 73.840 131.560 74.040 ;
        RECT 124.060 73.700 131.560 73.840 ;
        RECT 131.790 73.840 132.110 73.900 ;
        RECT 135.485 73.840 135.775 73.885 ;
        RECT 136.850 73.840 137.170 73.900 ;
        RECT 138.320 73.885 138.460 74.040 ;
        RECT 131.790 73.700 137.170 73.840 ;
        RECT 114.785 73.655 115.075 73.700 ;
        RECT 119.830 73.640 120.150 73.700 ;
        RECT 131.790 73.640 132.110 73.700 ;
        RECT 135.485 73.655 135.775 73.700 ;
        RECT 136.850 73.640 137.170 73.700 ;
        RECT 138.245 73.655 138.535 73.885 ;
        RECT 22.700 73.020 157.820 73.500 ;
        RECT 34.270 72.820 34.590 72.880 ;
        RECT 44.865 72.820 45.155 72.865 ;
        RECT 45.770 72.820 46.090 72.880 ;
        RECT 34.270 72.680 43.700 72.820 ;
        RECT 34.270 72.620 34.590 72.680 ;
        RECT 38.425 72.480 38.715 72.525 ;
        RECT 39.805 72.480 40.095 72.525 ;
        RECT 41.170 72.480 41.490 72.540 ;
        RECT 38.425 72.340 41.490 72.480 ;
        RECT 43.560 72.480 43.700 72.680 ;
        RECT 44.865 72.680 46.090 72.820 ;
        RECT 44.865 72.635 45.155 72.680 ;
        RECT 45.770 72.620 46.090 72.680 ;
        RECT 52.225 72.635 52.515 72.865 ;
        RECT 57.745 72.820 58.035 72.865 ;
        RECT 60.030 72.820 60.350 72.880 ;
        RECT 68.310 72.820 68.630 72.880 ;
        RECT 56.900 72.680 60.350 72.820 ;
        RECT 52.300 72.480 52.440 72.635 ;
        RECT 43.560 72.340 52.440 72.480 ;
        RECT 38.425 72.295 38.715 72.340 ;
        RECT 39.805 72.295 40.095 72.340 ;
        RECT 41.170 72.280 41.490 72.340 ;
        RECT 54.970 72.280 55.290 72.540 ;
        RECT 37.950 71.940 38.270 72.200 ;
        RECT 39.345 72.140 39.635 72.185 ;
        RECT 40.250 72.140 40.570 72.200 ;
        RECT 39.345 72.000 40.570 72.140 ;
        RECT 39.345 71.955 39.635 72.000 ;
        RECT 40.250 71.940 40.570 72.000 ;
        RECT 40.710 71.940 41.030 72.200 ;
        RECT 41.645 72.140 41.935 72.185 ;
        RECT 43.025 72.140 43.315 72.185 ;
        RECT 41.645 72.000 43.315 72.140 ;
        RECT 41.645 71.955 41.935 72.000 ;
        RECT 43.025 71.955 43.315 72.000 ;
        RECT 50.370 71.940 50.690 72.200 ;
        RECT 51.290 71.940 51.610 72.200 ;
        RECT 54.050 71.940 54.370 72.200 ;
        RECT 54.525 72.140 54.815 72.185 ;
        RECT 55.060 72.140 55.200 72.280 ;
        RECT 54.525 72.000 55.200 72.140 ;
        RECT 54.525 71.955 54.815 72.000 ;
        RECT 43.485 71.800 43.775 71.845 ;
        RECT 50.845 71.800 51.135 71.845 ;
        RECT 52.670 71.800 52.990 71.860 ;
        RECT 43.485 71.660 52.990 71.800 ;
        RECT 43.485 71.615 43.775 71.660 ;
        RECT 50.845 71.615 51.135 71.660 ;
        RECT 52.670 71.600 52.990 71.660 ;
        RECT 53.605 71.800 53.895 71.845 ;
        RECT 54.985 71.800 55.275 71.845 ;
        RECT 53.605 71.660 55.275 71.800 ;
        RECT 53.605 71.615 53.895 71.660 ;
        RECT 54.985 71.615 55.275 71.660 ;
        RECT 37.490 71.460 37.810 71.520 ;
        RECT 46.690 71.460 47.010 71.520 ;
        RECT 56.350 71.460 56.670 71.520 ;
        RECT 37.490 71.320 56.670 71.460 ;
        RECT 37.490 71.260 37.810 71.320 ;
        RECT 46.690 71.260 47.010 71.320 ;
        RECT 56.350 71.260 56.670 71.320 ;
        RECT 43.930 70.920 44.250 71.180 ;
        RECT 54.065 71.120 54.355 71.165 ;
        RECT 56.900 71.120 57.040 72.680 ;
        RECT 57.745 72.635 58.035 72.680 ;
        RECT 60.030 72.620 60.350 72.680 ;
        RECT 66.560 72.680 68.630 72.820 ;
        RECT 59.110 72.480 59.430 72.540 ;
        RECT 63.710 72.480 64.030 72.540 ;
        RECT 57.360 72.340 59.430 72.480 ;
        RECT 57.360 72.185 57.500 72.340 ;
        RECT 59.110 72.280 59.430 72.340 ;
        RECT 61.040 72.340 64.030 72.480 ;
        RECT 57.285 71.955 57.575 72.185 ;
        RECT 58.190 71.940 58.510 72.200 ;
        RECT 61.040 72.185 61.180 72.340 ;
        RECT 63.710 72.280 64.030 72.340 ;
        RECT 60.965 71.955 61.255 72.185 ;
        RECT 61.885 72.140 62.175 72.185 ;
        RECT 62.790 72.140 63.110 72.200 ;
        RECT 61.885 72.000 63.110 72.140 ;
        RECT 61.885 71.955 62.175 72.000 ;
        RECT 62.790 71.940 63.110 72.000 ;
        RECT 65.565 72.140 65.855 72.185 ;
        RECT 66.560 72.140 66.700 72.680 ;
        RECT 68.310 72.620 68.630 72.680 ;
        RECT 70.610 72.620 70.930 72.880 ;
        RECT 81.665 72.820 81.955 72.865 ;
        RECT 83.950 72.820 84.270 72.880 ;
        RECT 81.665 72.680 84.270 72.820 ;
        RECT 81.665 72.635 81.955 72.680 ;
        RECT 83.950 72.620 84.270 72.680 ;
        RECT 89.485 72.820 89.775 72.865 ;
        RECT 90.850 72.820 91.170 72.880 ;
        RECT 89.485 72.680 91.170 72.820 ;
        RECT 89.485 72.635 89.775 72.680 ;
        RECT 90.850 72.620 91.170 72.680 ;
        RECT 97.290 72.865 97.610 72.880 ;
        RECT 97.290 72.635 97.675 72.865 ;
        RECT 97.290 72.620 97.610 72.635 ;
        RECT 99.590 72.620 99.910 72.880 ;
        RECT 102.350 72.620 102.670 72.880 ;
        RECT 106.950 72.820 107.270 72.880 ;
        RECT 111.550 72.820 111.870 72.880 ;
        RECT 114.310 72.820 114.630 72.880 ;
        RECT 106.950 72.680 111.320 72.820 ;
        RECT 106.950 72.620 107.270 72.680 ;
        RECT 83.490 72.480 83.810 72.540 ;
        RECT 95.450 72.480 95.770 72.540 ;
        RECT 96.385 72.480 96.675 72.525 ;
        RECT 67.020 72.340 84.640 72.480 ;
        RECT 67.020 72.185 67.160 72.340 ;
        RECT 83.490 72.280 83.810 72.340 ;
        RECT 65.565 72.000 66.700 72.140 ;
        RECT 65.565 71.955 65.855 72.000 ;
        RECT 66.945 71.955 67.235 72.185 ;
        RECT 74.750 71.940 75.070 72.200 ;
        RECT 75.670 72.140 75.990 72.200 ;
        RECT 79.810 72.140 80.130 72.200 ;
        RECT 82.125 72.140 82.415 72.185 ;
        RECT 75.670 72.000 82.415 72.140 ;
        RECT 75.670 71.940 75.990 72.000 ;
        RECT 79.810 71.940 80.130 72.000 ;
        RECT 66.030 71.800 66.320 71.845 ;
        RECT 68.370 71.800 68.660 71.845 ;
        RECT 66.030 71.660 68.660 71.800 ;
        RECT 74.840 71.800 74.980 71.940 ;
        RECT 79.365 71.800 79.655 71.845 ;
        RECT 74.840 71.660 79.655 71.800 ;
        RECT 66.030 71.615 66.320 71.660 ;
        RECT 68.370 71.615 68.660 71.660 ;
        RECT 79.365 71.615 79.655 71.660 ;
        RECT 66.490 71.460 66.780 71.505 ;
        RECT 67.865 71.460 68.155 71.505 ;
        RECT 66.490 71.320 68.155 71.460 ;
        RECT 66.490 71.275 66.780 71.320 ;
        RECT 67.865 71.275 68.155 71.320 ;
        RECT 54.065 70.980 57.040 71.120 ;
        RECT 60.030 71.120 60.350 71.180 ;
        RECT 61.425 71.120 61.715 71.165 ;
        RECT 60.030 70.980 61.715 71.120 ;
        RECT 54.065 70.935 54.355 70.980 ;
        RECT 60.030 70.920 60.350 70.980 ;
        RECT 61.425 70.935 61.715 70.980 ;
        RECT 75.210 70.920 75.530 71.180 ;
        RECT 79.440 71.120 79.580 71.615 ;
        RECT 80.820 71.505 80.960 72.000 ;
        RECT 82.125 71.955 82.415 72.000 ;
        RECT 83.045 71.955 83.335 72.185 ;
        RECT 80.745 71.275 81.035 71.505 ;
        RECT 83.120 71.120 83.260 71.955 ;
        RECT 84.500 71.800 84.640 72.340 ;
        RECT 95.450 72.340 96.675 72.480 ;
        RECT 99.680 72.480 99.820 72.620 ;
        RECT 105.110 72.480 105.430 72.540 ;
        RECT 99.680 72.340 105.430 72.480 ;
        RECT 95.450 72.280 95.770 72.340 ;
        RECT 96.385 72.295 96.675 72.340 ;
        RECT 105.110 72.280 105.430 72.340 ;
        RECT 109.250 72.280 109.570 72.540 ;
        RECT 111.180 72.525 111.320 72.680 ;
        RECT 111.550 72.680 114.630 72.820 ;
        RECT 111.550 72.620 111.870 72.680 ;
        RECT 114.310 72.620 114.630 72.680 ;
        RECT 119.845 72.820 120.135 72.865 ;
        RECT 122.130 72.820 122.450 72.880 ;
        RECT 119.845 72.680 122.450 72.820 ;
        RECT 119.845 72.635 120.135 72.680 ;
        RECT 122.130 72.620 122.450 72.680 ;
        RECT 129.030 72.620 129.350 72.880 ;
        RECT 145.590 72.820 145.910 72.880 ;
        RECT 147.445 72.820 147.735 72.865 ;
        RECT 145.590 72.680 147.735 72.820 ;
        RECT 145.590 72.620 145.910 72.680 ;
        RECT 147.445 72.635 147.735 72.680 ;
        RECT 111.105 72.295 111.395 72.525 ;
        RECT 113.390 72.480 113.710 72.540 ;
        RECT 123.985 72.480 124.275 72.525 ;
        RECT 126.745 72.480 127.035 72.525 ;
        RECT 113.390 72.340 122.820 72.480 ;
        RECT 113.390 72.280 113.710 72.340 ;
        RECT 87.170 71.940 87.490 72.200 ;
        RECT 88.565 72.140 88.855 72.185 ;
        RECT 90.850 72.140 91.170 72.200 ;
        RECT 88.565 72.000 91.170 72.140 ;
        RECT 88.565 71.955 88.855 72.000 ;
        RECT 90.850 71.940 91.170 72.000 ;
        RECT 96.830 72.140 97.150 72.200 ;
        RECT 98.685 72.140 98.975 72.185 ;
        RECT 96.830 72.000 98.975 72.140 ;
        RECT 96.830 71.940 97.150 72.000 ;
        RECT 98.685 71.955 98.975 72.000 ;
        RECT 101.430 71.940 101.750 72.200 ;
        RECT 113.850 71.940 114.170 72.200 ;
        RECT 114.770 71.940 115.090 72.200 ;
        RECT 115.690 72.140 116.010 72.200 ;
        RECT 117.545 72.140 117.835 72.185 ;
        RECT 115.690 72.000 117.835 72.140 ;
        RECT 115.690 71.940 116.010 72.000 ;
        RECT 117.545 71.955 117.835 72.000 ;
        RECT 120.750 71.940 121.070 72.200 ;
        RECT 122.680 72.185 122.820 72.340 ;
        RECT 123.985 72.340 127.035 72.480 ;
        RECT 123.985 72.295 124.275 72.340 ;
        RECT 126.745 72.295 127.035 72.340 ;
        RECT 135.470 72.480 135.790 72.540 ;
        RECT 138.705 72.480 138.995 72.525 ;
        RECT 135.470 72.340 138.995 72.480 ;
        RECT 135.470 72.280 135.790 72.340 ;
        RECT 138.705 72.295 138.995 72.340 ;
        RECT 139.855 72.310 140.145 72.355 ;
        RECT 122.605 71.955 122.895 72.185 ;
        RECT 88.105 71.800 88.395 71.845 ;
        RECT 91.310 71.800 91.630 71.860 ;
        RECT 84.500 71.660 87.400 71.800 ;
        RECT 79.440 70.980 83.260 71.120 ;
        RECT 83.950 70.920 84.270 71.180 ;
        RECT 87.260 71.165 87.400 71.660 ;
        RECT 88.105 71.660 91.630 71.800 ;
        RECT 88.105 71.615 88.395 71.660 ;
        RECT 91.310 71.600 91.630 71.660 ;
        RECT 109.710 71.800 110.030 71.860 ;
        RECT 110.185 71.800 110.475 71.845 ;
        RECT 110.630 71.800 110.950 71.860 ;
        RECT 112.930 71.800 113.250 71.860 ;
        RECT 116.150 71.800 116.470 71.860 ;
        RECT 109.710 71.660 116.470 71.800 ;
        RECT 109.710 71.600 110.030 71.660 ;
        RECT 110.185 71.615 110.475 71.660 ;
        RECT 110.630 71.600 110.950 71.660 ;
        RECT 112.930 71.600 113.250 71.660 ;
        RECT 116.150 71.600 116.470 71.660 ;
        RECT 98.225 71.460 98.515 71.505 ;
        RECT 101.430 71.460 101.750 71.520 ;
        RECT 98.225 71.320 101.750 71.460 ;
        RECT 98.225 71.275 98.515 71.320 ;
        RECT 101.430 71.260 101.750 71.320 ;
        RECT 111.090 71.460 111.410 71.520 ;
        RECT 112.025 71.460 112.315 71.505 ;
        RECT 111.090 71.320 112.315 71.460 ;
        RECT 111.090 71.260 111.410 71.320 ;
        RECT 112.025 71.275 112.315 71.320 ;
        RECT 114.770 71.460 115.090 71.520 ;
        RECT 118.925 71.460 119.215 71.505 ;
        RECT 114.770 71.320 119.215 71.460 ;
        RECT 122.680 71.460 122.820 71.955 ;
        RECT 123.510 71.940 123.830 72.200 ;
        RECT 124.445 71.955 124.735 72.185 ;
        RECT 128.125 72.140 128.415 72.185 ;
        RECT 132.710 72.140 133.030 72.200 ;
        RECT 128.125 72.000 133.030 72.140 ;
        RECT 128.125 71.955 128.415 72.000 ;
        RECT 123.050 71.800 123.370 71.860 ;
        RECT 124.520 71.800 124.660 71.955 ;
        RECT 132.710 71.940 133.030 72.000 ;
        RECT 135.930 72.140 136.250 72.200 ;
        RECT 137.325 72.140 137.615 72.185 ;
        RECT 139.780 72.140 140.145 72.310 ;
        RECT 135.930 72.125 140.145 72.140 ;
        RECT 135.930 72.000 139.920 72.125 ;
        RECT 135.930 71.940 136.250 72.000 ;
        RECT 137.325 71.955 137.615 72.000 ;
        RECT 143.750 71.940 144.070 72.200 ;
        RECT 123.050 71.660 124.660 71.800 ;
        RECT 127.665 71.800 127.955 71.845 ;
        RECT 134.090 71.800 134.410 71.860 ;
        RECT 136.405 71.800 136.695 71.845 ;
        RECT 127.665 71.660 134.410 71.800 ;
        RECT 123.050 71.600 123.370 71.660 ;
        RECT 127.665 71.615 127.955 71.660 ;
        RECT 134.090 71.600 134.410 71.660 ;
        RECT 134.640 71.660 136.695 71.800 ;
        RECT 128.110 71.460 128.430 71.520 ;
        RECT 122.680 71.320 128.430 71.460 ;
        RECT 114.770 71.260 115.090 71.320 ;
        RECT 118.925 71.275 119.215 71.320 ;
        RECT 128.110 71.260 128.430 71.320 ;
        RECT 134.640 71.180 134.780 71.660 ;
        RECT 136.405 71.615 136.695 71.660 ;
        RECT 141.925 71.800 142.215 71.845 ;
        RECT 142.385 71.800 142.675 71.845 ;
        RECT 141.925 71.660 142.675 71.800 ;
        RECT 141.925 71.615 142.215 71.660 ;
        RECT 142.385 71.615 142.675 71.660 ;
        RECT 142.850 71.800 143.140 71.845 ;
        RECT 145.190 71.800 145.480 71.845 ;
        RECT 142.850 71.660 145.480 71.800 ;
        RECT 142.850 71.615 143.140 71.660 ;
        RECT 145.190 71.615 145.480 71.660 ;
        RECT 136.480 71.460 136.620 71.615 ;
        RECT 143.310 71.460 143.600 71.505 ;
        RECT 144.685 71.460 144.975 71.505 ;
        RECT 136.480 71.320 139.840 71.460 ;
        RECT 87.185 70.935 87.475 71.165 ;
        RECT 97.290 70.920 97.610 71.180 ;
        RECT 101.890 71.120 102.210 71.180 ;
        RECT 102.825 71.120 103.115 71.165 ;
        RECT 101.890 70.980 103.115 71.120 ;
        RECT 101.890 70.920 102.210 70.980 ;
        RECT 102.825 70.935 103.115 70.980 ;
        RECT 122.130 71.120 122.450 71.180 ;
        RECT 122.605 71.120 122.895 71.165 ;
        RECT 123.050 71.120 123.370 71.180 ;
        RECT 122.130 70.980 123.370 71.120 ;
        RECT 122.130 70.920 122.450 70.980 ;
        RECT 122.605 70.935 122.895 70.980 ;
        RECT 123.050 70.920 123.370 70.980 ;
        RECT 126.730 70.920 127.050 71.180 ;
        RECT 130.410 71.120 130.730 71.180 ;
        RECT 134.550 71.120 134.870 71.180 ;
        RECT 130.410 70.980 134.870 71.120 ;
        RECT 130.410 70.920 130.730 70.980 ;
        RECT 134.550 70.920 134.870 70.980 ;
        RECT 138.230 70.920 138.550 71.180 ;
        RECT 139.700 71.165 139.840 71.320 ;
        RECT 143.310 71.320 144.975 71.460 ;
        RECT 143.310 71.275 143.600 71.320 ;
        RECT 144.685 71.275 144.975 71.320 ;
        RECT 139.625 70.935 139.915 71.165 ;
        RECT 140.545 71.120 140.835 71.165 ;
        RECT 145.130 71.120 145.450 71.180 ;
        RECT 140.545 70.980 145.450 71.120 ;
        RECT 140.545 70.935 140.835 70.980 ;
        RECT 145.130 70.920 145.450 70.980 ;
        RECT 22.700 70.300 157.020 70.780 ;
        RECT 41.170 69.900 41.490 70.160 ;
        RECT 42.105 70.100 42.395 70.145 ;
        RECT 43.470 70.100 43.790 70.160 ;
        RECT 42.105 69.960 43.790 70.100 ;
        RECT 42.105 69.915 42.395 69.960 ;
        RECT 43.470 69.900 43.790 69.960 ;
        RECT 43.930 70.100 44.250 70.160 ;
        RECT 45.770 70.100 46.090 70.160 ;
        RECT 43.930 69.960 46.090 70.100 ;
        RECT 43.930 69.900 44.250 69.960 ;
        RECT 45.770 69.900 46.090 69.960 ;
        RECT 53.605 70.100 53.895 70.145 ;
        RECT 54.050 70.100 54.370 70.160 ;
        RECT 53.605 69.960 54.370 70.100 ;
        RECT 53.605 69.915 53.895 69.960 ;
        RECT 54.050 69.900 54.370 69.960 ;
        RECT 69.690 70.100 70.010 70.160 ;
        RECT 72.005 70.100 72.295 70.145 ;
        RECT 74.750 70.100 75.070 70.160 ;
        RECT 69.690 69.960 75.070 70.100 ;
        RECT 69.690 69.900 70.010 69.960 ;
        RECT 72.005 69.915 72.295 69.960 ;
        RECT 74.750 69.900 75.070 69.960 ;
        RECT 83.965 70.100 84.255 70.145 ;
        RECT 87.170 70.100 87.490 70.160 ;
        RECT 83.965 69.960 87.490 70.100 ;
        RECT 83.965 69.915 84.255 69.960 ;
        RECT 87.170 69.900 87.490 69.960 ;
        RECT 88.550 69.900 88.870 70.160 ;
        RECT 91.310 70.100 91.630 70.160 ;
        RECT 94.070 70.100 94.390 70.160 ;
        RECT 91.310 69.960 94.390 70.100 ;
        RECT 91.310 69.900 91.630 69.960 ;
        RECT 94.070 69.900 94.390 69.960 ;
        RECT 95.465 69.915 95.755 70.145 ;
        RECT 96.385 70.100 96.675 70.145 ;
        RECT 96.830 70.100 97.150 70.160 ;
        RECT 96.385 69.960 97.150 70.100 ;
        RECT 96.385 69.915 96.675 69.960 ;
        RECT 37.950 69.760 38.270 69.820 ;
        RECT 43.010 69.760 43.330 69.820 ;
        RECT 47.625 69.760 47.915 69.805 ;
        RECT 37.950 69.620 47.915 69.760 ;
        RECT 37.950 69.560 38.270 69.620 ;
        RECT 43.010 69.560 43.330 69.620 ;
        RECT 47.625 69.575 47.915 69.620 ;
        RECT 50.370 69.760 50.690 69.820 ;
        RECT 60.030 69.760 60.350 69.820 ;
        RECT 50.370 69.620 60.350 69.760 ;
        RECT 50.370 69.560 50.690 69.620 ;
        RECT 60.030 69.560 60.350 69.620 ;
        RECT 67.865 69.760 68.155 69.805 ;
        RECT 71.070 69.760 71.390 69.820 ;
        RECT 67.865 69.620 71.390 69.760 ;
        RECT 67.865 69.575 68.155 69.620 ;
        RECT 71.070 69.560 71.390 69.620 ;
        RECT 80.270 69.760 80.590 69.820 ;
        RECT 93.610 69.760 93.930 69.820 ;
        RECT 95.540 69.760 95.680 69.915 ;
        RECT 96.830 69.900 97.150 69.960 ;
        RECT 98.685 69.915 98.975 70.145 ;
        RECT 108.805 70.100 109.095 70.145 ;
        RECT 112.010 70.100 112.330 70.160 ;
        RECT 113.850 70.100 114.170 70.160 ;
        RECT 108.805 69.960 114.170 70.100 ;
        RECT 108.805 69.915 109.095 69.960 ;
        RECT 97.290 69.760 97.610 69.820 ;
        RECT 98.760 69.760 98.900 69.915 ;
        RECT 112.010 69.900 112.330 69.960 ;
        RECT 113.850 69.900 114.170 69.960 ;
        RECT 120.290 70.100 120.610 70.160 ;
        RECT 129.030 70.100 129.350 70.160 ;
        RECT 120.290 69.960 129.350 70.100 ;
        RECT 120.290 69.900 120.610 69.960 ;
        RECT 129.030 69.900 129.350 69.960 ;
        RECT 129.490 70.100 129.810 70.160 ;
        RECT 130.410 70.100 130.730 70.160 ;
        RECT 129.490 69.960 130.730 70.100 ;
        RECT 129.490 69.900 129.810 69.960 ;
        RECT 130.410 69.900 130.730 69.960 ;
        RECT 131.345 70.100 131.635 70.145 ;
        RECT 132.710 70.100 133.030 70.160 ;
        RECT 131.345 69.960 133.030 70.100 ;
        RECT 131.345 69.915 131.635 69.960 ;
        RECT 132.710 69.900 133.030 69.960 ;
        RECT 134.550 70.100 134.870 70.160 ;
        RECT 135.025 70.100 135.315 70.145 ;
        RECT 136.850 70.100 137.170 70.160 ;
        RECT 139.165 70.100 139.455 70.145 ;
        RECT 134.550 69.960 135.315 70.100 ;
        RECT 134.550 69.900 134.870 69.960 ;
        RECT 135.025 69.915 135.315 69.960 ;
        RECT 135.560 69.960 136.620 70.100 ;
        RECT 80.270 69.620 98.900 69.760 ;
        RECT 102.830 69.760 103.120 69.805 ;
        RECT 104.205 69.760 104.495 69.805 ;
        RECT 102.830 69.620 104.495 69.760 ;
        RECT 80.270 69.560 80.590 69.620 ;
        RECT 42.565 69.420 42.855 69.465 ;
        RECT 51.290 69.420 51.610 69.480 ;
        RECT 75.670 69.420 75.990 69.480 ;
        RECT 83.505 69.420 83.795 69.465 ;
        RECT 40.340 69.280 42.855 69.420 ;
        RECT 35.650 69.080 35.970 69.140 ;
        RECT 36.585 69.080 36.875 69.125 ;
        RECT 35.650 68.940 36.875 69.080 ;
        RECT 35.650 68.880 35.970 68.940 ;
        RECT 36.585 68.895 36.875 68.940 ;
        RECT 37.490 68.880 37.810 69.140 ;
        RECT 40.340 69.125 40.480 69.280 ;
        RECT 42.565 69.235 42.855 69.280 ;
        RECT 43.560 69.280 53.820 69.420 ;
        RECT 43.560 69.125 43.700 69.280 ;
        RECT 40.265 68.895 40.555 69.125 ;
        RECT 40.725 68.895 41.015 69.125 ;
        RECT 43.485 68.895 43.775 69.125 ;
        RECT 37.045 68.740 37.335 68.785 ;
        RECT 40.800 68.740 40.940 68.895 ;
        RECT 43.930 68.880 44.250 69.140 ;
        RECT 44.850 68.880 45.170 69.140 ;
        RECT 45.860 69.125 46.000 69.280 ;
        RECT 51.290 69.220 51.610 69.280 ;
        RECT 45.325 68.895 45.615 69.125 ;
        RECT 45.785 69.080 46.075 69.125 ;
        RECT 46.230 69.080 46.550 69.140 ;
        RECT 45.785 68.940 46.550 69.080 ;
        RECT 45.785 68.895 46.075 68.940 ;
        RECT 33.670 68.600 40.940 68.740 ;
        RECT 45.400 68.740 45.540 68.895 ;
        RECT 46.230 68.880 46.550 68.940 ;
        RECT 46.690 68.880 47.010 69.140 ;
        RECT 52.210 69.125 52.530 69.140 ;
        RECT 53.680 69.125 53.820 69.280 ;
        RECT 68.860 69.280 75.990 69.420 ;
        RECT 48.085 69.080 48.375 69.125 ;
        RECT 49.465 69.080 49.755 69.125 ;
        RECT 52.210 69.080 52.665 69.125 ;
        RECT 48.085 68.940 49.220 69.080 ;
        RECT 48.085 68.895 48.375 68.940 ;
        RECT 47.610 68.740 47.930 68.800 ;
        RECT 45.400 68.600 47.930 68.740 ;
        RECT 25.990 68.400 26.310 68.460 ;
        RECT 33.670 68.400 33.810 68.600 ;
        RECT 37.045 68.555 37.335 68.600 ;
        RECT 47.610 68.540 47.930 68.600 ;
        RECT 25.990 68.260 33.810 68.400 ;
        RECT 49.080 68.400 49.220 68.940 ;
        RECT 49.465 68.940 52.665 69.080 ;
        RECT 49.465 68.895 49.755 68.940 ;
        RECT 52.210 68.895 52.665 68.940 ;
        RECT 53.145 68.895 53.435 69.125 ;
        RECT 53.605 68.895 53.895 69.125 ;
        RECT 52.210 68.880 52.530 68.895 ;
        RECT 53.220 68.740 53.360 68.895 ;
        RECT 54.510 68.880 54.830 69.140 ;
        RECT 58.650 69.080 58.970 69.140 ;
        RECT 59.125 69.080 59.415 69.125 ;
        RECT 58.650 68.940 59.415 69.080 ;
        RECT 58.650 68.880 58.970 68.940 ;
        RECT 59.125 68.895 59.415 68.940 ;
        RECT 59.570 69.080 59.890 69.140 ;
        RECT 60.045 69.080 60.335 69.125 ;
        RECT 59.570 68.940 60.335 69.080 ;
        RECT 59.570 68.880 59.890 68.940 ;
        RECT 60.045 68.895 60.335 68.940 ;
        RECT 61.410 69.080 61.730 69.140 ;
        RECT 61.885 69.080 62.175 69.125 ;
        RECT 61.410 68.940 62.175 69.080 ;
        RECT 61.410 68.880 61.730 68.940 ;
        RECT 61.885 68.895 62.175 68.940 ;
        RECT 58.740 68.740 58.880 68.880 ;
        RECT 68.860 68.785 69.000 69.280 ;
        RECT 73.000 69.125 73.140 69.280 ;
        RECT 75.670 69.220 75.990 69.280 ;
        RECT 78.980 69.280 85.100 69.420 ;
        RECT 72.465 69.080 72.755 69.125 ;
        RECT 72.925 69.080 73.215 69.125 ;
        RECT 72.465 68.940 73.215 69.080 ;
        RECT 72.465 68.895 72.755 68.940 ;
        RECT 72.925 68.895 73.215 68.940 ;
        RECT 73.695 69.080 73.985 69.125 ;
        RECT 74.750 69.080 75.070 69.140 ;
        RECT 73.695 68.940 75.070 69.080 ;
        RECT 73.695 68.895 73.985 68.940 ;
        RECT 74.750 68.880 75.070 68.940 ;
        RECT 76.590 69.080 76.910 69.140 ;
        RECT 77.525 69.080 77.815 69.125 ;
        RECT 76.590 68.940 77.815 69.080 ;
        RECT 76.590 68.880 76.910 68.940 ;
        RECT 77.525 68.895 77.815 68.940 ;
        RECT 78.980 68.800 79.120 69.280 ;
        RECT 83.505 69.235 83.795 69.280 ;
        RECT 79.825 69.080 80.115 69.125 ;
        RECT 80.270 69.080 80.590 69.140 ;
        RECT 82.125 69.080 82.415 69.125 ;
        RECT 79.825 68.940 82.415 69.080 ;
        RECT 79.825 68.895 80.115 68.940 ;
        RECT 80.270 68.880 80.590 68.940 ;
        RECT 82.125 68.895 82.415 68.940 ;
        RECT 82.585 69.080 82.875 69.125 ;
        RECT 83.950 69.080 84.270 69.140 ;
        RECT 84.960 69.125 85.100 69.280 ;
        RECT 82.585 68.940 84.270 69.080 ;
        RECT 82.585 68.895 82.875 68.940 ;
        RECT 83.950 68.880 84.270 68.940 ;
        RECT 84.885 68.895 85.175 69.125 ;
        RECT 85.805 68.895 86.095 69.125 ;
        RECT 86.725 68.895 87.015 69.125 ;
        RECT 53.220 68.600 58.880 68.740 ;
        RECT 53.220 68.400 53.360 68.600 ;
        RECT 68.785 68.555 69.075 68.785 ;
        RECT 69.690 68.540 70.010 68.800 ;
        RECT 70.240 68.600 78.200 68.740 ;
        RECT 49.080 68.260 53.360 68.400 ;
        RECT 25.990 68.200 26.310 68.260 ;
        RECT 59.570 68.200 59.890 68.460 ;
        RECT 68.310 68.400 68.630 68.460 ;
        RECT 70.240 68.445 70.380 68.600 ;
        RECT 78.060 68.460 78.200 68.600 ;
        RECT 78.890 68.540 79.210 68.800 ;
        RECT 85.880 68.740 86.020 68.895 ;
        RECT 81.970 68.600 86.020 68.740 ;
        RECT 86.800 68.740 86.940 68.895 ;
        RECT 87.630 68.880 87.950 69.140 ;
        RECT 88.565 68.895 88.855 69.125 ;
        RECT 89.560 69.080 89.700 69.620 ;
        RECT 93.610 69.560 93.930 69.620 ;
        RECT 97.290 69.560 97.610 69.620 ;
        RECT 102.830 69.575 103.120 69.620 ;
        RECT 104.205 69.575 104.495 69.620 ;
        RECT 106.965 69.760 107.255 69.805 ;
        RECT 108.330 69.760 108.650 69.820 ;
        RECT 106.965 69.620 108.650 69.760 ;
        RECT 106.965 69.575 107.255 69.620 ;
        RECT 108.330 69.560 108.650 69.620 ;
        RECT 119.845 69.760 120.135 69.805 ;
        RECT 123.050 69.760 123.370 69.820 ;
        RECT 119.845 69.620 123.370 69.760 ;
        RECT 119.845 69.575 120.135 69.620 ;
        RECT 123.050 69.560 123.370 69.620 ;
        RECT 123.525 69.760 123.815 69.805 ;
        RECT 135.560 69.760 135.700 69.960 ;
        RECT 123.525 69.620 135.700 69.760 ;
        RECT 123.525 69.575 123.815 69.620 ;
        RECT 135.945 69.575 136.235 69.805 ;
        RECT 136.480 69.760 136.620 69.960 ;
        RECT 136.850 69.960 139.455 70.100 ;
        RECT 136.850 69.900 137.170 69.960 ;
        RECT 139.165 69.915 139.455 69.960 ;
        RECT 139.610 70.100 139.930 70.160 ;
        RECT 141.005 70.100 141.295 70.145 ;
        RECT 139.610 69.960 141.295 70.100 ;
        RECT 139.610 69.900 139.930 69.960 ;
        RECT 141.005 69.915 141.295 69.960 ;
        RECT 141.450 69.900 141.770 70.160 ;
        RECT 143.750 69.900 144.070 70.160 ;
        RECT 136.480 69.620 142.140 69.760 ;
        RECT 96.830 69.220 97.150 69.480 ;
        RECT 101.890 69.220 102.210 69.480 ;
        RECT 102.370 69.420 102.660 69.465 ;
        RECT 104.710 69.420 105.000 69.465 ;
        RECT 102.370 69.280 105.000 69.420 ;
        RECT 102.370 69.235 102.660 69.280 ;
        RECT 104.710 69.235 105.000 69.280 ;
        RECT 109.725 69.420 110.015 69.465 ;
        RECT 110.630 69.420 110.950 69.480 ;
        RECT 114.770 69.420 115.090 69.480 ;
        RECT 118.005 69.420 118.295 69.465 ;
        RECT 109.725 69.280 110.950 69.420 ;
        RECT 109.725 69.235 110.015 69.280 ;
        RECT 110.630 69.220 110.950 69.280 ;
        RECT 113.480 69.280 118.295 69.420 ;
        RECT 90.175 69.080 90.465 69.125 ;
        RECT 89.560 68.940 90.465 69.080 ;
        RECT 90.175 68.895 90.465 68.940 ;
        RECT 90.865 68.895 91.155 69.125 ;
        RECT 88.090 68.740 88.410 68.800 ;
        RECT 88.640 68.740 88.780 68.895 ;
        RECT 89.025 68.740 89.315 68.785 ;
        RECT 86.800 68.600 89.315 68.740 ;
        RECT 70.165 68.400 70.455 68.445 ;
        RECT 68.310 68.260 70.455 68.400 ;
        RECT 68.310 68.200 68.630 68.260 ;
        RECT 70.165 68.215 70.455 68.260 ;
        RECT 70.610 68.400 70.930 68.460 ;
        RECT 74.750 68.400 75.070 68.460 ;
        RECT 70.610 68.260 75.070 68.400 ;
        RECT 70.610 68.200 70.930 68.260 ;
        RECT 74.750 68.200 75.070 68.260 ;
        RECT 77.970 68.400 78.290 68.460 ;
        RECT 81.970 68.400 82.110 68.600 ;
        RECT 88.090 68.540 88.410 68.600 ;
        RECT 89.025 68.555 89.315 68.600 ;
        RECT 89.470 68.740 89.790 68.800 ;
        RECT 90.940 68.740 91.080 68.895 ;
        RECT 91.310 68.880 91.630 69.140 ;
        RECT 92.230 69.080 92.550 69.140 ;
        RECT 93.625 69.080 93.915 69.125 ;
        RECT 92.230 68.940 93.915 69.080 ;
        RECT 92.230 68.880 92.550 68.940 ;
        RECT 93.625 68.895 93.915 68.940 ;
        RECT 99.590 69.080 99.910 69.140 ;
        RECT 100.525 69.080 100.815 69.125 ;
        RECT 99.590 68.940 100.815 69.080 ;
        RECT 99.590 68.880 99.910 68.940 ;
        RECT 100.525 68.895 100.815 68.940 ;
        RECT 103.285 68.895 103.575 69.125 ;
        RECT 104.190 69.080 104.510 69.140 ;
        RECT 113.480 69.125 113.620 69.280 ;
        RECT 114.770 69.220 115.090 69.280 ;
        RECT 118.005 69.235 118.295 69.280 ;
        RECT 122.130 69.420 122.450 69.480 ;
        RECT 123.985 69.420 124.275 69.465 ;
        RECT 129.950 69.420 130.270 69.480 ;
        RECT 132.265 69.420 132.555 69.465 ;
        RECT 134.090 69.420 134.410 69.480 ;
        RECT 122.130 69.280 124.275 69.420 ;
        RECT 122.130 69.220 122.450 69.280 ;
        RECT 123.985 69.235 124.275 69.280 ;
        RECT 127.740 69.280 128.800 69.420 ;
        RECT 107.425 69.080 107.715 69.125 ;
        RECT 111.105 69.080 111.395 69.125 ;
        RECT 113.405 69.080 113.695 69.125 ;
        RECT 104.190 68.940 113.695 69.080 ;
        RECT 89.470 68.600 91.080 68.740 ;
        RECT 95.450 68.740 95.770 68.800 ;
        RECT 98.685 68.740 98.975 68.785 ;
        RECT 103.360 68.740 103.500 68.895 ;
        RECT 104.190 68.880 104.510 68.940 ;
        RECT 107.425 68.895 107.715 68.940 ;
        RECT 111.105 68.895 111.395 68.940 ;
        RECT 113.405 68.895 113.695 68.940 ;
        RECT 113.850 69.080 114.170 69.140 ;
        RECT 115.690 69.080 116.010 69.140 ;
        RECT 118.925 69.080 119.215 69.125 ;
        RECT 113.850 68.940 119.215 69.080 ;
        RECT 113.850 68.880 114.170 68.940 ;
        RECT 115.690 68.880 116.010 68.940 ;
        RECT 118.925 68.895 119.215 68.940 ;
        RECT 120.750 69.080 121.070 69.140 ;
        RECT 122.605 69.080 122.895 69.125 ;
        RECT 127.740 69.080 127.880 69.280 ;
        RECT 120.750 68.940 127.880 69.080 ;
        RECT 120.750 68.880 121.070 68.940 ;
        RECT 122.605 68.895 122.895 68.940 ;
        RECT 128.110 68.880 128.430 69.140 ;
        RECT 128.660 69.125 128.800 69.280 ;
        RECT 129.950 69.280 131.560 69.420 ;
        RECT 129.950 69.220 130.270 69.280 ;
        RECT 128.590 68.895 128.880 69.125 ;
        RECT 129.030 69.080 129.350 69.140 ;
        RECT 131.420 69.125 131.560 69.280 ;
        RECT 132.265 69.280 134.410 69.420 ;
        RECT 132.265 69.235 132.555 69.280 ;
        RECT 134.090 69.220 134.410 69.280 ;
        RECT 130.425 69.080 130.715 69.125 ;
        RECT 129.030 68.940 130.715 69.080 ;
        RECT 95.450 68.600 98.975 68.740 ;
        RECT 89.470 68.540 89.790 68.600 ;
        RECT 95.450 68.540 95.770 68.600 ;
        RECT 98.685 68.555 98.975 68.600 ;
        RECT 101.520 68.600 103.500 68.740 ;
        RECT 77.970 68.260 82.110 68.400 ;
        RECT 77.970 68.200 78.290 68.260 ;
        RECT 83.490 68.200 83.810 68.460 ;
        RECT 86.265 68.400 86.555 68.445 ;
        RECT 90.850 68.400 91.170 68.460 ;
        RECT 86.265 68.260 91.170 68.400 ;
        RECT 86.265 68.215 86.555 68.260 ;
        RECT 90.850 68.200 91.170 68.260 ;
        RECT 99.605 68.400 99.895 68.445 ;
        RECT 100.510 68.400 100.830 68.460 ;
        RECT 101.520 68.445 101.660 68.600 ;
        RECT 112.010 68.540 112.330 68.800 ;
        RECT 115.245 68.555 115.535 68.785 ;
        RECT 128.660 68.740 128.800 68.895 ;
        RECT 129.030 68.880 129.350 68.940 ;
        RECT 130.425 68.895 130.715 68.940 ;
        RECT 131.345 69.080 131.635 69.125 ;
        RECT 131.805 69.080 132.095 69.125 ;
        RECT 132.725 69.080 133.015 69.125 ;
        RECT 133.185 69.080 133.475 69.125 ;
        RECT 131.345 68.940 132.095 69.080 ;
        RECT 131.345 68.895 131.635 68.940 ;
        RECT 131.805 68.895 132.095 68.940 ;
        RECT 132.340 68.940 133.475 69.080 ;
        RECT 136.020 69.080 136.160 69.575 ;
        RECT 142.000 69.465 142.140 69.620 ;
        RECT 141.925 69.235 142.215 69.465 ;
        RECT 146.510 69.420 146.830 69.480 ;
        RECT 142.460 69.280 146.830 69.420 ;
        RECT 137.325 69.080 137.615 69.125 ;
        RECT 136.020 68.940 137.615 69.080 ;
        RECT 129.490 68.740 129.810 68.800 ;
        RECT 128.660 68.600 129.810 68.740 ;
        RECT 99.605 68.260 100.830 68.400 ;
        RECT 99.605 68.215 99.895 68.260 ;
        RECT 100.510 68.200 100.830 68.260 ;
        RECT 101.445 68.215 101.735 68.445 ;
        RECT 110.170 68.200 110.490 68.460 ;
        RECT 113.850 68.400 114.170 68.460 ;
        RECT 115.320 68.400 115.460 68.555 ;
        RECT 129.490 68.540 129.810 68.600 ;
        RECT 121.670 68.400 121.990 68.460 ;
        RECT 132.340 68.400 132.480 68.940 ;
        RECT 132.725 68.895 133.015 68.940 ;
        RECT 133.185 68.895 133.475 68.940 ;
        RECT 137.325 68.895 137.615 68.940 ;
        RECT 138.230 69.080 138.550 69.140 ;
        RECT 139.165 69.080 139.455 69.125 ;
        RECT 138.230 68.940 139.455 69.080 ;
        RECT 138.230 68.880 138.550 68.940 ;
        RECT 139.165 68.895 139.455 68.940 ;
        RECT 140.085 68.895 140.375 69.125 ;
        RECT 140.990 69.080 141.310 69.140 ;
        RECT 141.465 69.080 141.755 69.125 ;
        RECT 140.990 68.940 141.755 69.080 ;
        RECT 135.025 68.740 135.315 68.785 ;
        RECT 135.470 68.740 135.790 68.800 ;
        RECT 140.160 68.740 140.300 68.895 ;
        RECT 140.990 68.880 141.310 68.940 ;
        RECT 141.465 68.895 141.755 68.940 ;
        RECT 142.460 68.740 142.600 69.280 ;
        RECT 146.510 69.220 146.830 69.280 ;
        RECT 144.685 69.080 144.975 69.125 ;
        RECT 135.025 68.600 135.790 68.740 ;
        RECT 135.025 68.555 135.315 68.600 ;
        RECT 135.470 68.540 135.790 68.600 ;
        RECT 138.320 68.600 142.600 68.740 ;
        RECT 143.380 68.940 144.975 69.080 ;
        RECT 138.320 68.445 138.460 68.600 ;
        RECT 143.380 68.445 143.520 68.940 ;
        RECT 144.685 68.895 144.975 68.940 ;
        RECT 145.130 68.880 145.450 69.140 ;
        RECT 113.850 68.260 132.480 68.400 ;
        RECT 113.850 68.200 114.170 68.260 ;
        RECT 121.670 68.200 121.990 68.260 ;
        RECT 138.245 68.215 138.535 68.445 ;
        RECT 143.305 68.215 143.595 68.445 ;
        RECT 145.590 68.400 145.910 68.460 ;
        RECT 146.065 68.400 146.355 68.445 ;
        RECT 145.590 68.260 146.355 68.400 ;
        RECT 145.590 68.200 145.910 68.260 ;
        RECT 146.065 68.215 146.355 68.260 ;
        RECT 22.700 67.580 157.820 68.060 ;
        RECT 43.930 67.380 44.250 67.440 ;
        RECT 44.405 67.380 44.695 67.425 ;
        RECT 59.585 67.380 59.875 67.425 ;
        RECT 60.490 67.380 60.810 67.440 ;
        RECT 84.410 67.380 84.730 67.440 ;
        RECT 43.930 67.240 44.695 67.380 ;
        RECT 43.930 67.180 44.250 67.240 ;
        RECT 44.405 67.195 44.695 67.240 ;
        RECT 44.940 67.240 54.740 67.380 ;
        RECT 37.965 67.040 38.255 67.085 ;
        RECT 33.670 66.900 38.255 67.040 ;
        RECT 32.905 66.700 33.195 66.745 ;
        RECT 33.670 66.700 33.810 66.900 ;
        RECT 37.965 66.855 38.255 66.900 ;
        RECT 42.640 66.900 44.160 67.040 ;
        RECT 42.640 66.760 42.780 66.900 ;
        RECT 32.905 66.560 33.810 66.700 ;
        RECT 32.905 66.515 33.195 66.560 ;
        RECT 37.030 66.500 37.350 66.760 ;
        RECT 37.505 66.515 37.795 66.745 ;
        RECT 38.425 66.700 38.715 66.745 ;
        RECT 40.250 66.700 40.570 66.760 ;
        RECT 38.425 66.560 40.570 66.700 ;
        RECT 38.425 66.515 38.715 66.560 ;
        RECT 31.065 66.360 31.355 66.405 ;
        RECT 31.525 66.360 31.815 66.405 ;
        RECT 31.065 66.220 31.815 66.360 ;
        RECT 31.065 66.175 31.355 66.220 ;
        RECT 31.525 66.175 31.815 66.220 ;
        RECT 31.990 66.360 32.280 66.405 ;
        RECT 34.330 66.360 34.620 66.405 ;
        RECT 31.990 66.220 34.620 66.360 ;
        RECT 31.990 66.175 32.280 66.220 ;
        RECT 34.330 66.175 34.620 66.220 ;
        RECT 35.650 66.360 35.970 66.420 ;
        RECT 37.580 66.360 37.720 66.515 ;
        RECT 40.250 66.500 40.570 66.560 ;
        RECT 42.550 66.500 42.870 66.760 ;
        RECT 43.470 66.500 43.790 66.760 ;
        RECT 43.560 66.360 43.700 66.500 ;
        RECT 35.650 66.220 43.700 66.360 ;
        RECT 44.020 66.360 44.160 66.900 ;
        RECT 44.390 66.700 44.710 66.760 ;
        RECT 44.940 66.745 45.080 67.240 ;
        RECT 54.600 67.100 54.740 67.240 ;
        RECT 59.585 67.240 60.810 67.380 ;
        RECT 59.585 67.195 59.875 67.240 ;
        RECT 60.490 67.180 60.810 67.240 ;
        RECT 75.760 67.240 89.700 67.380 ;
        RECT 50.370 67.040 50.690 67.100 ;
        RECT 45.860 66.900 50.690 67.040 ;
        RECT 44.865 66.700 45.155 66.745 ;
        RECT 44.390 66.560 45.155 66.700 ;
        RECT 44.390 66.500 44.710 66.560 ;
        RECT 44.865 66.515 45.155 66.560 ;
        RECT 45.860 66.360 46.000 66.900 ;
        RECT 50.370 66.840 50.690 66.900 ;
        RECT 54.050 66.840 54.370 67.100 ;
        RECT 54.510 66.840 54.830 67.100 ;
        RECT 60.580 67.040 60.720 67.180 ;
        RECT 57.360 66.900 58.880 67.040 ;
        RECT 60.580 66.900 62.100 67.040 ;
        RECT 46.230 66.700 46.550 66.760 ;
        RECT 47.165 66.700 47.455 66.745 ;
        RECT 46.230 66.560 47.455 66.700 ;
        RECT 46.230 66.500 46.550 66.560 ;
        RECT 47.165 66.515 47.455 66.560 ;
        RECT 48.085 66.515 48.375 66.745 ;
        RECT 49.005 66.700 49.295 66.745 ;
        RECT 50.830 66.700 51.150 66.760 ;
        RECT 49.005 66.560 51.150 66.700 ;
        RECT 49.005 66.515 49.295 66.560 ;
        RECT 44.020 66.220 46.000 66.360 ;
        RECT 48.160 66.360 48.300 66.515 ;
        RECT 50.830 66.500 51.150 66.560 ;
        RECT 53.145 66.700 53.435 66.745 ;
        RECT 54.140 66.700 54.280 66.840 ;
        RECT 53.145 66.560 54.280 66.700 ;
        RECT 54.600 66.700 54.740 66.840 ;
        RECT 57.360 66.745 57.500 66.900 ;
        RECT 56.365 66.700 56.655 66.745 ;
        RECT 54.600 66.560 56.655 66.700 ;
        RECT 53.145 66.515 53.435 66.560 ;
        RECT 56.365 66.515 56.655 66.560 ;
        RECT 57.285 66.515 57.575 66.745 ;
        RECT 57.730 66.500 58.050 66.760 ;
        RECT 58.740 66.745 58.880 66.900 ;
        RECT 58.665 66.700 58.955 66.745 ;
        RECT 59.125 66.700 59.415 66.745 ;
        RECT 59.570 66.700 59.890 66.760 ;
        RECT 58.665 66.560 59.890 66.700 ;
        RECT 58.665 66.515 58.955 66.560 ;
        RECT 59.125 66.515 59.415 66.560 ;
        RECT 59.570 66.500 59.890 66.560 ;
        RECT 60.030 66.500 60.350 66.760 ;
        RECT 60.505 66.700 60.795 66.745 ;
        RECT 61.410 66.700 61.730 66.760 ;
        RECT 61.960 66.745 62.100 66.900 ;
        RECT 69.780 66.900 72.220 67.040 ;
        RECT 60.505 66.560 61.730 66.700 ;
        RECT 60.505 66.515 60.795 66.560 ;
        RECT 61.410 66.500 61.730 66.560 ;
        RECT 61.885 66.515 62.175 66.745 ;
        RECT 66.025 66.700 66.315 66.745 ;
        RECT 67.390 66.700 67.710 66.760 ;
        RECT 66.025 66.560 67.710 66.700 ;
        RECT 66.025 66.515 66.315 66.560 ;
        RECT 67.390 66.500 67.710 66.560 ;
        RECT 68.310 66.500 68.630 66.760 ;
        RECT 69.780 66.745 69.920 66.900 ;
        RECT 69.245 66.700 69.535 66.745 ;
        RECT 69.705 66.700 69.995 66.745 ;
        RECT 69.245 66.560 69.995 66.700 ;
        RECT 69.245 66.515 69.535 66.560 ;
        RECT 69.705 66.515 69.995 66.560 ;
        RECT 70.610 66.500 70.930 66.760 ;
        RECT 71.070 66.500 71.390 66.760 ;
        RECT 72.080 66.745 72.220 66.900 ;
        RECT 72.005 66.700 72.295 66.745 ;
        RECT 74.765 66.700 75.055 66.745 ;
        RECT 72.005 66.560 75.055 66.700 ;
        RECT 72.005 66.515 72.295 66.560 ;
        RECT 74.765 66.515 75.055 66.560 ;
        RECT 75.210 66.700 75.530 66.760 ;
        RECT 75.760 66.745 75.900 67.240 ;
        RECT 84.410 67.180 84.730 67.240 ;
        RECT 77.600 66.900 79.120 67.040 ;
        RECT 77.600 66.745 77.740 66.900 ;
        RECT 78.980 66.760 79.120 66.900 ;
        RECT 75.685 66.700 75.975 66.745 ;
        RECT 75.210 66.560 75.975 66.700 ;
        RECT 49.910 66.360 50.230 66.420 ;
        RECT 48.160 66.220 50.230 66.360 ;
        RECT 35.650 66.160 35.970 66.220 ;
        RECT 32.450 66.020 32.740 66.065 ;
        RECT 33.870 66.020 34.160 66.065 ;
        RECT 32.450 65.880 34.160 66.020 ;
        RECT 32.450 65.835 32.740 65.880 ;
        RECT 33.870 65.835 34.160 65.880 ;
        RECT 40.250 66.020 40.570 66.080 ;
        RECT 48.160 66.020 48.300 66.220 ;
        RECT 49.910 66.160 50.230 66.220 ;
        RECT 51.720 66.360 52.010 66.405 ;
        RECT 54.060 66.360 54.350 66.405 ;
        RECT 51.720 66.220 54.350 66.360 ;
        RECT 51.720 66.175 52.010 66.220 ;
        RECT 54.060 66.175 54.350 66.220 ;
        RECT 54.510 66.160 54.830 66.420 ;
        RECT 54.970 66.360 55.290 66.420 ;
        RECT 56.825 66.360 57.115 66.405 ;
        RECT 54.970 66.220 57.115 66.360 ;
        RECT 54.970 66.160 55.290 66.220 ;
        RECT 56.825 66.175 57.115 66.220 ;
        RECT 60.970 66.360 61.260 66.405 ;
        RECT 63.310 66.360 63.600 66.405 ;
        RECT 60.970 66.220 63.600 66.360 ;
        RECT 60.970 66.175 61.260 66.220 ;
        RECT 63.310 66.175 63.600 66.220 ;
        RECT 40.250 65.880 48.300 66.020 ;
        RECT 52.180 66.020 52.470 66.065 ;
        RECT 53.600 66.020 53.890 66.065 ;
        RECT 52.180 65.880 53.890 66.020 ;
        RECT 40.250 65.820 40.570 65.880 ;
        RECT 52.180 65.835 52.470 65.880 ;
        RECT 53.600 65.835 53.890 65.880 ;
        RECT 61.430 66.020 61.720 66.065 ;
        RECT 62.850 66.020 63.140 66.065 ;
        RECT 61.430 65.880 63.140 66.020 ;
        RECT 71.160 66.020 71.300 66.500 ;
        RECT 74.840 66.360 74.980 66.515 ;
        RECT 75.210 66.500 75.530 66.560 ;
        RECT 75.685 66.515 75.975 66.560 ;
        RECT 76.605 66.515 76.895 66.745 ;
        RECT 77.525 66.515 77.815 66.745 ;
        RECT 76.130 66.360 76.450 66.420 ;
        RECT 74.840 66.220 76.450 66.360 ;
        RECT 76.130 66.160 76.450 66.220 ;
        RECT 76.680 66.360 76.820 66.515 ;
        RECT 77.970 66.500 78.290 66.760 ;
        RECT 78.890 66.500 79.210 66.760 ;
        RECT 89.560 66.745 89.700 67.240 ;
        RECT 99.590 67.180 99.910 67.440 ;
        RECT 110.630 67.380 110.950 67.440 ;
        RECT 120.290 67.380 120.610 67.440 ;
        RECT 110.630 67.240 120.610 67.380 ;
        RECT 110.630 67.180 110.950 67.240 ;
        RECT 120.290 67.180 120.610 67.240 ;
        RECT 135.025 67.380 135.315 67.425 ;
        RECT 135.470 67.380 135.790 67.440 ;
        RECT 135.025 67.240 135.790 67.380 ;
        RECT 135.025 67.195 135.315 67.240 ;
        RECT 135.470 67.180 135.790 67.240 ;
        RECT 135.945 67.195 136.235 67.425 ;
        RECT 138.705 67.380 138.995 67.425 ;
        RECT 141.450 67.380 141.770 67.440 ;
        RECT 138.705 67.240 141.770 67.380 ;
        RECT 138.705 67.195 138.995 67.240 ;
        RECT 89.945 67.040 90.235 67.085 ;
        RECT 110.170 67.040 110.490 67.100 ;
        RECT 122.130 67.040 122.450 67.100 ;
        RECT 89.945 66.900 97.980 67.040 ;
        RECT 89.945 66.855 90.235 66.900 ;
        RECT 89.485 66.515 89.775 66.745 ;
        RECT 90.405 66.700 90.695 66.745 ;
        RECT 91.310 66.700 91.630 66.760 ;
        RECT 90.405 66.560 91.630 66.700 ;
        RECT 90.405 66.515 90.695 66.560 ;
        RECT 87.630 66.360 87.950 66.420 ;
        RECT 76.680 66.220 87.950 66.360 ;
        RECT 76.680 66.020 76.820 66.220 ;
        RECT 87.630 66.160 87.950 66.220 ;
        RECT 88.090 66.360 88.410 66.420 ;
        RECT 90.480 66.360 90.620 66.515 ;
        RECT 91.310 66.500 91.630 66.560 ;
        RECT 97.290 66.700 97.610 66.760 ;
        RECT 97.840 66.745 97.980 66.900 ;
        RECT 108.420 66.900 110.490 67.040 ;
        RECT 97.765 66.700 98.055 66.745 ;
        RECT 97.290 66.560 98.055 66.700 ;
        RECT 97.290 66.500 97.610 66.560 ;
        RECT 97.765 66.515 98.055 66.560 ;
        RECT 100.510 66.500 100.830 66.760 ;
        RECT 101.430 66.700 101.750 66.760 ;
        RECT 108.420 66.745 108.560 66.900 ;
        RECT 110.170 66.840 110.490 66.900 ;
        RECT 119.920 66.900 123.740 67.040 ;
        RECT 101.905 66.700 102.195 66.745 ;
        RECT 101.430 66.560 102.195 66.700 ;
        RECT 101.430 66.500 101.750 66.560 ;
        RECT 101.905 66.515 102.195 66.560 ;
        RECT 108.345 66.515 108.635 66.745 ;
        RECT 109.265 66.700 109.555 66.745 ;
        RECT 109.710 66.700 110.030 66.760 ;
        RECT 109.265 66.560 110.030 66.700 ;
        RECT 109.265 66.515 109.555 66.560 ;
        RECT 109.710 66.500 110.030 66.560 ;
        RECT 110.630 66.500 110.950 66.760 ;
        RECT 112.930 66.500 113.250 66.760 ;
        RECT 113.850 66.500 114.170 66.760 ;
        RECT 114.325 66.515 114.615 66.745 ;
        RECT 114.770 66.700 115.090 66.760 ;
        RECT 119.920 66.745 120.060 66.900 ;
        RECT 115.245 66.700 115.535 66.745 ;
        RECT 114.770 66.560 115.535 66.700 ;
        RECT 88.090 66.220 90.620 66.360 ;
        RECT 88.090 66.160 88.410 66.220 ;
        RECT 98.225 66.175 98.515 66.405 ;
        RECT 113.020 66.360 113.160 66.500 ;
        RECT 114.400 66.360 114.540 66.515 ;
        RECT 114.770 66.500 115.090 66.560 ;
        RECT 115.245 66.515 115.535 66.560 ;
        RECT 118.925 66.515 119.215 66.745 ;
        RECT 119.845 66.515 120.135 66.745 ;
        RECT 113.020 66.220 114.540 66.360 ;
        RECT 71.160 65.880 76.820 66.020 ;
        RECT 83.490 66.020 83.810 66.080 ;
        RECT 98.300 66.020 98.440 66.175 ;
        RECT 83.490 65.880 98.440 66.020 ;
        RECT 110.170 66.020 110.490 66.080 ;
        RECT 119.000 66.020 119.140 66.515 ;
        RECT 120.290 66.500 120.610 66.760 ;
        RECT 121.300 66.745 121.440 66.900 ;
        RECT 122.130 66.840 122.450 66.900 ;
        RECT 123.600 66.760 123.740 66.900 ;
        RECT 130.500 66.900 132.020 67.040 ;
        RECT 121.225 66.515 121.515 66.745 ;
        RECT 121.670 66.700 121.990 66.760 ;
        RECT 123.065 66.700 123.355 66.745 ;
        RECT 121.670 66.560 123.355 66.700 ;
        RECT 121.670 66.500 121.990 66.560 ;
        RECT 123.065 66.515 123.355 66.560 ;
        RECT 123.510 66.700 123.830 66.760 ;
        RECT 123.985 66.700 124.275 66.745 ;
        RECT 123.510 66.560 124.275 66.700 ;
        RECT 123.510 66.500 123.830 66.560 ;
        RECT 123.985 66.515 124.275 66.560 ;
        RECT 129.505 66.515 129.795 66.745 ;
        RECT 129.950 66.700 130.270 66.760 ;
        RECT 130.500 66.745 130.640 66.900 ;
        RECT 130.425 66.700 130.715 66.745 ;
        RECT 129.950 66.560 130.715 66.700 ;
        RECT 129.580 66.360 129.720 66.515 ;
        RECT 129.950 66.500 130.270 66.560 ;
        RECT 130.425 66.515 130.715 66.560 ;
        RECT 130.885 66.700 131.175 66.745 ;
        RECT 131.330 66.700 131.650 66.760 ;
        RECT 131.880 66.745 132.020 66.900 ;
        RECT 130.885 66.560 131.650 66.700 ;
        RECT 130.885 66.515 131.175 66.560 ;
        RECT 131.330 66.500 131.650 66.560 ;
        RECT 131.805 66.515 132.095 66.745 ;
        RECT 136.020 66.700 136.160 67.195 ;
        RECT 141.450 67.180 141.770 67.240 ;
        RECT 137.785 66.700 138.075 66.745 ;
        RECT 136.020 66.560 138.075 66.700 ;
        RECT 137.785 66.515 138.075 66.560 ;
        RECT 133.185 66.360 133.475 66.405 ;
        RECT 129.580 66.220 133.475 66.360 ;
        RECT 129.580 66.020 129.720 66.220 ;
        RECT 133.185 66.175 133.475 66.220 ;
        RECT 110.170 65.880 129.720 66.020 ;
        RECT 130.425 66.020 130.715 66.065 ;
        RECT 130.870 66.020 131.190 66.080 ;
        RECT 130.425 65.880 131.190 66.020 ;
        RECT 61.430 65.835 61.720 65.880 ;
        RECT 62.850 65.835 63.140 65.880 ;
        RECT 83.490 65.820 83.810 65.880 ;
        RECT 110.170 65.820 110.490 65.880 ;
        RECT 130.425 65.835 130.715 65.880 ;
        RECT 130.870 65.820 131.190 65.880 ;
        RECT 131.805 66.020 132.095 66.065 ;
        RECT 138.230 66.020 138.550 66.080 ;
        RECT 140.990 66.020 141.310 66.080 ;
        RECT 131.805 65.880 141.310 66.020 ;
        RECT 131.805 65.835 132.095 65.880 ;
        RECT 138.230 65.820 138.550 65.880 ;
        RECT 140.990 65.820 141.310 65.880 ;
        RECT 40.710 65.680 41.030 65.740 ;
        RECT 42.565 65.680 42.855 65.725 ;
        RECT 44.850 65.680 45.170 65.740 ;
        RECT 40.710 65.540 45.170 65.680 ;
        RECT 40.710 65.480 41.030 65.540 ;
        RECT 42.565 65.495 42.855 65.540 ;
        RECT 44.850 65.480 45.170 65.540 ;
        RECT 47.610 65.680 47.930 65.740 ;
        RECT 48.085 65.680 48.375 65.725 ;
        RECT 49.450 65.680 49.770 65.740 ;
        RECT 47.610 65.540 49.770 65.680 ;
        RECT 47.610 65.480 47.930 65.540 ;
        RECT 48.085 65.495 48.375 65.540 ;
        RECT 49.450 65.480 49.770 65.540 ;
        RECT 51.290 65.680 51.610 65.740 ;
        RECT 54.985 65.680 55.275 65.725 ;
        RECT 51.290 65.540 55.275 65.680 ;
        RECT 51.290 65.480 51.610 65.540 ;
        RECT 54.985 65.495 55.275 65.540 ;
        RECT 58.665 65.680 58.955 65.725 ;
        RECT 60.950 65.680 61.270 65.740 ;
        RECT 58.665 65.540 61.270 65.680 ;
        RECT 58.665 65.495 58.955 65.540 ;
        RECT 60.950 65.480 61.270 65.540 ;
        RECT 68.310 65.480 68.630 65.740 ;
        RECT 69.690 65.680 70.010 65.740 ;
        RECT 70.625 65.680 70.915 65.725 ;
        RECT 69.690 65.540 70.915 65.680 ;
        RECT 69.690 65.480 70.010 65.540 ;
        RECT 70.625 65.495 70.915 65.540 ;
        RECT 71.070 65.480 71.390 65.740 ;
        RECT 75.685 65.680 75.975 65.725 ;
        RECT 76.130 65.680 76.450 65.740 ;
        RECT 75.685 65.540 76.450 65.680 ;
        RECT 75.685 65.495 75.975 65.540 ;
        RECT 76.130 65.480 76.450 65.540 ;
        RECT 76.590 65.680 76.910 65.740 ;
        RECT 77.525 65.680 77.815 65.725 ;
        RECT 76.590 65.540 77.815 65.680 ;
        RECT 76.590 65.480 76.910 65.540 ;
        RECT 77.525 65.495 77.815 65.540 ;
        RECT 78.905 65.680 79.195 65.725 ;
        RECT 79.350 65.680 79.670 65.740 ;
        RECT 78.905 65.540 79.670 65.680 ;
        RECT 78.905 65.495 79.195 65.540 ;
        RECT 79.350 65.480 79.670 65.540 ;
        RECT 81.190 65.680 81.510 65.740 ;
        RECT 81.665 65.680 81.955 65.725 ;
        RECT 81.190 65.540 81.955 65.680 ;
        RECT 81.190 65.480 81.510 65.540 ;
        RECT 81.665 65.495 81.955 65.540 ;
        RECT 95.910 65.680 96.230 65.740 ;
        RECT 96.385 65.680 96.675 65.725 ;
        RECT 95.910 65.540 96.675 65.680 ;
        RECT 95.910 65.480 96.230 65.540 ;
        RECT 96.385 65.495 96.675 65.540 ;
        RECT 98.685 65.680 98.975 65.725 ;
        RECT 101.430 65.680 101.750 65.740 ;
        RECT 98.685 65.540 101.750 65.680 ;
        RECT 98.685 65.495 98.975 65.540 ;
        RECT 101.430 65.480 101.750 65.540 ;
        RECT 102.810 65.480 103.130 65.740 ;
        RECT 108.330 65.480 108.650 65.740 ;
        RECT 110.645 65.680 110.935 65.725 ;
        RECT 112.470 65.680 112.790 65.740 ;
        RECT 110.645 65.540 112.790 65.680 ;
        RECT 110.645 65.495 110.935 65.540 ;
        RECT 112.470 65.480 112.790 65.540 ;
        RECT 113.865 65.680 114.155 65.725 ;
        RECT 114.770 65.680 115.090 65.740 ;
        RECT 113.865 65.540 115.090 65.680 ;
        RECT 113.865 65.495 114.155 65.540 ;
        RECT 114.770 65.480 115.090 65.540 ;
        RECT 115.230 65.480 115.550 65.740 ;
        RECT 118.910 65.680 119.230 65.740 ;
        RECT 119.845 65.680 120.135 65.725 ;
        RECT 118.910 65.540 120.135 65.680 ;
        RECT 118.910 65.480 119.230 65.540 ;
        RECT 119.845 65.495 120.135 65.540 ;
        RECT 121.210 65.480 121.530 65.740 ;
        RECT 123.985 65.680 124.275 65.725 ;
        RECT 127.650 65.680 127.970 65.740 ;
        RECT 123.985 65.540 127.970 65.680 ;
        RECT 123.985 65.495 124.275 65.540 ;
        RECT 127.650 65.480 127.970 65.540 ;
        RECT 135.010 65.480 135.330 65.740 ;
        RECT 22.700 64.860 157.020 65.340 ;
        RECT 49.910 64.660 50.230 64.720 ;
        RECT 44.020 64.520 50.230 64.660 ;
        RECT 25.550 64.320 25.840 64.365 ;
        RECT 26.970 64.320 27.260 64.365 ;
        RECT 25.550 64.180 27.260 64.320 ;
        RECT 25.550 64.135 25.840 64.180 ;
        RECT 26.970 64.135 27.260 64.180 ;
        RECT 25.090 63.980 25.380 64.025 ;
        RECT 27.430 63.980 27.720 64.025 ;
        RECT 43.470 63.980 43.790 64.040 ;
        RECT 25.090 63.840 27.720 63.980 ;
        RECT 25.090 63.795 25.380 63.840 ;
        RECT 27.430 63.795 27.720 63.840 ;
        RECT 33.900 63.840 43.790 63.980 ;
        RECT 24.610 63.440 24.930 63.700 ;
        RECT 26.005 63.455 26.295 63.685 ;
        RECT 28.750 63.640 29.070 63.700 ;
        RECT 30.145 63.640 30.435 63.685 ;
        RECT 28.750 63.500 30.435 63.640 ;
        RECT 26.080 63.300 26.220 63.455 ;
        RECT 28.750 63.440 29.070 63.500 ;
        RECT 30.145 63.455 30.435 63.500 ;
        RECT 30.590 63.440 30.910 63.700 ;
        RECT 33.900 63.685 34.040 63.840 ;
        RECT 33.825 63.455 34.115 63.685 ;
        RECT 34.745 63.640 35.035 63.685 ;
        RECT 35.650 63.640 35.970 63.700 ;
        RECT 36.200 63.685 36.340 63.840 ;
        RECT 43.470 63.780 43.790 63.840 ;
        RECT 34.745 63.500 35.970 63.640 ;
        RECT 34.745 63.455 35.035 63.500 ;
        RECT 35.650 63.440 35.970 63.500 ;
        RECT 36.125 63.455 36.415 63.685 ;
        RECT 37.045 63.455 37.335 63.685 ;
        RECT 34.285 63.300 34.575 63.345 ;
        RECT 26.080 63.160 34.575 63.300 ;
        RECT 37.120 63.300 37.260 63.455 ;
        RECT 37.490 63.440 37.810 63.700 ;
        RECT 38.425 63.455 38.715 63.685 ;
        RECT 38.500 63.300 38.640 63.455 ;
        RECT 41.170 63.440 41.490 63.700 ;
        RECT 41.645 63.455 41.935 63.685 ;
        RECT 41.720 63.300 41.860 63.455 ;
        RECT 42.550 63.440 42.870 63.700 ;
        RECT 43.010 63.440 43.330 63.700 ;
        RECT 44.020 63.685 44.160 64.520 ;
        RECT 49.910 64.460 50.230 64.520 ;
        RECT 74.750 64.660 75.070 64.720 ;
        RECT 114.310 64.660 114.630 64.720 ;
        RECT 131.330 64.660 131.650 64.720 ;
        RECT 74.750 64.520 82.110 64.660 ;
        RECT 74.750 64.460 75.070 64.520 ;
        RECT 46.250 64.320 46.540 64.365 ;
        RECT 47.670 64.320 47.960 64.365 ;
        RECT 46.250 64.180 47.960 64.320 ;
        RECT 46.250 64.135 46.540 64.180 ;
        RECT 47.670 64.135 47.960 64.180 ;
        RECT 52.230 64.320 52.520 64.365 ;
        RECT 53.650 64.320 53.940 64.365 ;
        RECT 52.230 64.180 53.940 64.320 ;
        RECT 52.230 64.135 52.520 64.180 ;
        RECT 53.650 64.135 53.940 64.180 ;
        RECT 54.510 64.320 54.830 64.380 ;
        RECT 57.285 64.320 57.575 64.365 ;
        RECT 54.510 64.180 57.575 64.320 ;
        RECT 54.510 64.120 54.830 64.180 ;
        RECT 57.285 64.135 57.575 64.180 ;
        RECT 66.030 64.320 66.320 64.365 ;
        RECT 67.450 64.320 67.740 64.365 ;
        RECT 66.030 64.180 67.740 64.320 ;
        RECT 66.030 64.135 66.320 64.180 ;
        RECT 67.450 64.135 67.740 64.180 ;
        RECT 78.910 64.320 79.200 64.365 ;
        RECT 80.330 64.320 80.620 64.365 ;
        RECT 78.910 64.180 80.620 64.320 ;
        RECT 78.910 64.135 79.200 64.180 ;
        RECT 80.330 64.135 80.620 64.180 ;
        RECT 45.790 63.980 46.080 64.025 ;
        RECT 48.130 63.980 48.420 64.025 ;
        RECT 45.790 63.840 48.420 63.980 ;
        RECT 45.790 63.795 46.080 63.840 ;
        RECT 48.130 63.795 48.420 63.840 ;
        RECT 51.290 63.780 51.610 64.040 ;
        RECT 51.770 63.980 52.060 64.025 ;
        RECT 54.110 63.980 54.400 64.025 ;
        RECT 51.770 63.840 54.400 63.980 ;
        RECT 51.770 63.795 52.060 63.840 ;
        RECT 54.110 63.795 54.400 63.840 ;
        RECT 65.570 63.980 65.860 64.025 ;
        RECT 67.910 63.980 68.200 64.025 ;
        RECT 71.070 63.980 71.390 64.040 ;
        RECT 65.570 63.840 68.200 63.980 ;
        RECT 65.570 63.795 65.860 63.840 ;
        RECT 67.910 63.795 68.200 63.840 ;
        RECT 68.860 63.840 71.390 63.980 ;
        RECT 43.945 63.455 44.235 63.685 ;
        RECT 45.325 63.455 45.615 63.685 ;
        RECT 46.230 63.640 46.550 63.700 ;
        RECT 46.705 63.640 46.995 63.685 ;
        RECT 46.230 63.500 46.995 63.640 ;
        RECT 43.100 63.300 43.240 63.440 ;
        RECT 37.120 63.160 43.240 63.300 ;
        RECT 45.400 63.300 45.540 63.455 ;
        RECT 46.230 63.440 46.550 63.500 ;
        RECT 46.705 63.455 46.995 63.500 ;
        RECT 50.845 63.455 51.135 63.685 ;
        RECT 47.150 63.300 47.470 63.360 ;
        RECT 45.400 63.160 47.470 63.300 ;
        RECT 50.920 63.300 51.060 63.455 ;
        RECT 52.670 63.440 52.990 63.700 ;
        RECT 56.825 63.640 57.115 63.685 ;
        RECT 57.270 63.640 57.590 63.700 ;
        RECT 56.825 63.500 57.590 63.640 ;
        RECT 56.825 63.455 57.115 63.500 ;
        RECT 57.270 63.440 57.590 63.500 ;
        RECT 65.090 63.440 65.410 63.700 ;
        RECT 66.485 63.640 66.775 63.685 ;
        RECT 68.860 63.640 69.000 63.840 ;
        RECT 71.070 63.780 71.390 63.840 ;
        RECT 78.450 63.980 78.740 64.025 ;
        RECT 80.790 63.980 81.080 64.025 ;
        RECT 78.450 63.840 81.080 63.980 ;
        RECT 81.970 63.980 82.110 64.520 ;
        RECT 114.310 64.520 131.650 64.660 ;
        RECT 114.310 64.460 114.630 64.520 ;
        RECT 96.850 64.320 97.140 64.365 ;
        RECT 98.270 64.320 98.560 64.365 ;
        RECT 96.850 64.180 98.560 64.320 ;
        RECT 96.850 64.135 97.140 64.180 ;
        RECT 98.270 64.135 98.560 64.180 ;
        RECT 118.470 64.320 118.760 64.365 ;
        RECT 119.890 64.320 120.180 64.365 ;
        RECT 118.470 64.180 120.180 64.320 ;
        RECT 118.470 64.135 118.760 64.180 ;
        RECT 119.890 64.135 120.180 64.180 ;
        RECT 123.050 64.320 123.370 64.380 ;
        RECT 123.050 64.180 124.660 64.320 ;
        RECT 123.050 64.120 123.370 64.180 ;
        RECT 92.230 63.980 92.550 64.040 ;
        RECT 81.970 63.840 92.550 63.980 ;
        RECT 78.450 63.795 78.740 63.840 ;
        RECT 80.790 63.795 81.080 63.840 ;
        RECT 66.485 63.500 69.000 63.640 ;
        RECT 70.150 63.640 70.470 63.700 ;
        RECT 70.625 63.640 70.915 63.685 ;
        RECT 70.150 63.500 70.915 63.640 ;
        RECT 66.485 63.455 66.775 63.500 ;
        RECT 70.150 63.440 70.470 63.500 ;
        RECT 70.625 63.455 70.915 63.500 ;
        RECT 74.290 63.440 74.610 63.700 ;
        RECT 75.210 63.440 75.530 63.700 ;
        RECT 77.525 63.640 77.815 63.685 ;
        RECT 77.985 63.640 78.275 63.685 ;
        RECT 77.525 63.500 78.275 63.640 ;
        RECT 77.525 63.455 77.815 63.500 ;
        RECT 77.985 63.455 78.275 63.500 ;
        RECT 79.350 63.440 79.670 63.700 ;
        RECT 83.490 63.440 83.810 63.700 ;
        RECT 83.965 63.640 84.255 63.685 ;
        RECT 84.410 63.640 84.730 63.700 ;
        RECT 86.340 63.685 86.480 63.840 ;
        RECT 92.230 63.780 92.550 63.840 ;
        RECT 95.910 63.780 96.230 64.040 ;
        RECT 96.390 63.980 96.680 64.025 ;
        RECT 98.730 63.980 99.020 64.025 ;
        RECT 96.390 63.840 99.020 63.980 ;
        RECT 96.390 63.795 96.680 63.840 ;
        RECT 98.730 63.795 99.020 63.840 ;
        RECT 118.010 63.980 118.300 64.025 ;
        RECT 120.350 63.980 120.640 64.025 ;
        RECT 118.010 63.840 120.640 63.980 ;
        RECT 118.010 63.795 118.300 63.840 ;
        RECT 120.350 63.795 120.640 63.840 ;
        RECT 83.965 63.500 84.730 63.640 ;
        RECT 83.965 63.455 84.255 63.500 ;
        RECT 84.410 63.440 84.730 63.500 ;
        RECT 84.885 63.640 85.175 63.685 ;
        RECT 85.345 63.640 85.635 63.685 ;
        RECT 84.885 63.500 85.635 63.640 ;
        RECT 84.885 63.455 85.175 63.500 ;
        RECT 85.345 63.455 85.635 63.500 ;
        RECT 86.265 63.455 86.555 63.685 ;
        RECT 53.130 63.300 53.450 63.360 ;
        RECT 50.920 63.160 53.450 63.300 ;
        RECT 34.285 63.115 34.575 63.160 ;
        RECT 47.150 63.100 47.470 63.160 ;
        RECT 53.130 63.100 53.450 63.160 ;
        RECT 78.890 63.300 79.210 63.360 ;
        RECT 84.960 63.300 85.100 63.455 ;
        RECT 87.630 63.440 87.950 63.700 ;
        RECT 90.405 63.640 90.695 63.685 ;
        RECT 90.850 63.640 91.170 63.700 ;
        RECT 90.405 63.500 91.170 63.640 ;
        RECT 90.405 63.455 90.695 63.500 ;
        RECT 90.850 63.440 91.170 63.500 ;
        RECT 92.690 63.440 93.010 63.700 ;
        RECT 97.290 63.440 97.610 63.700 ;
        RECT 100.510 63.640 100.830 63.700 ;
        RECT 101.445 63.640 101.735 63.685 ;
        RECT 100.510 63.500 101.735 63.640 ;
        RECT 100.510 63.440 100.830 63.500 ;
        RECT 101.445 63.455 101.735 63.500 ;
        RECT 101.890 63.440 102.210 63.700 ;
        RECT 104.205 63.640 104.495 63.685 ;
        RECT 106.490 63.640 106.810 63.700 ;
        RECT 104.205 63.500 106.810 63.640 ;
        RECT 104.205 63.455 104.495 63.500 ;
        RECT 106.490 63.440 106.810 63.500 ;
        RECT 106.965 63.640 107.255 63.685 ;
        RECT 107.870 63.640 108.190 63.700 ;
        RECT 106.965 63.500 108.190 63.640 ;
        RECT 106.965 63.455 107.255 63.500 ;
        RECT 107.870 63.440 108.190 63.500 ;
        RECT 109.250 63.440 109.570 63.700 ;
        RECT 113.390 63.440 113.710 63.700 ;
        RECT 115.705 63.640 115.995 63.685 ;
        RECT 116.150 63.640 116.470 63.700 ;
        RECT 115.705 63.500 116.470 63.640 ;
        RECT 115.705 63.455 115.995 63.500 ;
        RECT 116.150 63.440 116.470 63.500 ;
        RECT 117.085 63.640 117.375 63.685 ;
        RECT 117.545 63.640 117.835 63.685 ;
        RECT 117.085 63.500 117.835 63.640 ;
        RECT 117.085 63.455 117.375 63.500 ;
        RECT 117.545 63.455 117.835 63.500 ;
        RECT 118.910 63.440 119.230 63.700 ;
        RECT 122.130 63.640 122.450 63.700 ;
        RECT 124.520 63.685 124.660 64.180 ;
        RECT 123.065 63.640 123.355 63.685 ;
        RECT 122.130 63.500 123.355 63.640 ;
        RECT 122.130 63.440 122.450 63.500 ;
        RECT 123.065 63.455 123.355 63.500 ;
        RECT 124.445 63.455 124.735 63.685 ;
        RECT 124.980 63.640 125.120 64.520 ;
        RECT 131.330 64.460 131.650 64.520 ;
        RECT 126.750 64.320 127.040 64.365 ;
        RECT 128.170 64.320 128.460 64.365 ;
        RECT 126.750 64.180 128.460 64.320 ;
        RECT 126.750 64.135 127.040 64.180 ;
        RECT 128.170 64.135 128.460 64.180 ;
        RECT 131.790 64.320 132.110 64.380 ;
        RECT 133.185 64.320 133.475 64.365 ;
        RECT 131.790 64.180 133.475 64.320 ;
        RECT 131.790 64.120 132.110 64.180 ;
        RECT 133.185 64.135 133.475 64.180 ;
        RECT 140.550 64.320 140.840 64.365 ;
        RECT 141.970 64.320 142.260 64.365 ;
        RECT 140.550 64.180 142.260 64.320 ;
        RECT 140.550 64.135 140.840 64.180 ;
        RECT 141.970 64.135 142.260 64.180 ;
        RECT 126.290 63.980 126.580 64.025 ;
        RECT 128.630 63.980 128.920 64.025 ;
        RECT 126.290 63.840 128.920 63.980 ;
        RECT 126.290 63.795 126.580 63.840 ;
        RECT 128.630 63.795 128.920 63.840 ;
        RECT 137.770 63.980 138.090 64.040 ;
        RECT 139.625 63.980 139.915 64.025 ;
        RECT 137.770 63.840 139.915 63.980 ;
        RECT 137.770 63.780 138.090 63.840 ;
        RECT 139.625 63.795 139.915 63.840 ;
        RECT 140.090 63.980 140.380 64.025 ;
        RECT 142.430 63.980 142.720 64.025 ;
        RECT 140.090 63.840 142.720 63.980 ;
        RECT 140.090 63.795 140.380 63.840 ;
        RECT 142.430 63.795 142.720 63.840 ;
        RECT 144.210 63.980 144.530 64.040 ;
        RECT 145.605 63.980 145.895 64.025 ;
        RECT 144.210 63.840 145.895 63.980 ;
        RECT 144.210 63.780 144.530 63.840 ;
        RECT 145.605 63.795 145.895 63.840 ;
        RECT 125.365 63.640 125.655 63.685 ;
        RECT 124.980 63.500 125.655 63.640 ;
        RECT 125.365 63.455 125.655 63.500 ;
        RECT 125.825 63.640 126.115 63.685 ;
        RECT 126.730 63.640 127.050 63.700 ;
        RECT 125.825 63.500 127.050 63.640 ;
        RECT 125.825 63.455 126.115 63.500 ;
        RECT 126.730 63.440 127.050 63.500 ;
        RECT 127.205 63.455 127.495 63.685 ;
        RECT 130.870 63.640 131.190 63.700 ;
        RECT 131.345 63.640 131.635 63.685 ;
        RECT 130.870 63.500 131.635 63.640 ;
        RECT 78.890 63.160 85.100 63.300 ;
        RECT 124.905 63.300 125.195 63.345 ;
        RECT 127.280 63.300 127.420 63.455 ;
        RECT 130.870 63.440 131.190 63.500 ;
        RECT 131.345 63.455 131.635 63.500 ;
        RECT 131.805 63.640 132.095 63.685 ;
        RECT 132.250 63.640 132.570 63.700 ;
        RECT 131.805 63.500 132.570 63.640 ;
        RECT 131.805 63.455 132.095 63.500 ;
        RECT 132.250 63.440 132.570 63.500 ;
        RECT 135.485 63.640 135.775 63.685 ;
        RECT 136.850 63.640 137.170 63.700 ;
        RECT 135.485 63.500 137.170 63.640 ;
        RECT 135.485 63.455 135.775 63.500 ;
        RECT 136.850 63.440 137.170 63.500 ;
        RECT 138.245 63.640 138.535 63.685 ;
        RECT 138.690 63.640 139.010 63.700 ;
        RECT 138.245 63.500 139.010 63.640 ;
        RECT 138.245 63.455 138.535 63.500 ;
        RECT 138.690 63.440 139.010 63.500 ;
        RECT 141.005 63.640 141.295 63.685 ;
        RECT 141.450 63.640 141.770 63.700 ;
        RECT 141.005 63.500 141.770 63.640 ;
        RECT 141.005 63.455 141.295 63.500 ;
        RECT 141.450 63.440 141.770 63.500 ;
        RECT 144.670 63.640 144.990 63.700 ;
        RECT 145.145 63.640 145.435 63.685 ;
        RECT 144.670 63.500 145.435 63.640 ;
        RECT 144.670 63.440 144.990 63.500 ;
        RECT 145.145 63.455 145.435 63.500 ;
        RECT 146.050 63.640 146.370 63.700 ;
        RECT 146.985 63.640 147.275 63.685 ;
        RECT 146.050 63.500 147.275 63.640 ;
        RECT 146.050 63.440 146.370 63.500 ;
        RECT 146.985 63.455 147.275 63.500 ;
        RECT 124.905 63.160 127.420 63.300 ;
        RECT 78.890 63.100 79.210 63.160 ;
        RECT 124.905 63.115 125.195 63.160 ;
        RECT 34.730 62.960 35.050 63.020 ;
        RECT 36.585 62.960 36.875 63.005 ;
        RECT 34.730 62.820 36.875 62.960 ;
        RECT 34.730 62.760 35.050 62.820 ;
        RECT 36.585 62.775 36.875 62.820 ;
        RECT 37.950 62.760 38.270 63.020 ;
        RECT 42.105 62.960 42.395 63.005 ;
        RECT 42.550 62.960 42.870 63.020 ;
        RECT 42.105 62.820 42.870 62.960 ;
        RECT 42.105 62.775 42.395 62.820 ;
        RECT 42.550 62.760 42.870 62.820 ;
        RECT 43.485 62.960 43.775 63.005 ;
        RECT 43.930 62.960 44.250 63.020 ;
        RECT 43.485 62.820 44.250 62.960 ;
        RECT 43.485 62.775 43.775 62.820 ;
        RECT 43.930 62.760 44.250 62.820 ;
        RECT 84.425 62.960 84.715 63.005 ;
        RECT 84.870 62.960 85.190 63.020 ;
        RECT 84.425 62.820 85.190 62.960 ;
        RECT 84.425 62.775 84.715 62.820 ;
        RECT 84.870 62.760 85.190 62.820 ;
        RECT 85.790 62.760 86.110 63.020 ;
        RECT 22.700 62.140 157.820 62.620 ;
        RECT 61.870 61.940 62.190 62.000 ;
        RECT 75.670 61.940 75.990 62.000 ;
        RECT 58.280 61.800 62.190 61.940 ;
        RECT 31.510 61.600 31.830 61.660 ;
        RECT 37.490 61.600 37.810 61.660 ;
        RECT 30.220 61.460 31.830 61.600 ;
        RECT 25.990 61.060 26.310 61.320 ;
        RECT 30.220 61.305 30.360 61.460 ;
        RECT 31.510 61.400 31.830 61.460 ;
        RECT 33.670 61.460 37.810 61.600 ;
        RECT 30.145 61.075 30.435 61.305 ;
        RECT 30.605 61.260 30.895 61.305 ;
        RECT 33.670 61.260 33.810 61.460 ;
        RECT 37.490 61.400 37.810 61.460 ;
        RECT 30.605 61.120 33.810 61.260 ;
        RECT 30.605 61.075 30.895 61.120 ;
        RECT 34.730 61.060 35.050 61.320 ;
        RECT 37.950 61.060 38.270 61.320 ;
        RECT 42.090 61.060 42.410 61.320 ;
        RECT 43.930 61.060 44.250 61.320 ;
        RECT 48.070 61.060 48.390 61.320 ;
        RECT 54.510 61.260 54.830 61.320 ;
        RECT 53.680 61.120 54.830 61.260 ;
        RECT 24.625 60.735 24.915 60.965 ;
        RECT 25.090 60.920 25.380 60.965 ;
        RECT 27.430 60.920 27.720 60.965 ;
        RECT 25.090 60.780 27.720 60.920 ;
        RECT 25.090 60.735 25.380 60.780 ;
        RECT 27.430 60.735 27.720 60.780 ;
        RECT 33.320 60.920 33.610 60.965 ;
        RECT 35.660 60.920 35.950 60.965 ;
        RECT 33.320 60.780 35.950 60.920 ;
        RECT 33.320 60.735 33.610 60.780 ;
        RECT 35.660 60.735 35.950 60.780 ;
        RECT 24.700 60.240 24.840 60.735 ;
        RECT 36.110 60.720 36.430 60.980 ;
        RECT 36.570 60.720 36.890 60.980 ;
        RECT 37.050 60.920 37.340 60.965 ;
        RECT 39.390 60.920 39.680 60.965 ;
        RECT 37.050 60.780 39.680 60.920 ;
        RECT 37.050 60.735 37.340 60.780 ;
        RECT 39.390 60.735 39.680 60.780 ;
        RECT 42.565 60.735 42.855 60.965 ;
        RECT 43.030 60.920 43.320 60.965 ;
        RECT 45.370 60.920 45.660 60.965 ;
        RECT 43.030 60.780 45.660 60.920 ;
        RECT 43.030 60.735 43.320 60.780 ;
        RECT 45.370 60.735 45.660 60.780 ;
        RECT 47.150 60.920 47.470 60.980 ;
        RECT 53.680 60.965 53.820 61.120 ;
        RECT 54.510 61.060 54.830 61.120 ;
        RECT 54.970 61.060 55.290 61.320 ;
        RECT 58.280 61.260 58.420 61.800 ;
        RECT 61.870 61.740 62.190 61.800 ;
        RECT 73.920 61.800 75.990 61.940 ;
        RECT 59.125 61.260 59.415 61.305 ;
        RECT 58.280 61.120 59.415 61.260 ;
        RECT 59.125 61.075 59.415 61.120 ;
        RECT 60.950 61.060 61.270 61.320 ;
        RECT 64.630 61.260 64.950 61.320 ;
        RECT 65.105 61.260 65.395 61.305 ;
        RECT 64.630 61.120 65.395 61.260 ;
        RECT 64.630 61.060 64.950 61.120 ;
        RECT 65.105 61.075 65.395 61.120 ;
        RECT 69.690 61.060 70.010 61.320 ;
        RECT 73.920 61.305 74.060 61.800 ;
        RECT 75.670 61.740 75.990 61.800 ;
        RECT 108.790 61.940 109.110 62.000 ;
        RECT 108.790 61.800 112.240 61.940 ;
        RECT 108.790 61.740 109.110 61.800 ;
        RECT 75.210 61.400 75.530 61.660 ;
        RECT 105.110 61.600 105.430 61.660 ;
        RECT 105.110 61.460 108.100 61.600 ;
        RECT 105.110 61.400 105.430 61.460 ;
        RECT 73.845 61.075 74.135 61.305 ;
        RECT 75.300 61.260 75.440 61.400 ;
        RECT 74.840 61.120 75.440 61.260 ;
        RECT 76.145 61.260 76.435 61.305 ;
        RECT 76.590 61.260 76.910 61.320 ;
        RECT 76.145 61.120 76.910 61.260 ;
        RECT 50.385 60.920 50.675 60.965 ;
        RECT 47.150 60.780 50.675 60.920 ;
        RECT 25.550 60.580 25.840 60.625 ;
        RECT 26.970 60.580 27.260 60.625 ;
        RECT 25.550 60.440 27.260 60.580 ;
        RECT 25.550 60.395 25.840 60.440 ;
        RECT 26.970 60.395 27.260 60.440 ;
        RECT 33.780 60.580 34.070 60.625 ;
        RECT 35.200 60.580 35.490 60.625 ;
        RECT 33.780 60.440 35.490 60.580 ;
        RECT 33.780 60.395 34.070 60.440 ;
        RECT 35.200 60.395 35.490 60.440 ;
        RECT 37.510 60.580 37.800 60.625 ;
        RECT 38.930 60.580 39.220 60.625 ;
        RECT 37.510 60.440 39.220 60.580 ;
        RECT 37.510 60.395 37.800 60.440 ;
        RECT 38.930 60.395 39.220 60.440 ;
        RECT 26.450 60.240 26.770 60.300 ;
        RECT 24.700 60.100 26.770 60.240 ;
        RECT 42.640 60.240 42.780 60.735 ;
        RECT 47.150 60.720 47.470 60.780 ;
        RECT 50.385 60.735 50.675 60.780 ;
        RECT 53.605 60.735 53.895 60.965 ;
        RECT 54.070 60.920 54.360 60.965 ;
        RECT 56.410 60.920 56.700 60.965 ;
        RECT 54.070 60.780 56.700 60.920 ;
        RECT 54.070 60.735 54.360 60.780 ;
        RECT 56.410 60.735 56.700 60.780 ;
        RECT 59.570 60.720 59.890 60.980 ;
        RECT 74.840 60.965 74.980 61.120 ;
        RECT 76.145 61.075 76.435 61.120 ;
        RECT 76.590 61.060 76.910 61.120 ;
        RECT 80.270 61.060 80.590 61.320 ;
        RECT 84.870 61.060 85.190 61.320 ;
        RECT 86.265 61.260 86.555 61.305 ;
        RECT 87.630 61.260 87.950 61.320 ;
        RECT 86.265 61.120 87.950 61.260 ;
        RECT 86.265 61.075 86.555 61.120 ;
        RECT 87.630 61.060 87.950 61.120 ;
        RECT 88.105 61.260 88.395 61.305 ;
        RECT 88.550 61.260 88.870 61.320 ;
        RECT 88.105 61.120 88.870 61.260 ;
        RECT 88.105 61.075 88.395 61.120 ;
        RECT 88.550 61.060 88.870 61.120 ;
        RECT 92.230 61.060 92.550 61.320 ;
        RECT 92.690 61.060 93.010 61.320 ;
        RECT 94.070 61.060 94.390 61.320 ;
        RECT 97.750 61.260 98.070 61.320 ;
        RECT 98.225 61.260 98.515 61.305 ;
        RECT 97.750 61.120 98.515 61.260 ;
        RECT 97.750 61.060 98.070 61.120 ;
        RECT 98.225 61.075 98.515 61.120 ;
        RECT 101.430 61.260 101.750 61.320 ;
        RECT 101.905 61.260 102.195 61.305 ;
        RECT 101.430 61.120 102.195 61.260 ;
        RECT 101.430 61.060 101.750 61.120 ;
        RECT 101.905 61.075 102.195 61.120 ;
        RECT 103.730 61.260 104.050 61.320 ;
        RECT 106.045 61.260 106.335 61.305 ;
        RECT 103.730 61.120 106.335 61.260 ;
        RECT 103.730 61.060 104.050 61.120 ;
        RECT 106.045 61.075 106.335 61.120 ;
        RECT 106.490 61.060 106.810 61.320 ;
        RECT 107.960 61.305 108.100 61.460 ;
        RECT 109.250 61.400 109.570 61.660 ;
        RECT 107.885 61.075 108.175 61.305 ;
        RECT 109.340 61.260 109.480 61.400 ;
        RECT 112.100 61.305 112.240 61.800 ;
        RECT 112.470 61.400 112.790 61.660 ;
        RECT 115.230 61.600 115.550 61.660 ;
        RECT 131.330 61.600 131.650 61.660 ;
        RECT 134.550 61.600 134.870 61.660 ;
        RECT 115.230 61.460 120.060 61.600 ;
        RECT 115.230 61.400 115.550 61.460 ;
        RECT 109.340 61.120 109.940 61.260 ;
        RECT 60.050 60.920 60.340 60.965 ;
        RECT 62.390 60.920 62.680 60.965 ;
        RECT 60.050 60.780 62.680 60.920 ;
        RECT 60.050 60.735 60.340 60.780 ;
        RECT 62.390 60.735 62.680 60.780 ;
        RECT 67.865 60.920 68.155 60.965 ;
        RECT 68.325 60.920 68.615 60.965 ;
        RECT 67.865 60.780 68.615 60.920 ;
        RECT 67.865 60.735 68.155 60.780 ;
        RECT 68.325 60.735 68.615 60.780 ;
        RECT 68.790 60.920 69.080 60.965 ;
        RECT 71.130 60.920 71.420 60.965 ;
        RECT 68.790 60.780 71.420 60.920 ;
        RECT 68.790 60.735 69.080 60.780 ;
        RECT 71.130 60.735 71.420 60.780 ;
        RECT 74.765 60.735 75.055 60.965 ;
        RECT 75.230 60.920 75.520 60.965 ;
        RECT 77.570 60.920 77.860 60.965 ;
        RECT 75.230 60.780 77.860 60.920 ;
        RECT 75.230 60.735 75.520 60.780 ;
        RECT 77.570 60.735 77.860 60.780 ;
        RECT 83.460 60.920 83.750 60.965 ;
        RECT 85.800 60.920 86.090 60.965 ;
        RECT 83.460 60.780 86.090 60.920 ;
        RECT 83.460 60.735 83.750 60.780 ;
        RECT 85.800 60.735 86.090 60.780 ;
        RECT 86.710 60.720 87.030 60.980 ;
        RECT 87.190 60.920 87.480 60.965 ;
        RECT 89.530 60.920 89.820 60.965 ;
        RECT 87.190 60.780 89.820 60.920 ;
        RECT 87.190 60.735 87.480 60.780 ;
        RECT 89.530 60.735 89.820 60.780 ;
        RECT 93.170 60.920 93.460 60.965 ;
        RECT 95.510 60.920 95.800 60.965 ;
        RECT 93.170 60.780 95.800 60.920 ;
        RECT 93.170 60.735 93.460 60.780 ;
        RECT 95.510 60.735 95.800 60.780 ;
        RECT 99.605 60.920 99.895 60.965 ;
        RECT 100.525 60.920 100.815 60.965 ;
        RECT 99.605 60.780 100.815 60.920 ;
        RECT 99.605 60.735 99.895 60.780 ;
        RECT 100.525 60.735 100.815 60.780 ;
        RECT 100.990 60.920 101.280 60.965 ;
        RECT 103.330 60.920 103.620 60.965 ;
        RECT 100.990 60.780 103.620 60.920 ;
        RECT 100.990 60.735 101.280 60.780 ;
        RECT 103.330 60.735 103.620 60.780 ;
        RECT 106.970 60.920 107.260 60.965 ;
        RECT 109.310 60.920 109.600 60.965 ;
        RECT 106.970 60.780 109.600 60.920 ;
        RECT 109.800 60.920 109.940 61.120 ;
        RECT 112.025 61.075 112.315 61.305 ;
        RECT 112.560 61.260 112.700 61.400 ;
        RECT 113.865 61.260 114.155 61.305 ;
        RECT 112.560 61.120 114.155 61.260 ;
        RECT 113.865 61.075 114.155 61.120 ;
        RECT 114.310 61.260 114.630 61.320 ;
        RECT 119.920 61.305 120.060 61.460 ;
        RECT 131.330 61.460 133.860 61.600 ;
        RECT 131.330 61.400 131.650 61.460 ;
        RECT 118.005 61.260 118.295 61.305 ;
        RECT 114.310 61.120 118.295 61.260 ;
        RECT 114.310 61.060 114.630 61.120 ;
        RECT 118.005 61.075 118.295 61.120 ;
        RECT 119.845 61.075 120.135 61.305 ;
        RECT 120.290 61.260 120.610 61.320 ;
        RECT 123.985 61.260 124.275 61.305 ;
        RECT 120.290 61.120 124.275 61.260 ;
        RECT 120.290 61.060 120.610 61.120 ;
        RECT 123.985 61.075 124.275 61.120 ;
        RECT 127.650 61.060 127.970 61.320 ;
        RECT 128.110 61.260 128.430 61.320 ;
        RECT 131.805 61.260 132.095 61.305 ;
        RECT 128.110 61.120 132.095 61.260 ;
        RECT 128.110 61.060 128.430 61.120 ;
        RECT 131.805 61.075 132.095 61.120 ;
        RECT 132.250 61.060 132.570 61.320 ;
        RECT 133.720 61.305 133.860 61.460 ;
        RECT 134.550 61.460 139.840 61.600 ;
        RECT 134.550 61.400 134.870 61.460 ;
        RECT 133.645 61.075 133.935 61.305 ;
        RECT 134.090 61.260 134.410 61.320 ;
        RECT 139.700 61.305 139.840 61.460 ;
        RECT 137.785 61.260 138.075 61.305 ;
        RECT 134.090 61.120 138.075 61.260 ;
        RECT 134.090 61.060 134.410 61.120 ;
        RECT 137.785 61.075 138.075 61.120 ;
        RECT 139.625 61.075 139.915 61.305 ;
        RECT 141.450 61.260 141.770 61.320 ;
        RECT 143.765 61.260 144.055 61.305 ;
        RECT 141.450 61.120 144.055 61.260 ;
        RECT 141.450 61.060 141.770 61.120 ;
        RECT 143.765 61.075 144.055 61.120 ;
        RECT 144.210 61.060 144.530 61.320 ;
        RECT 145.590 61.060 145.910 61.320 ;
        RECT 147.430 61.260 147.750 61.320 ;
        RECT 149.745 61.260 150.035 61.305 ;
        RECT 147.430 61.120 150.035 61.260 ;
        RECT 147.430 61.060 147.750 61.120 ;
        RECT 149.745 61.075 150.035 61.120 ;
        RECT 112.485 60.920 112.775 60.965 ;
        RECT 109.800 60.780 112.775 60.920 ;
        RECT 106.970 60.735 107.260 60.780 ;
        RECT 109.310 60.735 109.600 60.780 ;
        RECT 112.485 60.735 112.775 60.780 ;
        RECT 112.950 60.920 113.240 60.965 ;
        RECT 115.290 60.920 115.580 60.965 ;
        RECT 112.950 60.780 115.580 60.920 ;
        RECT 112.950 60.735 113.240 60.780 ;
        RECT 115.290 60.735 115.580 60.780 ;
        RECT 116.150 60.920 116.470 60.980 ;
        RECT 118.465 60.920 118.755 60.965 ;
        RECT 116.150 60.780 118.755 60.920 ;
        RECT 116.150 60.720 116.470 60.780 ;
        RECT 118.465 60.735 118.755 60.780 ;
        RECT 118.930 60.920 119.220 60.965 ;
        RECT 121.270 60.920 121.560 60.965 ;
        RECT 118.930 60.780 121.560 60.920 ;
        RECT 118.930 60.735 119.220 60.780 ;
        RECT 121.270 60.735 121.560 60.780 ;
        RECT 126.270 60.720 126.590 60.980 ;
        RECT 126.750 60.920 127.040 60.965 ;
        RECT 129.090 60.920 129.380 60.965 ;
        RECT 126.750 60.780 129.380 60.920 ;
        RECT 126.750 60.735 127.040 60.780 ;
        RECT 129.090 60.735 129.380 60.780 ;
        RECT 132.730 60.920 133.020 60.965 ;
        RECT 135.070 60.920 135.360 60.965 ;
        RECT 132.730 60.780 135.360 60.920 ;
        RECT 132.730 60.735 133.020 60.780 ;
        RECT 135.070 60.735 135.360 60.780 ;
        RECT 136.850 60.920 137.170 60.980 ;
        RECT 138.245 60.920 138.535 60.965 ;
        RECT 136.850 60.780 138.535 60.920 ;
        RECT 136.850 60.720 137.170 60.780 ;
        RECT 138.245 60.735 138.535 60.780 ;
        RECT 138.710 60.920 139.000 60.965 ;
        RECT 141.050 60.920 141.340 60.965 ;
        RECT 138.710 60.780 141.340 60.920 ;
        RECT 138.710 60.735 139.000 60.780 ;
        RECT 141.050 60.735 141.340 60.780 ;
        RECT 144.690 60.920 144.980 60.965 ;
        RECT 147.030 60.920 147.320 60.965 ;
        RECT 144.690 60.780 147.320 60.920 ;
        RECT 144.690 60.735 144.980 60.780 ;
        RECT 147.030 60.735 147.320 60.780 ;
        RECT 43.490 60.580 43.780 60.625 ;
        RECT 44.910 60.580 45.200 60.625 ;
        RECT 43.490 60.440 45.200 60.580 ;
        RECT 43.490 60.395 43.780 60.440 ;
        RECT 44.910 60.395 45.200 60.440 ;
        RECT 49.925 60.580 50.215 60.625 ;
        RECT 54.530 60.580 54.820 60.625 ;
        RECT 55.950 60.580 56.240 60.625 ;
        RECT 49.925 60.440 54.280 60.580 ;
        RECT 49.925 60.395 50.215 60.440 ;
        RECT 54.140 60.300 54.280 60.440 ;
        RECT 54.530 60.440 56.240 60.580 ;
        RECT 54.530 60.395 54.820 60.440 ;
        RECT 55.950 60.395 56.240 60.440 ;
        RECT 60.510 60.580 60.800 60.625 ;
        RECT 61.930 60.580 62.220 60.625 ;
        RECT 60.510 60.440 62.220 60.580 ;
        RECT 60.510 60.395 60.800 60.440 ;
        RECT 61.930 60.395 62.220 60.440 ;
        RECT 69.250 60.580 69.540 60.625 ;
        RECT 70.670 60.580 70.960 60.625 ;
        RECT 69.250 60.440 70.960 60.580 ;
        RECT 69.250 60.395 69.540 60.440 ;
        RECT 70.670 60.395 70.960 60.440 ;
        RECT 75.690 60.580 75.980 60.625 ;
        RECT 77.110 60.580 77.400 60.625 ;
        RECT 75.690 60.440 77.400 60.580 ;
        RECT 75.690 60.395 75.980 60.440 ;
        RECT 77.110 60.395 77.400 60.440 ;
        RECT 83.920 60.580 84.210 60.625 ;
        RECT 85.340 60.580 85.630 60.625 ;
        RECT 83.920 60.440 85.630 60.580 ;
        RECT 83.920 60.395 84.210 60.440 ;
        RECT 85.340 60.395 85.630 60.440 ;
        RECT 87.650 60.580 87.940 60.625 ;
        RECT 89.070 60.580 89.360 60.625 ;
        RECT 87.650 60.440 89.360 60.580 ;
        RECT 87.650 60.395 87.940 60.440 ;
        RECT 89.070 60.395 89.360 60.440 ;
        RECT 93.630 60.580 93.920 60.625 ;
        RECT 95.050 60.580 95.340 60.625 ;
        RECT 93.630 60.440 95.340 60.580 ;
        RECT 93.630 60.395 93.920 60.440 ;
        RECT 95.050 60.395 95.340 60.440 ;
        RECT 101.450 60.580 101.740 60.625 ;
        RECT 102.870 60.580 103.160 60.625 ;
        RECT 101.450 60.440 103.160 60.580 ;
        RECT 101.450 60.395 101.740 60.440 ;
        RECT 102.870 60.395 103.160 60.440 ;
        RECT 107.430 60.580 107.720 60.625 ;
        RECT 108.850 60.580 109.140 60.625 ;
        RECT 107.430 60.440 109.140 60.580 ;
        RECT 107.430 60.395 107.720 60.440 ;
        RECT 108.850 60.395 109.140 60.440 ;
        RECT 113.410 60.580 113.700 60.625 ;
        RECT 114.830 60.580 115.120 60.625 ;
        RECT 113.410 60.440 115.120 60.580 ;
        RECT 113.410 60.395 113.700 60.440 ;
        RECT 114.830 60.395 115.120 60.440 ;
        RECT 119.390 60.580 119.680 60.625 ;
        RECT 120.810 60.580 121.100 60.625 ;
        RECT 119.390 60.440 121.100 60.580 ;
        RECT 119.390 60.395 119.680 60.440 ;
        RECT 120.810 60.395 121.100 60.440 ;
        RECT 127.210 60.580 127.500 60.625 ;
        RECT 128.630 60.580 128.920 60.625 ;
        RECT 127.210 60.440 128.920 60.580 ;
        RECT 127.210 60.395 127.500 60.440 ;
        RECT 128.630 60.395 128.920 60.440 ;
        RECT 133.190 60.580 133.480 60.625 ;
        RECT 134.610 60.580 134.900 60.625 ;
        RECT 133.190 60.440 134.900 60.580 ;
        RECT 133.190 60.395 133.480 60.440 ;
        RECT 134.610 60.395 134.900 60.440 ;
        RECT 139.170 60.580 139.460 60.625 ;
        RECT 140.590 60.580 140.880 60.625 ;
        RECT 139.170 60.440 140.880 60.580 ;
        RECT 139.170 60.395 139.460 60.440 ;
        RECT 140.590 60.395 140.880 60.440 ;
        RECT 145.150 60.580 145.440 60.625 ;
        RECT 146.570 60.580 146.860 60.625 ;
        RECT 145.150 60.440 146.860 60.580 ;
        RECT 145.150 60.395 145.440 60.440 ;
        RECT 146.570 60.395 146.860 60.440 ;
        RECT 47.150 60.240 47.470 60.300 ;
        RECT 42.640 60.100 47.470 60.240 ;
        RECT 26.450 60.040 26.770 60.100 ;
        RECT 47.150 60.040 47.470 60.100 ;
        RECT 53.145 60.240 53.435 60.285 ;
        RECT 53.590 60.240 53.910 60.300 ;
        RECT 53.145 60.100 53.910 60.240 ;
        RECT 53.145 60.055 53.435 60.100 ;
        RECT 53.590 60.040 53.910 60.100 ;
        RECT 54.050 60.040 54.370 60.300 ;
        RECT 66.485 60.240 66.775 60.285 ;
        RECT 66.930 60.240 67.250 60.300 ;
        RECT 66.485 60.100 67.250 60.240 ;
        RECT 66.485 60.055 66.775 60.100 ;
        RECT 66.930 60.040 67.250 60.100 ;
        RECT 81.155 60.240 81.445 60.285 ;
        RECT 88.550 60.240 88.870 60.300 ;
        RECT 81.155 60.100 88.870 60.240 ;
        RECT 81.155 60.055 81.445 60.100 ;
        RECT 88.550 60.040 88.870 60.100 ;
        RECT 119.830 60.240 120.150 60.300 ;
        RECT 124.445 60.240 124.735 60.285 ;
        RECT 119.830 60.100 124.735 60.240 ;
        RECT 119.830 60.040 120.150 60.100 ;
        RECT 124.445 60.055 124.735 60.100 ;
        RECT 22.700 59.420 157.020 59.900 ;
        RECT 24.610 59.220 24.930 59.280 ;
        RECT 25.085 59.220 25.375 59.265 ;
        RECT 24.610 59.080 25.375 59.220 ;
        RECT 24.610 59.020 24.930 59.080 ;
        RECT 25.085 59.035 25.375 59.080 ;
        RECT 26.450 59.220 26.770 59.280 ;
        RECT 26.925 59.220 27.215 59.265 ;
        RECT 26.450 59.080 27.215 59.220 ;
        RECT 26.450 59.020 26.770 59.080 ;
        RECT 26.925 59.035 27.215 59.080 ;
        RECT 36.570 59.220 36.890 59.280 ;
        RECT 37.045 59.220 37.335 59.265 ;
        RECT 36.570 59.080 37.335 59.220 ;
        RECT 36.570 59.020 36.890 59.080 ;
        RECT 37.045 59.035 37.335 59.080 ;
        RECT 47.150 59.020 47.470 59.280 ;
        RECT 59.570 59.020 59.890 59.280 ;
        RECT 65.090 59.020 65.410 59.280 ;
        RECT 86.710 59.220 87.030 59.280 ;
        RECT 88.105 59.220 88.395 59.265 ;
        RECT 86.710 59.080 88.395 59.220 ;
        RECT 86.710 59.020 87.030 59.080 ;
        RECT 88.105 59.035 88.395 59.080 ;
        RECT 126.270 59.020 126.590 59.280 ;
        RECT 126.730 59.220 127.050 59.280 ;
        RECT 127.665 59.220 127.955 59.265 ;
        RECT 126.730 59.080 127.955 59.220 ;
        RECT 126.730 59.020 127.050 59.080 ;
        RECT 127.665 59.035 127.955 59.080 ;
        RECT 137.770 59.220 138.090 59.280 ;
        RECT 138.245 59.220 138.535 59.265 ;
        RECT 137.770 59.080 138.535 59.220 ;
        RECT 137.770 59.020 138.090 59.080 ;
        RECT 138.245 59.035 138.535 59.080 ;
        RECT 30.610 58.880 30.900 58.925 ;
        RECT 32.030 58.880 32.320 58.925 ;
        RECT 30.610 58.740 32.320 58.880 ;
        RECT 30.610 58.695 30.900 58.740 ;
        RECT 32.030 58.695 32.320 58.740 ;
        RECT 36.110 58.880 36.430 58.940 ;
        RECT 38.425 58.880 38.715 58.925 ;
        RECT 36.110 58.740 38.715 58.880 ;
        RECT 36.110 58.680 36.430 58.740 ;
        RECT 38.425 58.695 38.715 58.740 ;
        RECT 42.110 58.880 42.400 58.925 ;
        RECT 43.530 58.880 43.820 58.925 ;
        RECT 42.110 58.740 43.820 58.880 ;
        RECT 42.110 58.695 42.400 58.740 ;
        RECT 43.530 58.695 43.820 58.740 ;
        RECT 54.530 58.880 54.820 58.925 ;
        RECT 55.950 58.880 56.240 58.925 ;
        RECT 54.530 58.740 56.240 58.880 ;
        RECT 54.530 58.695 54.820 58.740 ;
        RECT 55.950 58.695 56.240 58.740 ;
        RECT 67.870 58.880 68.160 58.925 ;
        RECT 69.290 58.880 69.580 58.925 ;
        RECT 67.870 58.740 69.580 58.880 ;
        RECT 67.870 58.695 68.160 58.740 ;
        RECT 69.290 58.695 69.580 58.740 ;
        RECT 75.690 58.880 75.980 58.925 ;
        RECT 77.110 58.880 77.400 58.925 ;
        RECT 75.690 58.740 77.400 58.880 ;
        RECT 75.690 58.695 75.980 58.740 ;
        RECT 77.110 58.695 77.400 58.740 ;
        RECT 82.130 58.880 82.420 58.925 ;
        RECT 83.550 58.880 83.840 58.925 ;
        RECT 82.130 58.740 83.840 58.880 ;
        RECT 82.130 58.695 82.420 58.740 ;
        RECT 83.550 58.695 83.840 58.740 ;
        RECT 90.870 58.880 91.160 58.925 ;
        RECT 92.290 58.880 92.580 58.925 ;
        RECT 90.870 58.740 92.580 58.880 ;
        RECT 90.870 58.695 91.160 58.740 ;
        RECT 92.290 58.695 92.580 58.740 ;
        RECT 101.910 58.880 102.200 58.925 ;
        RECT 103.330 58.880 103.620 58.925 ;
        RECT 101.910 58.740 103.620 58.880 ;
        RECT 101.910 58.695 102.200 58.740 ;
        RECT 103.330 58.695 103.620 58.740 ;
        RECT 107.890 58.880 108.180 58.925 ;
        RECT 109.310 58.880 109.600 58.925 ;
        RECT 107.890 58.740 109.600 58.880 ;
        RECT 107.890 58.695 108.180 58.740 ;
        RECT 109.310 58.695 109.600 58.740 ;
        RECT 114.330 58.880 114.620 58.925 ;
        RECT 115.750 58.880 116.040 58.925 ;
        RECT 114.330 58.740 116.040 58.880 ;
        RECT 114.330 58.695 114.620 58.740 ;
        RECT 115.750 58.695 116.040 58.740 ;
        RECT 120.770 58.880 121.060 58.925 ;
        RECT 122.190 58.880 122.480 58.925 ;
        RECT 120.770 58.740 122.480 58.880 ;
        RECT 120.770 58.695 121.060 58.740 ;
        RECT 122.190 58.695 122.480 58.740 ;
        RECT 131.810 58.880 132.100 58.925 ;
        RECT 133.230 58.880 133.520 58.925 ;
        RECT 131.810 58.740 133.520 58.880 ;
        RECT 131.810 58.695 132.100 58.740 ;
        RECT 133.230 58.695 133.520 58.740 ;
        RECT 140.090 58.880 140.380 58.925 ;
        RECT 141.510 58.880 141.800 58.925 ;
        RECT 140.090 58.740 141.800 58.880 ;
        RECT 140.090 58.695 140.380 58.740 ;
        RECT 141.510 58.695 141.800 58.740 ;
        RECT 146.070 58.880 146.360 58.925 ;
        RECT 147.490 58.880 147.780 58.925 ;
        RECT 146.070 58.740 147.780 58.880 ;
        RECT 146.070 58.695 146.360 58.740 ;
        RECT 147.490 58.695 147.780 58.740 ;
        RECT 30.150 58.540 30.440 58.585 ;
        RECT 32.490 58.540 32.780 58.585 ;
        RECT 40.710 58.540 41.030 58.600 ;
        RECT 30.150 58.400 32.780 58.540 ;
        RECT 30.150 58.355 30.440 58.400 ;
        RECT 32.490 58.355 32.780 58.400 ;
        RECT 33.670 58.400 41.030 58.540 ;
        RECT 29.685 58.200 29.975 58.245 ;
        RECT 30.590 58.200 30.910 58.260 ;
        RECT 29.685 58.060 30.910 58.200 ;
        RECT 29.685 58.015 29.975 58.060 ;
        RECT 30.590 58.000 30.910 58.060 ;
        RECT 31.065 58.200 31.355 58.245 ;
        RECT 33.670 58.200 33.810 58.400 ;
        RECT 40.710 58.340 41.030 58.400 ;
        RECT 41.170 58.340 41.490 58.600 ;
        RECT 41.650 58.540 41.940 58.585 ;
        RECT 43.990 58.540 44.280 58.585 ;
        RECT 41.650 58.400 44.280 58.540 ;
        RECT 41.650 58.355 41.940 58.400 ;
        RECT 43.990 58.355 44.280 58.400 ;
        RECT 53.590 58.340 53.910 58.600 ;
        RECT 54.070 58.540 54.360 58.585 ;
        RECT 56.410 58.540 56.700 58.585 ;
        RECT 54.070 58.400 56.700 58.540 ;
        RECT 54.070 58.355 54.360 58.400 ;
        RECT 56.410 58.355 56.700 58.400 ;
        RECT 66.930 58.340 67.250 58.600 ;
        RECT 67.410 58.540 67.700 58.585 ;
        RECT 69.750 58.540 70.040 58.585 ;
        RECT 67.410 58.400 70.040 58.540 ;
        RECT 67.410 58.355 67.700 58.400 ;
        RECT 69.750 58.355 70.040 58.400 ;
        RECT 74.290 58.540 74.610 58.600 ;
        RECT 74.765 58.540 75.055 58.585 ;
        RECT 74.290 58.400 75.055 58.540 ;
        RECT 74.290 58.340 74.610 58.400 ;
        RECT 74.765 58.355 75.055 58.400 ;
        RECT 75.230 58.540 75.520 58.585 ;
        RECT 77.570 58.540 77.860 58.585 ;
        RECT 75.230 58.400 77.860 58.540 ;
        RECT 75.230 58.355 75.520 58.400 ;
        RECT 77.570 58.355 77.860 58.400 ;
        RECT 81.190 58.340 81.510 58.600 ;
        RECT 81.670 58.540 81.960 58.585 ;
        RECT 84.010 58.540 84.300 58.585 ;
        RECT 81.670 58.400 84.300 58.540 ;
        RECT 81.670 58.355 81.960 58.400 ;
        RECT 84.010 58.355 84.300 58.400 ;
        RECT 90.410 58.540 90.700 58.585 ;
        RECT 92.750 58.540 93.040 58.585 ;
        RECT 90.410 58.400 93.040 58.540 ;
        RECT 90.410 58.355 90.700 58.400 ;
        RECT 92.750 58.355 93.040 58.400 ;
        RECT 101.450 58.540 101.740 58.585 ;
        RECT 103.790 58.540 104.080 58.585 ;
        RECT 101.450 58.400 104.080 58.540 ;
        RECT 101.450 58.355 101.740 58.400 ;
        RECT 103.790 58.355 104.080 58.400 ;
        RECT 107.430 58.540 107.720 58.585 ;
        RECT 109.770 58.540 110.060 58.585 ;
        RECT 107.430 58.400 110.060 58.540 ;
        RECT 107.430 58.355 107.720 58.400 ;
        RECT 109.770 58.355 110.060 58.400 ;
        RECT 113.390 58.340 113.710 58.600 ;
        RECT 113.870 58.540 114.160 58.585 ;
        RECT 116.210 58.540 116.500 58.585 ;
        RECT 113.870 58.400 116.500 58.540 ;
        RECT 113.870 58.355 114.160 58.400 ;
        RECT 116.210 58.355 116.500 58.400 ;
        RECT 119.830 58.340 120.150 58.600 ;
        RECT 120.310 58.540 120.600 58.585 ;
        RECT 122.650 58.540 122.940 58.585 ;
        RECT 120.310 58.400 122.940 58.540 ;
        RECT 120.310 58.355 120.600 58.400 ;
        RECT 122.650 58.355 122.940 58.400 ;
        RECT 131.350 58.540 131.640 58.585 ;
        RECT 133.690 58.540 133.980 58.585 ;
        RECT 131.350 58.400 133.980 58.540 ;
        RECT 131.350 58.355 131.640 58.400 ;
        RECT 133.690 58.355 133.980 58.400 ;
        RECT 138.690 58.540 139.010 58.600 ;
        RECT 139.165 58.540 139.455 58.585 ;
        RECT 138.690 58.400 139.455 58.540 ;
        RECT 138.690 58.340 139.010 58.400 ;
        RECT 139.165 58.355 139.455 58.400 ;
        RECT 139.630 58.540 139.920 58.585 ;
        RECT 141.970 58.540 142.260 58.585 ;
        RECT 139.630 58.400 142.260 58.540 ;
        RECT 139.630 58.355 139.920 58.400 ;
        RECT 141.970 58.355 142.260 58.400 ;
        RECT 145.610 58.540 145.900 58.585 ;
        RECT 147.950 58.540 148.240 58.585 ;
        RECT 145.610 58.400 148.240 58.540 ;
        RECT 145.610 58.355 145.900 58.400 ;
        RECT 147.950 58.355 148.240 58.400 ;
        RECT 31.065 58.060 33.810 58.200 ;
        RECT 34.270 58.200 34.590 58.260 ;
        RECT 35.205 58.200 35.495 58.245 ;
        RECT 34.270 58.060 35.495 58.200 ;
        RECT 31.065 58.015 31.355 58.060 ;
        RECT 34.270 58.000 34.590 58.060 ;
        RECT 35.205 58.015 35.495 58.060 ;
        RECT 42.550 58.000 42.870 58.260 ;
        RECT 45.310 58.200 45.630 58.260 ;
        RECT 46.705 58.200 46.995 58.245 ;
        RECT 45.310 58.060 46.995 58.200 ;
        RECT 45.310 58.000 45.630 58.060 ;
        RECT 46.705 58.015 46.995 58.060 ;
        RECT 49.450 58.200 49.770 58.260 ;
        RECT 54.985 58.200 55.275 58.245 ;
        RECT 49.450 58.060 55.275 58.200 ;
        RECT 49.450 58.000 49.770 58.060 ;
        RECT 54.985 58.015 55.275 58.060 ;
        RECT 59.110 58.000 59.430 58.260 ;
        RECT 68.310 58.000 68.630 58.260 ;
        RECT 72.465 58.200 72.755 58.245 ;
        RECT 72.910 58.200 73.230 58.260 ;
        RECT 72.465 58.060 73.230 58.200 ;
        RECT 72.465 58.015 72.755 58.060 ;
        RECT 72.910 58.000 73.230 58.060 ;
        RECT 76.130 58.000 76.450 58.260 ;
        RECT 78.430 58.200 78.750 58.260 ;
        RECT 80.285 58.200 80.575 58.245 ;
        RECT 78.430 58.060 80.575 58.200 ;
        RECT 78.430 58.000 78.750 58.060 ;
        RECT 80.285 58.015 80.575 58.060 ;
        RECT 82.585 58.200 82.875 58.245 ;
        RECT 85.790 58.200 86.110 58.260 ;
        RECT 82.585 58.060 86.110 58.200 ;
        RECT 82.585 58.015 82.875 58.060 ;
        RECT 85.790 58.000 86.110 58.060 ;
        RECT 86.710 58.000 87.030 58.260 ;
        RECT 89.945 58.200 90.235 58.245 ;
        RECT 90.850 58.200 91.170 58.260 ;
        RECT 89.945 58.060 91.170 58.200 ;
        RECT 89.945 58.015 90.235 58.060 ;
        RECT 90.850 58.000 91.170 58.060 ;
        RECT 91.310 58.000 91.630 58.260 ;
        RECT 94.990 58.200 95.310 58.260 ;
        RECT 95.465 58.200 95.755 58.245 ;
        RECT 94.990 58.060 95.755 58.200 ;
        RECT 94.990 58.000 95.310 58.060 ;
        RECT 95.465 58.015 95.755 58.060 ;
        RECT 100.985 58.200 101.275 58.245 ;
        RECT 101.890 58.200 102.210 58.260 ;
        RECT 100.985 58.060 102.210 58.200 ;
        RECT 100.985 58.015 101.275 58.060 ;
        RECT 101.890 58.000 102.210 58.060 ;
        RECT 102.365 58.200 102.655 58.245 ;
        RECT 102.810 58.200 103.130 58.260 ;
        RECT 102.365 58.060 103.130 58.200 ;
        RECT 102.365 58.015 102.655 58.060 ;
        RECT 102.810 58.000 103.130 58.060 ;
        RECT 106.030 58.200 106.350 58.260 ;
        RECT 106.505 58.200 106.795 58.245 ;
        RECT 106.030 58.060 106.795 58.200 ;
        RECT 106.030 58.000 106.350 58.060 ;
        RECT 106.505 58.015 106.795 58.060 ;
        RECT 106.965 58.200 107.255 58.245 ;
        RECT 107.870 58.200 108.190 58.260 ;
        RECT 106.965 58.060 108.190 58.200 ;
        RECT 106.965 58.015 107.255 58.060 ;
        RECT 107.870 58.000 108.190 58.060 ;
        RECT 108.330 58.000 108.650 58.260 ;
        RECT 111.550 58.200 111.870 58.260 ;
        RECT 112.485 58.200 112.775 58.245 ;
        RECT 111.550 58.060 112.775 58.200 ;
        RECT 111.550 58.000 111.870 58.060 ;
        RECT 112.485 58.015 112.775 58.060 ;
        RECT 114.770 58.000 115.090 58.260 ;
        RECT 117.070 58.200 117.390 58.260 ;
        RECT 118.925 58.200 119.215 58.245 ;
        RECT 117.070 58.060 119.215 58.200 ;
        RECT 117.070 58.000 117.390 58.060 ;
        RECT 118.925 58.015 119.215 58.060 ;
        RECT 121.210 58.000 121.530 58.260 ;
        RECT 125.350 58.000 125.670 58.260 ;
        RECT 130.885 58.200 131.175 58.245 ;
        RECT 131.790 58.200 132.110 58.260 ;
        RECT 130.885 58.060 132.110 58.200 ;
        RECT 130.885 58.015 131.175 58.060 ;
        RECT 131.790 58.000 132.110 58.060 ;
        RECT 132.265 58.200 132.555 58.245 ;
        RECT 132.710 58.200 133.030 58.260 ;
        RECT 132.265 58.060 133.030 58.200 ;
        RECT 132.265 58.015 132.555 58.060 ;
        RECT 132.710 58.000 133.030 58.060 ;
        RECT 136.390 58.000 136.710 58.260 ;
        RECT 138.230 58.200 138.550 58.260 ;
        RECT 140.545 58.200 140.835 58.245 ;
        RECT 138.230 58.060 140.835 58.200 ;
        RECT 138.230 58.000 138.550 58.060 ;
        RECT 140.545 58.015 140.835 58.060 ;
        RECT 142.370 58.200 142.690 58.260 ;
        RECT 144.685 58.200 144.975 58.245 ;
        RECT 142.370 58.060 144.975 58.200 ;
        RECT 142.370 58.000 142.690 58.060 ;
        RECT 144.685 58.015 144.975 58.060 ;
        RECT 145.145 58.200 145.435 58.245 ;
        RECT 146.050 58.200 146.370 58.260 ;
        RECT 145.145 58.060 146.370 58.200 ;
        RECT 145.145 58.015 145.435 58.060 ;
        RECT 146.050 58.000 146.370 58.060 ;
        RECT 146.510 58.000 146.830 58.260 ;
        RECT 150.190 58.200 150.510 58.260 ;
        RECT 150.665 58.200 150.955 58.245 ;
        RECT 150.190 58.060 150.955 58.200 ;
        RECT 150.190 58.000 150.510 58.060 ;
        RECT 150.665 58.015 150.955 58.060 ;
        RECT 22.700 56.700 157.820 57.180 ;
        RECT 122.130 56.500 122.450 56.560 ;
        RECT 123.050 56.500 123.370 56.560 ;
        RECT 122.130 56.360 123.370 56.500 ;
        RECT 122.130 56.300 122.450 56.360 ;
        RECT 123.050 56.300 123.370 56.360 ;
        RECT 114.980 52.000 115.830 52.015 ;
        RECT 120.065 52.000 120.875 52.055 ;
        RECT 122.030 52.000 122.780 52.005 ;
        RECT 124.675 52.000 125.485 52.025 ;
        RECT 132.755 52.000 133.505 52.005 ;
        RECT 136.755 52.000 137.505 52.055 ;
        RECT 138.620 52.000 139.430 52.025 ;
        RECT 142.555 52.000 143.305 52.055 ;
        RECT 75.100 50.600 75.950 50.615 ;
        RECT 80.185 50.600 80.995 50.655 ;
        RECT 82.150 50.600 82.900 50.605 ;
        RECT 84.795 50.600 85.605 50.625 ;
        RECT 92.875 50.600 93.625 50.605 ;
        RECT 96.875 50.600 97.625 50.655 ;
        RECT 98.740 50.600 99.550 50.625 ;
        RECT 102.675 50.600 103.425 50.655 ;
        RECT 33.880 49.760 34.730 49.775 ;
        RECT 38.965 49.760 39.775 49.815 ;
        RECT 40.930 49.760 41.680 49.765 ;
        RECT 43.575 49.760 44.385 49.785 ;
        RECT 51.655 49.760 52.405 49.765 ;
        RECT 55.655 49.760 56.405 49.815 ;
        RECT 57.520 49.760 58.330 49.785 ;
        RECT 61.455 49.760 62.205 49.815 ;
        RECT 30.280 46.660 32.280 49.760 ;
        RECT 33.280 48.865 34.730 49.760 ;
        RECT 35.280 48.920 36.750 49.760 ;
        RECT 33.280 48.760 34.280 48.865 ;
        RECT 35.280 48.760 36.280 48.920 ;
        RECT 37.280 48.760 38.280 49.760 ;
        RECT 38.965 48.945 40.280 49.760 ;
        RECT 40.930 48.955 42.280 49.760 ;
        RECT 39.280 48.760 40.280 48.945 ;
        RECT 41.280 48.760 42.280 48.955 ;
        RECT 43.280 49.035 44.385 49.760 ;
        RECT 45.280 49.685 46.280 49.760 ;
        RECT 47.280 49.685 48.280 49.760 ;
        RECT 49.280 49.735 50.280 49.760 ;
        RECT 43.280 48.760 44.280 49.035 ;
        RECT 45.280 48.935 46.610 49.685 ;
        RECT 47.280 48.935 48.760 49.685 ;
        RECT 49.280 48.985 50.610 49.735 ;
        RECT 45.280 48.760 46.280 48.935 ;
        RECT 47.280 48.760 48.280 48.935 ;
        RECT 49.280 48.760 50.280 48.985 ;
        RECT 51.280 48.955 52.405 49.760 ;
        RECT 53.280 49.735 54.280 49.760 ;
        RECT 53.280 48.985 54.485 49.735 ;
        RECT 55.280 49.005 56.405 49.760 ;
        RECT 57.280 49.035 58.330 49.760 ;
        RECT 59.280 49.715 60.280 49.760 ;
        RECT 51.280 48.760 52.280 48.955 ;
        RECT 53.280 48.760 54.280 48.985 ;
        RECT 55.280 48.760 56.280 49.005 ;
        RECT 57.280 48.760 58.280 49.035 ;
        RECT 59.280 48.905 60.455 49.715 ;
        RECT 59.280 48.760 60.280 48.905 ;
        RECT 61.280 48.760 62.280 49.760 ;
        RECT 33.850 47.100 34.760 47.725 ;
        RECT 33.820 46.870 34.780 47.100 ;
        RECT 63.280 46.760 66.280 49.810 ;
        RECT 71.500 47.500 73.500 50.600 ;
        RECT 74.500 49.705 75.950 50.600 ;
        RECT 76.500 49.760 77.970 50.600 ;
        RECT 74.500 49.600 75.500 49.705 ;
        RECT 76.500 49.600 77.500 49.760 ;
        RECT 78.500 49.600 79.500 50.600 ;
        RECT 80.185 49.785 81.500 50.600 ;
        RECT 82.150 49.795 83.500 50.600 ;
        RECT 80.500 49.600 81.500 49.785 ;
        RECT 82.500 49.600 83.500 49.795 ;
        RECT 84.500 49.875 85.605 50.600 ;
        RECT 86.500 50.525 87.500 50.600 ;
        RECT 88.500 50.525 89.500 50.600 ;
        RECT 90.500 50.575 91.500 50.600 ;
        RECT 84.500 49.600 85.500 49.875 ;
        RECT 86.500 49.775 87.830 50.525 ;
        RECT 88.500 49.775 89.980 50.525 ;
        RECT 90.500 49.825 91.830 50.575 ;
        RECT 86.500 49.600 87.500 49.775 ;
        RECT 88.500 49.600 89.500 49.775 ;
        RECT 90.500 49.600 91.500 49.825 ;
        RECT 92.500 49.795 93.625 50.600 ;
        RECT 94.500 50.575 95.500 50.600 ;
        RECT 94.500 49.825 95.705 50.575 ;
        RECT 96.500 49.845 97.625 50.600 ;
        RECT 98.500 49.875 99.550 50.600 ;
        RECT 100.500 50.555 101.500 50.600 ;
        RECT 92.500 49.600 93.500 49.795 ;
        RECT 94.500 49.600 95.500 49.825 ;
        RECT 96.500 49.600 97.500 49.845 ;
        RECT 98.500 49.600 99.500 49.875 ;
        RECT 100.500 49.745 101.675 50.555 ;
        RECT 100.500 49.600 101.500 49.745 ;
        RECT 102.500 49.600 103.500 50.600 ;
        RECT 75.070 47.940 75.980 48.565 ;
        RECT 75.040 47.710 76.000 47.940 ;
        RECT 104.500 47.600 107.500 50.650 ;
        RECT 111.380 48.900 113.380 52.000 ;
        RECT 114.380 51.105 115.830 52.000 ;
        RECT 116.380 51.160 117.850 52.000 ;
        RECT 114.380 51.000 115.380 51.105 ;
        RECT 116.380 51.000 117.380 51.160 ;
        RECT 118.380 51.000 119.380 52.000 ;
        RECT 120.065 51.185 121.380 52.000 ;
        RECT 122.030 51.195 123.380 52.000 ;
        RECT 120.380 51.000 121.380 51.185 ;
        RECT 122.380 51.000 123.380 51.195 ;
        RECT 124.380 51.275 125.485 52.000 ;
        RECT 126.380 51.925 127.380 52.000 ;
        RECT 128.380 51.925 129.380 52.000 ;
        RECT 130.380 51.975 131.380 52.000 ;
        RECT 124.380 51.000 125.380 51.275 ;
        RECT 126.380 51.175 127.710 51.925 ;
        RECT 128.380 51.175 129.860 51.925 ;
        RECT 130.380 51.225 131.710 51.975 ;
        RECT 126.380 51.000 127.380 51.175 ;
        RECT 128.380 51.000 129.380 51.175 ;
        RECT 130.380 51.000 131.380 51.225 ;
        RECT 132.380 51.195 133.505 52.000 ;
        RECT 134.380 51.975 135.380 52.000 ;
        RECT 134.380 51.225 135.585 51.975 ;
        RECT 136.380 51.245 137.505 52.000 ;
        RECT 138.380 51.275 139.430 52.000 ;
        RECT 140.380 51.955 141.380 52.000 ;
        RECT 132.380 51.000 133.380 51.195 ;
        RECT 134.380 51.000 135.380 51.225 ;
        RECT 136.380 51.000 137.380 51.245 ;
        RECT 138.380 51.000 139.380 51.275 ;
        RECT 140.380 51.145 141.555 51.955 ;
        RECT 140.380 51.000 141.380 51.145 ;
        RECT 142.380 51.000 143.380 52.000 ;
        RECT 114.950 49.340 115.860 49.965 ;
        RECT 114.920 49.110 115.880 49.340 ;
        RECT 144.380 49.000 147.380 52.050 ;
        RECT 30.250 44.660 33.280 46.660 ;
        RECT 33.540 46.650 33.770 46.710 ;
        RECT 33.465 44.360 33.770 46.650 ;
        RECT 31.280 34.760 33.770 44.360 ;
        RECT 31.280 32.360 33.280 34.760 ;
        RECT 33.540 34.710 33.770 34.760 ;
        RECT 34.830 46.650 35.060 46.710 ;
        RECT 36.780 46.650 66.280 46.760 ;
        RECT 34.830 43.760 66.280 46.650 ;
        RECT 71.470 45.500 74.500 47.500 ;
        RECT 74.760 47.490 74.990 47.550 ;
        RECT 74.685 45.200 74.990 47.490 ;
        RECT 34.830 37.700 37.760 43.760 ;
        RECT 40.900 38.100 41.710 38.635 ;
        RECT 40.820 37.870 41.780 38.100 ;
        RECT 40.540 37.700 40.770 37.710 ;
        RECT 34.830 34.770 40.770 37.700 ;
        RECT 34.830 34.710 35.060 34.770 ;
        RECT 33.820 34.320 34.780 34.550 ;
        RECT 33.850 33.675 34.760 34.320 ;
        RECT 35.850 32.600 36.750 33.230 ;
        RECT 35.820 32.370 36.780 32.600 ;
        RECT 31.280 29.660 33.080 32.360 ;
        RECT 35.540 32.150 35.770 32.210 ;
        RECT 33.280 30.030 35.280 32.090 ;
        RECT 35.480 29.660 35.770 32.150 ;
        RECT 31.280 24.260 35.770 29.660 ;
        RECT 31.280 23.260 32.780 24.260 ;
        RECT 33.780 23.800 35.770 24.260 ;
        RECT 33.780 23.260 34.880 23.800 ;
        RECT 35.540 23.730 35.770 23.800 ;
        RECT 36.830 32.150 37.060 32.210 ;
        RECT 37.880 32.150 39.680 34.770 ;
        RECT 40.540 34.710 40.770 34.770 ;
        RECT 41.830 36.260 42.060 37.710 ;
        RECT 42.280 36.410 43.980 38.160 ;
        RECT 44.680 37.680 45.325 37.710 ;
        RECT 44.650 37.650 45.355 37.680 ;
        RECT 44.520 37.420 45.480 37.650 ;
        RECT 44.240 36.260 44.470 37.260 ;
        RECT 44.650 37.035 45.355 37.420 ;
        RECT 45.530 37.210 45.760 37.260 ;
        RECT 46.530 37.210 48.530 43.760 ;
        RECT 44.680 37.005 45.325 37.035 ;
        RECT 41.830 35.210 44.470 36.260 ;
        RECT 41.830 35.030 43.580 35.210 ;
        RECT 44.240 35.140 44.470 35.210 ;
        RECT 41.830 34.760 43.600 35.030 ;
        RECT 44.650 34.980 45.355 35.385 ;
        RECT 45.530 35.210 52.180 37.210 ;
        RECT 45.530 35.140 45.760 35.210 ;
        RECT 41.830 34.710 42.060 34.760 ;
        RECT 40.820 34.320 41.780 34.550 ;
        RECT 40.900 33.735 41.710 34.320 ;
        RECT 36.830 25.660 39.680 32.150 ;
        RECT 42.230 29.010 43.600 34.760 ;
        RECT 44.520 34.750 45.480 34.980 ;
        RECT 44.650 34.740 45.355 34.750 ;
        RECT 47.680 34.390 48.980 35.210 ;
        RECT 47.580 34.160 49.080 34.390 ;
        RECT 47.190 34.010 47.420 34.110 ;
        RECT 49.240 34.010 49.470 34.110 ;
        RECT 45.580 33.890 46.930 34.010 ;
        RECT 44.480 33.860 46.930 33.890 ;
        RECT 44.430 32.760 46.930 33.860 ;
        RECT 47.160 33.980 47.800 34.010 ;
        RECT 48.910 33.980 49.550 34.010 ;
        RECT 47.160 33.340 49.550 33.980 ;
        RECT 47.160 33.310 47.800 33.340 ;
        RECT 48.910 33.310 49.550 33.340 ;
        RECT 47.190 33.150 47.420 33.310 ;
        RECT 49.240 33.150 49.470 33.310 ;
        RECT 47.580 32.870 49.080 33.100 ;
        RECT 44.480 32.730 45.580 32.760 ;
        RECT 47.680 32.560 48.980 32.870 ;
        RECT 49.730 32.760 50.630 34.510 ;
        RECT 51.380 34.390 52.180 35.210 ;
        RECT 51.280 34.160 52.280 34.390 ;
        RECT 50.890 33.965 51.120 34.110 ;
        RECT 52.440 33.965 52.670 34.110 ;
        RECT 50.855 33.250 51.510 33.965 ;
        RECT 52.050 33.250 52.705 33.965 ;
        RECT 50.890 33.150 51.120 33.250 ;
        RECT 52.440 33.150 52.670 33.250 ;
        RECT 51.280 32.870 52.280 33.100 ;
        RECT 51.380 32.560 52.230 32.870 ;
        RECT 47.680 31.785 52.230 32.560 ;
        RECT 47.680 29.010 48.980 31.785 ;
        RECT 51.380 31.440 52.230 31.785 ;
        RECT 51.280 31.210 52.280 31.440 ;
        RECT 50.890 30.585 51.120 31.160 ;
        RECT 51.380 31.060 52.230 31.210 ;
        RECT 52.440 30.865 52.670 31.160 ;
        RECT 50.180 30.490 50.630 30.510 ;
        RECT 49.130 29.330 50.630 30.490 ;
        RECT 50.875 29.835 51.685 30.585 ;
        RECT 52.055 30.055 52.805 30.865 ;
        RECT 50.890 29.700 51.120 29.835 ;
        RECT 52.440 29.700 52.670 30.055 ;
        RECT 42.230 27.160 48.980 29.010 ;
        RECT 49.280 29.310 50.630 29.330 ;
        RECT 51.280 29.560 52.280 29.650 ;
        RECT 51.280 29.410 52.330 29.560 ;
        RECT 63.280 29.420 66.280 43.760 ;
        RECT 54.070 29.410 66.280 29.420 ;
        RECT 49.280 28.410 50.280 29.310 ;
        RECT 51.280 28.510 66.280 29.410 ;
        RECT 54.070 28.420 66.280 28.510 ;
        RECT 49.280 27.960 50.880 28.410 ;
        RECT 51.055 28.285 51.805 28.315 ;
        RECT 49.280 27.310 50.280 27.960 ;
        RECT 51.055 27.750 52.885 28.285 ;
        RECT 50.800 27.520 52.885 27.750 ;
        RECT 51.055 27.505 52.885 27.520 ;
        RECT 63.280 27.360 66.280 28.420 ;
        RECT 50.520 27.160 50.830 27.360 ;
        RECT 42.230 26.360 50.830 27.160 ;
        RECT 36.830 23.860 40.680 25.660 ;
        RECT 36.830 23.800 38.630 23.860 ;
        RECT 36.830 23.730 37.060 23.800 ;
        RECT 35.850 23.570 36.750 23.600 ;
        RECT 35.820 23.340 36.780 23.570 ;
        RECT 31.280 21.360 34.880 23.260 ;
        RECT 35.850 22.760 36.750 23.340 ;
        RECT 37.360 21.600 38.240 22.150 ;
        RECT 37.320 21.370 38.280 21.600 ;
        RECT 31.280 18.760 34.280 21.360 ;
        RECT 37.360 21.330 38.240 21.370 ;
        RECT 37.040 21.130 37.270 21.210 ;
        RECT 34.780 19.030 36.780 21.090 ;
        RECT 36.980 18.760 37.270 21.130 ;
        RECT 31.280 15.760 37.270 18.760 ;
        RECT 31.280 14.760 34.280 15.760 ;
        RECT 35.280 15.300 37.270 15.760 ;
        RECT 37.040 15.210 37.270 15.300 ;
        RECT 38.330 21.130 38.560 21.210 ;
        RECT 38.880 21.130 40.680 23.860 ;
        RECT 38.330 20.140 40.680 21.130 ;
        RECT 42.230 23.840 48.980 26.360 ;
        RECT 51.025 26.200 52.780 26.685 ;
        RECT 52.930 26.360 66.280 27.360 ;
        RECT 50.800 25.970 52.880 26.200 ;
        RECT 51.025 25.950 52.780 25.970 ;
        RECT 50.370 25.700 53.420 25.730 ;
        RECT 50.360 25.660 53.420 25.700 ;
        RECT 50.350 24.510 53.420 25.660 ;
        RECT 50.360 24.460 53.420 24.510 ;
        RECT 51.175 24.200 51.925 24.275 ;
        RECT 50.970 23.970 53.930 24.200 ;
        RECT 42.230 23.810 50.890 23.840 ;
        RECT 42.230 22.810 50.920 23.810 ;
        RECT 51.175 23.465 51.925 23.970 ;
        RECT 63.280 23.810 66.280 26.360 ;
        RECT 42.230 22.800 50.890 22.810 ;
        RECT 42.230 21.560 48.980 22.800 ;
        RECT 51.145 22.650 51.955 23.145 ;
        RECT 53.980 22.810 66.280 23.810 ;
        RECT 54.030 22.800 66.280 22.810 ;
        RECT 50.970 22.420 53.930 22.650 ;
        RECT 51.145 22.395 51.955 22.420 ;
        RECT 50.370 22.120 53.420 22.150 ;
        RECT 50.360 22.080 53.420 22.120 ;
        RECT 42.230 21.110 49.000 21.560 ;
        RECT 43.480 20.230 49.000 21.110 ;
        RECT 50.350 20.930 53.420 22.080 ;
        RECT 50.360 20.880 53.420 20.930 ;
        RECT 51.115 20.620 51.865 20.670 ;
        RECT 54.215 20.620 54.965 20.665 ;
        RECT 50.940 20.390 55.140 20.620 ;
        RECT 38.330 15.880 43.080 20.140 ;
        RECT 38.330 15.360 40.680 15.880 ;
        RECT 38.330 15.300 40.440 15.360 ;
        RECT 38.330 15.210 38.560 15.300 ;
        RECT 37.320 14.820 38.280 15.050 ;
        RECT 31.280 10.560 36.180 14.760 ;
        RECT 37.360 14.200 38.240 14.820 ;
        RECT 39.370 13.100 40.240 13.705 ;
        RECT 36.780 10.830 38.780 12.890 ;
        RECT 39.320 12.870 40.280 13.100 ;
        RECT 39.040 12.630 39.270 12.710 ;
        RECT 38.980 10.560 39.270 12.630 ;
        RECT 31.280 8.560 39.270 10.560 ;
        RECT 31.280 7.160 36.180 8.560 ;
        RECT 36.490 8.550 39.270 8.560 ;
        RECT 39.040 8.470 39.270 8.550 ;
        RECT 40.330 12.630 40.560 12.710 ;
        RECT 41.090 12.630 43.080 15.880 ;
        RECT 40.330 8.550 43.080 12.630 ;
        RECT 43.480 19.230 50.890 20.230 ;
        RECT 51.115 19.860 51.865 20.390 ;
        RECT 54.215 19.855 54.965 20.390 ;
        RECT 55.190 20.220 55.420 20.230 ;
        RECT 63.280 20.220 66.280 22.800 ;
        RECT 43.480 16.660 48.980 19.230 ;
        RECT 51.085 19.070 51.895 19.535 ;
        RECT 54.295 19.070 55.045 19.565 ;
        RECT 55.190 19.290 66.280 20.220 ;
        RECT 55.190 19.230 55.420 19.290 ;
        RECT 50.940 18.840 55.140 19.070 ;
        RECT 51.085 18.785 51.895 18.840 ;
        RECT 54.295 18.755 55.045 18.840 ;
        RECT 50.370 18.540 53.420 18.570 ;
        RECT 50.360 18.500 53.420 18.540 ;
        RECT 50.350 17.350 53.420 18.500 ;
        RECT 50.360 17.300 53.420 17.350 ;
        RECT 50.985 17.040 51.735 17.110 ;
        RECT 55.825 17.040 56.635 17.075 ;
        RECT 50.810 16.810 56.770 17.040 ;
        RECT 43.480 16.650 50.730 16.660 ;
        RECT 43.480 15.660 50.760 16.650 ;
        RECT 50.985 16.300 51.735 16.810 ;
        RECT 55.825 16.325 56.635 16.810 ;
        RECT 56.820 16.640 57.050 16.650 ;
        RECT 63.280 16.640 66.280 19.290 ;
        RECT 43.480 13.060 48.980 15.660 ;
        RECT 50.530 15.650 50.760 15.660 ;
        RECT 50.955 15.490 51.765 15.955 ;
        RECT 55.855 15.490 56.605 15.985 ;
        RECT 56.800 15.710 66.280 16.640 ;
        RECT 56.820 15.650 57.050 15.710 ;
        RECT 50.810 15.260 56.770 15.490 ;
        RECT 50.955 15.205 51.765 15.260 ;
        RECT 55.855 15.175 56.605 15.260 ;
        RECT 50.370 14.960 53.420 14.990 ;
        RECT 50.360 14.920 53.420 14.960 ;
        RECT 50.350 13.770 53.420 14.920 ;
        RECT 50.360 13.720 53.420 13.770 ;
        RECT 50.965 13.460 51.715 13.550 ;
        RECT 58.355 13.460 59.165 13.505 ;
        RECT 50.830 13.230 59.270 13.460 ;
        RECT 50.550 13.060 50.780 13.070 ;
        RECT 43.480 12.070 50.780 13.060 ;
        RECT 50.965 12.740 51.715 13.230 ;
        RECT 58.355 12.755 59.165 13.230 ;
        RECT 59.320 13.060 59.550 13.070 ;
        RECT 63.280 13.060 66.280 15.710 ;
        RECT 43.480 12.060 50.740 12.070 ;
        RECT 43.480 9.500 48.980 12.060 ;
        RECT 50.935 11.910 51.745 12.385 ;
        RECT 58.385 11.910 59.135 12.415 ;
        RECT 59.320 12.130 66.280 13.060 ;
        RECT 59.320 12.070 59.550 12.130 ;
        RECT 50.830 11.680 59.270 11.910 ;
        RECT 50.935 11.635 51.745 11.680 ;
        RECT 58.385 11.605 59.135 11.680 ;
        RECT 50.370 11.380 53.420 11.410 ;
        RECT 50.360 11.340 53.420 11.380 ;
        RECT 50.350 10.190 53.420 11.340 ;
        RECT 63.280 10.760 66.280 12.130 ;
        RECT 72.500 35.600 74.990 45.200 ;
        RECT 72.500 33.200 74.500 35.600 ;
        RECT 74.760 35.550 74.990 35.600 ;
        RECT 76.050 47.490 76.280 47.550 ;
        RECT 78.000 47.490 107.500 47.600 ;
        RECT 76.050 45.950 107.500 47.490 ;
        RECT 111.350 46.900 114.380 48.900 ;
        RECT 114.640 48.890 114.870 48.950 ;
        RECT 114.565 46.600 114.870 48.890 ;
        RECT 76.050 44.600 107.530 45.950 ;
        RECT 76.050 38.540 78.980 44.600 ;
        RECT 82.120 38.940 82.930 39.475 ;
        RECT 82.040 38.710 83.000 38.940 ;
        RECT 81.760 38.540 81.990 38.550 ;
        RECT 76.050 35.610 81.990 38.540 ;
        RECT 76.050 35.550 76.280 35.610 ;
        RECT 75.040 35.160 76.000 35.390 ;
        RECT 75.070 34.515 75.980 35.160 ;
        RECT 77.070 33.440 77.970 34.070 ;
        RECT 77.040 33.210 78.000 33.440 ;
        RECT 72.500 30.500 74.300 33.200 ;
        RECT 76.760 32.990 76.990 33.050 ;
        RECT 74.500 30.870 76.500 32.930 ;
        RECT 76.700 30.500 76.990 32.990 ;
        RECT 72.500 25.100 76.990 30.500 ;
        RECT 72.500 24.100 74.000 25.100 ;
        RECT 75.000 24.640 76.990 25.100 ;
        RECT 75.000 24.100 76.100 24.640 ;
        RECT 76.760 24.570 76.990 24.640 ;
        RECT 78.050 32.990 78.280 33.050 ;
        RECT 79.100 32.990 80.900 35.610 ;
        RECT 81.760 35.550 81.990 35.610 ;
        RECT 83.050 37.100 83.280 38.550 ;
        RECT 83.500 37.250 85.200 39.000 ;
        RECT 85.900 38.520 86.545 38.550 ;
        RECT 85.870 38.490 86.575 38.520 ;
        RECT 85.740 38.260 86.700 38.490 ;
        RECT 85.460 37.100 85.690 38.100 ;
        RECT 85.870 37.875 86.575 38.260 ;
        RECT 86.750 38.050 86.980 38.100 ;
        RECT 87.750 38.050 89.750 44.600 ;
        RECT 85.900 37.845 86.545 37.875 ;
        RECT 83.050 36.050 85.690 37.100 ;
        RECT 83.050 35.870 84.800 36.050 ;
        RECT 85.460 35.980 85.690 36.050 ;
        RECT 83.050 35.600 84.820 35.870 ;
        RECT 85.870 35.820 86.575 36.225 ;
        RECT 86.750 36.050 93.400 38.050 ;
        RECT 86.750 35.980 86.980 36.050 ;
        RECT 83.050 35.550 83.280 35.600 ;
        RECT 82.040 35.160 83.000 35.390 ;
        RECT 82.120 34.575 82.930 35.160 ;
        RECT 78.050 26.500 80.900 32.990 ;
        RECT 83.450 29.850 84.820 35.600 ;
        RECT 85.740 35.590 86.700 35.820 ;
        RECT 85.870 35.580 86.575 35.590 ;
        RECT 88.900 35.230 90.200 36.050 ;
        RECT 88.800 35.000 90.300 35.230 ;
        RECT 88.410 34.850 88.640 34.950 ;
        RECT 90.460 34.850 90.690 34.950 ;
        RECT 86.800 34.730 88.150 34.850 ;
        RECT 85.700 34.700 88.150 34.730 ;
        RECT 85.650 33.600 88.150 34.700 ;
        RECT 88.380 34.820 89.020 34.850 ;
        RECT 90.130 34.820 90.770 34.850 ;
        RECT 88.380 34.180 90.770 34.820 ;
        RECT 88.380 34.150 89.020 34.180 ;
        RECT 90.130 34.150 90.770 34.180 ;
        RECT 88.410 33.990 88.640 34.150 ;
        RECT 90.460 33.990 90.690 34.150 ;
        RECT 88.800 33.710 90.300 33.940 ;
        RECT 85.700 33.570 86.800 33.600 ;
        RECT 88.900 33.400 90.200 33.710 ;
        RECT 90.950 33.600 91.850 35.350 ;
        RECT 92.600 35.230 93.400 36.050 ;
        RECT 92.500 35.000 93.500 35.230 ;
        RECT 92.110 34.805 92.340 34.950 ;
        RECT 93.660 34.805 93.890 34.950 ;
        RECT 92.075 34.090 92.730 34.805 ;
        RECT 93.270 34.090 93.925 34.805 ;
        RECT 92.110 33.990 92.340 34.090 ;
        RECT 93.660 33.990 93.890 34.090 ;
        RECT 92.500 33.710 93.500 33.940 ;
        RECT 92.600 33.400 93.450 33.710 ;
        RECT 88.900 32.625 93.450 33.400 ;
        RECT 88.900 29.850 90.200 32.625 ;
        RECT 92.600 32.280 93.450 32.625 ;
        RECT 92.500 32.050 93.500 32.280 ;
        RECT 92.110 31.425 92.340 32.000 ;
        RECT 92.600 31.900 93.450 32.050 ;
        RECT 93.660 31.705 93.890 32.000 ;
        RECT 91.400 31.330 91.850 31.350 ;
        RECT 90.350 30.170 91.850 31.330 ;
        RECT 92.095 30.675 92.905 31.425 ;
        RECT 93.275 30.895 94.025 31.705 ;
        RECT 92.110 30.540 92.340 30.675 ;
        RECT 93.660 30.540 93.890 30.895 ;
        RECT 83.450 28.000 90.200 29.850 ;
        RECT 90.500 30.150 91.850 30.170 ;
        RECT 92.500 30.400 93.500 30.490 ;
        RECT 92.500 30.250 93.550 30.400 ;
        RECT 104.500 30.260 107.530 44.600 ;
        RECT 95.290 30.250 107.530 30.260 ;
        RECT 90.500 29.250 91.500 30.150 ;
        RECT 92.500 29.350 107.530 30.250 ;
        RECT 95.290 29.260 107.530 29.350 ;
        RECT 90.500 28.800 92.100 29.250 ;
        RECT 92.275 29.125 93.025 29.155 ;
        RECT 90.500 28.150 91.500 28.800 ;
        RECT 92.275 28.590 94.105 29.125 ;
        RECT 92.020 28.360 94.105 28.590 ;
        RECT 92.275 28.345 94.105 28.360 ;
        RECT 104.500 28.200 107.530 29.260 ;
        RECT 91.740 28.000 92.050 28.200 ;
        RECT 83.450 27.200 92.050 28.000 ;
        RECT 78.050 24.700 81.900 26.500 ;
        RECT 78.050 24.640 79.850 24.700 ;
        RECT 78.050 24.570 78.280 24.640 ;
        RECT 77.070 24.410 77.970 24.440 ;
        RECT 77.040 24.180 78.000 24.410 ;
        RECT 72.500 22.200 76.100 24.100 ;
        RECT 77.070 23.600 77.970 24.180 ;
        RECT 78.580 22.440 79.460 22.990 ;
        RECT 78.540 22.210 79.500 22.440 ;
        RECT 72.500 19.600 75.500 22.200 ;
        RECT 78.580 22.170 79.460 22.210 ;
        RECT 78.260 21.970 78.490 22.050 ;
        RECT 76.000 19.870 78.000 21.930 ;
        RECT 78.200 19.600 78.490 21.970 ;
        RECT 72.500 16.600 78.490 19.600 ;
        RECT 72.500 15.600 75.500 16.600 ;
        RECT 76.500 16.140 78.490 16.600 ;
        RECT 78.260 16.050 78.490 16.140 ;
        RECT 79.550 21.970 79.780 22.050 ;
        RECT 80.100 21.970 81.900 24.700 ;
        RECT 79.550 20.980 81.900 21.970 ;
        RECT 83.450 24.680 90.200 27.200 ;
        RECT 92.245 27.040 94.000 27.525 ;
        RECT 94.150 27.200 107.530 28.200 ;
        RECT 92.020 26.810 94.100 27.040 ;
        RECT 92.245 26.790 94.000 26.810 ;
        RECT 91.590 26.540 94.640 26.570 ;
        RECT 91.580 26.500 94.640 26.540 ;
        RECT 91.570 25.350 94.640 26.500 ;
        RECT 91.580 25.300 94.640 25.350 ;
        RECT 92.395 25.040 93.145 25.115 ;
        RECT 92.190 24.810 95.150 25.040 ;
        RECT 83.450 24.650 92.110 24.680 ;
        RECT 83.450 23.650 92.140 24.650 ;
        RECT 92.395 24.305 93.145 24.810 ;
        RECT 104.500 24.650 107.530 27.200 ;
        RECT 83.450 23.640 92.110 23.650 ;
        RECT 83.450 22.400 90.200 23.640 ;
        RECT 92.365 23.490 93.175 23.985 ;
        RECT 95.200 23.650 107.530 24.650 ;
        RECT 95.250 23.640 107.530 23.650 ;
        RECT 92.190 23.260 95.150 23.490 ;
        RECT 92.365 23.235 93.175 23.260 ;
        RECT 91.590 22.960 94.640 22.990 ;
        RECT 91.580 22.920 94.640 22.960 ;
        RECT 83.450 21.950 90.220 22.400 ;
        RECT 84.700 21.070 90.220 21.950 ;
        RECT 91.570 21.770 94.640 22.920 ;
        RECT 91.580 21.720 94.640 21.770 ;
        RECT 92.335 21.460 93.085 21.510 ;
        RECT 95.435 21.460 96.185 21.505 ;
        RECT 92.160 21.230 96.360 21.460 ;
        RECT 79.550 16.720 84.300 20.980 ;
        RECT 79.550 16.200 81.900 16.720 ;
        RECT 79.550 16.140 81.660 16.200 ;
        RECT 79.550 16.050 79.780 16.140 ;
        RECT 78.540 15.660 79.500 15.890 ;
        RECT 72.500 11.400 77.400 15.600 ;
        RECT 78.580 15.040 79.460 15.660 ;
        RECT 80.590 13.940 81.460 14.545 ;
        RECT 78.000 11.670 80.000 13.730 ;
        RECT 80.540 13.710 81.500 13.940 ;
        RECT 80.260 13.470 80.490 13.550 ;
        RECT 80.200 11.400 80.490 13.470 ;
        RECT 50.360 10.140 53.420 10.190 ;
        RECT 50.995 9.880 51.745 9.950 ;
        RECT 61.875 9.880 62.685 9.915 ;
        RECT 50.840 9.650 62.800 9.880 ;
        RECT 43.480 9.490 50.770 9.500 ;
        RECT 40.330 8.470 40.560 8.550 ;
        RECT 43.480 8.500 50.790 9.490 ;
        RECT 50.995 9.140 51.745 9.650 ;
        RECT 61.875 9.165 62.685 9.650 ;
        RECT 62.850 9.480 63.080 9.490 ;
        RECT 64.000 9.480 65.020 10.760 ;
        RECT 39.320 8.080 40.280 8.310 ;
        RECT 39.370 7.495 40.240 8.080 ;
        RECT 43.480 7.240 48.980 8.500 ;
        RECT 50.560 8.490 50.790 8.500 ;
        RECT 50.965 8.330 51.775 8.785 ;
        RECT 61.905 8.330 62.655 8.815 ;
        RECT 62.850 8.500 65.020 9.480 ;
        RECT 72.500 9.400 80.490 11.400 ;
        RECT 62.850 8.490 63.080 8.500 ;
        RECT 50.840 8.100 62.800 8.330 ;
        RECT 50.965 8.035 51.775 8.100 ;
        RECT 61.905 8.005 62.655 8.100 ;
        RECT 72.500 8.000 77.400 9.400 ;
        RECT 77.710 9.390 80.490 9.400 ;
        RECT 80.260 9.310 80.490 9.390 ;
        RECT 81.550 13.470 81.780 13.550 ;
        RECT 82.310 13.470 84.300 16.720 ;
        RECT 81.550 9.390 84.300 13.470 ;
        RECT 84.700 20.070 92.110 21.070 ;
        RECT 92.335 20.700 93.085 21.230 ;
        RECT 95.435 20.695 96.185 21.230 ;
        RECT 96.410 21.060 96.640 21.070 ;
        RECT 104.500 21.060 107.530 23.640 ;
        RECT 84.700 17.500 90.200 20.070 ;
        RECT 92.305 19.910 93.115 20.375 ;
        RECT 95.515 19.910 96.265 20.405 ;
        RECT 96.410 20.130 107.530 21.060 ;
        RECT 96.410 20.070 96.640 20.130 ;
        RECT 92.160 19.680 96.360 19.910 ;
        RECT 92.305 19.625 93.115 19.680 ;
        RECT 95.515 19.595 96.265 19.680 ;
        RECT 91.590 19.380 94.640 19.410 ;
        RECT 91.580 19.340 94.640 19.380 ;
        RECT 91.570 18.190 94.640 19.340 ;
        RECT 91.580 18.140 94.640 18.190 ;
        RECT 92.205 17.880 92.955 17.950 ;
        RECT 97.045 17.880 97.855 17.915 ;
        RECT 92.030 17.650 97.990 17.880 ;
        RECT 84.700 17.490 91.950 17.500 ;
        RECT 84.700 16.500 91.980 17.490 ;
        RECT 92.205 17.140 92.955 17.650 ;
        RECT 97.045 17.165 97.855 17.650 ;
        RECT 98.040 17.480 98.270 17.490 ;
        RECT 104.500 17.480 107.530 20.130 ;
        RECT 84.700 13.900 90.200 16.500 ;
        RECT 91.750 16.490 91.980 16.500 ;
        RECT 92.175 16.330 92.985 16.795 ;
        RECT 97.075 16.330 97.825 16.825 ;
        RECT 98.020 16.550 107.530 17.480 ;
        RECT 98.040 16.490 98.270 16.550 ;
        RECT 92.030 16.100 97.990 16.330 ;
        RECT 92.175 16.045 92.985 16.100 ;
        RECT 97.075 16.015 97.825 16.100 ;
        RECT 91.590 15.800 94.640 15.830 ;
        RECT 91.580 15.760 94.640 15.800 ;
        RECT 91.570 14.610 94.640 15.760 ;
        RECT 91.580 14.560 94.640 14.610 ;
        RECT 92.185 14.300 92.935 14.390 ;
        RECT 99.575 14.300 100.385 14.345 ;
        RECT 92.050 14.070 100.490 14.300 ;
        RECT 91.770 13.900 92.000 13.910 ;
        RECT 84.700 12.910 92.000 13.900 ;
        RECT 92.185 13.580 92.935 14.070 ;
        RECT 99.575 13.595 100.385 14.070 ;
        RECT 100.540 13.900 100.770 13.910 ;
        RECT 104.500 13.900 107.530 16.550 ;
        RECT 84.700 12.900 91.960 12.910 ;
        RECT 84.700 10.340 90.200 12.900 ;
        RECT 92.155 12.750 92.965 13.225 ;
        RECT 99.605 12.750 100.355 13.255 ;
        RECT 100.540 12.970 107.530 13.900 ;
        RECT 100.540 12.910 100.770 12.970 ;
        RECT 92.050 12.520 100.490 12.750 ;
        RECT 92.155 12.475 92.965 12.520 ;
        RECT 99.605 12.445 100.355 12.520 ;
        RECT 91.590 12.220 94.640 12.250 ;
        RECT 91.580 12.180 94.640 12.220 ;
        RECT 91.570 11.030 94.640 12.180 ;
        RECT 104.500 11.600 107.530 12.970 ;
        RECT 91.580 10.980 94.640 11.030 ;
        RECT 105.220 10.850 107.530 11.600 ;
        RECT 112.380 37.000 114.870 46.600 ;
        RECT 112.380 34.600 114.380 37.000 ;
        RECT 114.640 36.950 114.870 37.000 ;
        RECT 115.930 48.890 116.160 48.950 ;
        RECT 117.880 48.890 147.380 49.000 ;
        RECT 115.930 46.000 147.380 48.890 ;
        RECT 115.930 39.940 118.860 46.000 ;
        RECT 122.000 40.340 122.810 40.875 ;
        RECT 121.920 40.110 122.880 40.340 ;
        RECT 121.640 39.940 121.870 39.950 ;
        RECT 115.930 37.010 121.870 39.940 ;
        RECT 115.930 36.950 116.160 37.010 ;
        RECT 114.920 36.560 115.880 36.790 ;
        RECT 114.950 35.915 115.860 36.560 ;
        RECT 116.950 34.840 117.850 35.470 ;
        RECT 116.920 34.610 117.880 34.840 ;
        RECT 112.380 31.900 114.180 34.600 ;
        RECT 116.640 34.390 116.870 34.450 ;
        RECT 114.380 32.270 116.380 34.330 ;
        RECT 116.580 31.900 116.870 34.390 ;
        RECT 112.380 26.500 116.870 31.900 ;
        RECT 112.380 25.500 113.880 26.500 ;
        RECT 114.880 26.040 116.870 26.500 ;
        RECT 114.880 25.500 115.980 26.040 ;
        RECT 116.640 25.970 116.870 26.040 ;
        RECT 117.930 34.390 118.160 34.450 ;
        RECT 118.980 34.390 120.780 37.010 ;
        RECT 121.640 36.950 121.870 37.010 ;
        RECT 122.930 38.500 123.160 39.950 ;
        RECT 123.380 38.650 125.080 40.400 ;
        RECT 125.780 39.920 126.425 39.950 ;
        RECT 125.750 39.890 126.455 39.920 ;
        RECT 125.620 39.660 126.580 39.890 ;
        RECT 125.340 38.500 125.570 39.500 ;
        RECT 125.750 39.275 126.455 39.660 ;
        RECT 126.630 39.450 126.860 39.500 ;
        RECT 127.630 39.450 129.630 46.000 ;
        RECT 144.380 45.850 147.380 46.000 ;
        RECT 125.780 39.245 126.425 39.275 ;
        RECT 122.930 37.450 125.570 38.500 ;
        RECT 122.930 37.270 124.680 37.450 ;
        RECT 125.340 37.380 125.570 37.450 ;
        RECT 122.930 37.000 124.700 37.270 ;
        RECT 125.750 37.220 126.455 37.625 ;
        RECT 126.630 37.450 133.280 39.450 ;
        RECT 126.630 37.380 126.860 37.450 ;
        RECT 122.930 36.950 123.160 37.000 ;
        RECT 121.920 36.560 122.880 36.790 ;
        RECT 122.000 35.975 122.810 36.560 ;
        RECT 117.930 27.900 120.780 34.390 ;
        RECT 123.330 31.250 124.700 37.000 ;
        RECT 125.620 36.990 126.580 37.220 ;
        RECT 125.750 36.980 126.455 36.990 ;
        RECT 128.780 36.630 130.080 37.450 ;
        RECT 128.680 36.400 130.180 36.630 ;
        RECT 128.290 36.250 128.520 36.350 ;
        RECT 130.340 36.250 130.570 36.350 ;
        RECT 126.680 36.130 128.030 36.250 ;
        RECT 125.580 36.100 128.030 36.130 ;
        RECT 125.530 35.000 128.030 36.100 ;
        RECT 128.260 36.220 128.900 36.250 ;
        RECT 130.010 36.220 130.650 36.250 ;
        RECT 128.260 35.580 130.650 36.220 ;
        RECT 128.260 35.550 128.900 35.580 ;
        RECT 130.010 35.550 130.650 35.580 ;
        RECT 128.290 35.390 128.520 35.550 ;
        RECT 130.340 35.390 130.570 35.550 ;
        RECT 128.680 35.110 130.180 35.340 ;
        RECT 125.580 34.970 126.680 35.000 ;
        RECT 128.780 34.800 130.080 35.110 ;
        RECT 130.830 35.000 131.730 36.750 ;
        RECT 132.480 36.630 133.280 37.450 ;
        RECT 132.380 36.400 133.380 36.630 ;
        RECT 131.990 36.205 132.220 36.350 ;
        RECT 133.540 36.205 133.770 36.350 ;
        RECT 131.955 35.490 132.610 36.205 ;
        RECT 133.150 35.490 133.805 36.205 ;
        RECT 131.990 35.390 132.220 35.490 ;
        RECT 133.540 35.390 133.770 35.490 ;
        RECT 132.380 35.110 133.380 35.340 ;
        RECT 132.480 34.800 133.330 35.110 ;
        RECT 128.780 34.025 133.330 34.800 ;
        RECT 128.780 31.250 130.080 34.025 ;
        RECT 132.480 33.680 133.330 34.025 ;
        RECT 132.380 33.450 133.380 33.680 ;
        RECT 131.990 32.825 132.220 33.400 ;
        RECT 132.480 33.300 133.330 33.450 ;
        RECT 133.540 33.105 133.770 33.400 ;
        RECT 131.280 32.730 131.730 32.750 ;
        RECT 130.230 31.570 131.730 32.730 ;
        RECT 131.975 32.075 132.785 32.825 ;
        RECT 133.155 32.295 133.905 33.105 ;
        RECT 131.990 31.940 132.220 32.075 ;
        RECT 133.540 31.940 133.770 32.295 ;
        RECT 123.330 29.400 130.080 31.250 ;
        RECT 130.380 31.550 131.730 31.570 ;
        RECT 132.380 31.800 133.380 31.890 ;
        RECT 132.380 31.650 133.430 31.800 ;
        RECT 144.380 31.660 147.400 45.850 ;
        RECT 135.170 31.650 147.400 31.660 ;
        RECT 130.380 30.650 131.380 31.550 ;
        RECT 132.380 30.750 147.400 31.650 ;
        RECT 135.170 30.660 147.400 30.750 ;
        RECT 130.380 30.200 131.980 30.650 ;
        RECT 132.155 30.525 132.905 30.555 ;
        RECT 130.380 29.550 131.380 30.200 ;
        RECT 132.155 29.990 133.985 30.525 ;
        RECT 131.900 29.760 133.985 29.990 ;
        RECT 132.155 29.745 133.985 29.760 ;
        RECT 144.380 29.600 147.400 30.660 ;
        RECT 131.620 29.400 131.930 29.600 ;
        RECT 123.330 28.600 131.930 29.400 ;
        RECT 117.930 26.100 121.780 27.900 ;
        RECT 117.930 26.040 119.730 26.100 ;
        RECT 117.930 25.970 118.160 26.040 ;
        RECT 116.950 25.810 117.850 25.840 ;
        RECT 116.920 25.580 117.880 25.810 ;
        RECT 112.380 23.600 115.980 25.500 ;
        RECT 116.950 25.000 117.850 25.580 ;
        RECT 118.460 23.840 119.340 24.390 ;
        RECT 118.420 23.610 119.380 23.840 ;
        RECT 112.380 21.000 115.380 23.600 ;
        RECT 118.460 23.570 119.340 23.610 ;
        RECT 118.140 23.370 118.370 23.450 ;
        RECT 115.880 21.270 117.880 23.330 ;
        RECT 118.080 21.000 118.370 23.370 ;
        RECT 112.380 18.000 118.370 21.000 ;
        RECT 112.380 17.000 115.380 18.000 ;
        RECT 116.380 17.540 118.370 18.000 ;
        RECT 118.140 17.450 118.370 17.540 ;
        RECT 119.430 23.370 119.660 23.450 ;
        RECT 119.980 23.370 121.780 26.100 ;
        RECT 119.430 22.380 121.780 23.370 ;
        RECT 123.330 26.080 130.080 28.600 ;
        RECT 132.125 28.440 133.880 28.925 ;
        RECT 134.030 28.600 147.400 29.600 ;
        RECT 131.900 28.210 133.980 28.440 ;
        RECT 132.125 28.190 133.880 28.210 ;
        RECT 131.470 27.940 134.520 27.970 ;
        RECT 131.460 27.900 134.520 27.940 ;
        RECT 131.450 26.750 134.520 27.900 ;
        RECT 131.460 26.700 134.520 26.750 ;
        RECT 132.275 26.440 133.025 26.515 ;
        RECT 132.070 26.210 135.030 26.440 ;
        RECT 123.330 26.050 131.990 26.080 ;
        RECT 123.330 25.050 132.020 26.050 ;
        RECT 132.275 25.705 133.025 26.210 ;
        RECT 144.380 26.050 147.400 28.600 ;
        RECT 123.330 25.040 131.990 25.050 ;
        RECT 123.330 23.800 130.080 25.040 ;
        RECT 132.245 24.890 133.055 25.385 ;
        RECT 135.080 25.050 147.400 26.050 ;
        RECT 135.130 25.040 147.400 25.050 ;
        RECT 132.070 24.660 135.030 24.890 ;
        RECT 132.245 24.635 133.055 24.660 ;
        RECT 131.470 24.360 134.520 24.390 ;
        RECT 131.460 24.320 134.520 24.360 ;
        RECT 123.330 23.350 130.100 23.800 ;
        RECT 124.580 22.470 130.100 23.350 ;
        RECT 131.450 23.170 134.520 24.320 ;
        RECT 131.460 23.120 134.520 23.170 ;
        RECT 132.215 22.860 132.965 22.910 ;
        RECT 135.315 22.860 136.065 22.905 ;
        RECT 132.040 22.630 136.240 22.860 ;
        RECT 119.430 18.120 124.180 22.380 ;
        RECT 119.430 17.600 121.780 18.120 ;
        RECT 119.430 17.540 121.540 17.600 ;
        RECT 119.430 17.450 119.660 17.540 ;
        RECT 118.420 17.060 119.380 17.290 ;
        RECT 112.380 12.800 117.280 17.000 ;
        RECT 118.460 16.440 119.340 17.060 ;
        RECT 120.470 15.340 121.340 15.945 ;
        RECT 117.880 13.070 119.880 15.130 ;
        RECT 120.420 15.110 121.380 15.340 ;
        RECT 120.140 14.870 120.370 14.950 ;
        RECT 120.080 12.800 120.370 14.870 ;
        RECT 92.215 10.720 92.965 10.790 ;
        RECT 103.095 10.720 103.905 10.755 ;
        RECT 92.060 10.490 104.020 10.720 ;
        RECT 84.700 10.330 91.990 10.340 ;
        RECT 81.550 9.310 81.780 9.390 ;
        RECT 84.700 9.340 92.010 10.330 ;
        RECT 92.215 9.980 92.965 10.490 ;
        RECT 103.095 10.005 103.905 10.490 ;
        RECT 104.070 10.320 104.300 10.330 ;
        RECT 105.220 10.320 106.240 10.850 ;
        RECT 80.540 8.920 81.500 9.150 ;
        RECT 80.590 8.335 81.460 8.920 ;
        RECT 84.700 8.080 90.200 9.340 ;
        RECT 91.780 9.330 92.010 9.340 ;
        RECT 92.185 9.170 92.995 9.625 ;
        RECT 103.125 9.170 103.875 9.655 ;
        RECT 104.070 9.340 106.240 10.320 ;
        RECT 112.380 10.800 120.370 12.800 ;
        RECT 112.380 9.400 117.280 10.800 ;
        RECT 117.590 10.790 120.370 10.800 ;
        RECT 120.140 10.710 120.370 10.790 ;
        RECT 121.430 14.870 121.660 14.950 ;
        RECT 122.190 14.870 124.180 18.120 ;
        RECT 121.430 10.790 124.180 14.870 ;
        RECT 124.580 21.470 131.990 22.470 ;
        RECT 132.215 22.100 132.965 22.630 ;
        RECT 135.315 22.095 136.065 22.630 ;
        RECT 136.290 22.460 136.520 22.470 ;
        RECT 144.380 22.460 147.400 25.040 ;
        RECT 124.580 18.900 130.080 21.470 ;
        RECT 132.185 21.310 132.995 21.775 ;
        RECT 135.395 21.310 136.145 21.805 ;
        RECT 136.290 21.530 147.400 22.460 ;
        RECT 136.290 21.470 136.520 21.530 ;
        RECT 132.040 21.080 136.240 21.310 ;
        RECT 132.185 21.025 132.995 21.080 ;
        RECT 135.395 20.995 136.145 21.080 ;
        RECT 131.470 20.780 134.520 20.810 ;
        RECT 131.460 20.740 134.520 20.780 ;
        RECT 131.450 19.590 134.520 20.740 ;
        RECT 131.460 19.540 134.520 19.590 ;
        RECT 132.085 19.280 132.835 19.350 ;
        RECT 136.925 19.280 137.735 19.315 ;
        RECT 131.910 19.050 137.870 19.280 ;
        RECT 124.580 18.890 131.830 18.900 ;
        RECT 124.580 17.900 131.860 18.890 ;
        RECT 132.085 18.540 132.835 19.050 ;
        RECT 136.925 18.565 137.735 19.050 ;
        RECT 137.920 18.880 138.150 18.890 ;
        RECT 144.380 18.880 147.400 21.530 ;
        RECT 124.580 15.300 130.080 17.900 ;
        RECT 131.630 17.890 131.860 17.900 ;
        RECT 132.055 17.730 132.865 18.195 ;
        RECT 136.955 17.730 137.705 18.225 ;
        RECT 137.900 17.950 147.400 18.880 ;
        RECT 137.920 17.890 138.150 17.950 ;
        RECT 131.910 17.500 137.870 17.730 ;
        RECT 132.055 17.445 132.865 17.500 ;
        RECT 136.955 17.415 137.705 17.500 ;
        RECT 131.470 17.200 134.520 17.230 ;
        RECT 131.460 17.160 134.520 17.200 ;
        RECT 131.450 16.010 134.520 17.160 ;
        RECT 131.460 15.960 134.520 16.010 ;
        RECT 132.065 15.700 132.815 15.790 ;
        RECT 139.455 15.700 140.265 15.745 ;
        RECT 131.930 15.470 140.370 15.700 ;
        RECT 131.650 15.300 131.880 15.310 ;
        RECT 124.580 14.310 131.880 15.300 ;
        RECT 132.065 14.980 132.815 15.470 ;
        RECT 139.455 14.995 140.265 15.470 ;
        RECT 140.420 15.300 140.650 15.310 ;
        RECT 144.380 15.300 147.400 17.950 ;
        RECT 124.580 14.300 131.840 14.310 ;
        RECT 124.580 11.740 130.080 14.300 ;
        RECT 132.035 14.150 132.845 14.625 ;
        RECT 139.485 14.150 140.235 14.655 ;
        RECT 140.420 14.370 147.400 15.300 ;
        RECT 140.420 14.310 140.650 14.370 ;
        RECT 131.930 13.920 140.370 14.150 ;
        RECT 132.035 13.875 132.845 13.920 ;
        RECT 139.485 13.845 140.235 13.920 ;
        RECT 131.470 13.620 134.520 13.650 ;
        RECT 131.460 13.580 134.520 13.620 ;
        RECT 131.450 12.430 134.520 13.580 ;
        RECT 144.380 13.000 147.400 14.370 ;
        RECT 131.460 12.380 134.520 12.430 ;
        RECT 132.095 12.120 132.845 12.190 ;
        RECT 142.975 12.120 143.785 12.155 ;
        RECT 131.940 11.890 143.900 12.120 ;
        RECT 124.580 11.730 131.870 11.740 ;
        RECT 121.430 10.710 121.660 10.790 ;
        RECT 124.580 10.740 131.890 11.730 ;
        RECT 132.095 11.380 132.845 11.890 ;
        RECT 142.975 11.405 143.785 11.890 ;
        RECT 143.950 11.720 144.180 11.730 ;
        RECT 145.100 11.720 147.400 13.000 ;
        RECT 120.420 10.320 121.380 10.550 ;
        RECT 120.470 9.735 121.340 10.320 ;
        RECT 124.580 9.480 130.080 10.740 ;
        RECT 131.660 10.730 131.890 10.740 ;
        RECT 132.065 10.570 132.875 11.025 ;
        RECT 143.005 10.570 143.755 11.055 ;
        RECT 143.950 10.900 147.400 11.720 ;
        RECT 143.950 10.740 146.120 10.900 ;
        RECT 143.950 10.730 144.180 10.740 ;
        RECT 131.940 10.340 143.900 10.570 ;
        RECT 132.065 10.275 132.875 10.340 ;
        RECT 143.005 10.245 143.755 10.340 ;
        RECT 141.380 9.850 144.530 10.100 ;
        RECT 124.580 9.400 130.070 9.480 ;
        RECT 104.070 9.330 104.300 9.340 ;
        RECT 92.060 8.940 104.020 9.170 ;
        RECT 92.185 8.875 92.995 8.940 ;
        RECT 103.125 8.845 103.875 8.940 ;
        RECT 101.500 8.450 104.650 8.700 ;
        RECT 84.700 8.000 90.190 8.080 ;
        RECT 60.280 7.610 63.430 7.860 ;
        RECT 43.480 7.160 48.970 7.240 ;
        RECT 31.280 2.260 48.970 7.160 ;
        RECT 60.280 6.210 63.580 7.610 ;
        RECT 72.500 3.100 90.190 8.000 ;
        RECT 101.500 7.050 104.800 8.450 ;
        RECT 112.380 4.500 130.070 9.400 ;
        RECT 141.380 8.450 144.680 9.850 ;
        RECT 124.155 4.475 126.245 4.500 ;
        RECT 41.640 2.255 43.860 2.260 ;
      LAYER met2 ;
        RECT 78.460 220.900 78.740 220.935 ;
        RECT 26.950 217.940 27.250 217.950 ;
        RECT 26.915 217.660 27.285 217.940 ;
        RECT 26.950 215.690 27.250 217.660 ;
        RECT 34.300 217.240 34.600 217.250 ;
        RECT 34.265 216.960 34.635 217.240 ;
        RECT 26.930 215.100 27.250 215.690 ;
        RECT 34.300 215.290 34.600 216.960 ;
        RECT 41.650 216.540 41.950 216.550 ;
        RECT 41.615 216.260 41.985 216.540 ;
        RECT 26.930 212.220 27.210 215.100 ;
        RECT 34.290 214.650 34.600 215.290 ;
        RECT 41.650 214.700 41.950 216.260 ;
        RECT 63.700 214.940 64.000 214.950 ;
        RECT 49.010 214.900 49.290 214.935 ;
        RECT 34.290 212.220 34.570 214.650 ;
        RECT 41.650 212.220 41.930 214.700 ;
        RECT 49.000 213.700 49.300 214.900 ;
        RECT 56.350 214.890 56.650 214.900 ;
        RECT 56.315 214.610 56.685 214.890 ;
        RECT 63.665 214.660 64.035 214.940 ;
        RECT 71.050 214.890 71.350 214.900 ;
        RECT 56.350 213.700 56.650 214.610 ;
        RECT 63.700 214.220 64.000 214.660 ;
        RECT 71.015 214.610 71.385 214.890 ;
        RECT 71.050 214.220 71.350 214.610 ;
        RECT 78.450 214.600 78.750 220.900 ;
        RECT 85.800 220.190 86.100 220.200 ;
        RECT 85.765 219.910 86.135 220.190 ;
        RECT 63.700 213.800 64.010 214.220 ;
        RECT 49.010 212.220 49.290 213.700 ;
        RECT 56.370 212.220 56.650 213.700 ;
        RECT 56.900 212.250 57.960 212.390 ;
        RECT 27.000 203.470 27.140 212.220 ;
        RECT 34.360 204.910 34.500 212.220 ;
        RECT 38.720 206.355 40.260 206.725 ;
        RECT 41.720 205.850 41.860 212.220 ;
        RECT 48.100 207.910 48.360 208.230 ;
        RECT 41.660 205.530 41.920 205.850 ;
        RECT 33.840 204.510 34.100 204.830 ;
        RECT 34.360 204.770 34.960 204.910 ;
        RECT 36.140 204.850 36.400 205.170 ;
        RECT 47.640 204.850 47.900 205.170 ;
        RECT 26.940 203.150 27.200 203.470 ;
        RECT 32.460 201.450 32.720 201.770 ;
        RECT 29.240 191.590 29.500 191.910 ;
        RECT 24.180 188.530 24.440 188.850 ;
        RECT 24.240 181.030 24.380 188.530 ;
        RECT 29.300 188.510 29.440 191.590 ;
        RECT 30.160 190.910 30.420 191.230 ;
        RECT 25.560 188.190 25.820 188.510 ;
        RECT 27.400 188.190 27.660 188.510 ;
        RECT 29.240 188.190 29.500 188.510 ;
        RECT 25.620 187.150 25.760 188.190 ;
        RECT 25.560 186.830 25.820 187.150 ;
        RECT 24.180 180.710 24.440 181.030 ;
        RECT 25.560 180.710 25.820 181.030 ;
        RECT 25.620 178.990 25.760 180.710 ;
        RECT 25.560 178.670 25.820 178.990 ;
        RECT 27.460 171.850 27.600 188.190 ;
        RECT 29.240 182.410 29.500 182.730 ;
        RECT 29.300 177.630 29.440 182.410 ;
        RECT 29.700 178.670 29.960 178.990 ;
        RECT 29.240 177.310 29.500 177.630 ;
        RECT 29.240 174.480 29.500 174.570 ;
        RECT 29.760 174.480 29.900 178.670 ;
        RECT 30.220 177.630 30.360 190.910 ;
        RECT 32.000 188.530 32.260 188.850 ;
        RECT 31.080 187.850 31.340 188.170 ;
        RECT 31.540 187.850 31.800 188.170 ;
        RECT 31.140 187.150 31.280 187.850 ;
        RECT 31.080 186.830 31.340 187.150 ;
        RECT 31.600 186.470 31.740 187.850 ;
        RECT 31.540 186.150 31.800 186.470 ;
        RECT 32.060 185.790 32.200 188.530 ;
        RECT 32.000 185.470 32.260 185.790 ;
        RECT 32.060 183.750 32.200 185.470 ;
        RECT 32.000 183.430 32.260 183.750 ;
        RECT 32.060 181.030 32.200 183.430 ;
        RECT 32.000 180.710 32.260 181.030 ;
        RECT 30.620 180.370 30.880 180.690 ;
        RECT 30.160 177.310 30.420 177.630 ;
        RECT 29.240 174.340 29.900 174.480 ;
        RECT 29.240 174.250 29.500 174.340 ;
        RECT 29.300 172.190 29.440 174.250 ;
        RECT 30.220 173.630 30.360 177.310 ;
        RECT 30.680 175.250 30.820 180.370 ;
        RECT 31.080 179.690 31.340 180.010 ;
        RECT 31.140 177.970 31.280 179.690 ;
        RECT 31.080 177.650 31.340 177.970 ;
        RECT 31.540 175.500 31.800 175.590 ;
        RECT 32.060 175.500 32.200 180.710 ;
        RECT 31.540 175.360 32.200 175.500 ;
        RECT 31.540 175.270 31.800 175.360 ;
        RECT 30.620 174.930 30.880 175.250 ;
        RECT 29.760 173.490 30.360 173.630 ;
        RECT 29.240 171.870 29.500 172.190 ;
        RECT 25.560 171.530 25.820 171.850 ;
        RECT 27.400 171.530 27.660 171.850 ;
        RECT 25.620 170.150 25.760 171.530 ;
        RECT 25.560 169.830 25.820 170.150 ;
        RECT 24.180 169.490 24.440 169.810 ;
        RECT 24.240 161.650 24.380 169.490 ;
        RECT 26.940 163.370 27.200 163.690 ;
        RECT 24.180 161.330 24.440 161.650 ;
        RECT 24.240 158.930 24.380 161.330 ;
        RECT 24.640 160.990 24.900 161.310 ;
        RECT 24.700 159.950 24.840 160.990 ;
        RECT 27.000 159.950 27.140 163.370 ;
        RECT 24.640 159.630 24.900 159.950 ;
        RECT 26.940 159.630 27.200 159.950 ;
        RECT 24.180 158.610 24.440 158.930 ;
        RECT 24.240 153.490 24.380 158.610 ;
        RECT 26.020 155.210 26.280 155.530 ;
        RECT 25.560 153.510 25.820 153.830 ;
        RECT 24.180 153.170 24.440 153.490 ;
        RECT 24.240 142.950 24.380 153.170 ;
        RECT 25.620 151.790 25.760 153.510 ;
        RECT 25.560 151.470 25.820 151.790 ;
        RECT 26.080 150.770 26.220 155.210 ;
        RECT 27.460 151.790 27.600 171.530 ;
        RECT 29.760 162.670 29.900 173.490 ;
        RECT 30.160 172.890 30.420 173.210 ;
        RECT 27.860 162.350 28.120 162.670 ;
        RECT 29.700 162.350 29.960 162.670 ;
        RECT 27.920 159.610 28.060 162.350 ;
        RECT 30.220 162.330 30.360 172.890 ;
        RECT 30.680 172.190 30.820 174.930 ;
        RECT 31.600 173.550 31.740 175.270 ;
        RECT 32.520 174.990 32.660 201.450 ;
        RECT 33.380 193.290 33.640 193.610 ;
        RECT 33.440 190.890 33.580 193.290 ;
        RECT 33.380 190.570 33.640 190.890 ;
        RECT 33.900 190.630 34.040 204.510 ;
        RECT 34.820 204.490 34.960 204.770 ;
        RECT 34.760 204.170 35.020 204.490 ;
        RECT 36.200 203.130 36.340 204.850 ;
        RECT 41.660 204.510 41.920 204.830 ;
        RECT 37.060 204.170 37.320 204.490 ;
        RECT 36.140 202.810 36.400 203.130 ;
        RECT 36.600 202.470 36.860 202.790 ;
        RECT 36.660 198.030 36.800 202.470 ;
        RECT 35.220 197.710 35.480 198.030 ;
        RECT 36.600 197.710 36.860 198.030 ;
        RECT 34.300 196.010 34.560 196.330 ;
        RECT 34.360 193.610 34.500 196.010 ;
        RECT 34.300 193.290 34.560 193.610 ;
        RECT 35.280 191.570 35.420 197.710 ;
        RECT 36.140 193.970 36.400 194.290 ;
        RECT 35.680 193.630 35.940 193.950 ;
        RECT 35.740 191.990 35.880 193.630 ;
        RECT 36.200 192.590 36.340 193.970 ;
        RECT 36.600 193.290 36.860 193.610 ;
        RECT 36.140 192.270 36.400 192.590 ;
        RECT 35.740 191.910 36.340 191.990 ;
        RECT 35.740 191.850 36.400 191.910 ;
        RECT 36.140 191.590 36.400 191.850 ;
        RECT 35.220 191.250 35.480 191.570 ;
        RECT 33.900 190.490 34.960 190.630 ;
        RECT 35.680 190.570 35.940 190.890 ;
        RECT 33.840 189.550 34.100 189.870 ;
        RECT 33.900 187.150 34.040 189.550 ;
        RECT 33.840 186.830 34.100 187.150 ;
        RECT 33.840 183.770 34.100 184.090 ;
        RECT 33.380 183.430 33.640 183.750 ;
        RECT 32.920 182.410 33.180 182.730 ;
        RECT 32.980 178.990 33.120 182.410 ;
        RECT 33.440 181.710 33.580 183.430 ;
        RECT 33.380 181.390 33.640 181.710 ;
        RECT 33.380 179.690 33.640 180.010 ;
        RECT 32.920 178.670 33.180 178.990 ;
        RECT 32.920 177.990 33.180 178.310 ;
        RECT 32.980 175.930 33.120 177.990 ;
        RECT 33.440 177.630 33.580 179.690 ;
        RECT 33.900 178.310 34.040 183.770 ;
        RECT 34.300 183.090 34.560 183.410 ;
        RECT 34.360 178.990 34.500 183.090 ;
        RECT 34.300 178.670 34.560 178.990 ;
        RECT 33.840 177.990 34.100 178.310 ;
        RECT 33.380 177.310 33.640 177.630 ;
        RECT 32.920 175.610 33.180 175.930 ;
        RECT 32.060 174.850 32.660 174.990 ;
        RECT 31.540 173.230 31.800 173.550 ;
        RECT 30.620 171.870 30.880 172.190 ;
        RECT 31.540 171.530 31.800 171.850 ;
        RECT 31.600 168.110 31.740 171.530 ;
        RECT 31.540 167.790 31.800 168.110 ;
        RECT 32.060 167.510 32.200 174.850 ;
        RECT 32.980 173.550 33.120 175.610 ;
        RECT 34.300 175.270 34.560 175.590 ;
        RECT 33.380 174.250 33.640 174.570 ;
        RECT 33.840 174.250 34.100 174.570 ;
        RECT 32.920 173.230 33.180 173.550 ;
        RECT 32.460 171.530 32.720 171.850 ;
        RECT 30.680 167.370 32.200 167.510 ;
        RECT 30.160 162.010 30.420 162.330 ;
        RECT 27.860 159.290 28.120 159.610 ;
        RECT 27.920 155.870 28.060 159.290 ;
        RECT 30.220 156.550 30.360 162.010 ;
        RECT 30.160 156.230 30.420 156.550 ;
        RECT 27.860 155.550 28.120 155.870 ;
        RECT 27.400 151.470 27.660 151.790 ;
        RECT 26.020 150.450 26.280 150.770 ;
        RECT 26.480 145.010 26.740 145.330 ;
        RECT 25.560 144.330 25.820 144.650 ;
        RECT 25.620 143.290 25.760 144.330 ;
        RECT 25.560 142.970 25.820 143.290 ;
        RECT 24.180 142.630 24.440 142.950 ;
        RECT 26.540 140.910 26.680 145.010 ;
        RECT 27.460 140.910 27.600 151.470 ;
        RECT 26.480 140.590 26.740 140.910 ;
        RECT 27.400 140.590 27.660 140.910 ;
        RECT 27.920 138.190 28.060 155.550 ;
        RECT 29.240 155.210 29.500 155.530 ;
        RECT 29.300 150.770 29.440 155.210 ;
        RECT 30.220 153.830 30.360 156.230 ;
        RECT 30.160 153.510 30.420 153.830 ;
        RECT 30.160 151.130 30.420 151.450 ;
        RECT 29.240 150.450 29.500 150.770 ;
        RECT 30.220 145.330 30.360 151.130 ;
        RECT 30.160 145.010 30.420 145.330 ;
        RECT 29.240 144.330 29.500 144.650 ;
        RECT 29.700 144.330 29.960 144.650 ;
        RECT 29.300 140.570 29.440 144.330 ;
        RECT 29.240 140.250 29.500 140.570 ;
        RECT 29.300 139.210 29.440 140.250 ;
        RECT 29.760 139.550 29.900 144.330 ;
        RECT 29.700 139.230 29.960 139.550 ;
        RECT 29.240 138.890 29.500 139.210 ;
        RECT 27.860 137.870 28.120 138.190 ;
        RECT 29.300 135.550 29.440 138.890 ;
        RECT 29.300 135.410 29.900 135.550 ;
        RECT 29.240 134.470 29.500 134.790 ;
        RECT 27.400 133.450 27.660 133.770 ;
        RECT 27.460 132.070 27.600 133.450 ;
        RECT 27.400 131.750 27.660 132.070 ;
        RECT 28.310 131.895 28.590 132.265 ;
        RECT 29.300 132.070 29.440 134.470 ;
        RECT 29.760 134.450 29.900 135.410 ;
        RECT 29.700 134.130 29.960 134.450 ;
        RECT 28.320 131.750 28.580 131.895 ;
        RECT 29.240 131.750 29.500 132.070 ;
        RECT 26.940 131.070 27.200 131.390 ;
        RECT 26.020 130.730 26.280 131.050 ;
        RECT 26.080 128.670 26.220 130.730 ;
        RECT 27.000 129.010 27.140 131.070 ;
        RECT 26.940 128.690 27.200 129.010 ;
        RECT 26.020 128.350 26.280 128.670 ;
        RECT 27.000 123.570 27.140 128.690 ;
        RECT 28.380 126.970 28.520 131.750 ;
        RECT 29.300 128.070 29.440 131.750 ;
        RECT 29.300 127.930 29.900 128.070 ;
        RECT 28.320 126.650 28.580 126.970 ;
        RECT 27.860 125.290 28.120 125.610 ;
        RECT 26.940 123.250 27.200 123.570 ;
        RECT 26.480 122.910 26.740 123.230 ;
        RECT 26.540 121.870 26.680 122.910 ;
        RECT 26.480 121.550 26.740 121.870 ;
        RECT 27.000 116.090 27.140 123.250 ;
        RECT 27.920 118.130 28.060 125.290 ;
        RECT 28.780 122.570 29.040 122.890 ;
        RECT 28.320 118.490 28.580 118.810 ;
        RECT 27.860 117.810 28.120 118.130 ;
        RECT 26.940 115.770 27.200 116.090 ;
        RECT 25.560 115.430 25.820 115.750 ;
        RECT 25.620 113.710 25.760 115.430 ;
        RECT 25.560 113.390 25.820 113.710 ;
        RECT 26.940 112.370 27.200 112.690 ;
        RECT 27.000 110.990 27.140 112.370 ;
        RECT 26.940 110.670 27.200 110.990 ;
        RECT 28.380 110.310 28.520 118.490 ;
        RECT 28.840 118.470 28.980 122.570 ;
        RECT 29.240 120.530 29.500 120.850 ;
        RECT 29.300 119.150 29.440 120.530 ;
        RECT 29.240 118.830 29.500 119.150 ;
        RECT 29.760 118.550 29.900 127.930 ;
        RECT 30.160 126.990 30.420 127.310 ;
        RECT 30.220 118.810 30.360 126.990 ;
        RECT 29.300 118.470 29.900 118.550 ;
        RECT 30.160 118.490 30.420 118.810 ;
        RECT 28.780 118.150 29.040 118.470 ;
        RECT 29.240 118.410 29.900 118.470 ;
        RECT 29.240 118.150 29.500 118.410 ;
        RECT 30.680 116.430 30.820 167.370 ;
        RECT 31.080 164.690 31.340 164.710 ;
        RECT 32.520 164.690 32.660 171.530 ;
        RECT 32.980 170.150 33.120 173.230 ;
        RECT 33.440 172.190 33.580 174.250 ;
        RECT 33.900 172.870 34.040 174.250 ;
        RECT 33.840 172.550 34.100 172.870 ;
        RECT 33.380 171.870 33.640 172.190 ;
        RECT 33.900 170.490 34.040 172.550 ;
        RECT 34.360 172.190 34.500 175.270 ;
        RECT 34.300 171.870 34.560 172.190 ;
        RECT 34.360 170.830 34.500 171.870 ;
        RECT 34.300 170.510 34.560 170.830 ;
        RECT 33.840 170.170 34.100 170.490 ;
        RECT 32.920 169.830 33.180 170.150 ;
        RECT 32.980 167.090 33.120 169.830 ;
        RECT 34.360 167.090 34.500 170.510 ;
        RECT 32.920 166.770 33.180 167.090 ;
        RECT 34.300 166.770 34.560 167.090 ;
        RECT 33.380 166.090 33.640 166.410 ;
        RECT 31.080 164.550 32.660 164.690 ;
        RECT 31.080 164.390 31.340 164.550 ;
        RECT 32.000 157.930 32.260 158.250 ;
        RECT 31.540 156.910 31.800 157.230 ;
        RECT 31.080 155.890 31.340 156.210 ;
        RECT 31.140 154.510 31.280 155.890 ;
        RECT 31.600 154.510 31.740 156.910 ;
        RECT 32.060 156.210 32.200 157.930 ;
        RECT 32.000 155.890 32.260 156.210 ;
        RECT 32.520 155.530 32.660 164.550 ;
        RECT 32.920 164.690 33.180 164.710 ;
        RECT 33.440 164.690 33.580 166.090 ;
        RECT 32.920 164.550 33.580 164.690 ;
        RECT 32.920 164.390 33.180 164.550 ;
        RECT 32.980 160.970 33.120 164.390 ;
        RECT 34.820 162.070 34.960 190.490 ;
        RECT 35.220 188.870 35.480 189.190 ;
        RECT 35.280 186.470 35.420 188.870 ;
        RECT 35.740 186.470 35.880 190.570 ;
        RECT 36.200 189.190 36.340 191.590 ;
        RECT 36.660 191.570 36.800 193.290 ;
        RECT 36.600 191.250 36.860 191.570 ;
        RECT 36.140 188.870 36.400 189.190 ;
        RECT 35.220 186.150 35.480 186.470 ;
        RECT 35.680 186.150 35.940 186.470 ;
        RECT 36.660 185.790 36.800 191.250 ;
        RECT 36.600 185.470 36.860 185.790 ;
        RECT 36.140 182.750 36.400 183.070 ;
        RECT 35.220 182.410 35.480 182.730 ;
        RECT 35.280 181.030 35.420 182.410 ;
        RECT 35.220 180.710 35.480 181.030 ;
        RECT 35.220 177.990 35.480 178.310 ;
        RECT 35.280 170.150 35.420 177.990 ;
        RECT 35.220 169.830 35.480 170.150 ;
        RECT 35.680 166.430 35.940 166.750 ;
        RECT 35.740 164.370 35.880 166.430 ;
        RECT 35.680 164.050 35.940 164.370 ;
        RECT 34.820 161.930 35.880 162.070 ;
        RECT 34.760 160.990 35.020 161.310 ;
        RECT 32.920 160.650 33.180 160.970 ;
        RECT 33.380 160.650 33.640 160.970 ;
        RECT 34.300 160.650 34.560 160.970 ;
        RECT 32.980 156.630 33.120 160.650 ;
        RECT 33.440 157.230 33.580 160.650 ;
        RECT 34.360 159.270 34.500 160.650 ;
        RECT 34.300 158.950 34.560 159.270 ;
        RECT 33.840 158.610 34.100 158.930 ;
        RECT 33.380 156.910 33.640 157.230 ;
        RECT 32.980 156.490 33.580 156.630 ;
        RECT 33.440 156.210 33.580 156.490 ;
        RECT 33.380 155.890 33.640 156.210 ;
        RECT 33.900 155.870 34.040 158.610 ;
        RECT 34.820 158.590 34.960 160.990 ;
        RECT 34.760 158.270 35.020 158.590 ;
        RECT 33.840 155.550 34.100 155.870 ;
        RECT 32.460 155.210 32.720 155.530 ;
        RECT 31.080 154.190 31.340 154.510 ;
        RECT 31.540 154.190 31.800 154.510 ;
        RECT 33.380 153.510 33.640 153.830 ;
        RECT 33.840 153.510 34.100 153.830 ;
        RECT 32.460 150.110 32.720 150.430 ;
        RECT 32.520 149.070 32.660 150.110 ;
        RECT 33.440 150.090 33.580 153.510 ;
        RECT 33.900 151.790 34.040 153.510 ;
        RECT 34.760 152.490 35.020 152.810 ;
        RECT 33.840 151.470 34.100 151.790 ;
        RECT 33.380 149.770 33.640 150.090 ;
        RECT 32.460 148.750 32.720 149.070 ;
        RECT 34.820 148.730 34.960 152.490 ;
        RECT 34.760 148.410 35.020 148.730 ;
        RECT 31.080 145.010 31.340 145.330 ;
        RECT 31.140 143.630 31.280 145.010 ;
        RECT 33.380 144.670 33.640 144.990 ;
        RECT 31.080 143.310 31.340 143.630 ;
        RECT 33.440 142.610 33.580 144.670 ;
        RECT 35.220 142.630 35.480 142.950 ;
        RECT 32.460 142.290 32.720 142.610 ;
        RECT 33.380 142.290 33.640 142.610 ;
        RECT 32.520 140.990 32.660 142.290 ;
        RECT 34.300 141.610 34.560 141.930 ;
        RECT 31.080 140.820 31.340 140.910 ;
        RECT 32.060 140.850 32.660 140.990 ;
        RECT 32.060 140.820 32.200 140.850 ;
        RECT 31.080 140.680 32.200 140.820 ;
        RECT 31.080 140.590 31.340 140.680 ;
        RECT 31.140 135.130 31.280 140.590 ;
        RECT 32.460 140.250 32.720 140.570 ;
        RECT 32.000 137.870 32.260 138.190 ;
        RECT 31.080 134.810 31.340 135.130 ;
        RECT 32.060 134.450 32.200 137.870 ;
        RECT 32.520 137.510 32.660 140.250 ;
        RECT 33.380 139.910 33.640 140.230 ;
        RECT 33.440 138.190 33.580 139.910 ;
        RECT 34.360 139.550 34.500 141.610 ;
        RECT 35.280 140.910 35.420 142.630 ;
        RECT 35.220 140.590 35.480 140.910 ;
        RECT 35.740 140.310 35.880 161.930 ;
        RECT 36.200 159.950 36.340 182.750 ;
        RECT 36.600 169.490 36.860 169.810 ;
        RECT 36.660 168.110 36.800 169.490 ;
        RECT 36.600 167.790 36.860 168.110 ;
        RECT 37.120 164.690 37.260 204.170 ;
        RECT 41.720 203.470 41.860 204.510 ;
        RECT 41.660 203.150 41.920 203.470 ;
        RECT 47.700 203.130 47.840 204.850 ;
        RECT 37.520 202.810 37.780 203.130 ;
        RECT 47.640 202.810 47.900 203.130 ;
        RECT 37.580 200.070 37.720 202.810 ;
        RECT 40.740 202.470 41.000 202.790 ;
        RECT 37.980 201.450 38.240 201.770 ;
        RECT 37.520 199.750 37.780 200.070 ;
        RECT 37.580 197.690 37.720 199.750 ;
        RECT 38.040 199.730 38.180 201.450 ;
        RECT 38.720 200.915 40.260 201.285 ;
        RECT 37.980 199.410 38.240 199.730 ;
        RECT 40.800 198.030 40.940 202.470 ;
        RECT 48.160 199.730 48.300 207.910 ;
        RECT 49.080 204.830 49.220 212.220 ;
        RECT 56.440 211.710 56.580 212.220 ;
        RECT 56.900 211.710 57.040 212.250 ;
        RECT 56.440 211.570 57.040 211.710 ;
        RECT 55.510 209.075 57.050 209.445 ;
        RECT 57.820 208.230 57.960 212.250 ;
        RECT 63.730 212.220 64.010 213.800 ;
        RECT 71.050 213.700 71.370 214.220 ;
        RECT 71.090 212.220 71.370 213.700 ;
        RECT 78.450 212.220 78.730 214.600 ;
        RECT 85.800 213.700 86.100 219.910 ;
        RECT 93.160 219.550 93.440 219.585 ;
        RECT 93.150 213.700 93.450 219.550 ;
        RECT 100.560 218.850 100.840 218.885 ;
        RECT 100.550 214.220 100.850 218.850 ;
        RECT 107.910 218.150 108.190 218.185 ;
        RECT 107.900 214.220 108.200 218.150 ;
        RECT 115.260 217.400 115.540 217.435 ;
        RECT 85.810 212.220 86.090 213.700 ;
        RECT 93.170 212.220 93.450 213.700 ;
        RECT 100.530 213.700 100.850 214.220 ;
        RECT 107.890 213.700 108.200 214.220 ;
        RECT 115.250 213.700 115.550 217.400 ;
        RECT 122.610 216.750 122.890 216.785 ;
        RECT 122.600 213.700 122.900 216.750 ;
        RECT 129.950 216.090 130.250 216.100 ;
        RECT 129.915 215.810 130.285 216.090 ;
        RECT 129.950 213.700 130.250 215.810 ;
        RECT 137.300 215.460 137.580 215.495 ;
        RECT 137.290 214.220 137.590 215.460 ;
        RECT 144.690 214.790 144.970 214.825 ;
        RECT 137.290 213.700 137.610 214.220 ;
        RECT 144.680 213.700 144.980 214.790 ;
        RECT 152.050 214.140 152.330 214.220 ;
        RECT 152.570 214.140 152.850 214.175 ;
        RECT 152.040 213.840 152.860 214.140 ;
        RECT 152.040 213.700 152.340 213.840 ;
        RECT 152.570 213.805 152.850 213.840 ;
        RECT 100.530 212.220 100.810 213.700 ;
        RECT 107.890 212.220 108.170 213.700 ;
        RECT 108.420 212.250 109.940 212.390 ;
        RECT 63.800 208.230 63.940 212.220 ;
        RECT 70.640 208.250 70.900 208.570 ;
        RECT 57.760 207.910 58.020 208.230 ;
        RECT 63.740 207.910 64.000 208.230 ;
        RECT 54.540 207.630 54.800 207.890 ;
        RECT 54.140 207.570 54.800 207.630 ;
        RECT 60.060 207.570 60.320 207.890 ;
        RECT 51.780 207.230 52.040 207.550 ;
        RECT 54.140 207.490 54.740 207.570 ;
        RECT 51.320 206.890 51.580 207.210 ;
        RECT 49.020 204.510 49.280 204.830 ;
        RECT 50.400 204.170 50.660 204.490 ;
        RECT 49.940 202.470 50.200 202.790 ;
        RECT 49.020 202.130 49.280 202.450 ;
        RECT 48.560 200.090 48.820 200.410 ;
        RECT 48.620 199.730 48.760 200.090 ;
        RECT 48.100 199.410 48.360 199.730 ;
        RECT 48.560 199.410 48.820 199.730 ;
        RECT 46.720 199.070 46.980 199.390 ;
        RECT 44.880 198.730 45.140 199.050 ;
        RECT 44.940 198.030 45.080 198.730 ;
        RECT 40.740 197.710 41.000 198.030 ;
        RECT 44.880 197.710 45.140 198.030 ;
        RECT 37.520 197.370 37.780 197.690 ;
        RECT 46.780 197.350 46.920 199.070 ;
        RECT 47.640 198.730 47.900 199.050 ;
        RECT 48.100 198.730 48.360 199.050 ;
        RECT 37.980 197.030 38.240 197.350 ;
        RECT 46.720 197.030 46.980 197.350 ;
        RECT 38.040 195.310 38.180 197.030 ;
        RECT 38.720 195.475 40.260 195.845 ;
        RECT 37.980 194.990 38.240 195.310 ;
        RECT 46.780 194.290 46.920 197.030 ;
        RECT 40.740 193.970 41.000 194.290 ;
        RECT 46.720 193.970 46.980 194.290 ;
        RECT 39.360 193.290 39.620 193.610 ;
        RECT 39.420 192.250 39.560 193.290 ;
        RECT 39.360 191.930 39.620 192.250 ;
        RECT 37.980 191.590 38.240 191.910 ;
        RECT 37.520 185.810 37.780 186.130 ;
        RECT 37.580 177.970 37.720 185.810 ;
        RECT 38.040 183.070 38.180 191.590 ;
        RECT 38.720 190.035 40.260 190.405 ;
        RECT 40.800 189.870 40.940 193.970 ;
        RECT 46.780 191.910 46.920 193.970 ;
        RECT 46.720 191.590 46.980 191.910 ;
        RECT 44.420 190.570 44.680 190.890 ;
        RECT 45.800 190.570 46.060 190.890 ;
        RECT 40.740 189.550 41.000 189.870 ;
        RECT 44.480 188.760 44.620 190.570 ;
        RECT 45.860 189.530 46.000 190.570 ;
        RECT 45.800 189.210 46.060 189.530 ;
        RECT 46.780 189.190 46.920 191.590 ;
        RECT 46.720 188.870 46.980 189.190 ;
        RECT 44.880 188.760 45.140 188.850 ;
        RECT 44.480 188.620 45.140 188.760 ;
        RECT 41.660 186.150 41.920 186.470 ;
        RECT 40.740 185.470 41.000 185.790 ;
        RECT 38.720 184.595 40.260 184.965 ;
        RECT 40.800 183.830 40.940 185.470 ;
        RECT 40.340 183.690 40.940 183.830 ;
        RECT 37.980 182.750 38.240 183.070 ;
        RECT 38.040 181.370 38.180 182.750 ;
        RECT 37.980 181.050 38.240 181.370 ;
        RECT 37.520 177.650 37.780 177.970 ;
        RECT 38.040 174.910 38.180 181.050 ;
        RECT 40.340 179.920 40.480 183.690 ;
        RECT 41.200 182.410 41.460 182.730 ;
        RECT 40.340 179.780 40.940 179.920 ;
        RECT 38.720 179.155 40.260 179.525 ;
        RECT 40.800 178.990 40.940 179.780 ;
        RECT 40.740 178.670 41.000 178.990 ;
        RECT 37.980 174.590 38.240 174.910 ;
        RECT 40.740 174.250 41.000 174.570 ;
        RECT 38.720 173.715 40.260 174.085 ;
        RECT 38.900 172.385 39.160 172.530 ;
        RECT 39.360 172.440 39.620 172.530 ;
        RECT 40.800 172.440 40.940 174.250 ;
        RECT 38.440 171.870 38.700 172.190 ;
        RECT 38.890 172.015 39.170 172.385 ;
        RECT 39.360 172.300 40.940 172.440 ;
        RECT 39.360 172.210 39.620 172.300 ;
        RECT 38.500 170.150 38.640 171.870 ;
        RECT 38.960 170.830 39.100 172.015 ;
        RECT 38.900 170.510 39.160 170.830 ;
        RECT 40.800 170.490 40.940 172.300 ;
        RECT 40.740 170.170 41.000 170.490 ;
        RECT 38.440 169.830 38.700 170.150 ;
        RECT 37.980 169.490 38.240 169.810 ;
        RECT 37.520 169.150 37.780 169.470 ;
        RECT 37.580 165.390 37.720 169.150 ;
        RECT 38.040 168.110 38.180 169.490 ;
        RECT 38.720 168.275 40.260 168.645 ;
        RECT 37.980 167.790 38.240 168.110 ;
        RECT 41.260 166.410 41.400 182.410 ;
        RECT 41.720 172.530 41.860 186.150 ;
        RECT 43.040 185.130 43.300 185.450 ;
        RECT 42.120 183.090 42.380 183.410 ;
        RECT 42.180 181.710 42.320 183.090 ;
        RECT 42.120 181.390 42.380 181.710 ;
        RECT 43.100 180.010 43.240 185.130 ;
        RECT 44.480 180.690 44.620 188.620 ;
        RECT 44.880 188.530 45.140 188.620 ;
        RECT 47.700 188.170 47.840 198.730 ;
        RECT 48.160 196.330 48.300 198.730 ;
        RECT 48.100 196.010 48.360 196.330 ;
        RECT 48.620 194.290 48.760 199.410 ;
        RECT 49.080 198.030 49.220 202.130 ;
        RECT 49.020 197.710 49.280 198.030 ;
        RECT 48.560 193.970 48.820 194.290 ;
        RECT 48.620 192.250 48.760 193.970 ;
        RECT 49.480 193.290 49.740 193.610 ;
        RECT 48.560 191.930 48.820 192.250 ;
        RECT 48.100 191.250 48.360 191.570 ;
        RECT 48.160 189.870 48.300 191.250 ;
        RECT 48.620 189.870 48.760 191.930 ;
        RECT 49.540 191.910 49.680 193.290 ;
        RECT 49.480 191.590 49.740 191.910 ;
        RECT 49.020 190.570 49.280 190.890 ;
        RECT 48.100 189.550 48.360 189.870 ;
        RECT 48.560 189.550 48.820 189.870 ;
        RECT 47.640 187.850 47.900 188.170 ;
        RECT 48.160 187.150 48.300 189.550 ;
        RECT 48.560 188.190 48.820 188.510 ;
        RECT 48.100 186.830 48.360 187.150 ;
        RECT 47.180 186.380 47.440 186.470 ;
        RECT 47.180 186.240 47.840 186.380 ;
        RECT 47.180 186.150 47.440 186.240 ;
        RECT 44.880 185.130 45.140 185.450 ;
        RECT 44.940 183.750 45.080 185.130 ;
        RECT 44.880 183.430 45.140 183.750 ;
        RECT 45.340 183.090 45.600 183.410 ;
        RECT 45.800 183.090 46.060 183.410 ;
        RECT 45.400 181.030 45.540 183.090 ;
        RECT 44.880 180.710 45.140 181.030 ;
        RECT 45.340 180.710 45.600 181.030 ;
        RECT 44.420 180.370 44.680 180.690 ;
        RECT 43.040 179.690 43.300 180.010 ;
        RECT 44.480 177.970 44.620 180.370 ;
        RECT 44.940 178.310 45.080 180.710 ;
        RECT 45.400 178.990 45.540 180.710 ;
        RECT 45.340 178.670 45.600 178.990 ;
        RECT 44.880 177.990 45.140 178.310 ;
        RECT 44.420 177.650 44.680 177.970 ;
        RECT 43.960 175.270 44.220 175.590 ;
        RECT 44.020 173.550 44.160 175.270 ;
        RECT 44.420 174.250 44.680 174.570 ;
        RECT 43.960 173.230 44.220 173.550 ;
        RECT 42.580 172.550 42.840 172.870 ;
        RECT 41.660 172.210 41.920 172.530 ;
        RECT 41.720 170.150 41.860 172.210 ;
        RECT 42.640 172.190 42.780 172.550 ;
        RECT 44.480 172.530 44.620 174.250 ;
        RECT 45.860 173.550 46.000 183.090 ;
        RECT 47.700 181.710 47.840 186.240 ;
        RECT 47.640 181.390 47.900 181.710 ;
        RECT 46.720 180.370 46.980 180.690 ;
        RECT 46.780 178.990 46.920 180.370 ;
        RECT 46.720 178.670 46.980 178.990 ;
        RECT 48.620 176.350 48.760 188.190 ;
        RECT 49.080 186.470 49.220 190.570 ;
        RECT 49.480 187.850 49.740 188.170 ;
        RECT 49.020 186.150 49.280 186.470 ;
        RECT 49.540 185.985 49.680 187.850 ;
        RECT 49.470 185.615 49.750 185.985 ;
        RECT 47.700 176.210 48.760 176.350 ;
        RECT 47.180 174.590 47.440 174.910 ;
        RECT 45.800 173.230 46.060 173.550 ;
        RECT 46.720 173.230 46.980 173.550 ;
        RECT 44.420 172.210 44.680 172.530 ;
        RECT 44.880 172.385 45.140 172.530 ;
        RECT 42.580 172.100 42.840 172.190 ;
        RECT 42.180 171.960 42.840 172.100 ;
        RECT 44.870 172.015 45.150 172.385 ;
        RECT 45.340 172.210 45.600 172.530 ;
        RECT 41.660 169.830 41.920 170.150 ;
        RECT 42.180 169.810 42.320 171.960 ;
        RECT 42.580 171.870 42.840 171.960 ;
        RECT 43.040 171.760 43.300 171.850 ;
        RECT 43.040 171.620 44.160 171.760 ;
        RECT 43.040 171.530 43.300 171.620 ;
        RECT 44.020 170.150 44.160 171.620 ;
        RECT 45.400 170.830 45.540 172.210 ;
        RECT 45.340 170.510 45.600 170.830 ;
        RECT 43.960 169.830 44.220 170.150 ;
        RECT 42.120 169.490 42.380 169.810 ;
        RECT 42.580 168.810 42.840 169.130 ;
        RECT 42.640 167.090 42.780 168.810 ;
        RECT 46.260 167.790 46.520 168.110 ;
        RECT 43.040 167.450 43.300 167.770 ;
        RECT 42.580 166.770 42.840 167.090 ;
        RECT 41.200 166.090 41.460 166.410 ;
        RECT 37.520 165.070 37.780 165.390 ;
        RECT 37.120 164.550 37.720 164.690 ;
        RECT 36.600 164.050 36.860 164.370 ;
        RECT 36.660 160.970 36.800 164.050 ;
        RECT 36.600 160.650 36.860 160.970 ;
        RECT 36.140 159.630 36.400 159.950 ;
        RECT 36.660 159.270 36.800 160.650 ;
        RECT 36.600 158.950 36.860 159.270 ;
        RECT 36.600 155.890 36.860 156.210 ;
        RECT 36.660 153.830 36.800 155.890 ;
        RECT 36.600 153.510 36.860 153.830 ;
        RECT 36.660 151.790 36.800 153.510 ;
        RECT 36.600 151.470 36.860 151.790 ;
        RECT 36.140 141.950 36.400 142.270 ;
        RECT 36.200 140.910 36.340 141.950 ;
        RECT 36.600 141.610 36.860 141.930 ;
        RECT 36.140 140.590 36.400 140.910 ;
        RECT 35.280 140.170 35.880 140.310 ;
        RECT 34.300 139.230 34.560 139.550 ;
        RECT 33.380 137.870 33.640 138.190 ;
        RECT 32.460 137.190 32.720 137.510 ;
        RECT 32.920 136.510 33.180 136.830 ;
        RECT 32.460 136.170 32.720 136.490 ;
        RECT 32.520 135.130 32.660 136.170 ;
        RECT 32.460 134.810 32.720 135.130 ;
        RECT 32.520 134.450 32.660 134.810 ;
        RECT 32.000 134.130 32.260 134.450 ;
        RECT 32.460 134.130 32.720 134.450 ;
        RECT 32.520 130.030 32.660 134.130 ;
        RECT 32.980 132.070 33.120 136.510 ;
        RECT 32.920 131.750 33.180 132.070 ;
        RECT 32.980 131.050 33.120 131.750 ;
        RECT 32.920 130.730 33.180 131.050 ;
        RECT 32.460 129.710 32.720 130.030 ;
        RECT 31.080 125.290 31.340 125.610 ;
        RECT 34.760 125.520 35.020 125.610 ;
        RECT 34.360 125.380 35.020 125.520 ;
        RECT 31.140 124.590 31.280 125.290 ;
        RECT 31.080 124.270 31.340 124.590 ;
        RECT 31.540 120.190 31.800 120.510 ;
        RECT 31.600 118.130 31.740 120.190 ;
        RECT 33.380 119.850 33.640 120.170 ;
        RECT 31.540 117.810 31.800 118.130 ;
        RECT 31.080 117.130 31.340 117.450 ;
        RECT 30.620 116.110 30.880 116.430 ;
        RECT 31.140 114.730 31.280 117.130 ;
        RECT 31.080 114.410 31.340 114.730 ;
        RECT 31.140 113.030 31.280 114.410 ;
        RECT 31.080 112.710 31.340 113.030 ;
        RECT 29.240 111.690 29.500 112.010 ;
        RECT 29.300 110.310 29.440 111.690 ;
        RECT 28.320 109.990 28.580 110.310 ;
        RECT 29.240 109.990 29.500 110.310 ;
        RECT 31.600 109.970 31.740 117.810 ;
        RECT 32.920 117.130 33.180 117.450 ;
        RECT 32.980 116.090 33.120 117.130 ;
        RECT 32.920 115.770 33.180 116.090 ;
        RECT 31.540 109.650 31.800 109.970 ;
        RECT 33.440 109.290 33.580 119.850 ;
        RECT 33.840 117.810 34.100 118.130 ;
        RECT 33.900 109.630 34.040 117.810 ;
        RECT 34.360 117.790 34.500 125.380 ;
        RECT 34.760 125.290 35.020 125.380 ;
        RECT 34.760 118.490 35.020 118.810 ;
        RECT 34.300 117.470 34.560 117.790 ;
        RECT 33.840 109.310 34.100 109.630 ;
        RECT 32.460 108.970 32.720 109.290 ;
        RECT 33.380 108.970 33.640 109.290 ;
        RECT 31.540 106.250 31.800 106.570 ;
        RECT 31.600 104.530 31.740 106.250 ;
        RECT 31.540 104.385 31.800 104.530 ;
        RECT 31.530 104.015 31.810 104.385 ;
        RECT 32.520 101.810 32.660 108.970 ;
        RECT 34.820 107.590 34.960 118.490 ;
        RECT 34.760 107.270 35.020 107.590 ;
        RECT 32.920 106.930 33.180 107.250 ;
        RECT 33.840 106.930 34.100 107.250 ;
        RECT 32.980 104.870 33.120 106.930 ;
        RECT 33.900 105.630 34.040 106.930 ;
        RECT 34.760 106.250 35.020 106.570 ;
        RECT 35.280 106.310 35.420 140.170 ;
        RECT 36.660 137.510 36.800 141.610 ;
        RECT 36.600 137.190 36.860 137.510 ;
        RECT 36.600 134.130 36.860 134.450 ;
        RECT 36.660 132.750 36.800 134.130 ;
        RECT 36.600 132.430 36.860 132.750 ;
        RECT 36.660 127.310 36.800 132.430 ;
        RECT 36.600 126.990 36.860 127.310 ;
        RECT 36.660 126.630 36.800 126.990 ;
        RECT 35.680 126.310 35.940 126.630 ;
        RECT 36.600 126.310 36.860 126.630 ;
        RECT 35.740 124.590 35.880 126.310 ;
        RECT 35.680 124.270 35.940 124.590 ;
        RECT 35.740 121.190 35.880 124.270 ;
        RECT 36.660 121.870 36.800 126.310 ;
        RECT 37.060 123.250 37.320 123.570 ;
        RECT 36.600 121.550 36.860 121.870 ;
        RECT 37.120 121.190 37.260 123.250 ;
        RECT 35.680 120.870 35.940 121.190 ;
        RECT 37.060 120.870 37.320 121.190 ;
        RECT 36.140 117.130 36.400 117.450 ;
        RECT 36.200 110.990 36.340 117.130 ;
        RECT 37.060 115.430 37.320 115.750 ;
        RECT 37.120 112.690 37.260 115.430 ;
        RECT 37.060 112.370 37.320 112.690 ;
        RECT 37.060 111.690 37.320 112.010 ;
        RECT 36.140 110.670 36.400 110.990 ;
        RECT 37.120 109.970 37.260 111.690 ;
        RECT 37.060 109.650 37.320 109.970 ;
        RECT 37.580 108.270 37.720 164.550 ;
        RECT 38.720 162.835 40.260 163.205 ;
        RECT 41.200 162.350 41.460 162.670 ;
        RECT 40.740 160.990 41.000 161.310 ;
        RECT 40.800 158.930 40.940 160.990 ;
        RECT 40.740 158.610 41.000 158.930 ;
        RECT 38.720 157.395 40.260 157.765 ;
        RECT 40.800 156.550 40.940 158.610 ;
        RECT 40.740 156.230 41.000 156.550 ;
        RECT 41.260 156.210 41.400 162.350 ;
        RECT 41.660 158.610 41.920 158.930 ;
        RECT 42.120 158.610 42.380 158.930 ;
        RECT 42.580 158.610 42.840 158.930 ;
        RECT 41.720 156.890 41.860 158.610 ;
        RECT 41.660 156.570 41.920 156.890 ;
        RECT 41.200 155.890 41.460 156.210 ;
        RECT 38.900 155.210 39.160 155.530 ;
        RECT 38.440 154.080 38.700 154.170 ;
        RECT 38.040 153.940 38.700 154.080 ;
        RECT 38.040 151.110 38.180 153.940 ;
        RECT 38.440 153.850 38.700 153.940 ;
        RECT 38.960 153.830 39.100 155.210 ;
        RECT 42.180 154.510 42.320 158.610 ;
        RECT 42.640 157.230 42.780 158.610 ;
        RECT 42.580 156.910 42.840 157.230 ;
        RECT 42.120 154.190 42.380 154.510 ;
        RECT 38.900 153.510 39.160 153.830 ;
        RECT 42.120 153.170 42.380 153.490 ;
        RECT 41.200 152.830 41.460 153.150 ;
        RECT 38.720 151.955 40.260 152.325 ;
        RECT 41.260 151.790 41.400 152.830 ;
        RECT 42.180 151.790 42.320 153.170 ;
        RECT 41.200 151.470 41.460 151.790 ;
        RECT 42.120 151.470 42.380 151.790 ;
        RECT 37.980 150.790 38.240 151.110 ;
        RECT 43.100 150.770 43.240 167.450 ;
        RECT 45.800 167.110 46.060 167.430 ;
        RECT 44.880 166.770 45.140 167.090 ;
        RECT 44.940 165.390 45.080 166.770 ;
        RECT 45.860 165.390 46.000 167.110 ;
        RECT 46.320 167.090 46.460 167.790 ;
        RECT 46.780 167.430 46.920 173.230 ;
        RECT 47.240 172.870 47.380 174.590 ;
        RECT 47.180 172.550 47.440 172.870 ;
        RECT 46.720 167.110 46.980 167.430 ;
        RECT 46.260 166.770 46.520 167.090 ;
        RECT 44.880 165.070 45.140 165.390 ;
        RECT 45.800 165.070 46.060 165.390 ;
        RECT 43.960 164.390 44.220 164.710 ;
        RECT 45.340 164.390 45.600 164.710 ;
        RECT 43.500 160.650 43.760 160.970 ;
        RECT 43.560 153.830 43.700 160.650 ;
        RECT 44.020 159.610 44.160 164.390 ;
        RECT 44.420 160.650 44.680 160.970 ;
        RECT 43.960 159.290 44.220 159.610 ;
        RECT 44.480 158.590 44.620 160.650 ;
        RECT 44.420 158.270 44.680 158.590 ;
        RECT 44.420 155.890 44.680 156.210 ;
        RECT 43.500 153.510 43.760 153.830 ;
        RECT 44.480 153.490 44.620 155.890 ;
        RECT 45.400 153.830 45.540 164.390 ;
        RECT 46.720 164.225 46.980 164.370 ;
        RECT 46.710 163.855 46.990 164.225 ;
        RECT 47.700 164.030 47.840 176.210 ;
        RECT 49.540 170.150 49.680 185.615 ;
        RECT 49.480 170.060 49.740 170.150 ;
        RECT 49.080 169.920 49.740 170.060 ;
        RECT 48.100 166.770 48.360 167.090 ;
        RECT 46.260 159.290 46.520 159.610 ;
        RECT 46.320 157.230 46.460 159.290 ;
        RECT 46.780 158.250 46.920 163.855 ;
        RECT 47.640 163.710 47.900 164.030 ;
        RECT 47.180 163.370 47.440 163.690 ;
        RECT 47.240 159.270 47.380 163.370 ;
        RECT 47.700 162.330 47.840 163.710 ;
        RECT 47.640 162.010 47.900 162.330 ;
        RECT 47.640 160.650 47.900 160.970 ;
        RECT 47.180 158.950 47.440 159.270 ;
        RECT 46.720 157.930 46.980 158.250 ;
        RECT 46.260 156.910 46.520 157.230 ;
        RECT 47.240 156.550 47.380 158.950 ;
        RECT 47.180 156.230 47.440 156.550 ;
        RECT 47.700 155.870 47.840 160.650 ;
        RECT 48.160 159.350 48.300 166.770 ;
        RECT 48.560 166.090 48.820 166.410 ;
        RECT 48.620 159.860 48.760 166.090 ;
        RECT 49.080 160.710 49.220 169.920 ;
        RECT 49.480 169.830 49.740 169.920 ;
        RECT 49.480 166.430 49.740 166.750 ;
        RECT 49.540 162.670 49.680 166.430 ;
        RECT 49.480 162.350 49.740 162.670 ;
        RECT 49.080 160.570 49.680 160.710 ;
        RECT 48.620 159.720 49.220 159.860 ;
        RECT 48.160 159.210 48.760 159.350 ;
        RECT 48.620 158.930 48.760 159.210 ;
        RECT 48.560 158.610 48.820 158.930 ;
        RECT 48.620 156.210 48.760 158.610 ;
        RECT 48.560 155.890 48.820 156.210 ;
        RECT 47.640 155.550 47.900 155.870 ;
        RECT 45.340 153.510 45.600 153.830 ;
        RECT 44.420 153.170 44.680 153.490 ;
        RECT 43.040 150.450 43.300 150.770 ;
        RECT 43.040 149.770 43.300 150.090 ;
        RECT 38.720 146.515 40.260 146.885 ;
        RECT 42.580 145.010 42.840 145.330 ;
        RECT 42.640 143.630 42.780 145.010 ;
        RECT 42.580 143.310 42.840 143.630 ;
        RECT 42.580 142.630 42.840 142.950 ;
        RECT 40.740 142.290 41.000 142.610 ;
        RECT 38.720 141.075 40.260 141.445 ;
        RECT 40.800 139.210 40.940 142.290 ;
        RECT 41.660 141.610 41.920 141.930 ;
        RECT 41.720 139.890 41.860 141.610 ;
        RECT 41.660 139.570 41.920 139.890 ;
        RECT 40.740 138.890 41.000 139.210 ;
        RECT 40.800 136.490 40.940 138.890 ;
        RECT 41.660 137.870 41.920 138.190 ;
        RECT 40.740 136.170 41.000 136.490 ;
        RECT 38.720 135.635 40.260 136.005 ;
        RECT 41.720 135.470 41.860 137.870 ;
        RECT 42.640 136.490 42.780 142.630 ;
        RECT 42.580 136.170 42.840 136.490 ;
        RECT 41.660 135.150 41.920 135.470 ;
        RECT 43.100 134.450 43.240 149.770 ;
        RECT 44.880 147.050 45.140 147.370 ;
        RECT 44.940 145.330 45.080 147.050 ;
        RECT 45.400 146.350 45.540 153.510 ;
        RECT 48.620 153.490 48.760 155.890 ;
        RECT 48.560 153.170 48.820 153.490 ;
        RECT 48.100 152.490 48.360 152.810 ;
        RECT 48.160 151.110 48.300 152.490 ;
        RECT 48.100 150.790 48.360 151.110 ;
        RECT 48.100 150.340 48.360 150.430 ;
        RECT 47.240 150.200 48.360 150.340 ;
        RECT 45.340 146.030 45.600 146.350 ;
        RECT 46.260 145.350 46.520 145.670 ;
        RECT 44.880 145.010 45.140 145.330 ;
        RECT 43.960 144.670 44.220 144.990 ;
        RECT 44.020 143.630 44.160 144.670 ;
        RECT 43.960 143.310 44.220 143.630 ;
        RECT 45.800 142.630 46.060 142.950 ;
        RECT 45.860 140.910 46.000 142.630 ;
        RECT 46.320 140.910 46.460 145.350 ;
        RECT 47.240 144.650 47.380 150.200 ;
        RECT 48.100 150.110 48.360 150.200 ;
        RECT 48.620 148.390 48.760 153.170 ;
        RECT 49.080 151.450 49.220 159.720 ;
        RECT 49.020 151.130 49.280 151.450 ;
        RECT 49.020 150.450 49.280 150.770 ;
        RECT 49.080 149.070 49.220 150.450 ;
        RECT 49.540 150.090 49.680 160.570 ;
        RECT 49.480 149.770 49.740 150.090 ;
        RECT 49.020 148.750 49.280 149.070 ;
        RECT 50.000 148.980 50.140 202.470 ;
        RECT 50.460 199.730 50.600 204.170 ;
        RECT 51.380 202.790 51.520 206.890 ;
        RECT 51.840 204.490 51.980 207.230 ;
        RECT 54.140 205.590 54.280 207.490 ;
        RECT 54.540 206.890 54.800 207.210 ;
        RECT 52.240 205.190 52.500 205.510 ;
        RECT 53.220 205.450 54.280 205.590 ;
        RECT 51.780 204.170 52.040 204.490 ;
        RECT 51.320 202.470 51.580 202.790 ;
        RECT 51.840 200.410 51.980 204.170 ;
        RECT 51.780 200.090 52.040 200.410 ;
        RECT 50.400 199.410 50.660 199.730 ;
        RECT 52.300 197.010 52.440 205.190 ;
        RECT 52.700 202.470 52.960 202.790 ;
        RECT 52.240 196.690 52.500 197.010 ;
        RECT 50.400 194.990 50.660 195.310 ;
        RECT 50.460 192.590 50.600 194.990 ;
        RECT 50.860 193.630 51.120 193.950 ;
        RECT 50.400 192.270 50.660 192.590 ;
        RECT 50.460 188.850 50.600 192.270 ;
        RECT 50.920 191.910 51.060 193.630 ;
        RECT 50.860 191.820 51.120 191.910 ;
        RECT 50.860 191.680 51.520 191.820 ;
        RECT 50.860 191.590 51.120 191.680 ;
        RECT 50.860 190.570 51.120 190.890 ;
        RECT 50.400 188.530 50.660 188.850 ;
        RECT 50.400 187.850 50.660 188.170 ;
        RECT 50.460 186.470 50.600 187.850 ;
        RECT 50.920 187.150 51.060 190.570 ;
        RECT 51.380 188.170 51.520 191.680 ;
        RECT 51.780 188.870 52.040 189.190 ;
        RECT 51.320 187.850 51.580 188.170 ;
        RECT 50.860 186.830 51.120 187.150 ;
        RECT 50.920 186.470 51.060 186.830 ;
        RECT 50.400 186.150 50.660 186.470 ;
        RECT 50.860 186.150 51.120 186.470 ;
        RECT 51.840 186.380 51.980 188.870 ;
        RECT 52.300 186.470 52.440 196.690 ;
        RECT 51.380 186.240 51.980 186.380 ;
        RECT 51.380 183.410 51.520 186.240 ;
        RECT 52.240 186.150 52.500 186.470 ;
        RECT 51.780 185.470 52.040 185.790 ;
        RECT 51.320 183.090 51.580 183.410 ;
        RECT 50.860 177.310 51.120 177.630 ;
        RECT 50.920 176.270 51.060 177.310 ;
        RECT 51.320 176.970 51.580 177.290 ;
        RECT 51.380 176.270 51.520 176.970 ;
        RECT 50.860 175.950 51.120 176.270 ;
        RECT 51.320 175.950 51.580 176.270 ;
        RECT 50.400 170.170 50.660 170.490 ;
        RECT 50.460 161.650 50.600 170.170 ;
        RECT 50.850 169.975 51.130 170.345 ;
        RECT 50.860 169.830 51.120 169.975 ;
        RECT 51.320 169.490 51.580 169.810 ;
        RECT 50.860 164.050 51.120 164.370 ;
        RECT 50.400 161.330 50.660 161.650 ;
        RECT 50.920 159.270 51.060 164.050 ;
        RECT 51.380 161.650 51.520 169.490 ;
        RECT 51.840 167.090 51.980 185.470 ;
        RECT 52.240 171.870 52.500 172.190 ;
        RECT 52.300 170.830 52.440 171.870 ;
        RECT 52.240 170.510 52.500 170.830 ;
        RECT 51.780 166.770 52.040 167.090 ;
        RECT 52.760 164.690 52.900 202.470 ;
        RECT 53.220 199.390 53.360 205.450 ;
        RECT 54.600 205.170 54.740 206.890 ;
        RECT 60.120 206.190 60.260 207.570 ;
        RECT 63.740 207.230 64.000 207.550 ;
        RECT 60.060 205.870 60.320 206.190 ;
        RECT 54.540 204.850 54.800 205.170 ;
        RECT 55.510 203.635 57.050 204.005 ;
        RECT 55.000 202.470 55.260 202.790 ;
        RECT 54.080 202.130 54.340 202.450 ;
        RECT 53.160 199.070 53.420 199.390 ;
        RECT 53.220 196.330 53.360 199.070 ;
        RECT 54.140 198.030 54.280 202.130 ;
        RECT 55.060 200.750 55.200 202.470 ;
        RECT 55.000 200.430 55.260 200.750 ;
        RECT 55.510 198.195 57.050 198.565 ;
        RECT 54.080 197.710 54.340 198.030 ;
        RECT 53.620 197.030 53.880 197.350 ;
        RECT 53.160 196.010 53.420 196.330 ;
        RECT 53.220 193.950 53.360 196.010 ;
        RECT 53.680 195.310 53.820 197.030 ;
        RECT 53.620 194.990 53.880 195.310 ;
        RECT 54.140 194.290 54.280 197.710 ;
        RECT 59.140 197.030 59.400 197.350 ;
        RECT 57.300 196.350 57.560 196.670 ;
        RECT 57.360 194.290 57.500 196.350 ;
        RECT 59.200 196.330 59.340 197.030 ;
        RECT 60.120 197.010 60.260 205.870 ;
        RECT 62.360 205.190 62.620 205.510 ;
        RECT 61.440 204.850 61.700 205.170 ;
        RECT 61.500 199.390 61.640 204.850 ;
        RECT 61.900 201.680 62.160 201.770 ;
        RECT 62.420 201.680 62.560 205.190 ;
        RECT 62.820 204.170 63.080 204.490 ;
        RECT 63.280 204.170 63.540 204.490 ;
        RECT 61.900 201.540 62.560 201.680 ;
        RECT 61.900 201.450 62.160 201.540 ;
        RECT 61.440 199.070 61.700 199.390 ;
        RECT 60.520 197.370 60.780 197.690 ;
        RECT 60.060 196.690 60.320 197.010 ;
        RECT 59.140 196.010 59.400 196.330 ;
        RECT 59.200 194.290 59.340 196.010 ;
        RECT 54.080 193.970 54.340 194.290 ;
        RECT 57.300 193.970 57.560 194.290 ;
        RECT 59.140 193.970 59.400 194.290 ;
        RECT 53.160 193.630 53.420 193.950 ;
        RECT 53.220 171.025 53.360 193.630 ;
        RECT 53.620 193.290 53.880 193.610 ;
        RECT 53.680 185.985 53.820 193.290 ;
        RECT 54.140 192.250 54.280 193.970 ;
        RECT 60.120 193.950 60.260 196.690 ;
        RECT 60.580 195.310 60.720 197.370 ;
        RECT 61.500 196.670 61.640 199.070 ;
        RECT 61.440 196.350 61.700 196.670 ;
        RECT 61.960 196.070 62.100 201.450 ;
        RECT 62.880 200.750 63.020 204.170 ;
        RECT 63.340 202.790 63.480 204.170 ;
        RECT 63.280 202.470 63.540 202.790 ;
        RECT 62.820 200.430 63.080 200.750 ;
        RECT 63.800 199.050 63.940 207.230 ;
        RECT 68.340 206.890 68.600 207.210 ;
        RECT 68.400 205.590 68.540 206.890 ;
        RECT 67.020 205.450 68.540 205.590 ;
        RECT 67.020 205.170 67.160 205.450 ;
        RECT 64.200 204.850 64.460 205.170 ;
        RECT 65.580 204.850 65.840 205.170 ;
        RECT 66.960 204.850 67.220 205.170 ;
        RECT 64.260 200.410 64.400 204.850 ;
        RECT 65.640 203.470 65.780 204.850 ;
        RECT 66.500 204.170 66.760 204.490 ;
        RECT 65.580 203.150 65.840 203.470 ;
        RECT 64.660 202.810 64.920 203.130 ;
        RECT 64.200 200.090 64.460 200.410 ;
        RECT 62.820 198.730 63.080 199.050 ;
        RECT 63.740 198.730 64.000 199.050 ;
        RECT 62.880 197.690 63.020 198.730 ;
        RECT 62.820 197.370 63.080 197.690 ;
        RECT 62.360 196.350 62.620 196.670 ;
        RECT 62.420 196.070 62.560 196.350 ;
        RECT 61.960 195.930 62.560 196.070 ;
        RECT 60.520 194.990 60.780 195.310 ;
        RECT 61.960 194.290 62.100 195.930 ;
        RECT 61.900 193.970 62.160 194.290 ;
        RECT 60.060 193.630 60.320 193.950 ;
        RECT 55.510 192.755 57.050 193.125 ;
        RECT 60.120 192.590 60.260 193.630 ;
        RECT 54.540 192.270 54.800 192.590 ;
        RECT 60.060 192.270 60.320 192.590 ;
        RECT 54.080 191.930 54.340 192.250 ;
        RECT 54.600 189.190 54.740 192.270 ;
        RECT 55.000 191.590 55.260 191.910 ;
        RECT 54.540 188.870 54.800 189.190 ;
        RECT 54.540 188.190 54.800 188.510 ;
        RECT 54.080 187.850 54.340 188.170 ;
        RECT 53.610 185.615 53.890 185.985 ;
        RECT 54.140 185.450 54.280 187.850 ;
        RECT 54.080 185.130 54.340 185.450 ;
        RECT 54.600 183.750 54.740 188.190 ;
        RECT 55.060 184.430 55.200 191.590 ;
        RECT 61.960 191.570 62.100 193.970 ;
        RECT 62.360 193.630 62.620 193.950 ;
        RECT 62.420 191.570 62.560 193.630 ;
        RECT 62.880 193.610 63.020 197.370 ;
        RECT 64.720 193.950 64.860 202.810 ;
        RECT 66.560 199.730 66.700 204.170 ;
        RECT 70.700 203.470 70.840 208.250 ;
        RECT 71.160 208.230 71.300 212.220 ;
        RECT 78.520 208.230 78.660 212.220 ;
        RECT 71.100 207.910 71.360 208.230 ;
        RECT 78.460 207.910 78.720 208.230 ;
        RECT 80.300 207.910 80.560 208.230 ;
        RECT 76.160 207.230 76.420 207.550 ;
        RECT 71.560 206.890 71.820 207.210 ;
        RECT 75.240 206.890 75.500 207.210 ;
        RECT 71.620 203.470 71.760 206.890 ;
        RECT 72.300 206.355 73.840 206.725 ;
        RECT 75.300 205.170 75.440 206.890 ;
        RECT 76.220 205.170 76.360 207.230 ;
        RECT 78.460 206.890 78.720 207.210 ;
        RECT 76.620 205.190 76.880 205.510 ;
        RECT 75.240 204.850 75.500 205.170 ;
        RECT 76.160 204.850 76.420 205.170 ;
        RECT 72.940 204.170 73.200 204.490 ;
        RECT 74.320 204.170 74.580 204.490 ;
        RECT 70.640 203.150 70.900 203.470 ;
        RECT 71.560 203.150 71.820 203.470 ;
        RECT 70.180 202.130 70.440 202.450 ;
        RECT 70.240 200.410 70.380 202.130 ;
        RECT 70.180 200.090 70.440 200.410 ;
        RECT 66.500 199.410 66.760 199.730 ;
        RECT 69.720 199.410 69.980 199.730 ;
        RECT 66.560 196.750 66.700 199.410 ;
        RECT 66.960 198.730 67.220 199.050 ;
        RECT 67.020 197.690 67.160 198.730 ;
        RECT 66.960 197.370 67.220 197.690 ;
        RECT 68.800 197.030 69.060 197.350 ;
        RECT 66.560 196.610 67.160 196.750 ;
        RECT 64.660 193.630 64.920 193.950 ;
        RECT 62.820 193.290 63.080 193.610 ;
        RECT 61.900 191.250 62.160 191.570 ;
        RECT 62.360 191.250 62.620 191.570 ;
        RECT 60.520 188.530 60.780 188.850 ;
        RECT 57.300 187.850 57.560 188.170 ;
        RECT 55.510 187.315 57.050 187.685 ;
        RECT 55.000 184.110 55.260 184.430 ;
        RECT 54.540 183.430 54.800 183.750 ;
        RECT 54.600 181.370 54.740 183.430 ;
        RECT 57.360 183.410 57.500 187.850 ;
        RECT 60.580 187.150 60.720 188.530 ;
        RECT 60.520 186.830 60.780 187.150 ;
        RECT 61.440 186.150 61.700 186.470 ;
        RECT 61.500 183.410 61.640 186.150 ;
        RECT 61.960 183.410 62.100 191.250 ;
        RECT 62.420 188.850 62.560 191.250 ;
        RECT 66.500 190.910 66.760 191.230 ;
        RECT 65.120 190.570 65.380 190.890 ;
        RECT 65.580 190.570 65.840 190.890 ;
        RECT 62.360 188.530 62.620 188.850 ;
        RECT 65.180 188.760 65.320 190.570 ;
        RECT 65.640 189.530 65.780 190.570 ;
        RECT 66.560 189.870 66.700 190.910 ;
        RECT 66.500 189.550 66.760 189.870 ;
        RECT 65.580 189.210 65.840 189.530 ;
        RECT 65.580 188.760 65.840 188.850 ;
        RECT 65.180 188.620 65.840 188.760 ;
        RECT 65.580 188.530 65.840 188.620 ;
        RECT 67.020 188.510 67.160 196.610 ;
        RECT 68.860 191.570 69.000 197.030 ;
        RECT 69.780 195.310 69.920 199.410 ;
        RECT 69.720 194.990 69.980 195.310 ;
        RECT 70.240 194.290 70.380 200.090 ;
        RECT 71.620 200.070 71.760 203.150 ;
        RECT 73.000 202.790 73.140 204.170 ;
        RECT 72.940 202.470 73.200 202.790 ;
        RECT 72.300 200.915 73.840 201.285 ;
        RECT 71.560 199.750 71.820 200.070 ;
        RECT 71.100 199.410 71.360 199.730 ;
        RECT 70.640 198.730 70.900 199.050 ;
        RECT 70.700 195.310 70.840 198.730 ;
        RECT 71.160 197.010 71.300 199.410 ;
        RECT 71.620 198.030 71.760 199.750 ;
        RECT 71.560 197.710 71.820 198.030 ;
        RECT 71.100 196.690 71.360 197.010 ;
        RECT 71.160 196.330 71.300 196.690 ;
        RECT 71.560 196.350 71.820 196.670 ;
        RECT 71.100 196.010 71.360 196.330 ;
        RECT 70.640 194.990 70.900 195.310 ;
        RECT 71.620 194.630 71.760 196.350 ;
        RECT 72.300 195.475 73.840 195.845 ;
        RECT 71.560 194.310 71.820 194.630 ;
        RECT 74.380 194.290 74.520 204.170 ;
        RECT 75.300 203.470 75.440 204.850 ;
        RECT 75.240 203.150 75.500 203.470 ;
        RECT 76.220 203.130 76.360 204.850 ;
        RECT 76.160 202.810 76.420 203.130 ;
        RECT 76.680 199.470 76.820 205.190 ;
        RECT 77.080 204.510 77.340 204.830 ;
        RECT 77.140 200.750 77.280 204.510 ;
        RECT 77.080 200.430 77.340 200.750 ;
        RECT 78.520 199.730 78.660 206.890 ;
        RECT 80.360 206.190 80.500 207.910 ;
        RECT 83.520 207.570 83.780 207.890 ;
        RECT 83.580 206.190 83.720 207.570 ;
        RECT 80.300 205.870 80.560 206.190 ;
        RECT 83.520 205.870 83.780 206.190 ;
        RECT 83.580 203.470 83.720 205.870 ;
        RECT 85.880 205.170 86.020 212.220 ;
        RECT 89.090 209.075 90.630 209.445 ;
        RECT 93.240 208.230 93.380 212.220 ;
        RECT 100.600 208.570 100.740 212.220 ;
        RECT 107.960 211.710 108.100 212.220 ;
        RECT 108.420 211.710 108.560 212.250 ;
        RECT 107.960 211.570 108.560 211.710 ;
        RECT 103.300 209.610 103.560 209.930 ;
        RECT 100.540 208.250 100.800 208.570 ;
        RECT 103.360 208.230 103.500 209.610 ;
        RECT 109.800 208.570 109.940 212.250 ;
        RECT 115.250 212.220 115.530 213.700 ;
        RECT 115.780 212.250 116.840 212.390 ;
        RECT 115.320 211.710 115.460 212.220 ;
        RECT 115.780 211.710 115.920 212.250 ;
        RECT 115.320 211.570 115.920 211.710 ;
        RECT 116.700 208.570 116.840 212.250 ;
        RECT 122.610 212.220 122.890 213.700 ;
        RECT 123.140 212.250 124.660 212.390 ;
        RECT 122.680 211.710 122.820 212.220 ;
        RECT 123.140 211.710 123.280 212.250 ;
        RECT 122.680 211.570 123.280 211.710 ;
        RECT 117.100 209.610 117.360 209.930 ;
        RECT 117.160 208.910 117.300 209.610 ;
        RECT 122.670 209.075 124.210 209.445 ;
        RECT 117.100 208.590 117.360 208.910 ;
        RECT 124.520 208.570 124.660 212.250 ;
        RECT 129.970 212.220 130.250 213.700 ;
        RECT 137.330 212.220 137.610 213.700 ;
        RECT 144.690 212.220 144.970 213.700 ;
        RECT 152.050 212.220 152.330 213.700 ;
        RECT 130.040 208.990 130.180 212.220 ;
        RECT 130.040 208.850 130.640 208.990 ;
        RECT 130.500 208.570 130.640 208.850 ;
        RECT 90.880 207.910 91.140 208.230 ;
        RECT 93.180 207.910 93.440 208.230 ;
        RECT 103.300 207.910 103.560 208.230 ;
        RECT 108.350 208.055 108.630 208.425 ;
        RECT 109.740 208.250 110.000 208.570 ;
        RECT 108.360 207.910 108.620 208.055 ;
        RECT 108.820 207.910 109.080 208.230 ;
        RECT 110.200 207.910 110.460 208.230 ;
        RECT 113.880 207.910 114.140 208.230 ;
        RECT 115.250 208.140 115.530 208.425 ;
        RECT 115.720 208.250 115.980 208.570 ;
        RECT 116.640 208.250 116.900 208.570 ;
        RECT 124.460 208.250 124.720 208.570 ;
        RECT 130.440 208.250 130.700 208.570 ;
        RECT 114.860 208.055 115.530 208.140 ;
        RECT 114.860 208.000 115.520 208.055 ;
        RECT 88.120 206.890 88.380 207.210 ;
        RECT 89.960 206.890 90.220 207.210 ;
        RECT 85.820 204.850 86.080 205.170 ;
        RECT 85.820 204.170 86.080 204.490 ;
        RECT 87.660 204.170 87.920 204.490 ;
        RECT 83.520 203.150 83.780 203.470 ;
        RECT 82.600 202.130 82.860 202.450 ;
        RECT 83.060 202.130 83.320 202.450 ;
        RECT 81.220 201.450 81.480 201.770 ;
        RECT 74.780 199.070 75.040 199.390 ;
        RECT 75.700 199.070 75.960 199.390 ;
        RECT 76.680 199.330 77.280 199.470 ;
        RECT 78.460 199.410 78.720 199.730 ;
        RECT 74.840 196.670 74.980 199.070 ;
        RECT 74.780 196.350 75.040 196.670 ;
        RECT 74.840 194.970 74.980 196.350 ;
        RECT 75.240 196.010 75.500 196.330 ;
        RECT 74.780 194.650 75.040 194.970 ;
        RECT 70.180 193.970 70.440 194.290 ;
        RECT 74.320 193.970 74.580 194.290 ;
        RECT 71.560 193.630 71.820 193.950 ;
        RECT 68.800 191.250 69.060 191.570 ;
        RECT 69.260 190.570 69.520 190.890 ;
        RECT 68.800 188.530 69.060 188.850 ;
        RECT 66.960 188.190 67.220 188.510 ;
        RECT 66.040 186.150 66.300 186.470 ;
        RECT 62.820 185.130 63.080 185.450 ;
        RECT 63.280 185.130 63.540 185.450 ;
        RECT 62.880 184.430 63.020 185.130 ;
        RECT 62.820 184.110 63.080 184.430 ;
        RECT 63.340 183.410 63.480 185.130 ;
        RECT 55.000 183.090 55.260 183.410 ;
        RECT 57.300 183.090 57.560 183.410 ;
        RECT 61.440 183.090 61.700 183.410 ;
        RECT 61.900 183.090 62.160 183.410 ;
        RECT 63.280 183.090 63.540 183.410 ;
        RECT 54.540 181.050 54.800 181.370 ;
        RECT 54.600 180.690 54.740 181.050 ;
        RECT 55.060 181.030 55.200 183.090 ;
        RECT 59.140 182.750 59.400 183.070 ;
        RECT 55.510 181.875 57.050 182.245 ;
        RECT 59.200 181.710 59.340 182.750 ;
        RECT 59.600 182.410 59.860 182.730 ;
        RECT 59.140 181.390 59.400 181.710 ;
        RECT 55.000 180.710 55.260 181.030 ;
        RECT 58.220 180.710 58.480 181.030 ;
        RECT 54.540 180.370 54.800 180.690 ;
        RECT 53.620 176.970 53.880 177.290 ;
        RECT 53.680 175.590 53.820 176.970 ;
        RECT 54.600 175.930 54.740 180.370 ;
        RECT 54.540 175.610 54.800 175.930 ;
        RECT 53.620 175.270 53.880 175.590 ;
        RECT 54.080 175.270 54.340 175.590 ;
        RECT 54.140 173.550 54.280 175.270 ;
        RECT 54.080 173.230 54.340 173.550 ;
        RECT 53.150 170.655 53.430 171.025 ;
        RECT 54.600 170.490 54.740 175.610 ;
        RECT 55.060 174.910 55.200 180.710 ;
        RECT 57.760 179.690 58.020 180.010 ;
        RECT 57.300 177.650 57.560 177.970 ;
        RECT 55.510 176.435 57.050 176.805 ;
        RECT 55.920 175.270 56.180 175.590 ;
        RECT 55.980 174.910 56.120 175.270 ;
        RECT 57.360 175.250 57.500 177.650 ;
        RECT 57.820 175.930 57.960 179.690 ;
        RECT 57.760 175.610 58.020 175.930 ;
        RECT 56.840 174.930 57.100 175.250 ;
        RECT 57.300 174.930 57.560 175.250 ;
        RECT 55.000 174.590 55.260 174.910 ;
        RECT 55.920 174.590 56.180 174.910 ;
        RECT 55.980 173.210 56.120 174.590 ;
        RECT 55.920 172.890 56.180 173.210 ;
        RECT 56.900 171.850 57.040 174.930 ;
        RECT 57.760 172.890 58.020 173.210 ;
        RECT 55.000 171.530 55.260 171.850 ;
        RECT 56.840 171.530 57.100 171.850 ;
        RECT 54.540 170.170 54.800 170.490 ;
        RECT 55.060 170.150 55.200 171.530 ;
        RECT 55.510 170.995 57.050 171.365 ;
        RECT 57.820 170.830 57.960 172.890 ;
        RECT 57.760 170.510 58.020 170.830 ;
        RECT 57.820 170.150 57.960 170.510 ;
        RECT 53.620 170.060 53.880 170.150 ;
        RECT 53.220 169.920 53.880 170.060 ;
        RECT 53.220 169.470 53.360 169.920 ;
        RECT 53.620 169.830 53.880 169.920 ;
        RECT 55.000 169.830 55.260 170.150 ;
        RECT 55.460 169.830 55.720 170.150 ;
        RECT 57.760 169.830 58.020 170.150 ;
        RECT 53.160 169.150 53.420 169.470 ;
        RECT 51.840 164.550 52.900 164.690 ;
        RECT 51.320 161.330 51.580 161.650 ;
        RECT 50.860 158.950 51.120 159.270 ;
        RECT 51.840 149.830 51.980 164.550 ;
        RECT 52.240 163.370 52.500 163.690 ;
        RECT 52.300 161.650 52.440 163.370 ;
        RECT 52.240 161.330 52.500 161.650 ;
        RECT 49.540 148.840 50.140 148.980 ;
        RECT 50.920 149.690 51.980 149.830 ;
        RECT 52.240 149.770 52.500 150.090 ;
        RECT 48.560 148.070 48.820 148.390 ;
        RECT 48.100 145.350 48.360 145.670 ;
        RECT 47.640 145.010 47.900 145.330 ;
        RECT 47.180 144.330 47.440 144.650 ;
        RECT 45.800 140.590 46.060 140.910 ;
        RECT 46.260 140.590 46.520 140.910 ;
        RECT 44.420 139.570 44.680 139.890 ;
        RECT 44.880 139.570 45.140 139.890 ;
        RECT 44.480 136.830 44.620 139.570 ;
        RECT 44.940 138.190 45.080 139.570 ;
        RECT 44.880 137.870 45.140 138.190 ;
        RECT 46.320 137.510 46.460 140.590 ;
        RECT 47.240 140.570 47.380 144.330 ;
        RECT 47.700 143.290 47.840 145.010 ;
        RECT 47.640 142.970 47.900 143.290 ;
        RECT 48.160 142.350 48.300 145.350 ;
        RECT 47.700 142.210 48.300 142.350 ;
        RECT 47.700 141.930 47.840 142.210 ;
        RECT 47.640 141.610 47.900 141.930 ;
        RECT 48.100 141.610 48.360 141.930 ;
        RECT 47.180 140.250 47.440 140.570 ;
        RECT 46.720 139.910 46.980 140.230 ;
        RECT 46.780 139.210 46.920 139.910 ;
        RECT 48.160 139.890 48.300 141.610 ;
        RECT 48.100 139.570 48.360 139.890 ;
        RECT 46.720 138.890 46.980 139.210 ;
        RECT 47.180 138.890 47.440 139.210 ;
        RECT 47.240 138.190 47.380 138.890 ;
        RECT 47.180 137.870 47.440 138.190 ;
        RECT 46.260 137.190 46.520 137.510 ;
        RECT 44.420 136.510 44.680 136.830 ;
        RECT 49.020 134.470 49.280 134.790 ;
        RECT 43.040 134.360 43.300 134.450 ;
        RECT 43.040 134.220 43.700 134.360 ;
        RECT 43.040 134.130 43.300 134.220 ;
        RECT 40.740 133.790 41.000 134.110 ;
        RECT 37.980 132.090 38.240 132.410 ;
        RECT 38.040 130.030 38.180 132.090 ;
        RECT 38.720 130.195 40.260 130.565 ;
        RECT 37.980 129.710 38.240 130.030 ;
        RECT 40.800 129.350 40.940 133.790 ;
        RECT 43.040 133.450 43.300 133.770 ;
        RECT 42.580 130.730 42.840 131.050 ;
        RECT 40.740 129.030 41.000 129.350 ;
        RECT 42.640 129.010 42.780 130.730 ;
        RECT 43.100 129.350 43.240 133.450 ;
        RECT 43.560 129.350 43.700 134.220 ;
        RECT 43.960 134.130 44.220 134.450 ;
        RECT 44.020 131.050 44.160 134.130 ;
        RECT 45.340 131.750 45.600 132.070 ;
        RECT 43.960 130.730 44.220 131.050 ;
        RECT 43.040 129.030 43.300 129.350 ;
        RECT 43.500 129.030 43.760 129.350 ;
        RECT 42.580 128.690 42.840 129.010 ;
        RECT 42.640 126.290 42.780 128.690 ;
        RECT 44.020 126.630 44.160 130.730 ;
        RECT 45.400 126.970 45.540 131.750 ;
        RECT 49.080 131.050 49.220 134.470 ;
        RECT 45.800 130.730 46.060 131.050 ;
        RECT 49.020 130.730 49.280 131.050 ;
        RECT 45.860 128.670 46.000 130.730 ;
        RECT 45.800 128.350 46.060 128.670 ;
        RECT 45.340 126.650 45.600 126.970 ;
        RECT 49.080 126.710 49.220 130.730 ;
        RECT 47.240 126.630 49.220 126.710 ;
        RECT 43.960 126.310 44.220 126.630 ;
        RECT 47.180 126.570 49.220 126.630 ;
        RECT 47.180 126.310 47.440 126.570 ;
        RECT 42.580 125.970 42.840 126.290 ;
        RECT 38.720 124.755 40.260 125.125 ;
        RECT 42.640 123.570 42.780 125.970 ;
        RECT 42.580 123.250 42.840 123.570 ;
        RECT 45.800 123.250 46.060 123.570 ;
        RECT 47.180 123.250 47.440 123.570 ;
        RECT 40.740 122.910 41.000 123.230 ;
        RECT 39.360 122.570 39.620 122.890 ;
        RECT 39.420 121.190 39.560 122.570 ;
        RECT 40.800 121.870 40.940 122.910 ;
        RECT 40.740 121.550 41.000 121.870 ;
        RECT 39.360 120.870 39.620 121.190 ;
        RECT 42.640 120.170 42.780 123.250 ;
        RECT 43.500 122.910 43.760 123.230 ;
        RECT 43.040 122.570 43.300 122.890 ;
        RECT 42.580 119.850 42.840 120.170 ;
        RECT 38.720 119.315 40.260 119.685 ;
        RECT 42.580 118.830 42.840 119.150 ;
        RECT 38.440 118.490 38.700 118.810 ;
        RECT 37.980 117.470 38.240 117.790 ;
        RECT 38.040 115.750 38.180 117.470 ;
        RECT 38.500 116.430 38.640 118.490 ;
        RECT 42.640 118.470 42.780 118.830 ;
        RECT 42.580 118.150 42.840 118.470 ;
        RECT 41.660 117.810 41.920 118.130 ;
        RECT 41.200 117.130 41.460 117.450 ;
        RECT 38.440 116.110 38.700 116.430 ;
        RECT 37.980 115.430 38.240 115.750 ;
        RECT 38.500 115.150 38.640 116.110 ;
        RECT 41.260 115.750 41.400 117.130 ;
        RECT 41.720 116.430 41.860 117.810 ;
        RECT 41.660 116.110 41.920 116.430 ;
        RECT 41.200 115.430 41.460 115.750 ;
        RECT 38.040 115.010 38.640 115.150 ;
        RECT 38.040 113.710 38.180 115.010 ;
        RECT 40.740 114.410 41.000 114.730 ;
        RECT 38.720 113.875 40.260 114.245 ;
        RECT 37.980 113.390 38.240 113.710 ;
        RECT 40.800 112.430 40.940 114.410 ;
        RECT 41.720 113.710 41.860 116.110 ;
        RECT 43.100 115.750 43.240 122.570 ;
        RECT 43.560 118.130 43.700 122.910 ;
        RECT 45.860 119.150 46.000 123.250 ;
        RECT 46.720 120.190 46.980 120.510 ;
        RECT 45.800 118.830 46.060 119.150 ;
        RECT 43.500 117.810 43.760 118.130 ;
        RECT 43.040 115.430 43.300 115.750 ;
        RECT 41.660 113.390 41.920 113.710 ;
        RECT 40.340 112.350 40.940 112.430 ;
        RECT 40.280 112.290 40.940 112.350 ;
        RECT 40.280 112.030 40.540 112.290 ;
        RECT 41.720 110.310 41.860 113.390 ;
        RECT 41.660 109.990 41.920 110.310 ;
        RECT 38.720 108.435 40.260 108.805 ;
        RECT 37.520 107.950 37.780 108.270 ;
        RECT 37.060 106.930 37.320 107.250 ;
        RECT 33.440 105.490 34.040 105.630 ;
        RECT 32.920 104.550 33.180 104.870 ;
        RECT 31.540 101.490 31.800 101.810 ;
        RECT 32.460 101.490 32.720 101.810 ;
        RECT 32.980 101.550 33.120 104.550 ;
        RECT 33.440 104.530 33.580 105.490 ;
        RECT 34.300 105.065 34.560 105.210 ;
        RECT 34.290 104.695 34.570 105.065 ;
        RECT 33.380 104.440 33.640 104.530 ;
        RECT 33.380 104.300 34.040 104.440 ;
        RECT 33.380 104.210 33.640 104.300 ;
        RECT 33.380 103.530 33.640 103.850 ;
        RECT 33.440 102.150 33.580 103.530 ;
        RECT 33.380 101.830 33.640 102.150 ;
        RECT 29.700 101.150 29.960 101.470 ;
        RECT 26.940 99.790 27.200 100.110 ;
        RECT 25.560 99.110 25.820 99.430 ;
        RECT 25.620 97.390 25.760 99.110 ;
        RECT 25.560 97.070 25.820 97.390 ;
        RECT 25.560 92.650 25.820 92.970 ;
        RECT 25.620 90.590 25.760 92.650 ;
        RECT 27.000 90.930 27.140 99.790 ;
        RECT 29.760 99.090 29.900 101.150 ;
        RECT 31.600 99.430 31.740 101.490 ;
        RECT 32.980 101.410 33.580 101.550 ;
        RECT 33.900 101.470 34.040 104.300 ;
        RECT 34.820 102.490 34.960 106.250 ;
        RECT 35.280 106.170 36.340 106.310 ;
        RECT 35.670 104.015 35.950 104.385 ;
        RECT 34.760 102.170 35.020 102.490 ;
        RECT 34.300 101.490 34.560 101.810 ;
        RECT 33.440 99.770 33.580 101.410 ;
        RECT 33.840 101.150 34.100 101.470 ;
        RECT 34.360 99.770 34.500 101.490 ;
        RECT 34.760 100.810 35.020 101.130 ;
        RECT 33.380 99.450 33.640 99.770 ;
        RECT 34.300 99.450 34.560 99.770 ;
        RECT 31.540 99.110 31.800 99.430 ;
        RECT 29.700 98.770 29.960 99.090 ;
        RECT 30.620 98.430 30.880 98.750 ;
        RECT 30.680 96.370 30.820 98.430 ;
        RECT 30.620 96.050 30.880 96.370 ;
        RECT 30.620 91.630 30.880 91.950 ;
        RECT 26.940 90.610 27.200 90.930 ;
        RECT 28.320 90.610 28.580 90.930 ;
        RECT 25.560 90.270 25.820 90.590 ;
        RECT 25.560 81.770 25.820 82.090 ;
        RECT 25.620 77.670 25.760 81.770 ;
        RECT 28.380 80.390 28.520 90.610 ;
        RECT 30.680 89.230 30.820 91.630 ;
        RECT 31.080 89.930 31.340 90.250 ;
        RECT 30.620 88.910 30.880 89.230 ;
        RECT 31.140 88.550 31.280 89.930 ;
        RECT 30.620 88.230 30.880 88.550 ;
        RECT 31.080 88.230 31.340 88.550 ;
        RECT 28.320 80.070 28.580 80.390 ;
        RECT 26.940 79.050 27.200 79.370 ;
        RECT 27.000 77.670 27.140 79.050 ;
        RECT 30.680 78.350 30.820 88.230 ;
        RECT 30.620 78.030 30.880 78.350 ;
        RECT 25.560 77.350 25.820 77.670 ;
        RECT 26.940 77.350 27.200 77.670 ;
        RECT 31.600 73.930 31.740 99.110 ;
        RECT 32.460 98.090 32.720 98.410 ;
        RECT 32.920 98.090 33.180 98.410 ;
        RECT 32.520 96.710 32.660 98.090 ;
        RECT 32.980 97.390 33.120 98.090 ;
        RECT 32.920 97.070 33.180 97.390 ;
        RECT 32.460 96.390 32.720 96.710 ;
        RECT 32.920 96.050 33.180 96.370 ;
        RECT 32.980 91.950 33.120 96.050 ;
        RECT 33.440 96.030 33.580 99.450 ;
        RECT 33.840 98.430 34.100 98.750 ;
        RECT 33.900 97.390 34.040 98.430 ;
        RECT 33.840 97.070 34.100 97.390 ;
        RECT 33.380 95.710 33.640 96.030 ;
        RECT 33.900 95.430 34.040 97.070 ;
        RECT 33.440 95.290 34.040 95.430 ;
        RECT 32.920 91.630 33.180 91.950 ;
        RECT 32.920 90.610 33.180 90.930 ;
        RECT 32.980 88.890 33.120 90.610 ;
        RECT 32.920 88.570 33.180 88.890 ;
        RECT 33.440 88.210 33.580 95.290 ;
        RECT 34.360 92.970 34.500 99.450 ;
        RECT 34.820 99.090 34.960 100.810 ;
        RECT 35.740 99.430 35.880 104.015 ;
        RECT 35.680 99.110 35.940 99.430 ;
        RECT 34.760 98.770 35.020 99.090 ;
        RECT 35.220 98.090 35.480 98.410 ;
        RECT 35.280 97.050 35.420 98.090 ;
        RECT 36.200 97.390 36.340 106.170 ;
        RECT 36.600 105.230 36.860 105.550 ;
        RECT 36.660 102.830 36.800 105.230 ;
        RECT 36.600 102.510 36.860 102.830 ;
        RECT 37.120 101.130 37.260 106.930 ;
        RECT 37.520 106.590 37.780 106.910 ;
        RECT 37.580 103.850 37.720 106.590 ;
        RECT 37.980 106.250 38.240 106.570 ;
        RECT 37.520 103.530 37.780 103.850 ;
        RECT 38.040 101.810 38.180 106.250 ;
        RECT 41.190 104.695 41.470 105.065 ;
        RECT 41.260 104.530 41.400 104.695 ;
        RECT 41.200 104.210 41.460 104.530 ;
        RECT 38.720 102.995 40.260 103.365 ;
        RECT 41.260 102.590 41.400 104.210 ;
        RECT 40.800 102.450 41.400 102.590 ;
        RECT 37.980 101.490 38.240 101.810 ;
        RECT 37.060 100.810 37.320 101.130 ;
        RECT 36.140 97.070 36.400 97.390 ;
        RECT 35.220 96.730 35.480 97.050 ;
        RECT 35.280 96.370 35.420 96.730 ;
        RECT 35.220 96.050 35.480 96.370 ;
        RECT 35.680 93.670 35.940 93.990 ;
        RECT 34.300 92.650 34.560 92.970 ;
        RECT 34.760 88.230 35.020 88.550 ;
        RECT 33.380 87.890 33.640 88.210 ;
        RECT 34.820 85.150 34.960 88.230 ;
        RECT 35.740 87.870 35.880 93.670 ;
        RECT 36.140 93.330 36.400 93.650 ;
        RECT 36.200 91.950 36.340 93.330 ;
        RECT 36.140 91.630 36.400 91.950 ;
        RECT 36.600 90.950 36.860 91.270 ;
        RECT 36.140 90.270 36.400 90.590 ;
        RECT 36.200 88.550 36.340 90.270 ;
        RECT 36.660 88.890 36.800 90.950 ;
        RECT 36.600 88.570 36.860 88.890 ;
        RECT 36.140 88.230 36.400 88.550 ;
        RECT 35.680 87.550 35.940 87.870 ;
        RECT 34.760 84.830 35.020 85.150 ;
        RECT 32.000 81.770 32.260 82.090 ;
        RECT 32.060 80.050 32.200 81.770 ;
        RECT 32.000 79.730 32.260 80.050 ;
        RECT 34.820 78.350 34.960 84.830 ;
        RECT 35.220 82.790 35.480 83.110 ;
        RECT 35.280 81.070 35.420 82.790 ;
        RECT 35.680 82.000 35.940 82.090 ;
        RECT 36.200 82.000 36.340 88.230 ;
        RECT 37.120 83.790 37.260 100.810 ;
        RECT 40.800 100.110 40.940 102.450 ;
        RECT 40.740 99.790 41.000 100.110 ;
        RECT 38.720 97.555 40.260 97.925 ;
        RECT 40.800 96.370 40.940 99.790 ;
        RECT 40.740 96.050 41.000 96.370 ;
        RECT 41.200 95.710 41.460 96.030 ;
        RECT 41.260 93.310 41.400 95.710 ;
        RECT 42.120 93.670 42.380 93.990 ;
        RECT 41.200 92.990 41.460 93.310 ;
        RECT 38.720 92.115 40.260 92.485 ;
        RECT 42.180 91.950 42.320 93.670 ;
        RECT 42.120 91.630 42.380 91.950 ;
        RECT 37.520 90.840 37.780 90.930 ;
        RECT 37.520 90.700 38.180 90.840 ;
        RECT 37.520 90.610 37.780 90.700 ;
        RECT 38.040 88.550 38.180 90.700 ;
        RECT 43.040 90.610 43.300 90.930 ;
        RECT 40.280 90.270 40.540 90.590 ;
        RECT 37.980 88.230 38.240 88.550 ;
        RECT 37.520 87.210 37.780 87.530 ;
        RECT 37.580 85.490 37.720 87.210 ;
        RECT 38.040 86.170 38.180 88.230 ;
        RECT 40.340 87.950 40.480 90.270 ;
        RECT 41.200 89.930 41.460 90.250 ;
        RECT 41.260 88.550 41.400 89.930 ;
        RECT 41.200 88.230 41.460 88.550 ;
        RECT 43.100 88.210 43.240 90.610 ;
        RECT 43.560 90.250 43.700 117.810 ;
        RECT 43.960 117.470 44.220 117.790 ;
        RECT 44.020 115.410 44.160 117.470 ;
        RECT 45.860 116.430 46.000 118.830 ;
        RECT 45.800 116.110 46.060 116.430 ;
        RECT 46.780 115.750 46.920 120.190 ;
        RECT 47.240 120.170 47.380 123.250 ;
        RECT 49.080 120.850 49.220 126.570 ;
        RECT 49.540 125.610 49.680 148.840 ;
        RECT 49.940 148.070 50.200 148.390 ;
        RECT 50.400 148.070 50.660 148.390 ;
        RECT 50.000 144.650 50.140 148.070 ;
        RECT 50.460 146.350 50.600 148.070 ;
        RECT 50.400 146.030 50.660 146.350 ;
        RECT 49.940 144.330 50.200 144.650 ;
        RECT 50.920 140.140 51.060 149.690 ;
        RECT 51.780 148.750 52.040 149.070 ;
        RECT 51.840 145.330 51.980 148.750 ;
        RECT 52.300 147.710 52.440 149.770 ;
        RECT 52.700 148.410 52.960 148.730 ;
        RECT 52.240 147.390 52.500 147.710 ;
        RECT 52.300 146.010 52.440 147.390 ;
        RECT 52.240 145.690 52.500 146.010 ;
        RECT 51.780 145.010 52.040 145.330 ;
        RECT 51.320 144.330 51.580 144.650 ;
        RECT 51.380 140.910 51.520 144.330 ;
        RECT 52.300 142.950 52.440 145.690 ;
        RECT 52.760 145.670 52.900 148.410 ;
        RECT 52.700 145.350 52.960 145.670 ;
        RECT 52.240 142.630 52.500 142.950 ;
        RECT 52.240 141.610 52.500 141.930 ;
        RECT 51.320 140.590 51.580 140.910 ;
        RECT 50.000 140.000 51.060 140.140 ;
        RECT 49.480 125.290 49.740 125.610 ;
        RECT 49.020 120.530 49.280 120.850 ;
        RECT 47.180 119.850 47.440 120.170 ;
        RECT 47.240 118.810 47.380 119.850 ;
        RECT 47.180 118.490 47.440 118.810 ;
        RECT 50.000 117.450 50.140 140.000 ;
        RECT 52.300 139.890 52.440 141.610 ;
        RECT 52.760 140.230 52.900 145.350 ;
        RECT 52.700 139.910 52.960 140.230 ;
        RECT 53.220 139.890 53.360 169.150 ;
        RECT 55.520 167.770 55.660 169.830 ;
        RECT 55.460 167.450 55.720 167.770 ;
        RECT 57.820 167.430 57.960 169.830 ;
        RECT 57.760 167.110 58.020 167.430 ;
        RECT 57.300 166.770 57.560 167.090 ;
        RECT 54.540 166.090 54.800 166.410 ;
        RECT 55.000 166.090 55.260 166.410 ;
        RECT 54.600 164.710 54.740 166.090 ;
        RECT 53.620 164.390 53.880 164.710 ;
        RECT 54.540 164.390 54.800 164.710 ;
        RECT 53.680 162.330 53.820 164.390 ;
        RECT 53.620 162.010 53.880 162.330 ;
        RECT 55.060 161.990 55.200 166.090 ;
        RECT 55.510 165.555 57.050 165.925 ;
        RECT 57.360 165.390 57.500 166.770 ;
        RECT 57.760 166.430 58.020 166.750 ;
        RECT 57.300 165.070 57.560 165.390 ;
        RECT 57.820 162.670 57.960 166.430 ;
        RECT 58.280 164.370 58.420 180.710 ;
        RECT 59.140 177.650 59.400 177.970 ;
        RECT 59.200 176.270 59.340 177.650 ;
        RECT 59.140 175.950 59.400 176.270 ;
        RECT 59.140 172.210 59.400 172.530 ;
        RECT 58.680 171.530 58.940 171.850 ;
        RECT 58.740 170.345 58.880 171.530 ;
        RECT 58.670 169.975 58.950 170.345 ;
        RECT 58.220 164.050 58.480 164.370 ;
        RECT 57.760 162.350 58.020 162.670 ;
        RECT 55.000 161.670 55.260 161.990 ;
        RECT 53.620 161.330 53.880 161.650 ;
        RECT 53.680 159.610 53.820 161.330 ;
        RECT 55.000 160.990 55.260 161.310 ;
        RECT 53.620 159.290 53.880 159.610 ;
        RECT 53.680 157.230 53.820 159.290 ;
        RECT 54.080 158.950 54.340 159.270 ;
        RECT 53.620 156.910 53.880 157.230 ;
        RECT 53.620 153.510 53.880 153.830 ;
        RECT 53.680 151.790 53.820 153.510 ;
        RECT 53.620 151.470 53.880 151.790 ;
        RECT 52.240 139.570 52.500 139.890 ;
        RECT 53.160 139.570 53.420 139.890 ;
        RECT 50.400 139.230 50.660 139.550 ;
        RECT 50.460 137.510 50.600 139.230 ;
        RECT 51.780 138.890 52.040 139.210 ;
        RECT 51.840 137.510 51.980 138.890 ;
        RECT 54.140 137.510 54.280 158.950 ;
        RECT 55.060 158.590 55.200 160.990 ;
        RECT 57.300 160.650 57.560 160.970 ;
        RECT 55.510 160.115 57.050 160.485 ;
        RECT 55.000 158.270 55.260 158.590 ;
        RECT 57.360 156.210 57.500 160.650 ;
        RECT 57.300 155.890 57.560 156.210 ;
        RECT 55.510 154.675 57.050 155.045 ;
        RECT 57.360 153.830 57.500 155.890 ;
        RECT 57.300 153.510 57.560 153.830 ;
        RECT 57.360 151.190 57.500 153.510 ;
        RECT 55.980 151.050 57.960 151.190 ;
        RECT 55.980 150.770 56.120 151.050 ;
        RECT 55.920 150.450 56.180 150.770 ;
        RECT 57.300 149.770 57.560 150.090 ;
        RECT 55.510 149.235 57.050 149.605 ;
        RECT 56.380 148.070 56.640 148.390 ;
        RECT 56.440 146.350 56.580 148.070 ;
        RECT 56.380 146.030 56.640 146.350 ;
        RECT 55.510 143.795 57.050 144.165 ;
        RECT 56.380 143.540 56.640 143.630 ;
        RECT 55.060 143.400 56.640 143.540 ;
        RECT 54.540 143.200 54.800 143.290 ;
        RECT 55.060 143.200 55.200 143.400 ;
        RECT 56.380 143.310 56.640 143.400 ;
        RECT 57.360 143.290 57.500 149.770 ;
        RECT 57.820 145.670 57.960 151.050 ;
        RECT 58.740 150.770 58.880 169.975 ;
        RECT 59.200 169.470 59.340 172.210 ;
        RECT 59.140 169.150 59.400 169.470 ;
        RECT 59.140 161.670 59.400 161.990 ;
        RECT 58.680 150.450 58.940 150.770 ;
        RECT 58.220 149.770 58.480 150.090 ;
        RECT 57.760 145.350 58.020 145.670 ;
        RECT 54.540 143.060 55.200 143.200 ;
        RECT 54.540 142.970 54.800 143.060 ;
        RECT 57.300 142.970 57.560 143.290 ;
        RECT 57.300 142.290 57.560 142.610 ;
        RECT 55.510 138.355 57.050 138.725 ;
        RECT 57.360 138.190 57.500 142.290 ;
        RECT 57.820 139.890 57.960 145.350 ;
        RECT 58.280 145.330 58.420 149.770 ;
        RECT 58.220 145.010 58.480 145.330 ;
        RECT 59.200 144.650 59.340 161.670 ;
        RECT 59.660 155.530 59.800 182.410 ;
        RECT 61.440 181.050 61.700 181.370 ;
        RECT 61.500 175.590 61.640 181.050 ;
        RECT 61.960 178.310 62.100 183.090 ;
        RECT 66.100 183.070 66.240 186.150 ;
        RECT 67.020 183.750 67.160 188.190 ;
        RECT 67.880 186.150 68.140 186.470 ;
        RECT 66.960 183.430 67.220 183.750 ;
        RECT 66.040 182.750 66.300 183.070 ;
        RECT 66.960 182.410 67.220 182.730 ;
        RECT 64.200 180.370 64.460 180.690 ;
        RECT 61.900 177.990 62.160 178.310 ;
        RECT 63.740 177.540 64.000 177.630 ;
        RECT 64.260 177.540 64.400 180.370 ;
        RECT 63.740 177.400 64.400 177.540 ;
        RECT 63.740 177.310 64.000 177.400 ;
        RECT 64.260 176.270 64.400 177.400 ;
        RECT 66.500 177.310 66.760 177.630 ;
        RECT 66.560 176.270 66.700 177.310 ;
        RECT 64.200 175.950 64.460 176.270 ;
        RECT 66.500 175.950 66.760 176.270 ;
        RECT 67.020 175.590 67.160 182.410 ;
        RECT 67.940 181.030 68.080 186.150 ;
        RECT 68.340 185.130 68.600 185.450 ;
        RECT 68.400 181.030 68.540 185.130 ;
        RECT 68.860 184.430 69.000 188.530 ;
        RECT 68.800 184.110 69.060 184.430 ;
        RECT 69.320 183.660 69.460 190.570 ;
        RECT 70.180 189.550 70.440 189.870 ;
        RECT 69.720 186.490 69.980 186.810 ;
        RECT 68.860 183.520 69.460 183.660 ;
        RECT 67.880 180.710 68.140 181.030 ;
        RECT 68.340 180.710 68.600 181.030 ;
        RECT 67.940 178.990 68.080 180.710 ;
        RECT 68.340 180.030 68.600 180.350 ;
        RECT 67.880 178.670 68.140 178.990 ;
        RECT 67.420 177.650 67.680 177.970 ;
        RECT 60.060 175.270 60.320 175.590 ;
        RECT 61.440 175.270 61.700 175.590 ;
        RECT 66.960 175.270 67.220 175.590 ;
        RECT 59.600 155.210 59.860 155.530 ;
        RECT 59.140 144.330 59.400 144.650 ;
        RECT 59.140 141.950 59.400 142.270 ;
        RECT 57.760 139.570 58.020 139.890 ;
        RECT 57.300 137.870 57.560 138.190 ;
        RECT 57.820 137.850 57.960 139.570 ;
        RECT 58.220 139.230 58.480 139.550 ;
        RECT 58.280 138.190 58.420 139.230 ;
        RECT 58.220 137.870 58.480 138.190 ;
        RECT 57.760 137.530 58.020 137.850 ;
        RECT 59.200 137.510 59.340 141.950 ;
        RECT 60.120 138.190 60.260 175.270 ;
        RECT 63.740 174.250 64.000 174.570 ;
        RECT 62.820 170.510 63.080 170.830 ;
        RECT 61.440 170.170 61.700 170.490 ;
        RECT 60.520 158.950 60.780 159.270 ;
        RECT 60.580 157.230 60.720 158.950 ;
        RECT 60.520 156.910 60.780 157.230 ;
        RECT 60.520 151.470 60.780 151.790 ;
        RECT 60.580 141.930 60.720 151.470 ;
        RECT 61.500 144.650 61.640 170.170 ;
        RECT 62.360 166.090 62.620 166.410 ;
        RECT 61.900 160.650 62.160 160.970 ;
        RECT 62.420 160.880 62.560 166.090 ;
        RECT 62.880 164.710 63.020 170.510 ;
        RECT 63.800 170.490 63.940 174.250 ;
        RECT 67.480 172.870 67.620 177.650 ;
        RECT 68.400 175.590 68.540 180.030 ;
        RECT 68.340 175.270 68.600 175.590 ;
        RECT 67.420 172.550 67.680 172.870 ;
        RECT 63.740 170.170 64.000 170.490 ;
        RECT 67.480 170.150 67.620 172.550 ;
        RECT 67.420 169.830 67.680 170.150 ;
        RECT 68.340 169.490 68.600 169.810 ;
        RECT 65.580 168.810 65.840 169.130 ;
        RECT 65.640 168.110 65.780 168.810 ;
        RECT 65.580 167.790 65.840 168.110 ;
        RECT 63.740 166.430 64.000 166.750 ;
        RECT 64.200 166.430 64.460 166.750 ;
        RECT 63.800 165.390 63.940 166.430 ;
        RECT 63.740 165.070 64.000 165.390 ;
        RECT 62.820 164.390 63.080 164.710 ;
        RECT 64.260 164.370 64.400 166.430 ;
        RECT 65.640 164.690 65.780 167.790 ;
        RECT 65.180 164.550 65.780 164.690 ;
        RECT 64.200 164.050 64.460 164.370 ;
        RECT 63.280 162.350 63.540 162.670 ;
        RECT 62.820 160.880 63.080 160.970 ;
        RECT 62.420 160.740 63.080 160.880 ;
        RECT 62.820 160.650 63.080 160.740 ;
        RECT 61.960 156.210 62.100 160.650 ;
        RECT 62.360 159.290 62.620 159.610 ;
        RECT 62.420 157.230 62.560 159.290 ;
        RECT 62.880 159.270 63.020 160.650 ;
        RECT 62.820 158.950 63.080 159.270 ;
        RECT 63.340 158.250 63.480 162.350 ;
        RECT 63.740 158.950 64.000 159.270 ;
        RECT 63.280 157.930 63.540 158.250 ;
        RECT 62.360 156.910 62.620 157.230 ;
        RECT 61.900 155.890 62.160 156.210 ;
        RECT 62.420 155.870 62.560 156.910 ;
        RECT 62.360 155.550 62.620 155.870 ;
        RECT 61.900 152.490 62.160 152.810 ;
        RECT 61.960 150.430 62.100 152.490 ;
        RECT 61.900 150.110 62.160 150.430 ;
        RECT 62.820 150.110 63.080 150.430 ;
        RECT 62.880 149.070 63.020 150.110 ;
        RECT 63.800 150.090 63.940 158.950 ;
        RECT 64.260 158.930 64.400 164.050 ;
        RECT 65.180 162.670 65.320 164.550 ;
        RECT 66.960 164.390 67.220 164.710 ;
        RECT 67.420 164.690 67.680 164.710 ;
        RECT 68.400 164.690 68.540 169.490 ;
        RECT 68.860 168.110 69.000 183.520 ;
        RECT 69.260 182.750 69.520 183.070 ;
        RECT 68.800 167.790 69.060 168.110 ;
        RECT 69.320 164.690 69.460 182.750 ;
        RECT 69.780 181.620 69.920 186.490 ;
        RECT 70.240 186.470 70.380 189.550 ;
        RECT 70.640 188.190 70.900 188.510 ;
        RECT 70.180 186.150 70.440 186.470 ;
        RECT 70.240 182.730 70.380 186.150 ;
        RECT 70.700 183.410 70.840 188.190 ;
        RECT 71.100 187.850 71.360 188.170 ;
        RECT 71.160 186.470 71.300 187.850 ;
        RECT 71.100 186.150 71.360 186.470 ;
        RECT 71.100 185.470 71.360 185.790 ;
        RECT 71.160 184.430 71.300 185.470 ;
        RECT 71.100 184.110 71.360 184.430 ;
        RECT 70.640 183.090 70.900 183.410 ;
        RECT 70.180 182.410 70.440 182.730 ;
        RECT 70.180 181.620 70.440 181.710 ;
        RECT 69.780 181.480 70.440 181.620 ;
        RECT 69.780 176.270 69.920 181.480 ;
        RECT 70.180 181.390 70.440 181.480 ;
        RECT 70.700 181.030 70.840 183.090 ;
        RECT 70.640 180.710 70.900 181.030 ;
        RECT 70.700 178.990 70.840 180.710 ;
        RECT 70.640 178.670 70.900 178.990 ;
        RECT 70.180 177.990 70.440 178.310 ;
        RECT 69.720 175.950 69.980 176.270 ;
        RECT 70.240 175.590 70.380 177.990 ;
        RECT 70.180 175.270 70.440 175.590 ;
        RECT 69.720 171.870 69.980 172.190 ;
        RECT 69.780 170.830 69.920 171.870 ;
        RECT 70.240 171.850 70.380 175.270 ;
        RECT 71.160 175.250 71.300 184.110 ;
        RECT 71.620 183.070 71.760 193.630 ;
        RECT 74.380 191.910 74.520 193.970 ;
        RECT 74.320 191.590 74.580 191.910 ;
        RECT 74.320 190.570 74.580 190.890 ;
        RECT 72.300 190.035 73.840 190.405 ;
        RECT 72.480 188.530 72.740 188.850 ;
        RECT 73.860 188.760 74.120 188.850 ;
        RECT 74.380 188.760 74.520 190.570 ;
        RECT 75.300 188.850 75.440 196.010 ;
        RECT 75.760 194.970 75.900 199.070 ;
        RECT 76.620 198.730 76.880 199.050 ;
        RECT 76.160 196.350 76.420 196.670 ;
        RECT 75.700 194.650 75.960 194.970 ;
        RECT 75.760 192.250 75.900 194.650 ;
        RECT 76.220 194.290 76.360 196.350 ;
        RECT 76.680 196.330 76.820 198.730 ;
        RECT 76.620 196.010 76.880 196.330 ;
        RECT 77.140 194.710 77.280 199.330 ;
        RECT 80.760 199.070 81.020 199.390 ;
        RECT 77.540 197.370 77.800 197.690 ;
        RECT 76.680 194.630 77.280 194.710 ;
        RECT 76.620 194.570 77.280 194.630 ;
        RECT 76.620 194.310 76.880 194.570 ;
        RECT 76.160 193.970 76.420 194.290 ;
        RECT 77.600 193.610 77.740 197.370 ;
        RECT 78.920 196.010 79.180 196.330 ;
        RECT 78.000 193.630 78.260 193.950 ;
        RECT 77.540 193.290 77.800 193.610 ;
        RECT 78.060 192.590 78.200 193.630 ;
        RECT 78.000 192.270 78.260 192.590 ;
        RECT 75.700 191.930 75.960 192.250 ;
        RECT 78.980 191.910 79.120 196.010 ;
        RECT 78.920 191.590 79.180 191.910 ;
        RECT 79.840 190.570 80.100 190.890 ;
        RECT 79.900 188.850 80.040 190.570 ;
        RECT 73.860 188.620 74.520 188.760 ;
        RECT 73.860 188.530 74.120 188.620 ;
        RECT 72.540 185.790 72.680 188.530 ;
        RECT 72.480 185.470 72.740 185.790 ;
        RECT 72.300 184.595 73.840 184.965 ;
        RECT 74.380 183.750 74.520 188.620 ;
        RECT 75.240 188.530 75.500 188.850 ;
        RECT 75.700 188.530 75.960 188.850 ;
        RECT 79.840 188.530 80.100 188.850 ;
        RECT 75.760 188.170 75.900 188.530 ;
        RECT 75.700 188.080 75.960 188.170 ;
        RECT 75.700 187.940 76.360 188.080 ;
        RECT 75.700 187.850 75.960 187.940 ;
        RECT 74.780 185.130 75.040 185.450 ;
        RECT 74.840 184.090 74.980 185.130 ;
        RECT 74.780 183.770 75.040 184.090 ;
        RECT 75.240 183.770 75.500 184.090 ;
        RECT 74.320 183.430 74.580 183.750 ;
        RECT 71.560 182.750 71.820 183.070 ;
        RECT 71.560 180.030 71.820 180.350 ;
        RECT 71.620 177.630 71.760 180.030 ;
        RECT 74.840 180.010 74.980 183.770 ;
        RECT 75.300 181.370 75.440 183.770 ;
        RECT 75.700 183.430 75.960 183.750 ;
        RECT 75.240 181.050 75.500 181.370 ;
        RECT 75.760 181.030 75.900 183.430 ;
        RECT 76.220 183.410 76.360 187.940 ;
        RECT 77.080 187.850 77.340 188.170 ;
        RECT 78.000 187.850 78.260 188.170 ;
        RECT 77.140 187.150 77.280 187.850 ;
        RECT 77.080 186.830 77.340 187.150 ;
        RECT 78.060 186.470 78.200 187.850 ;
        RECT 78.460 186.490 78.720 186.810 ;
        RECT 78.000 186.150 78.260 186.470 ;
        RECT 77.080 185.810 77.340 186.130 ;
        RECT 76.160 183.090 76.420 183.410 ;
        RECT 75.700 180.710 75.960 181.030 ;
        RECT 74.780 179.690 75.040 180.010 ;
        RECT 72.300 179.155 73.840 179.525 ;
        RECT 71.560 177.310 71.820 177.630 ;
        RECT 71.560 175.950 71.820 176.270 ;
        RECT 71.100 174.930 71.360 175.250 ;
        RECT 70.640 174.250 70.900 174.570 ;
        RECT 70.180 171.530 70.440 171.850 ;
        RECT 69.720 170.510 69.980 170.830 ;
        RECT 70.240 169.810 70.380 171.530 ;
        RECT 70.700 170.150 70.840 174.250 ;
        RECT 71.160 173.550 71.300 174.930 ;
        RECT 71.100 173.230 71.360 173.550 ;
        RECT 71.620 170.910 71.760 175.950 ;
        RECT 74.840 175.500 74.980 179.690 ;
        RECT 75.760 178.310 75.900 180.710 ;
        RECT 76.220 178.990 76.360 183.090 ;
        RECT 76.160 178.670 76.420 178.990 ;
        RECT 75.700 177.990 75.960 178.310 ;
        RECT 75.760 177.290 75.900 177.990 ;
        RECT 75.700 176.970 75.960 177.290 ;
        RECT 74.380 175.360 74.980 175.500 ;
        RECT 74.380 174.570 74.520 175.360 ;
        RECT 75.700 175.270 75.960 175.590 ;
        RECT 74.780 174.590 75.040 174.910 ;
        RECT 74.320 174.250 74.580 174.570 ;
        RECT 72.300 173.715 73.840 174.085 ;
        RECT 74.380 172.870 74.520 174.250 ;
        RECT 72.480 172.550 72.740 172.870 ;
        RECT 74.320 172.550 74.580 172.870 ;
        RECT 71.160 170.770 71.760 170.910 ;
        RECT 70.640 169.830 70.900 170.150 ;
        RECT 70.180 169.490 70.440 169.810 ;
        RECT 70.640 166.090 70.900 166.410 ;
        RECT 70.700 165.050 70.840 166.090 ;
        RECT 71.160 165.390 71.300 170.770 ;
        RECT 71.550 169.975 71.830 170.345 ;
        RECT 71.560 169.830 71.820 169.975 ;
        RECT 72.540 169.550 72.680 172.550 ;
        RECT 71.620 169.410 72.680 169.550 ;
        RECT 71.100 165.070 71.360 165.390 ;
        RECT 70.640 164.730 70.900 165.050 ;
        RECT 67.420 164.550 68.540 164.690 ;
        RECT 68.860 164.550 69.460 164.690 ;
        RECT 67.420 164.390 67.680 164.550 ;
        RECT 67.020 163.690 67.160 164.390 ;
        RECT 66.960 163.370 67.220 163.690 ;
        RECT 65.120 162.350 65.380 162.670 ;
        RECT 64.660 162.010 64.920 162.330 ;
        RECT 64.720 161.310 64.860 162.010 ;
        RECT 64.660 160.990 64.920 161.310 ;
        RECT 68.860 159.950 69.000 164.550 ;
        RECT 70.640 164.050 70.900 164.370 ;
        RECT 69.720 163.370 69.980 163.690 ;
        RECT 68.800 159.630 69.060 159.950 ;
        RECT 68.330 159.095 68.610 159.465 ;
        RECT 68.340 158.950 68.600 159.095 ;
        RECT 64.200 158.610 64.460 158.930 ;
        RECT 67.880 158.610 68.140 158.930 ;
        RECT 64.200 157.930 64.460 158.250 ;
        RECT 64.260 153.830 64.400 157.930 ;
        RECT 67.940 156.120 68.080 158.610 ;
        RECT 68.340 158.270 68.600 158.590 ;
        RECT 68.400 156.745 68.540 158.270 ;
        RECT 68.330 156.375 68.610 156.745 ;
        RECT 68.340 156.120 68.600 156.210 ;
        RECT 67.940 155.980 68.600 156.120 ;
        RECT 65.120 155.550 65.380 155.870 ;
        RECT 65.180 154.510 65.320 155.550 ;
        RECT 65.120 154.190 65.380 154.510 ;
        RECT 64.200 153.510 64.460 153.830 ;
        RECT 67.420 150.110 67.680 150.430 ;
        RECT 63.740 149.770 64.000 150.090 ;
        RECT 64.660 149.770 64.920 150.090 ;
        RECT 62.820 148.750 63.080 149.070 ;
        RECT 62.820 148.070 63.080 148.390 ;
        RECT 61.900 147.050 62.160 147.370 ;
        RECT 61.440 144.330 61.700 144.650 ;
        RECT 61.960 143.710 62.100 147.050 ;
        RECT 62.880 146.350 63.020 148.070 ;
        RECT 62.820 146.030 63.080 146.350 ;
        RECT 64.720 145.330 64.860 149.770 ;
        RECT 64.660 145.010 64.920 145.330 ;
        RECT 67.480 144.990 67.620 150.110 ;
        RECT 67.940 148.050 68.080 155.980 ;
        RECT 68.340 155.890 68.600 155.980 ;
        RECT 68.860 150.430 69.000 159.630 ;
        RECT 69.260 159.290 69.520 159.610 ;
        RECT 69.320 153.830 69.460 159.290 ;
        RECT 69.260 153.510 69.520 153.830 ;
        RECT 68.800 150.110 69.060 150.430 ;
        RECT 67.880 147.730 68.140 148.050 ;
        RECT 67.940 144.990 68.080 147.730 ;
        RECT 67.420 144.670 67.680 144.990 ;
        RECT 67.880 144.670 68.140 144.990 ;
        RECT 61.500 143.570 62.100 143.710 ;
        RECT 60.520 141.610 60.780 141.930 ;
        RECT 60.060 137.870 60.320 138.190 ;
        RECT 50.400 137.190 50.660 137.510 ;
        RECT 51.780 137.190 52.040 137.510 ;
        RECT 53.160 137.190 53.420 137.510 ;
        RECT 54.080 137.190 54.340 137.510 ;
        RECT 59.140 137.190 59.400 137.510 ;
        RECT 50.460 129.010 50.600 137.190 ;
        RECT 52.240 134.130 52.500 134.450 ;
        RECT 52.300 132.750 52.440 134.130 ;
        RECT 52.700 133.450 52.960 133.770 ;
        RECT 52.240 132.430 52.500 132.750 ;
        RECT 50.860 132.090 51.120 132.410 ;
        RECT 50.400 128.690 50.660 129.010 ;
        RECT 50.920 128.670 51.060 132.090 ;
        RECT 51.320 131.410 51.580 131.730 ;
        RECT 51.380 131.050 51.520 131.410 ;
        RECT 51.320 130.730 51.580 131.050 ;
        RECT 52.760 129.010 52.900 133.450 ;
        RECT 52.700 128.690 52.960 129.010 ;
        RECT 50.860 128.350 51.120 128.670 ;
        RECT 50.920 125.610 51.060 128.350 ;
        RECT 50.860 125.290 51.120 125.610 ;
        RECT 51.320 125.290 51.580 125.610 ;
        RECT 51.380 121.190 51.520 125.290 ;
        RECT 53.220 123.570 53.360 137.190 ;
        RECT 55.510 132.915 57.050 133.285 ;
        RECT 55.000 132.430 55.260 132.750 ;
        RECT 54.540 129.710 54.800 130.030 ;
        RECT 54.600 125.610 54.740 129.710 ;
        RECT 55.060 125.950 55.200 132.430 ;
        RECT 55.920 130.730 56.180 131.050 ;
        RECT 58.680 130.730 58.940 131.050 ;
        RECT 55.980 130.030 56.120 130.730 ;
        RECT 55.920 129.710 56.180 130.030 ;
        RECT 58.740 129.010 58.880 130.730 ;
        RECT 60.580 130.030 60.720 141.610 ;
        RECT 60.980 131.980 61.240 132.070 ;
        RECT 61.500 131.980 61.640 143.570 ;
        RECT 63.280 142.290 63.540 142.610 ;
        RECT 63.340 140.910 63.480 142.290 ;
        RECT 65.120 141.610 65.380 141.930 ;
        RECT 63.280 140.590 63.540 140.910 ;
        RECT 65.180 139.890 65.320 141.610 ;
        RECT 61.900 139.570 62.160 139.890 ;
        RECT 65.120 139.570 65.380 139.890 ;
        RECT 60.980 131.840 61.640 131.980 ;
        RECT 60.980 131.750 61.240 131.840 ;
        RECT 60.520 129.710 60.780 130.030 ;
        RECT 58.680 128.690 58.940 129.010 ;
        RECT 59.600 128.690 59.860 129.010 ;
        RECT 58.680 128.010 58.940 128.330 ;
        RECT 55.510 127.475 57.050 127.845 ;
        RECT 58.740 126.630 58.880 128.010 ;
        RECT 59.660 126.970 59.800 128.690 ;
        RECT 59.600 126.650 59.860 126.970 ;
        RECT 58.220 126.310 58.480 126.630 ;
        RECT 58.680 126.310 58.940 126.630 ;
        RECT 57.300 125.970 57.560 126.290 ;
        RECT 55.000 125.630 55.260 125.950 ;
        RECT 54.540 125.290 54.800 125.610 ;
        RECT 52.700 123.250 52.960 123.570 ;
        RECT 53.160 123.250 53.420 123.570 ;
        RECT 54.080 123.250 54.340 123.570 ;
        RECT 52.760 121.870 52.900 123.250 ;
        RECT 53.620 122.570 53.880 122.890 ;
        RECT 52.700 121.550 52.960 121.870 ;
        RECT 53.680 121.190 53.820 122.570 ;
        RECT 50.860 120.870 51.120 121.190 ;
        RECT 51.320 120.870 51.580 121.190 ;
        RECT 51.780 120.870 52.040 121.190 ;
        RECT 53.620 120.870 53.880 121.190 ;
        RECT 50.400 120.530 50.660 120.850 ;
        RECT 49.940 117.130 50.200 117.450 ;
        RECT 46.720 115.430 46.980 115.750 ;
        RECT 49.480 115.430 49.740 115.750 ;
        RECT 43.960 115.090 44.220 115.410 ;
        RECT 44.020 113.710 44.160 115.090 ;
        RECT 43.960 113.390 44.220 113.710 ;
        RECT 46.780 112.690 46.920 115.430 ;
        RECT 49.540 113.710 49.680 115.430 ;
        RECT 49.480 113.390 49.740 113.710 ;
        RECT 46.720 112.370 46.980 112.690 ;
        RECT 50.460 109.970 50.600 120.530 ;
        RECT 50.920 117.450 51.060 120.870 ;
        RECT 50.860 117.130 51.120 117.450 ;
        RECT 51.380 116.510 51.520 120.870 ;
        RECT 51.840 118.130 51.980 120.870 ;
        RECT 54.140 119.150 54.280 123.250 ;
        RECT 55.510 122.035 57.050 122.405 ;
        RECT 54.540 121.210 54.800 121.530 ;
        RECT 54.080 118.830 54.340 119.150 ;
        RECT 51.780 117.810 52.040 118.130 ;
        RECT 52.700 117.810 52.960 118.130 ;
        RECT 52.760 116.510 52.900 117.810 ;
        RECT 51.380 116.370 52.900 116.510 ;
        RECT 52.760 112.350 52.900 116.370 ;
        RECT 53.160 112.710 53.420 113.030 ;
        RECT 52.700 112.030 52.960 112.350 ;
        RECT 53.220 110.310 53.360 112.710 ;
        RECT 53.620 112.370 53.880 112.690 ;
        RECT 53.680 110.990 53.820 112.370 ;
        RECT 53.620 110.670 53.880 110.990 ;
        RECT 54.140 110.310 54.280 118.830 ;
        RECT 54.600 113.710 54.740 121.210 ;
        RECT 55.510 116.595 57.050 116.965 ;
        RECT 55.000 114.750 55.260 115.070 ;
        RECT 54.540 113.390 54.800 113.710 ;
        RECT 54.540 111.690 54.800 112.010 ;
        RECT 54.600 110.990 54.740 111.690 ;
        RECT 54.540 110.670 54.800 110.990 ;
        RECT 53.160 109.990 53.420 110.310 ;
        RECT 54.080 109.990 54.340 110.310 ;
        RECT 50.400 109.650 50.660 109.970 ;
        RECT 53.220 109.710 53.360 109.990 ;
        RECT 43.960 106.930 44.220 107.250 ;
        RECT 49.940 107.160 50.200 107.250 ;
        RECT 50.460 107.160 50.600 109.650 ;
        RECT 53.220 109.570 53.820 109.710 ;
        RECT 50.860 108.970 51.120 109.290 ;
        RECT 50.920 108.270 51.060 108.970 ;
        RECT 50.860 107.950 51.120 108.270 ;
        RECT 49.940 107.020 50.600 107.160 ;
        RECT 49.940 106.930 50.200 107.020 ;
        RECT 53.160 106.930 53.420 107.250 ;
        RECT 53.680 107.160 53.820 109.570 ;
        RECT 54.080 107.160 54.340 107.250 ;
        RECT 53.680 107.020 54.340 107.160 ;
        RECT 54.080 106.930 54.340 107.020 ;
        RECT 44.020 105.550 44.160 106.930 ;
        RECT 45.340 106.250 45.600 106.570 ;
        RECT 51.320 106.250 51.580 106.570 ;
        RECT 43.960 105.230 44.220 105.550 ;
        RECT 44.020 101.810 44.160 105.230 ;
        RECT 44.420 104.550 44.680 104.870 ;
        RECT 44.480 102.830 44.620 104.550 ;
        RECT 44.420 102.510 44.680 102.830 ;
        RECT 45.400 101.810 45.540 106.250 ;
        RECT 51.380 104.870 51.520 106.250 ;
        RECT 53.220 105.550 53.360 106.930 ;
        RECT 53.160 105.230 53.420 105.550 ;
        RECT 51.320 104.550 51.580 104.870 ;
        RECT 54.140 104.530 54.280 106.930 ;
        RECT 54.600 104.870 54.740 110.670 ;
        RECT 55.060 110.310 55.200 114.750 ;
        RECT 57.360 113.710 57.500 125.970 ;
        RECT 57.760 114.410 58.020 114.730 ;
        RECT 57.300 113.390 57.560 113.710 ;
        RECT 57.820 112.690 57.960 114.410 ;
        RECT 57.760 112.370 58.020 112.690 ;
        RECT 55.510 111.155 57.050 111.525 ;
        RECT 57.820 110.310 57.960 112.370 ;
        RECT 55.000 109.990 55.260 110.310 ;
        RECT 57.760 109.990 58.020 110.310 ;
        RECT 55.000 109.310 55.260 109.630 ;
        RECT 55.060 107.590 55.200 109.310 ;
        RECT 55.000 107.270 55.260 107.590 ;
        RECT 54.540 104.550 54.800 104.870 ;
        RECT 54.080 104.210 54.340 104.530 ;
        RECT 54.540 103.530 54.800 103.850 ;
        RECT 43.960 101.490 44.220 101.810 ;
        RECT 45.340 101.490 45.600 101.810 ;
        RECT 54.600 101.470 54.740 103.530 ;
        RECT 54.540 101.150 54.800 101.470 ;
        RECT 55.060 99.090 55.200 107.270 ;
        RECT 58.280 106.910 58.420 126.310 ;
        RECT 60.580 123.570 60.720 129.710 ;
        RECT 61.960 129.010 62.100 139.570 ;
        RECT 67.480 137.705 67.620 144.670 ;
        RECT 67.410 137.335 67.690 137.705 ;
        RECT 65.580 136.850 65.840 137.170 ;
        RECT 65.640 131.730 65.780 136.850 ;
        RECT 66.500 136.170 66.760 136.490 ;
        RECT 66.560 132.410 66.700 136.170 ;
        RECT 66.500 132.090 66.760 132.410 ;
        RECT 65.580 131.410 65.840 131.730 ;
        RECT 66.040 131.410 66.300 131.730 ;
        RECT 62.360 130.730 62.620 131.050 ;
        RECT 63.740 130.730 64.000 131.050 ;
        RECT 61.900 128.690 62.160 129.010 ;
        RECT 60.980 126.310 61.240 126.630 ;
        RECT 60.520 123.250 60.780 123.570 ;
        RECT 59.600 122.570 59.860 122.890 ;
        RECT 58.680 115.770 58.940 116.090 ;
        RECT 58.220 106.590 58.480 106.910 ;
        RECT 57.300 106.250 57.560 106.570 ;
        RECT 55.510 105.715 57.050 106.085 ;
        RECT 57.360 105.550 57.500 106.250 ;
        RECT 57.300 105.230 57.560 105.550 ;
        RECT 58.280 105.210 58.420 106.590 ;
        RECT 58.220 104.890 58.480 105.210 ;
        RECT 57.760 102.510 58.020 102.830 ;
        RECT 57.300 100.810 57.560 101.130 ;
        RECT 55.510 100.275 57.050 100.645 ;
        RECT 57.360 99.430 57.500 100.810 ;
        RECT 57.300 99.110 57.560 99.430 ;
        RECT 55.000 98.770 55.260 99.090 ;
        RECT 45.340 97.070 45.600 97.390 ;
        RECT 44.420 96.050 44.680 96.370 ;
        RECT 44.480 94.330 44.620 96.050 ;
        RECT 44.420 94.010 44.680 94.330 ;
        RECT 44.420 90.950 44.680 91.270 ;
        RECT 43.960 90.610 44.220 90.930 ;
        RECT 43.500 89.930 43.760 90.250 ;
        RECT 44.020 88.210 44.160 90.610 ;
        RECT 44.480 88.550 44.620 90.950 ;
        RECT 44.880 90.610 45.140 90.930 ;
        RECT 44.940 88.550 45.080 90.610 ;
        RECT 45.400 88.550 45.540 97.070 ;
        RECT 52.700 96.730 52.960 97.050 ;
        RECT 49.020 95.710 49.280 96.030 ;
        RECT 49.080 93.310 49.220 95.710 ;
        RECT 49.940 93.670 50.200 93.990 ;
        RECT 49.020 92.990 49.280 93.310 ;
        RECT 50.000 91.950 50.140 93.670 ;
        RECT 51.320 92.990 51.580 93.310 ;
        RECT 49.940 91.630 50.200 91.950 ;
        RECT 51.380 91.270 51.520 92.990 ;
        RECT 51.320 90.950 51.580 91.270 ;
        RECT 49.940 90.610 50.200 90.930 ;
        RECT 52.240 90.610 52.500 90.930 ;
        RECT 49.480 89.930 49.740 90.250 ;
        RECT 49.540 89.230 49.680 89.930 ;
        RECT 49.480 88.910 49.740 89.230 ;
        RECT 50.000 88.550 50.140 90.610 ;
        RECT 52.300 88.550 52.440 90.610 ;
        RECT 44.420 88.230 44.680 88.550 ;
        RECT 44.880 88.230 45.140 88.550 ;
        RECT 45.340 88.230 45.600 88.550 ;
        RECT 46.260 88.230 46.520 88.550 ;
        RECT 49.940 88.230 50.200 88.550 ;
        RECT 52.240 88.230 52.500 88.550 ;
        RECT 52.760 88.460 52.900 96.730 ;
        RECT 54.540 96.050 54.800 96.370 ;
        RECT 53.160 94.010 53.420 94.330 ;
        RECT 53.220 91.950 53.360 94.010 ;
        RECT 54.600 93.310 54.740 96.050 ;
        RECT 55.000 95.370 55.260 95.690 ;
        RECT 55.060 94.330 55.200 95.370 ;
        RECT 55.510 94.835 57.050 95.205 ;
        RECT 55.000 94.010 55.260 94.330 ;
        RECT 54.540 92.990 54.800 93.310 ;
        RECT 53.160 91.630 53.420 91.950 ;
        RECT 54.540 90.950 54.800 91.270 ;
        RECT 53.620 90.610 53.880 90.930 ;
        RECT 54.080 90.610 54.340 90.930 ;
        RECT 53.160 88.460 53.420 88.550 ;
        RECT 52.760 88.320 53.420 88.460 ;
        RECT 40.340 87.810 40.940 87.950 ;
        RECT 43.040 87.890 43.300 88.210 ;
        RECT 43.960 87.890 44.220 88.210 ;
        RECT 38.720 86.675 40.260 87.045 ;
        RECT 40.800 86.420 40.940 87.810 ;
        RECT 43.100 86.510 43.240 87.890 ;
        RECT 40.340 86.280 40.940 86.420 ;
        RECT 37.980 85.850 38.240 86.170 ;
        RECT 37.520 85.170 37.780 85.490 ;
        RECT 38.040 85.150 38.180 85.850 ;
        RECT 40.340 85.150 40.480 86.280 ;
        RECT 43.040 86.190 43.300 86.510 ;
        RECT 45.400 85.830 45.540 88.230 ;
        RECT 46.320 86.170 46.460 88.230 ;
        RECT 50.000 86.510 50.140 88.230 ;
        RECT 49.940 86.190 50.200 86.510 ;
        RECT 46.260 85.850 46.520 86.170 ;
        RECT 45.340 85.510 45.600 85.830 ;
        RECT 42.580 85.170 42.840 85.490 ;
        RECT 43.500 85.230 43.760 85.490 ;
        RECT 43.500 85.170 44.160 85.230 ;
        RECT 44.420 85.170 44.680 85.490 ;
        RECT 48.100 85.170 48.360 85.490 ;
        RECT 50.860 85.170 51.120 85.490 ;
        RECT 37.980 84.830 38.240 85.150 ;
        RECT 40.280 84.830 40.540 85.150 ;
        RECT 38.440 84.490 38.700 84.810 ;
        RECT 37.060 83.470 37.320 83.790 ;
        RECT 38.500 83.450 38.640 84.490 ;
        RECT 38.440 83.130 38.700 83.450 ;
        RECT 42.640 83.110 42.780 85.170 ;
        RECT 43.560 85.090 44.160 85.170 ;
        RECT 40.740 82.790 41.000 83.110 ;
        RECT 41.200 82.790 41.460 83.110 ;
        RECT 42.580 82.790 42.840 83.110 ;
        RECT 35.680 81.860 36.340 82.000 ;
        RECT 35.680 81.770 35.940 81.860 ;
        RECT 35.220 80.750 35.480 81.070 ;
        RECT 35.280 80.050 35.420 80.750 ;
        RECT 35.220 79.730 35.480 80.050 ;
        RECT 34.760 78.030 35.020 78.350 ;
        RECT 35.740 77.670 35.880 81.770 ;
        RECT 38.720 81.235 40.260 81.605 ;
        RECT 40.800 80.470 40.940 82.790 ;
        RECT 41.260 81.070 41.400 82.790 ;
        RECT 41.200 80.750 41.460 81.070 ;
        RECT 44.020 80.730 44.160 85.090 ;
        RECT 44.480 83.790 44.620 85.170 ;
        RECT 48.160 83.790 48.300 85.170 ;
        RECT 44.420 83.470 44.680 83.790 ;
        RECT 48.100 83.470 48.360 83.790 ;
        RECT 50.920 83.110 51.060 85.170 ;
        RECT 52.760 85.150 52.900 88.320 ;
        RECT 53.160 88.230 53.420 88.320 ;
        RECT 53.680 88.210 53.820 90.610 ;
        RECT 54.140 89.230 54.280 90.610 ;
        RECT 54.600 89.230 54.740 90.950 ;
        RECT 55.000 89.930 55.260 90.250 ;
        RECT 54.080 88.910 54.340 89.230 ;
        RECT 54.540 88.910 54.800 89.230 ;
        RECT 55.060 88.890 55.200 89.930 ;
        RECT 55.510 89.395 57.050 89.765 ;
        RECT 55.000 88.570 55.260 88.890 ;
        RECT 54.080 88.230 54.340 88.550 ;
        RECT 53.620 87.890 53.880 88.210 ;
        RECT 54.140 85.830 54.280 88.230 ;
        RECT 54.080 85.510 54.340 85.830 ;
        RECT 57.300 85.170 57.560 85.490 ;
        RECT 52.700 84.830 52.960 85.150 ;
        RECT 55.000 84.830 55.260 85.150 ;
        RECT 44.420 82.790 44.680 83.110 ;
        RECT 50.860 82.790 51.120 83.110 ;
        RECT 51.320 82.790 51.580 83.110 ;
        RECT 40.800 80.330 41.400 80.470 ;
        RECT 43.960 80.410 44.220 80.730 ;
        RECT 41.260 79.710 41.400 80.330 ;
        RECT 36.600 79.390 36.860 79.710 ;
        RECT 41.200 79.390 41.460 79.710 ;
        RECT 36.660 78.350 36.800 79.390 ;
        RECT 37.980 79.050 38.240 79.370 ;
        RECT 36.600 78.030 36.860 78.350 ;
        RECT 38.040 78.010 38.180 79.050 ;
        RECT 37.980 77.690 38.240 78.010 ;
        RECT 35.680 77.350 35.940 77.670 ;
        RECT 34.760 76.330 35.020 76.650 ;
        RECT 34.820 74.950 34.960 76.330 ;
        RECT 38.720 75.795 40.260 76.165 ;
        RECT 41.260 75.630 41.400 79.390 ;
        RECT 44.480 78.350 44.620 82.790 ;
        RECT 51.380 81.070 51.520 82.790 ;
        RECT 55.060 82.430 55.200 84.830 ;
        RECT 55.510 83.955 57.050 84.325 ;
        RECT 55.000 82.110 55.260 82.430 ;
        RECT 55.920 82.110 56.180 82.430 ;
        RECT 51.320 80.750 51.580 81.070 ;
        RECT 52.240 80.750 52.500 81.070 ;
        RECT 50.400 80.070 50.660 80.390 ;
        RECT 44.880 79.730 45.140 80.050 ;
        RECT 46.260 79.730 46.520 80.050 ;
        RECT 49.480 79.730 49.740 80.050 ;
        RECT 44.940 78.350 45.080 79.730 ;
        RECT 44.420 78.030 44.680 78.350 ;
        RECT 44.880 78.030 45.140 78.350 ;
        RECT 43.500 77.350 43.760 77.670 ;
        RECT 45.800 77.350 46.060 77.670 ;
        RECT 41.200 75.310 41.460 75.630 ;
        RECT 34.760 74.630 35.020 74.950 ;
        RECT 34.300 74.290 34.560 74.610 ;
        RECT 37.060 74.290 37.320 74.610 ;
        RECT 31.540 73.610 31.800 73.930 ;
        RECT 34.360 72.910 34.500 74.290 ;
        RECT 36.140 73.840 36.400 73.930 ;
        RECT 37.120 73.840 37.260 74.290 ;
        RECT 40.740 73.950 41.000 74.270 ;
        RECT 36.140 73.700 37.260 73.840 ;
        RECT 36.140 73.610 36.400 73.700 ;
        RECT 34.300 72.590 34.560 72.910 ;
        RECT 40.800 72.230 40.940 73.950 ;
        RECT 41.200 72.250 41.460 72.570 ;
        RECT 37.980 71.910 38.240 72.230 ;
        RECT 40.280 71.910 40.540 72.230 ;
        RECT 40.740 71.910 41.000 72.230 ;
        RECT 37.520 71.230 37.780 71.550 ;
        RECT 37.580 69.170 37.720 71.230 ;
        RECT 38.040 69.850 38.180 71.910 ;
        RECT 40.340 71.120 40.480 71.910 ;
        RECT 40.340 70.980 40.940 71.120 ;
        RECT 38.720 70.355 40.260 70.725 ;
        RECT 37.980 69.530 38.240 69.850 ;
        RECT 40.800 69.590 40.940 70.980 ;
        RECT 41.260 70.190 41.400 72.250 ;
        RECT 43.560 70.190 43.700 77.350 ;
        RECT 44.420 74.970 44.680 75.290 ;
        RECT 43.960 70.890 44.220 71.210 ;
        RECT 44.020 70.190 44.160 70.890 ;
        RECT 41.200 69.870 41.460 70.190 ;
        RECT 43.500 69.870 43.760 70.190 ;
        RECT 43.960 69.870 44.220 70.190 ;
        RECT 40.340 69.450 40.940 69.590 ;
        RECT 43.040 69.530 43.300 69.850 ;
        RECT 44.480 69.590 44.620 74.970 ;
        RECT 45.860 72.910 46.000 77.350 ;
        RECT 46.320 75.290 46.460 79.730 ;
        RECT 49.540 78.350 49.680 79.730 ;
        RECT 49.480 78.030 49.740 78.350 ;
        RECT 49.940 77.690 50.200 78.010 ;
        RECT 46.260 74.970 46.520 75.290 ;
        RECT 50.000 73.930 50.140 77.690 ;
        RECT 50.460 76.650 50.600 80.070 ;
        RECT 50.860 79.730 51.120 80.050 ;
        RECT 50.920 79.370 51.060 79.730 ;
        RECT 50.860 79.050 51.120 79.370 ;
        RECT 50.400 76.330 50.660 76.650 ;
        RECT 50.920 74.610 51.060 79.050 ;
        RECT 52.300 78.010 52.440 80.750 ;
        RECT 54.540 80.410 54.800 80.730 ;
        RECT 52.240 77.690 52.500 78.010 ;
        RECT 50.860 74.290 51.120 74.610 ;
        RECT 49.940 73.610 50.200 73.930 ;
        RECT 45.800 72.590 46.060 72.910 ;
        RECT 46.720 71.230 46.980 71.550 ;
        RECT 45.800 69.870 46.060 70.190 ;
        RECT 35.680 68.850 35.940 69.170 ;
        RECT 37.520 68.850 37.780 69.170 ;
        RECT 26.020 68.170 26.280 68.490 ;
        RECT 24.640 63.410 24.900 63.730 ;
        RECT 24.700 59.310 24.840 63.410 ;
        RECT 26.080 61.350 26.220 68.170 ;
        RECT 35.740 66.450 35.880 68.850 ;
        RECT 37.060 66.470 37.320 66.790 ;
        RECT 35.680 66.130 35.940 66.450 ;
        RECT 35.740 63.730 35.880 66.130 ;
        RECT 28.780 63.410 29.040 63.730 ;
        RECT 30.620 63.410 30.880 63.730 ;
        RECT 35.680 63.410 35.940 63.730 ;
        RECT 26.020 61.030 26.280 61.350 ;
        RECT 26.480 60.010 26.740 60.330 ;
        RECT 26.540 59.310 26.680 60.010 ;
        RECT 24.640 58.990 24.900 59.310 ;
        RECT 26.480 58.990 26.740 59.310 ;
        RECT 28.840 56.220 28.980 63.410 ;
        RECT 30.680 58.290 30.820 63.410 ;
        RECT 34.760 62.730 35.020 63.050 ;
        RECT 31.540 61.370 31.800 61.690 ;
        RECT 30.620 57.970 30.880 58.290 ;
        RECT 31.600 56.220 31.740 61.370 ;
        RECT 34.820 61.350 34.960 62.730 ;
        RECT 34.760 61.030 35.020 61.350 ;
        RECT 36.140 60.690 36.400 61.010 ;
        RECT 36.600 60.690 36.860 61.010 ;
        RECT 36.200 58.970 36.340 60.690 ;
        RECT 36.660 59.310 36.800 60.690 ;
        RECT 36.600 58.990 36.860 59.310 ;
        RECT 36.140 58.650 36.400 58.970 ;
        RECT 34.300 57.970 34.560 58.290 ;
        RECT 34.360 56.220 34.500 57.970 ;
        RECT 37.120 56.220 37.260 66.470 ;
        RECT 37.580 63.730 37.720 68.850 ;
        RECT 40.340 66.790 40.480 69.450 ;
        RECT 40.280 66.470 40.540 66.790 ;
        RECT 42.580 66.470 42.840 66.790 ;
        RECT 40.340 66.110 40.480 66.470 ;
        RECT 40.280 65.790 40.540 66.110 ;
        RECT 40.740 65.450 41.000 65.770 ;
        RECT 38.720 64.915 40.260 65.285 ;
        RECT 37.520 63.410 37.780 63.730 ;
        RECT 37.980 62.730 38.240 63.050 ;
        RECT 37.520 61.370 37.780 61.690 ;
        RECT 28.770 49.740 29.050 56.220 ;
        RECT 31.530 51.790 31.810 56.220 ;
        RECT 34.290 52.390 34.570 56.220 ;
        RECT 37.050 52.890 37.330 56.220 ;
        RECT 37.580 55.990 37.720 61.370 ;
        RECT 38.040 61.350 38.180 62.730 ;
        RECT 37.980 61.030 38.240 61.350 ;
        RECT 38.720 59.475 40.260 59.845 ;
        RECT 40.800 58.630 40.940 65.450 ;
        RECT 42.640 63.730 42.780 66.470 ;
        RECT 43.100 63.730 43.240 69.530 ;
        RECT 43.560 69.450 44.620 69.590 ;
        RECT 43.560 66.790 43.700 69.450 ;
        RECT 43.960 68.850 44.220 69.170 ;
        RECT 44.880 68.850 45.140 69.170 ;
        RECT 44.020 67.470 44.160 68.850 ;
        RECT 43.960 67.150 44.220 67.470 ;
        RECT 43.500 66.470 43.760 66.790 ;
        RECT 44.420 66.470 44.680 66.790 ;
        RECT 44.480 64.150 44.620 66.470 ;
        RECT 44.940 65.770 45.080 68.850 ;
        RECT 44.880 65.450 45.140 65.770 ;
        RECT 43.560 64.070 44.620 64.150 ;
        RECT 43.500 64.010 44.620 64.070 ;
        RECT 43.500 63.750 43.760 64.010 ;
        RECT 41.200 63.410 41.460 63.730 ;
        RECT 42.580 63.410 42.840 63.730 ;
        RECT 43.040 63.410 43.300 63.730 ;
        RECT 45.860 63.640 46.000 69.870 ;
        RECT 46.780 69.170 46.920 71.230 ;
        RECT 46.260 68.850 46.520 69.170 ;
        RECT 46.720 68.850 46.980 69.170 ;
        RECT 46.320 66.790 46.460 68.850 ;
        RECT 47.640 68.510 47.900 68.830 ;
        RECT 46.260 66.470 46.520 66.790 ;
        RECT 47.700 65.770 47.840 68.510 ;
        RECT 50.000 66.450 50.140 73.610 ;
        RECT 50.400 71.910 50.660 72.230 ;
        RECT 51.320 71.910 51.580 72.230 ;
        RECT 50.460 69.850 50.600 71.910 ;
        RECT 50.400 69.530 50.660 69.850 ;
        RECT 50.460 67.130 50.600 69.530 ;
        RECT 51.380 69.510 51.520 71.910 ;
        RECT 51.320 69.190 51.580 69.510 ;
        RECT 52.300 69.170 52.440 77.690 ;
        RECT 54.600 76.990 54.740 80.410 ;
        RECT 55.980 80.390 56.120 82.110 ;
        RECT 57.360 82.090 57.500 85.170 ;
        RECT 57.300 81.770 57.560 82.090 ;
        RECT 55.920 80.070 56.180 80.390 ;
        RECT 57.360 80.050 57.500 81.770 ;
        RECT 57.300 79.730 57.560 80.050 ;
        RECT 57.820 79.710 57.960 102.510 ;
        RECT 58.740 102.490 58.880 115.770 ;
        RECT 58.680 102.170 58.940 102.490 ;
        RECT 59.140 101.490 59.400 101.810 ;
        RECT 59.200 98.750 59.340 101.490 ;
        RECT 59.660 98.830 59.800 122.570 ;
        RECT 61.040 112.690 61.180 126.310 ;
        RECT 61.960 121.530 62.100 128.690 ;
        RECT 62.420 128.670 62.560 130.730 ;
        RECT 62.360 128.350 62.620 128.670 ;
        RECT 63.800 126.290 63.940 130.730 ;
        RECT 63.740 125.970 64.000 126.290 ;
        RECT 66.100 125.950 66.240 131.410 ;
        RECT 67.480 127.310 67.620 137.335 ;
        RECT 67.940 134.020 68.080 144.670 ;
        RECT 68.340 134.020 68.600 134.110 ;
        RECT 67.940 133.880 68.600 134.020 ;
        RECT 67.940 129.010 68.080 133.880 ;
        RECT 68.340 133.790 68.600 133.880 ;
        RECT 67.880 128.690 68.140 129.010 ;
        RECT 67.880 128.010 68.140 128.330 ;
        RECT 67.420 126.990 67.680 127.310 ;
        RECT 67.940 126.630 68.080 128.010 ;
        RECT 67.880 126.310 68.140 126.630 ;
        RECT 66.040 125.630 66.300 125.950 ;
        RECT 62.360 123.930 62.620 124.250 ;
        RECT 61.900 121.210 62.160 121.530 ;
        RECT 62.420 116.390 62.560 123.930 ;
        RECT 69.780 123.310 69.920 163.370 ;
        RECT 70.170 159.095 70.450 159.465 ;
        RECT 70.240 153.490 70.380 159.095 ;
        RECT 70.700 158.930 70.840 164.050 ;
        RECT 71.620 163.690 71.760 169.410 ;
        RECT 72.300 168.275 73.840 168.645 ;
        RECT 72.020 166.090 72.280 166.410 ;
        RECT 72.080 164.710 72.220 166.090 ;
        RECT 72.020 164.390 72.280 164.710 ;
        RECT 71.560 163.370 71.820 163.690 ;
        RECT 72.300 162.835 73.840 163.205 ;
        RECT 70.640 158.610 70.900 158.930 ;
        RECT 70.180 153.170 70.440 153.490 ;
        RECT 70.170 143.455 70.450 143.825 ;
        RECT 70.180 143.310 70.440 143.455 ;
        RECT 70.700 143.030 70.840 158.610 ;
        RECT 71.100 157.930 71.360 158.250 ;
        RECT 71.160 156.210 71.300 157.930 ;
        RECT 72.300 157.395 73.840 157.765 ;
        RECT 71.100 155.890 71.360 156.210 ;
        RECT 74.840 154.510 74.980 174.590 ;
        RECT 75.760 172.530 75.900 175.270 ;
        RECT 75.700 172.210 75.960 172.530 ;
        RECT 76.620 172.210 76.880 172.530 ;
        RECT 76.680 169.470 76.820 172.210 ;
        RECT 77.140 169.810 77.280 185.810 ;
        RECT 78.520 184.430 78.660 186.490 ;
        RECT 80.300 186.150 80.560 186.470 ;
        RECT 79.380 185.130 79.640 185.450 ;
        RECT 78.460 184.110 78.720 184.430 ;
        RECT 79.440 181.370 79.580 185.130 ;
        RECT 80.360 181.710 80.500 186.150 ;
        RECT 80.300 181.390 80.560 181.710 ;
        RECT 79.380 181.050 79.640 181.370 ;
        RECT 78.460 174.590 78.720 174.910 ;
        RECT 77.080 169.490 77.340 169.810 ;
        RECT 77.540 169.490 77.800 169.810 ;
        RECT 76.620 169.150 76.880 169.470 ;
        RECT 76.680 168.020 76.820 169.150 ;
        RECT 76.680 167.880 77.280 168.020 ;
        RECT 76.620 167.110 76.880 167.430 ;
        RECT 76.160 166.090 76.420 166.410 ;
        RECT 76.220 164.905 76.360 166.090 ;
        RECT 76.150 164.535 76.430 164.905 ;
        RECT 76.680 164.710 76.820 167.110 ;
        RECT 76.620 164.390 76.880 164.710 ;
        RECT 75.230 163.855 75.510 164.225 ;
        RECT 75.300 161.310 75.440 163.855 ;
        RECT 76.160 163.370 76.420 163.690 ;
        RECT 76.220 161.650 76.360 163.370 ;
        RECT 76.680 162.670 76.820 164.390 ;
        RECT 76.620 162.350 76.880 162.670 ;
        RECT 77.140 161.650 77.280 167.880 ;
        RECT 77.600 167.430 77.740 169.490 ;
        RECT 78.520 169.130 78.660 174.590 ;
        RECT 78.920 171.870 79.180 172.190 ;
        RECT 79.380 171.870 79.640 172.190 ;
        RECT 78.980 170.490 79.120 171.870 ;
        RECT 78.920 170.170 79.180 170.490 ;
        RECT 79.440 170.150 79.580 171.870 ;
        RECT 80.300 171.530 80.560 171.850 ;
        RECT 80.360 170.150 80.500 171.530 ;
        RECT 79.380 169.830 79.640 170.150 ;
        RECT 80.300 169.830 80.560 170.150 ;
        RECT 80.820 169.550 80.960 199.070 ;
        RECT 79.900 169.410 80.960 169.550 ;
        RECT 78.460 168.810 78.720 169.130 ;
        RECT 78.920 168.810 79.180 169.130 ;
        RECT 77.540 167.110 77.800 167.430 ;
        RECT 77.600 164.690 77.740 167.110 ;
        RECT 78.980 166.750 79.120 168.810 ;
        RECT 79.380 166.770 79.640 167.090 ;
        RECT 78.920 166.430 79.180 166.750 ;
        RECT 77.600 164.550 78.660 164.690 ;
        RECT 77.540 162.010 77.800 162.330 ;
        RECT 76.160 161.330 76.420 161.650 ;
        RECT 77.080 161.330 77.340 161.650 ;
        RECT 75.240 160.990 75.500 161.310 ;
        RECT 77.600 160.880 77.740 162.010 ;
        RECT 77.140 160.740 77.740 160.880 ;
        RECT 77.140 159.270 77.280 160.740 ;
        RECT 77.080 158.950 77.340 159.270 ;
        RECT 76.620 158.610 76.880 158.930 ;
        RECT 76.680 157.230 76.820 158.610 ;
        RECT 76.620 156.910 76.880 157.230 ;
        RECT 74.780 154.190 75.040 154.510 ;
        RECT 77.140 154.420 77.280 158.950 ;
        RECT 78.520 158.930 78.660 164.550 ;
        RECT 78.920 164.390 79.180 164.710 ;
        RECT 78.980 161.990 79.120 164.390 ;
        RECT 78.920 161.670 79.180 161.990 ;
        RECT 79.440 161.310 79.580 166.770 ;
        RECT 79.380 160.990 79.640 161.310 ;
        RECT 79.440 159.610 79.580 160.990 ;
        RECT 79.380 159.290 79.640 159.610 ;
        RECT 78.460 158.610 78.720 158.930 ;
        RECT 79.900 156.745 80.040 169.410 ;
        RECT 81.280 167.430 81.420 201.450 ;
        RECT 82.660 200.410 82.800 202.130 ;
        RECT 82.600 200.090 82.860 200.410 ;
        RECT 81.680 199.750 81.940 200.070 ;
        RECT 81.740 170.150 81.880 199.750 ;
        RECT 82.140 186.150 82.400 186.470 ;
        RECT 82.200 171.850 82.340 186.150 ;
        RECT 83.120 183.750 83.260 202.130 ;
        RECT 85.360 199.070 85.620 199.390 ;
        RECT 84.900 197.030 85.160 197.350 ;
        RECT 84.960 195.310 85.100 197.030 ;
        RECT 84.900 194.990 85.160 195.310 ;
        RECT 85.420 194.290 85.560 199.070 ;
        RECT 85.360 193.970 85.620 194.290 ;
        RECT 83.520 193.290 83.780 193.610 ;
        RECT 83.580 192.250 83.720 193.290 ;
        RECT 83.520 191.930 83.780 192.250 ;
        RECT 84.900 190.570 85.160 190.890 ;
        RECT 83.980 188.870 84.240 189.190 ;
        RECT 83.520 187.850 83.780 188.170 ;
        RECT 83.580 186.470 83.720 187.850 ;
        RECT 83.520 186.150 83.780 186.470 ;
        RECT 83.060 183.430 83.320 183.750 ;
        RECT 84.040 183.410 84.180 188.870 ;
        RECT 84.960 188.850 85.100 190.570 ;
        RECT 84.440 188.530 84.700 188.850 ;
        RECT 84.900 188.530 85.160 188.850 ;
        RECT 83.980 183.090 84.240 183.410 ;
        RECT 84.040 180.430 84.180 183.090 ;
        RECT 83.580 180.290 84.180 180.430 ;
        RECT 83.580 180.010 83.720 180.290 ;
        RECT 83.520 179.690 83.780 180.010 ;
        RECT 83.060 177.310 83.320 177.630 ;
        RECT 83.120 176.270 83.260 177.310 ;
        RECT 83.060 175.950 83.320 176.270 ;
        RECT 83.520 175.950 83.780 176.270 ;
        RECT 82.590 172.015 82.870 172.385 ;
        RECT 82.140 171.530 82.400 171.850 ;
        RECT 82.660 170.490 82.800 172.015 ;
        RECT 83.580 170.830 83.720 175.950 ;
        RECT 84.500 173.550 84.640 188.530 ;
        RECT 84.900 187.850 85.160 188.170 ;
        RECT 84.960 186.470 85.100 187.850 ;
        RECT 84.900 186.150 85.160 186.470 ;
        RECT 84.900 182.410 85.160 182.730 ;
        RECT 84.960 181.370 85.100 182.410 ;
        RECT 84.900 181.050 85.160 181.370 ;
        RECT 85.880 176.180 86.020 204.170 ;
        RECT 87.720 203.130 87.860 204.170 ;
        RECT 87.660 202.810 87.920 203.130 ;
        RECT 86.740 201.450 87.000 201.770 ;
        RECT 86.800 199.730 86.940 201.450 ;
        RECT 88.180 200.070 88.320 206.890 ;
        RECT 88.580 204.850 88.840 205.170 ;
        RECT 88.120 199.750 88.380 200.070 ;
        RECT 86.740 199.410 87.000 199.730 ;
        RECT 86.280 198.730 86.540 199.050 ;
        RECT 86.340 196.330 86.480 198.730 ;
        RECT 86.280 196.010 86.540 196.330 ;
        RECT 86.800 195.310 86.940 199.410 ;
        RECT 88.640 198.030 88.780 204.850 ;
        RECT 90.020 204.830 90.160 206.890 ;
        RECT 89.960 204.510 90.220 204.830 ;
        RECT 89.090 203.635 90.630 204.005 ;
        RECT 89.090 198.195 90.630 198.565 ;
        RECT 88.580 197.710 88.840 198.030 ;
        RECT 89.500 196.690 89.760 197.010 ;
        RECT 89.560 195.310 89.700 196.690 ;
        RECT 86.740 194.990 87.000 195.310 ;
        RECT 89.500 194.990 89.760 195.310 ;
        RECT 86.800 191.910 86.940 194.990 ;
        RECT 88.120 193.630 88.380 193.950 ;
        RECT 88.180 191.910 88.320 193.630 ;
        RECT 89.090 192.755 90.630 193.125 ;
        RECT 86.740 191.590 87.000 191.910 ;
        RECT 88.120 191.590 88.380 191.910 ;
        RECT 89.040 190.570 89.300 190.890 ;
        RECT 89.100 188.850 89.240 190.570 ;
        RECT 89.040 188.530 89.300 188.850 ;
        RECT 86.740 188.190 87.000 188.510 ;
        RECT 86.800 178.310 86.940 188.190 ;
        RECT 89.090 187.315 90.630 187.685 ;
        RECT 90.940 186.665 91.080 207.910 ;
        RECT 108.880 207.210 109.020 207.910 ;
        RECT 93.640 206.890 93.900 207.210 ;
        RECT 103.760 206.890 104.020 207.210 ;
        RECT 107.900 206.890 108.160 207.210 ;
        RECT 108.820 207.120 109.080 207.210 ;
        RECT 108.420 206.980 109.080 207.120 ;
        RECT 92.720 204.170 92.980 204.490 ;
        RECT 92.780 203.470 92.920 204.170 ;
        RECT 92.720 203.150 92.980 203.470 ;
        RECT 92.780 202.790 92.920 203.150 ;
        RECT 92.720 202.470 92.980 202.790 ;
        RECT 93.700 200.070 93.840 206.890 ;
        RECT 100.080 205.530 100.340 205.850 ;
        RECT 96.860 204.850 97.120 205.170 ;
        RECT 96.920 203.470 97.060 204.850 ;
        RECT 95.480 203.150 95.740 203.470 ;
        RECT 96.860 203.150 97.120 203.470 ;
        RECT 93.640 199.750 93.900 200.070 ;
        RECT 93.180 197.030 93.440 197.350 ;
        RECT 91.340 196.010 91.600 196.330 ;
        RECT 91.400 191.910 91.540 196.010 ;
        RECT 93.240 195.310 93.380 197.030 ;
        RECT 93.180 194.990 93.440 195.310 ;
        RECT 92.260 193.630 92.520 193.950 ;
        RECT 92.320 192.590 92.460 193.630 ;
        RECT 92.260 192.270 92.520 192.590 ;
        RECT 91.340 191.590 91.600 191.910 ;
        RECT 91.340 188.530 91.600 188.850 ;
        RECT 91.400 187.150 91.540 188.530 ;
        RECT 91.340 186.830 91.600 187.150 ;
        RECT 90.870 186.295 91.150 186.665 ;
        RECT 93.700 186.470 93.840 199.750 ;
        RECT 95.540 196.330 95.680 203.150 ;
        RECT 95.940 202.870 96.200 203.130 ;
        RECT 95.940 202.810 97.060 202.870 ;
        RECT 96.000 202.730 97.060 202.810 ;
        RECT 96.920 202.450 97.060 202.730 ;
        RECT 95.940 202.130 96.200 202.450 ;
        RECT 96.860 202.130 97.120 202.450 ;
        RECT 96.000 198.030 96.140 202.130 ;
        RECT 96.400 201.790 96.660 202.110 ;
        RECT 96.460 199.730 96.600 201.790 ;
        RECT 96.400 199.410 96.660 199.730 ;
        RECT 95.940 197.710 96.200 198.030 ;
        RECT 96.000 197.010 96.140 197.710 ;
        RECT 96.920 197.010 97.060 202.130 ;
        RECT 98.240 201.450 98.500 201.770 ;
        RECT 98.300 200.750 98.440 201.450 ;
        RECT 98.240 200.430 98.500 200.750 ;
        RECT 100.140 199.730 100.280 205.530 ;
        RECT 100.540 204.850 100.800 205.170 ;
        RECT 100.600 203.470 100.740 204.850 ;
        RECT 100.540 203.150 100.800 203.470 ;
        RECT 103.820 203.130 103.960 206.890 ;
        RECT 105.880 206.355 107.420 206.725 ;
        RECT 104.220 204.510 104.480 204.830 ;
        RECT 103.760 202.810 104.020 203.130 ;
        RECT 104.280 202.110 104.420 204.510 ;
        RECT 107.960 202.790 108.100 206.890 ;
        RECT 107.900 202.470 108.160 202.790 ;
        RECT 102.840 201.790 103.100 202.110 ;
        RECT 104.220 201.790 104.480 202.110 ;
        RECT 102.900 199.730 103.040 201.790 ;
        RECT 103.300 200.430 103.560 200.750 ;
        RECT 97.320 199.410 97.580 199.730 ;
        RECT 100.080 199.410 100.340 199.730 ;
        RECT 102.840 199.410 103.100 199.730 ;
        RECT 97.380 197.350 97.520 199.410 ;
        RECT 99.160 199.070 99.420 199.390 ;
        RECT 99.220 197.690 99.360 199.070 ;
        RECT 101.460 198.730 101.720 199.050 ;
        RECT 101.520 198.030 101.660 198.730 ;
        RECT 101.460 197.710 101.720 198.030 ;
        RECT 102.900 197.690 103.040 199.410 ;
        RECT 103.360 199.390 103.500 200.430 ;
        RECT 103.760 199.410 104.020 199.730 ;
        RECT 103.300 199.070 103.560 199.390 ;
        RECT 99.160 197.370 99.420 197.690 ;
        RECT 102.840 197.370 103.100 197.690 ;
        RECT 97.320 197.030 97.580 197.350 ;
        RECT 98.700 197.030 98.960 197.350 ;
        RECT 95.940 196.690 96.200 197.010 ;
        RECT 96.860 196.690 97.120 197.010 ;
        RECT 95.480 196.010 95.740 196.330 ;
        RECT 95.540 191.910 95.680 196.010 ;
        RECT 97.380 191.910 97.520 197.030 ;
        RECT 98.240 193.970 98.500 194.290 ;
        RECT 98.300 192.590 98.440 193.970 ;
        RECT 98.240 192.270 98.500 192.590 ;
        RECT 95.480 191.590 95.740 191.910 ;
        RECT 97.320 191.590 97.580 191.910 ;
        RECT 94.560 190.570 94.820 190.890 ;
        RECT 98.240 190.570 98.500 190.890 ;
        RECT 94.620 188.850 94.760 190.570 ;
        RECT 97.780 189.210 98.040 189.530 ;
        RECT 97.840 188.850 97.980 189.210 ;
        RECT 98.300 188.850 98.440 190.570 ;
        RECT 94.100 188.530 94.360 188.850 ;
        RECT 94.560 188.530 94.820 188.850 ;
        RECT 97.780 188.530 98.040 188.850 ;
        RECT 98.240 188.530 98.500 188.850 ;
        RECT 88.120 182.750 88.380 183.070 ;
        RECT 88.180 181.710 88.320 182.750 ;
        RECT 89.090 181.875 90.630 182.245 ;
        RECT 88.120 181.390 88.380 181.710 ;
        RECT 89.960 180.710 90.220 181.030 ;
        RECT 86.740 177.990 87.000 178.310 ;
        RECT 86.800 177.290 86.940 177.990 ;
        RECT 90.020 177.970 90.160 180.710 ;
        RECT 89.960 177.650 90.220 177.970 ;
        RECT 86.740 176.970 87.000 177.290 ;
        RECT 87.200 176.970 87.460 177.290 ;
        RECT 85.880 176.040 86.480 176.180 ;
        RECT 85.360 175.270 85.620 175.590 ;
        RECT 84.900 174.250 85.160 174.570 ;
        RECT 84.440 173.230 84.700 173.550 ;
        RECT 83.980 172.210 84.240 172.530 ;
        RECT 83.520 170.510 83.780 170.830 ;
        RECT 82.600 170.170 82.860 170.490 ;
        RECT 81.680 169.830 81.940 170.150 ;
        RECT 81.680 169.150 81.940 169.470 ;
        RECT 81.220 167.110 81.480 167.430 ;
        RECT 81.280 164.710 81.420 167.110 ;
        RECT 81.740 165.050 81.880 169.150 ;
        RECT 81.680 164.730 81.940 165.050 ;
        RECT 81.220 164.620 81.480 164.710 ;
        RECT 80.820 164.480 81.480 164.620 ;
        RECT 80.300 161.670 80.560 161.990 ;
        RECT 80.360 158.250 80.500 161.670 ;
        RECT 80.820 161.650 80.960 164.480 ;
        RECT 81.220 164.390 81.480 164.480 ;
        RECT 81.680 164.050 81.940 164.370 ;
        RECT 81.220 163.370 81.480 163.690 ;
        RECT 80.760 161.330 81.020 161.650 ;
        RECT 80.820 159.610 80.960 161.330 ;
        RECT 80.760 159.290 81.020 159.610 ;
        RECT 80.300 157.930 80.560 158.250 ;
        RECT 79.830 156.375 80.110 156.745 ;
        RECT 76.680 154.280 77.280 154.420 ;
        RECT 74.320 153.170 74.580 153.490 ;
        RECT 72.300 151.955 73.840 152.325 ;
        RECT 72.300 146.515 73.840 146.885 ;
        RECT 70.240 142.890 70.840 143.030 ;
        RECT 70.240 124.250 70.380 142.890 ;
        RECT 71.100 142.630 71.360 142.950 ;
        RECT 70.640 138.890 70.900 139.210 ;
        RECT 70.700 138.190 70.840 138.890 ;
        RECT 71.160 138.190 71.300 142.630 ;
        RECT 72.300 141.075 73.840 141.445 ;
        RECT 71.560 138.890 71.820 139.210 ;
        RECT 73.400 138.890 73.660 139.210 ;
        RECT 70.640 137.870 70.900 138.190 ;
        RECT 71.100 137.870 71.360 138.190 ;
        RECT 71.620 137.510 71.760 138.890 ;
        RECT 73.460 137.850 73.600 138.890 ;
        RECT 73.400 137.530 73.660 137.850 ;
        RECT 71.560 137.190 71.820 137.510 ;
        RECT 71.620 132.750 71.760 137.190 ;
        RECT 72.300 135.635 73.840 136.005 ;
        RECT 71.560 132.430 71.820 132.750 ;
        RECT 72.300 130.195 73.840 130.565 ;
        RECT 72.300 124.755 73.840 125.125 ;
        RECT 74.380 124.590 74.520 153.170 ;
        RECT 75.240 150.110 75.500 150.430 ;
        RECT 75.300 149.070 75.440 150.110 ;
        RECT 75.240 148.750 75.500 149.070 ;
        RECT 75.240 147.730 75.500 148.050 ;
        RECT 75.300 147.370 75.440 147.730 ;
        RECT 75.240 147.050 75.500 147.370 ;
        RECT 74.780 144.670 75.040 144.990 ;
        RECT 74.840 143.630 74.980 144.670 ;
        RECT 74.780 143.310 75.040 143.630 ;
        RECT 75.300 139.890 75.440 147.050 ;
        RECT 76.160 145.010 76.420 145.330 ;
        RECT 75.700 144.670 75.960 144.990 ;
        RECT 75.760 142.950 75.900 144.670 ;
        RECT 75.700 142.630 75.960 142.950 ;
        RECT 76.220 142.350 76.360 145.010 ;
        RECT 75.760 142.270 76.360 142.350 ;
        RECT 75.700 142.210 76.360 142.270 ;
        RECT 75.700 141.950 75.960 142.210 ;
        RECT 75.240 139.570 75.500 139.890 ;
        RECT 75.760 137.170 75.900 141.950 ;
        RECT 76.680 138.190 76.820 154.280 ;
        RECT 77.080 153.510 77.340 153.830 ;
        RECT 77.140 148.390 77.280 153.510 ;
        RECT 80.300 152.830 80.560 153.150 ;
        RECT 78.460 152.490 78.720 152.810 ;
        RECT 77.540 150.450 77.800 150.770 ;
        RECT 77.600 148.730 77.740 150.450 ;
        RECT 77.540 148.410 77.800 148.730 ;
        RECT 78.520 148.390 78.660 152.490 ;
        RECT 77.080 148.070 77.340 148.390 ;
        RECT 78.460 148.070 78.720 148.390 ;
        RECT 78.000 147.390 78.260 147.710 ;
        RECT 77.080 144.330 77.340 144.650 ;
        RECT 77.140 142.950 77.280 144.330 ;
        RECT 77.080 142.630 77.340 142.950 ;
        RECT 77.540 142.860 77.800 142.950 ;
        RECT 78.060 142.860 78.200 147.390 ;
        RECT 80.360 145.330 80.500 152.830 ;
        RECT 81.280 151.190 81.420 163.370 ;
        RECT 81.740 161.310 81.880 164.050 ;
        RECT 81.680 160.990 81.940 161.310 ;
        RECT 82.660 160.970 82.800 170.170 ;
        RECT 84.040 166.410 84.180 172.210 ;
        RECT 84.440 169.830 84.700 170.150 ;
        RECT 84.500 167.430 84.640 169.830 ;
        RECT 84.960 169.550 85.100 174.250 ;
        RECT 85.420 171.850 85.560 175.270 ;
        RECT 86.340 172.385 86.480 176.040 ;
        RECT 87.260 175.930 87.400 176.970 ;
        RECT 89.090 176.435 90.630 176.805 ;
        RECT 90.940 176.270 91.080 186.295 ;
        RECT 93.640 186.150 93.900 186.470 ;
        RECT 94.160 184.430 94.300 188.530 ;
        RECT 96.850 185.615 97.130 185.985 ;
        RECT 94.100 184.110 94.360 184.430 ;
        RECT 94.160 183.750 94.300 184.110 ;
        RECT 94.100 183.430 94.360 183.750 ;
        RECT 95.020 182.410 95.280 182.730 ;
        RECT 95.080 181.710 95.220 182.410 ;
        RECT 95.020 181.390 95.280 181.710 ;
        RECT 94.560 180.710 94.820 181.030 ;
        RECT 92.720 178.670 92.980 178.990 ;
        RECT 92.260 177.650 92.520 177.970 ;
        RECT 90.880 175.950 91.140 176.270 ;
        RECT 87.200 175.610 87.460 175.930 ;
        RECT 88.580 174.250 88.840 174.570 ;
        RECT 88.640 173.550 88.780 174.250 ;
        RECT 88.580 173.230 88.840 173.550 ;
        RECT 90.880 172.890 91.140 173.210 ;
        RECT 86.270 172.015 86.550 172.385 ;
        RECT 86.740 172.210 87.000 172.530 ;
        RECT 85.360 171.530 85.620 171.850 ;
        RECT 84.960 169.410 85.560 169.550 ;
        RECT 84.900 168.810 85.160 169.130 ;
        RECT 84.960 167.770 85.100 168.810 ;
        RECT 84.900 167.450 85.160 167.770 ;
        RECT 84.440 167.110 84.700 167.430 ;
        RECT 83.980 166.090 84.240 166.410 ;
        RECT 84.500 164.690 84.640 167.110 ;
        RECT 84.900 166.770 85.160 167.090 ;
        RECT 83.580 164.550 84.640 164.690 ;
        RECT 82.600 160.650 82.860 160.970 ;
        RECT 82.140 157.930 82.400 158.250 ;
        RECT 82.200 154.170 82.340 157.930 ;
        RECT 83.060 155.210 83.320 155.530 ;
        RECT 82.600 154.190 82.860 154.510 ;
        RECT 82.140 153.850 82.400 154.170 ;
        RECT 81.680 153.510 81.940 153.830 ;
        RECT 80.820 151.050 81.420 151.190 ;
        RECT 80.300 145.010 80.560 145.330 ;
        RECT 80.300 144.330 80.560 144.650 ;
        RECT 80.360 143.630 80.500 144.330 ;
        RECT 80.300 143.310 80.560 143.630 ;
        RECT 77.540 142.720 78.200 142.860 ;
        RECT 77.540 142.630 77.800 142.720 ;
        RECT 77.140 140.230 77.280 142.630 ;
        RECT 77.080 139.910 77.340 140.230 ;
        RECT 76.620 137.870 76.880 138.190 ;
        RECT 77.080 137.190 77.340 137.510 ;
        RECT 75.700 136.850 75.960 137.170 ;
        RECT 75.240 136.170 75.500 136.490 ;
        RECT 75.300 135.470 75.440 136.170 ;
        RECT 75.240 135.150 75.500 135.470 ;
        RECT 75.760 129.010 75.900 136.850 ;
        RECT 76.160 133.450 76.420 133.770 ;
        RECT 76.220 132.070 76.360 133.450 ;
        RECT 77.140 132.750 77.280 137.190 ;
        RECT 77.080 132.430 77.340 132.750 ;
        RECT 76.160 131.750 76.420 132.070 ;
        RECT 77.600 131.730 77.740 142.630 ;
        RECT 79.380 142.290 79.640 142.610 ;
        RECT 79.440 134.450 79.580 142.290 ;
        RECT 79.380 134.130 79.640 134.450 ;
        RECT 76.620 131.410 76.880 131.730 ;
        RECT 77.540 131.410 77.800 131.730 ;
        RECT 76.150 129.855 76.430 130.225 ;
        RECT 75.700 128.690 75.960 129.010 ;
        RECT 76.220 126.630 76.360 129.855 ;
        RECT 76.680 126.970 76.820 131.410 ;
        RECT 80.820 128.670 80.960 151.050 ;
        RECT 81.220 150.110 81.480 150.430 ;
        RECT 81.280 148.730 81.420 150.110 ;
        RECT 81.220 148.410 81.480 148.730 ;
        RECT 81.740 129.350 81.880 153.510 ;
        RECT 82.140 152.490 82.400 152.810 ;
        RECT 82.200 148.390 82.340 152.490 ;
        RECT 82.140 148.070 82.400 148.390 ;
        RECT 82.140 142.630 82.400 142.950 ;
        RECT 82.200 140.910 82.340 142.630 ;
        RECT 82.140 140.590 82.400 140.910 ;
        RECT 82.660 139.210 82.800 154.190 ;
        RECT 83.120 148.390 83.260 155.210 ;
        RECT 83.580 153.490 83.720 164.550 ;
        RECT 84.960 159.270 85.100 166.770 ;
        RECT 85.420 164.690 85.560 169.410 ;
        RECT 85.820 168.810 86.080 169.130 ;
        RECT 85.880 167.090 86.020 168.810 ;
        RECT 85.820 166.770 86.080 167.090 ;
        RECT 86.280 166.770 86.540 167.090 ;
        RECT 85.420 164.550 86.020 164.690 ;
        RECT 85.360 160.650 85.620 160.970 ;
        RECT 85.420 159.270 85.560 160.650 ;
        RECT 84.900 158.950 85.160 159.270 ;
        RECT 85.360 158.950 85.620 159.270 ;
        RECT 83.980 153.850 84.240 154.170 ;
        RECT 83.520 153.170 83.780 153.490 ;
        RECT 84.040 150.090 84.180 153.850 ;
        RECT 84.440 153.170 84.700 153.490 ;
        RECT 84.500 151.790 84.640 153.170 ;
        RECT 85.880 152.810 86.020 164.550 ;
        RECT 86.340 163.690 86.480 166.770 ;
        RECT 86.800 166.750 86.940 172.210 ;
        RECT 89.090 170.995 90.630 171.365 ;
        RECT 88.580 170.510 88.840 170.830 ;
        RECT 86.740 166.430 87.000 166.750 ;
        RECT 86.800 165.390 86.940 166.430 ;
        RECT 86.740 165.070 87.000 165.390 ;
        RECT 86.740 164.050 87.000 164.370 ;
        RECT 86.280 163.370 86.540 163.690 ;
        RECT 86.800 159.270 86.940 164.050 ;
        RECT 87.200 163.710 87.460 164.030 ;
        RECT 87.260 161.505 87.400 163.710 ;
        RECT 88.640 163.690 88.780 170.510 ;
        RECT 90.940 170.490 91.080 172.890 ;
        RECT 91.340 172.210 91.600 172.530 ;
        RECT 90.880 170.170 91.140 170.490 ;
        RECT 91.400 168.110 91.540 172.210 ;
        RECT 92.320 171.850 92.460 177.650 ;
        RECT 92.780 173.550 92.920 178.670 ;
        RECT 93.180 177.650 93.440 177.970 ;
        RECT 93.240 173.550 93.380 177.650 ;
        RECT 94.100 176.970 94.360 177.290 ;
        RECT 94.160 175.590 94.300 176.970 ;
        RECT 94.100 175.270 94.360 175.590 ;
        RECT 92.720 173.230 92.980 173.550 ;
        RECT 93.180 173.230 93.440 173.550 ;
        RECT 92.260 171.530 92.520 171.850 ;
        RECT 91.800 169.830 92.060 170.150 ;
        RECT 91.340 167.790 91.600 168.110 ;
        RECT 89.090 165.555 90.630 165.925 ;
        RECT 90.880 164.730 91.140 165.050 ;
        RECT 88.580 163.370 88.840 163.690 ;
        RECT 88.640 162.670 88.780 163.370 ;
        RECT 88.580 162.350 88.840 162.670 ;
        RECT 88.580 161.670 88.840 161.990 ;
        RECT 87.190 161.135 87.470 161.505 ;
        RECT 86.740 158.950 87.000 159.270 ;
        RECT 86.800 156.550 86.940 158.950 ;
        RECT 86.740 156.230 87.000 156.550 ;
        RECT 85.820 152.490 86.080 152.810 ;
        RECT 85.880 151.790 86.020 152.490 ;
        RECT 84.440 151.470 84.700 151.790 ;
        RECT 85.820 151.470 86.080 151.790 ;
        RECT 83.980 149.770 84.240 150.090 ;
        RECT 83.060 148.070 83.320 148.390 ;
        RECT 84.040 144.990 84.180 149.770 ;
        RECT 85.360 148.070 85.620 148.390 ;
        RECT 83.980 144.670 84.240 144.990 ;
        RECT 83.520 139.230 83.780 139.550 ;
        RECT 82.600 138.890 82.860 139.210 ;
        RECT 83.580 137.850 83.720 139.230 ;
        RECT 84.040 138.190 84.180 144.670 ;
        RECT 85.420 139.890 85.560 148.070 ;
        RECT 85.880 146.350 86.020 151.470 ;
        RECT 86.800 150.770 86.940 156.230 ;
        RECT 86.740 150.450 87.000 150.770 ;
        RECT 86.740 149.770 87.000 150.090 ;
        RECT 86.800 148.390 86.940 149.770 ;
        RECT 87.260 148.730 87.400 161.135 ;
        RECT 88.120 158.950 88.380 159.270 ;
        RECT 87.660 157.930 87.920 158.250 ;
        RECT 87.720 156.210 87.860 157.930 ;
        RECT 88.180 157.230 88.320 158.950 ;
        RECT 88.640 158.250 88.780 161.670 ;
        RECT 89.090 160.115 90.630 160.485 ;
        RECT 88.580 157.930 88.840 158.250 ;
        RECT 88.120 156.910 88.380 157.230 ;
        RECT 87.660 155.890 87.920 156.210 ;
        RECT 88.120 153.170 88.380 153.490 ;
        RECT 87.660 149.770 87.920 150.090 ;
        RECT 87.720 148.730 87.860 149.770 ;
        RECT 87.200 148.410 87.460 148.730 ;
        RECT 87.660 148.410 87.920 148.730 ;
        RECT 88.180 148.390 88.320 153.170 ;
        RECT 86.740 148.070 87.000 148.390 ;
        RECT 88.120 148.070 88.380 148.390 ;
        RECT 85.820 146.030 86.080 146.350 ;
        RECT 85.360 139.570 85.620 139.890 ;
        RECT 83.980 137.870 84.240 138.190 ;
        RECT 83.520 137.530 83.780 137.850 ;
        RECT 83.060 136.170 83.320 136.490 ;
        RECT 82.140 133.790 82.400 134.110 ;
        RECT 82.200 132.750 82.340 133.790 ;
        RECT 82.140 132.430 82.400 132.750 ;
        RECT 83.120 132.070 83.260 136.170 ;
        RECT 82.140 131.750 82.400 132.070 ;
        RECT 83.060 131.750 83.320 132.070 ;
        RECT 84.900 131.980 85.160 132.070 ;
        RECT 85.420 131.980 85.560 139.570 ;
        RECT 85.880 136.490 86.020 146.030 ;
        RECT 86.740 145.010 87.000 145.330 ;
        RECT 86.800 143.630 86.940 145.010 ;
        RECT 88.120 144.330 88.380 144.650 ;
        RECT 86.740 143.310 87.000 143.630 ;
        RECT 88.180 140.230 88.320 144.330 ;
        RECT 88.120 139.910 88.380 140.230 ;
        RECT 87.660 139.570 87.920 139.890 ;
        RECT 87.200 138.890 87.460 139.210 ;
        RECT 85.820 136.170 86.080 136.490 ;
        RECT 85.880 135.470 86.020 136.170 ;
        RECT 85.820 135.150 86.080 135.470 ;
        RECT 86.740 133.450 87.000 133.770 ;
        RECT 86.800 132.070 86.940 133.450 ;
        RECT 84.900 131.840 85.560 131.980 ;
        RECT 84.900 131.750 85.160 131.840 ;
        RECT 86.740 131.750 87.000 132.070 ;
        RECT 81.680 129.030 81.940 129.350 ;
        RECT 80.760 128.350 81.020 128.670 ;
        RECT 78.460 128.010 78.720 128.330 ;
        RECT 76.620 126.650 76.880 126.970 ;
        RECT 78.520 126.630 78.660 128.010 ;
        RECT 76.160 126.310 76.420 126.630 ;
        RECT 78.460 126.310 78.720 126.630 ;
        RECT 79.380 126.310 79.640 126.630 ;
        RECT 80.300 126.310 80.560 126.630 ;
        RECT 74.320 124.270 74.580 124.590 ;
        RECT 70.180 123.930 70.440 124.250 ;
        RECT 69.780 123.170 70.380 123.310 ;
        RECT 64.660 122.570 64.920 122.890 ;
        RECT 69.720 122.570 69.980 122.890 ;
        RECT 64.720 120.510 64.860 122.570 ;
        RECT 69.780 121.190 69.920 122.570 ;
        RECT 67.880 120.870 68.140 121.190 ;
        RECT 69.260 120.870 69.520 121.190 ;
        RECT 69.720 120.870 69.980 121.190 ;
        RECT 64.660 120.190 64.920 120.510 ;
        RECT 64.720 118.470 64.860 120.190 ;
        RECT 66.500 119.850 66.760 120.170 ;
        RECT 66.560 118.470 66.700 119.850 ;
        RECT 67.940 118.810 68.080 120.870 ;
        RECT 67.880 118.490 68.140 118.810 ;
        RECT 68.340 118.490 68.600 118.810 ;
        RECT 64.660 118.150 64.920 118.470 ;
        RECT 66.500 118.150 66.760 118.470 ;
        RECT 67.420 118.150 67.680 118.470 ;
        RECT 64.200 117.470 64.460 117.790 ;
        RECT 62.420 116.250 63.020 116.390 ;
        RECT 60.980 112.370 61.240 112.690 ;
        RECT 61.040 109.970 61.180 112.370 ;
        RECT 60.980 109.650 61.240 109.970 ;
        RECT 60.060 104.210 60.320 104.530 ;
        RECT 60.120 99.430 60.260 104.210 ;
        RECT 62.360 103.870 62.620 104.190 ;
        RECT 61.900 103.530 62.160 103.850 ;
        RECT 60.060 99.110 60.320 99.430 ;
        RECT 59.140 98.430 59.400 98.750 ;
        RECT 59.660 98.690 60.260 98.830 ;
        RECT 60.120 95.690 60.260 98.690 ;
        RECT 61.440 98.090 61.700 98.410 ;
        RECT 60.060 95.370 60.320 95.690 ;
        RECT 60.120 91.610 60.260 95.370 ;
        RECT 60.520 92.650 60.780 92.970 ;
        RECT 60.980 92.650 61.240 92.970 ;
        RECT 60.060 91.290 60.320 91.610 ;
        RECT 58.220 90.950 58.480 91.270 ;
        RECT 58.280 89.230 58.420 90.950 ;
        RECT 58.680 90.270 58.940 90.590 ;
        RECT 58.220 88.910 58.480 89.230 ;
        RECT 58.740 87.530 58.880 90.270 ;
        RECT 59.140 89.930 59.400 90.250 ;
        RECT 59.200 87.870 59.340 89.930 ;
        RECT 59.140 87.550 59.400 87.870 ;
        RECT 58.680 87.210 58.940 87.530 ;
        RECT 59.200 86.590 59.340 87.550 ;
        RECT 58.740 86.450 59.340 86.590 ;
        RECT 58.740 84.810 58.880 86.450 ;
        RECT 60.580 85.490 60.720 92.650 ;
        RECT 61.040 90.930 61.180 92.650 ;
        RECT 60.980 90.610 61.240 90.930 ;
        RECT 60.520 85.170 60.780 85.490 ;
        RECT 58.680 84.490 58.940 84.810 ;
        RECT 59.600 84.490 59.860 84.810 ;
        RECT 58.740 81.070 58.880 84.490 ;
        RECT 58.680 80.750 58.940 81.070 ;
        RECT 59.140 80.410 59.400 80.730 ;
        RECT 55.000 79.390 55.260 79.710 ;
        RECT 57.760 79.390 58.020 79.710 ;
        RECT 54.540 76.670 54.800 76.990 ;
        RECT 55.060 74.610 55.200 79.390 ;
        RECT 55.510 78.515 57.050 78.885 ;
        RECT 58.680 78.030 58.940 78.350 ;
        RECT 57.760 77.350 58.020 77.670 ;
        RECT 55.460 76.670 55.720 76.990 ;
        RECT 55.000 74.290 55.260 74.610 ;
        RECT 54.540 73.950 54.800 74.270 ;
        RECT 54.080 71.910 54.340 72.230 ;
        RECT 52.700 71.570 52.960 71.890 ;
        RECT 52.240 68.850 52.500 69.170 ;
        RECT 50.400 66.810 50.660 67.130 ;
        RECT 50.860 66.470 51.120 66.790 ;
        RECT 49.940 66.130 50.200 66.450 ;
        RECT 47.640 65.450 47.900 65.770 ;
        RECT 49.480 65.450 49.740 65.770 ;
        RECT 46.260 63.640 46.520 63.730 ;
        RECT 45.860 63.500 46.520 63.640 ;
        RECT 46.260 63.410 46.520 63.500 ;
        RECT 41.260 58.630 41.400 63.410 ;
        RECT 47.180 63.070 47.440 63.390 ;
        RECT 42.580 62.730 42.840 63.050 ;
        RECT 43.960 62.730 44.220 63.050 ;
        RECT 42.120 61.030 42.380 61.350 ;
        RECT 40.740 58.310 41.000 58.630 ;
        RECT 41.200 58.310 41.460 58.630 ;
        RECT 42.180 57.350 42.320 61.030 ;
        RECT 42.640 58.290 42.780 62.730 ;
        RECT 44.020 61.350 44.160 62.730 ;
        RECT 43.960 61.030 44.220 61.350 ;
        RECT 47.240 61.010 47.380 63.070 ;
        RECT 48.100 61.030 48.360 61.350 ;
        RECT 47.180 60.690 47.440 61.010 ;
        RECT 47.180 60.010 47.440 60.330 ;
        RECT 47.240 59.310 47.380 60.010 ;
        RECT 47.180 58.990 47.440 59.310 ;
        RECT 42.580 57.970 42.840 58.290 ;
        RECT 45.340 57.970 45.600 58.290 ;
        RECT 42.180 57.210 42.780 57.350 ;
        RECT 39.420 56.530 40.020 56.670 ;
        RECT 39.420 55.990 39.560 56.530 ;
        RECT 39.880 56.220 40.020 56.530 ;
        RECT 42.640 56.220 42.780 57.210 ;
        RECT 45.400 56.220 45.540 57.970 ;
        RECT 48.160 56.220 48.300 61.030 ;
        RECT 49.540 58.290 49.680 65.450 ;
        RECT 50.000 64.750 50.140 66.130 ;
        RECT 49.940 64.430 50.200 64.750 ;
        RECT 49.480 57.970 49.740 58.290 ;
        RECT 50.920 56.220 51.060 66.470 ;
        RECT 51.320 65.450 51.580 65.770 ;
        RECT 51.380 64.070 51.520 65.450 ;
        RECT 51.320 63.750 51.580 64.070 ;
        RECT 52.760 63.730 52.900 71.570 ;
        RECT 54.140 70.190 54.280 71.910 ;
        RECT 54.080 69.870 54.340 70.190 ;
        RECT 54.140 67.130 54.280 69.870 ;
        RECT 54.600 69.170 54.740 73.950 ;
        RECT 55.520 73.840 55.660 76.670 ;
        RECT 57.820 75.630 57.960 77.350 ;
        RECT 57.760 75.310 58.020 75.630 ;
        RECT 58.220 74.290 58.480 74.610 ;
        RECT 55.060 73.700 55.660 73.840 ;
        RECT 55.060 72.570 55.200 73.700 ;
        RECT 57.760 73.610 58.020 73.930 ;
        RECT 55.510 73.075 57.050 73.445 ;
        RECT 55.000 72.250 55.260 72.570 ;
        RECT 57.820 71.630 57.960 73.610 ;
        RECT 58.280 72.230 58.420 74.290 ;
        RECT 58.220 71.910 58.480 72.230 ;
        RECT 56.440 71.550 57.960 71.630 ;
        RECT 56.380 71.490 57.960 71.550 ;
        RECT 56.380 71.230 56.640 71.490 ;
        RECT 54.540 68.850 54.800 69.170 ;
        RECT 54.600 67.130 54.740 68.850 ;
        RECT 55.510 67.635 57.050 68.005 ;
        RECT 54.080 66.810 54.340 67.130 ;
        RECT 54.540 66.810 54.800 67.130 ;
        RECT 57.820 66.790 57.960 71.490 ;
        RECT 58.740 69.170 58.880 78.030 ;
        RECT 59.200 74.610 59.340 80.410 ;
        RECT 59.660 80.050 59.800 84.490 ;
        RECT 60.980 82.790 61.240 83.110 ;
        RECT 61.040 81.070 61.180 82.790 ;
        RECT 60.980 80.750 61.240 81.070 ;
        RECT 61.500 80.730 61.640 98.090 ;
        RECT 61.440 80.410 61.700 80.730 ;
        RECT 59.600 79.730 59.860 80.050 ;
        RECT 61.440 78.260 61.700 78.350 ;
        RECT 61.960 78.260 62.100 103.530 ;
        RECT 62.420 97.050 62.560 103.870 ;
        RECT 62.360 96.730 62.620 97.050 ;
        RECT 62.880 91.350 63.020 116.250 ;
        RECT 64.260 110.650 64.400 117.470 ;
        RECT 65.580 114.410 65.840 114.730 ;
        RECT 65.640 110.990 65.780 114.410 ;
        RECT 66.960 111.690 67.220 112.010 ;
        RECT 65.580 110.670 65.840 110.990 ;
        RECT 64.200 110.330 64.460 110.650 ;
        RECT 64.660 109.310 64.920 109.630 ;
        RECT 64.720 107.250 64.860 109.310 ;
        RECT 65.640 109.290 65.780 110.670 ;
        RECT 66.040 109.650 66.300 109.970 ;
        RECT 65.580 108.970 65.840 109.290 ;
        RECT 65.640 107.250 65.780 108.970 ;
        RECT 66.100 107.250 66.240 109.650 ;
        RECT 66.500 108.970 66.760 109.290 ;
        RECT 66.560 107.250 66.700 108.970 ;
        RECT 64.660 106.930 64.920 107.250 ;
        RECT 65.580 106.930 65.840 107.250 ;
        RECT 66.040 106.930 66.300 107.250 ;
        RECT 66.500 106.930 66.760 107.250 ;
        RECT 64.200 106.250 64.460 106.570 ;
        RECT 64.660 106.250 64.920 106.570 ;
        RECT 63.280 104.550 63.540 104.870 ;
        RECT 63.340 101.130 63.480 104.550 ;
        RECT 63.740 104.210 64.000 104.530 ;
        RECT 63.800 101.810 63.940 104.210 ;
        RECT 63.740 101.490 64.000 101.810 ;
        RECT 63.280 100.810 63.540 101.130 ;
        RECT 63.340 99.090 63.480 100.810 ;
        RECT 63.280 98.770 63.540 99.090 ;
        RECT 64.260 93.900 64.400 106.250 ;
        RECT 64.720 104.870 64.860 106.250 ;
        RECT 65.640 104.870 65.780 106.930 ;
        RECT 64.660 104.550 64.920 104.870 ;
        RECT 65.580 104.550 65.840 104.870 ;
        RECT 65.120 103.530 65.380 103.850 ;
        RECT 64.660 100.810 64.920 101.130 ;
        RECT 63.800 93.760 64.400 93.900 ;
        RECT 62.880 91.210 63.480 91.350 ;
        RECT 62.820 90.270 63.080 90.590 ;
        RECT 62.880 78.350 63.020 90.270 ;
        RECT 63.340 88.890 63.480 91.210 ;
        RECT 63.280 88.570 63.540 88.890 ;
        RECT 63.340 85.150 63.480 88.570 ;
        RECT 63.280 84.830 63.540 85.150 ;
        RECT 61.440 78.120 62.100 78.260 ;
        RECT 61.440 78.030 61.700 78.120 ;
        RECT 62.820 78.030 63.080 78.350 ;
        RECT 63.800 74.610 63.940 93.760 ;
        RECT 64.200 92.990 64.460 93.310 ;
        RECT 64.260 91.610 64.400 92.990 ;
        RECT 64.200 91.290 64.460 91.610 ;
        RECT 64.200 82.790 64.460 83.110 ;
        RECT 64.260 81.070 64.400 82.790 ;
        RECT 64.200 80.750 64.460 81.070 ;
        RECT 59.140 74.290 59.400 74.610 ;
        RECT 60.060 74.290 60.320 74.610 ;
        RECT 60.520 74.290 60.780 74.610 ;
        RECT 63.740 74.290 64.000 74.610 ;
        RECT 64.720 74.520 64.860 100.810 ;
        RECT 65.180 99.430 65.320 103.530 ;
        RECT 65.640 101.810 65.780 104.550 ;
        RECT 66.040 104.440 66.300 104.530 ;
        RECT 66.560 104.440 66.700 106.930 ;
        RECT 67.020 104.950 67.160 111.690 ;
        RECT 67.480 107.250 67.620 118.150 ;
        RECT 68.400 117.790 68.540 118.490 ;
        RECT 69.320 118.470 69.460 120.870 ;
        RECT 69.260 118.150 69.520 118.470 ;
        RECT 68.340 117.470 68.600 117.790 ;
        RECT 68.400 116.390 68.540 117.470 ;
        RECT 68.800 117.130 69.060 117.450 ;
        RECT 67.940 116.250 68.540 116.390 ;
        RECT 67.940 116.090 68.080 116.250 ;
        RECT 68.860 116.090 69.000 117.130 ;
        RECT 67.880 115.770 68.140 116.090 ;
        RECT 68.800 115.770 69.060 116.090 ;
        RECT 67.880 115.090 68.140 115.410 ;
        RECT 67.940 113.710 68.080 115.090 ;
        RECT 67.880 113.390 68.140 113.710 ;
        RECT 67.940 110.650 68.080 113.390 ;
        RECT 67.880 110.330 68.140 110.650 ;
        RECT 68.860 109.630 69.000 115.770 ;
        RECT 69.320 110.310 69.460 118.150 ;
        RECT 69.780 116.390 69.920 120.870 ;
        RECT 70.240 118.810 70.380 123.170 ;
        RECT 71.560 122.910 71.820 123.230 ;
        RECT 71.620 119.150 71.760 122.910 ;
        RECT 74.380 121.190 74.520 124.270 ;
        RECT 74.780 123.250 75.040 123.570 ;
        RECT 74.320 120.870 74.580 121.190 ;
        RECT 74.320 119.850 74.580 120.170 ;
        RECT 72.300 119.315 73.840 119.685 ;
        RECT 74.380 119.150 74.520 119.850 ;
        RECT 71.560 118.830 71.820 119.150 ;
        RECT 74.320 118.830 74.580 119.150 ;
        RECT 70.180 118.490 70.440 118.810 ;
        RECT 73.860 118.490 74.120 118.810 ;
        RECT 73.920 117.790 74.060 118.490 ;
        RECT 73.860 117.470 74.120 117.790 ;
        RECT 74.840 117.450 74.980 123.250 ;
        RECT 71.560 117.130 71.820 117.450 ;
        RECT 74.780 117.130 75.040 117.450 ;
        RECT 69.780 116.250 70.380 116.390 ;
        RECT 69.720 115.770 69.980 116.090 ;
        RECT 69.780 110.990 69.920 115.770 ;
        RECT 69.720 110.670 69.980 110.990 ;
        RECT 69.260 109.990 69.520 110.310 ;
        RECT 68.800 109.310 69.060 109.630 ;
        RECT 68.800 107.610 69.060 107.930 ;
        RECT 67.420 106.930 67.680 107.250 ;
        RECT 67.020 104.810 67.620 104.950 ;
        RECT 66.040 104.300 66.700 104.440 ;
        RECT 66.040 104.210 66.300 104.300 ;
        RECT 66.960 104.210 67.220 104.530 ;
        RECT 65.580 101.490 65.840 101.810 ;
        RECT 66.100 99.430 66.240 104.210 ;
        RECT 67.020 102.150 67.160 104.210 ;
        RECT 66.960 102.060 67.220 102.150 ;
        RECT 66.560 101.920 67.220 102.060 ;
        RECT 65.120 99.110 65.380 99.430 ;
        RECT 66.040 99.110 66.300 99.430 ;
        RECT 66.560 99.090 66.700 101.920 ;
        RECT 66.960 101.830 67.220 101.920 ;
        RECT 67.480 101.720 67.620 104.810 ;
        RECT 68.860 103.850 69.000 107.610 ;
        RECT 69.320 107.590 69.460 109.990 ;
        RECT 69.260 107.270 69.520 107.590 ;
        RECT 70.240 104.870 70.380 116.250 ;
        RECT 71.620 114.730 71.760 117.130 ;
        RECT 71.100 114.410 71.360 114.730 ;
        RECT 71.560 114.410 71.820 114.730 ;
        RECT 71.160 110.310 71.300 114.410 ;
        RECT 72.300 113.875 73.840 114.245 ;
        RECT 72.020 112.030 72.280 112.350 ;
        RECT 72.080 110.990 72.220 112.030 ;
        RECT 72.020 110.670 72.280 110.990 ;
        RECT 71.100 109.990 71.360 110.310 ;
        RECT 74.840 109.630 74.980 117.130 ;
        RECT 71.560 109.310 71.820 109.630 ;
        RECT 74.780 109.310 75.040 109.630 ;
        RECT 71.620 107.670 71.760 109.310 ;
        RECT 72.300 108.435 73.840 108.805 ;
        RECT 76.220 107.930 76.360 126.310 ;
        RECT 77.540 122.910 77.800 123.230 ;
        RECT 77.600 121.190 77.740 122.910 ;
        RECT 79.440 122.890 79.580 126.310 ;
        RECT 80.360 124.590 80.500 126.310 ;
        RECT 80.300 124.270 80.560 124.590 ;
        RECT 80.820 123.230 80.960 128.350 ;
        RECT 82.200 128.070 82.340 131.750 ;
        RECT 84.960 130.030 85.100 131.750 ;
        RECT 84.900 129.710 85.160 130.030 ;
        RECT 83.060 128.690 83.320 129.010 ;
        RECT 81.740 127.930 82.340 128.070 ;
        RECT 80.760 122.910 81.020 123.230 ;
        RECT 79.380 122.570 79.640 122.890 ;
        RECT 77.540 120.870 77.800 121.190 ;
        RECT 76.620 119.850 76.880 120.170 ;
        RECT 76.680 117.450 76.820 119.850 ;
        RECT 79.440 118.130 79.580 122.570 ;
        RECT 80.760 118.830 81.020 119.150 ;
        RECT 79.380 117.810 79.640 118.130 ;
        RECT 77.540 117.470 77.800 117.790 ;
        RECT 76.620 117.360 76.880 117.450 ;
        RECT 76.620 117.220 77.280 117.360 ;
        RECT 76.620 117.130 76.880 117.220 ;
        RECT 77.140 115.750 77.280 117.220 ;
        RECT 77.600 116.430 77.740 117.470 ;
        RECT 78.460 117.130 78.720 117.450 ;
        RECT 77.540 116.110 77.800 116.430 ;
        RECT 78.520 115.750 78.660 117.130 ;
        RECT 76.620 115.430 76.880 115.750 ;
        RECT 77.080 115.430 77.340 115.750 ;
        RECT 78.460 115.430 78.720 115.750 ;
        RECT 76.680 112.010 76.820 115.430 ;
        RECT 79.440 115.410 79.580 117.810 ;
        RECT 80.820 115.750 80.960 118.830 ;
        RECT 81.220 116.390 81.480 116.430 ;
        RECT 81.740 116.390 81.880 127.930 ;
        RECT 83.120 123.570 83.260 128.690 ;
        RECT 84.440 128.010 84.700 128.330 ;
        RECT 83.060 123.250 83.320 123.570 ;
        RECT 82.140 122.570 82.400 122.890 ;
        RECT 82.200 121.870 82.340 122.570 ;
        RECT 82.140 121.550 82.400 121.870 ;
        RECT 83.120 119.150 83.260 123.250 ;
        RECT 84.500 122.890 84.640 128.010 ;
        RECT 87.260 125.610 87.400 138.890 ;
        RECT 87.720 132.070 87.860 139.570 ;
        RECT 88.640 139.120 88.780 157.930 ;
        RECT 89.090 154.675 90.630 155.045 ;
        RECT 89.040 152.490 89.300 152.810 ;
        RECT 90.420 152.490 90.680 152.810 ;
        RECT 89.100 151.790 89.240 152.490 ;
        RECT 89.040 151.470 89.300 151.790 ;
        RECT 90.480 150.770 90.620 152.490 ;
        RECT 90.940 151.305 91.080 164.730 ;
        RECT 91.860 161.990 92.000 169.830 ;
        RECT 92.320 167.770 92.460 171.530 ;
        RECT 92.720 170.170 92.980 170.490 ;
        RECT 92.260 167.450 92.520 167.770 ;
        RECT 92.260 165.070 92.520 165.390 ;
        RECT 91.800 161.670 92.060 161.990 ;
        RECT 90.870 150.935 91.150 151.305 ;
        RECT 90.420 150.450 90.680 150.770 ;
        RECT 89.090 149.235 90.630 149.605 ;
        RECT 91.800 148.070 92.060 148.390 ;
        RECT 91.860 145.330 92.000 148.070 ;
        RECT 91.800 145.010 92.060 145.330 ;
        RECT 90.880 144.330 91.140 144.650 ;
        RECT 91.340 144.330 91.600 144.650 ;
        RECT 89.090 143.795 90.630 144.165 ;
        RECT 90.940 142.950 91.080 144.330 ;
        RECT 91.400 143.630 91.540 144.330 ;
        RECT 91.340 143.310 91.600 143.630 ;
        RECT 90.880 142.630 91.140 142.950 ;
        RECT 89.040 139.120 89.300 139.210 ;
        RECT 88.640 138.980 89.300 139.120 ;
        RECT 88.640 138.950 88.780 138.980 ;
        RECT 88.180 138.810 88.780 138.950 ;
        RECT 89.040 138.890 89.300 138.980 ;
        RECT 88.180 137.510 88.320 138.810 ;
        RECT 89.090 138.355 90.630 138.725 ;
        RECT 92.320 138.190 92.460 165.070 ;
        RECT 92.780 162.330 92.920 170.170 ;
        RECT 94.620 167.430 94.760 180.710 ;
        RECT 95.020 180.370 95.280 180.690 ;
        RECT 95.080 175.590 95.220 180.370 ;
        RECT 95.480 176.970 95.740 177.290 ;
        RECT 95.020 175.270 95.280 175.590 ;
        RECT 95.080 173.210 95.220 175.270 ;
        RECT 95.020 172.890 95.280 173.210 ;
        RECT 95.540 172.870 95.680 176.970 ;
        RECT 95.480 172.550 95.740 172.870 ;
        RECT 96.400 172.550 96.660 172.870 ;
        RECT 95.020 171.530 95.280 171.850 ;
        RECT 95.080 170.830 95.220 171.530 ;
        RECT 95.020 170.510 95.280 170.830 ;
        RECT 94.560 167.110 94.820 167.430 ;
        RECT 93.640 166.770 93.900 167.090 ;
        RECT 93.700 162.330 93.840 166.770 ;
        RECT 94.620 164.690 94.760 167.110 ;
        RECT 96.460 167.090 96.600 172.550 ;
        RECT 96.920 171.590 97.060 185.615 ;
        RECT 97.320 183.090 97.580 183.410 ;
        RECT 97.380 178.990 97.520 183.090 ;
        RECT 97.320 178.670 97.580 178.990 ;
        RECT 97.840 178.310 97.980 188.530 ;
        RECT 98.240 187.850 98.500 188.170 ;
        RECT 98.300 186.470 98.440 187.850 ;
        RECT 98.240 186.150 98.500 186.470 ;
        RECT 98.760 183.750 98.900 197.030 ;
        RECT 99.220 191.910 99.360 197.370 ;
        RECT 103.360 191.910 103.500 199.070 ;
        RECT 103.820 196.330 103.960 199.410 ;
        RECT 104.280 197.350 104.420 201.790 ;
        RECT 104.680 201.450 104.940 201.770 ;
        RECT 104.220 197.030 104.480 197.350 ;
        RECT 103.760 196.010 104.020 196.330 ;
        RECT 104.280 194.290 104.420 197.030 ;
        RECT 104.220 193.970 104.480 194.290 ;
        RECT 103.760 191.930 104.020 192.250 ;
        RECT 99.160 191.590 99.420 191.910 ;
        RECT 103.300 191.590 103.560 191.910 ;
        RECT 101.460 189.550 101.720 189.870 ;
        RECT 99.160 188.530 99.420 188.850 ;
        RECT 99.220 184.430 99.360 188.530 ;
        RECT 101.520 186.470 101.660 189.550 ;
        RECT 103.820 188.170 103.960 191.930 ;
        RECT 104.220 190.910 104.480 191.230 ;
        RECT 103.760 187.850 104.020 188.170 ;
        RECT 102.840 186.830 103.100 187.150 ;
        RECT 103.300 186.830 103.560 187.150 ;
        RECT 101.460 186.150 101.720 186.470 ;
        RECT 100.080 185.470 100.340 185.790 ;
        RECT 99.160 184.110 99.420 184.430 ;
        RECT 98.700 183.430 98.960 183.750 ;
        RECT 100.140 183.410 100.280 185.470 ;
        RECT 101.920 185.130 102.180 185.450 ;
        RECT 101.980 184.430 102.120 185.130 ;
        RECT 101.920 184.110 102.180 184.430 ;
        RECT 102.900 183.410 103.040 186.830 ;
        RECT 103.360 186.470 103.500 186.830 ;
        RECT 103.300 186.150 103.560 186.470 ;
        RECT 103.360 185.985 103.500 186.150 ;
        RECT 103.290 185.615 103.570 185.985 ;
        RECT 103.300 183.945 103.560 184.090 ;
        RECT 103.290 183.575 103.570 183.945 ;
        RECT 103.820 183.750 103.960 187.850 ;
        RECT 103.760 183.430 104.020 183.750 ;
        RECT 100.080 183.090 100.340 183.410 ;
        RECT 102.840 183.090 103.100 183.410 ;
        RECT 104.280 183.150 104.420 190.910 ;
        RECT 104.740 189.190 104.880 201.450 ;
        RECT 105.880 200.915 107.420 201.285 ;
        RECT 105.600 200.090 105.860 200.410 ;
        RECT 105.140 198.730 105.400 199.050 ;
        RECT 105.200 197.350 105.340 198.730 ;
        RECT 105.140 197.030 105.400 197.350 ;
        RECT 105.660 196.240 105.800 200.090 ;
        RECT 107.900 197.030 108.160 197.350 ;
        RECT 105.200 196.100 105.800 196.240 ;
        RECT 105.200 194.710 105.340 196.100 ;
        RECT 105.880 195.475 107.420 195.845 ;
        RECT 105.200 194.570 105.800 194.710 ;
        RECT 105.140 193.970 105.400 194.290 ;
        RECT 105.200 191.570 105.340 193.970 ;
        RECT 105.140 191.250 105.400 191.570 ;
        RECT 104.680 188.870 104.940 189.190 ;
        RECT 104.680 185.810 104.940 186.130 ;
        RECT 98.700 178.670 98.960 178.990 ;
        RECT 97.780 177.990 98.040 178.310 ;
        RECT 97.840 176.270 97.980 177.990 ;
        RECT 98.240 177.650 98.500 177.970 ;
        RECT 98.300 176.270 98.440 177.650 ;
        RECT 97.780 175.950 98.040 176.270 ;
        RECT 98.240 175.950 98.500 176.270 ;
        RECT 98.240 171.870 98.500 172.190 ;
        RECT 96.920 171.450 97.980 171.590 ;
        RECT 96.850 169.975 97.130 170.345 ;
        RECT 96.400 167.000 96.660 167.090 ;
        RECT 96.000 166.860 96.660 167.000 ;
        RECT 94.620 164.550 95.680 164.690 ;
        RECT 92.720 162.010 92.980 162.330 ;
        RECT 93.640 162.010 93.900 162.330 ;
        RECT 95.540 161.310 95.680 164.550 ;
        RECT 96.000 164.370 96.140 166.860 ;
        RECT 96.400 166.770 96.660 166.860 ;
        RECT 96.920 166.320 97.060 169.975 ;
        RECT 97.320 168.810 97.580 169.130 ;
        RECT 97.380 167.090 97.520 168.810 ;
        RECT 97.320 166.770 97.580 167.090 ;
        RECT 97.320 166.320 97.580 166.410 ;
        RECT 96.920 166.180 97.580 166.320 ;
        RECT 97.320 166.090 97.580 166.180 ;
        RECT 96.400 164.730 96.660 165.050 ;
        RECT 95.940 164.050 96.200 164.370 ;
        RECT 96.000 161.990 96.140 164.050 ;
        RECT 95.940 161.670 96.200 161.990 ;
        RECT 96.460 161.650 96.600 164.730 ;
        RECT 96.400 161.330 96.660 161.650 ;
        RECT 95.480 160.990 95.740 161.310 ;
        RECT 96.460 159.950 96.600 161.330 ;
        RECT 96.400 159.630 96.660 159.950 ;
        RECT 97.380 159.270 97.520 166.090 ;
        RECT 96.400 158.950 96.660 159.270 ;
        RECT 96.860 158.950 97.120 159.270 ;
        RECT 97.320 158.950 97.580 159.270 ;
        RECT 95.020 158.610 95.280 158.930 ;
        RECT 94.100 155.890 94.360 156.210 ;
        RECT 94.160 154.510 94.300 155.890 ;
        RECT 94.100 154.190 94.360 154.510 ;
        RECT 93.180 153.170 93.440 153.490 ;
        RECT 93.240 151.450 93.380 153.170 ;
        RECT 95.080 152.810 95.220 158.610 ;
        RECT 96.460 155.530 96.600 158.950 ;
        RECT 96.920 157.230 97.060 158.950 ;
        RECT 96.860 156.910 97.120 157.230 ;
        RECT 96.400 155.210 96.660 155.530 ;
        RECT 96.460 154.170 96.600 155.210 ;
        RECT 96.860 154.190 97.120 154.510 ;
        RECT 96.400 153.850 96.660 154.170 ;
        RECT 95.020 152.490 95.280 152.810 ;
        RECT 93.180 151.130 93.440 151.450 ;
        RECT 96.460 150.770 96.600 153.850 ;
        RECT 95.940 150.450 96.200 150.770 ;
        RECT 96.400 150.450 96.660 150.770 ;
        RECT 95.020 149.770 95.280 150.090 ;
        RECT 95.080 145.330 95.220 149.770 ;
        RECT 96.000 148.730 96.140 150.450 ;
        RECT 95.940 148.410 96.200 148.730 ;
        RECT 96.460 147.960 96.600 150.450 ;
        RECT 96.000 147.820 96.600 147.960 ;
        RECT 95.020 145.010 95.280 145.330 ;
        RECT 95.480 145.185 95.740 145.330 ;
        RECT 95.470 144.815 95.750 145.185 ;
        RECT 96.000 144.650 96.140 147.820 ;
        RECT 96.920 144.650 97.060 154.190 ;
        RECT 97.380 150.430 97.520 158.950 ;
        RECT 97.840 153.740 97.980 171.450 ;
        RECT 98.300 160.970 98.440 171.870 ;
        RECT 98.760 170.150 98.900 178.670 ;
        RECT 99.620 177.650 99.880 177.970 ;
        RECT 99.680 175.930 99.820 177.650 ;
        RECT 99.620 175.610 99.880 175.930 ;
        RECT 99.160 171.530 99.420 171.850 ;
        RECT 98.700 169.830 98.960 170.150 ;
        RECT 98.760 164.030 98.900 169.830 ;
        RECT 99.220 169.665 99.360 171.530 ;
        RECT 99.150 169.295 99.430 169.665 ;
        RECT 98.700 163.710 98.960 164.030 ;
        RECT 98.240 160.650 98.500 160.970 ;
        RECT 98.700 159.630 98.960 159.950 ;
        RECT 98.240 158.610 98.500 158.930 ;
        RECT 98.300 154.510 98.440 158.610 ;
        RECT 98.760 158.250 98.900 159.630 ;
        RECT 98.700 157.930 98.960 158.250 ;
        RECT 98.700 156.910 98.960 157.230 ;
        RECT 98.240 154.190 98.500 154.510 ;
        RECT 98.760 153.830 98.900 156.910 ;
        RECT 99.220 156.890 99.360 169.295 ;
        RECT 99.620 160.650 99.880 160.970 ;
        RECT 99.160 156.570 99.420 156.890 ;
        RECT 98.240 153.740 98.500 153.830 ;
        RECT 97.840 153.600 98.500 153.740 ;
        RECT 98.240 153.510 98.500 153.600 ;
        RECT 98.700 153.510 98.960 153.830 ;
        RECT 98.300 153.345 98.440 153.510 ;
        RECT 98.230 152.975 98.510 153.345 ;
        RECT 98.760 152.810 98.900 153.510 ;
        RECT 98.700 152.490 98.960 152.810 ;
        RECT 99.160 152.490 99.420 152.810 ;
        RECT 98.760 150.770 98.900 152.490 ;
        RECT 99.220 150.770 99.360 152.490 ;
        RECT 98.700 150.450 98.960 150.770 ;
        RECT 99.160 150.450 99.420 150.770 ;
        RECT 97.320 150.110 97.580 150.430 ;
        RECT 98.700 149.770 98.960 150.090 ;
        RECT 98.760 145.670 98.900 149.770 ;
        RECT 98.700 145.350 98.960 145.670 ;
        RECT 95.940 144.330 96.200 144.650 ;
        RECT 96.400 144.330 96.660 144.650 ;
        RECT 96.860 144.330 97.120 144.650 ;
        RECT 96.460 143.290 96.600 144.330 ;
        RECT 96.400 142.970 96.660 143.290 ;
        RECT 95.480 142.630 95.740 142.950 ;
        RECT 93.640 141.610 93.900 141.930 ;
        RECT 88.580 137.870 88.840 138.190 ;
        RECT 92.260 137.870 92.520 138.190 ;
        RECT 88.120 137.190 88.380 137.510 ;
        RECT 87.660 131.750 87.920 132.070 ;
        RECT 87.720 128.670 87.860 131.750 ;
        RECT 88.180 129.350 88.320 137.190 ;
        RECT 88.640 134.110 88.780 137.870 ;
        RECT 90.880 137.530 91.140 137.850 ;
        RECT 89.040 136.850 89.300 137.170 ;
        RECT 89.100 134.450 89.240 136.850 ;
        RECT 89.040 134.130 89.300 134.450 ;
        RECT 88.580 133.790 88.840 134.110 ;
        RECT 89.090 132.915 90.630 133.285 ;
        RECT 88.120 129.030 88.380 129.350 ;
        RECT 90.940 129.010 91.080 137.530 ;
        RECT 93.700 137.510 93.840 141.610 ;
        RECT 92.260 137.190 92.520 137.510 ;
        RECT 93.640 137.190 93.900 137.510 ;
        RECT 92.320 134.110 92.460 137.190 ;
        RECT 95.540 137.170 95.680 142.630 ;
        RECT 96.920 142.610 97.060 144.330 ;
        RECT 98.240 143.310 98.500 143.630 ;
        RECT 96.860 142.290 97.120 142.610 ;
        RECT 96.400 141.950 96.660 142.270 ;
        RECT 96.460 140.570 96.600 141.950 ;
        RECT 96.920 140.910 97.060 142.290 ;
        RECT 96.860 140.590 97.120 140.910 ;
        RECT 95.940 140.250 96.200 140.570 ;
        RECT 96.400 140.250 96.660 140.570 ;
        RECT 96.000 137.510 96.140 140.250 ;
        RECT 96.460 138.190 96.600 140.250 ;
        RECT 96.400 137.870 96.660 138.190 ;
        RECT 96.460 137.510 96.600 137.870 ;
        RECT 95.940 137.190 96.200 137.510 ;
        RECT 96.400 137.190 96.660 137.510 ;
        RECT 97.780 137.190 98.040 137.510 ;
        RECT 95.480 136.850 95.740 137.170 ;
        RECT 95.540 135.470 95.680 136.850 ;
        RECT 95.480 135.150 95.740 135.470 ;
        RECT 96.000 134.450 96.140 137.190 ;
        RECT 97.840 135.470 97.980 137.190 ;
        RECT 97.780 135.150 98.040 135.470 ;
        RECT 98.300 134.450 98.440 143.310 ;
        RECT 98.760 142.860 98.900 145.350 ;
        RECT 99.220 144.990 99.360 150.450 ;
        RECT 99.680 147.710 99.820 160.650 ;
        RECT 99.620 147.390 99.880 147.710 ;
        RECT 99.160 144.670 99.420 144.990 ;
        RECT 99.160 142.860 99.420 142.950 ;
        RECT 98.760 142.720 99.420 142.860 ;
        RECT 99.160 142.630 99.420 142.720 ;
        RECT 98.700 141.610 98.960 141.930 ;
        RECT 98.760 140.230 98.900 141.610 ;
        RECT 98.700 139.910 98.960 140.230 ;
        RECT 99.220 137.850 99.360 142.630 ;
        RECT 99.160 137.530 99.420 137.850 ;
        RECT 99.610 137.335 99.890 137.705 ;
        RECT 99.620 137.190 99.880 137.335 ;
        RECT 98.700 136.170 98.960 136.490 ;
        RECT 95.940 134.130 96.200 134.450 ;
        RECT 98.240 134.130 98.500 134.450 ;
        RECT 92.260 133.790 92.520 134.110 ;
        RECT 92.320 132.750 92.460 133.790 ;
        RECT 92.260 132.430 92.520 132.750 ;
        RECT 97.780 131.980 98.040 132.070 ;
        RECT 98.760 131.980 98.900 136.170 ;
        RECT 97.780 131.840 98.900 131.980 ;
        RECT 97.780 131.750 98.040 131.840 ;
        RECT 95.940 131.410 96.200 131.730 ;
        RECT 94.100 129.370 94.360 129.690 ;
        RECT 90.880 128.690 91.140 129.010 ;
        RECT 91.340 128.690 91.600 129.010 ;
        RECT 87.660 128.350 87.920 128.670 ;
        RECT 89.090 127.475 90.630 127.845 ;
        RECT 85.820 125.290 86.080 125.610 ;
        RECT 86.280 125.290 86.540 125.610 ;
        RECT 87.200 125.290 87.460 125.610 ;
        RECT 84.900 122.910 85.160 123.230 ;
        RECT 84.440 122.570 84.700 122.890 ;
        RECT 83.980 119.850 84.240 120.170 ;
        RECT 84.040 119.150 84.180 119.850 ;
        RECT 83.060 119.060 83.320 119.150 ;
        RECT 82.660 118.920 83.320 119.060 ;
        RECT 82.140 117.470 82.400 117.790 ;
        RECT 81.220 116.250 81.880 116.390 ;
        RECT 81.220 116.110 81.480 116.250 ;
        RECT 80.760 115.660 81.020 115.750 ;
        RECT 79.900 115.520 81.020 115.660 ;
        RECT 79.380 115.090 79.640 115.410 ;
        RECT 79.440 113.030 79.580 115.090 ;
        RECT 79.380 112.710 79.640 113.030 ;
        RECT 76.620 111.690 76.880 112.010 ;
        RECT 79.380 110.670 79.640 110.990 ;
        RECT 78.000 109.990 78.260 110.310 ;
        RECT 76.620 107.950 76.880 108.270 ;
        RECT 71.620 107.530 72.220 107.670 ;
        RECT 76.160 107.610 76.420 107.930 ;
        RECT 71.560 106.930 71.820 107.250 ;
        RECT 70.640 106.250 70.900 106.570 ;
        RECT 70.700 105.210 70.840 106.250 ;
        RECT 71.620 105.550 71.760 106.930 ;
        RECT 71.560 105.230 71.820 105.550 ;
        RECT 72.080 105.210 72.220 107.530 ;
        RECT 74.320 106.930 74.580 107.250 ;
        RECT 76.160 106.930 76.420 107.250 ;
        RECT 70.640 104.890 70.900 105.210 ;
        RECT 72.020 104.890 72.280 105.210 ;
        RECT 70.180 104.550 70.440 104.870 ;
        RECT 74.380 103.850 74.520 106.930 ;
        RECT 75.240 106.250 75.500 106.570 ;
        RECT 75.700 106.250 75.960 106.570 ;
        RECT 68.800 103.530 69.060 103.850 ;
        RECT 71.560 103.530 71.820 103.850 ;
        RECT 74.320 103.530 74.580 103.850 ;
        RECT 67.880 101.720 68.140 101.810 ;
        RECT 67.480 101.580 68.140 101.720 ;
        RECT 67.880 101.490 68.140 101.580 ;
        RECT 66.500 98.770 66.760 99.090 ;
        RECT 66.560 96.710 66.700 98.770 ;
        RECT 67.940 98.750 68.080 101.490 ;
        RECT 67.880 98.430 68.140 98.750 ;
        RECT 66.500 96.390 66.760 96.710 ;
        RECT 66.560 93.990 66.700 96.390 ;
        RECT 67.880 96.050 68.140 96.370 ;
        RECT 66.500 93.670 66.760 93.990 ;
        RECT 65.580 93.330 65.840 93.650 ;
        RECT 65.640 91.950 65.780 93.330 ;
        RECT 65.580 91.630 65.840 91.950 ;
        RECT 66.560 88.550 66.700 93.670 ;
        RECT 67.940 91.950 68.080 96.050 ;
        RECT 68.860 93.990 69.000 103.530 ;
        RECT 71.620 101.810 71.760 103.530 ;
        RECT 72.300 102.995 73.840 103.365 ;
        RECT 75.300 102.150 75.440 106.250 ;
        RECT 75.760 103.850 75.900 106.250 ;
        RECT 75.700 103.530 75.960 103.850 ;
        RECT 75.240 101.830 75.500 102.150 ;
        RECT 71.560 101.490 71.820 101.810 ;
        RECT 74.320 99.450 74.580 99.770 ;
        RECT 71.560 99.110 71.820 99.430 ;
        RECT 71.100 98.090 71.360 98.410 ;
        RECT 71.160 96.030 71.300 98.090 ;
        RECT 71.620 96.030 71.760 99.110 ;
        RECT 72.300 97.555 73.840 97.925 ;
        RECT 72.480 96.730 72.740 97.050 ;
        RECT 72.540 96.030 72.680 96.730 ;
        RECT 72.940 96.050 73.200 96.370 ;
        RECT 71.100 95.710 71.360 96.030 ;
        RECT 71.560 95.710 71.820 96.030 ;
        RECT 72.480 95.710 72.740 96.030 ;
        RECT 68.800 93.670 69.060 93.990 ;
        RECT 67.880 91.630 68.140 91.950 ;
        RECT 66.960 90.950 67.220 91.270 ;
        RECT 66.500 88.230 66.760 88.550 ;
        RECT 65.120 87.210 65.380 87.530 ;
        RECT 65.180 85.490 65.320 87.210 ;
        RECT 66.040 85.850 66.300 86.170 ;
        RECT 65.120 85.170 65.380 85.490 ;
        RECT 66.100 80.050 66.240 85.850 ;
        RECT 66.560 83.450 66.700 88.230 ;
        RECT 67.020 85.150 67.160 90.950 ;
        RECT 68.860 90.930 69.000 93.670 ;
        RECT 71.160 91.950 71.300 95.710 ;
        RECT 72.540 94.670 72.680 95.710 ;
        RECT 73.000 94.670 73.140 96.050 ;
        RECT 72.480 94.350 72.740 94.670 ;
        RECT 72.940 94.350 73.200 94.670 ;
        RECT 74.380 93.990 74.520 99.450 ;
        RECT 75.700 97.070 75.960 97.390 ;
        RECT 75.760 96.030 75.900 97.070 ;
        RECT 75.700 95.710 75.960 96.030 ;
        RECT 74.320 93.670 74.580 93.990 ;
        RECT 72.300 92.115 73.840 92.485 ;
        RECT 71.100 91.630 71.360 91.950 ;
        RECT 68.340 90.610 68.600 90.930 ;
        RECT 68.800 90.610 69.060 90.930 ;
        RECT 68.400 90.250 68.540 90.610 ;
        RECT 68.340 89.930 68.600 90.250 ;
        RECT 71.560 89.930 71.820 90.250 ;
        RECT 69.720 86.190 69.980 86.510 ;
        RECT 69.780 85.490 69.920 86.190 ;
        RECT 71.620 86.170 71.760 89.930 ;
        RECT 72.300 86.675 73.840 87.045 ;
        RECT 71.560 85.850 71.820 86.170 ;
        RECT 69.260 85.170 69.520 85.490 ;
        RECT 69.720 85.170 69.980 85.490 ;
        RECT 70.180 85.170 70.440 85.490 ;
        RECT 72.480 85.170 72.740 85.490 ;
        RECT 66.960 84.830 67.220 85.150 ;
        RECT 69.320 84.810 69.460 85.170 ;
        RECT 69.260 84.490 69.520 84.810 ;
        RECT 70.240 83.790 70.380 85.170 ;
        RECT 72.540 83.790 72.680 85.170 ;
        RECT 70.180 83.470 70.440 83.790 ;
        RECT 72.480 83.470 72.740 83.790 ;
        RECT 66.500 83.130 66.760 83.450 ;
        RECT 70.640 82.790 70.900 83.110 ;
        RECT 66.040 79.730 66.300 80.050 ;
        RECT 66.960 76.330 67.220 76.650 ;
        RECT 68.340 76.330 68.600 76.650 ;
        RECT 67.020 74.950 67.160 76.330 ;
        RECT 66.960 74.630 67.220 74.950 ;
        RECT 65.120 74.520 65.380 74.610 ;
        RECT 64.720 74.380 65.380 74.520 ;
        RECT 65.120 74.290 65.380 74.380 ;
        RECT 59.200 72.570 59.340 74.290 ;
        RECT 60.120 72.910 60.260 74.290 ;
        RECT 60.060 72.590 60.320 72.910 ;
        RECT 59.140 72.250 59.400 72.570 ;
        RECT 58.680 68.850 58.940 69.170 ;
        RECT 59.200 69.080 59.340 72.250 ;
        RECT 60.060 70.890 60.320 71.210 ;
        RECT 60.120 69.850 60.260 70.890 ;
        RECT 60.060 69.530 60.320 69.850 ;
        RECT 59.600 69.080 59.860 69.170 ;
        RECT 59.200 68.940 59.860 69.080 ;
        RECT 59.600 68.850 59.860 68.940 ;
        RECT 59.600 68.170 59.860 68.490 ;
        RECT 59.660 66.790 59.800 68.170 ;
        RECT 60.120 66.790 60.260 69.530 ;
        RECT 60.580 67.470 60.720 74.290 ;
        RECT 62.820 73.950 63.080 74.270 ;
        RECT 62.880 72.230 63.020 73.950 ;
        RECT 63.800 72.570 63.940 74.290 ;
        RECT 68.400 72.910 68.540 76.330 ;
        RECT 70.700 72.910 70.840 82.790 ;
        RECT 72.300 81.235 73.840 81.605 ;
        RECT 73.860 79.730 74.120 80.050 ;
        RECT 73.920 78.350 74.060 79.730 ;
        RECT 73.860 78.030 74.120 78.350 ;
        RECT 72.300 75.795 73.840 76.165 ;
        RECT 74.380 73.930 74.520 93.670 ;
        RECT 76.220 78.260 76.360 106.930 ;
        RECT 76.680 105.210 76.820 107.950 ;
        RECT 78.060 105.550 78.200 109.990 ;
        RECT 79.440 105.550 79.580 110.670 ;
        RECT 78.000 105.230 78.260 105.550 ;
        RECT 79.380 105.230 79.640 105.550 ;
        RECT 76.620 104.890 76.880 105.210 ;
        RECT 79.900 104.870 80.040 115.520 ;
        RECT 80.760 115.430 81.020 115.520 ;
        RECT 81.280 114.730 81.420 116.110 ;
        RECT 82.200 115.830 82.340 117.470 ;
        RECT 81.740 115.690 82.340 115.830 ;
        RECT 81.220 114.410 81.480 114.730 ;
        RECT 81.220 107.670 81.480 107.930 ;
        RECT 80.360 107.610 81.480 107.670 ;
        RECT 80.360 107.530 81.420 107.610 ;
        RECT 80.360 106.910 80.500 107.530 ;
        RECT 80.760 107.105 81.020 107.250 ;
        RECT 80.300 106.590 80.560 106.910 ;
        RECT 80.750 106.735 81.030 107.105 ;
        RECT 81.220 106.250 81.480 106.570 ;
        RECT 79.380 104.550 79.640 104.870 ;
        RECT 79.840 104.550 80.100 104.870 ;
        RECT 78.460 101.490 78.720 101.810 ;
        RECT 76.620 100.810 76.880 101.130 ;
        RECT 76.680 99.770 76.820 100.810 ;
        RECT 76.620 99.450 76.880 99.770 ;
        RECT 78.520 97.390 78.660 101.490 ;
        RECT 78.460 97.070 78.720 97.390 ;
        RECT 79.440 96.030 79.580 104.550 ;
        RECT 79.900 101.810 80.040 104.550 ;
        RECT 81.280 103.850 81.420 106.250 ;
        RECT 81.740 105.210 81.880 115.690 ;
        RECT 82.660 112.690 82.800 118.920 ;
        RECT 83.060 118.830 83.320 118.920 ;
        RECT 83.980 118.830 84.240 119.150 ;
        RECT 84.500 117.790 84.640 122.570 ;
        RECT 84.960 117.790 85.100 122.910 ;
        RECT 85.360 120.530 85.620 120.850 ;
        RECT 85.420 118.810 85.560 120.530 ;
        RECT 85.360 118.490 85.620 118.810 ;
        RECT 85.420 118.130 85.560 118.490 ;
        RECT 85.360 117.810 85.620 118.130 ;
        RECT 84.440 117.470 84.700 117.790 ;
        RECT 84.900 117.470 85.160 117.790 ;
        RECT 83.520 115.430 83.780 115.750 ;
        RECT 83.580 113.710 83.720 115.430 ;
        RECT 83.520 113.390 83.780 113.710 ;
        RECT 82.600 112.370 82.860 112.690 ;
        RECT 84.500 112.350 84.640 117.470 ;
        RECT 84.960 112.350 85.100 117.470 ;
        RECT 85.360 117.130 85.620 117.450 ;
        RECT 84.440 112.030 84.700 112.350 ;
        RECT 84.900 112.030 85.160 112.350 ;
        RECT 82.600 111.690 82.860 112.010 ;
        RECT 82.660 110.990 82.800 111.690 ;
        RECT 82.600 110.670 82.860 110.990 ;
        RECT 84.440 108.970 84.700 109.290 ;
        RECT 84.500 107.590 84.640 108.970 ;
        RECT 84.960 108.270 85.100 112.030 ;
        RECT 84.900 107.950 85.160 108.270 ;
        RECT 84.960 107.590 85.100 107.950 ;
        RECT 83.980 107.270 84.240 107.590 ;
        RECT 84.440 107.270 84.700 107.590 ;
        RECT 84.900 107.270 85.160 107.590 ;
        RECT 82.130 106.735 82.410 107.105 ;
        RECT 81.680 104.890 81.940 105.210 ;
        RECT 81.670 104.015 81.950 104.385 ;
        RECT 81.220 103.530 81.480 103.850 ;
        RECT 80.300 102.345 80.560 102.490 ;
        RECT 80.290 101.975 80.570 102.345 ;
        RECT 80.760 102.170 81.020 102.490 ;
        RECT 80.820 101.810 80.960 102.170 ;
        RECT 81.740 102.150 81.880 104.015 ;
        RECT 82.200 102.830 82.340 106.735 ;
        RECT 84.040 105.210 84.180 107.270 ;
        RECT 83.980 104.890 84.240 105.210 ;
        RECT 84.900 104.550 85.160 104.870 ;
        RECT 82.600 104.210 82.860 104.530 ;
        RECT 82.140 102.510 82.400 102.830 ;
        RECT 81.680 101.830 81.940 102.150 ;
        RECT 82.200 101.810 82.340 102.510 ;
        RECT 79.840 101.490 80.100 101.810 ;
        RECT 80.760 101.490 81.020 101.810 ;
        RECT 82.140 101.490 82.400 101.810 ;
        RECT 79.840 100.810 80.100 101.130 ;
        RECT 79.380 95.710 79.640 96.030 ;
        RECT 76.620 92.650 76.880 92.970 ;
        RECT 76.680 90.930 76.820 92.650 ;
        RECT 76.620 90.610 76.880 90.930 ;
        RECT 76.620 89.930 76.880 90.250 ;
        RECT 78.460 89.930 78.720 90.250 ;
        RECT 76.680 88.890 76.820 89.930 ;
        RECT 78.520 89.230 78.660 89.930 ;
        RECT 78.460 88.910 78.720 89.230 ;
        RECT 76.620 88.570 76.880 88.890 ;
        RECT 77.540 88.230 77.800 88.550 ;
        RECT 77.600 86.510 77.740 88.230 ;
        RECT 77.540 86.190 77.800 86.510 ;
        RECT 77.600 85.490 77.740 86.190 ;
        RECT 77.540 85.170 77.800 85.490 ;
        RECT 78.920 85.170 79.180 85.490 ;
        RECT 78.980 83.790 79.120 85.170 ;
        RECT 78.920 83.470 79.180 83.790 ;
        RECT 78.980 81.070 79.120 83.470 ;
        RECT 78.920 80.750 79.180 81.070 ;
        RECT 79.380 80.410 79.640 80.730 ;
        RECT 76.620 79.390 76.880 79.710 ;
        RECT 75.760 78.120 76.360 78.260 ;
        RECT 75.760 77.670 75.900 78.120 ;
        RECT 75.700 77.350 75.960 77.670 ;
        RECT 76.160 77.580 76.420 77.670 ;
        RECT 76.680 77.580 76.820 79.390 ;
        RECT 79.440 78.010 79.580 80.410 ;
        RECT 79.900 80.050 80.040 100.810 ;
        RECT 80.820 100.110 80.960 101.490 ;
        RECT 80.760 99.790 81.020 100.110 ;
        RECT 82.660 98.830 82.800 104.210 ;
        RECT 83.050 104.015 83.330 104.385 ;
        RECT 83.120 99.625 83.260 104.015 ;
        RECT 84.440 103.530 84.700 103.850 ;
        RECT 84.500 101.810 84.640 103.530 ;
        RECT 84.960 101.810 85.100 104.550 ;
        RECT 85.420 102.150 85.560 117.130 ;
        RECT 85.880 104.870 86.020 125.290 ;
        RECT 86.340 124.590 86.480 125.290 ;
        RECT 86.280 124.270 86.540 124.590 ;
        RECT 86.740 123.250 87.000 123.570 ;
        RECT 86.800 121.530 86.940 123.250 ;
        RECT 87.260 121.870 87.400 125.290 ;
        RECT 88.570 123.735 88.850 124.105 ;
        RECT 90.940 123.910 91.080 128.690 ;
        RECT 91.400 126.290 91.540 128.690 ;
        RECT 94.160 128.670 94.300 129.370 ;
        RECT 96.000 128.670 96.140 131.410 ;
        RECT 94.100 128.350 94.360 128.670 ;
        RECT 95.940 128.350 96.200 128.670 ;
        RECT 92.720 126.310 92.980 126.630 ;
        RECT 91.340 125.970 91.600 126.290 ;
        RECT 91.400 123.910 91.540 125.970 ;
        RECT 92.780 124.590 92.920 126.310 ;
        RECT 92.260 124.270 92.520 124.590 ;
        RECT 92.720 124.270 92.980 124.590 ;
        RECT 88.640 123.570 88.780 123.735 ;
        RECT 90.880 123.590 91.140 123.910 ;
        RECT 91.340 123.590 91.600 123.910 ;
        RECT 88.580 123.250 88.840 123.570 ;
        RECT 87.200 121.550 87.460 121.870 ;
        RECT 86.740 121.210 87.000 121.530 ;
        RECT 87.200 117.810 87.460 118.130 ;
        RECT 87.260 116.430 87.400 117.810 ;
        RECT 87.200 116.110 87.460 116.430 ;
        RECT 87.260 113.710 87.400 116.110 ;
        RECT 88.120 114.750 88.380 115.070 ;
        RECT 86.280 113.390 86.540 113.710 ;
        RECT 87.200 113.390 87.460 113.710 ;
        RECT 86.340 107.250 86.480 113.390 ;
        RECT 88.180 112.350 88.320 114.750 ;
        RECT 88.120 112.030 88.380 112.350 ;
        RECT 88.120 110.330 88.380 110.650 ;
        RECT 87.200 109.990 87.460 110.310 ;
        RECT 87.260 108.270 87.400 109.990 ;
        RECT 87.200 107.950 87.460 108.270 ;
        RECT 86.280 106.930 86.540 107.250 ;
        RECT 86.340 105.210 86.480 106.930 ;
        RECT 86.280 104.890 86.540 105.210 ;
        RECT 85.820 104.550 86.080 104.870 ;
        RECT 86.280 103.530 86.540 103.850 ;
        RECT 85.820 102.510 86.080 102.830 ;
        RECT 85.360 101.830 85.620 102.150 ;
        RECT 85.880 101.810 86.020 102.510 ;
        RECT 86.340 101.810 86.480 103.530 ;
        RECT 88.180 101.810 88.320 110.330 ;
        RECT 84.440 101.490 84.700 101.810 ;
        RECT 84.900 101.490 85.160 101.810 ;
        RECT 85.820 101.490 86.080 101.810 ;
        RECT 86.280 101.490 86.540 101.810 ;
        RECT 88.120 101.490 88.380 101.810 ;
        RECT 84.960 101.130 85.100 101.490 ;
        RECT 83.520 100.810 83.780 101.130 ;
        RECT 83.980 100.810 84.240 101.130 ;
        RECT 84.900 100.810 85.160 101.130 ;
        RECT 83.050 99.255 83.330 99.625 ;
        RECT 81.280 98.690 82.800 98.830 ;
        RECT 81.280 96.370 81.420 98.690 ;
        RECT 81.680 98.090 81.940 98.410 ;
        RECT 82.140 98.090 82.400 98.410 ;
        RECT 81.740 96.370 81.880 98.090 ;
        RECT 81.220 96.050 81.480 96.370 ;
        RECT 81.680 96.050 81.940 96.370 ;
        RECT 81.680 93.330 81.940 93.650 ;
        RECT 81.220 92.990 81.480 93.310 ;
        RECT 80.300 92.650 80.560 92.970 ;
        RECT 80.360 90.930 80.500 92.650 ;
        RECT 81.280 91.610 81.420 92.990 ;
        RECT 81.220 91.290 81.480 91.610 ;
        RECT 80.300 90.610 80.560 90.930 ;
        RECT 80.760 87.890 81.020 88.210 ;
        RECT 80.820 84.810 80.960 87.890 ;
        RECT 81.280 85.490 81.420 91.290 ;
        RECT 81.740 90.590 81.880 93.330 ;
        RECT 81.680 90.270 81.940 90.590 ;
        RECT 81.740 88.210 81.880 90.270 ;
        RECT 81.680 87.890 81.940 88.210 ;
        RECT 81.680 87.210 81.940 87.530 ;
        RECT 81.740 86.170 81.880 87.210 ;
        RECT 81.680 85.850 81.940 86.170 ;
        RECT 81.220 85.170 81.480 85.490 ;
        RECT 81.680 85.170 81.940 85.490 ;
        RECT 80.760 84.490 81.020 84.810 ;
        RECT 81.740 83.790 81.880 85.170 ;
        RECT 81.680 83.470 81.940 83.790 ;
        RECT 82.200 81.150 82.340 98.090 ;
        RECT 82.600 90.610 82.860 90.930 ;
        RECT 82.660 89.230 82.800 90.610 ;
        RECT 82.600 88.910 82.860 89.230 ;
        RECT 82.600 88.230 82.860 88.550 ;
        RECT 82.660 86.510 82.800 88.230 ;
        RECT 82.600 86.190 82.860 86.510 ;
        RECT 82.600 81.770 82.860 82.090 ;
        RECT 81.740 81.010 82.340 81.150 ;
        RECT 81.740 80.730 81.880 81.010 ;
        RECT 81.680 80.410 81.940 80.730 ;
        RECT 82.660 80.050 82.800 81.770 ;
        RECT 83.580 80.050 83.720 100.810 ;
        RECT 84.040 99.430 84.180 100.810 ;
        RECT 83.980 99.110 84.240 99.430 ;
        RECT 84.960 96.370 85.100 100.810 ;
        RECT 85.360 99.110 85.620 99.430 ;
        RECT 85.420 97.390 85.560 99.110 ;
        RECT 85.880 99.090 86.020 101.490 ;
        RECT 87.660 100.810 87.920 101.130 ;
        RECT 87.720 100.110 87.860 100.810 ;
        RECT 87.660 99.790 87.920 100.110 ;
        RECT 85.820 98.770 86.080 99.090 ;
        RECT 85.360 97.070 85.620 97.390 ;
        RECT 88.180 96.710 88.320 101.490 ;
        RECT 88.640 97.050 88.780 123.250 ;
        RECT 89.090 122.035 90.630 122.405 ;
        RECT 90.940 121.530 91.080 123.590 ;
        RECT 91.800 121.550 92.060 121.870 ;
        RECT 90.880 121.210 91.140 121.530 ;
        RECT 91.340 119.850 91.600 120.170 ;
        RECT 90.880 117.470 91.140 117.790 ;
        RECT 89.090 116.595 90.630 116.965 ;
        RECT 90.940 116.430 91.080 117.470 ;
        RECT 91.400 116.430 91.540 119.850 ;
        RECT 90.880 116.110 91.140 116.430 ;
        RECT 91.340 116.110 91.600 116.430 ;
        RECT 91.340 115.430 91.600 115.750 ;
        RECT 89.090 111.155 90.630 111.525 ;
        RECT 91.400 110.650 91.540 115.430 ;
        RECT 91.860 112.010 92.000 121.550 ;
        RECT 92.320 115.750 92.460 124.270 ;
        RECT 93.180 123.590 93.440 123.910 ;
        RECT 92.720 122.910 92.980 123.230 ;
        RECT 92.780 121.530 92.920 122.910 ;
        RECT 92.720 121.210 92.980 121.530 ;
        RECT 92.260 115.430 92.520 115.750 ;
        RECT 92.780 112.690 92.920 121.210 ;
        RECT 93.240 118.130 93.380 123.590 ;
        RECT 93.180 117.810 93.440 118.130 ;
        RECT 94.160 116.090 94.300 128.350 ;
        RECT 97.840 126.970 97.980 131.750 ;
        RECT 97.780 126.650 98.040 126.970 ;
        RECT 95.020 125.290 95.280 125.610 ;
        RECT 95.080 124.590 95.220 125.290 ;
        RECT 95.020 124.270 95.280 124.590 ;
        RECT 95.080 122.890 95.220 124.270 ;
        RECT 95.480 123.930 95.740 124.250 ;
        RECT 95.540 123.570 95.680 123.930 ;
        RECT 95.480 123.250 95.740 123.570 ;
        RECT 95.020 122.570 95.280 122.890 ;
        RECT 95.940 122.800 96.200 122.890 ;
        RECT 95.540 122.660 96.200 122.800 ;
        RECT 95.540 121.870 95.680 122.660 ;
        RECT 95.940 122.570 96.200 122.660 ;
        RECT 95.480 121.550 95.740 121.870 ;
        RECT 100.140 121.190 100.280 183.090 ;
        RECT 101.000 175.270 101.260 175.590 ;
        RECT 101.060 164.905 101.200 175.270 ;
        RECT 101.920 174.930 102.180 175.250 ;
        RECT 101.460 171.870 101.720 172.190 ;
        RECT 101.520 170.150 101.660 171.870 ;
        RECT 101.460 169.830 101.720 170.150 ;
        RECT 101.980 169.470 102.120 174.930 ;
        RECT 102.380 174.250 102.640 174.570 ;
        RECT 101.920 169.150 102.180 169.470 ;
        RECT 101.980 167.770 102.120 169.150 ;
        RECT 101.920 167.450 102.180 167.770 ;
        RECT 100.990 164.535 101.270 164.905 ;
        RECT 102.440 164.690 102.580 174.250 ;
        RECT 102.900 170.490 103.040 183.090 ;
        RECT 103.820 183.010 104.420 183.150 ;
        RECT 103.300 170.510 103.560 170.830 ;
        RECT 102.840 170.170 103.100 170.490 ;
        RECT 102.900 168.110 103.040 170.170 ;
        RECT 102.840 167.790 103.100 168.110 ;
        RECT 103.360 165.390 103.500 170.510 ;
        RECT 103.300 165.070 103.560 165.390 ;
        RECT 101.980 164.550 102.580 164.690 ;
        RECT 100.540 163.710 100.800 164.030 ;
        RECT 100.600 161.650 100.740 163.710 ;
        RECT 100.540 161.330 100.800 161.650 ;
        RECT 101.000 161.505 101.260 161.650 ;
        RECT 100.600 151.190 100.740 161.330 ;
        RECT 100.990 161.135 101.270 161.505 ;
        RECT 101.980 160.970 102.120 164.550 ;
        RECT 102.380 163.370 102.640 163.690 ;
        RECT 101.920 160.650 102.180 160.970 ;
        RECT 101.000 158.950 101.260 159.270 ;
        RECT 101.060 151.790 101.200 158.950 ;
        RECT 101.460 157.930 101.720 158.250 ;
        RECT 101.520 156.210 101.660 157.930 ;
        RECT 101.460 155.890 101.720 156.210 ;
        RECT 102.440 153.490 102.580 163.370 ;
        RECT 102.380 153.170 102.640 153.490 ;
        RECT 101.000 151.470 101.260 151.790 ;
        RECT 100.600 151.050 101.200 151.190 ;
        RECT 100.540 150.450 100.800 150.770 ;
        RECT 100.600 147.710 100.740 150.450 ;
        RECT 100.540 147.390 100.800 147.710 ;
        RECT 100.600 145.185 100.740 147.390 ;
        RECT 100.530 144.815 100.810 145.185 ;
        RECT 100.540 144.670 100.800 144.815 ;
        RECT 101.060 129.010 101.200 151.050 ;
        RECT 101.460 145.690 101.720 146.010 ;
        RECT 101.520 145.330 101.660 145.690 ;
        RECT 101.460 145.010 101.720 145.330 ;
        RECT 102.440 137.510 102.580 153.170 ;
        RECT 103.360 151.870 103.500 165.070 ;
        RECT 103.820 164.710 103.960 183.010 ;
        RECT 104.740 177.290 104.880 185.810 ;
        RECT 105.200 180.690 105.340 191.250 ;
        RECT 105.660 191.230 105.800 194.570 ;
        RECT 107.960 192.250 108.100 197.030 ;
        RECT 107.900 191.930 108.160 192.250 ;
        RECT 105.600 190.910 105.860 191.230 ;
        RECT 105.880 190.035 107.420 190.405 ;
        RECT 105.600 188.530 105.860 188.850 ;
        RECT 105.660 185.790 105.800 188.530 ;
        RECT 107.440 188.190 107.700 188.510 ;
        RECT 105.600 185.470 105.860 185.790 ;
        RECT 107.500 185.390 107.640 188.190 ;
        RECT 107.500 185.250 108.100 185.390 ;
        RECT 105.880 184.595 107.420 184.965 ;
        RECT 107.960 183.945 108.100 185.250 ;
        RECT 107.890 183.575 108.170 183.945 ;
        RECT 108.420 183.150 108.560 206.980 ;
        RECT 108.820 206.890 109.080 206.980 ;
        RECT 110.260 205.850 110.400 207.910 ;
        RECT 113.940 207.630 114.080 207.910 ;
        RECT 113.480 207.490 114.080 207.630 ;
        RECT 113.480 207.210 113.620 207.490 ;
        RECT 113.420 206.890 113.680 207.210 ;
        RECT 110.200 205.530 110.460 205.850 ;
        RECT 112.500 204.850 112.760 205.170 ;
        RECT 112.560 203.470 112.700 204.850 ;
        RECT 112.500 203.150 112.760 203.470 ;
        RECT 112.500 199.750 112.760 200.070 ;
        RECT 112.040 197.030 112.300 197.350 ;
        RECT 109.280 196.010 109.540 196.330 ;
        RECT 108.820 191.590 109.080 191.910 ;
        RECT 108.880 191.425 109.020 191.590 ;
        RECT 108.810 191.055 109.090 191.425 ;
        RECT 108.820 188.530 109.080 188.850 ;
        RECT 108.880 183.320 109.020 188.530 ;
        RECT 109.340 186.470 109.480 196.010 ;
        RECT 112.100 195.310 112.240 197.030 ;
        RECT 112.040 194.990 112.300 195.310 ;
        RECT 112.040 193.970 112.300 194.290 ;
        RECT 111.580 193.630 111.840 193.950 ;
        RECT 109.740 191.590 110.000 191.910 ;
        RECT 109.800 189.870 109.940 191.590 ;
        RECT 109.740 189.550 110.000 189.870 ;
        RECT 111.640 189.530 111.780 193.630 ;
        RECT 111.580 189.210 111.840 189.530 ;
        RECT 110.660 188.530 110.920 188.850 ;
        RECT 109.280 186.150 109.540 186.470 ;
        RECT 109.730 186.295 110.010 186.665 ;
        RECT 110.720 186.380 110.860 188.530 ;
        RECT 111.120 188.190 111.380 188.510 ;
        RECT 111.180 188.025 111.320 188.190 ;
        RECT 111.110 187.655 111.390 188.025 ;
        RECT 111.120 186.380 111.380 186.470 ;
        RECT 111.640 186.380 111.780 189.210 ;
        RECT 112.100 188.850 112.240 193.970 ;
        RECT 112.040 188.530 112.300 188.850 ;
        RECT 112.100 186.470 112.240 188.530 ;
        RECT 112.560 188.025 112.700 199.750 ;
        RECT 113.480 194.710 113.620 206.890 ;
        RECT 114.340 202.470 114.600 202.790 ;
        RECT 114.400 200.750 114.540 202.470 ;
        RECT 114.340 200.430 114.600 200.750 ;
        RECT 114.860 200.070 115.000 208.000 ;
        RECT 115.260 207.910 115.520 208.000 ;
        RECT 114.800 199.980 115.060 200.070 ;
        RECT 114.400 199.840 115.060 199.980 ;
        RECT 113.880 197.030 114.140 197.350 ;
        RECT 113.940 195.310 114.080 197.030 ;
        RECT 113.880 194.990 114.140 195.310 ;
        RECT 113.480 194.570 114.080 194.710 ;
        RECT 113.420 191.590 113.680 191.910 ;
        RECT 112.490 187.655 112.770 188.025 ;
        RECT 109.800 186.130 109.940 186.295 ;
        RECT 110.720 186.240 111.780 186.380 ;
        RECT 109.740 185.810 110.000 186.130 ;
        RECT 110.720 183.410 110.860 186.240 ;
        RECT 111.120 186.150 111.380 186.240 ;
        RECT 112.040 186.150 112.300 186.470 ;
        RECT 111.120 185.470 111.380 185.790 ;
        RECT 111.180 183.410 111.320 185.470 ;
        RECT 112.100 183.750 112.240 186.150 ;
        RECT 112.040 183.430 112.300 183.750 ;
        RECT 109.280 183.320 109.540 183.410 ;
        RECT 108.880 183.180 109.540 183.320 ;
        RECT 107.960 183.010 108.560 183.150 ;
        RECT 109.280 183.090 109.540 183.180 ;
        RECT 110.660 183.090 110.920 183.410 ;
        RECT 111.120 183.090 111.380 183.410 ;
        RECT 105.140 180.370 105.400 180.690 ;
        RECT 105.200 177.970 105.340 180.370 ;
        RECT 105.880 179.155 107.420 179.525 ;
        RECT 105.140 177.650 105.400 177.970 ;
        RECT 104.680 176.970 104.940 177.290 ;
        RECT 106.980 176.970 107.240 177.290 ;
        RECT 107.040 176.270 107.180 176.970 ;
        RECT 106.980 175.950 107.240 176.270 ;
        RECT 107.960 174.990 108.100 183.010 ;
        RECT 108.360 182.410 108.620 182.730 ;
        RECT 108.420 181.370 108.560 182.410 ;
        RECT 108.360 181.050 108.620 181.370 ;
        RECT 108.820 180.370 109.080 180.690 ;
        RECT 108.360 179.690 108.620 180.010 ;
        RECT 108.420 178.650 108.560 179.690 ;
        RECT 108.880 178.650 109.020 180.370 ;
        RECT 108.360 178.330 108.620 178.650 ;
        RECT 108.820 178.330 109.080 178.650 ;
        RECT 107.960 174.850 108.560 174.990 ;
        RECT 107.900 174.250 108.160 174.570 ;
        RECT 105.880 173.715 107.420 174.085 ;
        RECT 104.220 172.210 104.480 172.530 ;
        RECT 104.280 170.830 104.420 172.210 ;
        RECT 107.960 170.830 108.100 174.250 ;
        RECT 104.220 170.510 104.480 170.830 ;
        RECT 107.900 170.510 108.160 170.830 ;
        RECT 108.420 170.490 108.560 174.850 ;
        RECT 108.880 172.870 109.020 178.330 ;
        RECT 109.340 177.880 109.480 183.090 ;
        RECT 109.740 182.750 110.000 183.070 ;
        RECT 109.800 182.585 109.940 182.750 ;
        RECT 109.730 182.215 110.010 182.585 ;
        RECT 110.720 178.650 110.860 183.090 ;
        RECT 110.660 178.330 110.920 178.650 ;
        RECT 109.740 177.880 110.000 177.970 ;
        RECT 109.340 177.740 110.000 177.880 ;
        RECT 109.740 177.650 110.000 177.740 ;
        RECT 108.820 172.550 109.080 172.870 ;
        RECT 108.360 170.170 108.620 170.490 ;
        RECT 105.880 168.275 107.420 168.645 ;
        RECT 109.800 167.430 109.940 177.650 ;
        RECT 112.040 177.310 112.300 177.630 ;
        RECT 110.660 174.930 110.920 175.250 ;
        RECT 110.720 173.550 110.860 174.930 ;
        RECT 110.660 173.230 110.920 173.550 ;
        RECT 111.580 172.210 111.840 172.530 ;
        RECT 111.640 170.830 111.780 172.210 ;
        RECT 111.580 170.510 111.840 170.830 ;
        RECT 110.660 169.830 110.920 170.150 ;
        RECT 109.740 167.110 110.000 167.430 ;
        RECT 108.820 166.770 109.080 167.090 ;
        RECT 104.680 166.430 104.940 166.750 ;
        RECT 106.060 166.430 106.320 166.750 ;
        RECT 103.760 164.390 104.020 164.710 ;
        RECT 104.740 164.690 104.880 166.430 ;
        RECT 105.140 164.730 105.400 165.050 ;
        RECT 104.280 164.550 104.880 164.690 ;
        RECT 104.280 162.330 104.420 164.550 ;
        RECT 104.220 162.010 104.480 162.330 ;
        RECT 104.280 153.230 104.420 162.010 ;
        RECT 105.200 159.465 105.340 164.730 ;
        RECT 106.120 163.690 106.260 166.430 ;
        RECT 108.880 165.050 109.020 166.770 ;
        RECT 108.820 164.730 109.080 165.050 ;
        RECT 110.720 164.905 110.860 169.830 ;
        RECT 110.650 164.535 110.930 164.905 ;
        RECT 112.100 164.690 112.240 177.310 ;
        RECT 111.640 164.550 112.240 164.690 ;
        RECT 108.810 163.855 109.090 164.225 ;
        RECT 108.820 163.710 109.080 163.855 ;
        RECT 106.060 163.370 106.320 163.690 ;
        RECT 105.880 162.835 107.420 163.205 ;
        RECT 106.980 160.990 107.240 161.310 ;
        RECT 109.740 160.990 110.000 161.310 ;
        RECT 107.040 159.950 107.180 160.990 ;
        RECT 106.980 159.630 107.240 159.950 ;
        RECT 105.130 159.095 105.410 159.465 ;
        RECT 109.800 159.270 109.940 160.990 ;
        RECT 105.140 158.950 105.400 159.095 ;
        RECT 108.360 158.950 108.620 159.270 ;
        RECT 108.820 158.950 109.080 159.270 ;
        RECT 109.740 158.950 110.000 159.270 ;
        RECT 105.880 157.395 107.420 157.765 ;
        RECT 107.900 153.510 108.160 153.830 ;
        RECT 104.280 153.090 105.340 153.230 ;
        RECT 104.220 152.490 104.480 152.810 ;
        RECT 102.900 151.730 103.500 151.870 ;
        RECT 102.900 145.670 103.040 151.730 ;
        RECT 104.280 150.770 104.420 152.490 ;
        RECT 103.750 150.255 104.030 150.625 ;
        RECT 104.220 150.450 104.480 150.770 ;
        RECT 103.300 148.070 103.560 148.390 ;
        RECT 103.360 146.350 103.500 148.070 ;
        RECT 103.300 146.030 103.560 146.350 ;
        RECT 102.840 145.350 103.100 145.670 ;
        RECT 103.820 142.350 103.960 150.255 ;
        RECT 104.680 142.630 104.940 142.950 ;
        RECT 102.900 142.210 103.960 142.350 ;
        RECT 102.380 137.190 102.640 137.510 ;
        RECT 102.900 132.410 103.040 142.210 ;
        RECT 104.220 141.950 104.480 142.270 ;
        RECT 103.760 141.610 104.020 141.930 ;
        RECT 103.300 140.590 103.560 140.910 ;
        RECT 103.360 137.850 103.500 140.590 ;
        RECT 103.300 137.530 103.560 137.850 ;
        RECT 102.840 132.090 103.100 132.410 ;
        RECT 101.000 128.690 101.260 129.010 ;
        RECT 101.460 125.970 101.720 126.290 ;
        RECT 100.540 125.290 100.800 125.610 ;
        RECT 100.600 124.590 100.740 125.290 ;
        RECT 100.540 124.270 100.800 124.590 ;
        RECT 101.000 122.570 101.260 122.890 ;
        RECT 101.060 121.530 101.200 122.570 ;
        RECT 101.000 121.210 101.260 121.530 ;
        RECT 98.240 120.870 98.500 121.190 ;
        RECT 100.080 120.870 100.340 121.190 ;
        RECT 96.860 120.530 97.120 120.850 ;
        RECT 96.920 117.450 97.060 120.530 ;
        RECT 97.780 120.190 98.040 120.510 ;
        RECT 97.320 119.850 97.580 120.170 ;
        RECT 97.380 117.790 97.520 119.850 ;
        RECT 97.840 119.150 97.980 120.190 ;
        RECT 97.780 118.830 98.040 119.150 ;
        RECT 97.320 117.470 97.580 117.790 ;
        RECT 96.860 117.130 97.120 117.450 ;
        RECT 94.100 115.770 94.360 116.090 ;
        RECT 97.840 115.410 97.980 118.830 ;
        RECT 98.300 116.430 98.440 120.870 ;
        RECT 99.160 117.130 99.420 117.450 ;
        RECT 98.240 116.110 98.500 116.430 ;
        RECT 97.780 115.090 98.040 115.410 ;
        RECT 98.240 113.390 98.500 113.710 ;
        RECT 92.720 112.370 92.980 112.690 ;
        RECT 93.640 112.030 93.900 112.350 ;
        RECT 96.860 112.030 97.120 112.350 ;
        RECT 91.800 111.690 92.060 112.010 ;
        RECT 91.340 110.330 91.600 110.650 ;
        RECT 89.950 107.415 90.230 107.785 ;
        RECT 90.020 107.250 90.160 107.415 ;
        RECT 91.400 107.250 91.540 110.330 ;
        RECT 89.960 106.930 90.220 107.250 ;
        RECT 91.340 106.930 91.600 107.250 ;
        RECT 90.020 106.480 90.160 106.930 ;
        RECT 90.020 106.340 91.080 106.480 ;
        RECT 89.090 105.715 90.630 106.085 ;
        RECT 90.940 105.550 91.080 106.340 ;
        RECT 90.880 105.230 91.140 105.550 ;
        RECT 90.870 101.975 91.150 102.345 ;
        RECT 89.090 100.275 90.630 100.645 ;
        RECT 90.940 100.110 91.080 101.975 ;
        RECT 90.880 99.790 91.140 100.110 ;
        RECT 90.870 99.255 91.150 99.625 ;
        RECT 91.400 99.340 91.540 106.930 ;
        RECT 91.860 106.570 92.000 111.690 ;
        RECT 93.180 108.970 93.440 109.290 ;
        RECT 93.240 108.270 93.380 108.970 ;
        RECT 93.180 107.950 93.440 108.270 ;
        RECT 93.700 107.250 93.840 112.030 ;
        RECT 96.920 110.990 97.060 112.030 ;
        RECT 97.780 111.690 98.040 112.010 ;
        RECT 96.400 110.670 96.660 110.990 ;
        RECT 96.860 110.670 97.120 110.990 ;
        RECT 96.460 109.970 96.600 110.670 ;
        RECT 97.840 110.310 97.980 111.690 ;
        RECT 97.780 109.990 98.040 110.310 ;
        RECT 96.400 109.650 96.660 109.970 ;
        RECT 93.640 106.930 93.900 107.250 ;
        RECT 92.720 106.590 92.980 106.910 ;
        RECT 91.800 106.250 92.060 106.570 ;
        RECT 91.860 101.470 92.000 106.250 ;
        RECT 92.780 104.530 92.920 106.590 ;
        RECT 96.460 105.210 96.600 109.650 ;
        RECT 98.300 107.250 98.440 113.390 ;
        RECT 99.220 107.250 99.360 117.130 ;
        RECT 100.140 115.410 100.280 120.870 ;
        RECT 100.540 117.470 100.800 117.790 ;
        RECT 100.080 115.090 100.340 115.410 ;
        RECT 100.600 110.310 100.740 117.470 ;
        RECT 101.060 115.750 101.200 121.210 ;
        RECT 101.000 115.430 101.260 115.750 ;
        RECT 101.000 113.390 101.260 113.710 ;
        RECT 101.060 110.310 101.200 113.390 ;
        RECT 100.540 109.990 100.800 110.310 ;
        RECT 101.000 109.990 101.260 110.310 ;
        RECT 100.540 108.970 100.800 109.290 ;
        RECT 96.860 106.990 97.120 107.250 ;
        RECT 96.860 106.930 97.520 106.990 ;
        RECT 98.240 106.930 98.500 107.250 ;
        RECT 99.160 106.930 99.420 107.250 ;
        RECT 96.920 106.850 97.520 106.930 ;
        RECT 96.860 106.250 97.120 106.570 ;
        RECT 96.400 104.890 96.660 105.210 ;
        RECT 93.180 104.550 93.440 104.870 ;
        RECT 92.720 104.210 92.980 104.530 ;
        RECT 93.240 102.830 93.380 104.550 ;
        RECT 94.560 103.530 94.820 103.850 ;
        RECT 95.940 103.530 96.200 103.850 ;
        RECT 93.180 102.510 93.440 102.830 ;
        RECT 91.800 101.150 92.060 101.470 ;
        RECT 91.800 99.340 92.060 99.430 ;
        RECT 90.880 99.110 91.140 99.255 ;
        RECT 91.400 99.200 92.060 99.340 ;
        RECT 91.800 99.110 92.060 99.200 ;
        RECT 90.880 97.070 91.140 97.390 ;
        RECT 88.580 96.730 88.840 97.050 ;
        RECT 88.120 96.390 88.380 96.710 ;
        RECT 84.900 96.050 85.160 96.370 ;
        RECT 85.820 94.010 86.080 94.330 ;
        RECT 85.880 93.650 86.020 94.010 ;
        RECT 88.180 93.990 88.320 96.390 ;
        RECT 89.090 94.835 90.630 95.205 ;
        RECT 88.120 93.670 88.380 93.990 ;
        RECT 89.500 93.670 89.760 93.990 ;
        RECT 85.820 93.330 86.080 93.650 ;
        RECT 86.740 93.330 87.000 93.650 ;
        RECT 85.880 91.950 86.020 93.330 ;
        RECT 85.820 91.630 86.080 91.950 ;
        RECT 85.360 89.930 85.620 90.250 ;
        RECT 85.420 88.550 85.560 89.930 ;
        RECT 86.800 89.230 86.940 93.330 ;
        RECT 89.560 91.950 89.700 93.670 ;
        RECT 89.960 92.650 90.220 92.970 ;
        RECT 89.500 91.630 89.760 91.950 ;
        RECT 90.020 91.270 90.160 92.650 ;
        RECT 90.940 91.950 91.080 97.070 ;
        RECT 93.180 96.390 93.440 96.710 ;
        RECT 91.340 95.710 91.600 96.030 ;
        RECT 91.400 94.330 91.540 95.710 ;
        RECT 91.800 95.370 92.060 95.690 ;
        RECT 91.340 94.010 91.600 94.330 ;
        RECT 90.880 91.630 91.140 91.950 ;
        RECT 89.960 90.950 90.220 91.270 ;
        RECT 91.860 90.930 92.000 95.370 ;
        RECT 92.720 92.650 92.980 92.970 ;
        RECT 92.780 91.270 92.920 92.650 ;
        RECT 92.720 90.950 92.980 91.270 ;
        RECT 91.800 90.610 92.060 90.930 ;
        RECT 89.090 89.395 90.630 89.765 ;
        RECT 86.740 88.910 87.000 89.230 ;
        RECT 85.360 88.230 85.620 88.550 ;
        RECT 90.880 88.230 91.140 88.550 ;
        RECT 86.280 87.210 86.540 87.530 ;
        RECT 86.340 85.830 86.480 87.210 ;
        RECT 86.280 85.510 86.540 85.830 ;
        RECT 85.820 85.170 86.080 85.490 ;
        RECT 85.880 83.790 86.020 85.170 ;
        RECT 87.660 84.490 87.920 84.810 ;
        RECT 85.820 83.470 86.080 83.790 ;
        RECT 87.720 83.450 87.860 84.490 ;
        RECT 89.090 83.955 90.630 84.325 ;
        RECT 90.940 83.790 91.080 88.230 ;
        RECT 93.240 87.870 93.380 96.390 ;
        RECT 94.100 96.225 94.360 96.370 ;
        RECT 94.090 95.855 94.370 96.225 ;
        RECT 93.640 95.370 93.900 95.690 ;
        RECT 93.700 93.310 93.840 95.370 ;
        RECT 93.640 92.990 93.900 93.310 ;
        RECT 93.180 87.550 93.440 87.870 ;
        RECT 90.880 83.470 91.140 83.790 ;
        RECT 87.660 83.130 87.920 83.450 ;
        RECT 92.720 83.130 92.980 83.450 ;
        RECT 92.780 81.070 92.920 83.130 ;
        RECT 92.720 80.750 92.980 81.070 ;
        RECT 79.840 79.730 80.100 80.050 ;
        RECT 82.600 79.730 82.860 80.050 ;
        RECT 83.060 79.730 83.320 80.050 ;
        RECT 83.520 79.730 83.780 80.050 ;
        RECT 87.200 79.730 87.460 80.050 ;
        RECT 88.580 79.730 88.840 80.050 ;
        RECT 79.900 78.010 80.040 79.730 ;
        RECT 83.120 78.350 83.260 79.730 ;
        RECT 83.520 79.050 83.780 79.370 ;
        RECT 83.060 78.030 83.320 78.350 ;
        RECT 83.580 78.010 83.720 79.050 ;
        RECT 79.380 77.690 79.640 78.010 ;
        RECT 79.840 77.690 80.100 78.010 ;
        RECT 83.520 77.690 83.780 78.010 ;
        RECT 76.160 77.440 76.820 77.580 ;
        RECT 76.160 77.350 76.420 77.440 ;
        RECT 75.240 76.670 75.500 76.990 ;
        RECT 75.300 75.630 75.440 76.670 ;
        RECT 75.240 75.310 75.500 75.630 ;
        RECT 75.760 74.950 75.900 77.350 ;
        RECT 76.160 76.670 76.420 76.990 ;
        RECT 76.220 75.630 76.360 76.670 ;
        RECT 76.160 75.310 76.420 75.630 ;
        RECT 75.700 74.630 75.960 74.950 ;
        RECT 75.760 74.350 75.900 74.630 ;
        RECT 74.840 74.210 75.900 74.350 ;
        RECT 76.160 74.290 76.420 74.610 ;
        RECT 74.320 73.610 74.580 73.930 ;
        RECT 68.340 72.590 68.600 72.910 ;
        RECT 70.640 72.590 70.900 72.910 ;
        RECT 63.740 72.250 64.000 72.570 ;
        RECT 74.840 72.230 74.980 74.210 ;
        RECT 75.700 73.840 75.960 73.930 ;
        RECT 75.300 73.700 75.960 73.840 ;
        RECT 62.820 71.910 63.080 72.230 ;
        RECT 74.780 71.910 75.040 72.230 ;
        RECT 72.300 70.355 73.840 70.725 ;
        RECT 74.840 70.190 74.980 71.910 ;
        RECT 75.300 71.210 75.440 73.700 ;
        RECT 75.700 73.610 75.960 73.700 ;
        RECT 75.700 71.910 75.960 72.230 ;
        RECT 75.240 70.890 75.500 71.210 ;
        RECT 69.720 69.870 69.980 70.190 ;
        RECT 74.780 69.870 75.040 70.190 ;
        RECT 61.440 68.850 61.700 69.170 ;
        RECT 60.520 67.150 60.780 67.470 ;
        RECT 61.500 66.790 61.640 68.850 ;
        RECT 69.780 68.830 69.920 69.870 ;
        RECT 71.100 69.530 71.360 69.850 ;
        RECT 69.720 68.510 69.980 68.830 ;
        RECT 68.340 68.170 68.600 68.490 ;
        RECT 70.640 68.170 70.900 68.490 ;
        RECT 68.400 66.790 68.540 68.170 ;
        RECT 70.700 66.790 70.840 68.170 ;
        RECT 71.160 66.790 71.300 69.530 ;
        RECT 74.840 69.170 74.980 69.870 ;
        RECT 74.780 68.850 75.040 69.170 ;
        RECT 74.780 68.170 75.040 68.490 ;
        RECT 57.760 66.470 58.020 66.790 ;
        RECT 59.600 66.470 59.860 66.790 ;
        RECT 60.060 66.470 60.320 66.790 ;
        RECT 61.440 66.470 61.700 66.790 ;
        RECT 67.420 66.470 67.680 66.790 ;
        RECT 68.340 66.470 68.600 66.790 ;
        RECT 70.640 66.470 70.900 66.790 ;
        RECT 71.100 66.470 71.360 66.790 ;
        RECT 54.540 66.130 54.800 66.450 ;
        RECT 55.000 66.130 55.260 66.450 ;
        RECT 54.600 64.830 54.740 66.130 ;
        RECT 54.140 64.690 54.740 64.830 ;
        RECT 52.700 63.410 52.960 63.730 ;
        RECT 53.160 63.070 53.420 63.390 ;
        RECT 53.220 58.030 53.360 63.070 ;
        RECT 54.140 60.330 54.280 64.690 ;
        RECT 54.540 64.090 54.800 64.410 ;
        RECT 54.600 61.350 54.740 64.090 ;
        RECT 55.060 61.350 55.200 66.130 ;
        RECT 60.980 65.450 61.240 65.770 ;
        RECT 57.300 63.410 57.560 63.730 ;
        RECT 55.510 62.195 57.050 62.565 ;
        RECT 54.540 61.030 54.800 61.350 ;
        RECT 55.000 61.030 55.260 61.350 ;
        RECT 53.620 60.010 53.880 60.330 ;
        RECT 54.080 60.010 54.340 60.330 ;
        RECT 53.680 58.630 53.820 60.010 ;
        RECT 53.620 58.310 53.880 58.630 ;
        RECT 53.220 57.890 53.820 58.030 ;
        RECT 53.680 56.220 53.820 57.890 ;
        RECT 55.510 56.755 57.050 57.125 ;
        RECT 57.360 56.500 57.500 63.410 ;
        RECT 61.040 61.350 61.180 65.450 ;
        RECT 65.120 63.410 65.380 63.730 ;
        RECT 61.900 61.710 62.160 62.030 ;
        RECT 60.980 61.030 61.240 61.350 ;
        RECT 59.600 60.690 59.860 61.010 ;
        RECT 59.660 59.310 59.800 60.690 ;
        RECT 59.600 58.990 59.860 59.310 ;
        RECT 59.140 57.970 59.400 58.290 ;
        RECT 56.440 56.360 57.500 56.500 ;
        RECT 56.440 56.220 56.580 56.360 ;
        RECT 59.200 56.220 59.340 57.970 ;
        RECT 61.960 56.220 62.100 61.710 ;
        RECT 64.660 61.030 64.920 61.350 ;
        RECT 64.720 56.220 64.860 61.030 ;
        RECT 65.180 59.310 65.320 63.410 ;
        RECT 66.960 60.010 67.220 60.330 ;
        RECT 65.120 58.990 65.380 59.310 ;
        RECT 67.020 58.630 67.160 60.010 ;
        RECT 66.960 58.310 67.220 58.630 ;
        RECT 67.480 56.220 67.620 66.470 ;
        RECT 68.340 65.450 68.600 65.770 ;
        RECT 69.720 65.450 69.980 65.770 ;
        RECT 71.100 65.450 71.360 65.770 ;
        RECT 68.400 58.290 68.540 65.450 ;
        RECT 69.780 61.350 69.920 65.450 ;
        RECT 71.160 64.070 71.300 65.450 ;
        RECT 72.300 64.915 73.840 65.285 ;
        RECT 74.840 64.750 74.980 68.170 ;
        RECT 75.300 66.790 75.440 70.890 ;
        RECT 75.760 69.510 75.900 71.910 ;
        RECT 75.700 69.190 75.960 69.510 ;
        RECT 75.240 66.470 75.500 66.790 ;
        RECT 76.220 66.450 76.360 74.290 ;
        RECT 76.680 69.170 76.820 77.440 ;
        RECT 77.540 77.350 77.800 77.670 ;
        RECT 77.600 75.290 77.740 77.350 ;
        RECT 79.440 77.330 79.580 77.690 ;
        RECT 87.260 77.670 87.400 79.730 ;
        RECT 88.640 78.350 88.780 79.730 ;
        RECT 93.240 79.710 93.380 87.550 ;
        RECT 93.180 79.390 93.440 79.710 ;
        RECT 89.090 78.515 90.630 78.885 ;
        RECT 94.160 78.350 94.300 95.855 ;
        RECT 88.580 78.030 88.840 78.350 ;
        RECT 94.100 78.030 94.360 78.350 ;
        RECT 85.820 77.350 86.080 77.670 ;
        RECT 87.200 77.350 87.460 77.670 ;
        RECT 92.260 77.350 92.520 77.670 ;
        RECT 78.920 77.010 79.180 77.330 ;
        RECT 79.380 77.010 79.640 77.330 ;
        RECT 77.540 74.970 77.800 75.290 ;
        RECT 78.980 74.610 79.120 77.010 ;
        RECT 78.920 74.290 79.180 74.610 ;
        RECT 79.440 72.310 79.580 77.010 ;
        RECT 81.680 76.670 81.940 76.990 ;
        RECT 80.300 74.970 80.560 75.290 ;
        RECT 79.440 72.230 80.040 72.310 ;
        RECT 79.440 72.170 80.100 72.230 ;
        RECT 79.840 71.910 80.100 72.170 ;
        RECT 80.360 69.850 80.500 74.970 ;
        RECT 81.740 74.610 81.880 76.670 ;
        RECT 85.880 75.630 86.020 77.350 ;
        RECT 92.320 75.630 92.460 77.350 ;
        RECT 85.820 75.310 86.080 75.630 ;
        RECT 92.260 75.310 92.520 75.630 ;
        RECT 81.680 74.290 81.940 74.610 ;
        RECT 83.980 74.290 84.240 74.610 ;
        RECT 90.880 74.290 91.140 74.610 ;
        RECT 93.640 74.290 93.900 74.610 ;
        RECT 84.040 73.930 84.180 74.290 ;
        RECT 88.580 73.950 88.840 74.270 ;
        RECT 83.520 73.610 83.780 73.930 ;
        RECT 83.980 73.610 84.240 73.930 ;
        RECT 83.580 72.570 83.720 73.610 ;
        RECT 84.040 72.910 84.180 73.610 ;
        RECT 83.980 72.590 84.240 72.910 ;
        RECT 83.520 72.250 83.780 72.570 ;
        RECT 87.200 71.910 87.460 72.230 ;
        RECT 83.980 70.890 84.240 71.210 ;
        RECT 80.300 69.530 80.560 69.850 ;
        RECT 80.360 69.170 80.500 69.530 ;
        RECT 84.040 69.170 84.180 70.890 ;
        RECT 87.260 70.190 87.400 71.910 ;
        RECT 88.640 70.190 88.780 73.950 ;
        RECT 89.090 73.075 90.630 73.445 ;
        RECT 90.940 72.910 91.080 74.290 ;
        RECT 90.880 72.590 91.140 72.910 ;
        RECT 90.880 71.910 91.140 72.230 ;
        RECT 87.200 69.870 87.460 70.190 ;
        RECT 88.580 69.870 88.840 70.190 ;
        RECT 87.650 69.335 87.930 69.705 ;
        RECT 87.720 69.170 87.860 69.335 ;
        RECT 76.620 69.025 76.880 69.170 ;
        RECT 76.610 68.655 76.890 69.025 ;
        RECT 80.300 68.850 80.560 69.170 ;
        RECT 83.980 68.850 84.240 69.170 ;
        RECT 87.660 68.850 87.920 69.170 ;
        RECT 78.920 68.510 79.180 68.830 ;
        RECT 78.000 68.170 78.260 68.490 ;
        RECT 78.060 66.790 78.200 68.170 ;
        RECT 78.980 66.790 79.120 68.510 ;
        RECT 83.520 68.170 83.780 68.490 ;
        RECT 78.000 66.470 78.260 66.790 ;
        RECT 78.920 66.470 79.180 66.790 ;
        RECT 76.160 66.130 76.420 66.450 ;
        RECT 76.160 65.450 76.420 65.770 ;
        RECT 76.620 65.450 76.880 65.770 ;
        RECT 74.780 64.430 75.040 64.750 ;
        RECT 71.100 63.750 71.360 64.070 ;
        RECT 70.180 63.410 70.440 63.730 ;
        RECT 74.320 63.410 74.580 63.730 ;
        RECT 75.240 63.410 75.500 63.730 ;
        RECT 69.720 61.030 69.980 61.350 ;
        RECT 68.340 57.970 68.600 58.290 ;
        RECT 70.240 56.220 70.380 63.410 ;
        RECT 72.300 59.475 73.840 59.845 ;
        RECT 74.380 58.630 74.520 63.410 ;
        RECT 75.300 61.690 75.440 63.410 ;
        RECT 75.700 61.710 75.960 62.030 ;
        RECT 75.240 61.370 75.500 61.690 ;
        RECT 74.320 58.310 74.580 58.630 ;
        RECT 72.940 57.970 73.200 58.290 ;
        RECT 73.000 56.220 73.140 57.970 ;
        RECT 75.760 56.220 75.900 61.710 ;
        RECT 76.220 58.290 76.360 65.450 ;
        RECT 76.680 61.350 76.820 65.450 ;
        RECT 78.980 63.390 79.120 66.470 ;
        RECT 83.580 66.110 83.720 68.170 ;
        RECT 84.440 67.150 84.700 67.470 ;
        RECT 83.520 65.790 83.780 66.110 ;
        RECT 79.380 65.450 79.640 65.770 ;
        RECT 81.220 65.450 81.480 65.770 ;
        RECT 79.440 63.730 79.580 65.450 ;
        RECT 79.380 63.410 79.640 63.730 ;
        RECT 78.920 63.070 79.180 63.390 ;
        RECT 76.620 61.030 76.880 61.350 ;
        RECT 80.300 61.030 80.560 61.350 ;
        RECT 76.160 57.970 76.420 58.290 ;
        RECT 78.460 57.970 78.720 58.290 ;
        RECT 80.360 58.030 80.500 61.030 ;
        RECT 81.280 58.630 81.420 65.450 ;
        RECT 84.500 63.730 84.640 67.150 ;
        RECT 87.720 66.450 87.860 68.850 ;
        RECT 88.120 68.510 88.380 68.830 ;
        RECT 88.180 66.450 88.320 68.510 ;
        RECT 87.660 66.130 87.920 66.450 ;
        RECT 88.120 66.130 88.380 66.450 ;
        RECT 83.520 63.640 83.780 63.730 ;
        RECT 83.520 63.500 84.180 63.640 ;
        RECT 83.520 63.410 83.780 63.500 ;
        RECT 81.220 58.310 81.480 58.630 ;
        RECT 78.520 56.220 78.660 57.970 ;
        RECT 80.360 57.890 81.420 58.030 ;
        RECT 81.280 56.220 81.420 57.890 ;
        RECT 84.040 56.220 84.180 63.500 ;
        RECT 84.440 63.410 84.700 63.730 ;
        RECT 87.660 63.410 87.920 63.730 ;
        RECT 84.900 62.730 85.160 63.050 ;
        RECT 85.820 62.730 86.080 63.050 ;
        RECT 84.960 61.350 85.100 62.730 ;
        RECT 84.900 61.030 85.160 61.350 ;
        RECT 85.880 58.290 86.020 62.730 ;
        RECT 87.720 61.350 87.860 63.410 ;
        RECT 88.640 61.350 88.780 69.870 ;
        RECT 89.490 68.655 89.770 69.025 ;
        RECT 89.500 68.510 89.760 68.655 ;
        RECT 90.940 68.490 91.080 71.910 ;
        RECT 91.340 71.570 91.600 71.890 ;
        RECT 91.400 70.190 91.540 71.570 ;
        RECT 91.340 69.870 91.600 70.190 ;
        RECT 93.700 69.850 93.840 74.290 ;
        RECT 94.620 73.670 94.760 103.530 ;
        RECT 96.000 102.830 96.140 103.530 ;
        RECT 96.920 102.830 97.060 106.250 ;
        RECT 95.940 102.510 96.200 102.830 ;
        RECT 96.860 102.510 97.120 102.830 ;
        RECT 96.860 101.380 97.120 101.470 ;
        RECT 97.380 101.380 97.520 106.850 ;
        RECT 98.300 104.950 98.440 106.930 ;
        RECT 99.220 105.550 99.360 106.930 ;
        RECT 100.080 106.590 100.340 106.910 ;
        RECT 100.140 105.550 100.280 106.590 ;
        RECT 99.160 105.230 99.420 105.550 ;
        RECT 100.080 105.230 100.340 105.550 ;
        RECT 97.840 104.810 98.440 104.950 ;
        RECT 97.840 104.530 97.980 104.810 ;
        RECT 97.780 104.210 98.040 104.530 ;
        RECT 98.240 104.210 98.500 104.530 ;
        RECT 97.840 102.150 97.980 104.210 ;
        RECT 98.300 102.490 98.440 104.210 ;
        RECT 98.240 102.170 98.500 102.490 ;
        RECT 97.780 101.830 98.040 102.150 ;
        RECT 96.860 101.240 97.520 101.380 ;
        RECT 96.860 101.150 97.120 101.240 ;
        RECT 95.020 100.810 95.280 101.130 ;
        RECT 95.080 99.770 95.220 100.810 ;
        RECT 96.920 99.770 97.060 101.150 ;
        RECT 95.020 99.450 95.280 99.770 ;
        RECT 96.860 99.450 97.120 99.770 ;
        RECT 97.840 99.340 97.980 101.830 ;
        RECT 99.220 101.720 99.360 105.230 ;
        RECT 100.080 104.780 100.340 104.870 ;
        RECT 100.600 104.780 100.740 108.970 ;
        RECT 101.000 106.930 101.260 107.250 ;
        RECT 101.060 104.870 101.200 106.930 ;
        RECT 100.080 104.640 100.740 104.780 ;
        RECT 100.080 104.550 100.340 104.640 ;
        RECT 101.000 104.550 101.260 104.870 ;
        RECT 101.520 102.150 101.660 125.970 ;
        RECT 101.920 120.530 102.180 120.850 ;
        RECT 101.980 118.470 102.120 120.530 ;
        RECT 101.920 118.150 102.180 118.470 ;
        RECT 101.980 113.030 102.120 118.150 ;
        RECT 101.920 112.710 102.180 113.030 ;
        RECT 102.900 110.650 103.040 132.090 ;
        RECT 103.360 131.050 103.500 137.530 ;
        RECT 103.820 136.490 103.960 141.610 ;
        RECT 104.280 139.890 104.420 141.950 ;
        RECT 104.220 139.570 104.480 139.890 ;
        RECT 104.220 138.890 104.480 139.210 ;
        RECT 103.760 136.170 104.020 136.490 ;
        RECT 104.280 132.070 104.420 138.890 ;
        RECT 104.740 138.190 104.880 142.630 ;
        RECT 104.680 137.870 104.940 138.190 ;
        RECT 105.200 132.070 105.340 153.090 ;
        RECT 105.880 151.955 107.420 152.325 ;
        RECT 107.960 151.790 108.100 153.510 ;
        RECT 107.900 151.470 108.160 151.790 ;
        RECT 106.520 151.130 106.780 151.450 ;
        RECT 106.580 150.770 106.720 151.130 ;
        RECT 106.050 150.255 106.330 150.625 ;
        RECT 106.520 150.450 106.780 150.770 ;
        RECT 107.890 150.255 108.170 150.625 ;
        RECT 106.060 150.110 106.320 150.255 ;
        RECT 107.900 150.110 108.160 150.255 ;
        RECT 108.420 149.150 108.560 158.950 ;
        RECT 108.880 158.590 109.020 158.950 ;
        RECT 109.280 158.610 109.540 158.930 ;
        RECT 108.820 158.270 109.080 158.590 ;
        RECT 108.880 156.890 109.020 158.270 ;
        RECT 108.820 156.570 109.080 156.890 ;
        RECT 108.880 151.450 109.020 156.570 ;
        RECT 109.340 156.210 109.480 158.610 ;
        RECT 109.740 156.230 110.000 156.550 ;
        RECT 109.280 155.890 109.540 156.210 ;
        RECT 108.820 151.130 109.080 151.450 ;
        RECT 107.960 149.010 108.560 149.150 ;
        RECT 107.960 147.790 108.100 149.010 ;
        RECT 108.360 148.070 108.620 148.390 ;
        RECT 107.500 147.650 108.100 147.790 ;
        RECT 107.500 147.370 107.640 147.650 ;
        RECT 107.440 147.050 107.700 147.370 ;
        RECT 105.880 146.515 107.420 146.885 ;
        RECT 107.960 144.650 108.100 147.650 ;
        RECT 108.420 146.350 108.560 148.070 ;
        RECT 108.360 146.030 108.620 146.350 ;
        RECT 108.350 145.495 108.630 145.865 ;
        RECT 108.420 145.330 108.560 145.495 ;
        RECT 108.880 145.330 109.020 151.130 ;
        RECT 109.340 151.110 109.480 155.890 ;
        RECT 109.800 154.170 109.940 156.230 ;
        RECT 110.200 155.210 110.460 155.530 ;
        RECT 109.740 153.850 110.000 154.170 ;
        RECT 109.280 150.790 109.540 151.110 ;
        RECT 109.340 145.670 109.480 150.790 ;
        RECT 110.260 150.770 110.400 155.210 ;
        RECT 110.200 150.450 110.460 150.770 ;
        RECT 109.280 145.350 109.540 145.670 ;
        RECT 110.720 145.330 110.860 164.535 ;
        RECT 111.110 156.375 111.390 156.745 ;
        RECT 108.360 145.010 108.620 145.330 ;
        RECT 108.820 145.010 109.080 145.330 ;
        RECT 109.740 145.010 110.000 145.330 ;
        RECT 110.660 145.010 110.920 145.330 ;
        RECT 107.900 144.330 108.160 144.650 ;
        RECT 108.820 144.330 109.080 144.650 ;
        RECT 107.900 141.610 108.160 141.930 ;
        RECT 105.880 141.075 107.420 141.445 ;
        RECT 107.960 139.890 108.100 141.610 ;
        RECT 107.900 139.570 108.160 139.890 ;
        RECT 106.060 138.890 106.320 139.210 ;
        RECT 106.120 137.510 106.260 138.890 ;
        RECT 108.360 137.870 108.620 138.190 ;
        RECT 106.060 137.190 106.320 137.510 ;
        RECT 107.900 137.190 108.160 137.510 ;
        RECT 105.880 135.635 107.420 136.005 ;
        RECT 107.960 135.470 108.100 137.190 ;
        RECT 107.900 135.150 108.160 135.470 ;
        RECT 108.420 134.450 108.560 137.870 ;
        RECT 108.360 134.130 108.620 134.450 ;
        RECT 108.420 132.750 108.560 134.130 ;
        RECT 108.880 134.110 109.020 144.330 ;
        RECT 109.800 143.630 109.940 145.010 ;
        RECT 109.740 143.310 110.000 143.630 ;
        RECT 109.280 142.970 109.540 143.290 ;
        RECT 109.340 139.550 109.480 142.970 ;
        RECT 111.180 142.950 111.320 156.375 ;
        RECT 111.640 155.870 111.780 164.550 ;
        RECT 112.040 160.650 112.300 160.970 ;
        RECT 111.580 155.550 111.840 155.870 ;
        RECT 111.120 142.630 111.380 142.950 ;
        RECT 111.580 142.290 111.840 142.610 ;
        RECT 110.200 140.590 110.460 140.910 ;
        RECT 109.740 140.250 110.000 140.570 ;
        RECT 109.280 139.230 109.540 139.550 ;
        RECT 109.340 134.450 109.480 139.230 ;
        RECT 109.800 137.850 109.940 140.250 ;
        RECT 110.260 139.890 110.400 140.590 ;
        RECT 111.640 139.890 111.780 142.290 ;
        RECT 110.200 139.570 110.460 139.890 ;
        RECT 111.580 139.570 111.840 139.890 ;
        RECT 111.120 139.230 111.380 139.550 ;
        RECT 109.740 137.530 110.000 137.850 ;
        RECT 109.280 134.130 109.540 134.450 ;
        RECT 108.820 133.790 109.080 134.110 ;
        RECT 108.360 132.430 108.620 132.750 ;
        RECT 104.220 131.750 104.480 132.070 ;
        RECT 105.140 131.750 105.400 132.070 ;
        RECT 107.900 131.070 108.160 131.390 ;
        RECT 103.300 130.730 103.560 131.050 ;
        RECT 105.140 130.730 105.400 131.050 ;
        RECT 104.220 128.350 104.480 128.670 ;
        RECT 104.280 127.310 104.420 128.350 ;
        RECT 104.220 126.990 104.480 127.310 ;
        RECT 105.200 126.630 105.340 130.730 ;
        RECT 105.880 130.195 107.420 130.565 ;
        RECT 107.440 128.010 107.700 128.330 ;
        RECT 107.500 126.970 107.640 128.010 ;
        RECT 107.440 126.650 107.700 126.970 ;
        RECT 105.140 126.310 105.400 126.630 ;
        RECT 105.880 124.755 107.420 125.125 ;
        RECT 107.960 123.570 108.100 131.070 ;
        RECT 103.760 123.250 104.020 123.570 ;
        RECT 107.900 123.250 108.160 123.570 ;
        RECT 103.820 119.150 103.960 123.250 ;
        RECT 104.680 122.570 104.940 122.890 ;
        RECT 104.740 121.530 104.880 122.570 ;
        RECT 104.680 121.210 104.940 121.530 ;
        RECT 108.360 120.190 108.620 120.510 ;
        RECT 107.900 119.850 108.160 120.170 ;
        RECT 105.880 119.315 107.420 119.685 ;
        RECT 103.760 118.830 104.020 119.150 ;
        RECT 105.140 118.830 105.400 119.150 ;
        RECT 104.680 112.030 104.940 112.350 ;
        RECT 104.740 110.990 104.880 112.030 ;
        RECT 104.680 110.670 104.940 110.990 ;
        RECT 102.840 110.330 103.100 110.650 ;
        RECT 105.200 107.930 105.340 118.830 ;
        RECT 107.960 118.130 108.100 119.850 ;
        RECT 108.420 118.130 108.560 120.190 ;
        RECT 107.900 117.810 108.160 118.130 ;
        RECT 108.360 117.810 108.620 118.130 ;
        RECT 105.880 113.875 107.420 114.245 ;
        RECT 105.600 111.690 105.860 112.010 ;
        RECT 105.660 110.310 105.800 111.690 ;
        RECT 105.600 109.990 105.860 110.310 ;
        RECT 105.880 108.435 107.420 108.805 ;
        RECT 108.880 108.465 109.020 133.790 ;
        RECT 109.340 132.410 109.480 134.130 ;
        RECT 109.280 132.090 109.540 132.410 ;
        RECT 109.740 131.410 110.000 131.730 ;
        RECT 109.800 129.010 109.940 131.410 ;
        RECT 109.740 128.690 110.000 129.010 ;
        RECT 109.740 128.010 110.000 128.330 ;
        RECT 109.800 126.630 109.940 128.010 ;
        RECT 109.740 126.310 110.000 126.630 ;
        RECT 110.660 126.310 110.920 126.630 ;
        RECT 110.720 124.590 110.860 126.310 ;
        RECT 110.660 124.270 110.920 124.590 ;
        RECT 110.200 122.910 110.460 123.230 ;
        RECT 110.260 121.870 110.400 122.910 ;
        RECT 110.200 121.550 110.460 121.870 ;
        RECT 109.740 117.470 110.000 117.790 ;
        RECT 109.280 115.090 109.540 115.410 ;
        RECT 109.340 113.710 109.480 115.090 ;
        RECT 109.280 113.390 109.540 113.710 ;
        RECT 109.340 110.310 109.480 113.390 ;
        RECT 109.280 109.990 109.540 110.310 ;
        RECT 109.800 109.290 109.940 117.470 ;
        RECT 110.660 114.410 110.920 114.730 ;
        RECT 110.720 113.710 110.860 114.410 ;
        RECT 110.660 113.390 110.920 113.710 ;
        RECT 109.280 108.970 109.540 109.290 ;
        RECT 109.740 108.970 110.000 109.290 ;
        RECT 111.180 109.030 111.320 139.230 ;
        RECT 111.640 138.190 111.780 139.570 ;
        RECT 112.100 139.550 112.240 160.650 ;
        RECT 112.560 150.430 112.700 187.655 ;
        RECT 112.960 185.130 113.220 185.450 ;
        RECT 113.020 183.410 113.160 185.130 ;
        RECT 113.480 183.750 113.620 191.590 ;
        RECT 113.420 183.430 113.680 183.750 ;
        RECT 112.960 183.090 113.220 183.410 ;
        RECT 113.940 170.150 114.080 194.570 ;
        RECT 114.400 194.290 114.540 199.840 ;
        RECT 114.800 199.750 115.060 199.840 ;
        RECT 115.780 199.730 115.920 208.250 ;
        RECT 137.400 208.230 137.540 212.220 ;
        RECT 134.580 207.910 134.840 208.230 ;
        RECT 137.340 207.910 137.600 208.230 ;
        RECT 122.160 207.570 122.420 207.890 ;
        RECT 117.100 207.230 117.360 207.550 ;
        RECT 116.180 206.890 116.440 207.210 ;
        RECT 116.240 204.830 116.380 206.890 ;
        RECT 116.180 204.510 116.440 204.830 ;
        RECT 116.640 204.510 116.900 204.830 ;
        RECT 115.720 199.410 115.980 199.730 ;
        RECT 114.800 196.010 115.060 196.330 ;
        RECT 114.860 194.290 115.000 196.010 ;
        RECT 115.780 194.290 115.920 199.410 ;
        RECT 116.700 197.350 116.840 204.510 ;
        RECT 117.160 199.390 117.300 207.230 ;
        RECT 122.220 205.510 122.360 207.570 ;
        RECT 131.820 206.890 132.080 207.210 ;
        RECT 132.740 206.890 133.000 207.210 ;
        RECT 127.680 205.530 127.940 205.850 ;
        RECT 122.160 205.190 122.420 205.510 ;
        RECT 122.220 202.790 122.360 205.190 ;
        RECT 127.740 204.830 127.880 205.530 ;
        RECT 129.060 205.190 129.320 205.510 ;
        RECT 127.680 204.510 127.940 204.830 ;
        RECT 126.760 204.170 127.020 204.490 ;
        RECT 127.220 204.170 127.480 204.490 ;
        RECT 122.670 203.635 124.210 204.005 ;
        RECT 126.820 203.130 126.960 204.170 ;
        RECT 126.760 202.810 127.020 203.130 ;
        RECT 122.160 202.470 122.420 202.790 ;
        RECT 120.320 201.790 120.580 202.110 ;
        RECT 120.380 199.730 120.520 201.790 ;
        RECT 121.240 201.450 121.500 201.770 ;
        RECT 121.300 200.070 121.440 201.450 ;
        RECT 121.700 200.430 121.960 200.750 ;
        RECT 121.240 199.750 121.500 200.070 ;
        RECT 120.320 199.410 120.580 199.730 ;
        RECT 117.100 199.300 117.360 199.390 ;
        RECT 117.100 199.160 117.760 199.300 ;
        RECT 117.100 199.070 117.360 199.160 ;
        RECT 116.640 197.030 116.900 197.350 ;
        RECT 114.340 193.970 114.600 194.290 ;
        RECT 114.800 193.970 115.060 194.290 ;
        RECT 115.720 193.970 115.980 194.290 ;
        RECT 114.860 181.030 115.000 193.970 ;
        RECT 116.700 191.910 116.840 197.030 ;
        RECT 116.640 191.590 116.900 191.910 ;
        RECT 117.100 191.590 117.360 191.910 ;
        RECT 116.180 190.570 116.440 190.890 ;
        RECT 116.240 188.850 116.380 190.570 ;
        RECT 117.160 189.870 117.300 191.590 ;
        RECT 117.100 189.550 117.360 189.870 ;
        RECT 116.180 188.530 116.440 188.850 ;
        RECT 116.640 185.810 116.900 186.130 ;
        RECT 116.700 181.710 116.840 185.810 ;
        RECT 116.640 181.390 116.900 181.710 ;
        RECT 114.800 180.710 115.060 181.030 ;
        RECT 114.860 175.250 115.000 180.710 ;
        RECT 115.260 177.650 115.520 177.970 ;
        RECT 115.320 176.270 115.460 177.650 ;
        RECT 115.260 175.950 115.520 176.270 ;
        RECT 114.800 174.930 115.060 175.250 ;
        RECT 114.340 174.250 114.600 174.570 ;
        RECT 114.400 170.830 114.540 174.250 ;
        RECT 114.340 170.510 114.600 170.830 ;
        RECT 113.880 169.830 114.140 170.150 ;
        RECT 116.640 169.490 116.900 169.810 ;
        RECT 114.340 168.810 114.600 169.130 ;
        RECT 114.400 164.710 114.540 168.810 ;
        RECT 116.700 167.430 116.840 169.490 ;
        RECT 116.640 167.110 116.900 167.430 ;
        RECT 117.620 166.750 117.760 199.160 ;
        RECT 118.480 196.690 118.740 197.010 ;
        RECT 118.540 194.290 118.680 196.690 ;
        RECT 120.380 195.310 120.520 199.410 ;
        RECT 121.760 199.390 121.900 200.430 ;
        RECT 126.820 200.070 126.960 202.810 ;
        RECT 127.280 202.790 127.420 204.170 ;
        RECT 127.740 203.470 127.880 204.510 ;
        RECT 127.680 203.150 127.940 203.470 ;
        RECT 129.120 202.790 129.260 205.190 ;
        RECT 131.360 204.850 131.620 205.170 ;
        RECT 129.980 204.170 130.240 204.490 ;
        RECT 127.220 202.470 127.480 202.790 ;
        RECT 129.060 202.470 129.320 202.790 ;
        RECT 130.040 201.770 130.180 204.170 ;
        RECT 127.220 201.450 127.480 201.770 ;
        RECT 129.980 201.450 130.240 201.770 ;
        RECT 130.900 201.450 131.160 201.770 ;
        RECT 127.280 200.750 127.420 201.450 ;
        RECT 127.220 200.430 127.480 200.750 ;
        RECT 127.680 200.090 127.940 200.410 ;
        RECT 124.460 199.750 124.720 200.070 ;
        RECT 126.760 199.750 127.020 200.070 ;
        RECT 121.700 199.070 121.960 199.390 ;
        RECT 120.320 194.990 120.580 195.310 ;
        RECT 121.760 194.290 121.900 199.070 ;
        RECT 122.670 198.195 124.210 198.565 ;
        RECT 124.520 194.970 124.660 199.750 ;
        RECT 126.300 199.410 126.560 199.730 ;
        RECT 126.360 195.310 126.500 199.410 ;
        RECT 126.300 194.990 126.560 195.310 ;
        RECT 124.460 194.650 124.720 194.970 ;
        RECT 118.480 193.970 118.740 194.290 ;
        RECT 121.700 193.970 121.960 194.290 ;
        RECT 124.520 193.950 124.660 194.650 ;
        RECT 124.460 193.630 124.720 193.950 ;
        RECT 126.300 193.630 126.560 193.950 ;
        RECT 122.670 192.755 124.210 193.125 ;
        RECT 125.840 190.910 126.100 191.230 ;
        RECT 123.540 190.570 123.800 190.890 ;
        RECT 123.600 188.170 123.740 190.570 ;
        RECT 125.900 188.850 126.040 190.910 ;
        RECT 126.360 189.190 126.500 193.630 ;
        RECT 127.220 193.290 127.480 193.610 ;
        RECT 126.760 192.270 127.020 192.590 ;
        RECT 126.300 188.870 126.560 189.190 ;
        RECT 124.460 188.530 124.720 188.850 ;
        RECT 125.380 188.530 125.640 188.850 ;
        RECT 125.840 188.530 126.100 188.850 ;
        RECT 123.540 187.850 123.800 188.170 ;
        RECT 122.670 187.315 124.210 187.685 ;
        RECT 123.080 186.150 123.340 186.470 ;
        RECT 124.520 186.380 124.660 188.530 ;
        RECT 125.440 186.810 125.580 188.530 ;
        RECT 125.380 186.490 125.640 186.810 ;
        RECT 124.060 186.240 124.660 186.380 ;
        RECT 121.700 185.810 121.960 186.130 ;
        RECT 118.480 185.470 118.740 185.790 ;
        RECT 118.020 169.830 118.280 170.150 ;
        RECT 118.080 168.110 118.220 169.830 ;
        RECT 118.020 167.790 118.280 168.110 ;
        RECT 117.560 166.430 117.820 166.750 ;
        RECT 117.620 165.390 117.760 166.430 ;
        RECT 117.560 165.070 117.820 165.390 ;
        RECT 114.340 164.620 114.600 164.710 ;
        RECT 114.340 164.480 115.000 164.620 ;
        RECT 114.340 164.390 114.600 164.480 ;
        RECT 114.340 160.650 114.600 160.970 ;
        RECT 114.400 159.610 114.540 160.650 ;
        RECT 114.340 159.290 114.600 159.610 ;
        RECT 113.420 159.180 113.680 159.270 ;
        RECT 113.020 159.040 113.680 159.180 ;
        RECT 112.500 150.110 112.760 150.430 ;
        RECT 113.020 146.350 113.160 159.040 ;
        RECT 113.420 158.950 113.680 159.040 ;
        RECT 114.860 158.930 115.000 164.480 ;
        RECT 114.800 158.610 115.060 158.930 ;
        RECT 113.420 156.230 113.680 156.550 ;
        RECT 113.480 154.510 113.620 156.230 ;
        RECT 113.420 154.190 113.680 154.510 ;
        RECT 114.860 153.490 115.000 158.610 ;
        RECT 118.540 156.210 118.680 185.470 ;
        RECT 120.780 185.130 121.040 185.450 ;
        RECT 120.840 182.730 120.980 185.130 ;
        RECT 121.240 183.090 121.500 183.410 ;
        RECT 120.780 182.410 121.040 182.730 ;
        RECT 121.300 181.710 121.440 183.090 ;
        RECT 121.760 183.070 121.900 185.810 ;
        RECT 123.140 183.410 123.280 186.150 ;
        RECT 124.060 184.430 124.200 186.240 ;
        RECT 124.920 186.150 125.180 186.470 ;
        RECT 124.460 185.130 124.720 185.450 ;
        RECT 124.000 184.110 124.260 184.430 ;
        RECT 124.520 183.410 124.660 185.130 ;
        RECT 124.980 184.430 125.120 186.150 ;
        RECT 124.920 184.110 125.180 184.430 ;
        RECT 124.980 183.410 125.120 184.110 ;
        RECT 123.080 183.090 123.340 183.410 ;
        RECT 124.460 183.090 124.720 183.410 ;
        RECT 124.920 183.090 125.180 183.410 ;
        RECT 121.700 182.750 121.960 183.070 ;
        RECT 122.670 181.875 124.210 182.245 ;
        RECT 126.820 181.710 126.960 192.270 ;
        RECT 127.280 189.870 127.420 193.290 ;
        RECT 127.740 191.570 127.880 200.090 ;
        RECT 128.140 196.690 128.400 197.010 ;
        RECT 128.200 195.310 128.340 196.690 ;
        RECT 128.140 194.990 128.400 195.310 ;
        RECT 130.440 194.990 130.700 195.310 ;
        RECT 130.500 192.670 130.640 194.990 ;
        RECT 130.960 194.970 131.100 201.450 ;
        RECT 131.420 199.585 131.560 204.850 ;
        RECT 131.350 199.215 131.630 199.585 ;
        RECT 131.420 197.350 131.560 199.215 ;
        RECT 131.360 197.030 131.620 197.350 ;
        RECT 131.880 196.670 132.020 206.890 ;
        RECT 132.800 205.170 132.940 206.890 ;
        RECT 132.740 204.850 133.000 205.170 ;
        RECT 132.280 202.810 132.540 203.130 ;
        RECT 133.660 202.810 133.920 203.130 ;
        RECT 132.340 199.730 132.480 202.810 ;
        RECT 133.200 202.470 133.460 202.790 ;
        RECT 132.740 201.790 133.000 202.110 ;
        RECT 132.800 200.070 132.940 201.790 ;
        RECT 132.740 199.750 133.000 200.070 ;
        RECT 132.280 199.410 132.540 199.730 ;
        RECT 132.740 198.730 133.000 199.050 ;
        RECT 131.820 196.350 132.080 196.670 ;
        RECT 131.360 196.010 131.620 196.330 ;
        RECT 130.900 194.650 131.160 194.970 ;
        RECT 130.900 193.290 131.160 193.610 ;
        RECT 130.040 192.530 130.640 192.670 ;
        RECT 127.680 191.250 127.940 191.570 ;
        RECT 127.680 190.570 127.940 190.890 ;
        RECT 127.220 189.550 127.480 189.870 ;
        RECT 127.740 186.470 127.880 190.570 ;
        RECT 129.520 188.870 129.780 189.190 ;
        RECT 129.060 188.190 129.320 188.510 ;
        RECT 128.140 186.830 128.400 187.150 ;
        RECT 127.680 186.150 127.940 186.470 ;
        RECT 127.220 185.810 127.480 186.130 ;
        RECT 127.280 184.090 127.420 185.810 ;
        RECT 127.220 183.770 127.480 184.090 ;
        RECT 121.240 181.390 121.500 181.710 ;
        RECT 126.760 181.390 127.020 181.710 ;
        RECT 126.300 180.710 126.560 181.030 ;
        RECT 124.460 176.970 124.720 177.290 ;
        RECT 122.670 176.435 124.210 176.805 ;
        RECT 124.520 175.590 124.660 176.970 ;
        RECT 122.160 175.270 122.420 175.590 ;
        RECT 124.460 175.270 124.720 175.590 ;
        RECT 124.920 175.270 125.180 175.590 ;
        RECT 118.940 174.930 119.200 175.250 ;
        RECT 120.320 174.930 120.580 175.250 ;
        RECT 119.000 173.210 119.140 174.930 ;
        RECT 118.940 172.890 119.200 173.210 ;
        RECT 120.380 167.430 120.520 174.930 ;
        RECT 121.700 172.890 121.960 173.210 ;
        RECT 120.780 171.530 121.040 171.850 ;
        RECT 120.320 167.110 120.580 167.430 ;
        RECT 120.840 166.750 120.980 171.530 ;
        RECT 121.760 169.130 121.900 172.890 ;
        RECT 122.220 172.530 122.360 175.270 ;
        RECT 124.000 174.930 124.260 175.250 ;
        RECT 124.060 173.550 124.200 174.930 ;
        RECT 124.000 173.230 124.260 173.550 ;
        RECT 124.520 172.870 124.660 175.270 ;
        RECT 124.460 172.550 124.720 172.870 ;
        RECT 124.980 172.530 125.120 175.270 ;
        RECT 126.360 173.210 126.500 180.710 ;
        RECT 126.760 177.310 127.020 177.630 ;
        RECT 126.820 173.210 126.960 177.310 ;
        RECT 126.300 172.890 126.560 173.210 ;
        RECT 126.760 172.890 127.020 173.210 ;
        RECT 128.200 172.950 128.340 186.830 ;
        RECT 129.120 186.470 129.260 188.190 ;
        RECT 129.580 188.170 129.720 188.870 ;
        RECT 129.520 187.850 129.780 188.170 ;
        RECT 129.060 186.150 129.320 186.470 ;
        RECT 130.040 185.390 130.180 192.530 ;
        RECT 130.440 191.930 130.700 192.250 ;
        RECT 130.500 189.870 130.640 191.930 ;
        RECT 130.960 191.910 131.100 193.290 ;
        RECT 130.900 191.590 131.160 191.910 ;
        RECT 130.440 189.550 130.700 189.870 ;
        RECT 130.440 188.530 130.700 188.850 ;
        RECT 130.500 188.170 130.640 188.530 ;
        RECT 130.440 187.850 130.700 188.170 ;
        RECT 130.960 185.790 131.100 191.590 ;
        RECT 131.420 190.890 131.560 196.010 ;
        RECT 131.360 190.570 131.620 190.890 ;
        RECT 132.280 189.210 132.540 189.530 ;
        RECT 131.360 185.810 131.620 186.130 ;
        RECT 130.900 185.470 131.160 185.790 ;
        RECT 130.040 185.250 130.640 185.390 ;
        RECT 129.980 184.110 130.240 184.430 ;
        RECT 130.040 181.370 130.180 184.110 ;
        RECT 130.500 181.710 130.640 185.250 ;
        RECT 130.440 181.390 130.700 181.710 ;
        RECT 129.980 181.050 130.240 181.370 ;
        RECT 131.420 181.030 131.560 185.810 ;
        RECT 132.340 181.030 132.480 189.210 ;
        RECT 132.800 187.150 132.940 198.730 ;
        RECT 133.260 195.310 133.400 202.470 ;
        RECT 133.720 200.410 133.860 202.810 ;
        RECT 134.640 201.770 134.780 207.910 ;
        RECT 137.800 207.570 138.060 207.890 ;
        RECT 135.960 204.170 136.220 204.490 ;
        RECT 134.580 201.450 134.840 201.770 ;
        RECT 135.500 201.450 135.760 201.770 ;
        RECT 135.560 200.750 135.700 201.450 ;
        RECT 135.500 200.430 135.760 200.750 ;
        RECT 133.660 200.090 133.920 200.410 ;
        RECT 136.020 199.730 136.160 204.170 ;
        RECT 137.340 202.470 137.600 202.790 ;
        RECT 136.880 201.790 137.140 202.110 ;
        RECT 136.420 200.265 136.680 200.410 ;
        RECT 136.410 199.895 136.690 200.265 ;
        RECT 134.580 199.640 134.840 199.730 ;
        RECT 135.960 199.640 136.220 199.730 ;
        RECT 134.580 199.500 136.220 199.640 ;
        RECT 134.580 199.410 134.840 199.500 ;
        RECT 135.960 199.410 136.220 199.500 ;
        RECT 136.940 199.050 137.080 201.790 ;
        RECT 134.580 198.730 134.840 199.050 ;
        RECT 136.880 198.730 137.140 199.050 ;
        RECT 134.640 197.350 134.780 198.730 ;
        RECT 136.940 197.350 137.080 198.730 ;
        RECT 134.580 197.030 134.840 197.350 ;
        RECT 136.880 197.030 137.140 197.350 ;
        RECT 133.200 194.990 133.460 195.310 ;
        RECT 134.640 194.630 134.780 197.030 ;
        RECT 137.400 195.390 137.540 202.470 ;
        RECT 137.860 201.770 138.000 207.570 ;
        RECT 139.460 206.355 141.000 206.725 ;
        RECT 138.260 205.530 138.520 205.850 ;
        RECT 138.320 203.470 138.460 205.530 ;
        RECT 141.940 205.190 142.200 205.510 ;
        RECT 140.560 204.850 140.820 205.170 ;
        RECT 140.620 203.470 140.760 204.850 ;
        RECT 138.260 203.150 138.520 203.470 ;
        RECT 140.560 203.150 140.820 203.470 ;
        RECT 137.800 201.450 138.060 201.770 ;
        RECT 137.800 200.430 138.060 200.750 ;
        RECT 137.860 200.265 138.000 200.430 ;
        RECT 137.790 199.895 138.070 200.265 ;
        RECT 138.320 197.350 138.460 203.150 ;
        RECT 141.480 202.130 141.740 202.450 ;
        RECT 138.720 201.450 138.980 201.770 ;
        RECT 138.780 198.030 138.920 201.450 ;
        RECT 139.460 200.915 141.000 201.285 ;
        RECT 141.540 200.150 141.680 202.130 ;
        RECT 140.100 199.750 140.360 200.070 ;
        RECT 140.620 200.010 141.680 200.150 ;
        RECT 140.160 199.585 140.300 199.750 ;
        RECT 140.620 199.730 140.760 200.010 ;
        RECT 140.090 199.215 140.370 199.585 ;
        RECT 140.560 199.410 140.820 199.730 ;
        RECT 142.000 199.390 142.140 205.190 ;
        RECT 142.400 202.130 142.660 202.450 ;
        RECT 141.480 199.070 141.740 199.390 ;
        RECT 141.940 199.070 142.200 199.390 ;
        RECT 141.540 198.030 141.680 199.070 ;
        RECT 138.720 197.710 138.980 198.030 ;
        RECT 141.480 197.710 141.740 198.030 ;
        RECT 138.260 197.030 138.520 197.350 ;
        RECT 141.480 197.030 141.740 197.350 ;
        RECT 139.460 195.475 141.000 195.845 ;
        RECT 137.400 195.250 138.920 195.390 ;
        RECT 141.540 195.310 141.680 197.030 ;
        RECT 134.580 194.310 134.840 194.630 ;
        RECT 133.660 193.970 133.920 194.290 ;
        RECT 135.040 193.970 135.300 194.290 ;
        RECT 137.400 194.030 137.540 195.250 ;
        RECT 137.800 194.650 138.060 194.970 ;
        RECT 137.860 194.290 138.000 194.650 ;
        RECT 133.200 193.630 133.460 193.950 ;
        RECT 133.260 191.910 133.400 193.630 ;
        RECT 133.720 191.910 133.860 193.970 ;
        RECT 135.100 191.910 135.240 193.970 ;
        RECT 136.940 193.950 137.540 194.030 ;
        RECT 137.800 193.970 138.060 194.290 ;
        RECT 136.880 193.890 137.540 193.950 ;
        RECT 136.880 193.630 137.140 193.890 ;
        RECT 137.400 191.910 137.540 193.890 ;
        RECT 137.860 192.590 138.000 193.970 ;
        RECT 138.780 193.950 138.920 195.250 ;
        RECT 141.020 194.990 141.280 195.310 ;
        RECT 141.480 194.990 141.740 195.310 ;
        RECT 141.080 194.710 141.220 194.990 ;
        RECT 142.000 194.710 142.140 199.070 ;
        RECT 140.620 194.570 142.140 194.710 ;
        RECT 138.720 193.630 138.980 193.950 ;
        RECT 138.260 193.290 138.520 193.610 ;
        RECT 139.180 193.290 139.440 193.610 ;
        RECT 137.800 192.270 138.060 192.590 ;
        RECT 138.320 192.250 138.460 193.290 ;
        RECT 138.260 191.930 138.520 192.250 ;
        RECT 133.200 191.590 133.460 191.910 ;
        RECT 133.660 191.590 133.920 191.910 ;
        RECT 134.120 191.590 134.380 191.910 ;
        RECT 135.040 191.590 135.300 191.910 ;
        RECT 137.340 191.590 137.600 191.910 ;
        RECT 133.260 189.190 133.400 191.590 ;
        RECT 133.720 189.870 133.860 191.590 ;
        RECT 133.660 189.550 133.920 189.870 ;
        RECT 133.200 188.870 133.460 189.190 ;
        RECT 134.180 188.850 134.320 191.590 ;
        RECT 134.120 188.530 134.380 188.850 ;
        RECT 135.100 188.170 135.240 191.590 ;
        RECT 139.240 191.310 139.380 193.290 ;
        RECT 140.620 192.250 140.760 194.570 ;
        RECT 141.020 193.630 141.280 193.950 ;
        RECT 141.080 192.590 141.220 193.630 ;
        RECT 141.020 192.270 141.280 192.590 ;
        RECT 140.560 191.930 140.820 192.250 ;
        RECT 138.780 191.230 139.380 191.310 ;
        RECT 138.780 191.170 139.440 191.230 ;
        RECT 138.780 188.850 138.920 191.170 ;
        RECT 139.180 190.910 139.440 191.170 ;
        RECT 139.460 190.035 141.000 190.405 ;
        RECT 138.720 188.530 138.980 188.850 ;
        RECT 135.040 187.850 135.300 188.170 ;
        RECT 138.780 187.150 138.920 188.530 ;
        RECT 140.100 188.190 140.360 188.510 ;
        RECT 132.740 186.830 133.000 187.150 ;
        RECT 138.720 186.830 138.980 187.150 ;
        RECT 138.720 186.150 138.980 186.470 ;
        RECT 136.880 185.130 137.140 185.450 ;
        RECT 136.940 183.410 137.080 185.130 ;
        RECT 138.780 184.430 138.920 186.150 ;
        RECT 140.160 185.450 140.300 188.190 ;
        RECT 141.480 185.470 141.740 185.790 ;
        RECT 140.100 185.130 140.360 185.450 ;
        RECT 139.460 184.595 141.000 184.965 ;
        RECT 138.720 184.110 138.980 184.430 ;
        RECT 140.100 184.110 140.360 184.430 ;
        RECT 136.880 183.090 137.140 183.410 ;
        RECT 136.880 182.410 137.140 182.730 ;
        RECT 136.940 181.710 137.080 182.410 ;
        RECT 133.660 181.390 133.920 181.710 ;
        RECT 136.880 181.390 137.140 181.710 ;
        RECT 131.360 180.710 131.620 181.030 ;
        RECT 132.280 180.710 132.540 181.030 ;
        RECT 128.600 180.370 128.860 180.690 ;
        RECT 131.820 180.370 132.080 180.690 ;
        RECT 128.660 177.630 128.800 180.370 ;
        RECT 131.880 178.990 132.020 180.370 ;
        RECT 131.820 178.670 132.080 178.990 ;
        RECT 130.900 178.330 131.160 178.650 ;
        RECT 128.600 177.310 128.860 177.630 ;
        RECT 130.960 176.270 131.100 178.330 ;
        RECT 130.900 175.950 131.160 176.270 ;
        RECT 129.060 175.610 129.320 175.930 ;
        RECT 128.200 172.810 128.800 172.950 ;
        RECT 122.160 172.210 122.420 172.530 ;
        RECT 124.920 172.210 125.180 172.530 ;
        RECT 125.380 172.210 125.640 172.530 ;
        RECT 124.460 171.870 124.720 172.190 ;
        RECT 122.670 170.995 124.210 171.365 ;
        RECT 124.520 169.470 124.660 171.870 ;
        RECT 124.980 170.830 125.120 172.210 ;
        RECT 125.440 171.850 125.580 172.210 ;
        RECT 128.140 171.870 128.400 172.190 ;
        RECT 125.380 171.530 125.640 171.850 ;
        RECT 124.920 170.510 125.180 170.830 ;
        RECT 128.200 169.810 128.340 171.870 ;
        RECT 128.140 169.490 128.400 169.810 ;
        RECT 124.460 169.150 124.720 169.470 ;
        RECT 121.700 168.810 121.960 169.130 ;
        RECT 120.780 166.430 121.040 166.750 ;
        RECT 122.670 165.555 124.210 165.925 ;
        RECT 128.660 165.050 128.800 172.810 ;
        RECT 129.120 172.530 129.260 175.610 ;
        RECT 130.900 175.270 131.160 175.590 ;
        RECT 130.440 174.930 130.700 175.250 ;
        RECT 129.060 172.210 129.320 172.530 ;
        RECT 129.520 171.530 129.780 171.850 ;
        RECT 129.580 170.830 129.720 171.530 ;
        RECT 129.520 170.510 129.780 170.830 ;
        RECT 130.500 170.150 130.640 174.930 ;
        RECT 130.960 171.850 131.100 175.270 ;
        RECT 133.200 174.250 133.460 174.570 ;
        RECT 133.260 172.190 133.400 174.250 ;
        RECT 133.200 171.870 133.460 172.190 ;
        RECT 130.900 171.530 131.160 171.850 ;
        RECT 130.960 170.490 131.100 171.530 ;
        RECT 130.900 170.170 131.160 170.490 ;
        RECT 130.440 169.830 130.700 170.150 ;
        RECT 131.360 169.830 131.620 170.150 ;
        RECT 131.420 169.130 131.560 169.830 ;
        RECT 131.360 168.810 131.620 169.130 ;
        RECT 131.820 166.770 132.080 167.090 ;
        RECT 132.740 166.770 133.000 167.090 ;
        RECT 128.600 164.730 128.860 165.050 ;
        RECT 120.780 164.390 121.040 164.710 ;
        RECT 131.360 164.390 131.620 164.710 ;
        RECT 120.840 162.670 120.980 164.390 ;
        RECT 127.220 164.050 127.480 164.370 ;
        RECT 124.000 163.370 124.260 163.690 ;
        RECT 120.780 162.350 121.040 162.670 ;
        RECT 121.700 161.670 121.960 161.990 ;
        RECT 120.780 161.330 121.040 161.650 ;
        RECT 118.940 160.650 119.200 160.970 ;
        RECT 119.000 158.250 119.140 160.650 ;
        RECT 120.840 159.950 120.980 161.330 ;
        RECT 120.780 159.630 121.040 159.950 ;
        RECT 121.760 158.590 121.900 161.670 ;
        RECT 124.060 161.650 124.200 163.370 ;
        RECT 122.160 161.330 122.420 161.650 ;
        RECT 124.000 161.330 124.260 161.650 ;
        RECT 125.380 161.330 125.640 161.650 ;
        RECT 126.300 161.330 126.560 161.650 ;
        RECT 122.220 159.270 122.360 161.330 ;
        RECT 124.920 160.990 125.180 161.310 ;
        RECT 122.670 160.115 124.210 160.485 ;
        RECT 124.980 159.950 125.120 160.990 ;
        RECT 125.440 159.950 125.580 161.330 ;
        RECT 124.920 159.630 125.180 159.950 ;
        RECT 125.380 159.630 125.640 159.950 ;
        RECT 126.360 159.860 126.500 161.330 ;
        RECT 126.760 159.860 127.020 159.950 ;
        RECT 126.360 159.720 127.020 159.860 ;
        RECT 126.760 159.630 127.020 159.720 ;
        RECT 122.160 158.950 122.420 159.270 ;
        RECT 121.700 158.270 121.960 158.590 ;
        RECT 118.940 157.930 119.200 158.250 ;
        RECT 118.480 155.890 118.740 156.210 ;
        RECT 119.000 155.870 119.140 157.930 ;
        RECT 119.400 157.140 119.660 157.230 ;
        RECT 119.400 157.000 120.520 157.140 ;
        RECT 119.400 156.910 119.660 157.000 ;
        RECT 116.180 155.550 116.440 155.870 ;
        RECT 118.940 155.550 119.200 155.870 ;
        RECT 114.800 153.170 115.060 153.490 ;
        RECT 114.860 150.770 115.000 153.170 ;
        RECT 116.240 151.020 116.380 155.550 ;
        RECT 117.100 155.210 117.360 155.530 ;
        RECT 116.240 150.880 116.840 151.020 ;
        RECT 114.800 150.450 115.060 150.770 ;
        RECT 114.340 147.110 114.600 147.370 ;
        RECT 114.860 147.110 115.000 150.450 ;
        RECT 115.260 150.110 115.520 150.430 ;
        RECT 115.320 148.390 115.460 150.110 ;
        RECT 115.260 148.070 115.520 148.390 ;
        RECT 114.340 147.050 115.000 147.110 ;
        RECT 114.400 146.970 115.000 147.050 ;
        RECT 112.960 146.030 113.220 146.350 ;
        RECT 112.040 139.230 112.300 139.550 ;
        RECT 111.580 137.870 111.840 138.190 ;
        RECT 113.020 131.980 113.160 146.030 ;
        RECT 114.860 145.330 115.000 146.970 ;
        RECT 114.800 145.010 115.060 145.330 ;
        RECT 114.860 139.890 115.000 145.010 ;
        RECT 114.800 139.570 115.060 139.890 ;
        RECT 115.320 139.120 115.460 148.070 ;
        RECT 115.720 147.050 115.980 147.370 ;
        RECT 115.780 142.950 115.920 147.050 ;
        RECT 116.700 143.710 116.840 150.880 ;
        RECT 117.160 144.990 117.300 155.210 ;
        RECT 119.000 154.510 119.140 155.550 ;
        RECT 118.940 154.190 119.200 154.510 ;
        RECT 117.100 144.670 117.360 144.990 ;
        RECT 116.700 143.570 117.300 143.710 ;
        RECT 115.720 142.630 115.980 142.950 ;
        RECT 116.640 142.180 116.900 142.270 ;
        RECT 117.160 142.180 117.300 143.570 ;
        RECT 119.460 142.950 119.600 156.910 ;
        RECT 120.380 156.550 120.520 157.000 ;
        RECT 120.320 156.230 120.580 156.550 ;
        RECT 120.780 155.890 121.040 156.210 ;
        RECT 120.840 151.790 120.980 155.890 ;
        RECT 122.220 155.870 122.360 158.950 ;
        RECT 127.280 158.590 127.420 164.050 ;
        RECT 130.440 163.710 130.700 164.030 ;
        RECT 130.900 163.710 131.160 164.030 ;
        RECT 129.520 162.010 129.780 162.330 ;
        RECT 129.580 161.310 129.720 162.010 ;
        RECT 129.980 161.330 130.240 161.650 ;
        RECT 130.500 161.390 130.640 163.710 ;
        RECT 130.960 162.330 131.100 163.710 ;
        RECT 130.900 162.010 131.160 162.330 ;
        RECT 129.520 160.990 129.780 161.310 ;
        RECT 127.220 158.270 127.480 158.590 ;
        RECT 128.600 156.230 128.860 156.550 ;
        RECT 125.380 155.950 125.640 156.210 ;
        RECT 125.380 155.890 126.500 155.950 ;
        RECT 127.220 155.890 127.480 156.210 ;
        RECT 128.140 155.890 128.400 156.210 ;
        RECT 125.440 155.870 126.500 155.890 ;
        RECT 122.160 155.550 122.420 155.870 ;
        RECT 125.440 155.810 126.560 155.870 ;
        RECT 126.300 155.550 126.560 155.810 ;
        RECT 124.920 155.210 125.180 155.530 ;
        RECT 125.380 155.210 125.640 155.530 ;
        RECT 122.670 154.675 124.210 155.045 ;
        RECT 124.980 154.170 125.120 155.210 ;
        RECT 125.440 154.510 125.580 155.210 ;
        RECT 125.380 154.190 125.640 154.510 ;
        RECT 124.920 153.850 125.180 154.170 ;
        RECT 120.780 151.470 121.040 151.790 ;
        RECT 125.840 150.450 126.100 150.770 ;
        RECT 125.380 150.110 125.640 150.430 ;
        RECT 122.160 149.770 122.420 150.090 ;
        RECT 122.220 149.070 122.360 149.770 ;
        RECT 122.670 149.235 124.210 149.605 ;
        RECT 122.160 148.750 122.420 149.070 ;
        RECT 124.460 147.730 124.720 148.050 ;
        RECT 124.520 147.370 124.660 147.730 ;
        RECT 125.440 147.370 125.580 150.110 ;
        RECT 124.460 147.050 124.720 147.370 ;
        RECT 125.380 147.050 125.640 147.370 ;
        RECT 124.520 145.330 124.660 147.050 ;
        RECT 125.900 146.350 126.040 150.450 ;
        RECT 126.300 148.750 126.560 149.070 ;
        RECT 126.760 148.750 127.020 149.070 ;
        RECT 125.840 146.030 126.100 146.350 ;
        RECT 124.460 145.010 124.720 145.330 ;
        RECT 125.840 145.010 126.100 145.330 ;
        RECT 122.670 143.795 124.210 144.165 ;
        RECT 125.900 143.290 126.040 145.010 ;
        RECT 125.840 142.970 126.100 143.290 ;
        RECT 118.480 142.630 118.740 142.950 ;
        RECT 119.400 142.630 119.660 142.950 ;
        RECT 121.700 142.630 121.960 142.950 ;
        RECT 124.920 142.630 125.180 142.950 ;
        RECT 116.640 142.040 117.300 142.180 ;
        RECT 116.640 141.950 116.900 142.040 ;
        RECT 116.180 139.230 116.440 139.550 ;
        RECT 114.860 138.980 115.460 139.120 ;
        RECT 113.880 136.170 114.140 136.490 ;
        RECT 113.940 134.450 114.080 136.170 ;
        RECT 113.880 134.130 114.140 134.450 ;
        RECT 113.420 131.980 113.680 132.070 ;
        RECT 113.020 131.840 113.680 131.980 ;
        RECT 113.020 124.250 113.160 131.840 ;
        RECT 113.420 131.750 113.680 131.840 ;
        RECT 114.340 130.730 114.600 131.050 ;
        RECT 113.420 125.290 113.680 125.610 ;
        RECT 112.960 123.930 113.220 124.250 ;
        RECT 113.480 123.570 113.620 125.290 ;
        RECT 112.500 123.250 112.760 123.570 ;
        RECT 113.420 123.480 113.680 123.570 ;
        RECT 113.020 123.340 113.680 123.480 ;
        RECT 112.560 115.750 112.700 123.250 ;
        RECT 113.020 118.130 113.160 123.340 ;
        RECT 113.420 123.250 113.680 123.340 ;
        RECT 114.400 122.890 114.540 130.730 ;
        RECT 114.860 123.570 115.000 138.980 ;
        RECT 116.240 134.450 116.380 139.230 ;
        RECT 116.640 136.170 116.900 136.490 ;
        RECT 116.180 134.130 116.440 134.450 ;
        RECT 116.240 132.070 116.380 134.130 ;
        RECT 116.700 132.070 116.840 136.170 ;
        RECT 117.160 133.680 117.300 142.040 ;
        RECT 117.560 141.610 117.820 141.930 ;
        RECT 117.620 134.450 117.760 141.610 ;
        RECT 117.560 134.130 117.820 134.450 ;
        RECT 117.160 133.540 117.760 133.680 ;
        RECT 116.180 131.750 116.440 132.070 ;
        RECT 116.640 131.750 116.900 132.070 ;
        RECT 117.620 124.250 117.760 133.540 ;
        RECT 117.560 123.930 117.820 124.250 ;
        RECT 114.800 123.250 115.060 123.570 ;
        RECT 115.260 122.910 115.520 123.230 ;
        RECT 114.340 122.570 114.600 122.890 ;
        RECT 114.400 121.870 114.540 122.570 ;
        RECT 114.340 121.550 114.600 121.870 ;
        RECT 112.960 117.810 113.220 118.130 ;
        RECT 112.500 115.660 112.760 115.750 ;
        RECT 112.100 115.520 112.760 115.660 ;
        RECT 111.580 112.030 111.840 112.350 ;
        RECT 108.810 108.095 109.090 108.465 ;
        RECT 105.140 107.610 105.400 107.930 ;
        RECT 108.820 107.270 109.080 107.590 ;
        RECT 105.140 106.930 105.400 107.250 ;
        RECT 105.200 105.550 105.340 106.930 ;
        RECT 106.050 106.735 106.330 107.105 ;
        RECT 106.120 106.570 106.260 106.735 ;
        RECT 106.060 106.250 106.320 106.570 ;
        RECT 105.140 105.230 105.400 105.550 ;
        RECT 108.880 104.530 109.020 107.270 ;
        RECT 109.340 107.250 109.480 108.970 ;
        RECT 109.800 107.930 109.940 108.970 ;
        RECT 110.720 108.890 111.320 109.030 ;
        RECT 109.740 107.610 110.000 107.930 ;
        RECT 109.280 106.930 109.540 107.250 ;
        RECT 109.740 106.250 110.000 106.570 ;
        RECT 109.800 105.210 109.940 106.250 ;
        RECT 109.740 104.890 110.000 105.210 ;
        RECT 110.720 104.870 110.860 108.890 ;
        RECT 111.110 108.095 111.390 108.465 ;
        RECT 111.180 107.250 111.320 108.095 ;
        RECT 111.120 106.930 111.380 107.250 ;
        RECT 111.640 105.550 111.780 112.030 ;
        RECT 112.100 109.970 112.240 115.520 ;
        RECT 112.500 115.430 112.760 115.520 ;
        RECT 114.400 112.010 114.540 121.550 ;
        RECT 115.320 121.530 115.460 122.910 ;
        RECT 115.260 121.210 115.520 121.530 ;
        RECT 114.800 115.430 115.060 115.750 ;
        RECT 114.860 113.710 115.000 115.430 ;
        RECT 114.800 113.390 115.060 113.710 ;
        RECT 115.320 112.690 115.460 121.210 ;
        RECT 116.640 120.190 116.900 120.510 ;
        RECT 116.700 118.130 116.840 120.190 ;
        RECT 116.640 117.810 116.900 118.130 ;
        RECT 116.180 117.470 116.440 117.790 ;
        RECT 116.240 116.430 116.380 117.470 ;
        RECT 116.180 116.110 116.440 116.430 ;
        RECT 118.540 116.090 118.680 142.630 ;
        RECT 121.760 138.190 121.900 142.630 ;
        RECT 124.980 139.890 125.120 142.630 ;
        RECT 124.920 139.570 125.180 139.890 ;
        RECT 124.980 139.210 125.120 139.570 ;
        RECT 124.920 138.890 125.180 139.210 ;
        RECT 122.670 138.355 124.210 138.725 ;
        RECT 121.700 137.870 121.960 138.190 ;
        RECT 124.980 137.850 125.120 138.890 ;
        RECT 124.920 137.530 125.180 137.850 ;
        RECT 118.940 137.190 119.200 137.510 ;
        RECT 119.000 134.450 119.140 137.190 ;
        RECT 121.240 136.850 121.500 137.170 ;
        RECT 125.380 136.850 125.640 137.170 ;
        RECT 118.940 134.130 119.200 134.450 ;
        RECT 121.300 132.750 121.440 136.850 ;
        RECT 125.440 134.450 125.580 136.850 ;
        RECT 125.380 134.130 125.640 134.450 ;
        RECT 125.840 134.130 126.100 134.450 ;
        RECT 125.440 133.770 125.580 134.130 ;
        RECT 125.380 133.450 125.640 133.770 ;
        RECT 122.670 132.915 124.210 133.285 ;
        RECT 121.240 132.430 121.500 132.750 ;
        RECT 125.440 132.070 125.580 133.450 ;
        RECT 125.380 131.750 125.640 132.070 ;
        RECT 125.900 131.730 126.040 134.130 ;
        RECT 125.840 131.410 126.100 131.730 ;
        RECT 125.380 128.350 125.640 128.670 ;
        RECT 122.670 127.475 124.210 127.845 ;
        RECT 125.440 126.630 125.580 128.350 ;
        RECT 126.360 126.630 126.500 148.750 ;
        RECT 126.820 148.390 126.960 148.750 ;
        RECT 127.280 148.390 127.420 155.890 ;
        RECT 127.680 155.210 127.940 155.530 ;
        RECT 126.760 148.070 127.020 148.390 ;
        RECT 127.220 148.070 127.480 148.390 ;
        RECT 127.740 148.300 127.880 155.210 ;
        RECT 128.200 154.510 128.340 155.890 ;
        RECT 128.140 154.190 128.400 154.510 ;
        RECT 128.660 154.170 128.800 156.230 ;
        RECT 129.580 156.210 129.720 160.990 ;
        RECT 130.040 159.610 130.180 161.330 ;
        RECT 130.500 161.250 131.100 161.390 ;
        RECT 129.980 159.290 130.240 159.610 ;
        RECT 130.040 156.210 130.180 159.290 ;
        RECT 130.440 156.910 130.700 157.230 ;
        RECT 129.520 155.890 129.780 156.210 ;
        RECT 129.980 155.890 130.240 156.210 ;
        RECT 128.600 153.850 128.860 154.170 ;
        RECT 130.500 153.830 130.640 156.910 ;
        RECT 130.440 153.510 130.700 153.830 ;
        RECT 130.500 151.450 130.640 153.510 ;
        RECT 130.440 151.130 130.700 151.450 ;
        RECT 129.060 149.770 129.320 150.090 ;
        RECT 128.600 148.410 128.860 148.730 ;
        RECT 128.140 148.300 128.400 148.390 ;
        RECT 127.740 148.160 128.400 148.300 ;
        RECT 128.140 148.070 128.400 148.160 ;
        RECT 127.680 146.260 127.940 146.350 ;
        RECT 127.680 146.120 128.340 146.260 ;
        RECT 127.680 146.030 127.940 146.120 ;
        RECT 127.220 145.690 127.480 146.010 ;
        RECT 126.760 145.010 127.020 145.330 ;
        RECT 126.820 143.630 126.960 145.010 ;
        RECT 126.760 143.310 127.020 143.630 ;
        RECT 127.280 139.890 127.420 145.690 ;
        RECT 128.200 142.950 128.340 146.120 ;
        RECT 128.660 144.990 128.800 148.410 ;
        RECT 129.120 148.390 129.260 149.770 ;
        RECT 129.060 148.070 129.320 148.390 ;
        RECT 129.060 145.350 129.320 145.670 ;
        RECT 128.600 144.670 128.860 144.990 ;
        RECT 127.680 142.630 127.940 142.950 ;
        RECT 128.140 142.630 128.400 142.950 ;
        RECT 127.740 140.230 127.880 142.630 ;
        RECT 127.680 139.910 127.940 140.230 ;
        RECT 127.220 139.570 127.480 139.890 ;
        RECT 127.740 137.510 127.880 139.910 ;
        RECT 129.120 137.590 129.260 145.350 ;
        RECT 130.440 144.330 130.700 144.650 ;
        RECT 129.520 142.630 129.780 142.950 ;
        RECT 129.580 138.190 129.720 142.630 ;
        RECT 130.500 142.270 130.640 144.330 ;
        RECT 130.960 142.950 131.100 161.250 ;
        RECT 131.420 159.610 131.560 164.390 ;
        RECT 131.880 162.670 132.020 166.770 ;
        RECT 132.280 166.090 132.540 166.410 ;
        RECT 132.340 162.670 132.480 166.090 ;
        RECT 132.800 165.390 132.940 166.770 ;
        RECT 133.200 166.090 133.460 166.410 ;
        RECT 132.740 165.070 133.000 165.390 ;
        RECT 132.800 164.030 132.940 165.070 ;
        RECT 133.260 165.050 133.400 166.090 ;
        RECT 133.720 165.050 133.860 181.390 ;
        RECT 135.500 180.370 135.760 180.690 ;
        RECT 138.720 180.370 138.980 180.690 ;
        RECT 135.560 177.970 135.700 180.370 ;
        RECT 138.260 179.690 138.520 180.010 ;
        RECT 135.500 177.650 135.760 177.970 ;
        RECT 134.580 166.770 134.840 167.090 ;
        RECT 133.200 164.730 133.460 165.050 ;
        RECT 133.660 164.730 133.920 165.050 ;
        RECT 132.740 163.710 133.000 164.030 ;
        RECT 131.820 162.350 132.080 162.670 ;
        RECT 132.280 162.350 132.540 162.670 ;
        RECT 133.260 161.310 133.400 164.730 ;
        RECT 134.640 164.370 134.780 166.770 ;
        RECT 135.040 166.090 135.300 166.410 ;
        RECT 135.100 165.050 135.240 166.090 ;
        RECT 135.040 164.730 135.300 165.050 ;
        RECT 134.580 164.050 134.840 164.370 ;
        RECT 133.660 163.370 133.920 163.690 ;
        RECT 133.720 162.330 133.860 163.370 ;
        RECT 133.660 162.010 133.920 162.330 ;
        RECT 133.200 160.990 133.460 161.310 ;
        RECT 131.820 160.650 132.080 160.970 ;
        RECT 131.360 159.290 131.620 159.610 ;
        RECT 131.880 156.210 132.020 160.650 ;
        RECT 133.260 158.930 133.400 160.990 ;
        RECT 133.200 158.610 133.460 158.930 ;
        RECT 132.280 157.930 132.540 158.250 ;
        RECT 132.340 156.550 132.480 157.930 ;
        RECT 132.280 156.230 132.540 156.550 ;
        RECT 133.720 156.210 133.860 162.010 ;
        RECT 131.820 155.890 132.080 156.210 ;
        RECT 132.740 155.890 133.000 156.210 ;
        RECT 133.660 156.120 133.920 156.210 ;
        RECT 133.260 155.980 133.920 156.120 ;
        RECT 132.800 154.510 132.940 155.890 ;
        RECT 132.740 154.190 133.000 154.510 ;
        RECT 133.260 154.170 133.400 155.980 ;
        RECT 133.660 155.890 133.920 155.980 ;
        RECT 134.120 155.550 134.380 155.870 ;
        RECT 133.660 155.210 133.920 155.530 ;
        RECT 131.820 153.850 132.080 154.170 ;
        RECT 133.200 153.850 133.460 154.170 ;
        RECT 131.360 150.790 131.620 151.110 ;
        RECT 131.420 148.730 131.560 150.790 ;
        RECT 131.880 150.770 132.020 153.850 ;
        RECT 133.200 152.490 133.460 152.810 ;
        RECT 133.260 151.790 133.400 152.490 ;
        RECT 133.200 151.470 133.460 151.790 ;
        RECT 131.820 150.450 132.080 150.770 ;
        RECT 132.280 149.770 132.540 150.090 ;
        RECT 131.360 148.410 131.620 148.730 ;
        RECT 132.340 148.390 132.480 149.770 ;
        RECT 132.280 148.070 132.540 148.390 ;
        RECT 132.740 147.730 133.000 148.050 ;
        RECT 132.280 147.050 132.540 147.370 ;
        RECT 132.340 146.350 132.480 147.050 ;
        RECT 132.280 146.030 132.540 146.350 ;
        RECT 132.340 145.580 132.480 146.030 ;
        RECT 132.800 145.670 132.940 147.730 ;
        RECT 131.420 145.440 132.480 145.580 ;
        RECT 130.900 142.630 131.160 142.950 ;
        RECT 130.440 141.950 130.700 142.270 ;
        RECT 130.500 140.910 130.640 141.950 ;
        RECT 130.440 140.590 130.700 140.910 ;
        RECT 131.420 139.890 131.560 145.440 ;
        RECT 132.740 145.350 133.000 145.670 ;
        RECT 133.260 145.070 133.400 151.470 ;
        RECT 133.720 150.770 133.860 155.210 ;
        RECT 134.180 152.810 134.320 155.550 ;
        RECT 135.040 152.830 135.300 153.150 ;
        RECT 134.120 152.490 134.380 152.810 ;
        RECT 135.100 151.790 135.240 152.830 ;
        RECT 135.040 151.470 135.300 151.790 ;
        RECT 134.120 150.790 134.380 151.110 ;
        RECT 133.660 150.450 133.920 150.770 ;
        RECT 133.660 148.070 133.920 148.390 ;
        RECT 133.720 145.580 133.860 148.070 ;
        RECT 134.180 147.370 134.320 150.790 ;
        RECT 135.040 150.450 135.300 150.770 ;
        RECT 134.580 150.110 134.840 150.430 ;
        RECT 134.640 148.730 134.780 150.110 ;
        RECT 135.100 149.070 135.240 150.450 ;
        RECT 135.040 148.750 135.300 149.070 ;
        RECT 134.580 148.410 134.840 148.730 ;
        RECT 134.120 147.050 134.380 147.370 ;
        RECT 133.720 145.440 134.780 145.580 ;
        RECT 131.880 144.990 134.320 145.070 ;
        RECT 131.820 144.930 134.380 144.990 ;
        RECT 131.820 144.670 132.080 144.930 ;
        RECT 134.120 144.670 134.380 144.930 ;
        RECT 134.640 142.270 134.780 145.440 ;
        RECT 132.280 141.950 132.540 142.270 ;
        RECT 134.580 141.950 134.840 142.270 ;
        RECT 131.360 139.570 131.620 139.890 ;
        RECT 129.980 139.230 130.240 139.550 ;
        RECT 130.040 138.190 130.180 139.230 ;
        RECT 131.820 138.890 132.080 139.210 ;
        RECT 129.520 137.870 129.780 138.190 ;
        RECT 129.980 137.870 130.240 138.190 ;
        RECT 127.680 137.190 127.940 137.510 ;
        RECT 129.120 137.450 129.720 137.590 ;
        RECT 131.880 137.510 132.020 138.890 ;
        RECT 127.220 136.850 127.480 137.170 ;
        RECT 127.280 134.790 127.420 136.850 ;
        RECT 128.140 136.510 128.400 136.830 ;
        RECT 128.200 134.790 128.340 136.510 ;
        RECT 127.220 134.470 127.480 134.790 ;
        RECT 128.140 134.470 128.400 134.790 ;
        RECT 128.600 134.130 128.860 134.450 ;
        RECT 129.060 134.130 129.320 134.450 ;
        RECT 128.660 132.945 128.800 134.130 ;
        RECT 128.590 132.575 128.870 132.945 ;
        RECT 128.660 131.730 128.800 132.575 ;
        RECT 129.120 132.410 129.260 134.130 ;
        RECT 129.060 132.090 129.320 132.410 ;
        RECT 128.600 131.410 128.860 131.730 ;
        RECT 129.120 130.030 129.260 132.090 ;
        RECT 129.060 129.710 129.320 130.030 ;
        RECT 129.580 129.350 129.720 137.450 ;
        RECT 131.360 137.190 131.620 137.510 ;
        RECT 131.820 137.190 132.080 137.510 ;
        RECT 131.420 134.110 131.560 137.190 ;
        RECT 131.880 135.470 132.020 137.190 ;
        RECT 131.820 135.150 132.080 135.470 ;
        RECT 131.360 133.790 131.620 134.110 ;
        RECT 129.980 132.430 130.240 132.750 ;
        RECT 130.430 132.575 130.710 132.945 ;
        RECT 130.040 131.050 130.180 132.430 ;
        RECT 130.500 132.410 130.640 132.575 ;
        RECT 130.440 132.090 130.700 132.410 ;
        RECT 132.340 132.070 132.480 141.950 ;
        RECT 134.580 139.570 134.840 139.890 ;
        RECT 134.640 137.850 134.780 139.570 ;
        RECT 134.580 137.530 134.840 137.850 ;
        RECT 134.120 137.190 134.380 137.510 ;
        RECT 133.200 136.850 133.460 137.170 ;
        RECT 133.260 134.110 133.400 136.850 ;
        RECT 133.200 133.790 133.460 134.110 ;
        RECT 133.260 132.750 133.400 133.790 ;
        RECT 133.200 132.430 133.460 132.750 ;
        RECT 133.660 132.150 133.920 132.410 ;
        RECT 133.260 132.090 133.920 132.150 ;
        RECT 132.280 131.750 132.540 132.070 ;
        RECT 133.260 132.010 133.860 132.090 ;
        RECT 129.980 130.730 130.240 131.050 ;
        RECT 129.520 129.030 129.780 129.350 ;
        RECT 125.380 126.310 125.640 126.630 ;
        RECT 126.300 126.310 126.560 126.630 ;
        RECT 123.540 125.290 123.800 125.610 ;
        RECT 123.600 123.910 123.740 125.290 ;
        RECT 125.440 124.250 125.580 126.310 ;
        RECT 128.600 125.970 128.860 126.290 ;
        RECT 128.660 124.590 128.800 125.970 ;
        RECT 126.760 124.270 127.020 124.590 ;
        RECT 128.600 124.270 128.860 124.590 ;
        RECT 124.920 123.930 125.180 124.250 ;
        RECT 125.380 123.930 125.640 124.250 ;
        RECT 123.540 123.590 123.800 123.910 ;
        RECT 121.700 123.250 121.960 123.570 ;
        RECT 121.760 119.150 121.900 123.250 ;
        RECT 122.670 122.035 124.210 122.405 ;
        RECT 124.980 121.190 125.120 123.930 ;
        RECT 126.300 122.910 126.560 123.230 ;
        RECT 126.360 121.870 126.500 122.910 ;
        RECT 126.300 121.550 126.560 121.870 ;
        RECT 124.920 120.870 125.180 121.190 ;
        RECT 123.540 120.530 123.800 120.850 ;
        RECT 121.700 118.830 121.960 119.150 ;
        RECT 123.600 118.470 123.740 120.530 ;
        RECT 123.540 118.150 123.800 118.470 ;
        RECT 120.320 117.130 120.580 117.450 ;
        RECT 118.480 115.770 118.740 116.090 ;
        RECT 120.380 115.410 120.520 117.130 ;
        RECT 122.670 116.595 124.210 116.965 ;
        RECT 118.480 115.090 118.740 115.410 ;
        RECT 120.320 115.090 120.580 115.410 ;
        RECT 115.720 114.410 115.980 114.730 ;
        RECT 115.780 113.710 115.920 114.410 ;
        RECT 115.720 113.390 115.980 113.710 ;
        RECT 118.540 112.690 118.680 115.090 ;
        RECT 124.920 113.050 125.180 113.370 ;
        RECT 115.260 112.370 115.520 112.690 ;
        RECT 118.480 112.370 118.740 112.690 ;
        RECT 119.860 112.370 120.120 112.690 ;
        RECT 114.340 111.690 114.600 112.010 ;
        RECT 118.020 111.690 118.280 112.010 ;
        RECT 112.040 109.650 112.300 109.970 ;
        RECT 112.100 107.250 112.240 109.650 ;
        RECT 114.400 108.270 114.540 111.690 ;
        RECT 118.080 110.650 118.220 111.690 ;
        RECT 119.920 110.990 120.060 112.370 ;
        RECT 121.700 111.690 121.960 112.010 ;
        RECT 124.460 111.690 124.720 112.010 ;
        RECT 119.860 110.670 120.120 110.990 ;
        RECT 118.020 110.330 118.280 110.650 ;
        RECT 120.320 109.990 120.580 110.310 ;
        RECT 120.380 108.270 120.520 109.990 ;
        RECT 114.340 107.950 114.600 108.270 ;
        RECT 120.320 107.950 120.580 108.270 ;
        RECT 112.040 106.930 112.300 107.250 ;
        RECT 111.580 105.230 111.840 105.550 ;
        RECT 112.100 105.210 112.240 106.930 ;
        RECT 112.500 106.590 112.760 106.910 ;
        RECT 112.040 104.890 112.300 105.210 ;
        RECT 110.660 104.550 110.920 104.870 ;
        RECT 108.820 104.210 109.080 104.530 ;
        RECT 101.920 103.870 102.180 104.190 ;
        RECT 101.460 101.830 101.720 102.150 ;
        RECT 101.980 101.810 102.120 103.870 ;
        RECT 105.140 103.530 105.400 103.850 ;
        RECT 99.620 101.720 99.880 101.810 ;
        RECT 99.220 101.580 99.880 101.720 ;
        RECT 98.700 100.810 98.960 101.130 ;
        RECT 98.240 99.340 98.500 99.430 ;
        RECT 97.840 99.200 98.500 99.340 ;
        RECT 98.240 99.110 98.500 99.200 ;
        RECT 98.760 99.090 98.900 100.810 ;
        RECT 99.220 99.430 99.360 101.580 ;
        RECT 99.620 101.490 99.880 101.580 ;
        RECT 101.920 101.490 102.180 101.810 ;
        RECT 104.680 101.150 104.940 101.470 ;
        RECT 99.620 100.810 99.880 101.130 ;
        RECT 99.680 99.430 99.820 100.810 ;
        RECT 101.460 99.450 101.720 99.770 ;
        RECT 99.160 99.110 99.420 99.430 ;
        RECT 99.620 99.110 99.880 99.430 ;
        RECT 98.700 98.770 98.960 99.090 ;
        RECT 95.480 96.730 95.740 97.050 ;
        RECT 95.540 93.990 95.680 96.730 ;
        RECT 96.400 96.050 96.660 96.370 ;
        RECT 96.860 96.225 97.120 96.370 ;
        RECT 96.460 93.990 96.600 96.050 ;
        RECT 96.850 95.855 97.130 96.225 ;
        RECT 97.780 96.050 98.040 96.370 ;
        RECT 97.840 94.580 97.980 96.050 ;
        RECT 97.380 94.440 97.980 94.580 ;
        RECT 95.480 93.670 95.740 93.990 ;
        RECT 96.400 93.670 96.660 93.990 ;
        RECT 95.020 90.840 95.280 90.930 ;
        RECT 95.540 90.840 95.680 93.670 ;
        RECT 95.020 90.700 95.680 90.840 ;
        RECT 95.940 90.840 96.200 90.930 ;
        RECT 96.460 90.840 96.600 93.670 ;
        RECT 97.380 93.310 97.520 94.440 ;
        RECT 97.780 93.670 98.040 93.990 ;
        RECT 98.240 93.670 98.500 93.990 ;
        RECT 97.320 92.990 97.580 93.310 ;
        RECT 97.840 90.930 97.980 93.670 ;
        RECT 98.300 91.950 98.440 93.670 ;
        RECT 101.520 91.950 101.660 99.450 ;
        RECT 103.760 98.770 104.020 99.090 ;
        RECT 102.380 96.050 102.640 96.370 ;
        RECT 101.920 95.370 102.180 95.690 ;
        RECT 101.980 93.990 102.120 95.370 ;
        RECT 101.920 93.670 102.180 93.990 ;
        RECT 102.440 91.950 102.580 96.050 ;
        RECT 98.240 91.630 98.500 91.950 ;
        RECT 101.460 91.630 101.720 91.950 ;
        RECT 102.380 91.630 102.640 91.950 ;
        RECT 95.940 90.700 96.600 90.840 ;
        RECT 95.020 90.610 95.280 90.700 ;
        RECT 95.940 90.610 96.200 90.700 ;
        RECT 97.780 90.610 98.040 90.930 ;
        RECT 101.000 89.930 101.260 90.250 ;
        RECT 101.060 89.230 101.200 89.930 ;
        RECT 101.000 88.910 101.260 89.230 ;
        RECT 101.520 86.510 101.660 91.630 ;
        RECT 103.300 90.270 103.560 90.590 ;
        RECT 103.360 88.550 103.500 90.270 ;
        RECT 103.300 88.230 103.560 88.550 ;
        RECT 101.460 86.190 101.720 86.510 ;
        RECT 98.700 85.850 98.960 86.170 ;
        RECT 96.400 84.830 96.660 85.150 ;
        RECT 97.320 84.830 97.580 85.150 ;
        RECT 95.940 84.490 96.200 84.810 ;
        RECT 96.000 81.070 96.140 84.490 ;
        RECT 95.940 80.750 96.200 81.070 ;
        RECT 96.460 80.470 96.600 84.830 ;
        RECT 97.380 83.790 97.520 84.830 ;
        RECT 97.780 84.490 98.040 84.810 ;
        RECT 97.320 83.470 97.580 83.790 ;
        RECT 97.840 83.450 97.980 84.490 ;
        RECT 97.780 83.130 98.040 83.450 ;
        RECT 97.320 82.790 97.580 83.110 ;
        RECT 97.380 81.070 97.520 82.790 ;
        RECT 97.320 80.750 97.580 81.070 ;
        RECT 96.000 80.330 96.600 80.470 ;
        RECT 97.840 80.390 97.980 83.130 ;
        RECT 98.760 82.770 98.900 85.850 ;
        RECT 102.840 85.170 103.100 85.490 ;
        RECT 100.080 84.490 100.340 84.810 ;
        RECT 102.380 84.490 102.640 84.810 ;
        RECT 100.140 83.110 100.280 84.490 ;
        RECT 102.440 83.790 102.580 84.490 ;
        RECT 102.380 83.470 102.640 83.790 ;
        RECT 100.080 82.790 100.340 83.110 ;
        RECT 98.700 82.450 98.960 82.770 ;
        RECT 98.760 81.070 98.900 82.450 ;
        RECT 102.900 82.090 103.040 85.170 ;
        RECT 101.460 81.770 101.720 82.090 ;
        RECT 102.840 81.770 103.100 82.090 ;
        RECT 98.700 80.750 98.960 81.070 ;
        RECT 96.000 79.370 96.140 80.330 ;
        RECT 97.780 80.070 98.040 80.390 ;
        RECT 101.520 80.050 101.660 81.770 ;
        RECT 101.460 79.730 101.720 80.050 ;
        RECT 95.940 79.050 96.200 79.370 ;
        RECT 101.460 76.330 101.720 76.650 ;
        RECT 101.520 74.950 101.660 76.330 ;
        RECT 101.460 74.630 101.720 74.950 ;
        RECT 103.820 74.610 103.960 98.770 ;
        RECT 104.220 98.090 104.480 98.410 ;
        RECT 97.320 74.290 97.580 74.610 ;
        RECT 99.620 74.290 99.880 74.610 ;
        RECT 102.380 74.290 102.640 74.610 ;
        RECT 103.760 74.290 104.020 74.610 ;
        RECT 95.940 73.670 96.200 73.930 ;
        RECT 94.620 73.610 96.200 73.670 ;
        RECT 94.620 73.530 96.140 73.610 ;
        RECT 97.380 72.910 97.520 74.290 ;
        RECT 99.680 72.910 99.820 74.290 ;
        RECT 101.460 73.610 101.720 73.930 ;
        RECT 97.320 72.590 97.580 72.910 ;
        RECT 99.620 72.590 99.880 72.910 ;
        RECT 95.480 72.250 95.740 72.570 ;
        RECT 94.100 69.870 94.360 70.190 ;
        RECT 93.640 69.530 93.900 69.850 ;
        RECT 91.340 68.850 91.600 69.170 ;
        RECT 92.260 68.850 92.520 69.170 ;
        RECT 90.880 68.170 91.140 68.490 ;
        RECT 89.090 67.635 90.630 68.005 ;
        RECT 90.940 64.150 91.080 68.170 ;
        RECT 91.400 66.790 91.540 68.850 ;
        RECT 91.340 66.470 91.600 66.790 ;
        RECT 90.940 64.010 91.540 64.150 ;
        RECT 92.320 64.070 92.460 68.850 ;
        RECT 90.880 63.410 91.140 63.730 ;
        RECT 89.090 62.195 90.630 62.565 ;
        RECT 87.660 61.030 87.920 61.350 ;
        RECT 88.580 61.030 88.840 61.350 ;
        RECT 86.740 60.690 87.000 61.010 ;
        RECT 86.800 59.310 86.940 60.690 ;
        RECT 88.580 60.010 88.840 60.330 ;
        RECT 86.740 58.990 87.000 59.310 ;
        RECT 85.820 57.970 86.080 58.290 ;
        RECT 86.740 57.970 87.000 58.290 ;
        RECT 86.800 56.220 86.940 57.970 ;
        RECT 88.640 56.500 88.780 60.010 ;
        RECT 90.940 58.290 91.080 63.410 ;
        RECT 91.400 58.290 91.540 64.010 ;
        RECT 92.260 63.750 92.520 64.070 ;
        RECT 92.720 63.410 92.980 63.730 ;
        RECT 92.780 61.350 92.920 63.410 ;
        RECT 94.160 61.350 94.300 69.870 ;
        RECT 95.540 69.025 95.680 72.250 ;
        RECT 101.520 72.230 101.660 73.610 ;
        RECT 102.440 72.910 102.580 74.290 ;
        RECT 102.380 72.590 102.640 72.910 ;
        RECT 96.860 71.910 97.120 72.230 ;
        RECT 101.460 71.910 101.720 72.230 ;
        RECT 96.920 70.190 97.060 71.910 ;
        RECT 101.460 71.230 101.720 71.550 ;
        RECT 97.320 70.890 97.580 71.210 ;
        RECT 96.860 69.870 97.120 70.190 ;
        RECT 97.380 69.850 97.520 70.890 ;
        RECT 96.850 69.335 97.130 69.705 ;
        RECT 97.320 69.530 97.580 69.850 ;
        RECT 96.860 69.190 97.120 69.335 ;
        RECT 95.470 68.655 95.750 69.025 ;
        RECT 99.620 68.850 99.880 69.170 ;
        RECT 95.480 68.510 95.740 68.655 ;
        RECT 99.680 67.470 99.820 68.850 ;
        RECT 100.540 68.170 100.800 68.490 ;
        RECT 99.620 67.150 99.880 67.470 ;
        RECT 100.600 66.790 100.740 68.170 ;
        RECT 101.520 66.790 101.660 71.230 ;
        RECT 101.920 70.890 102.180 71.210 ;
        RECT 101.980 69.510 102.120 70.890 ;
        RECT 101.920 69.190 102.180 69.510 ;
        RECT 104.280 69.170 104.420 98.090 ;
        RECT 104.740 96.710 104.880 101.150 ;
        RECT 105.200 99.090 105.340 103.530 ;
        RECT 105.880 102.995 107.420 103.365 ;
        RECT 110.720 99.625 110.860 104.550 ;
        RECT 112.560 104.530 112.700 106.590 ;
        RECT 114.400 105.550 114.540 107.950 ;
        RECT 119.400 106.590 119.660 106.910 ;
        RECT 114.340 105.230 114.600 105.550 ;
        RECT 112.500 104.210 112.760 104.530 ;
        RECT 111.120 102.510 111.380 102.830 ;
        RECT 107.900 99.110 108.160 99.430 ;
        RECT 110.650 99.255 110.930 99.625 ;
        RECT 105.140 98.770 105.400 99.090 ;
        RECT 104.680 96.390 104.940 96.710 ;
        RECT 105.200 94.330 105.340 98.770 ;
        RECT 105.880 97.555 107.420 97.925 ;
        RECT 107.960 97.390 108.100 99.110 ;
        RECT 107.900 97.070 108.160 97.390 ;
        RECT 109.740 96.960 110.000 97.050 ;
        RECT 109.340 96.820 110.000 96.960 ;
        RECT 105.140 94.010 105.400 94.330 ;
        RECT 108.360 93.330 108.620 93.650 ;
        RECT 105.880 92.115 107.420 92.485 ;
        RECT 104.680 90.610 104.940 90.930 ;
        RECT 105.140 90.610 105.400 90.930 ;
        RECT 105.600 90.610 105.860 90.930 ;
        RECT 104.740 88.550 104.880 90.610 ;
        RECT 105.200 88.550 105.340 90.610 ;
        RECT 104.680 88.230 104.940 88.550 ;
        RECT 105.140 88.230 105.400 88.550 ;
        RECT 105.200 85.490 105.340 88.230 ;
        RECT 105.660 88.210 105.800 90.610 ;
        RECT 108.420 88.890 108.560 93.330 ;
        RECT 108.820 92.650 109.080 92.970 ;
        RECT 108.880 90.590 109.020 92.650 ;
        RECT 109.340 91.610 109.480 96.820 ;
        RECT 109.740 96.730 110.000 96.820 ;
        RECT 110.660 92.990 110.920 93.310 ;
        RECT 109.280 91.290 109.540 91.610 ;
        RECT 109.740 91.290 110.000 91.610 ;
        RECT 108.820 90.270 109.080 90.590 ;
        RECT 108.360 88.570 108.620 88.890 ;
        RECT 108.880 88.550 109.020 90.270 ;
        RECT 109.800 88.550 109.940 91.290 ;
        RECT 110.720 90.930 110.860 92.990 ;
        RECT 111.180 91.350 111.320 102.510 ;
        RECT 113.420 101.490 113.680 101.810 ;
        RECT 117.560 101.490 117.820 101.810 ;
        RECT 113.480 99.770 113.620 101.490 ;
        RECT 113.880 100.810 114.140 101.130 ;
        RECT 113.420 99.450 113.680 99.770 ;
        RECT 113.480 97.390 113.620 99.450 ;
        RECT 113.420 97.070 113.680 97.390 ;
        RECT 113.420 96.050 113.680 96.370 ;
        RECT 111.580 95.710 111.840 96.030 ;
        RECT 111.640 94.670 111.780 95.710 ;
        RECT 111.580 94.350 111.840 94.670 ;
        RECT 112.040 92.650 112.300 92.970 ;
        RECT 112.100 91.950 112.240 92.650 ;
        RECT 112.040 91.630 112.300 91.950 ;
        RECT 111.180 91.210 111.780 91.350 ;
        RECT 110.660 90.610 110.920 90.930 ;
        RECT 111.120 90.610 111.380 90.930 ;
        RECT 111.180 90.160 111.320 90.610 ;
        RECT 110.260 90.020 111.320 90.160 ;
        RECT 108.820 88.230 109.080 88.550 ;
        RECT 109.740 88.230 110.000 88.550 ;
        RECT 110.260 88.210 110.400 90.020 ;
        RECT 105.600 87.890 105.860 88.210 ;
        RECT 108.360 87.890 108.620 88.210 ;
        RECT 110.200 87.890 110.460 88.210 ;
        RECT 110.660 87.890 110.920 88.210 ;
        RECT 107.900 87.550 108.160 87.870 ;
        RECT 105.880 86.675 107.420 87.045 ;
        RECT 105.140 85.170 105.400 85.490 ;
        RECT 105.600 85.170 105.860 85.490 ;
        RECT 105.660 84.720 105.800 85.170 ;
        RECT 107.960 84.810 108.100 87.550 ;
        RECT 105.200 84.580 105.800 84.720 ;
        RECT 105.200 73.930 105.340 84.580 ;
        RECT 106.060 84.490 106.320 84.810 ;
        RECT 107.900 84.490 108.160 84.810 ;
        RECT 106.120 83.450 106.260 84.490 ;
        RECT 106.060 83.130 106.320 83.450 ;
        RECT 105.880 81.235 107.420 81.605 ;
        RECT 105.880 75.795 107.420 76.165 ;
        RECT 106.980 73.950 107.240 74.270 ;
        RECT 105.140 73.610 105.400 73.930 ;
        RECT 107.040 72.910 107.180 73.950 ;
        RECT 106.980 72.590 107.240 72.910 ;
        RECT 105.140 72.250 105.400 72.570 ;
        RECT 104.220 68.850 104.480 69.170 ;
        RECT 97.320 66.470 97.580 66.790 ;
        RECT 100.540 66.470 100.800 66.790 ;
        RECT 101.460 66.470 101.720 66.790 ;
        RECT 95.940 65.450 96.200 65.770 ;
        RECT 96.000 64.070 96.140 65.450 ;
        RECT 95.940 63.750 96.200 64.070 ;
        RECT 97.380 63.730 97.520 66.470 ;
        RECT 101.460 65.450 101.720 65.770 ;
        RECT 102.840 65.450 103.100 65.770 ;
        RECT 97.320 63.410 97.580 63.730 ;
        RECT 100.540 63.410 100.800 63.730 ;
        RECT 92.260 61.030 92.520 61.350 ;
        RECT 92.720 61.030 92.980 61.350 ;
        RECT 94.100 61.030 94.360 61.350 ;
        RECT 97.780 61.030 98.040 61.350 ;
        RECT 90.880 57.970 91.140 58.290 ;
        RECT 91.340 57.970 91.600 58.290 ;
        RECT 89.090 56.755 90.630 57.125 ;
        RECT 88.640 56.360 89.700 56.500 ;
        RECT 89.560 56.220 89.700 56.360 ;
        RECT 92.320 56.220 92.460 61.030 ;
        RECT 95.020 57.970 95.280 58.290 ;
        RECT 95.080 56.220 95.220 57.970 ;
        RECT 97.840 56.220 97.980 61.030 ;
        RECT 100.600 56.220 100.740 63.410 ;
        RECT 101.520 61.350 101.660 65.450 ;
        RECT 101.920 63.410 102.180 63.730 ;
        RECT 101.460 61.030 101.720 61.350 ;
        RECT 101.980 58.290 102.120 63.410 ;
        RECT 102.900 58.290 103.040 65.450 ;
        RECT 105.200 61.690 105.340 72.250 ;
        RECT 105.880 70.355 107.420 70.725 ;
        RECT 108.420 69.850 108.560 87.890 ;
        RECT 109.280 85.170 109.540 85.490 ;
        RECT 108.820 84.830 109.080 85.150 ;
        RECT 108.880 83.450 109.020 84.830 ;
        RECT 109.340 83.450 109.480 85.170 ;
        RECT 108.820 83.130 109.080 83.450 ;
        RECT 109.280 83.130 109.540 83.450 ;
        RECT 109.340 80.730 109.480 83.130 ;
        RECT 109.740 82.110 110.000 82.430 ;
        RECT 109.280 80.410 109.540 80.730 ;
        RECT 109.800 77.670 109.940 82.110 ;
        RECT 110.720 81.070 110.860 87.890 ;
        RECT 110.660 80.750 110.920 81.070 ;
        RECT 111.640 80.390 111.780 91.210 ;
        RECT 112.040 88.230 112.300 88.550 ;
        RECT 112.100 87.530 112.240 88.230 ;
        RECT 112.040 87.210 112.300 87.530 ;
        RECT 111.580 80.070 111.840 80.390 ;
        RECT 110.660 79.730 110.920 80.050 ;
        RECT 110.200 79.050 110.460 79.370 ;
        RECT 110.260 77.670 110.400 79.050 ;
        RECT 109.740 77.350 110.000 77.670 ;
        RECT 110.200 77.350 110.460 77.670 ;
        RECT 109.280 73.610 109.540 73.930 ;
        RECT 109.340 72.570 109.480 73.610 ;
        RECT 109.280 72.250 109.540 72.570 ;
        RECT 110.720 71.890 110.860 79.730 ;
        RECT 111.640 74.950 111.780 80.070 ;
        RECT 113.480 78.350 113.620 96.050 ;
        RECT 113.940 93.650 114.080 100.810 ;
        RECT 115.260 98.770 115.520 99.090 ;
        RECT 116.180 98.770 116.440 99.090 ;
        RECT 117.100 98.770 117.360 99.090 ;
        RECT 114.340 98.090 114.600 98.410 ;
        RECT 114.400 96.370 114.540 98.090 ;
        RECT 115.320 96.370 115.460 98.770 ;
        RECT 116.240 97.050 116.380 98.770 ;
        RECT 116.180 96.730 116.440 97.050 ;
        RECT 117.160 96.710 117.300 98.770 ;
        RECT 117.620 97.390 117.760 101.490 ;
        RECT 118.020 100.810 118.280 101.130 ;
        RECT 118.080 99.770 118.220 100.810 ;
        RECT 118.020 99.450 118.280 99.770 ;
        RECT 117.560 97.070 117.820 97.390 ;
        RECT 117.100 96.390 117.360 96.710 ;
        RECT 118.080 96.370 118.220 99.450 ;
        RECT 119.460 99.090 119.600 106.590 ;
        RECT 120.380 104.870 120.520 107.950 ;
        RECT 121.760 107.250 121.900 111.690 ;
        RECT 122.670 111.155 124.210 111.525 ;
        RECT 122.160 110.670 122.420 110.990 ;
        RECT 122.220 109.290 122.360 110.670 ;
        RECT 124.000 110.560 124.260 110.650 ;
        RECT 124.520 110.560 124.660 111.690 ;
        RECT 124.000 110.420 124.660 110.560 ;
        RECT 124.000 110.330 124.260 110.420 ;
        RECT 122.160 108.970 122.420 109.290 ;
        RECT 122.220 107.930 122.360 108.970 ;
        RECT 122.160 107.610 122.420 107.930 ;
        RECT 124.980 107.250 125.120 113.050 ;
        RECT 125.380 112.710 125.640 113.030 ;
        RECT 125.440 108.270 125.580 112.710 ;
        RECT 125.380 107.950 125.640 108.270 ;
        RECT 121.700 106.930 121.960 107.250 ;
        RECT 124.920 106.930 125.180 107.250 ;
        RECT 122.670 105.715 124.210 106.085 ;
        RECT 120.320 104.550 120.580 104.870 ;
        RECT 124.920 101.490 125.180 101.810 ;
        RECT 119.860 101.150 120.120 101.470 ;
        RECT 119.920 100.110 120.060 101.150 ;
        RECT 122.670 100.275 124.210 100.645 ;
        RECT 119.860 99.790 120.120 100.110 ;
        RECT 124.980 99.770 125.120 101.490 ;
        RECT 126.820 101.130 126.960 124.270 ;
        RECT 129.580 123.570 129.720 129.030 ;
        RECT 130.440 128.690 130.700 129.010 ;
        RECT 130.500 126.970 130.640 128.690 ;
        RECT 130.440 126.650 130.700 126.970 ;
        RECT 129.980 125.630 130.240 125.950 ;
        RECT 129.520 123.250 129.780 123.570 ;
        RECT 127.220 120.870 127.480 121.190 ;
        RECT 127.680 120.870 127.940 121.190 ;
        RECT 127.280 118.130 127.420 120.870 ;
        RECT 127.220 117.810 127.480 118.130 ;
        RECT 127.740 110.650 127.880 120.870 ;
        RECT 129.060 117.810 129.320 118.130 ;
        RECT 128.140 115.430 128.400 115.750 ;
        RECT 127.680 110.330 127.940 110.650 ;
        RECT 127.740 105.210 127.880 110.330 ;
        RECT 128.200 109.290 128.340 115.430 ;
        RECT 129.120 113.710 129.260 117.810 ;
        RECT 130.040 116.390 130.180 125.630 ;
        RECT 130.500 124.590 130.640 126.650 ;
        RECT 130.440 124.270 130.700 124.590 ;
        RECT 130.500 120.850 130.640 124.270 ;
        RECT 130.900 122.910 131.160 123.230 ;
        RECT 130.960 121.870 131.100 122.910 ;
        RECT 130.900 121.550 131.160 121.870 ;
        RECT 132.340 121.190 132.480 131.750 ;
        RECT 132.740 130.730 133.000 131.050 ;
        RECT 132.800 128.670 132.940 130.730 ;
        RECT 132.740 128.350 133.000 128.670 ;
        RECT 133.260 126.630 133.400 132.010 ;
        RECT 134.180 129.010 134.320 137.190 ;
        RECT 134.640 131.390 134.780 137.530 ;
        RECT 135.040 137.190 135.300 137.510 ;
        RECT 135.100 135.470 135.240 137.190 ;
        RECT 135.040 135.150 135.300 135.470 ;
        RECT 134.580 131.070 134.840 131.390 ;
        RECT 134.120 128.690 134.380 129.010 ;
        RECT 135.040 126.650 135.300 126.970 ;
        RECT 133.200 126.310 133.460 126.630 ;
        RECT 132.280 120.870 132.540 121.190 ;
        RECT 130.440 120.530 130.700 120.850 ;
        RECT 133.260 118.470 133.400 126.310 ;
        RECT 133.660 121.210 133.920 121.530 ;
        RECT 133.200 118.150 133.460 118.470 ;
        RECT 133.720 117.790 133.860 121.210 ;
        RECT 135.100 120.510 135.240 126.650 ;
        RECT 135.040 120.190 135.300 120.510 ;
        RECT 135.100 119.150 135.240 120.190 ;
        RECT 134.120 118.830 134.380 119.150 ;
        RECT 135.040 118.830 135.300 119.150 ;
        RECT 133.660 117.470 133.920 117.790 ;
        RECT 133.200 117.130 133.460 117.450 ;
        RECT 133.260 116.430 133.400 117.130 ;
        RECT 129.580 116.250 130.180 116.390 ;
        RECT 129.060 113.390 129.320 113.710 ;
        RECT 128.600 112.370 128.860 112.690 ;
        RECT 128.660 110.990 128.800 112.370 ;
        RECT 128.600 110.670 128.860 110.990 ;
        RECT 128.140 108.970 128.400 109.290 ;
        RECT 127.680 104.890 127.940 105.210 ;
        RECT 129.580 101.470 129.720 116.250 ;
        RECT 133.200 116.110 133.460 116.430 ;
        RECT 132.280 115.430 132.540 115.750 ;
        RECT 130.440 115.090 130.700 115.410 ;
        RECT 130.500 113.030 130.640 115.090 ;
        RECT 130.440 112.710 130.700 113.030 ;
        RECT 129.980 112.030 130.240 112.350 ;
        RECT 130.040 110.990 130.180 112.030 ;
        RECT 129.980 110.670 130.240 110.990 ;
        RECT 129.980 109.990 130.240 110.310 ;
        RECT 130.040 107.250 130.180 109.990 ;
        RECT 130.500 107.590 130.640 112.710 ;
        RECT 131.360 112.370 131.620 112.690 ;
        RECT 131.820 112.370 132.080 112.690 ;
        RECT 130.900 108.970 131.160 109.290 ;
        RECT 130.440 107.270 130.700 107.590 ;
        RECT 129.980 106.930 130.240 107.250 ;
        RECT 129.520 101.150 129.780 101.470 ;
        RECT 126.760 100.810 127.020 101.130 ;
        RECT 124.920 99.450 125.180 99.770 ;
        RECT 126.300 99.450 126.560 99.770 ;
        RECT 120.780 99.110 121.040 99.430 ;
        RECT 122.160 99.110 122.420 99.430 ;
        RECT 119.400 98.770 119.660 99.090 ;
        RECT 120.320 98.770 120.580 99.090 ;
        RECT 119.400 98.090 119.660 98.410 ;
        RECT 119.460 96.370 119.600 98.090 ;
        RECT 120.380 96.370 120.520 98.770 ;
        RECT 120.840 96.710 120.980 99.110 ;
        RECT 122.220 97.390 122.360 99.110 ;
        RECT 124.000 98.430 124.260 98.750 ;
        RECT 122.160 97.070 122.420 97.390 ;
        RECT 120.780 96.390 121.040 96.710 ;
        RECT 114.340 96.050 114.600 96.370 ;
        RECT 115.260 96.050 115.520 96.370 ;
        RECT 118.020 96.050 118.280 96.370 ;
        RECT 119.400 96.050 119.660 96.370 ;
        RECT 120.320 96.050 120.580 96.370 ;
        RECT 118.020 93.670 118.280 93.990 ;
        RECT 113.880 93.330 114.140 93.650 ;
        RECT 113.940 91.270 114.080 93.330 ;
        RECT 117.560 92.990 117.820 93.310 ;
        RECT 114.340 92.650 114.600 92.970 ;
        RECT 114.400 91.950 114.540 92.650 ;
        RECT 117.620 91.950 117.760 92.990 ;
        RECT 114.340 91.630 114.600 91.950 ;
        RECT 117.560 91.630 117.820 91.950 ;
        RECT 113.880 90.950 114.140 91.270 ;
        RECT 115.260 90.270 115.520 90.590 ;
        RECT 115.320 89.230 115.460 90.270 ;
        RECT 117.620 90.250 117.760 91.630 ;
        RECT 118.080 91.610 118.220 93.670 ;
        RECT 118.480 93.330 118.740 93.650 ;
        RECT 118.020 91.290 118.280 91.610 ;
        RECT 117.560 89.930 117.820 90.250 ;
        RECT 118.080 89.230 118.220 91.290 ;
        RECT 118.540 90.930 118.680 93.330 ;
        RECT 118.480 90.610 118.740 90.930 ;
        RECT 118.540 89.230 118.680 90.610 ;
        RECT 115.260 88.910 115.520 89.230 ;
        RECT 118.020 88.910 118.280 89.230 ;
        RECT 118.480 88.910 118.740 89.230 ;
        RECT 118.480 82.450 118.740 82.770 ;
        RECT 114.340 81.770 114.600 82.090 ;
        RECT 116.640 81.770 116.900 82.090 ;
        RECT 114.400 80.390 114.540 81.770 ;
        RECT 114.340 80.070 114.600 80.390 ;
        RECT 115.720 79.730 115.980 80.050 ;
        RECT 115.780 78.350 115.920 79.730 ;
        RECT 113.420 78.030 113.680 78.350 ;
        RECT 115.720 78.030 115.980 78.350 ;
        RECT 116.700 78.010 116.840 81.770 ;
        RECT 118.540 80.730 118.680 82.450 ;
        RECT 118.480 80.410 118.740 80.730 ;
        RECT 119.460 79.370 119.600 96.050 ;
        RECT 120.380 93.990 120.520 96.050 ;
        RECT 120.840 94.070 120.980 96.390 ;
        RECT 124.060 96.370 124.200 98.430 ;
        RECT 124.000 96.280 124.260 96.370 ;
        RECT 124.000 96.140 124.660 96.280 ;
        RECT 124.000 96.050 124.260 96.140 ;
        RECT 122.670 94.835 124.210 95.205 ;
        RECT 124.520 94.670 124.660 96.140 ;
        RECT 124.460 94.350 124.720 94.670 ;
        RECT 120.840 93.990 121.440 94.070 ;
        RECT 120.320 93.670 120.580 93.990 ;
        RECT 120.840 93.930 121.500 93.990 ;
        RECT 121.240 93.670 121.500 93.930 ;
        RECT 124.460 93.670 124.720 93.990 ;
        RECT 119.860 93.330 120.120 93.650 ;
        RECT 119.920 90.930 120.060 93.330 ;
        RECT 120.380 90.930 120.520 93.670 ;
        RECT 124.520 93.310 124.660 93.670 ;
        RECT 126.360 93.650 126.500 99.450 ;
        RECT 126.820 99.430 126.960 100.810 ;
        RECT 126.760 99.110 127.020 99.430 ;
        RECT 129.060 99.110 129.320 99.430 ;
        RECT 128.140 96.050 128.400 96.370 ;
        RECT 128.600 96.050 128.860 96.370 ;
        RECT 126.760 95.370 127.020 95.690 ;
        RECT 127.680 95.370 127.940 95.690 ;
        RECT 126.820 93.990 126.960 95.370 ;
        RECT 127.740 93.990 127.880 95.370 ;
        RECT 126.760 93.670 127.020 93.990 ;
        RECT 127.680 93.670 127.940 93.990 ;
        RECT 126.300 93.330 126.560 93.650 ;
        RECT 124.460 92.990 124.720 93.310 ;
        RECT 124.520 91.950 124.660 92.990 ;
        RECT 124.460 91.630 124.720 91.950 ;
        RECT 119.860 90.610 120.120 90.930 ;
        RECT 120.320 90.610 120.580 90.930 ;
        RECT 125.840 90.270 126.100 90.590 ;
        RECT 122.670 89.395 124.210 89.765 ;
        RECT 125.900 88.890 126.040 90.270 ;
        RECT 125.840 88.570 126.100 88.890 ;
        RECT 121.240 88.230 121.500 88.550 ;
        RECT 119.860 82.790 120.120 83.110 ;
        RECT 119.400 79.050 119.660 79.370 ;
        RECT 116.640 77.690 116.900 78.010 ;
        RECT 114.800 77.350 115.060 77.670 ;
        RECT 114.860 75.630 115.000 77.350 ;
        RECT 114.800 75.310 115.060 75.630 ;
        RECT 116.180 74.970 116.440 75.290 ;
        RECT 111.580 74.630 111.840 74.950 ;
        RECT 111.120 74.350 111.380 74.610 ;
        RECT 111.120 74.290 112.700 74.350 ;
        RECT 113.420 74.290 113.680 74.610 ;
        RECT 113.880 74.290 114.140 74.610 ;
        RECT 114.800 74.290 115.060 74.610 ;
        RECT 111.180 74.270 112.700 74.290 ;
        RECT 111.180 74.210 112.760 74.270 ;
        RECT 109.740 71.570 110.000 71.890 ;
        RECT 110.660 71.570 110.920 71.890 ;
        RECT 108.360 69.530 108.620 69.850 ;
        RECT 109.800 66.790 109.940 71.570 ;
        RECT 111.180 71.550 111.320 74.210 ;
        RECT 112.500 73.950 112.760 74.210 ;
        RECT 111.580 73.610 111.840 73.930 ;
        RECT 111.640 72.910 111.780 73.610 ;
        RECT 111.580 72.590 111.840 72.910 ;
        RECT 113.480 72.570 113.620 74.290 ;
        RECT 113.420 72.250 113.680 72.570 ;
        RECT 113.940 72.230 114.080 74.290 ;
        RECT 114.340 72.590 114.600 72.910 ;
        RECT 113.880 71.910 114.140 72.230 ;
        RECT 112.960 71.570 113.220 71.890 ;
        RECT 111.120 71.230 111.380 71.550 ;
        RECT 112.040 69.870 112.300 70.190 ;
        RECT 110.660 69.190 110.920 69.510 ;
        RECT 110.200 68.170 110.460 68.490 ;
        RECT 110.260 67.130 110.400 68.170 ;
        RECT 110.720 67.470 110.860 69.190 ;
        RECT 112.100 68.830 112.240 69.870 ;
        RECT 112.040 68.510 112.300 68.830 ;
        RECT 110.660 67.150 110.920 67.470 ;
        RECT 110.200 66.810 110.460 67.130 ;
        RECT 109.740 66.470 110.000 66.790 ;
        RECT 110.260 66.110 110.400 66.810 ;
        RECT 110.720 66.790 110.860 67.150 ;
        RECT 113.020 66.790 113.160 71.570 ;
        RECT 113.940 70.190 114.080 71.910 ;
        RECT 113.880 69.870 114.140 70.190 ;
        RECT 113.940 69.170 114.080 69.870 ;
        RECT 113.880 68.850 114.140 69.170 ;
        RECT 113.880 68.170 114.140 68.490 ;
        RECT 113.940 66.790 114.080 68.170 ;
        RECT 110.660 66.470 110.920 66.790 ;
        RECT 112.960 66.470 113.220 66.790 ;
        RECT 113.880 66.470 114.140 66.790 ;
        RECT 114.400 66.700 114.540 72.590 ;
        RECT 114.860 72.230 115.000 74.290 ;
        RECT 114.800 71.910 115.060 72.230 ;
        RECT 115.720 71.910 115.980 72.230 ;
        RECT 114.860 71.550 115.000 71.910 ;
        RECT 114.800 71.230 115.060 71.550 ;
        RECT 114.860 69.510 115.000 71.230 ;
        RECT 114.800 69.190 115.060 69.510 ;
        RECT 115.780 69.170 115.920 71.910 ;
        RECT 116.240 71.890 116.380 74.970 ;
        RECT 119.920 73.930 120.060 82.790 ;
        RECT 121.300 78.350 121.440 88.230 ;
        RECT 126.360 85.830 126.500 93.330 ;
        RECT 128.200 91.950 128.340 96.050 ;
        RECT 128.660 91.950 128.800 96.050 ;
        RECT 129.120 96.030 129.260 99.110 ;
        RECT 129.060 95.710 129.320 96.030 ;
        RECT 129.580 94.330 129.720 101.150 ;
        RECT 130.040 99.770 130.180 106.930 ;
        RECT 130.440 103.530 130.700 103.850 ;
        RECT 130.500 101.810 130.640 103.530 ;
        RECT 130.440 101.490 130.700 101.810 ;
        RECT 130.960 101.130 131.100 108.970 ;
        RECT 131.420 104.870 131.560 112.370 ;
        RECT 131.880 110.390 132.020 112.370 ;
        RECT 132.340 110.990 132.480 115.430 ;
        RECT 132.740 114.410 133.000 114.730 ;
        RECT 132.800 112.690 132.940 114.410 ;
        RECT 132.740 112.370 133.000 112.690 ;
        RECT 134.180 112.010 134.320 118.830 ;
        RECT 135.560 113.370 135.700 177.650 ;
        RECT 136.880 176.970 137.140 177.290 ;
        RECT 136.940 175.930 137.080 176.970 ;
        RECT 136.880 175.610 137.140 175.930 ;
        RECT 138.320 175.590 138.460 179.690 ;
        RECT 138.780 178.990 138.920 180.370 ;
        RECT 140.160 180.010 140.300 184.110 ;
        RECT 141.540 184.090 141.680 185.470 ;
        RECT 141.480 183.770 141.740 184.090 ;
        RECT 141.540 181.710 141.680 183.770 ;
        RECT 141.480 181.390 141.740 181.710 ;
        RECT 141.540 181.030 141.680 181.390 ;
        RECT 141.480 180.710 141.740 181.030 ;
        RECT 140.100 179.690 140.360 180.010 ;
        RECT 139.460 179.155 141.000 179.525 ;
        RECT 138.720 178.670 138.980 178.990 ;
        RECT 141.540 178.390 141.680 180.710 ;
        RECT 142.460 179.070 142.600 202.130 ;
        RECT 144.240 197.370 144.500 197.690 ;
        RECT 142.860 194.310 143.120 194.630 ;
        RECT 142.920 190.890 143.060 194.310 ;
        RECT 142.860 190.570 143.120 190.890 ;
        RECT 143.320 185.130 143.580 185.450 ;
        RECT 143.380 184.430 143.520 185.130 ;
        RECT 143.320 184.110 143.580 184.430 ;
        RECT 144.300 183.945 144.440 197.370 ;
        RECT 144.230 183.575 144.510 183.945 ;
        RECT 143.320 182.410 143.580 182.730 ;
        RECT 143.380 181.370 143.520 182.410 ;
        RECT 144.300 181.370 144.440 183.575 ;
        RECT 143.320 181.050 143.580 181.370 ;
        RECT 144.240 181.050 144.500 181.370 ;
        RECT 142.460 178.930 143.060 179.070 ;
        RECT 140.160 178.250 141.680 178.390 ;
        RECT 140.160 177.630 140.300 178.250 ;
        RECT 142.400 177.990 142.660 178.310 ;
        RECT 141.940 177.650 142.200 177.970 ;
        RECT 138.720 177.310 138.980 177.630 ;
        RECT 140.100 177.310 140.360 177.630 ;
        RECT 138.260 175.270 138.520 175.590 ;
        RECT 138.780 175.250 138.920 177.310 ;
        RECT 141.480 176.970 141.740 177.290 ;
        RECT 141.540 176.270 141.680 176.970 ;
        RECT 142.000 176.270 142.140 177.650 ;
        RECT 141.480 175.950 141.740 176.270 ;
        RECT 141.940 175.950 142.200 176.270 ;
        RECT 142.460 175.930 142.600 177.990 ;
        RECT 142.400 175.610 142.660 175.930 ;
        RECT 138.720 174.930 138.980 175.250 ;
        RECT 142.460 174.990 142.600 175.610 ;
        RECT 136.420 174.250 136.680 174.570 ;
        RECT 136.480 170.830 136.620 174.250 ;
        RECT 138.780 173.550 138.920 174.930 ;
        RECT 142.000 174.850 142.600 174.990 ;
        RECT 139.460 173.715 141.000 174.085 ;
        RECT 142.000 173.550 142.140 174.850 ;
        RECT 142.400 174.250 142.660 174.570 ;
        RECT 138.720 173.230 138.980 173.550 ;
        RECT 139.180 173.230 139.440 173.550 ;
        RECT 141.940 173.230 142.200 173.550 ;
        RECT 136.420 170.510 136.680 170.830 ;
        RECT 139.240 170.150 139.380 173.230 ;
        RECT 139.180 169.830 139.440 170.150 ;
        RECT 142.460 169.130 142.600 174.250 ;
        RECT 142.920 169.810 143.060 178.930 ;
        RECT 143.320 177.650 143.580 177.970 ;
        RECT 144.240 177.650 144.500 177.970 ;
        RECT 143.380 170.830 143.520 177.650 ;
        RECT 143.780 176.970 144.040 177.290 ;
        RECT 143.840 172.190 143.980 176.970 ;
        RECT 144.300 175.930 144.440 177.650 ;
        RECT 144.240 175.610 144.500 175.930 ;
        RECT 143.780 171.870 144.040 172.190 ;
        RECT 143.320 170.510 143.580 170.830 ;
        RECT 142.860 169.490 143.120 169.810 ;
        RECT 142.400 168.810 142.660 169.130 ;
        RECT 139.460 168.275 141.000 168.645 ;
        RECT 135.960 166.770 136.220 167.090 ;
        RECT 137.340 166.770 137.600 167.090 ;
        RECT 136.020 165.390 136.160 166.770 ;
        RECT 135.960 165.070 136.220 165.390 ;
        RECT 136.420 164.730 136.680 165.050 ;
        RECT 136.480 160.970 136.620 164.730 ;
        RECT 137.400 162.670 137.540 166.770 ;
        RECT 139.640 166.090 139.900 166.410 ;
        RECT 144.240 166.090 144.500 166.410 ;
        RECT 139.700 164.710 139.840 166.090 ;
        RECT 139.640 164.390 139.900 164.710 ;
        RECT 139.460 162.835 141.000 163.205 ;
        RECT 137.340 162.350 137.600 162.670 ;
        RECT 144.300 161.310 144.440 166.090 ;
        RECT 144.240 160.990 144.500 161.310 ;
        RECT 136.420 160.650 136.680 160.970 ;
        RECT 136.480 159.610 136.620 160.650 ;
        RECT 136.420 159.290 136.680 159.610 ;
        RECT 137.340 159.290 137.600 159.610 ;
        RECT 135.960 158.950 136.220 159.270 ;
        RECT 136.020 155.870 136.160 158.950 ;
        RECT 136.480 158.590 136.620 159.290 ;
        RECT 136.420 158.270 136.680 158.590 ;
        RECT 135.960 155.550 136.220 155.870 ;
        RECT 135.960 154.190 136.220 154.510 ;
        RECT 136.020 153.150 136.160 154.190 ;
        RECT 135.960 152.830 136.220 153.150 ;
        RECT 136.480 150.770 136.620 158.270 ;
        RECT 137.400 157.230 137.540 159.290 ;
        RECT 137.800 157.930 138.060 158.250 ;
        RECT 138.720 157.930 138.980 158.250 ;
        RECT 137.340 156.910 137.600 157.230 ;
        RECT 137.860 155.530 138.000 157.930 ;
        RECT 138.780 156.210 138.920 157.930 ;
        RECT 139.460 157.395 141.000 157.765 ;
        RECT 138.720 155.890 138.980 156.210 ;
        RECT 137.800 155.210 138.060 155.530 ;
        RECT 136.880 153.850 137.140 154.170 ;
        RECT 136.420 150.450 136.680 150.770 ;
        RECT 136.940 150.430 137.080 153.850 ;
        RECT 137.860 153.490 138.000 155.210 ;
        RECT 137.800 153.170 138.060 153.490 ;
        RECT 139.460 151.955 141.000 152.325 ;
        RECT 136.880 150.110 137.140 150.430 ;
        RECT 136.420 149.770 136.680 150.090 ;
        RECT 143.780 149.770 144.040 150.090 ;
        RECT 135.960 148.070 136.220 148.390 ;
        RECT 136.020 145.670 136.160 148.070 ;
        RECT 136.480 146.350 136.620 149.770 ;
        RECT 136.880 148.410 137.140 148.730 ;
        RECT 136.940 146.350 137.080 148.410 ;
        RECT 139.460 146.515 141.000 146.885 ;
        RECT 136.420 146.030 136.680 146.350 ;
        RECT 136.880 146.030 137.140 146.350 ;
        RECT 141.940 145.690 142.200 146.010 ;
        RECT 135.960 145.350 136.220 145.670 ;
        RECT 136.020 143.630 136.160 145.350 ;
        RECT 142.000 145.330 142.140 145.690 ;
        RECT 143.840 145.330 143.980 149.770 ;
        RECT 144.760 147.710 144.900 212.220 ;
        RECT 152.120 208.230 152.260 212.220 ;
        RECT 156.250 209.075 157.790 209.445 ;
        RECT 152.060 207.910 152.320 208.230 ;
        RECT 147.460 204.850 147.720 205.170 ;
        RECT 145.160 202.810 145.420 203.130 ;
        RECT 145.220 197.010 145.360 202.810 ;
        RECT 147.000 201.790 147.260 202.110 ;
        RECT 147.060 197.350 147.200 201.790 ;
        RECT 147.520 199.730 147.660 204.850 ;
        RECT 156.250 203.635 157.790 204.005 ;
        RECT 154.820 202.130 155.080 202.450 ;
        RECT 154.880 200.750 155.020 202.130 ;
        RECT 154.820 200.430 155.080 200.750 ;
        RECT 147.460 199.410 147.720 199.730 ;
        RECT 150.680 199.410 150.940 199.730 ;
        RECT 147.920 199.070 148.180 199.390 ;
        RECT 147.980 198.030 148.120 199.070 ;
        RECT 147.920 197.710 148.180 198.030 ;
        RECT 147.000 197.030 147.260 197.350 ;
        RECT 145.160 196.690 145.420 197.010 ;
        RECT 145.220 193.950 145.360 196.690 ;
        RECT 145.620 193.970 145.880 194.290 ;
        RECT 145.160 193.630 145.420 193.950 ;
        RECT 145.220 192.250 145.360 193.630 ;
        RECT 145.160 191.930 145.420 192.250 ;
        RECT 145.220 189.270 145.360 191.930 ;
        RECT 145.680 191.230 145.820 193.970 ;
        RECT 146.540 193.290 146.800 193.610 ;
        RECT 146.600 192.250 146.740 193.290 ;
        RECT 146.540 191.930 146.800 192.250 ;
        RECT 150.740 191.910 150.880 199.410 ;
        RECT 156.250 198.195 157.790 198.565 ;
        RECT 156.250 192.755 157.790 193.125 ;
        RECT 150.680 191.590 150.940 191.910 ;
        RECT 145.620 190.910 145.880 191.230 ;
        RECT 145.220 189.130 145.820 189.270 ;
        RECT 145.160 188.530 145.420 188.850 ;
        RECT 145.220 186.810 145.360 188.530 ;
        RECT 145.680 188.170 145.820 189.130 ;
        RECT 150.740 188.850 150.880 191.590 ;
        RECT 146.540 188.530 146.800 188.850 ;
        RECT 150.680 188.530 150.940 188.850 ;
        RECT 145.620 187.850 145.880 188.170 ;
        RECT 145.160 186.490 145.420 186.810 ;
        RECT 145.160 185.810 145.420 186.130 ;
        RECT 145.220 184.430 145.360 185.810 ;
        RECT 145.160 184.110 145.420 184.430 ;
        RECT 145.680 183.410 145.820 187.850 ;
        RECT 146.600 183.750 146.740 188.530 ;
        RECT 149.300 188.190 149.560 188.510 ;
        RECT 147.920 187.850 148.180 188.170 ;
        RECT 147.980 186.470 148.120 187.850 ;
        RECT 149.360 187.150 149.500 188.190 ;
        RECT 156.250 187.315 157.790 187.685 ;
        RECT 149.300 186.830 149.560 187.150 ;
        RECT 147.920 186.150 148.180 186.470 ;
        RECT 146.540 183.430 146.800 183.750 ;
        RECT 145.620 183.090 145.880 183.410 ;
        RECT 145.160 182.750 145.420 183.070 ;
        RECT 145.220 181.030 145.360 182.750 ;
        RECT 145.680 181.710 145.820 183.090 ;
        RECT 146.080 182.750 146.340 183.070 ;
        RECT 146.140 181.710 146.280 182.750 ;
        RECT 145.620 181.390 145.880 181.710 ;
        RECT 146.080 181.390 146.340 181.710 ;
        RECT 145.160 180.710 145.420 181.030 ;
        RECT 145.680 177.710 145.820 181.390 ;
        RECT 146.600 180.600 146.740 183.430 ;
        RECT 156.250 181.875 157.790 182.245 ;
        RECT 149.300 180.710 149.560 181.030 ;
        RECT 147.000 180.600 147.260 180.690 ;
        RECT 146.600 180.460 147.260 180.600 ;
        RECT 147.000 180.370 147.260 180.460 ;
        RECT 147.060 177.970 147.200 180.370 ;
        RECT 145.680 177.570 146.280 177.710 ;
        RECT 146.540 177.650 146.800 177.970 ;
        RECT 147.000 177.650 147.260 177.970 ;
        RECT 145.620 176.970 145.880 177.290 ;
        RECT 145.680 175.590 145.820 176.970 ;
        RECT 146.140 175.930 146.280 177.570 ;
        RECT 146.080 175.610 146.340 175.930 ;
        RECT 146.600 175.590 146.740 177.650 ;
        RECT 145.620 175.270 145.880 175.590 ;
        RECT 146.540 175.270 146.800 175.590 ;
        RECT 145.680 170.490 145.820 175.270 ;
        RECT 147.060 172.530 147.200 177.650 ;
        RECT 148.840 176.970 149.100 177.290 ;
        RECT 147.920 175.610 148.180 175.930 ;
        RECT 147.980 172.870 148.120 175.610 ;
        RECT 148.900 174.570 149.040 176.970 ;
        RECT 148.840 174.250 149.100 174.570 ;
        RECT 147.920 172.550 148.180 172.870 ;
        RECT 147.000 172.210 147.260 172.530 ;
        RECT 145.620 170.170 145.880 170.490 ;
        RECT 145.160 169.490 145.420 169.810 ;
        RECT 145.220 167.430 145.360 169.490 ;
        RECT 147.060 167.430 147.200 172.210 ;
        RECT 147.980 170.150 148.120 172.550 ;
        RECT 148.840 171.530 149.100 171.850 ;
        RECT 147.920 169.830 148.180 170.150 ;
        RECT 145.160 167.110 145.420 167.430 ;
        RECT 147.000 167.110 147.260 167.430 ;
        RECT 145.220 158.930 145.360 167.110 ;
        RECT 147.060 164.690 147.200 167.110 ;
        RECT 148.900 167.090 149.040 171.530 ;
        RECT 148.840 166.770 149.100 167.090 ;
        RECT 147.060 164.550 148.120 164.690 ;
        RECT 147.980 164.370 148.120 164.550 ;
        RECT 147.920 164.050 148.180 164.370 ;
        RECT 147.980 162.670 148.120 164.050 ;
        RECT 147.920 162.350 148.180 162.670 ;
        RECT 147.920 160.990 148.180 161.310 ;
        RECT 147.980 159.950 148.120 160.990 ;
        RECT 147.920 159.630 148.180 159.950 ;
        RECT 145.160 158.610 145.420 158.930 ;
        RECT 149.360 156.210 149.500 180.710 ;
        RECT 150.220 177.310 150.480 177.630 ;
        RECT 150.280 176.270 150.420 177.310 ;
        RECT 154.360 176.970 154.620 177.290 ;
        RECT 149.760 175.950 150.020 176.270 ;
        RECT 150.220 175.950 150.480 176.270 ;
        RECT 149.820 172.530 149.960 175.950 ;
        RECT 154.420 175.590 154.560 176.970 ;
        RECT 156.250 176.435 157.790 176.805 ;
        RECT 154.360 175.270 154.620 175.590 ;
        RECT 149.760 172.210 150.020 172.530 ;
        RECT 153.440 172.210 153.700 172.530 ;
        RECT 153.500 170.830 153.640 172.210 ;
        RECT 156.250 170.995 157.790 171.365 ;
        RECT 153.440 170.510 153.700 170.830 ;
        RECT 154.360 169.490 154.620 169.810 ;
        RECT 154.420 168.110 154.560 169.490 ;
        RECT 154.360 167.790 154.620 168.110 ;
        RECT 156.250 165.555 157.790 165.925 ;
        RECT 154.820 160.650 155.080 160.970 ;
        RECT 154.880 159.270 155.020 160.650 ;
        RECT 156.250 160.115 157.790 160.485 ;
        RECT 154.820 158.950 155.080 159.270 ;
        RECT 149.300 155.890 149.560 156.210 ;
        RECT 155.280 155.550 155.540 155.870 ;
        RECT 155.340 153.490 155.480 155.550 ;
        RECT 156.250 154.675 157.790 155.045 ;
        RECT 155.280 153.170 155.540 153.490 ;
        RECT 155.340 150.770 155.480 153.170 ;
        RECT 145.620 150.450 145.880 150.770 ;
        RECT 155.280 150.450 155.540 150.770 ;
        RECT 144.700 147.390 144.960 147.710 ;
        RECT 144.240 145.690 144.500 146.010 ;
        RECT 141.940 145.010 142.200 145.330 ;
        RECT 143.780 145.010 144.040 145.330 ;
        RECT 139.640 144.330 139.900 144.650 ;
        RECT 135.960 143.310 136.220 143.630 ;
        RECT 139.700 142.950 139.840 144.330 ;
        RECT 142.000 143.630 142.140 145.010 ;
        RECT 141.940 143.310 142.200 143.630 ;
        RECT 143.840 143.290 143.980 145.010 ;
        RECT 144.300 143.630 144.440 145.690 ;
        RECT 145.680 144.990 145.820 150.450 ;
        RECT 148.840 150.110 149.100 150.430 ;
        RECT 148.900 149.070 149.040 150.110 ;
        RECT 148.840 148.750 149.100 149.070 ;
        RECT 147.460 148.070 147.720 148.390 ;
        RECT 147.520 146.350 147.660 148.070 ;
        RECT 147.460 146.030 147.720 146.350 ;
        RECT 155.340 145.330 155.480 150.450 ;
        RECT 156.250 149.235 157.790 149.605 ;
        RECT 155.280 145.010 155.540 145.330 ;
        RECT 145.620 144.670 145.880 144.990 ;
        RECT 147.460 144.670 147.720 144.990 ;
        RECT 152.980 144.670 153.240 144.990 ;
        RECT 144.240 143.310 144.500 143.630 ;
        RECT 143.780 142.970 144.040 143.290 ;
        RECT 139.640 142.630 139.900 142.950 ;
        RECT 143.320 142.630 143.580 142.950 ;
        RECT 141.480 141.610 141.740 141.930 ;
        RECT 139.460 141.075 141.000 141.445 ;
        RECT 135.960 139.570 136.220 139.890 ;
        RECT 140.560 139.570 140.820 139.890 ;
        RECT 136.020 132.750 136.160 139.570 ;
        RECT 137.800 139.230 138.060 139.550 ;
        RECT 137.860 134.790 138.000 139.230 ;
        RECT 140.620 138.190 140.760 139.570 ;
        RECT 140.560 137.870 140.820 138.190 ;
        RECT 141.540 137.850 141.680 141.610 ;
        RECT 141.940 138.890 142.200 139.210 ;
        RECT 141.480 137.530 141.740 137.850 ;
        RECT 139.460 135.635 141.000 136.005 ;
        RECT 137.800 134.470 138.060 134.790 ;
        RECT 141.020 134.360 141.280 134.450 ;
        RECT 141.540 134.360 141.680 137.530 ;
        RECT 142.000 137.510 142.140 138.890 ;
        RECT 143.380 138.190 143.520 142.630 ;
        RECT 143.320 137.870 143.580 138.190 ;
        RECT 142.860 137.530 143.120 137.850 ;
        RECT 141.940 137.190 142.200 137.510 ;
        RECT 142.920 134.450 143.060 137.530 ;
        RECT 144.300 137.510 144.440 143.310 ;
        RECT 144.700 141.950 144.960 142.270 ;
        RECT 145.160 141.950 145.420 142.270 ;
        RECT 144.760 139.550 144.900 141.950 ;
        RECT 145.220 139.890 145.360 141.950 ;
        RECT 147.520 141.930 147.660 144.670 ;
        RECT 148.840 144.330 149.100 144.650 ;
        RECT 150.680 144.330 150.940 144.650 ;
        RECT 148.900 142.950 149.040 144.330 ;
        RECT 150.740 142.950 150.880 144.330 ;
        RECT 153.040 143.630 153.180 144.670 ;
        RECT 152.980 143.310 153.240 143.630 ;
        RECT 155.340 143.290 155.480 145.010 ;
        RECT 156.250 143.795 157.790 144.165 ;
        RECT 155.280 142.970 155.540 143.290 ;
        RECT 148.380 142.630 148.640 142.950 ;
        RECT 148.840 142.630 149.100 142.950 ;
        RECT 149.760 142.630 150.020 142.950 ;
        RECT 150.680 142.630 150.940 142.950 ;
        RECT 152.060 142.630 152.320 142.950 ;
        RECT 148.440 142.350 148.580 142.630 ;
        RECT 149.820 142.350 149.960 142.630 ;
        RECT 148.440 142.210 149.960 142.350 ;
        RECT 152.120 141.930 152.260 142.630 ;
        RECT 147.460 141.610 147.720 141.930 ;
        RECT 152.060 141.610 152.320 141.930 ;
        RECT 145.160 139.570 145.420 139.890 ;
        RECT 144.700 139.230 144.960 139.550 ;
        RECT 146.540 138.890 146.800 139.210 ;
        RECT 146.600 138.190 146.740 138.890 ;
        RECT 146.540 137.870 146.800 138.190 ;
        RECT 144.240 137.190 144.500 137.510 ;
        RECT 147.520 136.490 147.660 141.610 ;
        RECT 148.380 139.570 148.640 139.890 ;
        RECT 144.240 136.170 144.500 136.490 ;
        RECT 147.460 136.170 147.720 136.490 ;
        RECT 144.300 134.790 144.440 136.170 ;
        RECT 144.240 134.470 144.500 134.790 ;
        RECT 148.440 134.450 148.580 139.570 ;
        RECT 150.220 139.230 150.480 139.550 ;
        RECT 150.280 138.190 150.420 139.230 ;
        RECT 156.250 138.355 157.790 138.725 ;
        RECT 150.220 137.870 150.480 138.190 ;
        RECT 141.020 134.220 141.680 134.360 ;
        RECT 141.020 134.130 141.280 134.220 ;
        RECT 142.400 134.130 142.660 134.450 ;
        RECT 142.860 134.130 143.120 134.450 ;
        RECT 143.320 134.130 143.580 134.450 ;
        RECT 148.380 134.130 148.640 134.450 ;
        RECT 141.940 133.450 142.200 133.770 ;
        RECT 135.960 132.430 136.220 132.750 ;
        RECT 142.000 132.070 142.140 133.450 ;
        RECT 142.460 132.750 142.600 134.130 ;
        RECT 142.400 132.430 142.660 132.750 ;
        RECT 142.920 132.070 143.060 134.130 ;
        RECT 143.380 132.070 143.520 134.130 ;
        RECT 141.940 131.750 142.200 132.070 ;
        RECT 142.860 131.750 143.120 132.070 ;
        RECT 143.320 131.750 143.580 132.070 ;
        RECT 144.700 131.750 144.960 132.070 ;
        RECT 138.260 131.410 138.520 131.730 ;
        RECT 138.320 130.030 138.460 131.410 ;
        RECT 139.460 130.195 141.000 130.565 ;
        RECT 138.260 129.710 138.520 130.030 ;
        RECT 144.760 128.670 144.900 131.750 ;
        RECT 148.440 129.350 148.580 134.130 ;
        RECT 151.140 133.450 151.400 133.770 ;
        RECT 151.200 131.730 151.340 133.450 ;
        RECT 156.250 132.915 157.790 133.285 ;
        RECT 152.980 131.750 153.240 132.070 ;
        RECT 151.140 131.410 151.400 131.730 ;
        RECT 151.600 129.710 151.860 130.030 ;
        RECT 145.160 129.030 145.420 129.350 ;
        RECT 148.380 129.030 148.640 129.350 ;
        RECT 136.420 128.350 136.680 128.670 ;
        RECT 144.700 128.350 144.960 128.670 ;
        RECT 136.480 126.630 136.620 128.350 ;
        RECT 136.880 128.010 137.140 128.330 ;
        RECT 136.420 126.310 136.680 126.630 ;
        RECT 136.940 125.610 137.080 128.010 ;
        RECT 145.220 127.310 145.360 129.030 ;
        RECT 138.720 126.990 138.980 127.310 ;
        RECT 145.160 126.990 145.420 127.310 ;
        RECT 137.340 125.970 137.600 126.290 ;
        RECT 136.880 125.290 137.140 125.610 ;
        RECT 135.960 123.930 136.220 124.250 ;
        RECT 136.020 116.090 136.160 123.930 ;
        RECT 136.940 123.570 137.080 125.290 ;
        RECT 136.880 123.250 137.140 123.570 ;
        RECT 136.420 122.570 136.680 122.890 ;
        RECT 136.480 121.190 136.620 122.570 ;
        RECT 136.420 120.870 136.680 121.190 ;
        RECT 136.420 120.190 136.680 120.510 ;
        RECT 136.880 120.190 137.140 120.510 ;
        RECT 136.480 118.470 136.620 120.190 ;
        RECT 136.420 118.150 136.680 118.470 ;
        RECT 136.480 117.450 136.620 118.150 ;
        RECT 136.420 117.130 136.680 117.450 ;
        RECT 136.940 116.430 137.080 120.190 ;
        RECT 137.400 116.430 137.540 125.970 ;
        RECT 137.800 125.860 138.060 125.950 ;
        RECT 138.780 125.860 138.920 126.990 ;
        RECT 144.700 125.970 144.960 126.290 ;
        RECT 137.800 125.720 138.920 125.860 ;
        RECT 137.800 125.630 138.060 125.720 ;
        RECT 139.460 124.755 141.000 125.125 ;
        RECT 138.720 123.250 138.980 123.570 ;
        RECT 144.240 123.250 144.500 123.570 ;
        RECT 137.800 122.570 138.060 122.890 ;
        RECT 137.860 121.530 138.000 122.570 ;
        RECT 137.800 121.210 138.060 121.530 ;
        RECT 138.780 118.810 138.920 123.250 ;
        RECT 141.940 122.910 142.200 123.230 ;
        RECT 141.480 119.850 141.740 120.170 ;
        RECT 139.460 119.315 141.000 119.685 ;
        RECT 138.720 118.490 138.980 118.810 ;
        RECT 136.880 116.110 137.140 116.430 ;
        RECT 137.340 116.110 137.600 116.430 ;
        RECT 141.540 116.090 141.680 119.850 ;
        RECT 135.960 115.770 136.220 116.090 ;
        RECT 141.480 115.770 141.740 116.090 ;
        RECT 142.000 115.750 142.140 122.910 ;
        RECT 142.860 122.570 143.120 122.890 ;
        RECT 141.940 115.430 142.200 115.750 ;
        RECT 142.920 115.070 143.060 122.570 ;
        RECT 144.300 120.850 144.440 123.250 ;
        RECT 144.760 121.530 144.900 125.970 ;
        RECT 145.220 123.570 145.360 126.990 ;
        RECT 148.440 126.970 148.580 129.030 ;
        RECT 151.660 128.750 151.800 129.710 ;
        RECT 151.200 128.610 151.800 128.750 ;
        RECT 148.380 126.650 148.640 126.970 ;
        RECT 148.440 125.950 148.580 126.650 ;
        RECT 148.380 125.630 148.640 125.950 ;
        RECT 145.160 123.250 145.420 123.570 ;
        RECT 147.920 123.480 148.180 123.570 ;
        RECT 148.440 123.480 148.580 125.630 ;
        RECT 148.840 125.290 149.100 125.610 ;
        RECT 148.900 123.570 149.040 125.290 ;
        RECT 147.920 123.340 148.580 123.480 ;
        RECT 147.920 123.250 148.180 123.340 ;
        RECT 148.840 123.250 149.100 123.570 ;
        RECT 147.000 121.550 147.260 121.870 ;
        RECT 144.700 121.210 144.960 121.530 ;
        RECT 144.240 120.530 144.500 120.850 ;
        RECT 144.300 119.150 144.440 120.530 ;
        RECT 144.700 119.850 144.960 120.170 ;
        RECT 145.160 119.850 145.420 120.170 ;
        RECT 144.240 118.830 144.500 119.150 ;
        RECT 144.760 118.130 144.900 119.850 ;
        RECT 144.700 117.810 144.960 118.130 ;
        RECT 145.220 116.430 145.360 119.850 ;
        RECT 146.080 117.470 146.340 117.790 ;
        RECT 146.140 116.430 146.280 117.470 ;
        RECT 145.160 116.110 145.420 116.430 ;
        RECT 146.080 116.110 146.340 116.430 ;
        RECT 147.060 116.090 147.200 121.550 ;
        RECT 147.980 118.470 148.120 123.250 ;
        RECT 148.380 121.210 148.640 121.530 ;
        RECT 147.920 118.150 148.180 118.470 ;
        RECT 147.000 115.770 147.260 116.090 ;
        RECT 142.860 114.750 143.120 115.070 ;
        RECT 135.960 114.410 136.220 114.730 ;
        RECT 135.500 113.050 135.760 113.370 ;
        RECT 136.020 112.350 136.160 114.410 ;
        RECT 139.460 113.875 141.000 114.245 ;
        RECT 143.780 113.620 144.040 113.710 ;
        RECT 144.300 113.650 145.360 113.790 ;
        RECT 144.300 113.620 144.440 113.650 ;
        RECT 143.780 113.480 144.440 113.620 ;
        RECT 143.780 113.390 144.040 113.480 ;
        RECT 144.700 112.600 144.960 112.690 ;
        RECT 143.840 112.460 144.960 112.600 ;
        RECT 135.960 112.030 136.220 112.350 ;
        RECT 138.260 112.030 138.520 112.350 ;
        RECT 134.120 111.690 134.380 112.010 ;
        RECT 135.040 111.690 135.300 112.010 ;
        RECT 132.280 110.670 132.540 110.990 ;
        RECT 135.100 110.650 135.240 111.690 ;
        RECT 136.020 110.990 136.160 112.030 ;
        RECT 137.340 111.750 137.600 112.010 ;
        RECT 137.340 111.690 138.000 111.750 ;
        RECT 137.400 111.610 138.000 111.690 ;
        RECT 137.860 110.990 138.000 111.610 ;
        RECT 135.960 110.670 136.220 110.990 ;
        RECT 137.340 110.670 137.600 110.990 ;
        RECT 137.800 110.670 138.060 110.990 ;
        RECT 131.880 110.250 132.480 110.390 ;
        RECT 135.040 110.330 135.300 110.650 ;
        RECT 131.820 109.650 132.080 109.970 ;
        RECT 131.360 104.550 131.620 104.870 ;
        RECT 131.420 102.830 131.560 104.550 ;
        RECT 131.360 102.510 131.620 102.830 ;
        RECT 131.880 102.490 132.020 109.650 ;
        RECT 132.340 107.590 132.480 110.250 ;
        RECT 132.280 107.270 132.540 107.590 ;
        RECT 134.120 107.270 134.380 107.590 ;
        RECT 134.180 104.870 134.320 107.270 ;
        RECT 136.420 106.930 136.680 107.250 ;
        RECT 136.480 105.550 136.620 106.930 ;
        RECT 137.400 105.550 137.540 110.670 ;
        RECT 137.800 109.310 138.060 109.630 ;
        RECT 137.860 107.250 138.000 109.310 ;
        RECT 138.320 109.290 138.460 112.030 ;
        RECT 142.400 111.690 142.660 112.010 ;
        RECT 142.860 111.690 143.120 112.010 ;
        RECT 138.260 108.970 138.520 109.290 ;
        RECT 137.800 106.930 138.060 107.250 ;
        RECT 136.420 105.230 136.680 105.550 ;
        RECT 137.340 105.230 137.600 105.550 ;
        RECT 132.740 104.550 133.000 104.870 ;
        RECT 134.120 104.550 134.380 104.870 ;
        RECT 135.040 104.550 135.300 104.870 ;
        RECT 136.880 104.550 137.140 104.870 ;
        RECT 131.820 102.170 132.080 102.490 ;
        RECT 130.900 100.810 131.160 101.130 ;
        RECT 129.980 99.450 130.240 99.770 ;
        RECT 132.800 97.390 132.940 104.550 ;
        RECT 133.200 101.490 133.460 101.810 ;
        RECT 133.260 100.110 133.400 101.490 ;
        RECT 133.200 99.790 133.460 100.110 ;
        RECT 132.740 97.070 133.000 97.390 ;
        RECT 135.100 94.670 135.240 104.550 ;
        RECT 136.940 96.370 137.080 104.550 ;
        RECT 136.880 96.050 137.140 96.370 ;
        RECT 137.400 96.110 137.540 105.230 ;
        RECT 137.860 102.150 138.000 106.930 ;
        RECT 138.320 102.830 138.460 108.970 ;
        RECT 139.460 108.435 141.000 108.805 ;
        RECT 141.480 107.270 141.740 107.590 ;
        RECT 139.180 106.590 139.440 106.910 ;
        RECT 139.240 104.190 139.380 106.590 ;
        RECT 141.540 104.870 141.680 107.270 ;
        RECT 142.460 104.870 142.600 111.690 ;
        RECT 142.920 110.990 143.060 111.690 ;
        RECT 142.860 110.670 143.120 110.990 ;
        RECT 142.920 104.870 143.060 110.670 ;
        RECT 143.840 107.590 143.980 112.460 ;
        RECT 144.700 112.370 144.960 112.460 ;
        RECT 143.780 107.270 144.040 107.590 ;
        RECT 143.780 106.590 144.040 106.910 ;
        RECT 141.480 104.550 141.740 104.870 ;
        RECT 142.400 104.550 142.660 104.870 ;
        RECT 142.860 104.550 143.120 104.870 ;
        RECT 139.180 103.870 139.440 104.190 ;
        RECT 138.720 103.530 138.980 103.850 ;
        RECT 138.260 102.510 138.520 102.830 ;
        RECT 137.800 101.830 138.060 102.150 ;
        RECT 138.780 99.430 138.920 103.530 ;
        RECT 139.460 102.995 141.000 103.365 ;
        RECT 141.540 102.150 141.680 104.550 ;
        RECT 142.920 104.190 143.060 104.550 ;
        RECT 142.860 103.870 143.120 104.190 ;
        RECT 140.560 101.830 140.820 102.150 ;
        RECT 141.480 101.830 141.740 102.150 ;
        RECT 140.620 99.430 140.760 101.830 ;
        RECT 142.920 100.110 143.060 103.870 ;
        RECT 143.320 101.490 143.580 101.810 ;
        RECT 143.380 101.130 143.520 101.490 ;
        RECT 143.320 100.810 143.580 101.130 ;
        RECT 142.860 99.790 143.120 100.110 ;
        RECT 138.720 99.110 138.980 99.430 ;
        RECT 140.560 99.110 140.820 99.430 ;
        RECT 141.480 99.110 141.740 99.430 ;
        RECT 140.620 98.410 140.760 99.110 ;
        RECT 140.560 98.090 140.820 98.410 ;
        RECT 139.460 97.555 141.000 97.925 ;
        RECT 140.100 96.390 140.360 96.710 ;
        RECT 137.400 96.030 138.000 96.110 ;
        RECT 137.400 95.970 138.060 96.030 ;
        RECT 137.800 95.710 138.060 95.970 ;
        RECT 137.340 95.370 137.600 95.690 ;
        RECT 135.040 94.350 135.300 94.670 ;
        RECT 129.520 94.010 129.780 94.330 ;
        RECT 137.400 93.990 137.540 95.370 ;
        RECT 137.860 93.990 138.000 95.710 ;
        RECT 140.160 94.670 140.300 96.390 ;
        RECT 140.560 95.710 140.820 96.030 ;
        RECT 140.100 94.350 140.360 94.670 ;
        RECT 140.620 94.330 140.760 95.710 ;
        RECT 141.540 94.670 141.680 99.110 ;
        RECT 143.380 99.090 143.520 100.810 ;
        RECT 143.320 98.770 143.580 99.090 ;
        RECT 141.940 96.050 142.200 96.370 ;
        RECT 141.480 94.350 141.740 94.670 ;
        RECT 140.560 94.010 140.820 94.330 ;
        RECT 136.880 93.670 137.140 93.990 ;
        RECT 137.340 93.670 137.600 93.990 ;
        RECT 137.800 93.670 138.060 93.990 ;
        RECT 140.100 93.670 140.360 93.990 ;
        RECT 136.940 93.390 137.080 93.670 ;
        RECT 140.160 93.390 140.300 93.670 ;
        RECT 136.940 93.250 140.300 93.390 ;
        RECT 129.520 92.650 129.780 92.970 ;
        RECT 128.140 91.630 128.400 91.950 ;
        RECT 128.600 91.630 128.860 91.950 ;
        RECT 129.580 91.270 129.720 92.650 ;
        RECT 129.520 90.950 129.780 91.270 ;
        RECT 129.580 90.250 129.720 90.950 ;
        RECT 129.980 90.610 130.240 90.930 ;
        RECT 135.040 90.610 135.300 90.930 ;
        RECT 136.420 90.610 136.680 90.930 ;
        RECT 137.800 90.610 138.060 90.930 ;
        RECT 129.520 89.930 129.780 90.250 ;
        RECT 130.040 88.890 130.180 90.610 ;
        RECT 132.740 89.930 133.000 90.250 ;
        RECT 127.220 88.570 127.480 88.890 ;
        RECT 129.980 88.570 130.240 88.890 ;
        RECT 126.300 85.510 126.560 85.830 ;
        RECT 122.670 83.955 124.210 84.325 ;
        RECT 127.280 83.190 127.420 88.570 ;
        RECT 132.800 87.870 132.940 89.930 ;
        RECT 135.100 87.870 135.240 90.610 ;
        RECT 136.480 88.550 136.620 90.610 ;
        RECT 137.860 88.550 138.000 90.610 ;
        RECT 136.420 88.230 136.680 88.550 ;
        RECT 137.800 88.230 138.060 88.550 ;
        RECT 132.740 87.550 133.000 87.870 ;
        RECT 135.040 87.550 135.300 87.870 ;
        RECT 128.140 87.210 128.400 87.530 ;
        RECT 128.200 85.490 128.340 87.210 ;
        RECT 128.140 85.170 128.400 85.490 ;
        RECT 134.580 85.170 134.840 85.490 ;
        RECT 129.060 83.470 129.320 83.790 ;
        RECT 127.680 83.190 127.940 83.450 ;
        RECT 127.280 83.130 127.940 83.190 ;
        RECT 127.280 83.050 127.880 83.130 ;
        RECT 128.600 82.790 128.860 83.110 ;
        RECT 124.460 81.770 124.720 82.090 ;
        RECT 124.520 80.050 124.660 81.770 ;
        RECT 128.660 81.070 128.800 82.790 ;
        RECT 129.120 81.070 129.260 83.470 ;
        RECT 129.520 83.130 129.780 83.450 ;
        RECT 128.600 80.750 128.860 81.070 ;
        RECT 129.060 80.750 129.320 81.070 ;
        RECT 128.660 80.050 128.800 80.750 ;
        RECT 129.580 80.050 129.720 83.130 ;
        RECT 134.640 83.110 134.780 85.170 ;
        RECT 135.100 83.790 135.240 87.550 ;
        RECT 136.480 86.510 136.620 88.230 ;
        RECT 136.420 86.190 136.680 86.510 ;
        RECT 137.860 85.830 138.000 88.230 ;
        RECT 137.800 85.510 138.060 85.830 ;
        RECT 135.500 84.490 135.760 84.810 ;
        RECT 135.040 83.470 135.300 83.790 ;
        RECT 135.560 83.110 135.700 84.490 ;
        RECT 134.580 82.790 134.840 83.110 ;
        RECT 135.500 82.790 135.760 83.110 ;
        RECT 132.740 81.770 133.000 82.090 ;
        RECT 132.800 80.390 132.940 81.770 ;
        RECT 132.740 80.070 133.000 80.390 ;
        RECT 124.460 79.730 124.720 80.050 ;
        RECT 128.600 79.730 128.860 80.050 ;
        RECT 129.520 79.730 129.780 80.050 ;
        RECT 130.440 79.730 130.700 80.050 ;
        RECT 122.670 78.515 124.210 78.885 ;
        RECT 121.240 78.030 121.500 78.350 ;
        RECT 123.540 77.350 123.800 77.670 ;
        RECT 129.060 77.350 129.320 77.670 ;
        RECT 123.600 74.950 123.740 77.350 ;
        RECT 123.540 74.630 123.800 74.950 ;
        RECT 126.760 74.630 127.020 74.950 ;
        RECT 120.780 73.950 121.040 74.270 ;
        RECT 122.160 73.950 122.420 74.270 ;
        RECT 119.860 73.610 120.120 73.930 ;
        RECT 120.840 72.230 120.980 73.950 ;
        RECT 122.220 72.910 122.360 73.950 ;
        RECT 122.670 73.075 124.210 73.445 ;
        RECT 122.160 72.590 122.420 72.910 ;
        RECT 120.780 71.910 121.040 72.230 ;
        RECT 123.540 71.910 123.800 72.230 ;
        RECT 116.180 71.570 116.440 71.890 ;
        RECT 120.320 69.870 120.580 70.190 ;
        RECT 115.720 68.850 115.980 69.170 ;
        RECT 120.380 67.470 120.520 69.870 ;
        RECT 120.840 69.170 120.980 71.910 ;
        RECT 123.080 71.570 123.340 71.890 ;
        RECT 123.140 71.210 123.280 71.570 ;
        RECT 122.160 70.890 122.420 71.210 ;
        RECT 123.080 70.890 123.340 71.210 ;
        RECT 122.220 69.510 122.360 70.890 ;
        RECT 123.600 70.270 123.740 71.910 ;
        RECT 126.820 71.210 126.960 74.630 ;
        RECT 129.120 72.910 129.260 77.350 ;
        RECT 130.500 77.330 130.640 79.730 ;
        RECT 134.640 78.350 134.780 82.790 ;
        RECT 138.320 80.730 138.460 93.250 ;
        RECT 139.460 92.115 141.000 92.485 ;
        RECT 138.720 90.270 138.980 90.590 ;
        RECT 138.780 88.550 138.920 90.270 ;
        RECT 138.720 88.230 138.980 88.550 ;
        RECT 139.460 86.675 141.000 87.045 ;
        RECT 142.000 86.510 142.140 96.050 ;
        RECT 143.840 95.690 143.980 106.590 ;
        RECT 144.240 106.250 144.500 106.570 ;
        RECT 144.700 106.250 144.960 106.570 ;
        RECT 144.300 105.210 144.440 106.250 ;
        RECT 144.240 104.890 144.500 105.210 ;
        RECT 144.760 101.470 144.900 106.250 ;
        RECT 145.220 101.810 145.360 113.650 ;
        RECT 147.980 113.030 148.120 118.150 ;
        RECT 148.440 115.750 148.580 121.210 ;
        RECT 151.200 120.170 151.340 128.610 ;
        RECT 152.060 128.350 152.320 128.670 ;
        RECT 151.140 119.850 151.400 120.170 ;
        RECT 151.200 118.130 151.340 119.850 ;
        RECT 151.140 117.810 151.400 118.130 ;
        RECT 150.220 117.130 150.480 117.450 ;
        RECT 150.280 115.750 150.420 117.130 ;
        RECT 152.120 116.430 152.260 128.350 ;
        RECT 153.040 126.630 153.180 131.750 ;
        RECT 154.820 131.410 155.080 131.730 ;
        RECT 153.900 131.070 154.160 131.390 ;
        RECT 153.440 130.730 153.700 131.050 ;
        RECT 152.980 126.310 153.240 126.630 ;
        RECT 153.040 121.870 153.180 126.310 ;
        RECT 152.980 121.550 153.240 121.870 ;
        RECT 152.980 120.870 153.240 121.190 ;
        RECT 152.060 116.110 152.320 116.430 ;
        RECT 148.380 115.430 148.640 115.750 ;
        RECT 150.220 115.430 150.480 115.750 ;
        RECT 148.440 115.070 148.580 115.430 ;
        RECT 150.680 115.090 150.940 115.410 ;
        RECT 148.380 114.750 148.640 115.070 ;
        RECT 148.440 113.710 148.580 114.750 ;
        RECT 148.380 113.390 148.640 113.710 ;
        RECT 147.920 112.710 148.180 113.030 ;
        RECT 145.620 112.370 145.880 112.690 ;
        RECT 145.680 105.210 145.820 112.370 ;
        RECT 150.740 110.990 150.880 115.090 ;
        RECT 153.040 113.710 153.180 120.870 ;
        RECT 153.500 115.750 153.640 130.730 ;
        RECT 153.960 116.390 154.100 131.070 ;
        RECT 154.880 130.030 155.020 131.410 ;
        RECT 154.820 129.710 155.080 130.030 ;
        RECT 154.360 128.010 154.620 128.330 ;
        RECT 154.420 126.630 154.560 128.010 ;
        RECT 156.250 127.475 157.790 127.845 ;
        RECT 154.360 126.310 154.620 126.630 ;
        RECT 154.820 126.310 155.080 126.630 ;
        RECT 154.360 122.570 154.620 122.890 ;
        RECT 154.420 121.190 154.560 122.570 ;
        RECT 154.360 120.870 154.620 121.190 ;
        RECT 153.960 116.250 154.560 116.390 ;
        RECT 154.420 115.750 154.560 116.250 ;
        RECT 154.880 116.090 155.020 126.310 ;
        RECT 156.250 122.035 157.790 122.405 ;
        RECT 155.280 120.530 155.540 120.850 ;
        RECT 155.340 119.150 155.480 120.530 ;
        RECT 155.280 118.830 155.540 119.150 ;
        RECT 154.820 115.770 155.080 116.090 ;
        RECT 153.440 115.430 153.700 115.750 ;
        RECT 154.360 115.430 154.620 115.750 ;
        RECT 152.980 113.390 153.240 113.710 ;
        RECT 154.820 113.390 155.080 113.710 ;
        RECT 152.060 112.370 152.320 112.690 ;
        RECT 150.680 110.670 150.940 110.990 ;
        RECT 147.920 109.650 148.180 109.970 ;
        RECT 150.220 109.650 150.480 109.970 ;
        RECT 147.000 108.970 147.260 109.290 ;
        RECT 147.060 108.270 147.200 108.970 ;
        RECT 147.000 107.950 147.260 108.270 ;
        RECT 147.980 107.250 148.120 109.650 ;
        RECT 146.540 106.930 146.800 107.250 ;
        RECT 147.920 106.930 148.180 107.250 ;
        RECT 145.620 104.890 145.880 105.210 ;
        RECT 145.620 104.210 145.880 104.530 ;
        RECT 145.680 102.830 145.820 104.210 ;
        RECT 145.620 102.510 145.880 102.830 ;
        RECT 145.160 101.490 145.420 101.810 ;
        RECT 145.620 101.490 145.880 101.810 ;
        RECT 146.080 101.490 146.340 101.810 ;
        RECT 144.700 101.150 144.960 101.470 ;
        RECT 145.680 101.130 145.820 101.490 ;
        RECT 145.620 100.810 145.880 101.130 ;
        RECT 145.680 100.110 145.820 100.810 ;
        RECT 145.620 99.790 145.880 100.110 ;
        RECT 146.140 99.770 146.280 101.490 ;
        RECT 144.240 99.450 144.500 99.770 ;
        RECT 146.080 99.450 146.340 99.770 ;
        RECT 143.780 95.370 144.040 95.690 ;
        RECT 142.400 94.010 142.660 94.330 ;
        RECT 142.460 89.230 142.600 94.010 ;
        RECT 143.840 93.990 143.980 95.370 ;
        RECT 144.300 94.670 144.440 99.450 ;
        RECT 144.700 98.090 144.960 98.410 ;
        RECT 144.760 96.370 144.900 98.090 ;
        RECT 144.700 96.050 144.960 96.370 ;
        RECT 145.160 95.710 145.420 96.030 ;
        RECT 144.240 94.350 144.500 94.670 ;
        RECT 143.780 93.670 144.040 93.990 ;
        RECT 142.860 90.610 143.120 90.930 ;
        RECT 142.400 88.910 142.660 89.230 ;
        RECT 142.920 86.510 143.060 90.610 ;
        RECT 145.220 90.590 145.360 95.710 ;
        RECT 146.600 95.690 146.740 106.930 ;
        RECT 147.460 106.250 147.720 106.570 ;
        RECT 147.520 102.830 147.660 106.250 ;
        RECT 147.460 102.510 147.720 102.830 ;
        RECT 147.980 101.810 148.120 106.930 ;
        RECT 150.280 104.190 150.420 109.650 ;
        RECT 150.740 105.550 150.880 110.670 ;
        RECT 152.120 105.550 152.260 112.370 ;
        RECT 154.360 107.950 154.620 108.270 ;
        RECT 150.680 105.230 150.940 105.550 ;
        RECT 152.060 105.230 152.320 105.550 ;
        RECT 150.220 103.870 150.480 104.190 ;
        RECT 147.920 101.490 148.180 101.810 ;
        RECT 151.140 101.490 151.400 101.810 ;
        RECT 147.980 96.370 148.120 101.490 ;
        RECT 148.840 101.150 149.100 101.470 ;
        RECT 148.900 100.110 149.040 101.150 ;
        RECT 150.220 100.810 150.480 101.130 ;
        RECT 148.840 99.790 149.100 100.110 ;
        RECT 149.760 99.790 150.020 100.110 ;
        RECT 147.920 96.050 148.180 96.370 ;
        RECT 148.380 95.710 148.640 96.030 ;
        RECT 146.540 95.370 146.800 95.690 ;
        RECT 146.600 94.330 146.740 95.370 ;
        RECT 148.440 94.670 148.580 95.710 ;
        RECT 148.380 94.350 148.640 94.670 ;
        RECT 146.540 94.010 146.800 94.330 ;
        RECT 149.300 93.670 149.560 93.990 ;
        RECT 149.360 91.950 149.500 93.670 ;
        RECT 149.300 91.630 149.560 91.950 ;
        RECT 145.160 90.270 145.420 90.590 ;
        RECT 143.780 88.230 144.040 88.550 ;
        RECT 143.840 87.530 143.980 88.230 ;
        RECT 143.780 87.210 144.040 87.530 ;
        RECT 141.940 86.190 142.200 86.510 ;
        RECT 142.860 86.190 143.120 86.510 ;
        RECT 141.480 82.110 141.740 82.430 ;
        RECT 139.460 81.235 141.000 81.605 ;
        RECT 141.540 81.070 141.680 82.110 ;
        RECT 141.480 80.750 141.740 81.070 ;
        RECT 138.260 80.410 138.520 80.730 ;
        RECT 135.960 79.730 136.220 80.050 ;
        RECT 142.000 79.790 142.140 86.190 ;
        RECT 143.320 83.130 143.580 83.450 ;
        RECT 142.860 81.770 143.120 82.090 ;
        RECT 142.920 80.050 143.060 81.770 ;
        RECT 143.380 80.390 143.520 83.130 ;
        RECT 143.840 82.090 143.980 87.210 ;
        RECT 143.780 81.770 144.040 82.090 ;
        RECT 143.320 80.070 143.580 80.390 ;
        RECT 136.020 78.350 136.160 79.730 ;
        RECT 142.000 79.650 142.600 79.790 ;
        RECT 142.860 79.730 143.120 80.050 ;
        RECT 141.940 79.050 142.200 79.370 ;
        RECT 142.000 78.350 142.140 79.050 ;
        RECT 134.580 78.030 134.840 78.350 ;
        RECT 135.960 78.030 136.220 78.350 ;
        RECT 141.940 78.030 142.200 78.350 ;
        RECT 136.880 77.350 137.140 77.670 ;
        RECT 130.440 77.010 130.700 77.330 ;
        RECT 136.940 75.630 137.080 77.350 ;
        RECT 142.460 76.650 142.600 79.650 ;
        RECT 142.920 78.350 143.060 79.730 ;
        RECT 142.860 78.030 143.120 78.350 ;
        RECT 143.840 77.670 143.980 81.770 ;
        RECT 145.220 80.390 145.360 90.270 ;
        RECT 146.540 88.570 146.800 88.890 ;
        RECT 145.620 88.230 145.880 88.550 ;
        RECT 146.080 88.230 146.340 88.550 ;
        RECT 145.680 87.530 145.820 88.230 ;
        RECT 146.140 87.870 146.280 88.230 ;
        RECT 146.080 87.550 146.340 87.870 ;
        RECT 145.620 87.210 145.880 87.530 ;
        RECT 145.620 85.170 145.880 85.490 ;
        RECT 145.160 80.070 145.420 80.390 ;
        RECT 143.780 77.350 144.040 77.670 ;
        RECT 142.400 76.330 142.660 76.650 ;
        RECT 139.460 75.795 141.000 76.165 ;
        RECT 131.820 75.310 132.080 75.630 ;
        RECT 136.880 75.310 137.140 75.630 ;
        RECT 130.900 74.290 131.160 74.610 ;
        RECT 129.060 72.590 129.320 72.910 ;
        RECT 128.140 71.230 128.400 71.550 ;
        RECT 126.760 70.890 127.020 71.210 ;
        RECT 123.140 70.130 123.740 70.270 ;
        RECT 123.140 69.850 123.280 70.130 ;
        RECT 123.080 69.530 123.340 69.850 ;
        RECT 122.160 69.190 122.420 69.510 ;
        RECT 120.780 68.850 121.040 69.170 ;
        RECT 121.700 68.170 121.960 68.490 ;
        RECT 120.320 67.150 120.580 67.470 ;
        RECT 120.380 66.790 120.520 67.150 ;
        RECT 121.760 66.790 121.900 68.170 ;
        RECT 122.220 67.130 122.360 69.190 ;
        RECT 128.200 69.170 128.340 71.230 ;
        RECT 130.440 70.890 130.700 71.210 ;
        RECT 130.500 70.190 130.640 70.890 ;
        RECT 129.060 69.870 129.320 70.190 ;
        RECT 129.520 69.870 129.780 70.190 ;
        RECT 130.440 69.870 130.700 70.190 ;
        RECT 129.120 69.170 129.260 69.870 ;
        RECT 128.140 69.025 128.400 69.170 ;
        RECT 128.130 68.655 128.410 69.025 ;
        RECT 129.060 68.850 129.320 69.170 ;
        RECT 129.580 68.830 129.720 69.870 ;
        RECT 129.980 69.190 130.240 69.510 ;
        RECT 129.520 68.510 129.780 68.830 ;
        RECT 122.670 67.635 124.210 68.005 ;
        RECT 122.160 66.810 122.420 67.130 ;
        RECT 130.040 66.790 130.180 69.190 ;
        RECT 114.800 66.700 115.060 66.790 ;
        RECT 114.400 66.560 115.060 66.700 ;
        RECT 110.200 65.790 110.460 66.110 ;
        RECT 108.360 65.450 108.620 65.770 ;
        RECT 112.500 65.450 112.760 65.770 ;
        RECT 105.880 64.915 107.420 65.285 ;
        RECT 106.520 63.410 106.780 63.730 ;
        RECT 107.900 63.410 108.160 63.730 ;
        RECT 105.140 61.370 105.400 61.690 ;
        RECT 106.580 61.350 106.720 63.410 ;
        RECT 103.760 61.260 104.020 61.350 ;
        RECT 103.360 61.120 104.020 61.260 ;
        RECT 101.920 57.970 102.180 58.290 ;
        RECT 102.840 57.970 103.100 58.290 ;
        RECT 103.360 56.220 103.500 61.120 ;
        RECT 103.760 61.030 104.020 61.120 ;
        RECT 106.520 61.030 106.780 61.350 ;
        RECT 105.880 59.475 107.420 59.845 ;
        RECT 107.960 58.290 108.100 63.410 ;
        RECT 108.420 58.290 108.560 65.450 ;
        RECT 109.280 63.410 109.540 63.730 ;
        RECT 108.820 61.710 109.080 62.030 ;
        RECT 106.060 57.970 106.320 58.290 ;
        RECT 107.900 57.970 108.160 58.290 ;
        RECT 108.360 57.970 108.620 58.290 ;
        RECT 106.120 56.220 106.260 57.970 ;
        RECT 108.880 56.220 109.020 61.710 ;
        RECT 109.340 61.690 109.480 63.410 ;
        RECT 112.560 61.690 112.700 65.450 ;
        RECT 114.400 64.750 114.540 66.560 ;
        RECT 114.800 66.470 115.060 66.560 ;
        RECT 120.320 66.470 120.580 66.790 ;
        RECT 121.700 66.470 121.960 66.790 ;
        RECT 123.540 66.700 123.800 66.790 ;
        RECT 123.140 66.560 123.800 66.700 ;
        RECT 114.800 65.450 115.060 65.770 ;
        RECT 115.260 65.450 115.520 65.770 ;
        RECT 118.940 65.450 119.200 65.770 ;
        RECT 121.240 65.450 121.500 65.770 ;
        RECT 114.340 64.430 114.600 64.750 ;
        RECT 113.420 63.410 113.680 63.730 ;
        RECT 109.280 61.370 109.540 61.690 ;
        RECT 112.500 61.370 112.760 61.690 ;
        RECT 113.480 58.630 113.620 63.410 ;
        RECT 114.340 61.030 114.600 61.350 ;
        RECT 113.420 58.310 113.680 58.630 ;
        RECT 111.580 57.970 111.840 58.290 ;
        RECT 111.640 56.220 111.780 57.970 ;
        RECT 114.400 56.220 114.540 61.030 ;
        RECT 114.860 58.290 115.000 65.450 ;
        RECT 115.320 61.690 115.460 65.450 ;
        RECT 119.000 63.730 119.140 65.450 ;
        RECT 116.180 63.410 116.440 63.730 ;
        RECT 118.940 63.410 119.200 63.730 ;
        RECT 115.260 61.370 115.520 61.690 ;
        RECT 116.240 61.010 116.380 63.410 ;
        RECT 120.320 61.030 120.580 61.350 ;
        RECT 116.180 60.690 116.440 61.010 ;
        RECT 119.860 60.010 120.120 60.330 ;
        RECT 119.920 58.630 120.060 60.010 ;
        RECT 119.860 58.310 120.120 58.630 ;
        RECT 114.800 57.970 115.060 58.290 ;
        RECT 117.100 57.970 117.360 58.290 ;
        RECT 120.380 58.030 120.520 61.030 ;
        RECT 121.300 58.290 121.440 65.450 ;
        RECT 123.140 64.410 123.280 66.560 ;
        RECT 123.540 66.470 123.800 66.560 ;
        RECT 129.980 66.470 130.240 66.790 ;
        RECT 130.960 66.110 131.100 74.290 ;
        RECT 131.880 73.930 132.020 75.310 ;
        RECT 134.580 74.290 134.840 74.610 ;
        RECT 135.960 74.290 136.220 74.610 ;
        RECT 138.720 74.290 138.980 74.610 ;
        RECT 131.820 73.610 132.080 73.930 ;
        RECT 132.740 71.910 133.000 72.230 ;
        RECT 132.800 70.190 132.940 71.910 ;
        RECT 134.120 71.570 134.380 71.890 ;
        RECT 132.740 69.870 133.000 70.190 ;
        RECT 131.360 66.470 131.620 66.790 ;
        RECT 130.900 65.790 131.160 66.110 ;
        RECT 127.680 65.450 127.940 65.770 ;
        RECT 123.080 64.090 123.340 64.410 ;
        RECT 122.160 63.410 122.420 63.730 ;
        RECT 126.760 63.410 127.020 63.730 ;
        RECT 117.160 56.220 117.300 57.970 ;
        RECT 119.920 57.890 120.520 58.030 ;
        RECT 121.240 57.970 121.500 58.290 ;
        RECT 119.920 56.220 120.060 57.890 ;
        RECT 122.220 56.590 122.360 63.410 ;
        RECT 122.670 62.195 124.210 62.565 ;
        RECT 126.300 60.690 126.560 61.010 ;
        RECT 126.360 59.310 126.500 60.690 ;
        RECT 126.820 59.310 126.960 63.410 ;
        RECT 127.740 61.350 127.880 65.450 ;
        RECT 130.960 64.150 131.100 65.790 ;
        RECT 131.420 64.750 131.560 66.470 ;
        RECT 131.360 64.430 131.620 64.750 ;
        RECT 130.960 64.010 131.560 64.150 ;
        RECT 131.820 64.090 132.080 64.410 ;
        RECT 130.900 63.410 131.160 63.730 ;
        RECT 127.680 61.030 127.940 61.350 ;
        RECT 128.140 61.030 128.400 61.350 ;
        RECT 126.300 58.990 126.560 59.310 ;
        RECT 126.760 58.990 127.020 59.310 ;
        RECT 125.380 57.970 125.640 58.290 ;
        RECT 122.670 56.755 124.210 57.125 ;
        RECT 122.160 56.270 122.420 56.590 ;
        RECT 123.080 56.500 123.340 56.590 ;
        RECT 122.680 56.360 123.340 56.500 ;
        RECT 122.680 56.220 122.820 56.360 ;
        RECT 123.080 56.270 123.340 56.360 ;
        RECT 125.440 56.220 125.580 57.970 ;
        RECT 128.200 56.220 128.340 61.030 ;
        RECT 130.960 56.220 131.100 63.410 ;
        RECT 131.420 61.690 131.560 64.010 ;
        RECT 131.360 61.370 131.620 61.690 ;
        RECT 131.880 58.290 132.020 64.090 ;
        RECT 132.280 63.410 132.540 63.730 ;
        RECT 132.340 61.350 132.480 63.410 ;
        RECT 132.280 61.030 132.540 61.350 ;
        RECT 132.800 58.290 132.940 69.870 ;
        RECT 134.180 69.510 134.320 71.570 ;
        RECT 134.640 71.210 134.780 74.290 ;
        RECT 135.500 72.250 135.760 72.570 ;
        RECT 134.580 70.890 134.840 71.210 ;
        RECT 134.640 70.190 134.780 70.890 ;
        RECT 134.580 69.870 134.840 70.190 ;
        RECT 134.120 69.190 134.380 69.510 ;
        RECT 134.180 68.090 134.320 69.190 ;
        RECT 134.640 68.910 134.780 69.870 ;
        RECT 135.560 69.025 135.700 72.250 ;
        RECT 136.020 72.230 136.160 74.290 ;
        RECT 136.880 73.610 137.140 73.930 ;
        RECT 135.960 71.910 136.220 72.230 ;
        RECT 136.940 70.190 137.080 73.610 ;
        RECT 138.260 70.890 138.520 71.210 ;
        RECT 136.880 69.870 137.140 70.190 ;
        RECT 138.320 69.170 138.460 70.890 ;
        RECT 138.780 70.100 138.920 74.290 ;
        RECT 145.680 72.910 145.820 85.170 ;
        RECT 146.140 83.790 146.280 87.550 ;
        RECT 146.600 86.510 146.740 88.570 ;
        RECT 149.820 88.550 149.960 99.790 ;
        RECT 150.280 98.750 150.420 100.810 ;
        RECT 151.200 99.430 151.340 101.490 ;
        RECT 154.420 99.430 154.560 107.950 ;
        RECT 154.880 104.870 155.020 113.390 ;
        RECT 155.340 110.310 155.480 118.830 ;
        RECT 156.250 116.595 157.790 116.965 ;
        RECT 156.250 111.155 157.790 111.525 ;
        RECT 155.280 109.990 155.540 110.310 ;
        RECT 155.280 108.970 155.540 109.290 ;
        RECT 154.820 104.550 155.080 104.870 ;
        RECT 155.340 102.490 155.480 108.970 ;
        RECT 156.250 105.715 157.790 106.085 ;
        RECT 155.280 102.170 155.540 102.490 ;
        RECT 150.680 99.110 150.940 99.430 ;
        RECT 151.140 99.110 151.400 99.430 ;
        RECT 154.360 99.110 154.620 99.430 ;
        RECT 150.220 98.430 150.480 98.750 ;
        RECT 150.280 94.670 150.420 98.430 ;
        RECT 150.220 94.350 150.480 94.670 ;
        RECT 150.220 89.930 150.480 90.250 ;
        RECT 147.000 88.230 147.260 88.550 ;
        RECT 149.760 88.230 150.020 88.550 ;
        RECT 147.060 86.510 147.200 88.230 ;
        RECT 148.380 87.210 148.640 87.530 ;
        RECT 146.540 86.190 146.800 86.510 ;
        RECT 147.000 86.190 147.260 86.510 ;
        RECT 148.440 85.150 148.580 87.210 ;
        RECT 149.760 85.510 150.020 85.830 ;
        RECT 149.820 85.150 149.960 85.510 ;
        RECT 150.280 85.490 150.420 89.930 ;
        RECT 150.740 88.550 150.880 99.110 ;
        RECT 151.200 93.990 151.340 99.110 ;
        RECT 152.060 98.090 152.320 98.410 ;
        RECT 152.120 94.670 152.260 98.090 ;
        RECT 154.360 95.370 154.620 95.690 ;
        RECT 152.060 94.350 152.320 94.670 ;
        RECT 151.140 93.670 151.400 93.990 ;
        RECT 152.120 89.230 152.260 94.350 ;
        RECT 153.900 93.330 154.160 93.650 ;
        RECT 152.060 88.910 152.320 89.230 ;
        RECT 153.960 88.550 154.100 93.330 ;
        RECT 154.420 91.270 154.560 95.370 ;
        RECT 155.340 93.990 155.480 102.170 ;
        RECT 156.250 100.275 157.790 100.645 ;
        RECT 156.250 94.835 157.790 95.205 ;
        RECT 155.280 93.670 155.540 93.990 ;
        RECT 154.360 90.950 154.620 91.270 ;
        RECT 156.250 89.395 157.790 89.765 ;
        RECT 150.680 88.230 150.940 88.550 ;
        RECT 153.900 88.230 154.160 88.550 ;
        RECT 150.220 85.170 150.480 85.490 ;
        RECT 148.380 84.830 148.640 85.150 ;
        RECT 149.760 84.830 150.020 85.150 ;
        RECT 156.250 83.955 157.790 84.325 ;
        RECT 146.080 83.470 146.340 83.790 ;
        RECT 146.080 82.790 146.340 83.110 ;
        RECT 147.000 82.790 147.260 83.110 ;
        RECT 148.380 82.790 148.640 83.110 ;
        RECT 146.140 76.990 146.280 82.790 ;
        RECT 146.540 81.770 146.800 82.090 ;
        RECT 146.600 80.050 146.740 81.770 ;
        RECT 146.540 79.730 146.800 80.050 ;
        RECT 147.060 78.010 147.200 82.790 ;
        RECT 148.440 79.370 148.580 82.790 ;
        RECT 148.380 79.050 148.640 79.370 ;
        RECT 148.440 78.010 148.580 79.050 ;
        RECT 156.250 78.515 157.790 78.885 ;
        RECT 147.000 77.690 147.260 78.010 ;
        RECT 148.380 77.690 148.640 78.010 ;
        RECT 146.080 76.670 146.340 76.990 ;
        RECT 147.060 75.630 147.200 77.690 ;
        RECT 147.000 75.310 147.260 75.630 ;
        RECT 156.250 73.075 157.790 73.445 ;
        RECT 145.620 72.590 145.880 72.910 ;
        RECT 143.780 71.910 144.040 72.230 ;
        RECT 139.460 70.355 141.000 70.725 ;
        RECT 143.840 70.190 143.980 71.910 ;
        RECT 145.160 70.890 145.420 71.210 ;
        RECT 139.640 70.100 139.900 70.190 ;
        RECT 138.780 69.960 139.900 70.100 ;
        RECT 139.640 69.870 139.900 69.960 ;
        RECT 141.480 69.870 141.740 70.190 ;
        RECT 143.780 69.870 144.040 70.190 ;
        RECT 134.640 68.770 135.240 68.910 ;
        RECT 134.180 67.950 134.780 68.090 ;
        RECT 134.640 61.690 134.780 67.950 ;
        RECT 135.100 65.770 135.240 68.770 ;
        RECT 135.490 68.655 135.770 69.025 ;
        RECT 138.260 68.850 138.520 69.170 ;
        RECT 141.020 68.850 141.280 69.170 ;
        RECT 135.500 68.510 135.760 68.655 ;
        RECT 135.560 67.470 135.700 68.510 ;
        RECT 135.500 67.150 135.760 67.470 ;
        RECT 141.080 66.110 141.220 68.850 ;
        RECT 141.540 67.470 141.680 69.870 ;
        RECT 145.220 69.170 145.360 70.890 ;
        RECT 146.540 69.190 146.800 69.510 ;
        RECT 145.160 68.850 145.420 69.170 ;
        RECT 145.620 68.170 145.880 68.490 ;
        RECT 141.480 67.150 141.740 67.470 ;
        RECT 138.260 65.790 138.520 66.110 ;
        RECT 141.020 65.790 141.280 66.110 ;
        RECT 135.040 65.450 135.300 65.770 ;
        RECT 137.800 63.750 138.060 64.070 ;
        RECT 136.880 63.410 137.140 63.730 ;
        RECT 134.580 61.370 134.840 61.690 ;
        RECT 134.120 61.260 134.380 61.350 ;
        RECT 133.720 61.120 134.380 61.260 ;
        RECT 131.820 57.970 132.080 58.290 ;
        RECT 132.740 57.970 133.000 58.290 ;
        RECT 133.720 56.220 133.860 61.120 ;
        RECT 134.120 61.030 134.380 61.120 ;
        RECT 136.940 61.010 137.080 63.410 ;
        RECT 136.880 60.690 137.140 61.010 ;
        RECT 137.860 59.310 138.000 63.750 ;
        RECT 137.800 58.990 138.060 59.310 ;
        RECT 138.320 58.290 138.460 65.790 ;
        RECT 139.460 64.915 141.000 65.285 ;
        RECT 141.540 63.730 141.680 67.150 ;
        RECT 144.240 63.750 144.500 64.070 ;
        RECT 138.720 63.410 138.980 63.730 ;
        RECT 141.480 63.410 141.740 63.730 ;
        RECT 138.780 58.630 138.920 63.410 ;
        RECT 144.300 61.350 144.440 63.750 ;
        RECT 144.700 63.410 144.960 63.730 ;
        RECT 141.480 61.030 141.740 61.350 ;
        RECT 144.240 61.030 144.500 61.350 ;
        RECT 139.460 59.475 141.000 59.845 ;
        RECT 138.720 58.310 138.980 58.630 ;
        RECT 136.420 57.970 136.680 58.290 ;
        RECT 138.260 57.970 138.520 58.290 ;
        RECT 136.480 56.220 136.620 57.970 ;
        RECT 139.240 56.530 139.840 56.670 ;
        RECT 139.240 56.220 139.380 56.530 ;
        RECT 37.580 55.850 39.560 55.990 ;
        RECT 39.810 53.440 40.090 56.220 ;
        RECT 42.570 53.990 42.850 56.220 ;
        RECT 42.570 53.710 43.840 53.990 ;
        RECT 39.810 53.160 41.240 53.440 ;
        RECT 37.050 52.610 39.240 52.890 ;
        RECT 34.290 52.110 37.640 52.390 ;
        RECT 31.530 51.510 36.140 51.790 ;
        RECT 35.860 49.790 36.140 51.510 ;
        RECT 33.850 49.740 34.760 49.745 ;
        RECT 28.770 49.460 34.760 49.740 ;
        RECT 33.850 48.895 34.760 49.460 ;
        RECT 35.860 48.910 36.720 49.790 ;
        RECT 37.360 49.770 37.640 52.110 ;
        RECT 38.960 49.785 39.240 52.610 ;
        RECT 37.360 48.910 38.210 49.770 ;
        RECT 38.935 48.975 39.805 49.785 ;
        RECT 40.960 49.735 41.240 53.160 ;
        RECT 43.560 49.815 43.840 53.710 ;
        RECT 40.900 48.985 41.710 49.735 ;
        RECT 43.560 49.060 44.355 49.815 ;
        RECT 38.960 48.960 39.775 48.975 ;
        RECT 30.280 32.060 32.280 46.760 ;
        RECT 33.880 33.205 34.730 48.895 ;
        RECT 30.280 30.060 35.310 32.060 ;
        RECT 30.280 21.060 32.280 30.060 ;
        RECT 35.880 22.725 36.720 48.910 ;
        RECT 30.280 19.060 36.810 21.060 ;
        RECT 30.280 12.860 32.280 19.060 ;
        RECT 37.390 14.080 38.210 48.910 ;
        RECT 38.965 32.585 39.775 48.960 ;
        RECT 40.930 33.705 41.680 48.985 ;
        RECT 43.605 47.785 44.355 49.060 ;
        RECT 45.330 49.240 45.610 56.220 ;
        RECT 48.090 49.760 48.370 56.220 ;
        RECT 45.830 49.240 46.580 49.760 ;
        RECT 45.330 48.960 46.580 49.240 ;
        RECT 43.605 47.035 45.380 47.785 ;
        RECT 42.430 33.860 43.830 38.040 ;
        RECT 44.630 34.585 45.380 47.035 ;
        RECT 45.830 33.980 46.580 48.960 ;
        RECT 47.980 38.135 48.730 49.760 ;
        RECT 49.830 49.240 50.580 49.765 ;
        RECT 50.850 49.240 51.130 56.220 ;
        RECT 53.610 50.340 53.890 56.220 ;
        RECT 56.370 51.990 56.650 56.220 ;
        RECT 52.160 50.060 53.890 50.340 ;
        RECT 54.210 51.710 56.650 51.990 ;
        RECT 52.160 49.760 52.440 50.060 ;
        RECT 54.210 49.765 54.490 51.710 ;
        RECT 59.130 51.490 59.410 56.220 ;
        RECT 56.160 51.210 59.410 51.490 ;
        RECT 56.160 49.785 56.440 51.210 ;
        RECT 61.890 50.940 62.170 56.220 ;
        RECT 58.010 50.660 62.170 50.940 ;
        RECT 58.010 49.815 58.290 50.660 ;
        RECT 64.650 50.390 64.930 56.220 ;
        RECT 60.200 50.110 64.930 50.390 ;
        RECT 51.630 49.735 52.955 49.760 ;
        RECT 49.810 48.960 51.130 49.240 ;
        RECT 51.625 48.985 52.955 49.735 ;
        RECT 49.830 39.635 50.580 48.960 ;
        RECT 52.205 41.185 52.955 48.985 ;
        RECT 53.705 49.010 54.490 49.765 ;
        RECT 55.625 49.035 57.040 49.785 ;
        RECT 53.705 42.885 54.455 49.010 ;
        RECT 53.705 42.135 55.780 42.885 ;
        RECT 52.205 40.435 54.805 41.185 ;
        RECT 49.830 38.885 53.755 39.635 ;
        RECT 47.980 37.385 50.880 38.135 ;
        RECT 42.430 32.760 45.610 33.860 ;
        RECT 45.830 33.340 49.580 33.980 ;
        RECT 50.105 33.935 50.855 37.385 ;
        RECT 45.830 33.335 46.580 33.340 ;
        RECT 50.105 33.280 52.735 33.935 ;
        RECT 50.105 33.235 50.855 33.280 ;
        RECT 38.965 31.775 40.210 32.585 ;
        RECT 30.280 10.860 38.810 12.860 ;
        RECT 30.280 7.050 32.280 10.860 ;
        RECT 39.400 7.335 40.210 31.775 ;
        RECT 42.430 30.460 43.830 32.760 ;
        RECT 53.005 31.035 53.755 38.885 ;
        RECT 42.430 29.360 50.260 30.460 ;
        RECT 50.905 29.785 53.755 31.035 ;
        RECT 42.430 7.060 43.830 29.360 ;
        RECT 47.600 25.460 49.000 29.360 ;
        RECT 52.005 28.285 52.655 28.315 ;
        RECT 54.055 28.285 54.805 40.435 ;
        RECT 50.955 27.535 54.805 28.285 ;
        RECT 50.955 26.685 52.780 27.535 ;
        RECT 50.955 25.950 52.730 26.685 ;
        RECT 47.600 24.710 51.705 25.460 ;
        RECT 47.600 21.880 49.000 24.710 ;
        RECT 55.030 24.260 55.780 42.135 ;
        RECT 51.035 23.510 55.780 24.260 ;
        RECT 51.035 23.495 53.815 23.510 ;
        RECT 51.035 23.125 51.925 23.495 ;
        RECT 53.065 23.125 53.815 23.495 ;
        RECT 55.030 23.485 55.780 23.510 ;
        RECT 51.035 22.375 53.815 23.125 ;
        RECT 51.175 22.365 51.925 22.375 ;
        RECT 47.600 21.130 51.705 21.880 ;
        RECT 47.600 18.300 49.000 21.130 ;
        RECT 56.290 20.640 57.040 49.035 ;
        RECT 51.035 19.890 57.040 20.640 ;
        RECT 51.115 19.535 51.865 19.890 ;
        RECT 52.715 19.885 55.045 19.890 ;
        RECT 54.295 19.535 55.045 19.885 ;
        RECT 51.115 18.785 55.075 19.535 ;
        RECT 51.115 18.755 51.865 18.785 ;
        RECT 47.600 17.550 51.705 18.300 ;
        RECT 47.600 14.720 49.000 17.550 ;
        RECT 55.855 17.080 56.605 17.105 ;
        RECT 57.550 17.080 58.300 49.815 ;
        RECT 60.200 49.685 60.480 50.110 ;
        RECT 61.425 49.780 63.905 49.785 ;
        RECT 67.410 49.780 67.690 56.220 ;
        RECT 70.170 52.190 70.450 56.220 ;
        RECT 72.930 52.790 73.210 56.220 ;
        RECT 75.690 53.440 75.970 56.220 ;
        RECT 78.450 53.940 78.730 56.220 ;
        RECT 78.450 53.660 80.490 53.940 ;
        RECT 75.690 53.160 78.840 53.440 ;
        RECT 72.930 52.510 77.340 52.790 ;
        RECT 70.170 51.910 75.390 52.190 ;
        RECT 75.110 50.585 75.390 51.910 ;
        RECT 77.060 50.630 77.340 52.510 ;
        RECT 59.675 48.935 60.880 49.685 ;
        RECT 61.425 49.500 67.690 49.780 ;
        RECT 75.070 49.735 75.980 50.585 ;
        RECT 77.060 49.760 77.940 50.630 ;
        RECT 78.560 50.610 78.840 53.160 ;
        RECT 80.210 50.625 80.490 53.660 ;
        RECT 81.210 52.740 81.490 56.220 ;
        RECT 81.210 52.460 82.440 52.740 ;
        RECT 78.560 49.760 79.430 50.610 ;
        RECT 80.155 49.815 81.025 50.625 ;
        RECT 82.160 50.575 82.440 52.460 ;
        RECT 82.120 49.825 82.930 50.575 ;
        RECT 83.970 50.140 84.250 56.220 ;
        RECT 86.730 51.940 87.010 56.220 ;
        RECT 86.730 51.660 87.340 51.940 ;
        RECT 84.825 50.140 85.575 50.655 ;
        RECT 87.060 50.600 87.340 51.660 ;
        RECT 89.490 50.600 89.770 56.220 ;
        RECT 92.250 52.490 92.530 56.220 ;
        RECT 95.010 53.140 95.290 56.220 ;
        RECT 91.560 52.210 92.530 52.490 ;
        RECT 93.360 52.860 95.290 53.140 ;
        RECT 91.560 50.605 91.840 52.210 ;
        RECT 83.970 49.860 85.590 50.140 ;
        RECT 61.425 49.035 63.905 49.500 ;
        RECT 50.955 16.330 58.300 17.080 ;
        RECT 50.985 15.955 51.735 16.330 ;
        RECT 55.855 15.955 56.605 16.330 ;
        RECT 50.985 15.205 56.635 15.955 ;
        RECT 50.985 15.175 51.735 15.205 ;
        RECT 47.600 13.970 51.705 14.720 ;
        RECT 47.600 11.140 49.000 13.970 ;
        RECT 58.385 13.520 59.135 13.535 ;
        RECT 60.130 13.520 60.880 48.935 ;
        RECT 50.935 12.770 60.880 13.520 ;
        RECT 50.965 12.385 51.715 12.770 ;
        RECT 58.385 12.385 59.135 12.770 ;
        RECT 50.965 11.635 59.165 12.385 ;
        RECT 50.965 11.605 51.715 11.635 ;
        RECT 47.600 10.390 51.705 11.140 ;
        RECT 47.600 7.060 49.000 10.390 ;
        RECT 61.905 9.920 62.655 9.945 ;
        RECT 63.155 9.920 63.905 49.035 ;
        RECT 64.450 43.250 65.950 45.780 ;
        RECT 64.420 41.750 65.980 43.250 ;
        RECT 64.450 26.300 65.950 41.750 ;
        RECT 71.500 32.900 73.500 47.600 ;
        RECT 75.100 34.045 75.950 49.735 ;
        RECT 71.500 30.900 76.530 32.900 ;
        RECT 64.420 24.800 65.980 26.300 ;
        RECT 64.450 13.450 65.950 24.800 ;
        RECT 71.500 21.900 73.500 30.900 ;
        RECT 77.100 23.565 77.940 49.760 ;
        RECT 71.500 19.900 78.030 21.900 ;
        RECT 71.500 13.700 73.500 19.900 ;
        RECT 78.610 14.920 79.430 49.760 ;
        RECT 80.185 33.425 80.995 49.815 ;
        RECT 82.150 34.545 82.900 49.825 ;
        RECT 84.825 48.625 85.575 49.860 ;
        RECT 84.825 47.875 86.600 48.625 ;
        RECT 83.650 34.700 85.050 38.880 ;
        RECT 85.850 35.425 86.600 47.875 ;
        RECT 87.050 34.820 87.800 50.600 ;
        RECT 89.200 38.975 89.950 50.600 ;
        RECT 91.050 49.810 91.840 50.605 ;
        RECT 93.360 50.600 93.640 52.860 ;
        RECT 97.770 52.590 98.050 56.220 ;
        RECT 95.410 52.310 98.050 52.590 ;
        RECT 95.410 50.605 95.690 52.310 ;
        RECT 100.530 52.090 100.810 56.220 ;
        RECT 97.360 51.810 100.810 52.090 ;
        RECT 97.360 50.625 97.640 51.810 ;
        RECT 103.290 51.570 103.570 56.220 ;
        RECT 99.260 51.290 103.570 51.570 ;
        RECT 99.260 50.655 99.540 51.290 ;
        RECT 106.050 51.110 106.330 56.220 ;
        RECT 92.850 50.575 94.175 50.600 ;
        RECT 92.845 49.825 94.175 50.575 ;
        RECT 93.360 49.810 94.175 49.825 ;
        RECT 91.050 40.475 91.800 49.810 ;
        RECT 93.425 42.025 94.175 49.810 ;
        RECT 94.925 49.810 95.690 50.605 ;
        RECT 96.845 49.875 98.260 50.625 ;
        RECT 97.360 49.860 98.260 49.875 ;
        RECT 94.925 43.725 95.675 49.810 ;
        RECT 94.925 42.975 97.000 43.725 ;
        RECT 93.425 41.275 96.025 42.025 ;
        RECT 91.050 39.725 94.975 40.475 ;
        RECT 89.200 38.225 92.100 38.975 ;
        RECT 83.650 33.600 86.830 34.700 ;
        RECT 87.050 34.180 90.800 34.820 ;
        RECT 91.325 34.775 92.075 38.225 ;
        RECT 87.050 34.175 87.800 34.180 ;
        RECT 91.325 34.120 93.955 34.775 ;
        RECT 91.325 34.075 92.075 34.120 ;
        RECT 80.185 32.615 81.430 33.425 ;
        RECT 64.420 11.950 65.980 13.450 ;
        RECT 64.450 11.000 65.950 11.950 ;
        RECT 71.500 11.700 80.030 13.700 ;
        RECT 50.965 9.170 63.990 9.920 ;
        RECT 50.995 8.785 51.745 9.170 ;
        RECT 61.905 8.785 62.655 9.170 ;
        RECT 50.995 8.035 62.685 8.785 ;
        RECT 50.995 8.005 51.745 8.035 ;
        RECT 71.500 7.890 73.500 11.700 ;
        RECT 80.620 8.175 81.430 32.615 ;
        RECT 83.650 31.300 85.050 33.600 ;
        RECT 94.225 31.875 94.975 39.725 ;
        RECT 83.650 30.200 91.480 31.300 ;
        RECT 92.125 30.625 94.975 31.875 ;
        RECT 83.650 7.900 85.050 30.200 ;
        RECT 88.820 26.300 90.220 30.200 ;
        RECT 93.225 29.125 93.875 29.155 ;
        RECT 95.275 29.125 96.025 41.275 ;
        RECT 92.175 28.375 96.025 29.125 ;
        RECT 92.175 27.525 94.000 28.375 ;
        RECT 92.175 26.790 93.950 27.525 ;
        RECT 88.820 25.550 92.925 26.300 ;
        RECT 88.820 22.720 90.220 25.550 ;
        RECT 96.250 25.100 97.000 42.975 ;
        RECT 92.255 24.350 97.000 25.100 ;
        RECT 92.255 24.335 95.035 24.350 ;
        RECT 92.255 23.965 93.145 24.335 ;
        RECT 94.285 23.965 95.035 24.335 ;
        RECT 96.250 24.325 97.000 24.350 ;
        RECT 92.255 23.215 95.035 23.965 ;
        RECT 92.395 23.205 93.145 23.215 ;
        RECT 88.820 21.970 92.925 22.720 ;
        RECT 88.820 19.140 90.220 21.970 ;
        RECT 97.510 21.480 98.260 49.860 ;
        RECT 92.255 20.730 98.260 21.480 ;
        RECT 98.770 49.860 99.540 50.655 ;
        RECT 101.400 50.830 106.330 51.110 ;
        RECT 101.400 50.525 101.680 50.830 ;
        RECT 92.335 20.375 93.085 20.730 ;
        RECT 93.935 20.725 96.265 20.730 ;
        RECT 95.515 20.375 96.265 20.725 ;
        RECT 92.335 19.625 96.295 20.375 ;
        RECT 92.335 19.595 93.085 19.625 ;
        RECT 88.820 18.390 92.925 19.140 ;
        RECT 88.820 15.560 90.220 18.390 ;
        RECT 97.075 17.920 97.825 17.945 ;
        RECT 98.770 17.920 99.520 49.860 ;
        RECT 100.895 49.775 102.100 50.525 ;
        RECT 102.645 50.460 105.125 50.625 ;
        RECT 108.810 50.460 109.090 56.220 ;
        RECT 111.570 52.890 111.850 56.220 ;
        RECT 114.330 53.340 114.610 56.220 ;
        RECT 117.090 53.340 117.370 56.220 ;
        RECT 119.850 53.390 120.130 56.220 ;
        RECT 114.330 53.060 116.740 53.340 ;
        RECT 117.090 53.060 119.290 53.340 ;
        RECT 119.850 53.110 120.840 53.390 ;
        RECT 111.570 52.610 115.240 52.890 ;
        RECT 114.960 51.985 115.240 52.610 ;
        RECT 114.950 51.135 115.860 51.985 ;
        RECT 116.460 51.440 116.740 53.060 ;
        RECT 116.980 51.440 117.820 52.030 ;
        RECT 119.010 52.010 119.290 53.060 ;
        RECT 120.560 52.025 120.840 53.110 ;
        RECT 116.460 51.160 117.840 51.440 ;
        RECT 102.645 50.180 109.090 50.460 ;
        RECT 102.645 49.875 105.125 50.180 ;
        RECT 92.175 17.170 99.520 17.920 ;
        RECT 92.205 16.795 92.955 17.170 ;
        RECT 97.075 16.795 97.825 17.170 ;
        RECT 92.205 16.045 97.855 16.795 ;
        RECT 92.205 16.015 92.955 16.045 ;
        RECT 88.820 14.810 92.925 15.560 ;
        RECT 88.820 11.980 90.220 14.810 ;
        RECT 99.605 14.360 100.355 14.375 ;
        RECT 101.350 14.360 102.100 49.775 ;
        RECT 92.155 13.610 102.100 14.360 ;
        RECT 92.185 13.225 92.935 13.610 ;
        RECT 99.605 13.225 100.355 13.610 ;
        RECT 92.185 12.475 100.385 13.225 ;
        RECT 92.185 12.445 92.935 12.475 ;
        RECT 88.820 11.230 92.925 11.980 ;
        RECT 88.820 7.900 90.220 11.230 ;
        RECT 103.125 10.760 103.875 10.785 ;
        RECT 104.375 10.760 105.125 49.875 ;
        RECT 105.700 43.300 107.200 45.830 ;
        RECT 105.670 41.800 107.230 43.300 ;
        RECT 105.700 26.350 107.200 41.800 ;
        RECT 111.380 34.300 113.380 49.000 ;
        RECT 114.980 35.445 115.830 51.135 ;
        RECT 111.380 32.300 116.410 34.300 ;
        RECT 105.670 24.850 107.230 26.350 ;
        RECT 105.700 13.500 107.200 24.850 ;
        RECT 111.380 23.300 113.380 32.300 ;
        RECT 116.980 24.965 117.820 51.160 ;
        RECT 111.380 21.300 117.910 23.300 ;
        RECT 111.380 15.100 113.380 21.300 ;
        RECT 118.490 16.320 119.310 52.010 ;
        RECT 120.035 51.215 120.905 52.025 ;
        RECT 122.610 51.975 122.890 56.220 ;
        RECT 125.370 52.055 125.650 56.220 ;
        RECT 128.130 52.590 128.410 56.220 ;
        RECT 130.890 52.590 131.170 56.220 ;
        RECT 133.650 53.040 133.930 56.220 ;
        RECT 136.410 53.440 136.690 56.220 ;
        RECT 139.170 53.990 139.450 56.220 ;
        RECT 139.700 55.990 139.840 56.530 ;
        RECT 141.540 55.990 141.680 61.030 ;
        RECT 142.400 58.200 142.660 58.290 ;
        RECT 142.000 58.060 142.660 58.200 ;
        RECT 142.000 56.220 142.140 58.060 ;
        RECT 142.400 57.970 142.660 58.060 ;
        RECT 144.760 56.220 144.900 63.410 ;
        RECT 145.680 61.350 145.820 68.170 ;
        RECT 146.080 63.410 146.340 63.730 ;
        RECT 145.620 61.030 145.880 61.350 ;
        RECT 146.140 58.290 146.280 63.410 ;
        RECT 146.600 58.290 146.740 69.190 ;
        RECT 156.250 67.635 157.790 68.005 ;
        RECT 156.250 62.195 157.790 62.565 ;
        RECT 147.460 61.030 147.720 61.350 ;
        RECT 146.080 57.970 146.340 58.290 ;
        RECT 146.540 57.970 146.800 58.290 ;
        RECT 147.520 56.220 147.660 61.030 ;
        RECT 150.220 57.970 150.480 58.290 ;
        RECT 150.280 56.220 150.420 57.970 ;
        RECT 156.250 56.755 157.790 57.125 ;
        RECT 139.700 55.850 141.680 55.990 ;
        RECT 122.000 51.225 122.890 51.975 ;
        RECT 120.065 34.825 120.875 51.215 ;
        RECT 122.030 51.210 122.890 51.225 ;
        RECT 124.705 51.260 125.650 52.055 ;
        RECT 127.410 52.310 128.410 52.590 ;
        RECT 129.560 52.310 131.170 52.590 ;
        RECT 131.410 52.760 133.930 53.040 ;
        RECT 134.610 53.160 136.690 53.440 ;
        RECT 138.110 53.710 139.450 53.990 ;
        RECT 127.410 52.000 127.690 52.310 ;
        RECT 129.560 52.000 129.840 52.310 ;
        RECT 131.410 52.005 131.690 52.760 ;
        RECT 134.610 52.590 134.890 53.160 ;
        RECT 138.110 52.990 138.390 53.710 ;
        RECT 141.930 53.490 142.210 56.220 ;
        RECT 122.030 35.945 122.780 51.210 ;
        RECT 124.705 50.025 125.455 51.260 ;
        RECT 126.930 51.210 127.690 52.000 ;
        RECT 124.705 49.275 126.480 50.025 ;
        RECT 123.530 36.100 124.930 40.280 ;
        RECT 125.730 36.825 126.480 49.275 ;
        RECT 126.930 36.220 127.680 51.210 ;
        RECT 129.080 51.160 129.840 52.000 ;
        RECT 130.930 51.260 131.690 52.005 ;
        RECT 133.160 52.310 134.890 52.590 ;
        RECT 135.210 52.710 138.390 52.990 ;
        RECT 138.910 53.210 142.210 53.490 ;
        RECT 133.160 52.000 133.440 52.310 ;
        RECT 135.210 52.005 135.490 52.710 ;
        RECT 138.910 52.490 139.190 53.210 ;
        RECT 144.690 52.990 144.970 56.220 ;
        RECT 137.210 52.210 139.190 52.490 ;
        RECT 139.710 52.710 144.970 52.990 ;
        RECT 137.210 52.025 137.490 52.210 ;
        RECT 132.730 51.975 134.055 52.000 ;
        RECT 129.080 40.375 129.830 51.160 ;
        RECT 130.930 41.875 131.680 51.260 ;
        RECT 132.725 51.225 134.055 51.975 ;
        RECT 133.305 43.425 134.055 51.225 ;
        RECT 134.805 45.125 135.555 52.005 ;
        RECT 136.725 51.275 138.140 52.025 ;
        RECT 134.805 44.375 136.880 45.125 ;
        RECT 133.305 42.675 135.905 43.425 ;
        RECT 130.930 41.125 134.855 41.875 ;
        RECT 129.080 39.625 131.980 40.375 ;
        RECT 123.530 35.000 126.710 36.100 ;
        RECT 126.930 35.580 130.680 36.220 ;
        RECT 131.205 36.175 131.955 39.625 ;
        RECT 126.930 35.575 127.680 35.580 ;
        RECT 131.205 35.520 133.835 36.175 ;
        RECT 131.205 35.475 131.955 35.520 ;
        RECT 120.065 34.015 121.310 34.825 ;
        RECT 105.670 12.000 107.230 13.500 ;
        RECT 111.380 13.100 119.910 15.100 ;
        RECT 105.700 11.050 107.200 12.000 ;
        RECT 92.185 10.010 105.210 10.760 ;
        RECT 92.215 9.625 92.965 10.010 ;
        RECT 103.125 9.625 103.875 10.010 ;
        RECT 92.215 8.875 103.905 9.625 ;
        RECT 111.380 9.290 113.380 13.100 ;
        RECT 120.500 9.575 121.310 34.015 ;
        RECT 123.530 32.700 124.930 35.000 ;
        RECT 134.105 33.275 134.855 41.125 ;
        RECT 123.530 31.600 131.360 32.700 ;
        RECT 132.005 32.025 134.855 33.275 ;
        RECT 123.530 9.300 124.930 31.600 ;
        RECT 128.700 27.700 130.100 31.600 ;
        RECT 133.105 30.525 133.755 30.555 ;
        RECT 135.155 30.525 135.905 42.675 ;
        RECT 132.055 29.775 135.905 30.525 ;
        RECT 132.055 28.925 133.880 29.775 ;
        RECT 132.055 28.190 133.830 28.925 ;
        RECT 128.700 26.950 132.805 27.700 ;
        RECT 128.700 24.120 130.100 26.950 ;
        RECT 136.130 26.500 136.880 44.375 ;
        RECT 132.135 25.750 136.880 26.500 ;
        RECT 132.135 25.735 134.915 25.750 ;
        RECT 132.135 25.365 133.025 25.735 ;
        RECT 134.165 25.365 134.915 25.735 ;
        RECT 136.130 25.725 136.880 25.750 ;
        RECT 132.135 24.615 134.915 25.365 ;
        RECT 132.275 24.605 133.025 24.615 ;
        RECT 128.700 23.370 132.805 24.120 ;
        RECT 128.700 20.540 130.100 23.370 ;
        RECT 137.390 22.880 138.140 51.275 ;
        RECT 132.135 22.130 138.140 22.880 ;
        RECT 138.650 51.940 139.400 52.055 ;
        RECT 139.710 51.940 139.990 52.710 ;
        RECT 147.450 52.490 147.730 56.220 ;
        RECT 138.650 51.660 139.990 51.940 ;
        RECT 141.310 52.210 147.730 52.490 ;
        RECT 141.310 51.925 141.590 52.210 ;
        RECT 132.215 21.775 132.965 22.130 ;
        RECT 133.815 22.125 136.145 22.130 ;
        RECT 135.395 21.775 136.145 22.125 ;
        RECT 132.215 21.025 136.175 21.775 ;
        RECT 132.215 20.995 132.965 21.025 ;
        RECT 128.700 19.790 132.805 20.540 ;
        RECT 128.700 16.960 130.100 19.790 ;
        RECT 136.955 19.320 137.705 19.345 ;
        RECT 138.650 19.320 139.400 51.660 ;
        RECT 140.775 51.175 141.980 51.925 ;
        RECT 142.525 51.490 145.005 52.025 ;
        RECT 150.210 51.490 150.490 56.220 ;
        RECT 142.525 51.275 150.490 51.490 ;
        RECT 142.610 51.210 150.490 51.275 ;
        RECT 132.055 18.570 139.400 19.320 ;
        RECT 132.085 18.195 132.835 18.570 ;
        RECT 136.955 18.195 137.705 18.570 ;
        RECT 132.085 17.445 137.735 18.195 ;
        RECT 132.085 17.415 132.835 17.445 ;
        RECT 128.700 16.210 132.805 16.960 ;
        RECT 128.700 13.380 130.100 16.210 ;
        RECT 139.485 15.760 140.235 15.775 ;
        RECT 141.230 15.760 141.980 51.175 ;
        RECT 132.035 15.010 141.980 15.760 ;
        RECT 132.065 14.625 132.815 15.010 ;
        RECT 139.485 14.625 140.235 15.010 ;
        RECT 132.065 13.875 140.265 14.625 ;
        RECT 132.065 13.845 132.815 13.875 ;
        RECT 128.700 12.630 132.805 13.380 ;
        RECT 128.700 9.300 130.100 12.630 ;
        RECT 143.005 12.160 143.755 12.185 ;
        RECT 144.255 12.160 145.005 51.210 ;
        RECT 145.650 43.250 147.150 45.780 ;
        RECT 145.620 41.750 147.180 43.250 ;
        RECT 145.650 26.300 147.150 41.750 ;
        RECT 145.620 24.800 147.180 26.300 ;
        RECT 145.650 13.450 147.150 24.800 ;
        RECT 132.065 11.410 145.090 12.160 ;
        RECT 145.620 11.950 147.180 13.450 ;
        RECT 132.095 11.025 132.845 11.410 ;
        RECT 143.005 11.025 143.755 11.410 ;
        RECT 132.095 10.275 143.785 11.025 ;
        RECT 145.650 11.000 147.150 11.950 ;
        RECT 132.095 10.245 132.845 10.275 ;
        RECT 123.530 9.290 130.100 9.300 ;
        RECT 142.830 9.290 144.230 9.880 ;
        RECT 92.215 8.845 92.965 8.875 ;
        RECT 83.650 7.890 90.220 7.900 ;
        RECT 102.950 7.890 104.350 8.480 ;
        RECT 42.430 7.050 49.000 7.060 ;
        RECT 61.730 7.050 63.130 7.640 ;
        RECT 30.280 5.050 63.180 7.050 ;
        RECT 71.500 5.890 104.400 7.890 ;
        RECT 111.380 7.290 144.280 9.290 ;
        RECT 127.830 6.595 129.870 6.615 ;
        RECT 87.465 5.515 89.740 5.535 ;
        RECT 44.415 4.505 46.585 4.525 ;
        RECT 41.610 2.285 46.610 4.505 ;
        RECT 84.360 3.190 89.765 5.515 ;
        RECT 124.125 4.505 129.895 6.595 ;
        RECT 127.830 4.485 129.870 4.505 ;
        RECT 87.465 3.170 89.740 3.190 ;
        RECT 44.415 2.265 46.585 2.285 ;
      LAYER met3 ;
        RECT 81.230 223.890 81.610 224.210 ;
        RECT 84.910 223.890 85.290 224.210 ;
        RECT 88.590 223.890 88.970 224.210 ;
        RECT 78.435 220.900 78.765 220.915 ;
        RECT 79.190 220.900 79.510 220.940 ;
        RECT 78.435 220.600 79.510 220.900 ;
        RECT 78.435 220.585 78.765 220.600 ;
        RECT 79.190 220.560 79.510 220.600 ;
        RECT 26.935 217.950 27.265 217.965 ;
        RECT 81.270 217.950 81.570 223.890 ;
        RECT 26.935 217.650 81.570 217.950 ;
        RECT 26.935 217.635 27.265 217.650 ;
        RECT 34.285 217.250 34.615 217.265 ;
        RECT 84.950 217.250 85.250 223.890 ;
        RECT 85.785 220.200 86.115 220.215 ;
        RECT 86.590 220.200 86.910 220.240 ;
        RECT 85.785 219.900 86.910 220.200 ;
        RECT 85.785 219.885 86.115 219.900 ;
        RECT 86.590 219.860 86.910 219.900 ;
        RECT 34.285 216.950 85.250 217.250 ;
        RECT 34.285 216.935 34.615 216.950 ;
        RECT 41.635 216.550 41.965 216.565 ;
        RECT 88.630 216.550 88.930 223.890 ;
        RECT 93.135 219.550 93.465 219.565 ;
        RECT 94.040 219.550 94.360 219.590 ;
        RECT 93.135 219.250 94.360 219.550 ;
        RECT 93.135 219.235 93.465 219.250 ;
        RECT 94.040 219.210 94.360 219.250 ;
        RECT 100.535 218.850 100.865 218.865 ;
        RECT 101.490 218.850 101.810 218.890 ;
        RECT 100.535 218.550 101.810 218.850 ;
        RECT 100.535 218.535 100.865 218.550 ;
        RECT 101.490 218.510 101.810 218.550 ;
        RECT 107.885 218.150 108.215 218.165 ;
        RECT 108.690 218.150 109.010 218.190 ;
        RECT 107.885 217.850 109.010 218.150 ;
        RECT 107.885 217.835 108.215 217.850 ;
        RECT 108.690 217.810 109.010 217.850 ;
        RECT 115.235 217.400 115.565 217.415 ;
        RECT 116.040 217.400 116.360 217.440 ;
        RECT 115.235 217.100 116.360 217.400 ;
        RECT 115.235 217.085 115.565 217.100 ;
        RECT 116.040 217.060 116.360 217.100 ;
        RECT 41.635 216.250 88.930 216.550 ;
        RECT 122.585 216.750 122.915 216.765 ;
        RECT 123.390 216.750 123.710 216.790 ;
        RECT 122.585 216.450 123.710 216.750 ;
        RECT 122.585 216.435 122.915 216.450 ;
        RECT 123.390 216.410 123.710 216.450 ;
        RECT 41.635 216.235 41.965 216.250 ;
        RECT 129.935 216.100 130.265 216.115 ;
        RECT 130.840 216.100 131.160 216.140 ;
        RECT 48.960 215.540 49.340 215.860 ;
        RECT 49.000 214.915 49.300 215.540 ;
        RECT 56.340 215.510 56.660 215.890 ;
        RECT 63.690 215.510 64.010 215.890 ;
        RECT 129.935 215.800 131.160 216.100 ;
        RECT 129.935 215.785 130.265 215.800 ;
        RECT 130.840 215.760 131.160 215.800 ;
        RECT 56.350 214.915 56.650 215.510 ;
        RECT 63.700 214.965 64.000 215.510 ;
        RECT 137.275 215.460 137.605 215.475 ;
        RECT 138.560 215.460 138.880 215.500 ;
        RECT 137.275 215.160 138.880 215.460 ;
        RECT 137.275 215.145 137.605 215.160 ;
        RECT 138.560 215.120 138.880 215.160 ;
        RECT 48.985 214.585 49.315 214.915 ;
        RECT 56.335 214.585 56.665 214.915 ;
        RECT 63.685 214.635 64.015 214.965 ;
        RECT 71.050 214.915 71.350 214.950 ;
        RECT 71.035 214.900 71.365 214.915 ;
        RECT 71.940 214.900 72.260 214.940 ;
        RECT 71.035 214.600 72.260 214.900 ;
        RECT 71.035 214.585 71.365 214.600 ;
        RECT 71.940 214.560 72.260 214.600 ;
        RECT 144.665 214.790 144.995 214.805 ;
        RECT 145.870 214.790 146.190 214.830 ;
        RECT 144.665 214.490 146.190 214.790 ;
        RECT 144.665 214.475 144.995 214.490 ;
        RECT 145.870 214.450 146.190 214.490 ;
        RECT 152.545 214.140 152.875 214.155 ;
        RECT 153.500 214.140 153.820 214.180 ;
        RECT 152.545 213.840 153.820 214.140 ;
        RECT 152.545 213.825 152.875 213.840 ;
        RECT 153.500 213.800 153.820 213.840 ;
        RECT 55.490 209.095 57.070 209.425 ;
        RECT 89.070 209.095 90.650 209.425 ;
        RECT 122.650 209.095 124.230 209.425 ;
        RECT 156.230 209.095 157.810 209.425 ;
        RECT 108.325 208.390 108.655 208.405 ;
        RECT 115.225 208.390 115.555 208.405 ;
        RECT 108.325 208.090 115.555 208.390 ;
        RECT 108.325 208.075 108.655 208.090 ;
        RECT 115.225 208.075 115.555 208.090 ;
        RECT 38.700 206.375 40.280 206.705 ;
        RECT 72.280 206.375 73.860 206.705 ;
        RECT 105.860 206.375 107.440 206.705 ;
        RECT 139.440 206.375 141.020 206.705 ;
        RECT 55.490 203.655 57.070 203.985 ;
        RECT 89.070 203.655 90.650 203.985 ;
        RECT 122.650 203.655 124.230 203.985 ;
        RECT 156.230 203.655 157.810 203.985 ;
        RECT 38.700 200.935 40.280 201.265 ;
        RECT 72.280 200.935 73.860 201.265 ;
        RECT 105.860 200.935 107.440 201.265 ;
        RECT 139.440 200.935 141.020 201.265 ;
        RECT 136.385 200.230 136.715 200.245 ;
        RECT 137.765 200.230 138.095 200.245 ;
        RECT 136.385 199.930 138.095 200.230 ;
        RECT 136.385 199.915 136.715 199.930 ;
        RECT 137.765 199.915 138.095 199.930 ;
        RECT 131.325 199.550 131.655 199.565 ;
        RECT 140.065 199.550 140.395 199.565 ;
        RECT 131.325 199.250 140.395 199.550 ;
        RECT 131.325 199.235 131.655 199.250 ;
        RECT 140.065 199.235 140.395 199.250 ;
        RECT 55.490 198.215 57.070 198.545 ;
        RECT 89.070 198.215 90.650 198.545 ;
        RECT 122.650 198.215 124.230 198.545 ;
        RECT 156.230 198.215 157.810 198.545 ;
        RECT 38.700 195.495 40.280 195.825 ;
        RECT 72.280 195.495 73.860 195.825 ;
        RECT 105.860 195.495 107.440 195.825 ;
        RECT 139.440 195.495 141.020 195.825 ;
        RECT 55.490 192.775 57.070 193.105 ;
        RECT 89.070 192.775 90.650 193.105 ;
        RECT 122.650 192.775 124.230 193.105 ;
        RECT 156.230 192.775 157.810 193.105 ;
        RECT 108.785 191.400 109.115 191.405 ;
        RECT 108.530 191.390 109.115 191.400 ;
        RECT 108.530 191.090 109.340 191.390 ;
        RECT 108.530 191.080 109.115 191.090 ;
        RECT 108.785 191.075 109.115 191.080 ;
        RECT 38.700 190.055 40.280 190.385 ;
        RECT 72.280 190.055 73.860 190.385 ;
        RECT 105.860 190.055 107.440 190.385 ;
        RECT 139.440 190.055 141.020 190.385 ;
        RECT 111.085 187.990 111.415 188.005 ;
        RECT 112.465 187.990 112.795 188.005 ;
        RECT 111.085 187.690 112.795 187.990 ;
        RECT 111.085 187.675 111.415 187.690 ;
        RECT 112.465 187.675 112.795 187.690 ;
        RECT 55.490 187.335 57.070 187.665 ;
        RECT 89.070 187.335 90.650 187.665 ;
        RECT 122.650 187.335 124.230 187.665 ;
        RECT 156.230 187.335 157.810 187.665 ;
        RECT 90.845 186.630 91.175 186.645 ;
        RECT 109.705 186.630 110.035 186.645 ;
        RECT 90.845 186.330 110.035 186.630 ;
        RECT 90.845 186.315 91.175 186.330 ;
        RECT 109.705 186.315 110.035 186.330 ;
        RECT 49.445 185.950 49.775 185.965 ;
        RECT 53.585 185.950 53.915 185.965 ;
        RECT 96.825 185.950 97.155 185.965 ;
        RECT 103.265 185.950 103.595 185.965 ;
        RECT 49.445 185.650 103.595 185.950 ;
        RECT 49.445 185.635 49.775 185.650 ;
        RECT 53.585 185.635 53.915 185.650 ;
        RECT 96.825 185.635 97.155 185.650 ;
        RECT 103.265 185.635 103.595 185.650 ;
        RECT 38.700 184.615 40.280 184.945 ;
        RECT 72.280 184.615 73.860 184.945 ;
        RECT 105.860 184.615 107.440 184.945 ;
        RECT 139.440 184.615 141.020 184.945 ;
        RECT 103.265 183.920 103.595 183.925 ;
        RECT 103.010 183.910 103.595 183.920 ;
        RECT 107.865 183.910 108.195 183.925 ;
        RECT 102.810 183.610 108.195 183.910 ;
        RECT 103.010 183.600 103.595 183.610 ;
        RECT 103.265 183.595 103.595 183.600 ;
        RECT 107.865 183.595 108.195 183.610 ;
        RECT 108.530 183.910 108.910 183.920 ;
        RECT 144.205 183.910 144.535 183.925 ;
        RECT 108.530 183.610 144.535 183.910 ;
        RECT 108.530 183.600 108.910 183.610 ;
        RECT 144.205 183.595 144.535 183.610 ;
        RECT 109.705 182.560 110.035 182.565 ;
        RECT 109.450 182.550 110.035 182.560 ;
        RECT 109.450 182.250 110.260 182.550 ;
        RECT 109.450 182.240 110.035 182.250 ;
        RECT 109.705 182.235 110.035 182.240 ;
        RECT 55.490 181.895 57.070 182.225 ;
        RECT 89.070 181.895 90.650 182.225 ;
        RECT 122.650 181.895 124.230 182.225 ;
        RECT 156.230 181.895 157.810 182.225 ;
        RECT 38.700 179.175 40.280 179.505 ;
        RECT 72.280 179.175 73.860 179.505 ;
        RECT 105.860 179.175 107.440 179.505 ;
        RECT 139.440 179.175 141.020 179.505 ;
        RECT 55.490 176.455 57.070 176.785 ;
        RECT 89.070 176.455 90.650 176.785 ;
        RECT 122.650 176.455 124.230 176.785 ;
        RECT 156.230 176.455 157.810 176.785 ;
        RECT 38.700 173.735 40.280 174.065 ;
        RECT 72.280 173.735 73.860 174.065 ;
        RECT 105.860 173.735 107.440 174.065 ;
        RECT 139.440 173.735 141.020 174.065 ;
        RECT 38.865 172.350 39.195 172.365 ;
        RECT 44.845 172.350 45.175 172.365 ;
        RECT 38.865 172.050 45.175 172.350 ;
        RECT 38.865 172.035 39.195 172.050 ;
        RECT 44.845 172.035 45.175 172.050 ;
        RECT 82.565 172.350 82.895 172.365 ;
        RECT 86.245 172.350 86.575 172.365 ;
        RECT 109.450 172.350 109.830 172.360 ;
        RECT 82.565 172.050 109.830 172.350 ;
        RECT 82.565 172.035 82.895 172.050 ;
        RECT 86.245 172.035 86.575 172.050 ;
        RECT 109.450 172.040 109.830 172.050 ;
        RECT 55.490 171.015 57.070 171.345 ;
        RECT 89.070 171.015 90.650 171.345 ;
        RECT 122.650 171.015 124.230 171.345 ;
        RECT 156.230 171.015 157.810 171.345 ;
        RECT 53.125 170.990 53.455 171.005 ;
        RECT 53.125 170.675 53.670 170.990 ;
        RECT 50.825 170.310 51.155 170.325 ;
        RECT 53.370 170.310 53.670 170.675 ;
        RECT 57.970 170.690 82.190 170.990 ;
        RECT 57.970 170.310 58.270 170.690 ;
        RECT 50.825 170.010 58.270 170.310 ;
        RECT 58.645 170.310 58.975 170.325 ;
        RECT 71.525 170.310 71.855 170.325 ;
        RECT 81.890 170.310 82.190 170.690 ;
        RECT 96.825 170.310 97.155 170.325 ;
        RECT 58.645 170.010 72.070 170.310 ;
        RECT 81.890 170.010 97.155 170.310 ;
        RECT 50.825 169.995 51.155 170.010 ;
        RECT 58.645 169.995 58.975 170.010 ;
        RECT 71.525 169.995 72.070 170.010 ;
        RECT 96.825 169.995 97.155 170.010 ;
        RECT 71.770 169.630 72.070 169.995 ;
        RECT 99.125 169.630 99.455 169.645 ;
        RECT 71.770 169.330 99.455 169.630 ;
        RECT 99.125 169.315 99.455 169.330 ;
        RECT 38.700 168.295 40.280 168.625 ;
        RECT 72.280 168.295 73.860 168.625 ;
        RECT 105.860 168.295 107.440 168.625 ;
        RECT 139.440 168.295 141.020 168.625 ;
        RECT 55.490 165.575 57.070 165.905 ;
        RECT 89.070 165.575 90.650 165.905 ;
        RECT 122.650 165.575 124.230 165.905 ;
        RECT 156.230 165.575 157.810 165.905 ;
        RECT 75.410 164.870 75.790 164.880 ;
        RECT 76.125 164.870 76.455 164.885 ;
        RECT 100.965 164.870 101.295 164.885 ;
        RECT 110.625 164.870 110.955 164.885 ;
        RECT 75.410 164.570 110.955 164.870 ;
        RECT 75.410 164.560 75.790 164.570 ;
        RECT 76.125 164.555 76.455 164.570 ;
        RECT 100.965 164.555 101.295 164.570 ;
        RECT 110.625 164.555 110.955 164.570 ;
        RECT 45.970 164.190 46.350 164.200 ;
        RECT 46.685 164.190 47.015 164.205 ;
        RECT 45.970 163.890 47.015 164.190 ;
        RECT 45.970 163.880 46.350 163.890 ;
        RECT 46.685 163.875 47.015 163.890 ;
        RECT 75.205 164.190 75.535 164.205 ;
        RECT 76.330 164.190 76.710 164.200 ;
        RECT 108.785 164.190 109.115 164.205 ;
        RECT 75.205 163.890 109.115 164.190 ;
        RECT 75.205 163.875 75.535 163.890 ;
        RECT 76.330 163.880 76.710 163.890 ;
        RECT 108.785 163.875 109.115 163.890 ;
        RECT 38.700 162.855 40.280 163.185 ;
        RECT 72.280 162.855 73.860 163.185 ;
        RECT 105.860 162.855 107.440 163.185 ;
        RECT 139.440 162.855 141.020 163.185 ;
        RECT 87.165 161.470 87.495 161.485 ;
        RECT 100.965 161.470 101.295 161.485 ;
        RECT 87.165 161.170 101.295 161.470 ;
        RECT 87.165 161.155 87.495 161.170 ;
        RECT 100.965 161.155 101.295 161.170 ;
        RECT 55.490 160.135 57.070 160.465 ;
        RECT 89.070 160.135 90.650 160.465 ;
        RECT 122.650 160.135 124.230 160.465 ;
        RECT 156.230 160.135 157.810 160.465 ;
        RECT 68.305 159.430 68.635 159.445 ;
        RECT 70.145 159.430 70.475 159.445 ;
        RECT 105.105 159.430 105.435 159.445 ;
        RECT 68.305 159.130 105.435 159.430 ;
        RECT 68.305 159.115 68.635 159.130 ;
        RECT 70.145 159.115 70.475 159.130 ;
        RECT 105.105 159.115 105.435 159.130 ;
        RECT 38.700 157.415 40.280 157.745 ;
        RECT 72.280 157.415 73.860 157.745 ;
        RECT 105.860 157.415 107.440 157.745 ;
        RECT 139.440 157.415 141.020 157.745 ;
        RECT 68.305 156.710 68.635 156.725 ;
        RECT 79.805 156.710 80.135 156.725 ;
        RECT 111.085 156.710 111.415 156.725 ;
        RECT 68.305 156.410 111.415 156.710 ;
        RECT 68.305 156.395 68.635 156.410 ;
        RECT 79.805 156.395 80.135 156.410 ;
        RECT 111.085 156.395 111.415 156.410 ;
        RECT 55.490 154.695 57.070 155.025 ;
        RECT 89.070 154.695 90.650 155.025 ;
        RECT 122.650 154.695 124.230 155.025 ;
        RECT 156.230 154.695 157.810 155.025 ;
        RECT 98.205 153.310 98.535 153.325 ;
        RECT 100.250 153.310 100.630 153.320 ;
        RECT 98.205 153.010 100.630 153.310 ;
        RECT 98.205 152.995 98.535 153.010 ;
        RECT 100.250 153.000 100.630 153.010 ;
        RECT 38.700 151.975 40.280 152.305 ;
        RECT 72.280 151.975 73.860 152.305 ;
        RECT 105.860 151.975 107.440 152.305 ;
        RECT 139.440 151.975 141.020 152.305 ;
        RECT 82.770 151.270 83.150 151.280 ;
        RECT 90.845 151.270 91.175 151.285 ;
        RECT 82.770 150.970 91.175 151.270 ;
        RECT 82.770 150.960 83.150 150.970 ;
        RECT 90.845 150.955 91.175 150.970 ;
        RECT 103.010 150.590 103.390 150.600 ;
        RECT 103.725 150.590 104.055 150.605 ;
        RECT 106.025 150.590 106.355 150.605 ;
        RECT 103.010 150.290 106.355 150.590 ;
        RECT 103.010 150.280 103.390 150.290 ;
        RECT 103.725 150.275 104.055 150.290 ;
        RECT 106.025 150.275 106.355 150.290 ;
        RECT 107.865 150.590 108.195 150.605 ;
        RECT 108.530 150.590 108.910 150.600 ;
        RECT 107.865 150.290 108.910 150.590 ;
        RECT 107.865 150.275 108.195 150.290 ;
        RECT 108.530 150.280 108.910 150.290 ;
        RECT 55.490 149.255 57.070 149.585 ;
        RECT 89.070 149.255 90.650 149.585 ;
        RECT 122.650 149.255 124.230 149.585 ;
        RECT 156.230 149.255 157.810 149.585 ;
        RECT 38.700 146.535 40.280 146.865 ;
        RECT 72.280 146.535 73.860 146.865 ;
        RECT 105.860 146.535 107.440 146.865 ;
        RECT 139.440 146.535 141.020 146.865 ;
        RECT 108.325 145.830 108.655 145.845 ;
        RECT 109.450 145.830 109.830 145.840 ;
        RECT 108.325 145.530 109.830 145.830 ;
        RECT 108.325 145.515 108.655 145.530 ;
        RECT 109.450 145.520 109.830 145.530 ;
        RECT 95.445 145.150 95.775 145.165 ;
        RECT 100.505 145.150 100.835 145.165 ;
        RECT 95.445 144.850 100.835 145.150 ;
        RECT 95.445 144.835 95.775 144.850 ;
        RECT 100.505 144.835 100.835 144.850 ;
        RECT 55.490 143.815 57.070 144.145 ;
        RECT 89.070 143.815 90.650 144.145 ;
        RECT 122.650 143.815 124.230 144.145 ;
        RECT 156.230 143.815 157.810 144.145 ;
        RECT 70.145 143.790 70.475 143.805 ;
        RECT 75.410 143.790 75.790 143.800 ;
        RECT 70.145 143.490 75.790 143.790 ;
        RECT 70.145 143.475 70.475 143.490 ;
        RECT 75.410 143.480 75.790 143.490 ;
        RECT 38.700 141.095 40.280 141.425 ;
        RECT 72.280 141.095 73.860 141.425 ;
        RECT 105.860 141.095 107.440 141.425 ;
        RECT 139.440 141.095 141.020 141.425 ;
        RECT 55.490 138.375 57.070 138.705 ;
        RECT 89.070 138.375 90.650 138.705 ;
        RECT 122.650 138.375 124.230 138.705 ;
        RECT 156.230 138.375 157.810 138.705 ;
        RECT 67.385 137.670 67.715 137.685 ;
        RECT 82.770 137.670 83.150 137.680 ;
        RECT 67.385 137.370 83.150 137.670 ;
        RECT 67.385 137.355 67.715 137.370 ;
        RECT 82.770 137.360 83.150 137.370 ;
        RECT 99.585 137.670 99.915 137.685 ;
        RECT 100.250 137.670 100.630 137.680 ;
        RECT 99.585 137.370 100.630 137.670 ;
        RECT 99.585 137.355 99.915 137.370 ;
        RECT 100.250 137.360 100.630 137.370 ;
        RECT 38.700 135.655 40.280 135.985 ;
        RECT 72.280 135.655 73.860 135.985 ;
        RECT 105.860 135.655 107.440 135.985 ;
        RECT 139.440 135.655 141.020 135.985 ;
        RECT 55.490 132.935 57.070 133.265 ;
        RECT 89.070 132.935 90.650 133.265 ;
        RECT 122.650 132.935 124.230 133.265 ;
        RECT 156.230 132.935 157.810 133.265 ;
        RECT 128.565 132.910 128.895 132.925 ;
        RECT 130.405 132.910 130.735 132.925 ;
        RECT 128.565 132.610 130.735 132.910 ;
        RECT 128.565 132.595 128.895 132.610 ;
        RECT 130.405 132.595 130.735 132.610 ;
        RECT 28.285 132.230 28.615 132.245 ;
        RECT 45.970 132.230 46.350 132.240 ;
        RECT 28.285 131.930 46.350 132.230 ;
        RECT 28.285 131.915 28.615 131.930 ;
        RECT 45.970 131.920 46.350 131.930 ;
        RECT 38.700 130.215 40.280 130.545 ;
        RECT 72.280 130.215 73.860 130.545 ;
        RECT 105.860 130.215 107.440 130.545 ;
        RECT 139.440 130.215 141.020 130.545 ;
        RECT 76.125 130.200 76.455 130.205 ;
        RECT 76.125 130.190 76.710 130.200 ;
        RECT 76.125 129.890 76.910 130.190 ;
        RECT 76.125 129.880 76.710 129.890 ;
        RECT 76.125 129.875 76.455 129.880 ;
        RECT 55.490 127.495 57.070 127.825 ;
        RECT 89.070 127.495 90.650 127.825 ;
        RECT 122.650 127.495 124.230 127.825 ;
        RECT 156.230 127.495 157.810 127.825 ;
        RECT 38.700 124.775 40.280 125.105 ;
        RECT 72.280 124.775 73.860 125.105 ;
        RECT 105.860 124.775 107.440 125.105 ;
        RECT 139.440 124.775 141.020 125.105 ;
        RECT 82.770 124.070 83.150 124.080 ;
        RECT 88.545 124.070 88.875 124.085 ;
        RECT 82.770 123.770 88.875 124.070 ;
        RECT 82.770 123.760 83.150 123.770 ;
        RECT 88.545 123.755 88.875 123.770 ;
        RECT 55.490 122.055 57.070 122.385 ;
        RECT 89.070 122.055 90.650 122.385 ;
        RECT 122.650 122.055 124.230 122.385 ;
        RECT 156.230 122.055 157.810 122.385 ;
        RECT 38.700 119.335 40.280 119.665 ;
        RECT 72.280 119.335 73.860 119.665 ;
        RECT 105.860 119.335 107.440 119.665 ;
        RECT 139.440 119.335 141.020 119.665 ;
        RECT 55.490 116.615 57.070 116.945 ;
        RECT 89.070 116.615 90.650 116.945 ;
        RECT 122.650 116.615 124.230 116.945 ;
        RECT 156.230 116.615 157.810 116.945 ;
        RECT 38.700 113.895 40.280 114.225 ;
        RECT 72.280 113.895 73.860 114.225 ;
        RECT 105.860 113.895 107.440 114.225 ;
        RECT 139.440 113.895 141.020 114.225 ;
        RECT 55.490 111.175 57.070 111.505 ;
        RECT 89.070 111.175 90.650 111.505 ;
        RECT 122.650 111.175 124.230 111.505 ;
        RECT 156.230 111.175 157.810 111.505 ;
        RECT 38.700 108.455 40.280 108.785 ;
        RECT 72.280 108.455 73.860 108.785 ;
        RECT 105.860 108.455 107.440 108.785 ;
        RECT 139.440 108.455 141.020 108.785 ;
        RECT 108.785 108.430 109.115 108.445 ;
        RECT 111.085 108.430 111.415 108.445 ;
        RECT 108.570 108.130 111.415 108.430 ;
        RECT 108.570 108.115 109.115 108.130 ;
        RECT 111.085 108.115 111.415 108.130 ;
        RECT 89.925 107.750 90.255 107.765 ;
        RECT 108.570 107.750 108.870 108.115 ;
        RECT 89.925 107.450 108.870 107.750 ;
        RECT 89.925 107.435 90.255 107.450 ;
        RECT 80.725 107.070 81.055 107.085 ;
        RECT 82.105 107.070 82.435 107.085 ;
        RECT 106.025 107.070 106.355 107.085 ;
        RECT 80.725 106.770 106.355 107.070 ;
        RECT 80.725 106.755 81.055 106.770 ;
        RECT 82.105 106.755 82.435 106.770 ;
        RECT 106.025 106.755 106.355 106.770 ;
        RECT 55.490 105.735 57.070 106.065 ;
        RECT 89.070 105.735 90.650 106.065 ;
        RECT 122.650 105.735 124.230 106.065 ;
        RECT 156.230 105.735 157.810 106.065 ;
        RECT 34.265 105.030 34.595 105.045 ;
        RECT 41.165 105.030 41.495 105.045 ;
        RECT 34.265 104.730 41.495 105.030 ;
        RECT 34.265 104.715 34.595 104.730 ;
        RECT 41.165 104.715 41.495 104.730 ;
        RECT 31.505 104.350 31.835 104.365 ;
        RECT 35.645 104.350 35.975 104.365 ;
        RECT 31.505 104.050 35.975 104.350 ;
        RECT 31.505 104.035 31.835 104.050 ;
        RECT 35.645 104.035 35.975 104.050 ;
        RECT 81.645 104.350 81.975 104.365 ;
        RECT 83.025 104.350 83.355 104.365 ;
        RECT 81.645 104.050 83.355 104.350 ;
        RECT 81.645 104.035 81.975 104.050 ;
        RECT 83.025 104.035 83.355 104.050 ;
        RECT 38.700 103.015 40.280 103.345 ;
        RECT 72.280 103.015 73.860 103.345 ;
        RECT 105.860 103.015 107.440 103.345 ;
        RECT 139.440 103.015 141.020 103.345 ;
        RECT 80.265 102.310 80.595 102.325 ;
        RECT 90.845 102.310 91.175 102.325 ;
        RECT 80.265 102.010 91.175 102.310 ;
        RECT 80.265 101.995 80.595 102.010 ;
        RECT 90.845 101.995 91.175 102.010 ;
        RECT 55.490 100.295 57.070 100.625 ;
        RECT 89.070 100.295 90.650 100.625 ;
        RECT 122.650 100.295 124.230 100.625 ;
        RECT 156.230 100.295 157.810 100.625 ;
        RECT 83.025 99.590 83.355 99.605 ;
        RECT 90.845 99.590 91.175 99.605 ;
        RECT 110.625 99.590 110.955 99.605 ;
        RECT 83.025 99.290 110.955 99.590 ;
        RECT 83.025 99.275 83.355 99.290 ;
        RECT 90.845 99.275 91.175 99.290 ;
        RECT 110.625 99.275 110.955 99.290 ;
        RECT 38.700 97.575 40.280 97.905 ;
        RECT 72.280 97.575 73.860 97.905 ;
        RECT 105.860 97.575 107.440 97.905 ;
        RECT 139.440 97.575 141.020 97.905 ;
        RECT 94.065 96.190 94.395 96.205 ;
        RECT 96.825 96.190 97.155 96.205 ;
        RECT 94.065 95.890 97.155 96.190 ;
        RECT 94.065 95.875 94.395 95.890 ;
        RECT 96.825 95.875 97.155 95.890 ;
        RECT 55.490 94.855 57.070 95.185 ;
        RECT 89.070 94.855 90.650 95.185 ;
        RECT 122.650 94.855 124.230 95.185 ;
        RECT 156.230 94.855 157.810 95.185 ;
        RECT 38.700 92.135 40.280 92.465 ;
        RECT 72.280 92.135 73.860 92.465 ;
        RECT 105.860 92.135 107.440 92.465 ;
        RECT 139.440 92.135 141.020 92.465 ;
        RECT 55.490 89.415 57.070 89.745 ;
        RECT 89.070 89.415 90.650 89.745 ;
        RECT 122.650 89.415 124.230 89.745 ;
        RECT 156.230 89.415 157.810 89.745 ;
        RECT 38.700 86.695 40.280 87.025 ;
        RECT 72.280 86.695 73.860 87.025 ;
        RECT 105.860 86.695 107.440 87.025 ;
        RECT 139.440 86.695 141.020 87.025 ;
        RECT 55.490 83.975 57.070 84.305 ;
        RECT 89.070 83.975 90.650 84.305 ;
        RECT 122.650 83.975 124.230 84.305 ;
        RECT 156.230 83.975 157.810 84.305 ;
        RECT 38.700 81.255 40.280 81.585 ;
        RECT 72.280 81.255 73.860 81.585 ;
        RECT 105.860 81.255 107.440 81.585 ;
        RECT 139.440 81.255 141.020 81.585 ;
        RECT 55.490 78.535 57.070 78.865 ;
        RECT 89.070 78.535 90.650 78.865 ;
        RECT 122.650 78.535 124.230 78.865 ;
        RECT 156.230 78.535 157.810 78.865 ;
        RECT 38.700 75.815 40.280 76.145 ;
        RECT 72.280 75.815 73.860 76.145 ;
        RECT 105.860 75.815 107.440 76.145 ;
        RECT 139.440 75.815 141.020 76.145 ;
        RECT 55.490 73.095 57.070 73.425 ;
        RECT 89.070 73.095 90.650 73.425 ;
        RECT 122.650 73.095 124.230 73.425 ;
        RECT 156.230 73.095 157.810 73.425 ;
        RECT 38.700 70.375 40.280 70.705 ;
        RECT 72.280 70.375 73.860 70.705 ;
        RECT 105.860 70.375 107.440 70.705 ;
        RECT 139.440 70.375 141.020 70.705 ;
        RECT 87.625 69.670 87.955 69.685 ;
        RECT 96.825 69.670 97.155 69.685 ;
        RECT 87.625 69.370 97.155 69.670 ;
        RECT 87.625 69.355 87.955 69.370 ;
        RECT 96.825 69.355 97.155 69.370 ;
        RECT 76.585 68.990 76.915 69.005 ;
        RECT 89.465 68.990 89.795 69.005 ;
        RECT 95.445 68.990 95.775 69.005 ;
        RECT 76.585 68.690 95.775 68.990 ;
        RECT 76.585 68.675 76.915 68.690 ;
        RECT 89.465 68.675 89.795 68.690 ;
        RECT 95.445 68.675 95.775 68.690 ;
        RECT 128.105 68.990 128.435 69.005 ;
        RECT 135.465 68.990 135.795 69.005 ;
        RECT 128.105 68.690 135.795 68.990 ;
        RECT 128.105 68.675 128.435 68.690 ;
        RECT 135.465 68.675 135.795 68.690 ;
        RECT 55.490 67.655 57.070 67.985 ;
        RECT 89.070 67.655 90.650 67.985 ;
        RECT 122.650 67.655 124.230 67.985 ;
        RECT 156.230 67.655 157.810 67.985 ;
        RECT 38.700 64.935 40.280 65.265 ;
        RECT 72.280 64.935 73.860 65.265 ;
        RECT 105.860 64.935 107.440 65.265 ;
        RECT 139.440 64.935 141.020 65.265 ;
        RECT 55.490 62.215 57.070 62.545 ;
        RECT 89.070 62.215 90.650 62.545 ;
        RECT 122.650 62.215 124.230 62.545 ;
        RECT 156.230 62.215 157.810 62.545 ;
        RECT 38.700 59.495 40.280 59.825 ;
        RECT 72.280 59.495 73.860 59.825 ;
        RECT 105.860 59.495 107.440 59.825 ;
        RECT 139.440 59.495 141.020 59.825 ;
        RECT 55.490 56.775 57.070 57.105 ;
        RECT 89.070 56.775 90.650 57.105 ;
        RECT 122.650 56.775 124.230 57.105 ;
        RECT 156.230 56.775 157.810 57.105 ;
        RECT 26.955 46.400 28.445 46.425 ;
        RECT 26.950 44.900 32.100 46.400 ;
        RECT 26.955 44.875 28.445 44.900 ;
        RECT 5.005 40.400 6.495 40.425 ;
        RECT 38.750 40.400 40.250 54.010 ;
        RECT 72.280 52.410 77.970 53.910 ;
        RECT 68.300 47.095 73.350 47.100 ;
        RECT 68.275 45.605 73.350 47.095 ;
        RECT 68.300 45.600 73.350 45.605 ;
        RECT 76.470 40.400 77.970 52.410 ;
        RECT 105.980 40.450 107.480 53.940 ;
        RECT 109.155 48.650 110.645 48.675 ;
        RECT 109.150 47.150 113.100 48.650 ;
        RECT 109.155 47.125 110.645 47.150 ;
        RECT 105.550 40.400 107.550 40.450 ;
        RECT 139.480 40.400 140.980 53.940 ;
        RECT 5.000 38.900 147.400 40.400 ;
        RECT 5.005 38.875 6.495 38.900 ;
        RECT 127.805 6.305 133.445 6.595 ;
        RECT 149.450 6.305 150.950 6.330 ;
        RECT 87.440 5.095 93.665 5.515 ;
        RECT 102.710 5.095 104.190 5.120 ;
        RECT 44.390 4.170 51.510 4.505 ;
        RECT 52.235 4.170 53.770 4.195 ;
        RECT 44.390 2.625 53.775 4.170 ;
        RECT 87.440 3.605 104.195 5.095 ;
        RECT 127.805 4.795 150.955 6.305 ;
        RECT 127.805 4.505 133.445 4.795 ;
        RECT 149.450 4.770 150.950 4.795 ;
        RECT 87.440 3.190 93.665 3.605 ;
        RECT 102.710 3.580 104.190 3.605 ;
        RECT 44.390 2.285 51.510 2.625 ;
        RECT 52.235 2.600 53.770 2.625 ;
      LAYER met4 ;
        RECT 3.990 224.500 4.290 224.760 ;
        RECT 3.950 224.000 4.350 224.500 ;
        RECT 7.670 224.000 7.970 224.760 ;
        RECT 11.350 224.000 11.650 224.760 ;
        RECT 15.030 224.000 15.330 224.760 ;
        RECT 18.710 224.000 19.010 224.760 ;
        RECT 22.390 224.000 22.690 224.760 ;
        RECT 26.070 224.000 26.370 224.760 ;
        RECT 29.750 224.000 30.050 224.760 ;
        RECT 33.430 224.000 33.730 224.760 ;
        RECT 37.110 224.000 37.410 224.760 ;
        RECT 40.790 224.000 41.090 224.760 ;
        RECT 44.470 224.000 44.770 224.760 ;
        RECT 48.150 224.000 48.450 224.760 ;
        RECT 51.830 224.000 52.130 224.760 ;
        RECT 55.510 224.000 55.810 224.760 ;
        RECT 59.190 224.000 59.490 224.760 ;
        RECT 62.870 224.000 63.170 224.760 ;
        RECT 66.550 224.000 66.850 224.760 ;
        RECT 70.230 224.000 70.530 224.760 ;
        RECT 73.910 224.000 74.210 224.760 ;
        RECT 77.590 224.000 77.890 224.760 ;
        RECT 81.270 224.215 81.570 224.760 ;
        RECT 84.950 224.215 85.250 224.760 ;
        RECT 88.630 224.215 88.930 224.760 ;
        RECT 92.310 224.300 92.610 224.760 ;
        RECT 95.990 224.300 96.290 224.760 ;
        RECT 99.670 224.300 99.970 224.760 ;
        RECT 103.350 224.300 103.650 224.760 ;
        RECT 3.950 223.700 77.890 224.000 ;
        RECT 81.255 223.885 81.585 224.215 ;
        RECT 84.935 223.885 85.265 224.215 ;
        RECT 88.615 223.885 88.945 224.215 ;
        RECT 3.950 223.600 74.200 223.700 ;
        RECT 7.650 222.500 74.200 223.600 ;
        RECT 107.030 223.400 107.330 224.760 ;
        RECT 75.150 223.100 107.330 223.400 ;
        RECT 9.000 220.760 10.500 222.500 ;
        RECT 75.150 219.200 75.450 223.100 ;
        RECT 110.710 222.800 111.010 224.760 ;
        RECT 49.000 218.900 75.450 219.200 ;
        RECT 75.950 222.500 111.010 222.800 ;
        RECT 49.000 215.865 49.300 218.900 ;
        RECT 75.950 218.550 76.250 222.500 ;
        RECT 114.390 222.200 114.690 224.760 ;
        RECT 56.350 218.250 76.250 218.550 ;
        RECT 76.750 221.900 114.690 222.200 ;
        RECT 56.350 215.865 56.650 218.250 ;
        RECT 63.700 215.865 64.000 215.900 ;
        RECT 48.985 215.535 49.315 215.865 ;
        RECT 56.335 215.535 56.665 215.865 ;
        RECT 63.685 215.850 64.015 215.865 ;
        RECT 70.250 215.850 70.550 215.900 ;
        RECT 76.750 215.850 77.050 221.900 ;
        RECT 118.070 221.550 118.370 224.760 ;
        RECT 77.600 221.250 118.370 221.550 ;
        RECT 77.600 215.850 77.900 221.250 ;
        RECT 79.185 220.900 79.515 220.915 ;
        RECT 121.750 220.900 122.050 224.760 ;
        RECT 79.185 220.600 122.050 220.900 ;
        RECT 79.185 220.585 79.515 220.600 ;
        RECT 86.585 220.200 86.915 220.215 ;
        RECT 125.430 220.200 125.730 224.760 ;
        RECT 86.585 219.900 125.730 220.200 ;
        RECT 86.585 219.885 86.915 219.900 ;
        RECT 94.035 219.550 94.365 219.565 ;
        RECT 129.110 219.550 129.410 224.760 ;
        RECT 94.035 219.250 129.410 219.550 ;
        RECT 94.035 219.235 94.365 219.250 ;
        RECT 101.485 218.850 101.815 218.865 ;
        RECT 132.790 218.850 133.090 224.760 ;
        RECT 101.485 218.550 133.090 218.850 ;
        RECT 101.485 218.535 101.815 218.550 ;
        RECT 108.685 218.150 109.015 218.165 ;
        RECT 136.470 218.150 136.770 224.760 ;
        RECT 108.685 217.850 136.770 218.150 ;
        RECT 108.685 217.835 109.015 217.850 ;
        RECT 116.035 217.400 116.365 217.415 ;
        RECT 140.150 217.400 140.450 224.760 ;
        RECT 116.035 217.100 140.450 217.400 ;
        RECT 116.035 217.085 116.365 217.100 ;
        RECT 123.385 216.750 123.715 216.765 ;
        RECT 143.830 216.750 144.130 224.760 ;
        RECT 123.385 216.450 144.130 216.750 ;
        RECT 123.385 216.435 123.715 216.450 ;
        RECT 63.685 215.550 77.050 215.850 ;
        RECT 77.550 215.550 77.900 215.850 ;
        RECT 130.835 216.100 131.165 216.115 ;
        RECT 147.510 216.100 147.810 224.760 ;
        RECT 130.835 215.800 147.810 216.100 ;
        RECT 130.835 215.785 131.165 215.800 ;
        RECT 63.685 215.535 64.015 215.550 ;
        RECT 71.935 214.900 72.265 214.915 ;
        RECT 77.600 214.900 77.900 215.550 ;
        RECT 138.555 215.460 138.885 215.475 ;
        RECT 151.190 215.460 151.490 224.760 ;
        RECT 138.555 215.160 151.490 215.460 ;
        RECT 138.555 215.145 138.885 215.160 ;
        RECT 71.935 214.600 77.900 214.900 ;
        RECT 145.865 214.790 146.195 214.805 ;
        RECT 154.870 214.790 155.170 224.760 ;
        RECT 71.935 214.585 72.265 214.600 ;
        RECT 145.865 214.490 155.170 214.790 ;
        RECT 145.865 214.475 146.195 214.490 ;
        RECT 153.495 214.140 153.825 214.155 ;
        RECT 158.550 214.140 158.850 224.760 ;
        RECT 153.495 213.840 158.850 214.140 ;
        RECT 153.495 213.825 153.825 213.840 ;
        RECT 38.690 56.700 40.290 209.500 ;
        RECT 45.995 163.875 46.325 164.205 ;
        RECT 46.010 132.245 46.310 163.875 ;
        RECT 45.995 131.915 46.325 132.245 ;
        RECT 55.480 56.700 57.080 209.500 ;
        RECT 72.270 56.700 73.870 209.500 ;
        RECT 75.435 164.555 75.765 164.885 ;
        RECT 75.450 143.805 75.750 164.555 ;
        RECT 76.355 163.875 76.685 164.205 ;
        RECT 75.435 143.475 75.765 143.805 ;
        RECT 76.370 130.205 76.670 163.875 ;
        RECT 82.795 150.955 83.125 151.285 ;
        RECT 82.810 137.685 83.110 150.955 ;
        RECT 82.795 137.355 83.125 137.685 ;
        RECT 76.355 129.875 76.685 130.205 ;
        RECT 82.810 124.085 83.110 137.355 ;
        RECT 82.795 123.755 83.125 124.085 ;
        RECT 89.060 56.700 90.660 209.500 ;
        RECT 103.035 183.595 103.365 183.925 ;
        RECT 100.275 152.995 100.605 153.325 ;
        RECT 100.290 137.685 100.590 152.995 ;
        RECT 103.050 150.605 103.350 183.595 ;
        RECT 103.035 150.275 103.365 150.605 ;
        RECT 100.275 137.355 100.605 137.685 ;
        RECT 105.850 63.040 107.450 209.500 ;
        RECT 108.555 191.075 108.885 191.405 ;
        RECT 108.570 183.925 108.870 191.075 ;
        RECT 108.555 183.595 108.885 183.925 ;
        RECT 108.570 150.605 108.870 183.595 ;
        RECT 109.475 182.235 109.805 182.565 ;
        RECT 109.490 172.365 109.790 182.235 ;
        RECT 109.475 172.035 109.805 172.365 ;
        RECT 108.555 150.275 108.885 150.605 ;
        RECT 109.490 145.845 109.790 172.035 ;
        RECT 109.475 145.515 109.805 145.845 ;
        RECT 122.640 63.040 124.240 209.500 ;
        RECT 105.850 56.700 107.480 63.040 ;
        RECT 122.640 56.700 124.270 63.040 ;
        RECT 139.430 56.700 141.030 209.500 ;
        RECT 156.220 56.700 157.820 209.500 ;
        RECT 38.750 53.985 40.250 56.700 ;
        RECT 38.745 52.475 40.255 53.985 ;
        RECT 55.490 48.650 56.990 56.700 ;
        RECT 72.310 53.915 73.810 56.700 ;
        RECT 72.305 52.405 73.815 53.915 ;
        RECT 89.130 48.650 90.630 56.700 ;
        RECT 105.980 53.915 107.480 56.700 ;
        RECT 105.975 52.405 107.485 53.915 ;
        RECT 122.770 48.650 124.270 56.700 ;
        RECT 139.480 53.915 140.980 56.700 ;
        RECT 139.475 52.405 140.985 53.915 ;
        RECT 156.250 48.650 157.750 56.700 ;
        RECT 10.500 47.150 157.750 48.650 ;
        RECT 26.950 44.900 28.450 47.150 ;
        RECT 68.300 45.600 69.800 47.150 ;
        RECT 2.500 38.900 6.500 40.400 ;
        RECT 149.445 6.300 157.300 6.305 ;
        RECT 108.150 5.095 109.850 5.100 ;
        RECT 60.880 4.170 64.470 4.175 ;
        RECT 52.230 2.625 64.470 4.170 ;
        RECT 102.705 3.900 109.850 5.095 ;
        RECT 149.445 4.795 157.310 6.300 ;
        RECT 102.705 3.605 135.230 3.900 ;
        RECT 108.100 3.000 135.230 3.605 ;
        RECT 62.925 2.280 64.470 2.625 ;
        RECT 62.925 1.430 113.150 2.280 ;
        RECT 63.200 1.380 113.150 1.430 ;
        RECT 112.250 1.000 113.150 1.380 ;
        RECT 134.330 1.000 135.230 3.000 ;
        RECT 156.410 1.000 157.310 4.795 ;
  END
END tt_um_rejunity_ay8913
END LIBRARY

