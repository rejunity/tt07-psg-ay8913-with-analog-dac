magic
tech sky130A
magscale 1 2
timestamp 1717176801
<< viali >>
rect 8401 30889 8435 30923
rect 11989 30889 12023 30923
rect 26525 30889 26559 30923
rect 10133 30821 10167 30855
rect 10333 30821 10367 30855
rect 17877 30821 17911 30855
rect 18337 30821 18371 30855
rect 18889 30821 18923 30855
rect 20453 30821 20487 30855
rect 20821 30821 20855 30855
rect 22293 30821 22327 30855
rect 5825 30753 5859 30787
rect 6377 30753 6411 30787
rect 6561 30753 6595 30787
rect 7021 30753 7055 30787
rect 7481 30753 7515 30787
rect 8585 30753 8619 30787
rect 8861 30753 8895 30787
rect 10425 30753 10459 30787
rect 11805 30753 11839 30787
rect 12173 30753 12207 30787
rect 12357 30753 12391 30787
rect 12541 30753 12575 30787
rect 14289 30753 14323 30787
rect 14749 30753 14783 30787
rect 16681 30753 16715 30787
rect 16773 30753 16807 30787
rect 17693 30753 17727 30787
rect 17785 30753 17819 30787
rect 18061 30753 18095 30787
rect 18705 30753 18739 30787
rect 18981 30753 19015 30787
rect 19073 30753 19107 30787
rect 22937 30753 22971 30787
rect 23857 30753 23891 30787
rect 26709 30753 26743 30787
rect 6929 30685 6963 30719
rect 8033 30685 8067 30719
rect 13093 30685 13127 30719
rect 13921 30685 13955 30719
rect 16405 30685 16439 30719
rect 19533 30685 19567 30719
rect 20177 30685 20211 30719
rect 24133 30685 24167 30719
rect 6653 30617 6687 30651
rect 9045 30617 9079 30651
rect 14124 30617 14158 30651
rect 16129 30617 16163 30651
rect 20637 30617 20671 30651
rect 6101 30549 6135 30583
rect 6285 30549 6319 30583
rect 6469 30549 6503 30583
rect 9965 30549 9999 30583
rect 10149 30549 10183 30583
rect 10609 30549 10643 30583
rect 12265 30549 12299 30583
rect 13645 30549 13679 30583
rect 14013 30549 14047 30583
rect 14933 30549 14967 30583
rect 16589 30549 16623 30583
rect 16957 30549 16991 30583
rect 17509 30549 17543 30583
rect 18245 30549 18279 30583
rect 19257 30549 19291 30583
rect 20361 30549 20395 30583
rect 22201 30549 22235 30583
rect 22753 30549 22787 30583
rect 8033 30345 8067 30379
rect 11161 30345 11195 30379
rect 12725 30345 12759 30379
rect 4629 30277 4663 30311
rect 16037 30277 16071 30311
rect 17877 30277 17911 30311
rect 20269 30277 20303 30311
rect 21189 30277 21223 30311
rect 21925 30277 21959 30311
rect 24133 30277 24167 30311
rect 6653 30209 6687 30243
rect 9505 30209 9539 30243
rect 11345 30209 11379 30243
rect 20453 30209 20487 30243
rect 20913 30209 20947 30243
rect 3065 30141 3099 30175
rect 3249 30141 3283 30175
rect 4813 30141 4847 30175
rect 6561 30141 6595 30175
rect 6920 30141 6954 30175
rect 8401 30141 8435 30175
rect 8585 30141 8619 30175
rect 8861 30141 8895 30175
rect 9137 30141 9171 30175
rect 9229 30141 9263 30175
rect 11069 30141 11103 30175
rect 11253 30141 11287 30175
rect 13093 30141 13127 30175
rect 13737 30141 13771 30175
rect 15301 30141 15335 30175
rect 15577 30141 15611 30175
rect 15761 30141 15795 30175
rect 17417 30141 17451 30175
rect 18521 30141 18555 30175
rect 18889 30141 18923 30175
rect 20545 30141 20579 30175
rect 21465 30141 21499 30175
rect 22293 30141 22327 30175
rect 22560 30141 22594 30175
rect 23857 30141 23891 30175
rect 25513 30141 25547 30175
rect 2798 30073 2832 30107
rect 3516 30073 3550 30107
rect 5058 30073 5092 30107
rect 9750 30073 9784 30107
rect 11590 30073 11624 30107
rect 15056 30073 15090 30107
rect 17150 30073 17184 30107
rect 19156 30073 19190 30107
rect 21557 30073 21591 30107
rect 25246 30073 25280 30107
rect 1685 30005 1719 30039
rect 6193 30005 6227 30039
rect 6377 30005 6411 30039
rect 8585 30005 8619 30039
rect 8677 30005 8711 30039
rect 9045 30005 9079 30039
rect 9413 30005 9447 30039
rect 10885 30005 10919 30039
rect 13277 30005 13311 30039
rect 13553 30005 13587 30039
rect 13921 30005 13955 30039
rect 15393 30005 15427 30039
rect 15945 30005 15979 30039
rect 21005 30005 21039 30039
rect 22017 30005 22051 30039
rect 23673 30005 23707 30039
rect 24041 30005 24075 30039
rect 949 29801 983 29835
rect 4353 29801 4387 29835
rect 9413 29801 9447 29835
rect 10149 29801 10183 29835
rect 10609 29801 10643 29835
rect 11897 29801 11931 29835
rect 11989 29801 12023 29835
rect 15393 29801 15427 29835
rect 16129 29801 16163 29835
rect 18705 29801 18739 29835
rect 24133 29801 24167 29835
rect 4629 29733 4663 29767
rect 11621 29733 11655 29767
rect 12992 29733 13026 29767
rect 14381 29733 14415 29767
rect 15209 29733 15243 29767
rect 16313 29733 16347 29767
rect 16865 29733 16899 29767
rect 22293 29733 22327 29767
rect 22477 29733 22511 29767
rect 22569 29733 22603 29767
rect 23121 29733 23155 29767
rect 23949 29733 23983 29767
rect 2073 29665 2107 29699
rect 2329 29665 2363 29699
rect 3801 29665 3835 29699
rect 3985 29665 4019 29699
rect 4169 29665 4203 29699
rect 5365 29665 5399 29699
rect 6009 29665 6043 29699
rect 6285 29665 6319 29699
rect 6561 29665 6595 29699
rect 7021 29665 7055 29699
rect 8300 29665 8334 29699
rect 10333 29665 10367 29699
rect 10517 29665 10551 29699
rect 10609 29665 10643 29699
rect 10793 29665 10827 29699
rect 11345 29665 11379 29699
rect 12081 29665 12115 29699
rect 14565 29665 14599 29699
rect 15669 29665 15703 29699
rect 15761 29665 15795 29699
rect 17592 29665 17626 29699
rect 18797 29665 18831 29699
rect 19053 29665 19087 29699
rect 21465 29665 21499 29699
rect 21833 29665 21867 29699
rect 21925 29665 21959 29699
rect 22661 29665 22695 29699
rect 22845 29665 22879 29699
rect 23581 29665 23615 29699
rect 24777 29665 24811 29699
rect 26433 29665 26467 29699
rect 6837 29597 6871 29631
rect 8033 29597 8067 29631
rect 12725 29597 12759 29631
rect 17325 29597 17359 29631
rect 20821 29597 20855 29631
rect 21373 29597 21407 29631
rect 21557 29597 21591 29631
rect 24685 29597 24719 29631
rect 26985 29597 27019 29631
rect 14841 29529 14875 29563
rect 15485 29529 15519 29563
rect 16681 29529 16715 29563
rect 20177 29529 20211 29563
rect 23489 29529 23523 29563
rect 25145 29529 25179 29563
rect 2605 29461 2639 29495
rect 3893 29461 3927 29495
rect 12265 29461 12299 29495
rect 14105 29461 14139 29495
rect 14749 29461 14783 29495
rect 15209 29461 15243 29495
rect 16313 29461 16347 29495
rect 16957 29461 16991 29495
rect 20269 29461 20303 29495
rect 21741 29461 21775 29495
rect 22017 29461 22051 29495
rect 22201 29461 22235 29495
rect 22937 29461 22971 29495
rect 23121 29461 23155 29495
rect 23949 29461 23983 29495
rect 6009 29257 6043 29291
rect 8585 29257 8619 29291
rect 11437 29257 11471 29291
rect 15669 29257 15703 29291
rect 16313 29257 16347 29291
rect 18705 29257 18739 29291
rect 20361 29257 20395 29291
rect 21465 29257 21499 29291
rect 22569 29257 22603 29291
rect 23121 29257 23155 29291
rect 26893 29257 26927 29291
rect 5917 29189 5951 29223
rect 8401 29189 8435 29223
rect 8953 29189 8987 29223
rect 9045 29189 9079 29223
rect 21649 29189 21683 29223
rect 3525 29121 3559 29155
rect 20545 29121 20579 29155
rect 21373 29121 21407 29155
rect 24041 29121 24075 29155
rect 3781 29053 3815 29087
rect 5181 29053 5215 29087
rect 5457 29053 5491 29087
rect 5549 29053 5583 29087
rect 6101 29053 6135 29087
rect 6193 29053 6227 29087
rect 9045 29053 9079 29087
rect 9229 29053 9263 29087
rect 9597 29053 9631 29087
rect 10057 29053 10091 29087
rect 10241 29053 10275 29087
rect 11621 29053 11655 29087
rect 11713 29053 11747 29087
rect 13185 29053 13219 29087
rect 15301 29053 15335 29087
rect 15485 29053 15519 29087
rect 16589 29053 16623 29087
rect 16773 29053 16807 29087
rect 16865 29053 16899 29087
rect 18889 29053 18923 29087
rect 19073 29053 19107 29087
rect 19257 29053 19291 29087
rect 20085 29053 20119 29087
rect 21281 29053 21315 29087
rect 23029 29053 23063 29087
rect 23305 29053 23339 29087
rect 23581 29053 23615 29087
rect 25513 29053 25547 29087
rect 5365 28985 5399 29019
rect 6377 28985 6411 29019
rect 10977 28985 11011 29019
rect 11161 28985 11195 29019
rect 11437 28985 11471 29019
rect 13001 28985 13035 29019
rect 16129 28985 16163 29019
rect 16681 28985 16715 29019
rect 18981 28985 19015 29019
rect 22385 28985 22419 29019
rect 23489 28985 23523 29019
rect 24308 28985 24342 29019
rect 25758 28985 25792 29019
rect 4905 28917 4939 28951
rect 4997 28917 5031 28951
rect 6101 28917 6135 28951
rect 8585 28917 8619 28951
rect 9413 28917 9447 28951
rect 10149 28917 10183 28951
rect 11345 28917 11379 28951
rect 13369 28917 13403 28951
rect 16329 28917 16363 28951
rect 16497 28917 16531 28951
rect 17049 28917 17083 28951
rect 22585 28917 22619 28951
rect 22753 28917 22787 28951
rect 22937 28917 22971 28951
rect 25421 28917 25455 28951
rect 4445 28713 4479 28747
rect 4613 28713 4647 28747
rect 5825 28713 5859 28747
rect 13277 28713 13311 28747
rect 13461 28713 13495 28747
rect 15225 28713 15259 28747
rect 15393 28713 15427 28747
rect 16497 28713 16531 28747
rect 23765 28713 23799 28747
rect 24225 28713 24259 28747
rect 25605 28713 25639 28747
rect 4813 28645 4847 28679
rect 8109 28645 8143 28679
rect 8309 28645 8343 28679
rect 9220 28645 9254 28679
rect 11621 28645 11655 28679
rect 14197 28645 14231 28679
rect 15025 28645 15059 28679
rect 16129 28645 16163 28679
rect 22201 28645 22235 28679
rect 3626 28577 3660 28611
rect 3893 28577 3927 28611
rect 6193 28577 6227 28611
rect 6736 28577 6770 28611
rect 8401 28577 8435 28611
rect 8493 28577 8527 28611
rect 8677 28577 8711 28611
rect 10413 28577 10447 28611
rect 10609 28577 10643 28611
rect 10977 28577 11011 28611
rect 12909 28577 12943 28611
rect 14473 28577 14507 28611
rect 14657 28577 14691 28611
rect 15577 28577 15611 28611
rect 16313 28577 16347 28611
rect 16773 28577 16807 28611
rect 17040 28577 17074 28611
rect 18337 28577 18371 28611
rect 18429 28577 18463 28611
rect 18705 28577 18739 28611
rect 18961 28577 18995 28611
rect 21373 28577 21407 28611
rect 22477 28577 22511 28611
rect 22661 28577 22695 28611
rect 23397 28577 23431 28611
rect 23581 28577 23615 28611
rect 24041 28577 24075 28611
rect 25421 28577 25455 28611
rect 25605 28577 25639 28611
rect 6285 28509 6319 28543
rect 6469 28509 6503 28543
rect 8953 28509 8987 28543
rect 13829 28509 13863 28543
rect 20177 28509 20211 28543
rect 20729 28509 20763 28543
rect 7941 28441 7975 28475
rect 8401 28441 8435 28475
rect 10333 28441 10367 28475
rect 10609 28441 10643 28475
rect 11253 28441 11287 28475
rect 14841 28441 14875 28475
rect 15761 28441 15795 28475
rect 20085 28441 20119 28475
rect 2513 28373 2547 28407
rect 4629 28373 4663 28407
rect 7849 28373 7883 28407
rect 8125 28373 8159 28407
rect 11069 28373 11103 28407
rect 11621 28373 11655 28407
rect 11805 28373 11839 28407
rect 13277 28373 13311 28407
rect 14197 28373 14231 28407
rect 14381 28373 14415 28407
rect 15209 28373 15243 28407
rect 18153 28373 18187 28407
rect 22293 28373 22327 28407
rect 3433 28169 3467 28203
rect 6101 28169 6135 28203
rect 6929 28169 6963 28203
rect 8125 28169 8159 28203
rect 9965 28169 9999 28203
rect 10149 28169 10183 28203
rect 13001 28169 13035 28203
rect 13737 28169 13771 28203
rect 13921 28169 13955 28203
rect 14013 28169 14047 28203
rect 18429 28169 18463 28203
rect 18705 28169 18739 28203
rect 20269 28169 20303 28203
rect 21097 28169 21131 28203
rect 21649 28169 21683 28203
rect 24041 28169 24075 28203
rect 24317 28169 24351 28203
rect 24501 28169 24535 28203
rect 10517 28101 10551 28135
rect 11161 28101 11195 28135
rect 17693 28101 17727 28135
rect 11345 28033 11379 28067
rect 13369 28033 13403 28067
rect 15393 28033 15427 28067
rect 17785 28033 17819 28067
rect 20637 28033 20671 28067
rect 21373 28033 21407 28067
rect 21465 28033 21499 28067
rect 23121 28033 23155 28067
rect 3249 27965 3283 27999
rect 4077 27965 4111 27999
rect 5549 27965 5583 27999
rect 5825 27965 5859 27999
rect 6469 27965 6503 27999
rect 7113 27965 7147 27999
rect 7665 27965 7699 27999
rect 7941 27965 7975 27999
rect 9689 27965 9723 27999
rect 10793 27965 10827 27999
rect 10885 27965 10919 27999
rect 10977 27965 11011 27999
rect 13185 27965 13219 27999
rect 15669 27965 15703 27999
rect 16313 27965 16347 27999
rect 18889 27965 18923 27999
rect 18981 27965 19015 27999
rect 19073 27965 19107 27999
rect 19257 27965 19291 27999
rect 20177 27965 20211 27999
rect 20821 27965 20855 27999
rect 21741 27965 21775 27999
rect 22201 27965 22235 27999
rect 22385 27965 22419 27999
rect 23029 27965 23063 27999
rect 23213 27965 23247 27999
rect 23673 27965 23707 27999
rect 25145 27965 25179 27999
rect 2789 27897 2823 27931
rect 2973 27897 3007 27931
rect 5641 27897 5675 27931
rect 7757 27897 7791 27931
rect 8953 27897 8987 27931
rect 10609 27897 10643 27931
rect 11612 27897 11646 27931
rect 13553 27897 13587 27931
rect 15126 27897 15160 27931
rect 16221 27897 16255 27931
rect 16558 27897 16592 27931
rect 20913 27897 20947 27931
rect 21097 27897 21131 27931
rect 21281 27897 21315 27931
rect 23305 27897 23339 27931
rect 23489 27897 23523 27931
rect 24009 27897 24043 27931
rect 24225 27897 24259 27931
rect 24469 27897 24503 27931
rect 24685 27897 24719 27931
rect 2605 27829 2639 27863
rect 3893 27829 3927 27863
rect 6285 27829 6319 27863
rect 6745 27829 6779 27863
rect 10149 27829 10183 27863
rect 12725 27829 12759 27863
rect 13753 27829 13787 27863
rect 22293 27829 22327 27863
rect 23857 27829 23891 27863
rect 25329 27829 25363 27863
rect 2881 27625 2915 27659
rect 6377 27625 6411 27659
rect 11621 27625 11655 27659
rect 14473 27625 14507 27659
rect 16405 27625 16439 27659
rect 23489 27625 23523 27659
rect 24869 27625 24903 27659
rect 2697 27557 2731 27591
rect 3792 27557 3826 27591
rect 5273 27557 5307 27591
rect 8585 27557 8619 27591
rect 16497 27557 16531 27591
rect 21465 27557 21499 27591
rect 22385 27557 22419 27591
rect 24593 27557 24627 27591
rect 25982 27557 26016 27591
rect 1869 27489 1903 27523
rect 3157 27489 3191 27523
rect 3525 27489 3559 27523
rect 5365 27489 5399 27523
rect 5457 27489 5491 27523
rect 5917 27489 5951 27523
rect 6285 27489 6319 27523
rect 7490 27489 7524 27523
rect 10701 27489 10735 27523
rect 11805 27489 11839 27523
rect 12081 27489 12115 27523
rect 13185 27489 13219 27523
rect 13737 27489 13771 27523
rect 14289 27489 14323 27523
rect 14933 27489 14967 27523
rect 15669 27489 15703 27523
rect 16129 27489 16163 27523
rect 16589 27489 16623 27523
rect 17785 27489 17819 27523
rect 17877 27489 17911 27523
rect 18133 27489 18167 27523
rect 19349 27489 19383 27523
rect 19605 27489 19639 27523
rect 21373 27489 21407 27523
rect 21649 27489 21683 27523
rect 21925 27489 21959 27523
rect 22661 27489 22695 27523
rect 22753 27489 22787 27523
rect 22845 27489 22879 27523
rect 23029 27489 23063 27523
rect 23397 27489 23431 27523
rect 23581 27489 23615 27523
rect 23857 27489 23891 27523
rect 26249 27489 26283 27523
rect 3341 27421 3375 27455
rect 6009 27421 6043 27455
rect 7757 27421 7791 27455
rect 9597 27421 9631 27455
rect 17049 27421 17083 27455
rect 22017 27421 22051 27455
rect 23765 27421 23799 27455
rect 2053 27353 2087 27387
rect 2329 27353 2363 27387
rect 5089 27353 5123 27387
rect 8953 27353 8987 27387
rect 9321 27353 9355 27387
rect 22477 27353 22511 27387
rect 24225 27353 24259 27387
rect 24777 27353 24811 27387
rect 2697 27285 2731 27319
rect 2973 27285 3007 27319
rect 4905 27285 4939 27319
rect 5641 27285 5675 27319
rect 5825 27285 5859 27319
rect 6193 27285 6227 27319
rect 9045 27285 9079 27319
rect 9137 27285 9171 27319
rect 10609 27285 10643 27319
rect 11989 27285 12023 27319
rect 13093 27285 13127 27319
rect 13645 27285 13679 27319
rect 14841 27285 14875 27319
rect 15577 27285 15611 27319
rect 19257 27285 19291 27319
rect 20729 27285 20763 27319
rect 21649 27285 21683 27319
rect 21741 27285 21775 27319
rect 22293 27285 22327 27319
rect 24593 27285 24627 27319
rect 2513 27081 2547 27115
rect 3985 27081 4019 27115
rect 4169 27081 4203 27115
rect 5641 27081 5675 27115
rect 5825 27081 5859 27115
rect 7573 27081 7607 27115
rect 8769 27081 8803 27115
rect 14565 27081 14599 27115
rect 17785 27081 17819 27115
rect 18521 27081 18555 27115
rect 21465 27081 21499 27115
rect 21833 27081 21867 27115
rect 23213 27081 23247 27115
rect 24225 27081 24259 27115
rect 25145 27081 25179 27115
rect 4537 27013 4571 27047
rect 10333 27013 10367 27047
rect 15117 27013 15151 27047
rect 21649 27013 21683 27047
rect 3617 26945 3651 26979
rect 4813 26945 4847 26979
rect 6929 26945 6963 26979
rect 11713 26945 11747 26979
rect 13185 26945 13219 26979
rect 19809 26945 19843 26979
rect 21281 26945 21315 26979
rect 857 26877 891 26911
rect 2881 26877 2915 26911
rect 4721 26877 4755 26911
rect 4905 26877 4939 26911
rect 4997 26877 5031 26911
rect 6101 26877 6135 26911
rect 6193 26877 6227 26911
rect 6469 26877 6503 26911
rect 6561 26877 6595 26911
rect 8125 26877 8159 26911
rect 8493 26877 8527 26911
rect 9045 26877 9079 26911
rect 9138 26877 9172 26911
rect 9551 26877 9585 26911
rect 9781 26877 9815 26911
rect 10057 26877 10091 26911
rect 10517 26877 10551 26911
rect 10609 26877 10643 26911
rect 10885 26877 10919 26911
rect 11437 26877 11471 26911
rect 11529 26877 11563 26911
rect 11805 26877 11839 26911
rect 11989 26877 12023 26911
rect 12173 26877 12207 26911
rect 12357 26877 12391 26911
rect 12909 26877 12943 26911
rect 13001 26877 13035 26911
rect 13277 26877 13311 26911
rect 13737 26877 13771 26911
rect 13829 26877 13863 26911
rect 14105 26877 14139 26911
rect 14289 26877 14323 26911
rect 14841 26877 14875 26911
rect 14933 26877 14967 26911
rect 15209 26877 15243 26911
rect 15577 26877 15611 26911
rect 15669 26877 15703 26911
rect 15853 26877 15887 26911
rect 15945 26877 15979 26911
rect 17233 26877 17267 26911
rect 17417 26877 17451 26911
rect 17601 26877 17635 26911
rect 17969 26877 18003 26911
rect 18153 26877 18187 26911
rect 18337 26877 18371 26911
rect 19349 26877 19383 26911
rect 20453 26877 20487 26911
rect 20913 26877 20947 26911
rect 21097 26877 21131 26911
rect 21189 26877 21223 26911
rect 21465 26877 21499 26911
rect 22017 26877 22051 26911
rect 22201 26877 22235 26911
rect 23305 26877 23339 26911
rect 23857 26877 23891 26911
rect 24409 26877 24443 26911
rect 24501 26877 24535 26911
rect 24685 26877 24719 26911
rect 24777 26877 24811 26911
rect 25605 26877 25639 26911
rect 1124 26809 1158 26843
rect 2513 26809 2547 26843
rect 3985 26809 4019 26843
rect 6377 26809 6411 26843
rect 9321 26809 9355 26843
rect 9413 26809 9447 26843
rect 10701 26809 10735 26843
rect 12265 26809 12299 26843
rect 13921 26809 13955 26843
rect 14565 26809 14599 26843
rect 15393 26809 15427 26843
rect 17509 26809 17543 26843
rect 18245 26809 18279 26843
rect 21005 26809 21039 26843
rect 24041 26809 24075 26843
rect 25872 26809 25906 26843
rect 2237 26741 2271 26775
rect 2329 26741 2363 26775
rect 6745 26741 6779 26775
rect 7481 26741 7515 26775
rect 8953 26741 8987 26775
rect 9689 26741 9723 26775
rect 9873 26741 9907 26775
rect 10241 26741 10275 26775
rect 11253 26741 11287 26775
rect 12541 26741 12575 26775
rect 12725 26741 12759 26775
rect 13553 26741 13587 26775
rect 14381 26741 14415 26775
rect 14657 26741 14691 26775
rect 18705 26741 18739 26775
rect 25145 26741 25179 26775
rect 25329 26741 25363 26775
rect 26985 26741 27019 26775
rect 1133 26537 1167 26571
rect 2789 26537 2823 26571
rect 5549 26537 5583 26571
rect 8033 26537 8067 26571
rect 9597 26537 9631 26571
rect 11437 26537 11471 26571
rect 13185 26537 13219 26571
rect 24015 26537 24049 26571
rect 25789 26537 25823 26571
rect 2497 26469 2531 26503
rect 2697 26469 2731 26503
rect 2973 26469 3007 26503
rect 8401 26469 8435 26503
rect 8617 26469 8651 26503
rect 10577 26469 10611 26503
rect 10793 26469 10827 26503
rect 11805 26469 11839 26503
rect 12817 26469 12851 26503
rect 15945 26469 15979 26503
rect 19625 26469 19659 26503
rect 20453 26469 20487 26503
rect 21281 26469 21315 26503
rect 24225 26469 24259 26503
rect 24869 26469 24903 26503
rect 25053 26469 25087 26503
rect 1317 26401 1351 26435
rect 3157 26401 3191 26435
rect 3249 26401 3283 26435
rect 3341 26401 3375 26435
rect 5365 26401 5399 26435
rect 5641 26401 5675 26435
rect 5825 26401 5859 26435
rect 5917 26401 5951 26435
rect 6101 26401 6135 26435
rect 6193 26401 6227 26435
rect 6653 26401 6687 26435
rect 6909 26401 6943 26435
rect 9045 26401 9079 26435
rect 9229 26401 9263 26435
rect 9321 26401 9355 26435
rect 10149 26401 10183 26435
rect 11345 26401 11379 26435
rect 11621 26401 11655 26435
rect 12081 26401 12115 26435
rect 12265 26401 12299 26435
rect 12357 26401 12391 26435
rect 12725 26401 12759 26435
rect 13001 26401 13035 26435
rect 15669 26401 15703 26435
rect 15761 26401 15795 26435
rect 16129 26401 16163 26435
rect 16313 26401 16347 26435
rect 16681 26401 16715 26435
rect 17325 26401 17359 26435
rect 17785 26401 17819 26435
rect 18061 26401 18095 26435
rect 18245 26401 18279 26435
rect 18337 26401 18371 26435
rect 18429 26401 18463 26435
rect 20637 26401 20671 26435
rect 20729 26401 20763 26435
rect 21005 26401 21039 26435
rect 21557 26401 21591 26435
rect 21833 26401 21867 26435
rect 23121 26401 23155 26435
rect 25605 26401 25639 26435
rect 3985 26333 4019 26367
rect 15945 26333 15979 26367
rect 17049 26333 17083 26367
rect 17693 26333 17727 26367
rect 19349 26333 19383 26367
rect 20269 26333 20303 26367
rect 21465 26333 21499 26367
rect 2329 26265 2363 26299
rect 4261 26265 4295 26299
rect 6377 26265 6411 26299
rect 8769 26265 8803 26299
rect 16313 26265 16347 26299
rect 16773 26265 16807 26299
rect 17417 26265 17451 26299
rect 18705 26265 18739 26299
rect 21373 26265 21407 26299
rect 21649 26265 21683 26299
rect 23857 26265 23891 26299
rect 2513 26197 2547 26231
rect 4445 26197 4479 26231
rect 5181 26197 5215 26231
rect 8585 26197 8619 26231
rect 8861 26197 8895 26231
rect 10425 26197 10459 26231
rect 10609 26197 10643 26231
rect 11897 26197 11931 26231
rect 16957 26197 16991 26231
rect 18613 26197 18647 26231
rect 20913 26197 20947 26231
rect 23305 26197 23339 26231
rect 24041 26197 24075 26231
rect 24685 26197 24719 26231
rect 7021 25993 7055 26027
rect 8033 25993 8067 26027
rect 9965 25993 9999 26027
rect 10425 25993 10459 26027
rect 11897 25993 11931 26027
rect 14933 25993 14967 26027
rect 16405 25993 16439 26027
rect 20453 25993 20487 26027
rect 22293 25993 22327 26027
rect 23857 25993 23891 26027
rect 24041 25993 24075 26027
rect 24685 25993 24719 26027
rect 24961 25993 24995 26027
rect 20729 25925 20763 25959
rect 24317 25925 24351 25959
rect 4997 25857 5031 25891
rect 11713 25857 11747 25891
rect 13553 25857 13587 25891
rect 15393 25857 15427 25891
rect 15853 25857 15887 25891
rect 16773 25857 16807 25891
rect 18705 25857 18739 25891
rect 21281 25857 21315 25891
rect 23673 25857 23707 25891
rect 2329 25789 2363 25823
rect 2513 25789 2547 25823
rect 2605 25789 2639 25823
rect 2789 25789 2823 25823
rect 2881 25789 2915 25823
rect 4905 25789 4939 25823
rect 5089 25789 5123 25823
rect 5181 25789 5215 25823
rect 7205 25789 7239 25823
rect 7389 25789 7423 25823
rect 7573 25789 7607 25823
rect 8401 25789 8435 25823
rect 8668 25789 8702 25823
rect 10149 25789 10183 25823
rect 10241 25789 10275 25823
rect 10517 25789 10551 25823
rect 12449 25789 12483 25823
rect 12817 25789 12851 25823
rect 15209 25789 15243 25823
rect 15485 25789 15519 25823
rect 15669 25789 15703 25823
rect 16589 25789 16623 25823
rect 17877 25789 17911 25823
rect 18061 25789 18095 25823
rect 18245 25789 18279 25823
rect 18961 25789 18995 25823
rect 20177 25789 20211 25823
rect 20913 25789 20947 25823
rect 21005 25789 21039 25823
rect 21189 25789 21223 25823
rect 23406 25789 23440 25823
rect 26341 25789 26375 25823
rect 2697 25721 2731 25755
rect 3249 25721 3283 25755
rect 3985 25721 4019 25755
rect 7297 25721 7331 25755
rect 7849 25721 7883 25755
rect 8049 25721 8083 25755
rect 10885 25721 10919 25755
rect 13798 25721 13832 25755
rect 17969 25721 18003 25755
rect 20453 25721 20487 25755
rect 24225 25721 24259 25755
rect 26074 25721 26108 25755
rect 2329 25653 2363 25687
rect 3065 25653 3099 25687
rect 4721 25653 4755 25687
rect 8217 25653 8251 25687
rect 9781 25653 9815 25687
rect 13369 25653 13403 25687
rect 15025 25653 15059 25687
rect 17693 25653 17727 25687
rect 20085 25653 20119 25687
rect 20269 25653 20303 25687
rect 24015 25653 24049 25687
rect 24685 25653 24719 25687
rect 24869 25653 24903 25687
rect 4169 25449 4203 25483
rect 4445 25449 4479 25483
rect 5641 25449 5675 25483
rect 9965 25449 9999 25483
rect 12633 25449 12667 25483
rect 13921 25449 13955 25483
rect 14381 25449 14415 25483
rect 14841 25449 14875 25483
rect 19165 25449 19199 25483
rect 20269 25449 20303 25483
rect 21373 25449 21407 25483
rect 23397 25449 23431 25483
rect 24777 25449 24811 25483
rect 25237 25449 25271 25483
rect 7941 25381 7975 25415
rect 9505 25381 9539 25415
rect 11428 25381 11462 25415
rect 12785 25381 12819 25415
rect 13001 25381 13035 25415
rect 18030 25381 18064 25415
rect 23765 25381 23799 25415
rect 24685 25381 24719 25415
rect 857 25313 891 25347
rect 1124 25313 1158 25347
rect 2329 25313 2363 25347
rect 2513 25313 2547 25347
rect 2789 25313 2823 25347
rect 3056 25313 3090 25347
rect 4997 25313 5031 25347
rect 5089 25313 5123 25347
rect 7021 25313 7055 25347
rect 7297 25313 7331 25347
rect 7757 25313 7791 25347
rect 7849 25313 7883 25347
rect 8125 25313 8159 25347
rect 8493 25313 8527 25347
rect 9413 25313 9447 25347
rect 9689 25313 9723 25347
rect 10517 25313 10551 25347
rect 11161 25313 11195 25347
rect 14105 25313 14139 25347
rect 14749 25313 14783 25347
rect 20177 25313 20211 25347
rect 21833 25313 21867 25347
rect 22293 25313 22327 25347
rect 22477 25313 22511 25347
rect 22937 25313 22971 25347
rect 23581 25313 23615 25347
rect 23857 25313 23891 25347
rect 24041 25313 24075 25347
rect 25053 25313 25087 25347
rect 25329 25313 25363 25347
rect 4721 25245 4755 25279
rect 5365 25245 5399 25279
rect 6929 25245 6963 25279
rect 9045 25245 9079 25279
rect 15025 25245 15059 25279
rect 17785 25245 17819 25279
rect 21741 25245 21775 25279
rect 22017 25245 22051 25279
rect 22201 25245 22235 25279
rect 22385 25245 22419 25279
rect 22661 25245 22695 25279
rect 22753 25245 22787 25279
rect 26065 25245 26099 25279
rect 9873 25177 9907 25211
rect 2237 25109 2271 25143
rect 2697 25109 2731 25143
rect 4629 25109 4663 25143
rect 5181 25109 5215 25143
rect 7573 25109 7607 25143
rect 12541 25109 12575 25143
rect 12817 25109 12851 25143
rect 23121 25109 23155 25143
rect 23949 25109 23983 25143
rect 1041 24905 1075 24939
rect 1869 24905 1903 24939
rect 2605 24905 2639 24939
rect 2789 24905 2823 24939
rect 4169 24905 4203 24939
rect 4537 24905 4571 24939
rect 5273 24905 5307 24939
rect 10057 24905 10091 24939
rect 11529 24905 11563 24939
rect 14565 24905 14599 24939
rect 22109 24905 22143 24939
rect 23121 24905 23155 24939
rect 24041 24905 24075 24939
rect 18061 24837 18095 24871
rect 22017 24837 22051 24871
rect 24225 24837 24259 24871
rect 2973 24769 3007 24803
rect 4997 24769 5031 24803
rect 11989 24769 12023 24803
rect 13645 24769 13679 24803
rect 14289 24769 14323 24803
rect 15485 24769 15519 24803
rect 19349 24769 19383 24803
rect 23305 24769 23339 24803
rect 1225 24701 1259 24735
rect 2881 24701 2915 24735
rect 4077 24701 4111 24735
rect 4905 24701 4939 24735
rect 7113 24701 7147 24735
rect 7849 24701 7883 24735
rect 8677 24701 8711 24735
rect 10149 24701 10183 24735
rect 10416 24701 10450 24735
rect 15025 24701 15059 24735
rect 15301 24701 15335 24735
rect 15669 24701 15703 24735
rect 15945 24701 15979 24735
rect 17601 24701 17635 24735
rect 17693 24701 17727 24735
rect 18061 24701 18095 24735
rect 18337 24701 18371 24735
rect 19073 24701 19107 24735
rect 23029 24701 23063 24735
rect 24317 24701 24351 24735
rect 24593 24701 24627 24735
rect 24859 24701 24893 24735
rect 25053 24701 25087 24735
rect 25145 24701 25179 24735
rect 25329 24701 25363 24735
rect 25697 24701 25731 24735
rect 14519 24667 14553 24701
rect 1853 24633 1887 24667
rect 2053 24633 2087 24667
rect 2421 24633 2455 24667
rect 2637 24633 2671 24667
rect 6846 24633 6880 24667
rect 8944 24633 8978 24667
rect 12256 24633 12290 24667
rect 14749 24633 14783 24667
rect 16190 24633 16224 24667
rect 19594 24633 19628 24667
rect 21649 24633 21683 24667
rect 23857 24633 23891 24667
rect 24057 24633 24091 24667
rect 25964 24633 25998 24667
rect 1685 24565 1719 24599
rect 5733 24565 5767 24599
rect 7205 24565 7239 24599
rect 13369 24565 13403 24599
rect 14381 24565 14415 24599
rect 14841 24565 14875 24599
rect 15117 24565 15151 24599
rect 15853 24565 15887 24599
rect 17325 24565 17359 24599
rect 17417 24565 17451 24599
rect 19257 24565 19291 24599
rect 20729 24565 20763 24599
rect 23581 24565 23615 24599
rect 24409 24565 24443 24599
rect 24777 24565 24811 24599
rect 25053 24565 25087 24599
rect 25329 24565 25363 24599
rect 27077 24565 27111 24599
rect 6193 24361 6227 24395
rect 8861 24361 8895 24395
rect 9321 24361 9355 24395
rect 10307 24361 10341 24395
rect 12633 24361 12667 24395
rect 13001 24361 13035 24395
rect 15577 24361 15611 24395
rect 16129 24361 16163 24395
rect 16589 24361 16623 24395
rect 19533 24361 19567 24395
rect 22109 24361 22143 24395
rect 23581 24361 23615 24395
rect 24409 24361 24443 24395
rect 25513 24361 25547 24395
rect 25805 24361 25839 24395
rect 26065 24361 26099 24395
rect 6561 24293 6595 24327
rect 7021 24293 7055 24327
rect 7113 24293 7147 24327
rect 7726 24293 7760 24327
rect 10517 24293 10551 24327
rect 10977 24293 11011 24327
rect 23397 24293 23431 24327
rect 24685 24293 24719 24327
rect 24869 24293 24903 24327
rect 25605 24293 25639 24327
rect 26801 24293 26835 24327
rect 1777 24225 1811 24259
rect 1961 24225 1995 24259
rect 2237 24225 2271 24259
rect 2881 24225 2915 24259
rect 4813 24225 4847 24259
rect 6377 24225 6411 24259
rect 6469 24225 6503 24259
rect 6745 24225 6779 24259
rect 6837 24225 6871 24259
rect 7205 24225 7239 24259
rect 9505 24225 9539 24259
rect 9689 24225 9723 24259
rect 9781 24225 9815 24259
rect 11897 24225 11931 24259
rect 12817 24225 12851 24259
rect 13093 24225 13127 24259
rect 14197 24225 14231 24259
rect 14464 24225 14498 24259
rect 16497 24225 16531 24259
rect 17785 24225 17819 24259
rect 19073 24225 19107 24259
rect 19901 24225 19935 24259
rect 19993 24225 20027 24259
rect 20361 24225 20395 24259
rect 20545 24225 20579 24259
rect 20729 24225 20763 24259
rect 21373 24225 21407 24259
rect 21557 24225 21591 24259
rect 21649 24225 21683 24259
rect 21925 24225 21959 24259
rect 23673 24225 23707 24259
rect 25145 24225 25179 24259
rect 25329 24225 25363 24259
rect 26249 24225 26283 24259
rect 26893 24225 26927 24259
rect 2421 24157 2455 24191
rect 7481 24157 7515 24191
rect 11529 24157 11563 24191
rect 16681 24157 16715 24191
rect 17969 24157 18003 24191
rect 19257 24157 19291 24191
rect 20085 24157 20119 24191
rect 21741 24157 21775 24191
rect 23305 24157 23339 24191
rect 23765 24157 23799 24191
rect 11713 24089 11747 24123
rect 23397 24089 23431 24123
rect 25973 24089 26007 24123
rect 1869 24021 1903 24055
rect 2053 24021 2087 24055
rect 2789 24021 2823 24055
rect 4353 24021 4387 24055
rect 4721 24021 4755 24055
rect 7389 24021 7423 24055
rect 10149 24021 10183 24055
rect 10333 24021 10367 24055
rect 17601 24021 17635 24055
rect 18889 24021 18923 24055
rect 22661 24021 22695 24055
rect 24501 24021 24535 24055
rect 25789 24021 25823 24055
rect 1225 23817 1259 23851
rect 1593 23817 1627 23851
rect 2329 23817 2363 23851
rect 2789 23817 2823 23851
rect 4905 23817 4939 23851
rect 4997 23817 5031 23851
rect 5365 23817 5399 23851
rect 8401 23817 8435 23851
rect 10885 23817 10919 23851
rect 12725 23817 12759 23851
rect 13737 23817 13771 23851
rect 14657 23817 14691 23851
rect 18153 23817 18187 23851
rect 20821 23817 20855 23851
rect 23673 23817 23707 23851
rect 24041 23817 24075 23851
rect 1409 23749 1443 23783
rect 2513 23749 2547 23783
rect 14013 23749 14047 23783
rect 20085 23749 20119 23783
rect 21281 23749 21315 23783
rect 21373 23749 21407 23783
rect 5457 23681 5491 23715
rect 9505 23681 9539 23715
rect 10977 23681 11011 23715
rect 15117 23681 15151 23715
rect 15209 23681 15243 23715
rect 16773 23681 16807 23715
rect 18705 23681 18739 23715
rect 25513 23681 25547 23715
rect 857 23613 891 23647
rect 1133 23613 1167 23647
rect 1317 23613 1351 23647
rect 1961 23613 1995 23647
rect 3433 23613 3467 23647
rect 3801 23613 3835 23647
rect 3893 23613 3927 23647
rect 3985 23613 4019 23647
rect 4077 23613 4111 23647
rect 4353 23613 4387 23647
rect 4629 23613 4663 23647
rect 4721 23613 4755 23647
rect 4997 23613 5031 23647
rect 5089 23613 5123 23647
rect 7757 23613 7791 23647
rect 8953 23613 8987 23647
rect 11161 23613 11195 23647
rect 11345 23613 11379 23647
rect 12817 23613 12851 23647
rect 13093 23613 13127 23647
rect 14197 23613 14231 23647
rect 16497 23613 16531 23647
rect 18337 23613 18371 23647
rect 20361 23613 20395 23647
rect 20545 23613 20579 23647
rect 20729 23613 20763 23647
rect 21005 23613 21039 23647
rect 21097 23613 21131 23647
rect 21511 23613 21545 23647
rect 21741 23613 21775 23647
rect 21869 23613 21903 23647
rect 22017 23613 22051 23647
rect 22293 23613 22327 23647
rect 25421 23613 25455 23647
rect 25973 23613 26007 23647
rect 26709 23613 26743 23647
rect 2145 23545 2179 23579
rect 2757 23545 2791 23579
rect 2973 23545 3007 23579
rect 3525 23545 3559 23579
rect 4537 23545 4571 23579
rect 5724 23545 5758 23579
rect 9772 23545 9806 23579
rect 11612 23545 11646 23579
rect 13921 23545 13955 23579
rect 16037 23545 16071 23579
rect 17018 23545 17052 23579
rect 18950 23545 18984 23579
rect 21649 23545 21683 23579
rect 22560 23545 22594 23579
rect 25154 23545 25188 23579
rect 25881 23545 25915 23579
rect 26617 23545 26651 23579
rect 1041 23477 1075 23511
rect 1593 23477 1627 23511
rect 2345 23477 2379 23511
rect 2605 23477 2639 23511
rect 4261 23477 4295 23511
rect 6837 23477 6871 23511
rect 7205 23477 7239 23511
rect 12909 23477 12943 23511
rect 13553 23477 13587 23511
rect 13721 23477 13755 23511
rect 15025 23477 15059 23511
rect 16129 23477 16163 23511
rect 16681 23477 16715 23511
rect 18521 23477 18555 23511
rect 20177 23477 20211 23511
rect 25789 23477 25823 23511
rect 2237 23273 2271 23307
rect 2973 23273 3007 23307
rect 3617 23273 3651 23307
rect 4077 23273 4111 23307
rect 6469 23273 6503 23307
rect 7665 23273 7699 23307
rect 9965 23273 9999 23307
rect 12817 23273 12851 23307
rect 14749 23273 14783 23307
rect 17049 23273 17083 23307
rect 17509 23273 17543 23307
rect 18429 23273 18463 23307
rect 18889 23273 18923 23307
rect 19625 23273 19659 23307
rect 21281 23273 21315 23307
rect 21925 23273 21959 23307
rect 24685 23273 24719 23307
rect 26433 23273 26467 23307
rect 3341 23205 3375 23239
rect 7297 23205 7331 23239
rect 7389 23205 7423 23239
rect 8870 23205 8904 23239
rect 11805 23205 11839 23239
rect 12173 23205 12207 23239
rect 13636 23205 13670 23239
rect 17417 23205 17451 23239
rect 19962 23205 19996 23239
rect 22201 23205 22235 23239
rect 24317 23205 24351 23239
rect 24533 23205 24567 23239
rect 1124 23137 1158 23171
rect 2513 23137 2547 23171
rect 3065 23137 3099 23171
rect 3249 23137 3283 23171
rect 3433 23137 3467 23171
rect 4261 23137 4295 23171
rect 4537 23137 4571 23171
rect 4629 23137 4663 23171
rect 4813 23137 4847 23171
rect 5917 23137 5951 23171
rect 6193 23137 6227 23171
rect 6653 23137 6687 23171
rect 6745 23137 6779 23171
rect 6837 23137 6871 23171
rect 7021 23137 7055 23171
rect 7113 23137 7147 23171
rect 7481 23137 7515 23171
rect 9137 23137 9171 23171
rect 10149 23137 10183 23171
rect 10333 23137 10367 23171
rect 10425 23137 10459 23171
rect 11989 23137 12023 23171
rect 12265 23137 12299 23171
rect 12909 23137 12943 23171
rect 15485 23137 15519 23171
rect 15669 23137 15703 23171
rect 15761 23137 15795 23171
rect 16497 23137 16531 23171
rect 18797 23137 18831 23171
rect 19441 23137 19475 23171
rect 21465 23137 21499 23171
rect 21557 23137 21591 23171
rect 21833 23137 21867 23171
rect 22109 23137 22143 23171
rect 22293 23137 22327 23171
rect 22477 23137 22511 23171
rect 23857 23137 23891 23171
rect 857 23069 891 23103
rect 4077 23069 4111 23103
rect 4169 23069 4203 23103
rect 4445 23069 4479 23103
rect 12725 23069 12759 23103
rect 13369 23069 13403 23103
rect 15945 23069 15979 23103
rect 16589 23069 16623 23103
rect 16681 23069 16715 23103
rect 17693 23069 17727 23103
rect 19073 23069 19107 23103
rect 19717 23069 19751 23103
rect 23765 23069 23799 23103
rect 26985 23069 27019 23103
rect 7757 23001 7791 23035
rect 16129 23001 16163 23035
rect 21097 23001 21131 23035
rect 2789 22933 2823 22967
rect 4721 22933 4755 22967
rect 13277 22933 13311 22967
rect 15301 22933 15335 22967
rect 21741 22933 21775 22967
rect 24501 22933 24535 22967
rect 2421 22729 2455 22763
rect 3525 22729 3559 22763
rect 3709 22729 3743 22763
rect 5273 22729 5307 22763
rect 7205 22729 7239 22763
rect 9873 22729 9907 22763
rect 11989 22729 12023 22763
rect 13369 22729 13403 22763
rect 16589 22729 16623 22763
rect 19625 22729 19659 22763
rect 26893 22729 26927 22763
rect 5089 22661 5123 22695
rect 7481 22661 7515 22695
rect 13829 22661 13863 22695
rect 14381 22661 14415 22695
rect 16681 22661 16715 22695
rect 17509 22661 17543 22695
rect 5365 22593 5399 22627
rect 10701 22593 10735 22627
rect 11345 22593 11379 22627
rect 11529 22593 11563 22627
rect 12541 22593 12575 22627
rect 17969 22593 18003 22627
rect 20177 22593 20211 22627
rect 25513 22593 25547 22627
rect 2605 22525 2639 22559
rect 2697 22525 2731 22559
rect 3249 22525 3283 22559
rect 4537 22525 4571 22559
rect 4813 22525 4847 22559
rect 5457 22525 5491 22559
rect 5549 22525 5583 22559
rect 8033 22525 8067 22559
rect 8493 22525 8527 22559
rect 12173 22525 12207 22559
rect 13001 22525 13035 22559
rect 13185 22525 13219 22559
rect 13553 22525 13587 22559
rect 13737 22525 13771 22559
rect 15209 22525 15243 22559
rect 15476 22525 15510 22559
rect 17141 22525 17175 22559
rect 17601 22525 17635 22559
rect 17785 22525 17819 22559
rect 22385 22525 22419 22559
rect 22569 22525 22603 22559
rect 22661 22525 22695 22559
rect 22937 22525 22971 22559
rect 23213 22525 23247 22559
rect 23857 22525 23891 22559
rect 25780 22525 25814 22559
rect 2973 22457 3007 22491
rect 5816 22457 5850 22491
rect 7389 22457 7423 22491
rect 8760 22457 8794 22491
rect 14013 22457 14047 22491
rect 14197 22457 14231 22491
rect 16865 22457 16899 22491
rect 17049 22457 17083 22491
rect 17325 22457 17359 22491
rect 19993 22457 20027 22491
rect 20085 22457 20119 22491
rect 2789 22389 2823 22423
rect 4629 22389 4663 22423
rect 4997 22389 5031 22423
rect 6929 22389 6963 22423
rect 7021 22389 7055 22423
rect 7189 22389 7223 22423
rect 10149 22389 10183 22423
rect 10885 22389 10919 22423
rect 11253 22389 11287 22423
rect 12357 22389 12391 22423
rect 22477 22389 22511 22423
rect 22753 22389 22787 22423
rect 23121 22389 23155 22423
rect 23397 22389 23431 22423
rect 24041 22389 24075 22423
rect 4997 22185 5031 22219
rect 7481 22185 7515 22219
rect 9045 22185 9079 22219
rect 9949 22185 9983 22219
rect 13369 22185 13403 22219
rect 16313 22185 16347 22219
rect 22109 22185 22143 22219
rect 23213 22185 23247 22219
rect 1777 22117 1811 22151
rect 10149 22117 10183 22151
rect 13921 22117 13955 22151
rect 15761 22117 15795 22151
rect 21833 22117 21867 22151
rect 22017 22117 22051 22151
rect 22477 22117 22511 22151
rect 22845 22117 22879 22151
rect 23045 22117 23079 22151
rect 1961 22049 1995 22083
rect 3065 22049 3099 22083
rect 4905 22049 4939 22083
rect 5089 22049 5123 22083
rect 5641 22049 5675 22083
rect 6285 22049 6319 22083
rect 6929 22049 6963 22083
rect 8594 22049 8628 22083
rect 9229 22049 9263 22083
rect 9413 22049 9447 22083
rect 9505 22049 9539 22083
rect 10425 22049 10459 22083
rect 10609 22049 10643 22083
rect 10977 22049 11011 22083
rect 11805 22049 11839 22083
rect 12449 22049 12483 22083
rect 12633 22049 12667 22083
rect 13829 22049 13863 22083
rect 15025 22049 15059 22083
rect 15577 22049 15611 22083
rect 15945 22049 15979 22083
rect 16129 22049 16163 22083
rect 17141 22049 17175 22083
rect 17877 22049 17911 22083
rect 18797 22049 18831 22083
rect 19064 22049 19098 22083
rect 22109 22049 22143 22083
rect 22385 22049 22419 22083
rect 22569 22049 22603 22083
rect 24418 22049 24452 22083
rect 5365 21981 5399 22015
rect 6101 21981 6135 22015
rect 8861 21981 8895 22015
rect 10241 21981 10275 22015
rect 14749 21981 14783 22015
rect 15301 21981 15335 22015
rect 20361 21981 20395 22015
rect 24685 21981 24719 22015
rect 9781 21913 9815 21947
rect 17325 21913 17359 21947
rect 17785 21913 17819 21947
rect 20177 21913 20211 21947
rect 22201 21913 22235 21947
rect 23305 21913 23339 21947
rect 1593 21845 1627 21879
rect 3157 21845 3191 21879
rect 6377 21845 6411 21879
rect 9965 21845 9999 21879
rect 11161 21845 11195 21879
rect 12173 21845 12207 21879
rect 13737 21845 13771 21879
rect 15393 21845 15427 21879
rect 20913 21845 20947 21879
rect 22753 21845 22787 21879
rect 23029 21845 23063 21879
rect 2697 21641 2731 21675
rect 4905 21641 4939 21675
rect 5917 21641 5951 21675
rect 7205 21641 7239 21675
rect 8585 21641 8619 21675
rect 10149 21641 10183 21675
rect 20269 21641 20303 21675
rect 22293 21641 22327 21675
rect 23121 21641 23155 21675
rect 23305 21641 23339 21675
rect 2329 21573 2363 21607
rect 14749 21573 14783 21607
rect 18521 21573 18555 21607
rect 22753 21573 22787 21607
rect 23857 21573 23891 21607
rect 3249 21505 3283 21539
rect 13093 21505 13127 21539
rect 14197 21505 14231 21539
rect 17141 21505 17175 21539
rect 19257 21505 19291 21539
rect 25237 21505 25271 21539
rect 25329 21505 25363 21539
rect 857 21437 891 21471
rect 5549 21437 5583 21471
rect 5825 21437 5859 21471
rect 6101 21437 6135 21471
rect 6285 21437 6319 21471
rect 6469 21437 6503 21471
rect 6653 21437 6687 21471
rect 7297 21437 7331 21471
rect 11262 21437 11296 21471
rect 11529 21437 11563 21471
rect 12173 21437 12207 21471
rect 12541 21437 12575 21471
rect 13277 21437 13311 21471
rect 13921 21437 13955 21471
rect 14013 21437 14047 21471
rect 14565 21437 14599 21471
rect 14749 21437 14783 21471
rect 16129 21437 16163 21471
rect 20177 21437 20211 21471
rect 20453 21437 20487 21471
rect 20821 21437 20855 21471
rect 21097 21437 21131 21471
rect 21245 21437 21279 21471
rect 21603 21437 21637 21471
rect 22193 21437 22227 21471
rect 1102 21369 1136 21403
rect 3494 21369 3528 21403
rect 5089 21369 5123 21403
rect 5733 21369 5767 21403
rect 6193 21369 6227 21403
rect 7941 21369 7975 21403
rect 8769 21369 8803 21403
rect 16589 21369 16623 21403
rect 17408 21369 17442 21403
rect 18705 21369 18739 21403
rect 20545 21369 20579 21403
rect 20637 21369 20671 21403
rect 21373 21369 21407 21403
rect 21465 21369 21499 21403
rect 24970 21369 25004 21403
rect 25596 21369 25630 21403
rect 2237 21301 2271 21335
rect 2697 21301 2731 21335
rect 2881 21301 2915 21335
rect 4629 21301 4663 21335
rect 4721 21301 4755 21335
rect 4889 21301 4923 21335
rect 5365 21301 5399 21335
rect 8401 21301 8435 21335
rect 8569 21301 8603 21335
rect 13553 21301 13587 21335
rect 16313 21301 16347 21335
rect 16865 21301 16899 21335
rect 19533 21301 19567 21335
rect 21741 21301 21775 21335
rect 23121 21301 23155 21335
rect 26709 21301 26743 21335
rect 949 21097 983 21131
rect 1225 21097 1259 21131
rect 1393 21097 1427 21131
rect 14749 21097 14783 21131
rect 17417 21097 17451 21131
rect 18981 21097 19015 21131
rect 20453 21097 20487 21131
rect 21005 21097 21039 21131
rect 21281 21097 21315 21131
rect 21833 21097 21867 21131
rect 25605 21097 25639 21131
rect 1593 21029 1627 21063
rect 2605 21029 2639 21063
rect 4813 21029 4847 21063
rect 5181 21029 5215 21063
rect 5273 21029 5307 21063
rect 6929 21029 6963 21063
rect 8493 21029 8527 21063
rect 9505 21029 9539 21063
rect 11897 21029 11931 21063
rect 19318 21029 19352 21063
rect 23305 21029 23339 21063
rect 23505 21029 23539 21063
rect 26433 21029 26467 21063
rect 8723 20995 8757 21029
rect 12127 20995 12161 21029
rect 1133 20961 1167 20995
rect 2697 20961 2731 20995
rect 3249 20961 3283 20995
rect 3709 20961 3743 20995
rect 5089 20961 5123 20995
rect 5457 20961 5491 20995
rect 8134 20961 8168 20995
rect 9321 20961 9355 20995
rect 9689 20961 9723 20995
rect 10333 20961 10367 20995
rect 10517 20961 10551 20995
rect 10793 20961 10827 20995
rect 11437 20961 11471 20995
rect 12357 20961 12391 20995
rect 13001 20961 13035 20995
rect 13093 20961 13127 20995
rect 13369 20961 13403 20995
rect 13636 20961 13670 20995
rect 15209 20961 15243 20995
rect 15393 20961 15427 20995
rect 15485 20961 15519 20995
rect 16221 20961 16255 20995
rect 16405 20961 16439 20995
rect 16957 20961 16991 20995
rect 17141 20961 17175 20995
rect 17601 20961 17635 20995
rect 17693 20961 17727 20995
rect 17785 20961 17819 20995
rect 17969 20961 18003 20995
rect 18429 20961 18463 20995
rect 18613 20961 18647 20995
rect 18705 20961 18739 20995
rect 18797 20961 18831 20995
rect 20545 20961 20579 20995
rect 21741 20961 21775 20995
rect 22569 20961 22603 20995
rect 24869 20961 24903 20995
rect 25421 20961 25455 20995
rect 25605 20961 25639 20995
rect 26985 20961 27019 20995
rect 1777 20893 1811 20927
rect 3157 20893 3191 20927
rect 4169 20893 4203 20927
rect 4353 20893 4387 20927
rect 4445 20893 4479 20927
rect 4537 20893 4571 20927
rect 4629 20893 4663 20927
rect 6101 20893 6135 20927
rect 8401 20893 8435 20927
rect 10149 20893 10183 20927
rect 11529 20893 11563 20927
rect 11713 20893 11747 20927
rect 15025 20893 15059 20927
rect 17325 20893 17359 20927
rect 19073 20893 19107 20927
rect 22293 20893 22327 20927
rect 24961 20893 24995 20927
rect 2881 20825 2915 20859
rect 4905 20825 4939 20859
rect 7021 20825 7055 20859
rect 11069 20825 11103 20859
rect 12265 20825 12299 20859
rect 21373 20825 21407 20859
rect 21925 20825 21959 20859
rect 25237 20825 25271 20859
rect 1409 20757 1443 20791
rect 3985 20757 4019 20791
rect 8677 20757 8711 20791
rect 8861 20757 8895 20791
rect 10609 20757 10643 20791
rect 12081 20757 12115 20791
rect 12449 20757 12483 20791
rect 13277 20757 13311 20791
rect 16313 20757 16347 20791
rect 20637 20757 20671 20791
rect 22477 20757 22511 20791
rect 23489 20757 23523 20791
rect 23673 20757 23707 20791
rect 1869 20553 1903 20587
rect 2513 20553 2547 20587
rect 3893 20553 3927 20587
rect 4445 20553 4479 20587
rect 5089 20553 5123 20587
rect 7021 20553 7055 20587
rect 7941 20553 7975 20587
rect 8401 20553 8435 20587
rect 11345 20553 11379 20587
rect 13737 20553 13771 20587
rect 15945 20553 15979 20587
rect 23397 20553 23431 20587
rect 4721 20485 4755 20519
rect 17877 20485 17911 20519
rect 24225 20485 24259 20519
rect 2789 20417 2823 20451
rect 4077 20417 4111 20451
rect 5181 20417 5215 20451
rect 14289 20417 14323 20451
rect 17325 20417 17359 20451
rect 19349 20417 19383 20451
rect 20361 20417 20395 20451
rect 20913 20417 20947 20451
rect 21741 20417 21775 20451
rect 2145 20349 2179 20383
rect 2329 20349 2363 20383
rect 2421 20349 2455 20383
rect 2605 20349 2639 20383
rect 2697 20349 2731 20383
rect 2881 20349 2915 20383
rect 3617 20349 3651 20383
rect 4353 20349 4387 20383
rect 4537 20349 4571 20383
rect 4905 20349 4939 20383
rect 5641 20349 5675 20383
rect 7481 20349 7515 20383
rect 7757 20349 7791 20383
rect 9781 20349 9815 20383
rect 9965 20349 9999 20383
rect 10232 20349 10266 20383
rect 13553 20349 13587 20383
rect 14013 20349 14047 20383
rect 17058 20349 17092 20383
rect 17693 20349 17727 20383
rect 17877 20349 17911 20383
rect 19625 20349 19659 20383
rect 19717 20349 19751 20383
rect 19993 20349 20027 20383
rect 21189 20349 21223 20383
rect 21557 20349 21591 20383
rect 21649 20349 21683 20383
rect 21925 20349 21959 20383
rect 22017 20349 22051 20383
rect 22201 20349 22235 20383
rect 22293 20349 22327 20383
rect 22385 20349 22419 20383
rect 22569 20349 22603 20383
rect 23029 20349 23063 20383
rect 23489 20349 23523 20383
rect 23673 20349 23707 20383
rect 23949 20349 23983 20383
rect 25605 20349 25639 20383
rect 25973 20349 26007 20383
rect 2053 20281 2087 20315
rect 5886 20281 5920 20315
rect 9514 20281 9548 20315
rect 14534 20281 14568 20315
rect 19809 20281 19843 20315
rect 21281 20281 21315 20315
rect 21373 20281 21407 20315
rect 23213 20281 23247 20315
rect 25338 20281 25372 20315
rect 26801 20281 26835 20315
rect 1685 20213 1719 20247
rect 1853 20213 1887 20247
rect 2145 20213 2179 20247
rect 7573 20213 7607 20247
rect 14197 20213 14231 20247
rect 15669 20213 15703 20247
rect 18705 20213 18739 20247
rect 19441 20213 19475 20247
rect 21005 20213 21039 20247
rect 22753 20213 22787 20247
rect 23581 20213 23615 20247
rect 24133 20213 24167 20247
rect 2237 20009 2271 20043
rect 2329 20009 2363 20043
rect 4169 20009 4203 20043
rect 9045 20009 9079 20043
rect 14841 20009 14875 20043
rect 15025 20009 15059 20043
rect 15777 20009 15811 20043
rect 18705 20009 18739 20043
rect 21833 20009 21867 20043
rect 23581 20009 23615 20043
rect 24133 20009 24167 20043
rect 2513 19941 2547 19975
rect 3893 19941 3927 19975
rect 8677 19941 8711 19975
rect 12709 19941 12743 19975
rect 12909 19941 12943 19975
rect 13001 19941 13035 19975
rect 15577 19941 15611 19975
rect 19432 19941 19466 19975
rect 21465 19941 21499 19975
rect 22721 19941 22755 19975
rect 22937 19941 22971 19975
rect 23397 19941 23431 19975
rect 25338 19941 25372 19975
rect 1124 19873 1158 19907
rect 2697 19873 2731 19907
rect 2789 19873 2823 19907
rect 3341 19873 3375 19907
rect 3433 19873 3467 19907
rect 3617 19873 3651 19907
rect 3801 19873 3835 19907
rect 3985 19873 4019 19907
rect 4629 19873 4663 19907
rect 4721 19873 4755 19907
rect 4997 19873 5031 19907
rect 6184 19873 6218 19907
rect 8585 19873 8619 19907
rect 8861 19873 8895 19907
rect 9505 19873 9539 19907
rect 9689 19873 9723 19907
rect 11345 19873 11379 19907
rect 11805 19873 11839 19907
rect 12081 19873 12115 19907
rect 13921 19873 13955 19907
rect 16221 19873 16255 19907
rect 17325 19873 17359 19907
rect 17592 19873 17626 19907
rect 21281 19873 21315 19907
rect 21557 19873 21591 19907
rect 21649 19873 21683 19907
rect 22293 19873 22327 19907
rect 22477 19873 22511 19907
rect 23857 19873 23891 19907
rect 23949 19873 23983 19907
rect 857 19805 891 19839
rect 4905 19805 4939 19839
rect 5917 19805 5951 19839
rect 7757 19805 7791 19839
rect 9321 19805 9355 19839
rect 11161 19805 11195 19839
rect 11253 19805 11287 19839
rect 13553 19805 13587 19839
rect 14657 19805 14691 19839
rect 19165 19805 19199 19839
rect 25605 19805 25639 19839
rect 7297 19737 7331 19771
rect 12081 19737 12115 19771
rect 15393 19737 15427 19771
rect 20545 19737 20579 19771
rect 22385 19737 22419 19771
rect 23029 19737 23063 19771
rect 23765 19737 23799 19771
rect 24225 19737 24259 19771
rect 2973 19669 3007 19703
rect 5089 19669 5123 19703
rect 8401 19669 8435 19703
rect 11713 19669 11747 19703
rect 12541 19669 12575 19703
rect 12725 19669 12759 19703
rect 13829 19669 13863 19703
rect 14013 19669 14047 19703
rect 15025 19669 15059 19703
rect 15761 19669 15795 19703
rect 15945 19669 15979 19703
rect 16865 19669 16899 19703
rect 22569 19669 22603 19703
rect 22753 19669 22787 19703
rect 23397 19669 23431 19703
rect 1041 19465 1075 19499
rect 2421 19465 2455 19499
rect 2605 19465 2639 19499
rect 2881 19465 2915 19499
rect 4261 19465 4295 19499
rect 4445 19465 4479 19499
rect 6745 19465 6779 19499
rect 7481 19465 7515 19499
rect 7941 19465 7975 19499
rect 8769 19465 8803 19499
rect 12909 19465 12943 19499
rect 13185 19465 13219 19499
rect 15485 19465 15519 19499
rect 16221 19465 16255 19499
rect 16957 19465 16991 19499
rect 20637 19465 20671 19499
rect 2053 19397 2087 19431
rect 2697 19397 2731 19431
rect 7757 19397 7791 19431
rect 14933 19397 14967 19431
rect 3341 19329 3375 19363
rect 5641 19329 5675 19363
rect 16405 19329 16439 19363
rect 22201 19329 22235 19363
rect 1225 19261 1259 19295
rect 1777 19261 1811 19295
rect 1961 19261 1995 19295
rect 3433 19261 3467 19295
rect 3985 19261 4019 19295
rect 4905 19261 4939 19295
rect 4997 19261 5031 19295
rect 5549 19261 5583 19295
rect 5825 19261 5859 19295
rect 5917 19261 5951 19295
rect 6929 19261 6963 19295
rect 7113 19261 7147 19295
rect 7205 19261 7239 19295
rect 11529 19261 11563 19295
rect 13553 19261 13587 19295
rect 15209 19261 15243 19295
rect 15301 19261 15335 19295
rect 15577 19261 15611 19295
rect 15853 19261 15887 19295
rect 16037 19261 16071 19295
rect 16497 19261 16531 19295
rect 17141 19261 17175 19295
rect 17325 19261 17359 19295
rect 17509 19261 17543 19295
rect 18429 19261 18463 19295
rect 19165 19261 19199 19295
rect 21189 19261 21223 19295
rect 21373 19261 21407 19295
rect 22109 19261 22143 19295
rect 22385 19261 22419 19295
rect 22477 19261 22511 19295
rect 22753 19261 22787 19295
rect 23029 19261 23063 19295
rect 23581 19261 23615 19295
rect 26985 19261 27019 19295
rect 3065 19193 3099 19227
rect 5457 19193 5491 19227
rect 7297 19193 7331 19227
rect 7909 19193 7943 19227
rect 8125 19193 8159 19227
rect 8585 19193 8619 19227
rect 9505 19193 9539 19227
rect 11069 19193 11103 19227
rect 11796 19193 11830 19227
rect 13001 19193 13035 19227
rect 13798 19193 13832 19227
rect 17233 19193 17267 19227
rect 17601 19193 17635 19227
rect 19432 19193 19466 19227
rect 23397 19193 23431 19227
rect 26718 19193 26752 19227
rect 1961 19125 1995 19159
rect 2421 19125 2455 19159
rect 2855 19125 2889 19159
rect 4721 19125 4755 19159
rect 5365 19125 5399 19159
rect 7497 19125 7531 19159
rect 7665 19125 7699 19159
rect 8785 19125 8819 19159
rect 8953 19125 8987 19159
rect 13201 19125 13235 19159
rect 13369 19125 13403 19159
rect 15025 19125 15059 19159
rect 15669 19125 15703 19159
rect 20545 19125 20579 19159
rect 22017 19125 22051 19159
rect 22661 19125 22695 19159
rect 22845 19125 22879 19159
rect 23213 19125 23247 19159
rect 25605 19125 25639 19159
rect 2513 18921 2547 18955
rect 6101 18921 6135 18955
rect 7941 18921 7975 18955
rect 14381 18921 14415 18955
rect 20545 18921 20579 18955
rect 21925 18921 21959 18955
rect 25789 18921 25823 18955
rect 3626 18853 3660 18887
rect 12265 18853 12299 18887
rect 13185 18853 13219 18887
rect 13553 18853 13587 18887
rect 13737 18853 13771 18887
rect 15669 18853 15703 18887
rect 19257 18853 19291 18887
rect 21557 18853 21591 18887
rect 22293 18853 22327 18887
rect 22937 18853 22971 18887
rect 3893 18785 3927 18819
rect 5825 18785 5859 18819
rect 6009 18785 6043 18819
rect 6101 18785 6135 18819
rect 6285 18785 6319 18819
rect 7582 18785 7616 18819
rect 7849 18785 7883 18819
rect 9054 18785 9088 18819
rect 10537 18785 10571 18819
rect 10793 18785 10827 18819
rect 11253 18785 11287 18819
rect 11437 18785 11471 18819
rect 11713 18785 11747 18819
rect 12449 18785 12483 18819
rect 12633 18785 12667 18819
rect 12725 18785 12759 18819
rect 13093 18785 13127 18819
rect 13369 18785 13403 18819
rect 13645 18785 13679 18819
rect 17242 18785 17276 18819
rect 17857 18785 17891 18819
rect 21465 18785 21499 18819
rect 21649 18785 21683 18819
rect 21833 18785 21867 18819
rect 22109 18785 22143 18819
rect 22201 18785 22235 18819
rect 22477 18785 22511 18819
rect 22753 18785 22787 18819
rect 23213 18785 23247 18819
rect 25605 18785 25639 18819
rect 9321 18717 9355 18751
rect 11069 18717 11103 18751
rect 17509 18717 17543 18751
rect 17601 18717 17635 18751
rect 22569 18717 22603 18751
rect 23121 18717 23155 18751
rect 6469 18649 6503 18683
rect 11529 18649 11563 18683
rect 16129 18649 16163 18683
rect 5917 18581 5951 18615
rect 9413 18581 9447 18615
rect 18981 18581 19015 18615
rect 21281 18581 21315 18615
rect 5273 18377 5307 18411
rect 6101 18377 6135 18411
rect 7297 18377 7331 18411
rect 8585 18377 8619 18411
rect 13829 18377 13863 18411
rect 15761 18377 15795 18411
rect 16405 18377 16439 18411
rect 16681 18377 16715 18411
rect 17417 18377 17451 18411
rect 18429 18377 18463 18411
rect 20361 18377 20395 18411
rect 21189 18377 21223 18411
rect 22753 18377 22787 18411
rect 24225 18377 24259 18411
rect 25053 18377 25087 18411
rect 25329 18377 25363 18411
rect 25513 18377 25547 18411
rect 15945 18309 15979 18343
rect 21373 18309 21407 18343
rect 23121 18309 23155 18343
rect 23581 18309 23615 18343
rect 25697 18309 25731 18343
rect 4629 18241 4663 18275
rect 12173 18241 12207 18275
rect 12265 18241 12299 18275
rect 13277 18241 13311 18275
rect 15393 18241 15427 18275
rect 23213 18241 23247 18275
rect 1317 18173 1351 18207
rect 2053 18173 2087 18207
rect 2237 18173 2271 18207
rect 2513 18173 2547 18207
rect 4537 18173 4571 18207
rect 4997 18173 5031 18207
rect 5457 18173 5491 18207
rect 5550 18173 5584 18207
rect 5733 18173 5767 18207
rect 5963 18173 5997 18207
rect 6377 18173 6411 18207
rect 6469 18173 6503 18207
rect 7481 18173 7515 18207
rect 7757 18173 7791 18207
rect 8769 18173 8803 18207
rect 9045 18173 9079 18207
rect 10241 18173 10275 18207
rect 13369 18173 13403 18207
rect 14376 18173 14410 18207
rect 14565 18173 14599 18207
rect 14748 18173 14782 18207
rect 14841 18173 14875 18207
rect 15117 18173 15151 18207
rect 16497 18173 16531 18207
rect 17233 18173 17267 18207
rect 17601 18173 17635 18207
rect 17693 18173 17727 18207
rect 17785 18173 17819 18207
rect 17969 18173 18003 18207
rect 18153 18173 18187 18207
rect 18981 18173 19015 18207
rect 20913 18173 20947 18207
rect 21005 18173 21039 18207
rect 21235 18173 21269 18207
rect 21373 18173 21407 18207
rect 21649 18173 21683 18207
rect 22017 18173 22051 18207
rect 22293 18173 22327 18207
rect 23397 18173 23431 18207
rect 23857 18173 23891 18207
rect 24317 18173 24351 18207
rect 24409 18173 24443 18207
rect 24593 18173 24627 18207
rect 24869 18173 24903 18207
rect 27077 18173 27111 18207
rect 2697 18105 2731 18139
rect 4813 18105 4847 18139
rect 5825 18105 5859 18139
rect 6561 18105 6595 18139
rect 9229 18105 9263 18139
rect 9965 18105 9999 18139
rect 10508 18105 10542 18139
rect 13797 18105 13831 18139
rect 14013 18105 14047 18139
rect 14473 18105 14507 18139
rect 14933 18105 14967 18139
rect 16037 18105 16071 18139
rect 16221 18105 16255 18139
rect 19248 18105 19282 18139
rect 22477 18105 22511 18139
rect 22753 18105 22787 18139
rect 24685 18105 24719 18139
rect 25145 18105 25179 18139
rect 26810 18105 26844 18139
rect 1133 18037 1167 18071
rect 1869 18037 1903 18071
rect 2329 18037 2363 18071
rect 4905 18037 4939 18071
rect 6285 18037 6319 18071
rect 7665 18037 7699 18071
rect 8953 18037 8987 18071
rect 11621 18037 11655 18071
rect 11713 18037 11747 18071
rect 12081 18037 12115 18071
rect 13645 18037 13679 18071
rect 14197 18037 14231 18071
rect 15301 18037 15335 18071
rect 15761 18037 15795 18071
rect 17141 18037 17175 18071
rect 20729 18037 20763 18071
rect 21557 18037 21591 18071
rect 22109 18037 22143 18071
rect 22569 18037 22603 18071
rect 24041 18037 24075 18071
rect 24593 18037 24627 18071
rect 25345 18037 25379 18071
rect 2237 17833 2271 17867
rect 4445 17833 4479 17867
rect 4905 17833 4939 17867
rect 6637 17833 6671 17867
rect 8125 17833 8159 17867
rect 10057 17833 10091 17867
rect 10977 17833 11011 17867
rect 11713 17833 11747 17867
rect 13553 17833 13587 17867
rect 14473 17833 14507 17867
rect 15577 17833 15611 17867
rect 18521 17833 18555 17867
rect 21281 17833 21315 17867
rect 22845 17833 22879 17867
rect 24501 17833 24535 17867
rect 24685 17833 24719 17867
rect 25513 17833 25547 17867
rect 26065 17833 26099 17867
rect 26617 17833 26651 17867
rect 1124 17765 1158 17799
rect 4721 17765 4755 17799
rect 6837 17765 6871 17799
rect 6929 17765 6963 17799
rect 7129 17765 7163 17799
rect 14749 17765 14783 17799
rect 17877 17765 17911 17799
rect 19809 17765 19843 17799
rect 24593 17765 24627 17799
rect 857 17697 891 17731
rect 2605 17697 2639 17731
rect 4077 17697 4111 17731
rect 4353 17697 4387 17731
rect 4629 17697 4663 17731
rect 5089 17697 5123 17731
rect 5181 17697 5215 17731
rect 5457 17697 5491 17731
rect 6285 17697 6319 17731
rect 7389 17697 7423 17731
rect 9413 17697 9447 17731
rect 9965 17697 9999 17731
rect 11161 17697 11195 17731
rect 11437 17697 11471 17731
rect 11529 17697 11563 17731
rect 12440 17697 12474 17731
rect 13829 17697 13863 17731
rect 14565 17697 14599 17731
rect 14841 17697 14875 17731
rect 14933 17697 14967 17731
rect 15669 17697 15703 17731
rect 15761 17697 15795 17731
rect 15945 17697 15979 17731
rect 16313 17697 16347 17731
rect 16865 17697 16899 17731
rect 17049 17697 17083 17731
rect 17785 17697 17819 17731
rect 17969 17697 18003 17731
rect 19165 17697 19199 17731
rect 19625 17697 19659 17731
rect 19717 17697 19751 17731
rect 19993 17697 20027 17731
rect 21419 17697 21453 17731
rect 21557 17697 21591 17731
rect 21649 17697 21683 17731
rect 21777 17697 21811 17731
rect 21925 17697 21959 17731
rect 22017 17697 22051 17731
rect 22171 17697 22205 17731
rect 23958 17697 23992 17731
rect 25789 17697 25823 17731
rect 25973 17697 26007 17731
rect 26065 17697 26099 17731
rect 26249 17697 26283 17731
rect 26433 17697 26467 17731
rect 2421 17629 2455 17663
rect 2513 17629 2547 17663
rect 2697 17629 2731 17663
rect 3985 17629 4019 17663
rect 7941 17629 7975 17663
rect 8677 17629 8711 17663
rect 10149 17629 10183 17663
rect 12173 17629 12207 17663
rect 15209 17629 15243 17663
rect 24225 17629 24259 17663
rect 7297 17561 7331 17595
rect 9597 17561 9631 17595
rect 22385 17561 22419 17595
rect 24869 17561 24903 17595
rect 25145 17561 25179 17595
rect 25789 17561 25823 17595
rect 2881 17493 2915 17527
rect 3341 17493 3375 17527
rect 4261 17493 4295 17527
rect 5365 17493 5399 17527
rect 5825 17493 5859 17527
rect 6009 17493 6043 17527
rect 6469 17493 6503 17527
rect 6653 17493 6687 17527
rect 7113 17493 7147 17527
rect 9229 17493 9263 17527
rect 15117 17493 15151 17527
rect 15393 17493 15427 17527
rect 15853 17493 15887 17527
rect 17233 17493 17267 17527
rect 19441 17493 19475 17527
rect 24317 17493 24351 17527
rect 25513 17493 25547 17527
rect 25697 17493 25731 17527
rect 1317 17289 1351 17323
rect 1501 17289 1535 17323
rect 2237 17289 2271 17323
rect 2881 17289 2915 17323
rect 3065 17289 3099 17323
rect 3249 17289 3283 17323
rect 4997 17289 5031 17323
rect 5825 17289 5859 17323
rect 6837 17289 6871 17323
rect 12633 17289 12667 17323
rect 20361 17289 20395 17323
rect 21741 17289 21775 17323
rect 1869 17221 1903 17255
rect 2421 17221 2455 17255
rect 2513 17221 2547 17255
rect 15117 17221 15151 17255
rect 16313 17221 16347 17255
rect 5181 17153 5215 17187
rect 5917 17153 5951 17187
rect 11161 17153 11195 17187
rect 15761 17153 15795 17187
rect 17693 17153 17727 17187
rect 23949 17153 23983 17187
rect 4362 17085 4396 17119
rect 4629 17085 4663 17119
rect 4905 17085 4939 17119
rect 5457 17085 5491 17119
rect 5641 17085 5675 17119
rect 6469 17085 6503 17119
rect 6653 17085 6687 17119
rect 6745 17085 6779 17119
rect 8217 17085 8251 17119
rect 8769 17085 8803 17119
rect 9036 17085 9070 17119
rect 10241 17085 10275 17119
rect 11069 17085 11103 17119
rect 12817 17085 12851 17119
rect 13093 17085 13127 17119
rect 13737 17085 13771 17119
rect 17437 17085 17471 17119
rect 17969 17085 18003 17119
rect 18337 17085 18371 17119
rect 18889 17085 18923 17119
rect 21005 17085 21039 17119
rect 21465 17085 21499 17119
rect 22753 17085 22787 17119
rect 23121 17085 23155 17119
rect 23213 17085 23247 17119
rect 24041 17085 24075 17119
rect 24225 17085 24259 17119
rect 25053 17085 25087 17119
rect 25697 17085 25731 17119
rect 1501 17017 1535 17051
rect 2053 17017 2087 17051
rect 2881 17017 2915 17051
rect 7950 17017 7984 17051
rect 14004 17017 14038 17051
rect 15209 17017 15243 17051
rect 18153 17017 18187 17051
rect 18245 17017 18279 17051
rect 19134 17017 19168 17051
rect 21741 17017 21775 17051
rect 25237 17017 25271 17051
rect 25964 17017 25998 17051
rect 2253 16949 2287 16983
rect 5549 16949 5583 16983
rect 6285 16949 6319 16983
rect 10149 16949 10183 16983
rect 10333 16949 10367 16983
rect 10701 16949 10735 16983
rect 13001 16949 13035 16983
rect 18521 16949 18555 16983
rect 20269 16949 20303 16983
rect 21557 16949 21591 16983
rect 23029 16949 23063 16983
rect 24869 16949 24903 16983
rect 25421 16949 25455 16983
rect 27077 16949 27111 16983
rect 4905 16745 4939 16779
rect 5457 16745 5491 16779
rect 7481 16745 7515 16779
rect 7665 16745 7699 16779
rect 8033 16745 8067 16779
rect 9689 16745 9723 16779
rect 10241 16745 10275 16779
rect 11529 16745 11563 16779
rect 12975 16745 13009 16779
rect 14013 16745 14047 16779
rect 16497 16745 16531 16779
rect 16789 16745 16823 16779
rect 16957 16745 16991 16779
rect 17141 16745 17175 16779
rect 18705 16745 18739 16779
rect 20361 16745 20395 16779
rect 21925 16745 21959 16779
rect 22017 16745 22051 16779
rect 24133 16745 24167 16779
rect 24777 16745 24811 16779
rect 25329 16745 25363 16779
rect 25513 16745 25547 16779
rect 26065 16745 26099 16779
rect 2942 16677 2976 16711
rect 9781 16677 9815 16711
rect 13185 16677 13219 16711
rect 13277 16677 13311 16711
rect 14197 16677 14231 16711
rect 14565 16677 14599 16711
rect 16129 16677 16163 16711
rect 16313 16677 16347 16711
rect 16589 16677 16623 16711
rect 2329 16609 2363 16643
rect 2513 16609 2547 16643
rect 2605 16609 2639 16643
rect 4445 16609 4479 16643
rect 4997 16609 5031 16643
rect 6101 16609 6135 16643
rect 6368 16609 6402 16643
rect 7849 16609 7883 16643
rect 8125 16609 8159 16643
rect 10149 16609 10183 16643
rect 10333 16609 10367 16643
rect 11437 16609 11471 16643
rect 14381 16609 14415 16643
rect 14473 16609 14507 16643
rect 14749 16609 14783 16643
rect 14933 16609 14967 16643
rect 15025 16609 15059 16643
rect 15301 16609 15335 16643
rect 15577 16609 15611 16643
rect 17049 16609 17083 16643
rect 17233 16609 17267 16643
rect 17325 16609 17359 16643
rect 17592 16609 17626 16643
rect 19441 16609 19475 16643
rect 21649 16609 21683 16643
rect 21741 16609 21775 16643
rect 22201 16609 22235 16643
rect 22293 16609 22327 16643
rect 22385 16609 22419 16643
rect 22569 16609 22603 16643
rect 22753 16609 22787 16643
rect 23020 16609 23054 16643
rect 24409 16609 24443 16643
rect 24869 16609 24903 16643
rect 24961 16609 24995 16643
rect 25881 16609 25915 16643
rect 2145 16541 2179 16575
rect 2697 16541 2731 16575
rect 9873 16541 9907 16575
rect 11621 16541 11655 16575
rect 13829 16541 13863 16575
rect 15117 16541 15151 16575
rect 15853 16541 15887 16575
rect 20269 16541 20303 16575
rect 21005 16541 21039 16575
rect 21281 16541 21315 16575
rect 21373 16541 21407 16575
rect 24317 16541 24351 16575
rect 4077 16405 4111 16439
rect 4537 16405 4571 16439
rect 5089 16405 5123 16439
rect 9321 16405 9355 16439
rect 11069 16405 11103 16439
rect 12817 16405 12851 16439
rect 13001 16405 13035 16439
rect 15485 16405 15519 16439
rect 15669 16405 15703 16439
rect 15761 16405 15795 16439
rect 16773 16405 16807 16439
rect 18797 16405 18831 16439
rect 19625 16405 19659 16439
rect 25329 16405 25363 16439
rect 1409 16201 1443 16235
rect 2053 16201 2087 16235
rect 4353 16201 4387 16235
rect 13737 16201 13771 16235
rect 14197 16201 14231 16235
rect 15485 16201 15519 16235
rect 17509 16201 17543 16235
rect 22201 16201 22235 16235
rect 23029 16201 23063 16235
rect 22109 16133 22143 16167
rect 22293 16133 22327 16167
rect 3249 16065 3283 16099
rect 4721 16065 4755 16099
rect 15301 16065 15335 16099
rect 20821 16065 20855 16099
rect 21649 16065 21683 16099
rect 23581 16065 23615 16099
rect 1593 15997 1627 16031
rect 1777 15997 1811 16031
rect 2329 15997 2363 16031
rect 2513 15997 2547 16031
rect 3801 15997 3835 16031
rect 4537 15997 4571 16031
rect 5365 15997 5399 16031
rect 7113 15997 7147 16031
rect 10149 15997 10183 16031
rect 10425 15997 10459 16031
rect 11897 15997 11931 16031
rect 14105 15997 14139 16031
rect 15209 15997 15243 16031
rect 15485 15997 15519 16031
rect 15669 15997 15703 16031
rect 17693 15997 17727 16031
rect 17877 15997 17911 16031
rect 18061 15997 18095 16031
rect 19257 15997 19291 16031
rect 19524 15997 19558 16031
rect 20729 15997 20763 16031
rect 21097 15997 21131 16031
rect 21281 15997 21315 16031
rect 21373 15997 21407 16031
rect 21557 15997 21591 16031
rect 21741 15997 21775 16031
rect 21925 15997 21959 16031
rect 23857 15997 23891 16031
rect 24041 15997 24075 16031
rect 24317 15997 24351 16031
rect 24501 15997 24535 16031
rect 24593 15997 24627 16031
rect 24685 15997 24719 16031
rect 25053 15997 25087 16031
rect 2237 15929 2271 15963
rect 10670 15929 10704 15963
rect 12164 15929 12198 15963
rect 13721 15929 13755 15963
rect 13921 15929 13955 15963
rect 17785 15929 17819 15963
rect 22661 15929 22695 15963
rect 24961 15929 24995 15963
rect 25298 15929 25332 15963
rect 1869 15861 1903 15895
rect 2037 15861 2071 15895
rect 2421 15861 2455 15895
rect 4813 15861 4847 15895
rect 6561 15861 6595 15895
rect 10333 15861 10367 15895
rect 11805 15861 11839 15895
rect 13277 15861 13311 15895
rect 13553 15861 13587 15895
rect 20637 15861 20671 15895
rect 21281 15861 21315 15895
rect 24225 15861 24259 15895
rect 26433 15861 26467 15895
rect 1777 15657 1811 15691
rect 3341 15657 3375 15691
rect 6469 15657 6503 15691
rect 6561 15657 6595 15691
rect 9045 15657 9079 15691
rect 9413 15657 9447 15691
rect 11621 15657 11655 15691
rect 12449 15657 12483 15691
rect 13093 15657 13127 15691
rect 14933 15657 14967 15691
rect 19165 15657 19199 15691
rect 20637 15657 20671 15691
rect 23029 15657 23063 15691
rect 24225 15657 24259 15691
rect 24685 15657 24719 15691
rect 3862 15589 3896 15623
rect 8769 15589 8803 15623
rect 8953 15589 8987 15623
rect 12817 15589 12851 15623
rect 13461 15589 13495 15623
rect 13798 15589 13832 15623
rect 17509 15589 17543 15623
rect 18797 15589 18831 15623
rect 19502 15589 19536 15623
rect 21833 15589 21867 15623
rect 22109 15589 22143 15623
rect 22937 15589 22971 15623
rect 1409 15521 1443 15555
rect 1685 15521 1719 15555
rect 1869 15521 1903 15555
rect 2217 15521 2251 15555
rect 5273 15521 5307 15555
rect 6653 15521 6687 15555
rect 6929 15521 6963 15555
rect 7297 15521 7331 15555
rect 8309 15521 8343 15555
rect 11253 15521 11287 15555
rect 11437 15521 11471 15555
rect 12633 15521 12667 15555
rect 12909 15521 12943 15555
rect 13001 15521 13035 15555
rect 13277 15521 13311 15555
rect 13553 15521 13587 15555
rect 15577 15521 15611 15555
rect 16865 15521 16899 15555
rect 17141 15521 17175 15555
rect 17325 15521 17359 15555
rect 18613 15521 18647 15555
rect 18889 15521 18923 15555
rect 18981 15521 19015 15555
rect 19257 15521 19291 15555
rect 21557 15521 21591 15555
rect 22017 15521 22051 15555
rect 22845 15521 22879 15555
rect 23305 15521 23339 15555
rect 24133 15521 24167 15555
rect 24225 15521 24259 15555
rect 24409 15521 24443 15555
rect 24593 15521 24627 15555
rect 24777 15521 24811 15555
rect 25145 15521 25179 15555
rect 25329 15521 25363 15555
rect 1961 15453 1995 15487
rect 3617 15453 3651 15487
rect 6193 15453 6227 15487
rect 6837 15453 6871 15487
rect 9505 15453 9539 15487
rect 9597 15453 9631 15487
rect 15393 15453 15427 15487
rect 21465 15453 21499 15487
rect 21925 15453 21959 15487
rect 23581 15453 23615 15487
rect 25605 15453 25639 15487
rect 26249 15453 26283 15487
rect 26985 15453 27019 15487
rect 17141 15385 17175 15419
rect 23213 15385 23247 15419
rect 25513 15385 25547 15419
rect 1225 15317 1259 15351
rect 4997 15317 5031 15351
rect 5089 15317 5123 15351
rect 7205 15317 7239 15351
rect 7481 15317 7515 15351
rect 8493 15317 8527 15351
rect 8585 15317 8619 15351
rect 15761 15317 15795 15351
rect 17693 15317 17727 15351
rect 21281 15317 21315 15351
rect 22569 15317 22603 15351
rect 26433 15317 26467 15351
rect 2237 15113 2271 15147
rect 4077 15113 4111 15147
rect 6193 15113 6227 15147
rect 12909 15113 12943 15147
rect 23673 15113 23707 15147
rect 27077 15113 27111 15147
rect 11253 15045 11287 15079
rect 4629 14977 4663 15011
rect 4721 14977 4755 15011
rect 11345 14977 11379 15011
rect 24869 14977 24903 15011
rect 25697 14977 25731 15011
rect 857 14909 891 14943
rect 4261 14909 4295 14943
rect 4353 14909 4387 14943
rect 4813 14909 4847 14943
rect 6285 14909 6319 14943
rect 6552 14909 6586 14943
rect 7757 14909 7791 14943
rect 7941 14909 7975 14943
rect 8401 14909 8435 14943
rect 9873 14909 9907 14943
rect 10140 14909 10174 14943
rect 12265 14909 12299 14943
rect 12541 14909 12575 14943
rect 12633 14909 12667 14943
rect 12725 14909 12759 14943
rect 12909 14909 12943 14943
rect 13093 14909 13127 14943
rect 15669 14909 15703 14943
rect 17233 14909 17267 14943
rect 17877 14909 17911 14943
rect 18061 14909 18095 14943
rect 18245 14909 18279 14943
rect 18337 14909 18371 14943
rect 22293 14909 22327 14943
rect 25145 14909 25179 14943
rect 1124 14841 1158 14875
rect 5080 14841 5114 14875
rect 7849 14841 7883 14875
rect 8646 14841 8680 14875
rect 12449 14841 12483 14875
rect 15117 14841 15151 14875
rect 15301 14841 15335 14875
rect 15936 14841 15970 14875
rect 22560 14841 22594 14875
rect 24225 14841 24259 14875
rect 24961 14841 24995 14875
rect 25964 14841 25998 14875
rect 7665 14773 7699 14807
rect 9781 14773 9815 14807
rect 11989 14773 12023 14807
rect 12081 14773 12115 14807
rect 17049 14773 17083 14807
rect 17785 14773 17819 14807
rect 18521 14773 18555 14807
rect 25329 14773 25363 14807
rect 16865 14569 16899 14603
rect 22477 14569 22511 14603
rect 23581 14569 23615 14603
rect 25053 14569 25087 14603
rect 1685 14501 1719 14535
rect 1869 14501 1903 14535
rect 2697 14501 2731 14535
rect 2913 14501 2947 14535
rect 3709 14501 3743 14535
rect 5089 14501 5123 14535
rect 6193 14501 6227 14535
rect 6469 14501 6503 14535
rect 8401 14501 8435 14535
rect 11345 14501 11379 14535
rect 17417 14501 17451 14535
rect 17509 14501 17543 14535
rect 22109 14501 22143 14535
rect 25329 14501 25363 14535
rect 26065 14501 26099 14535
rect 1961 14433 1995 14467
rect 3157 14433 3191 14467
rect 3341 14433 3375 14467
rect 4813 14433 4847 14467
rect 4905 14433 4939 14467
rect 6929 14433 6963 14467
rect 7757 14433 7791 14467
rect 8861 14433 8895 14467
rect 9597 14433 9631 14467
rect 11437 14433 11471 14467
rect 11713 14433 11747 14467
rect 11805 14433 11839 14467
rect 12072 14433 12106 14467
rect 14556 14433 14590 14467
rect 17049 14433 17083 14467
rect 17141 14433 17175 14467
rect 18714 14433 18748 14467
rect 18981 14433 19015 14467
rect 19073 14433 19107 14467
rect 19329 14433 19363 14467
rect 20637 14433 20671 14467
rect 21281 14433 21315 14467
rect 22293 14433 22327 14467
rect 22937 14433 22971 14467
rect 23121 14433 23155 14467
rect 23213 14433 23247 14467
rect 23305 14433 23339 14467
rect 23929 14433 23963 14467
rect 26709 14433 26743 14467
rect 26801 14433 26835 14467
rect 26893 14433 26927 14467
rect 27077 14433 27111 14467
rect 4537 14365 4571 14399
rect 6837 14365 6871 14399
rect 8769 14365 8803 14399
rect 13829 14365 13863 14399
rect 14289 14365 14323 14399
rect 16681 14365 16715 14399
rect 23673 14365 23707 14399
rect 5825 14297 5859 14331
rect 7113 14297 7147 14331
rect 9229 14297 9263 14331
rect 9413 14297 9447 14331
rect 15669 14297 15703 14331
rect 1685 14229 1719 14263
rect 2881 14229 2915 14263
rect 3065 14229 3099 14263
rect 3157 14229 3191 14263
rect 3525 14229 3559 14263
rect 6193 14229 6227 14263
rect 6377 14229 6411 14263
rect 6837 14229 6871 14263
rect 13185 14229 13219 14263
rect 13277 14229 13311 14263
rect 16129 14229 16163 14263
rect 17601 14229 17635 14263
rect 20453 14229 20487 14263
rect 20729 14229 20763 14263
rect 21097 14229 21131 14263
rect 26433 14229 26467 14263
rect 2237 14025 2271 14059
rect 3249 14025 3283 14059
rect 12173 14025 12207 14059
rect 12909 14025 12943 14059
rect 14749 14025 14783 14059
rect 15485 14025 15519 14059
rect 18061 14025 18095 14059
rect 19349 14025 19383 14059
rect 19625 14025 19659 14059
rect 20085 14025 20119 14059
rect 20729 14025 20763 14059
rect 21741 14025 21775 14059
rect 24777 14025 24811 14059
rect 8585 13957 8619 13991
rect 12725 13957 12759 13991
rect 13369 13957 13403 13991
rect 15301 13957 15335 13991
rect 19441 13957 19475 13991
rect 20545 13957 20579 13991
rect 21557 13957 21591 13991
rect 23213 13957 23247 13991
rect 11161 13889 11195 13923
rect 14565 13889 14599 13923
rect 21281 13889 21315 13923
rect 21833 13889 21867 13923
rect 24409 13889 24443 13923
rect 857 13821 891 13855
rect 2973 13821 3007 13855
rect 4629 13821 4663 13855
rect 5089 13821 5123 13855
rect 5273 13821 5307 13855
rect 6561 13821 6595 13855
rect 6745 13821 6779 13855
rect 8217 13821 8251 13855
rect 8401 13821 8435 13855
rect 8769 13821 8803 13855
rect 11069 13821 11103 13855
rect 11345 13821 11379 13855
rect 12357 13821 12391 13855
rect 12633 13821 12667 13855
rect 13185 13821 13219 13855
rect 13369 13821 13403 13855
rect 13737 13821 13771 13855
rect 14933 13821 14967 13855
rect 15209 13821 15243 13855
rect 16773 13821 16807 13855
rect 17141 13821 17175 13855
rect 17325 13821 17359 13855
rect 17417 13821 17451 13855
rect 18245 13821 18279 13855
rect 18521 13821 18555 13855
rect 18705 13821 18739 13855
rect 19993 13821 20027 13855
rect 20361 13821 20395 13855
rect 20913 13821 20947 13855
rect 23489 13821 23523 13855
rect 24777 13821 24811 13855
rect 24869 13821 24903 13855
rect 25053 13821 25087 13855
rect 25513 13821 25547 13855
rect 25780 13821 25814 13855
rect 1124 13753 1158 13787
rect 4362 13753 4396 13787
rect 10802 13753 10836 13787
rect 11529 13753 11563 13787
rect 13093 13753 13127 13787
rect 15669 13753 15703 13787
rect 18429 13753 18463 13787
rect 19809 13753 19843 13787
rect 22100 13753 22134 13787
rect 23673 13753 23707 13787
rect 2329 13685 2363 13719
rect 4905 13685 4939 13719
rect 6653 13685 6687 13719
rect 8033 13685 8067 13719
rect 8953 13685 8987 13719
rect 9689 13685 9723 13719
rect 12541 13685 12575 13719
rect 12893 13685 12927 13719
rect 15117 13685 15151 13719
rect 15459 13685 15493 13719
rect 16221 13685 16255 13719
rect 16957 13685 16991 13719
rect 19599 13685 19633 13719
rect 23305 13685 23339 13719
rect 23857 13685 23891 13719
rect 24593 13685 24627 13719
rect 26893 13685 26927 13719
rect 1317 13481 1351 13515
rect 3341 13481 3375 13515
rect 3709 13481 3743 13515
rect 6101 13481 6135 13515
rect 7849 13481 7883 13515
rect 14105 13481 14139 13515
rect 14365 13481 14399 13515
rect 18705 13481 18739 13515
rect 18873 13481 18907 13515
rect 20821 13481 20855 13515
rect 21281 13481 21315 13515
rect 22017 13481 22051 13515
rect 26433 13481 26467 13515
rect 2697 13413 2731 13447
rect 2973 13413 3007 13447
rect 3985 13413 4019 13447
rect 4414 13413 4448 13447
rect 9781 13413 9815 13447
rect 13737 13413 13771 13447
rect 13921 13413 13955 13447
rect 14565 13413 14599 13447
rect 15853 13413 15887 13447
rect 16672 13413 16706 13447
rect 19073 13413 19107 13447
rect 20484 13413 20518 13447
rect 21741 13413 21775 13447
rect 3157 13345 3191 13379
rect 3433 13345 3467 13379
rect 3525 13345 3559 13379
rect 3893 13345 3927 13379
rect 4077 13345 4111 13379
rect 6285 13345 6319 13379
rect 6377 13345 6411 13379
rect 6736 13345 6770 13379
rect 7941 13345 7975 13379
rect 8208 13345 8242 13379
rect 9413 13345 9447 13379
rect 9597 13345 9631 13379
rect 9873 13345 9907 13379
rect 9965 13345 9999 13379
rect 10977 13345 11011 13379
rect 11161 13345 11195 13379
rect 15669 13345 15703 13379
rect 15945 13345 15979 13379
rect 21005 13345 21039 13379
rect 21281 13345 21315 13379
rect 21465 13345 21499 13379
rect 21557 13345 21591 13379
rect 23029 13345 23063 13379
rect 23121 13345 23155 13379
rect 23213 13345 23247 13379
rect 23397 13345 23431 13379
rect 23489 13345 23523 13379
rect 23673 13345 23707 13379
rect 23765 13345 23799 13379
rect 23857 13345 23891 13379
rect 25881 13345 25915 13379
rect 26157 13345 26191 13379
rect 26985 13345 27019 13379
rect 1869 13277 1903 13311
rect 4169 13277 4203 13311
rect 6101 13277 6135 13311
rect 6469 13277 6503 13311
rect 13277 13277 13311 13311
rect 15393 13277 15427 13311
rect 16405 13277 16439 13311
rect 17969 13277 18003 13311
rect 20729 13277 20763 13311
rect 22661 13277 22695 13311
rect 22753 13277 22787 13311
rect 24869 13277 24903 13311
rect 25513 13277 25547 13311
rect 26065 13277 26099 13311
rect 2329 13209 2363 13243
rect 2881 13209 2915 13243
rect 17785 13209 17819 13243
rect 18613 13209 18647 13243
rect 19349 13209 19383 13243
rect 21925 13209 21959 13243
rect 24133 13209 24167 13243
rect 2697 13141 2731 13175
rect 5549 13141 5583 13175
rect 9321 13141 9355 13175
rect 10609 13141 10643 13175
rect 11161 13141 11195 13175
rect 12725 13141 12759 13175
rect 14197 13141 14231 13175
rect 14381 13141 14415 13175
rect 14749 13141 14783 13175
rect 15485 13141 15519 13175
rect 18889 13141 18923 13175
rect 24225 13141 24259 13175
rect 24961 13141 24995 13175
rect 25697 13141 25731 13175
rect 26157 13141 26191 13175
rect 1409 12937 1443 12971
rect 4813 12937 4847 12971
rect 6745 12937 6779 12971
rect 8953 12937 8987 12971
rect 9229 12937 9263 12971
rect 10425 12937 10459 12971
rect 10701 12937 10735 12971
rect 12817 12937 12851 12971
rect 16589 12937 16623 12971
rect 20361 12937 20395 12971
rect 22845 12937 22879 12971
rect 23857 12937 23891 12971
rect 27077 12937 27111 12971
rect 1961 12869 1995 12903
rect 6929 12869 6963 12903
rect 9137 12869 9171 12903
rect 12541 12869 12575 12903
rect 22109 12869 22143 12903
rect 1777 12801 1811 12835
rect 1869 12801 1903 12835
rect 4537 12801 4571 12835
rect 4905 12801 4939 12835
rect 5549 12801 5583 12835
rect 6193 12801 6227 12835
rect 7113 12801 7147 12835
rect 9781 12801 9815 12835
rect 18705 12801 18739 12835
rect 20729 12801 20763 12835
rect 23581 12801 23615 12835
rect 25237 12801 25271 12835
rect 25697 12801 25731 12835
rect 1593 12733 1627 12767
rect 1961 12733 1995 12767
rect 2237 12733 2271 12767
rect 2789 12733 2823 12767
rect 3433 12733 3467 12767
rect 3709 12733 3743 12767
rect 4353 12733 4387 12767
rect 4445 12733 4479 12767
rect 4629 12733 4663 12767
rect 5089 12733 5123 12767
rect 6377 12733 6411 12767
rect 6561 12733 6595 12767
rect 6837 12733 6871 12767
rect 9965 12733 9999 12767
rect 10241 12733 10275 12767
rect 11161 12733 11195 12767
rect 13093 12733 13127 12767
rect 13277 12733 13311 12767
rect 13553 12733 13587 12767
rect 15209 12733 15243 12767
rect 17601 12733 17635 12767
rect 17693 12733 17727 12767
rect 18521 12733 18555 12767
rect 20177 12733 20211 12767
rect 20361 12733 20395 12767
rect 22477 12733 22511 12767
rect 22937 12733 22971 12767
rect 23029 12733 23063 12767
rect 24970 12733 25004 12767
rect 3617 12665 3651 12699
rect 4813 12665 4847 12699
rect 8769 12665 8803 12699
rect 10885 12665 10919 12699
rect 11428 12665 11462 12699
rect 12785 12665 12819 12699
rect 13001 12665 13035 12699
rect 13820 12665 13854 12699
rect 15476 12665 15510 12699
rect 17969 12665 18003 12699
rect 18061 12665 18095 12699
rect 18429 12665 18463 12699
rect 18972 12665 19006 12699
rect 20996 12665 21030 12699
rect 22201 12665 22235 12699
rect 22569 12665 22603 12699
rect 25942 12665 25976 12699
rect 2145 12597 2179 12631
rect 2605 12597 2639 12631
rect 3249 12597 3283 12631
rect 4169 12597 4203 12631
rect 5273 12597 5307 12631
rect 7113 12597 7147 12631
rect 8979 12597 9013 12631
rect 10057 12597 10091 12631
rect 10517 12597 10551 12631
rect 10685 12597 10719 12631
rect 12633 12597 12667 12631
rect 13185 12597 13219 12631
rect 14933 12597 14967 12631
rect 17417 12597 17451 12631
rect 20085 12597 20119 12631
rect 22661 12597 22695 12631
rect 3709 12393 3743 12427
rect 10977 12393 11011 12427
rect 11529 12393 11563 12427
rect 11897 12393 11931 12427
rect 13461 12393 13495 12427
rect 13829 12393 13863 12427
rect 15669 12393 15703 12427
rect 19257 12393 19291 12427
rect 21465 12393 21499 12427
rect 22477 12393 22511 12427
rect 23397 12393 23431 12427
rect 23857 12393 23891 12427
rect 25237 12393 25271 12427
rect 26433 12393 26467 12427
rect 2596 12325 2630 12359
rect 9260 12325 9294 12359
rect 9597 12325 9631 12359
rect 9797 12325 9831 12359
rect 14841 12325 14875 12359
rect 18889 12325 18923 12359
rect 23213 12325 23247 12359
rect 24041 12325 24075 12359
rect 857 12257 891 12291
rect 1124 12257 1158 12291
rect 2329 12257 2363 12291
rect 4261 12257 4295 12291
rect 4537 12257 4571 12291
rect 4721 12257 4755 12291
rect 4905 12257 4939 12291
rect 5825 12257 5859 12291
rect 6081 12257 6115 12291
rect 9505 12257 9539 12291
rect 11161 12257 11195 12291
rect 11345 12257 11379 12291
rect 11437 12257 11471 12291
rect 11713 12257 11747 12291
rect 11989 12257 12023 12291
rect 12348 12257 12382 12291
rect 14013 12257 14047 12291
rect 14197 12257 14231 12291
rect 14289 12257 14323 12291
rect 15945 12257 15979 12291
rect 18797 12257 18831 12291
rect 19073 12257 19107 12291
rect 21833 12257 21867 12291
rect 21925 12257 21959 12291
rect 22753 12257 22787 12291
rect 22937 12257 22971 12291
rect 23029 12257 23063 12291
rect 23581 12257 23615 12291
rect 24225 12257 24259 12291
rect 25605 12257 25639 12291
rect 25697 12257 25731 12291
rect 25789 12257 25823 12291
rect 25973 12257 26007 12291
rect 26709 12257 26743 12291
rect 26801 12257 26835 12291
rect 26893 12257 26927 12291
rect 27077 12257 27111 12291
rect 5457 12189 5491 12223
rect 7849 12189 7883 12223
rect 10609 12189 10643 12223
rect 12081 12189 12115 12223
rect 15669 12189 15703 12223
rect 15853 12189 15887 12223
rect 18061 12189 18095 12223
rect 20269 12189 20303 12223
rect 21741 12189 21775 12223
rect 22201 12189 22235 12223
rect 24685 12189 24719 12223
rect 25329 12189 25363 12223
rect 7297 12121 7331 12155
rect 10057 12121 10091 12155
rect 14657 12121 14691 12155
rect 2237 12053 2271 12087
rect 4077 12053 4111 12087
rect 7205 12053 7239 12087
rect 8125 12053 8159 12087
rect 9781 12053 9815 12087
rect 9965 12053 9999 12087
rect 18705 12053 18739 12087
rect 19717 12053 19751 12087
rect 21833 12053 21867 12087
rect 22293 12053 22327 12087
rect 22569 12053 22603 12087
rect 23673 12053 23707 12087
rect 1317 11849 1351 11883
rect 3433 11849 3467 11883
rect 5089 11849 5123 11883
rect 5641 11849 5675 11883
rect 7205 11849 7239 11883
rect 7481 11849 7515 11883
rect 9597 11849 9631 11883
rect 12173 11849 12207 11883
rect 12909 11849 12943 11883
rect 14473 11849 14507 11883
rect 16129 11849 16163 11883
rect 17877 11849 17911 11883
rect 18153 11849 18187 11883
rect 18981 11849 19015 11883
rect 19165 11849 19199 11883
rect 21833 11849 21867 11883
rect 22293 11849 22327 11883
rect 27077 11849 27111 11883
rect 3249 11781 3283 11815
rect 20913 11781 20947 11815
rect 2605 11713 2639 11747
rect 10977 11713 11011 11747
rect 14749 11713 14783 11747
rect 16497 11713 16531 11747
rect 20729 11713 20763 11747
rect 25697 11713 25731 11747
rect 1869 11645 1903 11679
rect 3709 11645 3743 11679
rect 5457 11645 5491 11679
rect 5641 11645 5675 11679
rect 6285 11645 6319 11679
rect 6837 11645 6871 11679
rect 7481 11645 7515 11679
rect 7573 11645 7607 11679
rect 7757 11645 7791 11679
rect 8493 11645 8527 11679
rect 8677 11645 8711 11679
rect 12357 11645 12391 11679
rect 12633 11645 12667 11679
rect 19717 11645 19751 11679
rect 19993 11645 20027 11679
rect 21005 11645 21039 11679
rect 21741 11645 21775 11679
rect 21833 11645 21867 11679
rect 22385 11645 22419 11679
rect 22569 11645 22603 11679
rect 22661 11645 22695 11679
rect 22753 11645 22787 11679
rect 23857 11645 23891 11679
rect 24409 11645 24443 11679
rect 24869 11645 24903 11679
rect 24961 11645 24995 11679
rect 25145 11645 25179 11679
rect 25237 11645 25271 11679
rect 25329 11645 25363 11679
rect 3617 11577 3651 11611
rect 3976 11577 4010 11611
rect 7173 11577 7207 11611
rect 7389 11577 7423 11611
rect 10710 11577 10744 11611
rect 12893 11577 12927 11611
rect 13093 11577 13127 11611
rect 14289 11577 14323 11611
rect 15016 11577 15050 11611
rect 16764 11577 16798 11611
rect 18337 11577 18371 11611
rect 19349 11577 19383 11611
rect 21557 11577 21591 11611
rect 21925 11577 21959 11611
rect 22109 11577 22143 11611
rect 23213 11577 23247 11611
rect 23397 11577 23431 11611
rect 25605 11577 25639 11611
rect 25942 11577 25976 11611
rect 2053 11509 2087 11543
rect 3417 11509 3451 11543
rect 7021 11509 7055 11543
rect 9505 11509 9539 11543
rect 12541 11509 12575 11543
rect 12725 11509 12759 11543
rect 14489 11509 14523 11543
rect 14657 11509 14691 11543
rect 17969 11509 18003 11543
rect 18137 11509 18171 11543
rect 19139 11509 19173 11543
rect 19625 11509 19659 11543
rect 20637 11509 20671 11543
rect 20729 11509 20763 11543
rect 23029 11509 23063 11543
rect 23581 11509 23615 11543
rect 24685 11509 24719 11543
rect 1409 11305 1443 11339
rect 2605 11305 2639 11339
rect 6745 11305 6779 11339
rect 9413 11305 9447 11339
rect 10425 11305 10459 11339
rect 14565 11305 14599 11339
rect 15393 11305 15427 11339
rect 15761 11305 15795 11339
rect 16957 11305 16991 11339
rect 19717 11305 19751 11339
rect 22477 11305 22511 11339
rect 26433 11305 26467 11339
rect 6561 11237 6595 11271
rect 9045 11237 9079 11271
rect 9245 11237 9279 11271
rect 10057 11237 10091 11271
rect 17325 11237 17359 11271
rect 19625 11237 19659 11271
rect 20830 11237 20864 11271
rect 22836 11237 22870 11271
rect 25176 11237 25210 11271
rect 25513 11237 25547 11271
rect 1593 11169 1627 11203
rect 1869 11169 1903 11203
rect 2973 11169 3007 11203
rect 6377 11169 6411 11203
rect 6929 11169 6963 11203
rect 7021 11169 7055 11203
rect 7297 11169 7331 11203
rect 9505 11169 9539 11203
rect 9689 11169 9723 11203
rect 9965 11169 9999 11203
rect 10241 11169 10275 11203
rect 11069 11169 11103 11203
rect 11336 11169 11370 11203
rect 13185 11169 13219 11203
rect 13452 11169 13486 11203
rect 15577 11169 15611 11203
rect 15853 11169 15887 11203
rect 16129 11169 16163 11203
rect 16313 11169 16347 11203
rect 17141 11169 17175 11203
rect 17417 11169 17451 11203
rect 17693 11169 17727 11203
rect 19145 11169 19179 11203
rect 19257 11169 19291 11203
rect 21097 11169 21131 11203
rect 22569 11169 22603 11203
rect 27077 11169 27111 11203
rect 1777 11101 1811 11135
rect 6745 11101 6779 11135
rect 7205 11101 7239 11135
rect 9597 11101 9631 11135
rect 15301 11101 15335 11135
rect 19533 11101 19567 11135
rect 21925 11101 21959 11135
rect 25421 11101 25455 11135
rect 26065 11101 26099 11135
rect 2421 11033 2455 11067
rect 7665 11033 7699 11067
rect 18981 11033 19015 11067
rect 24041 11033 24075 11067
rect 2605 10965 2639 10999
rect 6193 10965 6227 10999
rect 9229 10965 9263 10999
rect 12449 10965 12483 10999
rect 14657 10965 14691 10999
rect 16129 10965 16163 10999
rect 17601 10965 17635 10999
rect 23949 10965 23983 10999
rect 3525 10761 3559 10795
rect 5365 10761 5399 10795
rect 13645 10761 13679 10795
rect 14381 10761 14415 10795
rect 16221 10761 16255 10795
rect 16497 10761 16531 10795
rect 20085 10761 20119 10795
rect 20177 10761 20211 10795
rect 25421 10761 25455 10795
rect 26893 10761 26927 10795
rect 6009 10693 6043 10727
rect 20637 10693 20671 10727
rect 5641 10625 5675 10659
rect 6193 10625 6227 10659
rect 7021 10625 7055 10659
rect 12909 10625 12943 10659
rect 17417 10625 17451 10659
rect 18705 10625 18739 10659
rect 22109 10625 22143 10659
rect 2513 10557 2547 10591
rect 2789 10557 2823 10591
rect 3249 10557 3283 10591
rect 3985 10557 4019 10591
rect 4169 10557 4203 10591
rect 4261 10557 4295 10591
rect 4813 10557 4847 10591
rect 5825 10557 5859 10591
rect 6101 10557 6135 10591
rect 6653 10557 6687 10591
rect 7113 10557 7147 10591
rect 8953 10557 8987 10591
rect 9045 10557 9079 10591
rect 9229 10557 9263 10591
rect 9321 10557 9355 10591
rect 9413 10557 9447 10591
rect 9597 10557 9631 10591
rect 10333 10557 10367 10591
rect 10609 10557 10643 10591
rect 10885 10557 10919 10591
rect 11713 10557 11747 10591
rect 11897 10557 11931 10591
rect 11989 10557 12023 10591
rect 12173 10557 12207 10591
rect 12277 10557 12311 10591
rect 13093 10557 13127 10591
rect 13277 10557 13311 10591
rect 13829 10557 13863 10591
rect 14013 10557 14047 10591
rect 14105 10557 14139 10591
rect 15577 10557 15611 10591
rect 15669 10557 15703 10591
rect 15853 10557 15887 10591
rect 15945 10557 15979 10591
rect 17049 10557 17083 10591
rect 17509 10557 17543 10591
rect 17877 10557 17911 10591
rect 18153 10557 18187 10591
rect 18337 10557 18371 10591
rect 18429 10557 18463 10591
rect 20361 10557 20395 10591
rect 20453 10557 20487 10591
rect 22017 10557 22051 10591
rect 22753 10557 22787 10591
rect 23121 10557 23155 10591
rect 23213 10557 23247 10591
rect 23305 10557 23339 10591
rect 23489 10557 23523 10591
rect 24225 10557 24259 10591
rect 25145 10557 25179 10591
rect 25237 10557 25271 10591
rect 25513 10557 25547 10591
rect 3525 10489 3559 10523
rect 5349 10489 5383 10523
rect 5549 10489 5583 10523
rect 6561 10489 6595 10523
rect 13185 10489 13219 10523
rect 14565 10489 14599 10523
rect 16037 10489 16071 10523
rect 17785 10489 17819 10523
rect 18950 10489 18984 10523
rect 20177 10489 20211 10523
rect 21772 10489 21806 10523
rect 22845 10489 22879 10523
rect 25421 10489 25455 10523
rect 25758 10489 25792 10523
rect 2605 10421 2639 10455
rect 2973 10421 3007 10455
rect 3341 10421 3375 10455
rect 3985 10421 4019 10455
rect 5181 10421 5215 10455
rect 6469 10421 6503 10455
rect 7481 10421 7515 10455
rect 8769 10421 8803 10455
rect 9505 10421 9539 10455
rect 10149 10421 10183 10455
rect 10517 10421 10551 10455
rect 11529 10421 11563 10455
rect 12357 10421 12391 10455
rect 14197 10421 14231 10455
rect 14365 10421 14399 10455
rect 15393 10421 15427 10455
rect 16237 10421 16271 10455
rect 16405 10421 16439 10455
rect 17233 10421 17267 10455
rect 17969 10421 18003 10455
rect 24869 10421 24903 10455
rect 24961 10421 24995 10455
rect 4169 10217 4203 10251
rect 7021 10217 7055 10251
rect 10977 10217 11011 10251
rect 11529 10217 11563 10251
rect 11897 10217 11931 10251
rect 16405 10217 16439 10251
rect 18781 10217 18815 10251
rect 22017 10217 22051 10251
rect 26433 10217 26467 10251
rect 3056 10149 3090 10183
rect 7297 10149 7331 10183
rect 9680 10149 9714 10183
rect 11129 10149 11163 10183
rect 11345 10149 11379 10183
rect 12249 10149 12283 10183
rect 12449 10149 12483 10183
rect 17540 10149 17574 10183
rect 18981 10149 19015 10183
rect 21649 10149 21683 10183
rect 21833 10149 21867 10183
rect 25789 10149 25823 10183
rect 25973 10149 26007 10183
rect 2421 10081 2455 10115
rect 2789 10081 2823 10115
rect 4528 10081 4562 10115
rect 6285 10081 6319 10115
rect 6929 10081 6963 10115
rect 7113 10081 7147 10115
rect 7389 10081 7423 10115
rect 7481 10081 7515 10115
rect 8585 10081 8619 10115
rect 8677 10081 8711 10115
rect 8861 10081 8895 10115
rect 8953 10081 8987 10115
rect 9137 10081 9171 10115
rect 9321 10081 9355 10115
rect 11713 10081 11747 10115
rect 11989 10081 12023 10115
rect 13001 10081 13035 10115
rect 13185 10081 13219 10115
rect 14657 10081 14691 10115
rect 14749 10081 14783 10115
rect 14933 10081 14967 10115
rect 15025 10081 15059 10115
rect 16129 10081 16163 10115
rect 16221 10081 16255 10115
rect 16313 10081 16347 10115
rect 18061 10081 18095 10115
rect 18153 10081 18187 10115
rect 18337 10081 18371 10115
rect 20085 10081 20119 10115
rect 22385 10081 22419 10115
rect 22477 10081 22511 10115
rect 22569 10081 22603 10115
rect 22753 10081 22787 10115
rect 22845 10081 22879 10115
rect 23029 10081 23063 10115
rect 23121 10081 23155 10115
rect 23213 10081 23247 10115
rect 24317 10081 24351 10115
rect 24501 10081 24535 10115
rect 24593 10081 24627 10115
rect 24685 10081 24719 10115
rect 26157 10081 26191 10115
rect 26985 10081 27019 10115
rect 2237 10013 2271 10047
rect 2329 10013 2363 10047
rect 2513 10013 2547 10047
rect 4261 10013 4295 10047
rect 8033 10013 8067 10047
rect 9413 10013 9447 10047
rect 15669 10013 15703 10047
rect 17785 10013 17819 10047
rect 18521 10013 18555 10047
rect 23489 10013 23523 10047
rect 23581 10013 23615 10047
rect 25053 10013 25087 10047
rect 25605 10013 25639 10047
rect 5641 9945 5675 9979
rect 12081 9945 12115 9979
rect 18613 9945 18647 9979
rect 24961 9945 24995 9979
rect 2697 9877 2731 9911
rect 6837 9877 6871 9911
rect 8401 9877 8435 9911
rect 9321 9877 9355 9911
rect 10793 9877 10827 9911
rect 11161 9877 11195 9911
rect 12265 9877 12299 9911
rect 13001 9877 13035 9911
rect 14473 9877 14507 9911
rect 15117 9877 15151 9911
rect 18797 9877 18831 9911
rect 19441 9877 19475 9911
rect 22109 9877 22143 9911
rect 24225 9877 24259 9911
rect 3249 9673 3283 9707
rect 4905 9673 4939 9707
rect 7665 9673 7699 9707
rect 15209 9673 15243 9707
rect 22477 9673 22511 9707
rect 23673 9673 23707 9707
rect 25513 9673 25547 9707
rect 2973 9605 3007 9639
rect 14933 9605 14967 9639
rect 22385 9605 22419 9639
rect 27077 9605 27111 9639
rect 2605 9537 2639 9571
rect 3065 9537 3099 9571
rect 7297 9537 7331 9571
rect 23029 9537 23063 9571
rect 23581 9537 23615 9571
rect 2145 9469 2179 9503
rect 3433 9469 3467 9503
rect 3985 9469 4019 9503
rect 4169 9469 4203 9503
rect 4261 9469 4295 9503
rect 4629 9469 4663 9503
rect 5089 9469 5123 9503
rect 7849 9469 7883 9503
rect 7941 9469 7975 9503
rect 8125 9469 8159 9503
rect 8217 9469 8251 9503
rect 8769 9469 8803 9503
rect 9045 9469 9079 9503
rect 9229 9469 9263 9503
rect 9597 9469 9631 9503
rect 9689 9469 9723 9503
rect 9873 9469 9907 9503
rect 11529 9469 11563 9503
rect 11805 9469 11839 9503
rect 12173 9469 12207 9503
rect 12265 9469 12299 9503
rect 12449 9469 12483 9503
rect 12541 9469 12575 9503
rect 12909 9469 12943 9503
rect 13001 9469 13035 9503
rect 13185 9469 13219 9503
rect 13277 9469 13311 9503
rect 13553 9469 13587 9503
rect 15761 9469 15795 9503
rect 15853 9469 15887 9503
rect 16037 9469 16071 9503
rect 16129 9469 16163 9503
rect 16221 9469 16255 9503
rect 16405 9469 16439 9503
rect 16497 9469 16531 9503
rect 16681 9469 16715 9503
rect 18705 9469 18739 9503
rect 18889 9469 18923 9503
rect 20545 9469 20579 9503
rect 21005 9469 21039 9503
rect 21272 9469 21306 9503
rect 23397 9469 23431 9503
rect 23857 9469 23891 9503
rect 24593 9469 24627 9503
rect 24869 9469 24903 9503
rect 25053 9469 25087 9503
rect 25145 9469 25179 9503
rect 25237 9469 25271 9503
rect 25697 9469 25731 9503
rect 1961 9401 1995 9435
rect 4077 9401 4111 9435
rect 4445 9401 4479 9435
rect 7030 9401 7064 9435
rect 9781 9401 9815 9435
rect 13820 9401 13854 9435
rect 15177 9401 15211 9435
rect 15393 9401 15427 9435
rect 16313 9401 16347 9435
rect 20278 9401 20312 9435
rect 23673 9401 23707 9435
rect 25942 9401 25976 9435
rect 2329 9333 2363 9367
rect 5917 9333 5951 9367
rect 8861 9333 8895 9367
rect 11345 9333 11379 9367
rect 11713 9333 11747 9367
rect 11989 9333 12023 9367
rect 12725 9333 12759 9367
rect 15025 9333 15059 9367
rect 15577 9333 15611 9367
rect 16589 9333 16623 9367
rect 18797 9333 18831 9367
rect 19165 9333 19199 9367
rect 23213 9333 23247 9367
rect 7665 9129 7699 9163
rect 13921 9129 13955 9163
rect 19533 9129 19567 9163
rect 19993 9129 20027 9163
rect 22661 9129 22695 9163
rect 25605 9129 25639 9163
rect 2681 9061 2715 9095
rect 2881 9061 2915 9095
rect 3525 9061 3559 9095
rect 11244 9061 11278 9095
rect 26433 9061 26467 9095
rect 857 8993 891 9027
rect 1124 8993 1158 9027
rect 3160 8993 3194 9027
rect 3433 8993 3467 9027
rect 3617 8993 3651 9027
rect 7297 8993 7331 9027
rect 8769 8993 8803 9027
rect 8861 8993 8895 9027
rect 9045 8993 9079 9027
rect 9137 8993 9171 9027
rect 10241 8993 10275 9027
rect 10425 8993 10459 9027
rect 12725 8993 12759 9027
rect 12817 8993 12851 9027
rect 13001 8993 13035 9027
rect 13093 8993 13127 9027
rect 14105 8993 14139 9027
rect 14289 8993 14323 9027
rect 14381 8993 14415 9027
rect 15577 8993 15611 9027
rect 15669 8993 15703 9027
rect 15853 8993 15887 9027
rect 15945 8993 15979 9027
rect 17316 8993 17350 9027
rect 19533 8993 19567 9027
rect 20177 8993 20211 9027
rect 20453 8993 20487 9027
rect 20821 8993 20855 9027
rect 21741 8993 21775 9027
rect 23774 8993 23808 9027
rect 24133 8993 24167 9027
rect 24317 8993 24351 9027
rect 24409 8993 24443 9027
rect 24501 8993 24535 9027
rect 25881 8993 25915 9027
rect 25973 8993 26007 9027
rect 26065 8993 26099 9027
rect 26249 8993 26283 9027
rect 26985 8993 27019 9027
rect 2973 8925 3007 8959
rect 7205 8925 7239 8959
rect 10977 8925 11011 8959
rect 17049 8925 17083 8959
rect 19165 8925 19199 8959
rect 19349 8925 19383 8959
rect 19901 8925 19935 8959
rect 20269 8925 20303 8959
rect 20637 8925 20671 8959
rect 21005 8925 21039 8959
rect 24041 8925 24075 8959
rect 24777 8925 24811 8959
rect 24869 8925 24903 8959
rect 18429 8857 18463 8891
rect 20361 8857 20395 8891
rect 2237 8789 2271 8823
rect 2513 8789 2547 8823
rect 2697 8789 2731 8823
rect 3341 8789 3375 8823
rect 8585 8789 8619 8823
rect 10333 8789 10367 8823
rect 12357 8789 12391 8823
rect 12541 8789 12575 8823
rect 15393 8789 15427 8823
rect 18613 8789 18647 8823
rect 21925 8789 21959 8823
rect 25513 8789 25547 8823
rect 1133 8585 1167 8619
rect 2145 8585 2179 8619
rect 2789 8585 2823 8619
rect 4813 8585 4847 8619
rect 11713 8585 11747 8619
rect 11897 8585 11931 8619
rect 12173 8585 12207 8619
rect 12909 8585 12943 8619
rect 14197 8585 14231 8619
rect 17509 8585 17543 8619
rect 18797 8585 18831 8619
rect 19533 8585 19567 8619
rect 20545 8585 20579 8619
rect 23213 8585 23247 8619
rect 2421 8517 2455 8551
rect 6285 8517 6319 8551
rect 15485 8517 15519 8551
rect 18061 8517 18095 8551
rect 9137 8449 9171 8483
rect 11253 8449 11287 8483
rect 17877 8449 17911 8483
rect 19717 8449 19751 8483
rect 1317 8381 1351 8415
rect 1961 8381 1995 8415
rect 2145 8381 2179 8415
rect 2789 8381 2823 8415
rect 3065 8381 3099 8415
rect 3433 8381 3467 8415
rect 4905 8381 4939 8415
rect 7113 8381 7147 8415
rect 9505 8381 9539 8415
rect 9689 8381 9723 8415
rect 9873 8381 9907 8415
rect 12725 8381 12759 8415
rect 12909 8381 12943 8415
rect 13093 8381 13127 8415
rect 15301 8381 15335 8415
rect 15393 8383 15427 8417
rect 15577 8381 15611 8415
rect 16497 8381 16531 8415
rect 17693 8381 17727 8415
rect 18705 8381 18739 8415
rect 18889 8381 18923 8415
rect 19165 8381 19199 8415
rect 19625 8381 19659 8415
rect 19809 8381 19843 8415
rect 20085 8381 20119 8415
rect 20269 8381 20303 8415
rect 20453 8381 20487 8415
rect 20729 8381 20763 8415
rect 20821 8381 20855 8415
rect 21465 8381 21499 8415
rect 21557 8381 21591 8415
rect 21741 8381 21775 8415
rect 23397 8381 23431 8415
rect 24970 8381 25004 8415
rect 25237 8381 25271 8415
rect 25605 8381 25639 8415
rect 3700 8313 3734 8347
rect 5172 8313 5206 8347
rect 9229 8313 9263 8347
rect 10425 8313 10459 8347
rect 10517 8313 10551 8347
rect 11881 8313 11915 8347
rect 12081 8313 12115 8347
rect 14013 8313 14047 8347
rect 14229 8313 14263 8347
rect 14933 8313 14967 8347
rect 15117 8313 15151 8347
rect 18337 8313 18371 8347
rect 19349 8313 19383 8347
rect 20545 8313 20579 8347
rect 23581 8313 23615 8347
rect 25850 8313 25884 8347
rect 2513 8245 2547 8279
rect 7297 8245 7331 8279
rect 14381 8245 14415 8279
rect 16313 8245 16347 8279
rect 21373 8245 21407 8279
rect 21649 8245 21683 8279
rect 23857 8245 23891 8279
rect 26985 8245 27019 8279
rect 10609 8041 10643 8075
rect 18613 8041 18647 8075
rect 21005 8041 21039 8075
rect 22661 8041 22695 8075
rect 23305 8041 23339 8075
rect 24041 8041 24075 8075
rect 24777 8041 24811 8075
rect 24869 8041 24903 8075
rect 25605 8041 25639 8075
rect 26433 8041 26467 8075
rect 4169 7973 4203 8007
rect 6653 7973 6687 8007
rect 7174 7973 7208 8007
rect 9474 7973 9508 8007
rect 10977 7973 11011 8007
rect 12817 7973 12851 8007
rect 15209 7973 15243 8007
rect 18521 7973 18555 8007
rect 23121 7973 23155 8007
rect 24409 7973 24443 8007
rect 24593 7973 24627 8007
rect 2513 7905 2547 7939
rect 2697 7905 2731 7939
rect 3433 7905 3467 7939
rect 4445 7905 4479 7939
rect 6009 7905 6043 7939
rect 6929 7905 6963 7939
rect 8401 7905 8435 7939
rect 9229 7905 9263 7939
rect 11161 7905 11195 7939
rect 12173 7905 12207 7939
rect 12633 7905 12667 7939
rect 12909 7905 12943 7939
rect 13277 7905 13311 7939
rect 13645 7905 13679 7939
rect 13912 7905 13946 7939
rect 15117 7905 15151 7939
rect 15301 7905 15335 7939
rect 15577 7905 15611 7939
rect 15853 7905 15887 7939
rect 16129 7905 16163 7939
rect 16396 7905 16430 7939
rect 19073 7905 19107 7939
rect 19533 7905 19567 7939
rect 19625 7905 19659 7939
rect 19809 7905 19843 7939
rect 19901 7905 19935 7939
rect 20361 7905 20395 7939
rect 20637 7905 20671 7939
rect 20821 7905 20855 7939
rect 20913 7905 20947 7939
rect 21097 7905 21131 7939
rect 21548 7905 21582 7939
rect 22753 7905 22787 7939
rect 22937 7905 22971 7939
rect 23489 7905 23523 7939
rect 23673 7905 23707 7939
rect 23765 7905 23799 7939
rect 23949 7905 23983 7939
rect 24041 7905 24075 7939
rect 24225 7905 24259 7939
rect 25421 7905 25455 7939
rect 25881 7905 25915 7939
rect 25973 7905 26007 7939
rect 26065 7905 26099 7939
rect 26249 7905 26283 7939
rect 27077 7905 27111 7939
rect 8677 7837 8711 7871
rect 9137 7837 9171 7871
rect 12357 7837 12391 7871
rect 13093 7837 13127 7871
rect 13185 7837 13219 7871
rect 13369 7837 13403 7871
rect 17693 7837 17727 7871
rect 18797 7837 18831 7871
rect 18889 7837 18923 7871
rect 18981 7837 19015 7871
rect 20177 7837 20211 7871
rect 21281 7837 21315 7871
rect 4261 7769 4295 7803
rect 5825 7769 5859 7803
rect 6285 7769 6319 7803
rect 6837 7769 6871 7803
rect 8861 7769 8895 7803
rect 12449 7769 12483 7803
rect 15025 7769 15059 7803
rect 23857 7769 23891 7803
rect 2513 7701 2547 7735
rect 6653 7701 6687 7735
rect 8309 7701 8343 7735
rect 8585 7701 8619 7735
rect 11345 7701 11379 7735
rect 11989 7701 12023 7735
rect 13553 7701 13587 7735
rect 17509 7701 17543 7735
rect 19349 7701 19383 7735
rect 2605 7497 2639 7531
rect 3249 7497 3283 7531
rect 4261 7497 4295 7531
rect 4445 7497 4479 7531
rect 5917 7497 5951 7531
rect 6101 7497 6135 7531
rect 7297 7497 7331 7531
rect 9321 7497 9355 7531
rect 9965 7497 9999 7531
rect 14105 7497 14139 7531
rect 14841 7497 14875 7531
rect 15669 7497 15703 7531
rect 16221 7497 16255 7531
rect 16405 7497 16439 7531
rect 18337 7497 18371 7531
rect 18889 7497 18923 7531
rect 19533 7497 19567 7531
rect 21649 7497 21683 7531
rect 21741 7497 21775 7531
rect 26341 7497 26375 7531
rect 4537 7429 4571 7463
rect 13645 7429 13679 7463
rect 15853 7429 15887 7463
rect 16681 7429 16715 7463
rect 17693 7429 17727 7463
rect 18705 7429 18739 7463
rect 19441 7429 19475 7463
rect 2973 7361 3007 7395
rect 3433 7361 3467 7395
rect 5549 7361 5583 7395
rect 6193 7361 6227 7395
rect 7481 7361 7515 7395
rect 8125 7361 8159 7395
rect 9597 7361 9631 7395
rect 12357 7361 12391 7395
rect 12633 7361 12667 7395
rect 14013 7361 14047 7395
rect 21925 7361 21959 7395
rect 22201 7361 22235 7395
rect 26893 7361 26927 7395
rect 857 7293 891 7327
rect 2513 7293 2547 7327
rect 3525 7293 3559 7327
rect 3617 7293 3651 7327
rect 3709 7293 3743 7327
rect 4721 7293 4755 7327
rect 4813 7293 4847 7327
rect 4997 7293 5031 7327
rect 5089 7293 5123 7327
rect 5457 7293 5491 7327
rect 6469 7293 6503 7327
rect 6561 7293 6595 7327
rect 6653 7293 6687 7327
rect 6837 7293 6871 7327
rect 7205 7293 7239 7327
rect 7573 7293 7607 7327
rect 8033 7293 8067 7327
rect 8217 7293 8251 7327
rect 8401 7293 8435 7327
rect 9505 7293 9539 7327
rect 9689 7293 9723 7327
rect 9781 7293 9815 7327
rect 10149 7293 10183 7327
rect 10425 7293 10459 7327
rect 10517 7293 10551 7327
rect 10701 7293 10735 7327
rect 11805 7293 11839 7327
rect 12081 7293 12115 7327
rect 12265 7293 12299 7327
rect 12541 7293 12575 7327
rect 12725 7293 12759 7327
rect 12817 7293 12851 7327
rect 14289 7293 14323 7327
rect 15025 7293 15059 7327
rect 15117 7293 15151 7327
rect 15301 7293 15335 7327
rect 15393 7293 15427 7327
rect 15761 7293 15795 7327
rect 16957 7293 16991 7327
rect 17049 7293 17083 7327
rect 17141 7293 17175 7327
rect 17325 7293 17359 7327
rect 17877 7293 17911 7327
rect 18153 7293 18187 7327
rect 18245 7293 18279 7327
rect 18429 7293 18463 7327
rect 19717 7293 19751 7327
rect 19993 7293 20027 7327
rect 20177 7293 20211 7327
rect 21373 7293 21407 7327
rect 21465 7293 21499 7327
rect 22017 7293 22051 7327
rect 22109 7293 22143 7327
rect 23213 7293 23247 7327
rect 23305 7293 23339 7327
rect 23489 7293 23523 7327
rect 23581 7293 23615 7327
rect 24409 7293 24443 7327
rect 24685 7293 24719 7327
rect 1124 7225 1158 7259
rect 4077 7225 4111 7259
rect 5365 7225 5399 7259
rect 7113 7225 7147 7259
rect 8585 7225 8619 7259
rect 10609 7225 10643 7259
rect 19073 7225 19107 7259
rect 21649 7225 21683 7259
rect 24930 7225 24964 7259
rect 2237 7157 2271 7191
rect 4277 7157 4311 7191
rect 5917 7157 5951 7191
rect 7941 7157 7975 7191
rect 8769 7157 8803 7191
rect 10333 7157 10367 7191
rect 11621 7157 11655 7191
rect 13553 7157 13587 7191
rect 16221 7157 16255 7191
rect 18061 7157 18095 7191
rect 18873 7157 18907 7191
rect 23029 7157 23063 7191
rect 24593 7157 24627 7191
rect 26065 7157 26099 7191
rect 2145 6953 2179 6987
rect 6009 6953 6043 6987
rect 7481 6953 7515 6987
rect 7665 6953 7699 6987
rect 12817 6953 12851 6987
rect 13645 6953 13679 6987
rect 16497 6953 16531 6987
rect 19625 6953 19659 6987
rect 20177 6953 20211 6987
rect 2421 6885 2455 6919
rect 3341 6885 3375 6919
rect 4537 6885 4571 6919
rect 11244 6885 11278 6919
rect 17233 6885 17267 6919
rect 21373 6885 21407 6919
rect 21589 6885 21623 6919
rect 26617 6885 26651 6919
rect 2053 6817 2087 6851
rect 2237 6817 2271 6851
rect 2329 6817 2363 6851
rect 2513 6817 2547 6851
rect 2861 6817 2895 6851
rect 2973 6817 3007 6851
rect 3065 6817 3099 6851
rect 3249 6817 3283 6851
rect 3525 6817 3559 6851
rect 3617 6817 3651 6851
rect 4261 6817 4295 6851
rect 4905 6817 4939 6851
rect 4997 6817 5031 6851
rect 5089 6817 5123 6851
rect 5273 6817 5307 6851
rect 6193 6817 6227 6851
rect 6285 6817 6319 6851
rect 6469 6817 6503 6851
rect 6561 6817 6595 6851
rect 6653 6817 6687 6851
rect 6837 6817 6871 6851
rect 10977 6817 11011 6851
rect 12449 6817 12483 6851
rect 12633 6817 12667 6851
rect 13093 6817 13127 6851
rect 13553 6817 13587 6851
rect 13737 6817 13771 6851
rect 16681 6817 16715 6851
rect 16773 6817 16807 6851
rect 16957 6817 16991 6851
rect 17049 6817 17083 6851
rect 17325 6817 17359 6851
rect 17601 6817 17635 6851
rect 17785 6817 17819 6851
rect 17877 6817 17911 6851
rect 18409 6817 18443 6851
rect 19809 6817 19843 6851
rect 19993 6817 20027 6851
rect 20085 6817 20119 6851
rect 20269 6817 20303 6851
rect 23121 6817 23155 6851
rect 23305 6817 23339 6851
rect 23581 6817 23615 6851
rect 23765 6817 23799 6851
rect 24133 6817 24167 6851
rect 24225 6817 24259 6851
rect 24685 6817 24719 6851
rect 24777 6817 24811 6851
rect 24869 6817 24903 6851
rect 25053 6817 25087 6851
rect 25145 6817 25179 6851
rect 25237 6817 25271 6851
rect 25421 6817 25455 6851
rect 25513 6817 25547 6851
rect 25789 6817 25823 6851
rect 25973 6817 26007 6851
rect 26157 6817 26191 6851
rect 26433 6817 26467 6851
rect 26801 6817 26835 6851
rect 2605 6749 2639 6783
rect 4445 6749 4479 6783
rect 4629 6749 4663 6783
rect 4721 6749 4755 6783
rect 5457 6749 5491 6783
rect 7021 6749 7055 6783
rect 17417 6749 17451 6783
rect 18153 6749 18187 6783
rect 24409 6749 24443 6783
rect 3341 6681 3375 6715
rect 8033 6681 8067 6715
rect 19533 6681 19567 6715
rect 23029 6681 23063 6715
rect 4077 6613 4111 6647
rect 7665 6613 7699 6647
rect 12357 6613 12391 6647
rect 13277 6613 13311 6647
rect 18061 6613 18095 6647
rect 21557 6613 21591 6647
rect 21741 6613 21775 6647
rect 25697 6613 25731 6647
rect 2973 6409 3007 6443
rect 3893 6409 3927 6443
rect 4721 6409 4755 6443
rect 6009 6409 6043 6443
rect 7481 6409 7515 6443
rect 7757 6409 7791 6443
rect 9137 6409 9171 6443
rect 9413 6409 9447 6443
rect 11529 6409 11563 6443
rect 12541 6409 12575 6443
rect 16221 6409 16255 6443
rect 23581 6409 23615 6443
rect 24409 6409 24443 6443
rect 24593 6409 24627 6443
rect 25329 6409 25363 6443
rect 25789 6409 25823 6443
rect 3617 6341 3651 6375
rect 9321 6341 9355 6375
rect 11989 6341 12023 6375
rect 14933 6273 14967 6307
rect 21741 6273 21775 6307
rect 24041 6273 24075 6307
rect 2881 6205 2915 6239
rect 3065 6205 3099 6239
rect 3249 6205 3283 6239
rect 3433 6205 3467 6239
rect 4353 6205 4387 6239
rect 4629 6205 4663 6239
rect 4813 6205 4847 6239
rect 4905 6205 4939 6239
rect 5917 6205 5951 6239
rect 6101 6205 6135 6239
rect 6377 6205 6411 6239
rect 7113 6205 7147 6239
rect 9597 6205 9631 6239
rect 9689 6205 9723 6239
rect 9873 6205 9907 6239
rect 9965 6205 9999 6239
rect 10057 6205 10091 6239
rect 10333 6205 10367 6239
rect 10609 6205 10643 6239
rect 10885 6205 10919 6239
rect 11713 6205 11747 6239
rect 11805 6205 11839 6239
rect 12265 6205 12299 6239
rect 12357 6205 12391 6239
rect 12541 6205 12575 6239
rect 13185 6205 13219 6239
rect 13369 6205 13403 6239
rect 14666 6205 14700 6239
rect 15577 6205 15611 6239
rect 15761 6205 15795 6239
rect 16589 6205 16623 6239
rect 17233 6205 17267 6239
rect 17417 6205 17451 6239
rect 21465 6205 21499 6239
rect 23397 6205 23431 6239
rect 25237 6205 25271 6239
rect 25421 6205 25455 6239
rect 26157 6205 26191 6239
rect 3861 6137 3895 6171
rect 4077 6137 4111 6171
rect 7297 6137 7331 6171
rect 7573 6137 7607 6171
rect 8953 6137 8987 6171
rect 9169 6137 9203 6171
rect 10149 6137 10183 6171
rect 11989 6137 12023 6171
rect 15301 6137 15335 6171
rect 15485 6137 15519 6171
rect 21986 6137 22020 6171
rect 23213 6137 23247 6171
rect 24409 6137 24443 6171
rect 25973 6137 26007 6171
rect 3709 6069 3743 6103
rect 7773 6069 7807 6103
rect 7941 6069 7975 6103
rect 12173 6069 12207 6103
rect 13185 6069 13219 6103
rect 13553 6069 13587 6103
rect 15117 6069 15151 6103
rect 15577 6069 15611 6103
rect 16037 6069 16071 6103
rect 16221 6069 16255 6103
rect 17233 6069 17267 6103
rect 21649 6069 21683 6103
rect 23121 6069 23155 6103
rect 3525 5865 3559 5899
rect 5641 5865 5675 5899
rect 9965 5865 9999 5899
rect 10057 5865 10091 5899
rect 10517 5865 10551 5899
rect 14197 5865 14231 5899
rect 14381 5865 14415 5899
rect 16497 5865 16531 5899
rect 17141 5865 17175 5899
rect 21281 5865 21315 5899
rect 21449 5865 21483 5899
rect 23029 5865 23063 5899
rect 25053 5865 25087 5899
rect 10425 5797 10459 5831
rect 13829 5797 13863 5831
rect 14013 5797 14047 5831
rect 17417 5797 17451 5831
rect 17877 5797 17911 5831
rect 21649 5797 21683 5831
rect 21925 5797 21959 5831
rect 24685 5797 24719 5831
rect 2605 5729 2639 5763
rect 3065 5729 3099 5763
rect 3249 5729 3283 5763
rect 4261 5729 4295 5763
rect 4537 5729 4571 5763
rect 4629 5729 4663 5763
rect 4905 5729 4939 5763
rect 6009 5729 6043 5763
rect 6285 5729 6319 5763
rect 8226 5729 8260 5763
rect 8493 5729 8527 5763
rect 8585 5729 8619 5763
rect 8852 5729 8886 5763
rect 10241 5729 10275 5763
rect 10517 5729 10551 5763
rect 10701 5729 10735 5763
rect 15494 5729 15528 5763
rect 16221 5729 16255 5763
rect 16681 5729 16715 5763
rect 18061 5729 18095 5763
rect 19993 5729 20027 5763
rect 21097 5729 21131 5763
rect 21741 5729 21775 5763
rect 22937 5729 22971 5763
rect 23121 5729 23155 5763
rect 25145 5729 25179 5763
rect 25237 5729 25271 5763
rect 25513 5729 25547 5763
rect 25697 5729 25731 5763
rect 15761 5661 15795 5695
rect 16773 5661 16807 5695
rect 17785 5661 17819 5695
rect 19717 5661 19751 5695
rect 25605 5661 25639 5695
rect 7021 5593 7055 5627
rect 18337 5593 18371 5627
rect 20729 5593 20763 5627
rect 24317 5593 24351 5627
rect 1225 5525 1259 5559
rect 2421 5525 2455 5559
rect 3157 5525 3191 5559
rect 7113 5525 7147 5559
rect 12449 5525 12483 5559
rect 16405 5525 16439 5559
rect 17233 5525 17267 5559
rect 17417 5525 17451 5559
rect 18245 5525 18279 5559
rect 18981 5525 19015 5559
rect 19349 5525 19383 5559
rect 20913 5525 20947 5559
rect 21465 5525 21499 5559
rect 22109 5525 22143 5559
rect 22569 5525 22603 5559
rect 24685 5525 24719 5559
rect 24869 5525 24903 5559
rect 25421 5525 25455 5559
rect 3065 5321 3099 5355
rect 5457 5321 5491 5355
rect 6285 5321 6319 5355
rect 7573 5321 7607 5355
rect 8033 5321 8067 5355
rect 9045 5321 9079 5355
rect 11621 5321 11655 5355
rect 14565 5321 14599 5355
rect 15301 5321 15335 5355
rect 15577 5321 15611 5355
rect 21649 5321 21683 5355
rect 21833 5321 21867 5355
rect 5181 5253 5215 5287
rect 17601 5253 17635 5287
rect 19993 5253 20027 5287
rect 23581 5253 23615 5287
rect 1685 5185 1719 5219
rect 6101 5185 6135 5219
rect 6469 5185 6503 5219
rect 6653 5185 6687 5219
rect 6745 5185 6779 5219
rect 7021 5185 7055 5219
rect 16221 5185 16255 5219
rect 18889 5185 18923 5219
rect 20269 5185 20303 5219
rect 22569 5185 22603 5219
rect 24225 5185 24259 5219
rect 24685 5185 24719 5219
rect 25053 5185 25087 5219
rect 1593 5117 1627 5151
rect 1952 5117 1986 5151
rect 3249 5117 3283 5151
rect 4077 5117 4111 5151
rect 4169 5117 4203 5151
rect 4445 5117 4479 5151
rect 5273 5117 5307 5151
rect 5457 5117 5491 5151
rect 6009 5119 6043 5153
rect 6193 5117 6227 5151
rect 6561 5117 6595 5151
rect 6929 5117 6963 5151
rect 7113 5117 7147 5151
rect 7481 5117 7515 5151
rect 7665 5117 7699 5151
rect 7849 5117 7883 5151
rect 9229 5117 9263 5151
rect 10517 5117 10551 5151
rect 10609 5117 10643 5151
rect 10885 5117 10919 5151
rect 11897 5117 11931 5151
rect 12357 5117 12391 5151
rect 12633 5117 12667 5151
rect 13553 5117 13587 5151
rect 13829 5117 13863 5151
rect 15761 5117 15795 5151
rect 16477 5117 16511 5151
rect 17969 5117 18003 5151
rect 18153 5117 18187 5151
rect 19165 5117 19199 5151
rect 20536 5117 20570 5151
rect 21741 5117 21775 5151
rect 21925 5117 21959 5151
rect 22201 5117 22235 5151
rect 22845 5117 22879 5151
rect 24593 5117 24627 5151
rect 25320 5117 25354 5151
rect 3433 5049 3467 5083
rect 12081 5049 12115 5083
rect 15117 5049 15151 5083
rect 15333 5049 15367 5083
rect 1409 4981 1443 5015
rect 3617 4981 3651 5015
rect 12265 4981 12299 5015
rect 13369 4981 13403 5015
rect 15485 4981 15519 5015
rect 18061 4981 18095 5015
rect 19901 4981 19935 5015
rect 24869 4981 24903 5015
rect 26433 4981 26467 5015
rect 2145 4777 2179 4811
rect 2973 4777 3007 4811
rect 4905 4777 4939 4811
rect 4997 4777 5031 4811
rect 5825 4777 5859 4811
rect 8401 4777 8435 4811
rect 10793 4777 10827 4811
rect 12173 4777 12207 4811
rect 13369 4777 13403 4811
rect 15209 4777 15243 4811
rect 18797 4777 18831 4811
rect 19165 4777 19199 4811
rect 20269 4777 20303 4811
rect 22017 4777 22051 4811
rect 23121 4777 23155 4811
rect 23213 4777 23247 4811
rect 24409 4777 24443 4811
rect 25145 4777 25179 4811
rect 6009 4709 6043 4743
rect 6469 4709 6503 4743
rect 6653 4709 6687 4743
rect 12357 4709 12391 4743
rect 12725 4709 12759 4743
rect 25329 4709 25363 4743
rect 25513 4709 25547 4743
rect 1133 4641 1167 4675
rect 1409 4641 1443 4675
rect 2973 4641 3007 4675
rect 3157 4641 3191 4675
rect 4721 4641 4755 4675
rect 5181 4641 5215 4675
rect 6377 4641 6411 4675
rect 6837 4641 6871 4675
rect 7113 4641 7147 4675
rect 7389 4641 7423 4675
rect 7665 4641 7699 4675
rect 8493 4641 8527 4675
rect 10609 4641 10643 4675
rect 11069 4641 11103 4675
rect 11253 4641 11287 4675
rect 11345 4641 11379 4675
rect 11529 4641 11563 4675
rect 12541 4641 12575 4675
rect 13185 4641 13219 4675
rect 13461 4641 13495 4675
rect 14473 4641 14507 4675
rect 17785 4641 17819 4675
rect 18061 4641 18095 4675
rect 18981 4641 19015 4675
rect 19257 4641 19291 4675
rect 19533 4641 19567 4675
rect 21833 4641 21867 4675
rect 22385 4641 22419 4675
rect 23397 4641 23431 4675
rect 24041 4641 24075 4675
rect 11437 4573 11471 4607
rect 11713 4573 11747 4607
rect 11805 4573 11839 4607
rect 11897 4573 11931 4607
rect 11989 4573 12023 4607
rect 14105 4573 14139 4607
rect 14197 4573 14231 4607
rect 22109 4573 22143 4607
rect 6929 4505 6963 4539
rect 11161 4505 11195 4539
rect 12909 4505 12943 4539
rect 24593 4505 24627 4539
rect 2697 4437 2731 4471
rect 6009 4437 6043 4471
rect 9413 4437 9447 4471
rect 9689 4437 9723 4471
rect 16405 4437 16439 4471
rect 24409 4437 24443 4471
rect 4261 4233 4295 4267
rect 7573 4233 7607 4267
rect 11069 4233 11103 4267
rect 11253 4233 11287 4267
rect 13645 4233 13679 4267
rect 14013 4233 14047 4267
rect 14289 4233 14323 4267
rect 15853 4233 15887 4267
rect 18337 4233 18371 4267
rect 18521 4233 18555 4267
rect 22385 4233 22419 4267
rect 22569 4233 22603 4267
rect 25329 4233 25363 4267
rect 11621 4165 11655 4199
rect 15209 4165 15243 4199
rect 18797 4165 18831 4199
rect 3249 4097 3283 4131
rect 8953 4097 8987 4131
rect 9413 4097 9447 4131
rect 15301 4097 15335 4131
rect 16313 4097 16347 4131
rect 19165 4097 19199 4131
rect 19340 4097 19374 4131
rect 19434 4097 19468 4131
rect 19717 4097 19751 4131
rect 20729 4097 20763 4131
rect 21649 4097 21683 4131
rect 22293 4097 22327 4131
rect 1501 4029 1535 4063
rect 1593 4029 1627 4063
rect 1869 4029 1903 4063
rect 2881 4029 2915 4063
rect 3525 4029 3559 4063
rect 4353 4029 4387 4063
rect 4537 4029 4571 4063
rect 6101 4029 6135 4063
rect 6285 4029 6319 4063
rect 7297 4029 7331 4063
rect 7757 4029 7791 4063
rect 7849 4029 7883 4063
rect 8033 4029 8067 4063
rect 8125 4029 8159 4063
rect 8769 4029 8803 4063
rect 8861 4029 8895 4063
rect 9045 4029 9079 4063
rect 9689 4029 9723 4063
rect 10517 4029 10551 4063
rect 10701 4029 10735 4063
rect 12633 4029 12667 4063
rect 12817 4029 12851 4063
rect 13185 4029 13219 4063
rect 13277 4029 13311 4063
rect 13829 4029 13863 4063
rect 14013 4029 14047 4063
rect 14105 4029 14139 4063
rect 15025 4029 15059 4063
rect 15209 4029 15243 4063
rect 15485 4029 15519 4063
rect 15669 4029 15703 4063
rect 15853 4029 15887 4063
rect 15945 4029 15979 4063
rect 16589 4029 16623 4063
rect 17601 4029 17635 4063
rect 17969 4029 18003 4063
rect 18705 4029 18739 4063
rect 18889 4029 18923 4063
rect 19257 4029 19291 4063
rect 19625 4029 19659 4063
rect 19809 4029 19843 4063
rect 20637 4029 20671 4063
rect 20821 4029 20855 4063
rect 21557 4029 21591 4063
rect 22201 4029 22235 4063
rect 23029 4029 23063 4063
rect 23213 4029 23247 4063
rect 23489 4029 23523 4063
rect 24225 4029 24259 4063
rect 24317 4029 24351 4063
rect 24593 4029 24627 4063
rect 4445 3961 4479 3995
rect 7113 3961 7147 3995
rect 7481 3961 7515 3995
rect 8585 3961 8619 3995
rect 10609 3961 10643 3995
rect 17417 3961 17451 3995
rect 2605 3893 2639 3927
rect 3065 3893 3099 3927
rect 6193 3893 6227 3927
rect 8401 3893 8435 3927
rect 10425 3893 10459 3927
rect 11253 3893 11287 3927
rect 12725 3893 12759 3927
rect 16221 3893 16255 3927
rect 17325 3893 17359 3927
rect 17785 3893 17819 3927
rect 18337 3893 18371 3927
rect 18981 3893 19015 3927
rect 23121 3893 23155 3927
rect 23673 3893 23707 3927
rect 4997 3689 5031 3723
rect 6469 3689 6503 3723
rect 7573 3689 7607 3723
rect 10149 3689 10183 3723
rect 12357 3689 12391 3723
rect 13921 3689 13955 3723
rect 15501 3689 15535 3723
rect 15945 3689 15979 3723
rect 16497 3689 16531 3723
rect 18889 3689 18923 3723
rect 19993 3689 20027 3723
rect 21833 3689 21867 3723
rect 25513 3689 25547 3723
rect 3709 3621 3743 3655
rect 3985 3621 4019 3655
rect 15301 3621 15335 3655
rect 17877 3621 17911 3655
rect 18245 3621 18279 3655
rect 20821 3621 20855 3655
rect 21373 3621 21407 3655
rect 23765 3621 23799 3655
rect 23995 3587 24029 3621
rect 3617 3553 3651 3587
rect 3893 3553 3927 3587
rect 4169 3553 4203 3587
rect 4353 3553 4387 3587
rect 4629 3553 4663 3587
rect 6101 3553 6135 3587
rect 6285 3553 6319 3587
rect 6837 3553 6871 3587
rect 6929 3553 6963 3587
rect 7481 3553 7515 3587
rect 7665 3553 7699 3587
rect 8217 3553 8251 3587
rect 8401 3553 8435 3587
rect 9137 3553 9171 3587
rect 9413 3553 9447 3587
rect 10977 3553 11011 3587
rect 11161 3553 11195 3587
rect 12449 3553 12483 3587
rect 12633 3553 12667 3587
rect 13461 3553 13495 3587
rect 13737 3553 13771 3587
rect 15761 3553 15795 3587
rect 16313 3553 16347 3587
rect 18797 3553 18831 3587
rect 18981 3553 19015 3587
rect 19533 3553 19567 3587
rect 20177 3553 20211 3587
rect 20545 3553 20579 3587
rect 20729 3553 20763 3587
rect 20913 3553 20947 3587
rect 21649 3553 21683 3587
rect 23489 3553 23523 3587
rect 24777 3553 24811 3587
rect 4721 3485 4755 3519
rect 6193 3485 6227 3519
rect 6745 3485 6779 3519
rect 7021 3485 7055 3519
rect 11897 3485 11931 3519
rect 13645 3485 13679 3519
rect 18061 3485 18095 3519
rect 21557 3485 21591 3519
rect 23305 3485 23339 3519
rect 24409 3485 24443 3519
rect 24501 3485 24535 3519
rect 12173 3417 12207 3451
rect 15669 3417 15703 3451
rect 18429 3417 18463 3451
rect 19809 3417 19843 3451
rect 4813 3349 4847 3383
rect 6837 3349 6871 3383
rect 8309 3349 8343 3383
rect 11069 3349 11103 3383
rect 12817 3349 12851 3383
rect 13461 3349 13495 3383
rect 15485 3349 15519 3383
rect 16589 3349 16623 3383
rect 20545 3349 20579 3383
rect 21373 3349 21407 3383
rect 23673 3349 23707 3383
rect 23949 3349 23983 3383
rect 24133 3349 24167 3383
rect 4261 3145 4295 3179
rect 4445 3145 4479 3179
rect 5181 3145 5215 3179
rect 6745 3145 6779 3179
rect 10425 3145 10459 3179
rect 12817 3145 12851 3179
rect 13737 3145 13771 3179
rect 14289 3145 14323 3179
rect 15117 3145 15151 3179
rect 15301 3145 15335 3179
rect 15761 3145 15795 3179
rect 17785 3145 17819 3179
rect 22293 3145 22327 3179
rect 23029 3145 23063 3179
rect 23857 3145 23891 3179
rect 24225 3145 24259 3179
rect 24317 3145 24351 3179
rect 24777 3145 24811 3179
rect 5549 3077 5583 3111
rect 9597 3077 9631 3111
rect 17417 3077 17451 3111
rect 19993 3077 20027 3111
rect 20637 3077 20671 3111
rect 20729 3077 20763 3111
rect 23213 3077 23247 3111
rect 4537 3009 4571 3043
rect 6285 3009 6319 3043
rect 12725 3009 12759 3043
rect 15393 3009 15427 3043
rect 16405 3009 16439 3043
rect 17969 3009 18003 3043
rect 19625 3009 19659 3043
rect 20821 3009 20855 3043
rect 22017 3009 22051 3043
rect 22477 3009 22511 3043
rect 24409 3009 24443 3043
rect 3341 2941 3375 2975
rect 3525 2941 3559 2975
rect 4077 2941 4111 2975
rect 4169 2941 4203 2975
rect 4721 2941 4755 2975
rect 4813 2941 4847 2975
rect 4997 2941 5031 2975
rect 5089 2941 5123 2975
rect 5181 2941 5215 2975
rect 5365 2941 5399 2975
rect 5641 2941 5675 2975
rect 5917 2941 5951 2975
rect 6499 2941 6533 2975
rect 6653 2941 6687 2975
rect 6745 2941 6779 2975
rect 6929 2941 6963 2975
rect 7849 2941 7883 2975
rect 8033 2941 8067 2975
rect 8401 2941 8435 2975
rect 10517 2941 10551 2975
rect 10609 2941 10643 2975
rect 10763 2941 10797 2975
rect 11529 2941 11563 2975
rect 11989 2941 12023 2975
rect 12449 2941 12483 2975
rect 12541 2941 12575 2975
rect 12817 2941 12851 2975
rect 13001 2941 13035 2975
rect 13185 2941 13219 2975
rect 13369 2941 13403 2975
rect 13553 2941 13587 2975
rect 13737 2941 13771 2975
rect 14059 2941 14093 2975
rect 14197 2941 14231 2975
rect 14289 2941 14323 2975
rect 14473 2941 14507 2975
rect 14749 2941 14783 2975
rect 16129 2941 16163 2975
rect 16681 2941 16715 2975
rect 17509 2941 17543 2975
rect 18245 2941 18279 2975
rect 18705 2941 18739 2975
rect 18798 2941 18832 2975
rect 19809 2941 19843 2975
rect 20545 2941 20579 2975
rect 21649 2941 21683 2975
rect 21742 2941 21776 2975
rect 22109 2941 22143 2975
rect 22293 2941 22327 2975
rect 22385 2941 22419 2975
rect 22569 2941 22603 2975
rect 22661 2941 22695 2975
rect 23489 2941 23523 2975
rect 23857 2941 23891 2975
rect 24041 2941 24075 2975
rect 24317 2941 24351 2975
rect 24961 2941 24995 2975
rect 25053 2941 25087 2975
rect 3433 2873 3467 2907
rect 9781 2873 9815 2907
rect 9965 2873 9999 2907
rect 11805 2873 11839 2907
rect 13829 2873 13863 2907
rect 15117 2873 15151 2907
rect 15761 2873 15795 2907
rect 18429 2873 18463 2907
rect 19073 2873 19107 2907
rect 23029 2873 23063 2907
rect 7941 2805 7975 2839
rect 10057 2805 10091 2839
rect 10977 2805 11011 2839
rect 12725 2805 12759 2839
rect 13277 2805 13311 2839
rect 15945 2805 15979 2839
rect 16313 2805 16347 2839
rect 18061 2805 18095 2839
rect 23673 2805 23707 2839
rect 24685 2805 24719 2839
rect 25237 2805 25271 2839
rect 4905 2601 4939 2635
rect 7941 2601 7975 2635
rect 15945 2601 15979 2635
rect 23029 2601 23063 2635
rect 23213 2601 23247 2635
rect 23765 2601 23799 2635
rect 3617 2533 3651 2567
rect 14013 2533 14047 2567
rect 2605 2465 2639 2499
rect 3433 2465 3467 2499
rect 3525 2465 3559 2499
rect 3709 2465 3743 2499
rect 4537 2465 4571 2499
rect 4721 2465 4755 2499
rect 4997 2465 5031 2499
rect 5457 2465 5491 2499
rect 5641 2465 5675 2499
rect 5825 2465 5859 2499
rect 6653 2465 6687 2499
rect 7297 2465 7331 2499
rect 7481 2465 7515 2499
rect 7573 2465 7607 2499
rect 7757 2465 7791 2499
rect 7849 2465 7883 2499
rect 8033 2465 8067 2499
rect 8125 2465 8159 2499
rect 8401 2465 8435 2499
rect 9229 2465 9263 2499
rect 9689 2465 9723 2499
rect 9873 2465 9907 2499
rect 9965 2465 9999 2499
rect 10149 2465 10183 2499
rect 10241 2465 10275 2499
rect 10425 2465 10459 2499
rect 10977 2465 11011 2499
rect 11161 2465 11195 2499
rect 11345 2465 11379 2499
rect 11529 2465 11563 2499
rect 11621 2465 11655 2499
rect 11805 2465 11839 2499
rect 13921 2465 13955 2499
rect 14105 2465 14139 2499
rect 15577 2465 15611 2499
rect 16129 2465 16163 2499
rect 16405 2465 16439 2499
rect 17693 2465 17727 2499
rect 17877 2465 17911 2499
rect 17969 2465 18003 2499
rect 18153 2465 18187 2499
rect 18613 2465 18647 2499
rect 18797 2465 18831 2499
rect 18889 2465 18923 2499
rect 19073 2465 19107 2499
rect 19809 2465 19843 2499
rect 19993 2465 20027 2499
rect 20085 2465 20119 2499
rect 20269 2465 20303 2499
rect 20637 2465 20671 2499
rect 20821 2465 20855 2499
rect 21925 2465 21959 2499
rect 22109 2465 22143 2499
rect 22201 2465 22235 2499
rect 22385 2465 22419 2499
rect 23581 2465 23615 2499
rect 2237 2397 2271 2431
rect 2329 2397 2363 2431
rect 6929 2397 6963 2431
rect 7389 2397 7423 2431
rect 15669 2397 15703 2431
rect 22661 2397 22695 2431
rect 22109 2329 22143 2363
rect 22385 2329 22419 2363
rect 4537 2261 4571 2295
rect 5641 2261 5675 2295
rect 7021 2261 7055 2295
rect 7757 2261 7791 2295
rect 9689 2261 9723 2295
rect 10149 2261 10183 2295
rect 10241 2261 10275 2295
rect 11161 2261 11195 2295
rect 11529 2261 11563 2295
rect 11805 2261 11839 2295
rect 12357 2261 12391 2295
rect 15301 2261 15335 2295
rect 15761 2261 15795 2295
rect 16313 2261 16347 2295
rect 16589 2261 16623 2295
rect 17693 2261 17727 2295
rect 18153 2261 18187 2295
rect 18797 2261 18831 2295
rect 19073 2261 19107 2295
rect 19993 2261 20027 2295
rect 20269 2261 20303 2295
rect 20821 2261 20855 2295
rect 23029 2261 23063 2295
rect 7481 1989 7515 2023
rect 22661 1989 22695 2023
rect 6285 1921 6319 1955
rect 15209 1921 15243 1955
rect 23949 1921 23983 1955
rect 25145 1921 25179 1955
rect 949 1853 983 1887
rect 1225 1853 1259 1887
rect 2053 1853 2087 1887
rect 2145 1853 2179 1887
rect 2789 1853 2823 1887
rect 2973 1853 3007 1887
rect 3249 1853 3283 1887
rect 3433 1853 3467 1887
rect 3525 1853 3559 1887
rect 3709 1853 3743 1887
rect 4261 1853 4295 1887
rect 4353 1853 4387 1887
rect 4537 1853 4571 1887
rect 4629 1853 4663 1887
rect 4813 1853 4847 1887
rect 5089 1853 5123 1887
rect 5365 1853 5399 1887
rect 6193 1853 6227 1887
rect 6561 1853 6595 1887
rect 7389 1853 7423 1887
rect 9045 1853 9079 1887
rect 9321 1853 9355 1887
rect 10149 1853 10183 1887
rect 10885 1853 10919 1887
rect 11069 1853 11103 1887
rect 11529 1853 11563 1887
rect 11621 1853 11655 1887
rect 11897 1853 11931 1887
rect 12725 1853 12759 1887
rect 12817 1853 12851 1887
rect 13001 1853 13035 1887
rect 13093 1853 13127 1887
rect 13277 1853 13311 1887
rect 13553 1853 13587 1887
rect 14105 1853 14139 1887
rect 14565 1853 14599 1887
rect 15485 1853 15519 1887
rect 16313 1853 16347 1887
rect 16405 1853 16439 1887
rect 16865 1853 16899 1887
rect 17417 1853 17451 1887
rect 17877 1853 17911 1887
rect 18705 1853 18739 1887
rect 19165 1853 19199 1887
rect 19441 1853 19475 1887
rect 19533 1853 19567 1887
rect 19809 1853 19843 1887
rect 20637 1853 20671 1887
rect 20913 1853 20947 1887
rect 21097 1853 21131 1887
rect 21189 1853 21223 1887
rect 21465 1853 21499 1887
rect 22293 1853 22327 1887
rect 22385 1853 22419 1887
rect 23121 1853 23155 1887
rect 23673 1853 23707 1887
rect 24225 1853 24259 1887
rect 25053 1853 25087 1887
rect 25421 1853 25455 1887
rect 2881 1785 2915 1819
rect 21005 1785 21039 1819
rect 3341 1717 3375 1751
rect 3617 1717 3651 1751
rect 4445 1717 4479 1751
rect 4721 1717 4755 1751
rect 12909 1717 12943 1751
rect 13185 1717 13219 1751
rect 1225 1377 1259 1411
rect 2053 1377 2087 1411
rect 2145 1377 2179 1411
rect 2973 1377 3007 1411
rect 3617 1377 3651 1411
rect 4445 1377 4479 1411
rect 4813 1377 4847 1411
rect 5641 1377 5675 1411
rect 7021 1377 7055 1411
rect 7849 1377 7883 1411
rect 8217 1377 8251 1411
rect 9045 1377 9079 1411
rect 9965 1377 9999 1411
rect 10793 1377 10827 1411
rect 11253 1377 11287 1411
rect 12081 1377 12115 1411
rect 13001 1377 13035 1411
rect 13277 1377 13311 1411
rect 13645 1377 13679 1411
rect 14473 1377 14507 1411
rect 14565 1377 14599 1411
rect 14841 1377 14875 1411
rect 15669 1377 15703 1411
rect 16405 1377 16439 1411
rect 17233 1377 17267 1411
rect 17325 1377 17359 1411
rect 17601 1377 17635 1411
rect 18429 1377 18463 1411
rect 18797 1377 18831 1411
rect 19625 1377 19659 1411
rect 19993 1377 20027 1411
rect 20821 1377 20855 1411
rect 21557 1377 21591 1411
rect 22385 1377 22419 1411
rect 22477 1377 22511 1411
rect 22753 1377 22787 1411
rect 23581 1377 23615 1411
rect 23949 1377 23983 1411
rect 24777 1377 24811 1411
rect 24869 1377 24903 1411
rect 25145 1377 25179 1411
rect 25973 1377 26007 1411
rect 949 1309 983 1343
rect 3249 1309 3283 1343
rect 3341 1309 3375 1343
rect 4537 1309 4571 1343
rect 6101 1309 6135 1343
rect 6745 1309 6779 1343
rect 7941 1309 7975 1343
rect 9597 1309 9631 1343
rect 9689 1309 9723 1343
rect 10977 1309 11011 1343
rect 13369 1309 13403 1343
rect 15945 1309 15979 1343
rect 16129 1309 16163 1343
rect 18521 1309 18555 1343
rect 19717 1309 19751 1343
rect 21281 1309 21315 1343
rect 23673 1309 23707 1343
rect 6009 1241 6043 1275
rect 6653 1173 6687 1207
rect 9321 1173 9355 1207
rect 12255 1173 12289 1207
rect 20913 1173 20947 1207
rect 1041 969 1075 1003
rect 1409 969 1443 1003
rect 3433 969 3467 1003
rect 5457 969 5491 1003
rect 7941 969 7975 1003
rect 9045 969 9079 1003
rect 13645 969 13679 1003
rect 21281 969 21315 1003
rect 21557 969 21591 1003
rect 23673 969 23707 1003
rect 3709 901 3743 935
rect 4261 833 4295 867
rect 6745 833 6779 867
rect 9413 833 9447 867
rect 10977 833 11011 867
rect 12265 833 12299 867
rect 18705 833 18739 867
rect 19993 833 20027 867
rect 23857 833 23891 867
rect 1961 765 1995 799
rect 2237 765 2271 799
rect 3065 765 3099 799
rect 4537 765 4571 799
rect 5365 765 5399 799
rect 7021 765 7055 799
rect 7849 765 7883 799
rect 9689 765 9723 799
rect 10517 765 10551 799
rect 11253 765 11287 799
rect 12081 765 12115 799
rect 12541 765 12575 799
rect 13369 765 13403 799
rect 14013 765 14047 799
rect 14289 765 14323 799
rect 15117 765 15151 799
rect 16221 765 16255 799
rect 16497 765 16531 799
rect 17325 765 17359 799
rect 17417 765 17451 799
rect 17693 765 17727 799
rect 18521 765 18555 799
rect 18981 765 19015 799
rect 19809 765 19843 799
rect 20269 765 20303 799
rect 21097 765 21131 799
rect 22201 765 22235 799
rect 22477 765 22511 799
rect 23305 765 23339 799
rect 24133 765 24167 799
rect 24961 765 24995 799
rect 25053 765 25087 799
rect 25329 765 25363 799
rect 26157 765 26191 799
<< metal1 >>
rect 16666 31084 16672 31136
rect 16724 31124 16730 31136
rect 19426 31124 19432 31136
rect 16724 31096 19432 31124
rect 16724 31084 16730 31096
rect 19426 31084 19432 31096
rect 19484 31084 19490 31136
rect 552 31034 27576 31056
rect 552 30982 7114 31034
rect 7166 30982 7178 31034
rect 7230 30982 7242 31034
rect 7294 30982 7306 31034
rect 7358 30982 7370 31034
rect 7422 30982 13830 31034
rect 13882 30982 13894 31034
rect 13946 30982 13958 31034
rect 14010 30982 14022 31034
rect 14074 30982 14086 31034
rect 14138 30982 20546 31034
rect 20598 30982 20610 31034
rect 20662 30982 20674 31034
rect 20726 30982 20738 31034
rect 20790 30982 20802 31034
rect 20854 30982 27262 31034
rect 27314 30982 27326 31034
rect 27378 30982 27390 31034
rect 27442 30982 27454 31034
rect 27506 30982 27518 31034
rect 27570 30982 27576 31034
rect 552 30960 27576 30982
rect 8389 30923 8447 30929
rect 8389 30889 8401 30923
rect 8435 30889 8447 30923
rect 8389 30883 8447 30889
rect 11977 30923 12035 30929
rect 11977 30889 11989 30923
rect 12023 30920 12035 30923
rect 12023 30892 13952 30920
rect 12023 30889 12035 30892
rect 11977 30883 12035 30889
rect 8404 30852 8432 30883
rect 10134 30861 10140 30864
rect 5828 30824 8432 30852
rect 10121 30855 10140 30861
rect 5626 30744 5632 30796
rect 5684 30784 5690 30796
rect 5828 30793 5856 30824
rect 10121 30821 10133 30855
rect 10121 30815 10140 30821
rect 10134 30812 10140 30815
rect 10192 30812 10198 30864
rect 10321 30855 10379 30861
rect 10321 30821 10333 30855
rect 10367 30852 10379 30855
rect 10367 30824 10548 30852
rect 10367 30821 10379 30824
rect 10321 30815 10379 30821
rect 5813 30787 5871 30793
rect 5813 30784 5825 30787
rect 5684 30756 5825 30784
rect 5684 30744 5690 30756
rect 5813 30753 5825 30756
rect 5859 30753 5871 30787
rect 5813 30747 5871 30753
rect 6365 30787 6423 30793
rect 6365 30753 6377 30787
rect 6411 30753 6423 30787
rect 6365 30747 6423 30753
rect 6549 30787 6607 30793
rect 6549 30753 6561 30787
rect 6595 30784 6607 30787
rect 7009 30787 7067 30793
rect 6595 30756 6868 30784
rect 6595 30753 6607 30756
rect 6549 30747 6607 30753
rect 6380 30716 6408 30747
rect 6380 30688 6684 30716
rect 6362 30648 6368 30660
rect 6104 30620 6368 30648
rect 6104 30589 6132 30620
rect 6362 30608 6368 30620
rect 6420 30608 6426 30660
rect 6656 30657 6684 30688
rect 6641 30651 6699 30657
rect 6641 30617 6653 30651
rect 6687 30617 6699 30651
rect 6840 30648 6868 30756
rect 7009 30753 7021 30787
rect 7055 30784 7067 30787
rect 7469 30787 7527 30793
rect 7469 30784 7481 30787
rect 7055 30756 7481 30784
rect 7055 30753 7067 30756
rect 7009 30747 7067 30753
rect 7469 30753 7481 30756
rect 7515 30753 7527 30787
rect 7469 30747 7527 30753
rect 7558 30744 7564 30796
rect 7616 30784 7622 30796
rect 8573 30787 8631 30793
rect 8573 30784 8585 30787
rect 7616 30756 8585 30784
rect 7616 30744 7622 30756
rect 8573 30753 8585 30756
rect 8619 30753 8631 30787
rect 8573 30747 8631 30753
rect 8754 30744 8760 30796
rect 8812 30784 8818 30796
rect 8849 30787 8907 30793
rect 8849 30784 8861 30787
rect 8812 30756 8861 30784
rect 8812 30744 8818 30756
rect 8849 30753 8861 30756
rect 8895 30753 8907 30787
rect 8849 30747 8907 30753
rect 10226 30744 10232 30796
rect 10284 30784 10290 30796
rect 10413 30787 10471 30793
rect 10413 30784 10425 30787
rect 10284 30756 10425 30784
rect 10284 30744 10290 30756
rect 10413 30753 10425 30756
rect 10459 30753 10471 30787
rect 10413 30747 10471 30753
rect 6914 30676 6920 30728
rect 6972 30676 6978 30728
rect 8018 30676 8024 30728
rect 8076 30676 8082 30728
rect 10520 30716 10548 30824
rect 11698 30744 11704 30796
rect 11756 30784 11762 30796
rect 11793 30787 11851 30793
rect 11793 30784 11805 30787
rect 11756 30756 11805 30784
rect 11756 30744 11762 30756
rect 11793 30753 11805 30756
rect 11839 30753 11851 30787
rect 11793 30747 11851 30753
rect 12066 30744 12072 30796
rect 12124 30784 12130 30796
rect 12161 30787 12219 30793
rect 12161 30784 12173 30787
rect 12124 30756 12173 30784
rect 12124 30744 12130 30756
rect 12161 30753 12173 30756
rect 12207 30753 12219 30787
rect 12161 30747 12219 30753
rect 12345 30787 12403 30793
rect 12345 30753 12357 30787
rect 12391 30784 12403 30787
rect 12529 30787 12587 30793
rect 12529 30784 12541 30787
rect 12391 30756 12541 30784
rect 12391 30753 12403 30756
rect 12345 30747 12403 30753
rect 12529 30753 12541 30756
rect 12575 30753 12587 30787
rect 12529 30747 12587 30753
rect 8772 30688 10548 30716
rect 8772 30660 8800 30688
rect 8754 30648 8760 30660
rect 6840 30620 8760 30648
rect 6641 30611 6699 30617
rect 8754 30608 8760 30620
rect 8812 30608 8818 30660
rect 9033 30651 9091 30657
rect 9033 30617 9045 30651
rect 9079 30648 9091 30651
rect 11238 30648 11244 30660
rect 9079 30620 11244 30648
rect 9079 30617 9091 30620
rect 9033 30611 9091 30617
rect 11238 30608 11244 30620
rect 11296 30608 11302 30660
rect 12176 30648 12204 30747
rect 12710 30676 12716 30728
rect 12768 30716 12774 30728
rect 13924 30725 13952 30892
rect 17880 30892 18460 30920
rect 16114 30812 16120 30864
rect 16172 30852 16178 30864
rect 17880 30861 17908 30892
rect 17865 30855 17923 30861
rect 16172 30824 16804 30852
rect 16172 30812 16178 30824
rect 14182 30744 14188 30796
rect 14240 30744 14246 30796
rect 14277 30787 14335 30793
rect 14277 30753 14289 30787
rect 14323 30753 14335 30787
rect 14277 30747 14335 30753
rect 13081 30719 13139 30725
rect 13081 30716 13093 30719
rect 12768 30688 13093 30716
rect 12768 30676 12774 30688
rect 13081 30685 13093 30688
rect 13127 30685 13139 30719
rect 13081 30679 13139 30685
rect 13909 30719 13967 30725
rect 13909 30685 13921 30719
rect 13955 30716 13967 30719
rect 14200 30716 14228 30744
rect 13955 30688 14228 30716
rect 14292 30716 14320 30747
rect 14642 30744 14648 30796
rect 14700 30784 14706 30796
rect 14737 30787 14795 30793
rect 14737 30784 14749 30787
rect 14700 30756 14749 30784
rect 14700 30744 14706 30756
rect 14737 30753 14749 30756
rect 14783 30753 14795 30787
rect 14737 30747 14795 30753
rect 16666 30744 16672 30796
rect 16724 30744 16730 30796
rect 16776 30793 16804 30824
rect 17865 30821 17877 30855
rect 17911 30821 17923 30855
rect 17865 30815 17923 30821
rect 17954 30812 17960 30864
rect 18012 30852 18018 30864
rect 18325 30855 18383 30861
rect 18325 30852 18337 30855
rect 18012 30824 18337 30852
rect 18012 30812 18018 30824
rect 18325 30821 18337 30824
rect 18371 30821 18383 30855
rect 18432 30852 18460 30892
rect 19426 30880 19432 30932
rect 19484 30920 19490 30932
rect 26513 30923 26571 30929
rect 26513 30920 26525 30923
rect 19484 30892 26525 30920
rect 19484 30880 19490 30892
rect 26513 30889 26525 30892
rect 26559 30889 26571 30923
rect 26513 30883 26571 30889
rect 18877 30855 18935 30861
rect 18877 30852 18889 30855
rect 18432 30824 18889 30852
rect 18325 30815 18383 30821
rect 18877 30821 18889 30824
rect 18923 30852 18935 30855
rect 19150 30852 19156 30864
rect 18923 30824 19156 30852
rect 18923 30821 18935 30824
rect 18877 30815 18935 30821
rect 19150 30812 19156 30824
rect 19208 30812 19214 30864
rect 19334 30812 19340 30864
rect 19392 30852 19398 30864
rect 20441 30855 20499 30861
rect 20441 30852 20453 30855
rect 19392 30824 20453 30852
rect 19392 30812 19398 30824
rect 20441 30821 20453 30824
rect 20487 30821 20499 30855
rect 20441 30815 20499 30821
rect 20809 30855 20867 30861
rect 20809 30821 20821 30855
rect 20855 30852 20867 30855
rect 20898 30852 20904 30864
rect 20855 30824 20904 30852
rect 20855 30821 20867 30824
rect 20809 30815 20867 30821
rect 20898 30812 20904 30824
rect 20956 30812 20962 30864
rect 22094 30812 22100 30864
rect 22152 30852 22158 30864
rect 22281 30855 22339 30861
rect 22281 30852 22293 30855
rect 22152 30824 22293 30852
rect 22152 30812 22158 30824
rect 22281 30821 22293 30824
rect 22327 30821 22339 30855
rect 22281 30815 22339 30821
rect 16761 30787 16819 30793
rect 16761 30753 16773 30787
rect 16807 30753 16819 30787
rect 16761 30747 16819 30753
rect 17678 30744 17684 30796
rect 17736 30744 17742 30796
rect 17770 30744 17776 30796
rect 17828 30744 17834 30796
rect 18046 30744 18052 30796
rect 18104 30744 18110 30796
rect 18693 30787 18751 30793
rect 18693 30753 18705 30787
rect 18739 30753 18751 30787
rect 18693 30747 18751 30753
rect 16393 30719 16451 30725
rect 14292 30688 16160 30716
rect 13955 30685 13967 30688
rect 13909 30679 13967 30685
rect 16132 30657 16160 30688
rect 16393 30685 16405 30719
rect 16439 30685 16451 30719
rect 18708 30716 18736 30747
rect 18782 30744 18788 30796
rect 18840 30784 18846 30796
rect 18969 30787 19027 30793
rect 18969 30784 18981 30787
rect 18840 30756 18981 30784
rect 18840 30744 18846 30756
rect 18969 30753 18981 30756
rect 19015 30753 19027 30787
rect 18969 30747 19027 30753
rect 19058 30744 19064 30796
rect 19116 30744 19122 30796
rect 22922 30744 22928 30796
rect 22980 30744 22986 30796
rect 23474 30744 23480 30796
rect 23532 30784 23538 30796
rect 23845 30787 23903 30793
rect 23845 30784 23857 30787
rect 23532 30756 23857 30784
rect 23532 30744 23538 30756
rect 23845 30753 23857 30756
rect 23891 30753 23903 30787
rect 23845 30747 23903 30753
rect 26418 30744 26424 30796
rect 26476 30784 26482 30796
rect 26697 30787 26755 30793
rect 26697 30784 26709 30787
rect 26476 30756 26709 30784
rect 26476 30744 26482 30756
rect 26697 30753 26709 30756
rect 26743 30753 26755 30787
rect 26697 30747 26755 30753
rect 19521 30719 19579 30725
rect 19521 30716 19533 30719
rect 18708 30688 19533 30716
rect 16393 30679 16451 30685
rect 19521 30685 19533 30688
rect 19567 30685 19579 30719
rect 19521 30679 19579 30685
rect 20165 30719 20223 30725
rect 20165 30685 20177 30719
rect 20211 30716 20223 30719
rect 20438 30716 20444 30728
rect 20211 30688 20444 30716
rect 20211 30685 20223 30688
rect 20165 30679 20223 30685
rect 14112 30651 14170 30657
rect 14112 30648 14124 30651
rect 12176 30620 14124 30648
rect 14112 30617 14124 30620
rect 14158 30617 14170 30651
rect 14112 30611 14170 30617
rect 16117 30651 16175 30657
rect 16117 30617 16129 30651
rect 16163 30617 16175 30651
rect 16117 30611 16175 30617
rect 6089 30583 6147 30589
rect 6089 30549 6101 30583
rect 6135 30549 6147 30583
rect 6089 30543 6147 30549
rect 6270 30540 6276 30592
rect 6328 30540 6334 30592
rect 6457 30583 6515 30589
rect 6457 30549 6469 30583
rect 6503 30580 6515 30583
rect 6914 30580 6920 30592
rect 6503 30552 6920 30580
rect 6503 30549 6515 30552
rect 6457 30543 6515 30549
rect 6914 30540 6920 30552
rect 6972 30540 6978 30592
rect 9674 30540 9680 30592
rect 9732 30580 9738 30592
rect 9953 30583 10011 30589
rect 9953 30580 9965 30583
rect 9732 30552 9965 30580
rect 9732 30540 9738 30552
rect 9953 30549 9965 30552
rect 9999 30549 10011 30583
rect 9953 30543 10011 30549
rect 10137 30583 10195 30589
rect 10137 30549 10149 30583
rect 10183 30580 10195 30583
rect 10318 30580 10324 30592
rect 10183 30552 10324 30580
rect 10183 30549 10195 30552
rect 10137 30543 10195 30549
rect 10318 30540 10324 30552
rect 10376 30540 10382 30592
rect 10597 30583 10655 30589
rect 10597 30549 10609 30583
rect 10643 30580 10655 30583
rect 11054 30580 11060 30592
rect 10643 30552 11060 30580
rect 10643 30549 10655 30552
rect 10597 30543 10655 30549
rect 11054 30540 11060 30552
rect 11112 30540 11118 30592
rect 11698 30540 11704 30592
rect 11756 30580 11762 30592
rect 12253 30583 12311 30589
rect 12253 30580 12265 30583
rect 11756 30552 12265 30580
rect 11756 30540 11762 30552
rect 12253 30549 12265 30552
rect 12299 30549 12311 30583
rect 12253 30543 12311 30549
rect 13630 30540 13636 30592
rect 13688 30540 13694 30592
rect 13998 30540 14004 30592
rect 14056 30540 14062 30592
rect 14734 30540 14740 30592
rect 14792 30580 14798 30592
rect 14921 30583 14979 30589
rect 14921 30580 14933 30583
rect 14792 30552 14933 30580
rect 14792 30540 14798 30552
rect 14921 30549 14933 30552
rect 14967 30580 14979 30583
rect 16408 30580 16436 30679
rect 20438 30676 20444 30688
rect 20496 30676 20502 30728
rect 23566 30676 23572 30728
rect 23624 30716 23630 30728
rect 24121 30719 24179 30725
rect 24121 30716 24133 30719
rect 23624 30688 24133 30716
rect 23624 30676 23630 30688
rect 24121 30685 24133 30688
rect 24167 30685 24179 30719
rect 24121 30679 24179 30685
rect 19168 30620 19380 30648
rect 14967 30552 16436 30580
rect 16577 30583 16635 30589
rect 14967 30549 14979 30552
rect 14921 30543 14979 30549
rect 16577 30549 16589 30583
rect 16623 30580 16635 30583
rect 16758 30580 16764 30592
rect 16623 30552 16764 30580
rect 16623 30549 16635 30552
rect 16577 30543 16635 30549
rect 16758 30540 16764 30552
rect 16816 30580 16822 30592
rect 16945 30583 17003 30589
rect 16945 30580 16957 30583
rect 16816 30552 16957 30580
rect 16816 30540 16822 30552
rect 16945 30549 16957 30552
rect 16991 30549 17003 30583
rect 16945 30543 17003 30549
rect 17497 30583 17555 30589
rect 17497 30549 17509 30583
rect 17543 30580 17555 30583
rect 17586 30580 17592 30592
rect 17543 30552 17592 30580
rect 17543 30549 17555 30552
rect 17497 30543 17555 30549
rect 17586 30540 17592 30552
rect 17644 30540 17650 30592
rect 17770 30540 17776 30592
rect 17828 30580 17834 30592
rect 18233 30583 18291 30589
rect 18233 30580 18245 30583
rect 17828 30552 18245 30580
rect 17828 30540 17834 30552
rect 18233 30549 18245 30552
rect 18279 30549 18291 30583
rect 18233 30543 18291 30549
rect 18690 30540 18696 30592
rect 18748 30580 18754 30592
rect 19168 30580 19196 30620
rect 18748 30552 19196 30580
rect 18748 30540 18754 30552
rect 19242 30540 19248 30592
rect 19300 30540 19306 30592
rect 19352 30580 19380 30620
rect 19426 30608 19432 30660
rect 19484 30648 19490 30660
rect 20625 30651 20683 30657
rect 20625 30648 20637 30651
rect 19484 30620 20637 30648
rect 19484 30608 19490 30620
rect 20625 30617 20637 30620
rect 20671 30617 20683 30651
rect 20625 30611 20683 30617
rect 20349 30583 20407 30589
rect 20349 30580 20361 30583
rect 19352 30552 20361 30580
rect 20349 30549 20361 30552
rect 20395 30549 20407 30583
rect 20349 30543 20407 30549
rect 22189 30583 22247 30589
rect 22189 30549 22201 30583
rect 22235 30580 22247 30583
rect 22370 30580 22376 30592
rect 22235 30552 22376 30580
rect 22235 30549 22247 30552
rect 22189 30543 22247 30549
rect 22370 30540 22376 30552
rect 22428 30540 22434 30592
rect 22554 30540 22560 30592
rect 22612 30580 22618 30592
rect 22741 30583 22799 30589
rect 22741 30580 22753 30583
rect 22612 30552 22753 30580
rect 22612 30540 22618 30552
rect 22741 30549 22753 30552
rect 22787 30549 22799 30583
rect 22741 30543 22799 30549
rect 552 30490 27416 30512
rect 552 30438 3756 30490
rect 3808 30438 3820 30490
rect 3872 30438 3884 30490
rect 3936 30438 3948 30490
rect 4000 30438 4012 30490
rect 4064 30438 10472 30490
rect 10524 30438 10536 30490
rect 10588 30438 10600 30490
rect 10652 30438 10664 30490
rect 10716 30438 10728 30490
rect 10780 30438 17188 30490
rect 17240 30438 17252 30490
rect 17304 30438 17316 30490
rect 17368 30438 17380 30490
rect 17432 30438 17444 30490
rect 17496 30438 23904 30490
rect 23956 30438 23968 30490
rect 24020 30438 24032 30490
rect 24084 30438 24096 30490
rect 24148 30438 24160 30490
rect 24212 30438 27416 30490
rect 552 30416 27416 30438
rect 8018 30336 8024 30388
rect 8076 30336 8082 30388
rect 11149 30379 11207 30385
rect 11149 30345 11161 30379
rect 11195 30376 11207 30379
rect 12066 30376 12072 30388
rect 11195 30348 12072 30376
rect 11195 30345 11207 30348
rect 11149 30339 11207 30345
rect 12066 30336 12072 30348
rect 12124 30336 12130 30388
rect 12710 30336 12716 30388
rect 12768 30336 12774 30388
rect 4338 30268 4344 30320
rect 4396 30308 4402 30320
rect 4617 30311 4675 30317
rect 4617 30308 4629 30311
rect 4396 30280 4629 30308
rect 4396 30268 4402 30280
rect 4617 30277 4629 30280
rect 4663 30277 4675 30311
rect 4617 30271 4675 30277
rect 16022 30268 16028 30320
rect 16080 30268 16086 30320
rect 17865 30311 17923 30317
rect 17865 30277 17877 30311
rect 17911 30308 17923 30311
rect 18046 30308 18052 30320
rect 17911 30280 18052 30308
rect 17911 30277 17923 30280
rect 17865 30271 17923 30277
rect 18046 30268 18052 30280
rect 18104 30268 18110 30320
rect 20257 30311 20315 30317
rect 20257 30277 20269 30311
rect 20303 30277 20315 30311
rect 20257 30271 20315 30277
rect 21177 30311 21235 30317
rect 21177 30277 21189 30311
rect 21223 30308 21235 30311
rect 21542 30308 21548 30320
rect 21223 30280 21548 30308
rect 21223 30277 21235 30280
rect 21177 30271 21235 30277
rect 6454 30200 6460 30252
rect 6512 30240 6518 30252
rect 6641 30243 6699 30249
rect 6641 30240 6653 30243
rect 6512 30212 6653 30240
rect 6512 30200 6518 30212
rect 6641 30209 6653 30212
rect 6687 30209 6699 30243
rect 6641 30203 6699 30209
rect 8478 30200 8484 30252
rect 8536 30240 8542 30252
rect 9493 30243 9551 30249
rect 9493 30240 9505 30243
rect 8536 30212 9505 30240
rect 8536 30200 8542 30212
rect 9493 30209 9505 30212
rect 9539 30209 9551 30243
rect 11330 30240 11336 30252
rect 9493 30203 9551 30209
rect 10980 30212 11336 30240
rect 3053 30175 3111 30181
rect 3053 30141 3065 30175
rect 3099 30172 3111 30175
rect 3234 30172 3240 30184
rect 3099 30144 3240 30172
rect 3099 30141 3111 30144
rect 3053 30135 3111 30141
rect 3234 30132 3240 30144
rect 3292 30132 3298 30184
rect 4801 30175 4859 30181
rect 4801 30141 4813 30175
rect 4847 30172 4859 30175
rect 5534 30172 5540 30184
rect 4847 30144 5540 30172
rect 4847 30141 4859 30144
rect 4801 30135 4859 30141
rect 5534 30132 5540 30144
rect 5592 30172 5598 30184
rect 6472 30172 6500 30200
rect 6914 30181 6920 30184
rect 5592 30144 6500 30172
rect 6549 30175 6607 30181
rect 5592 30132 5598 30144
rect 6549 30141 6561 30175
rect 6595 30141 6607 30175
rect 6908 30172 6920 30181
rect 6875 30144 6920 30172
rect 6549 30135 6607 30141
rect 6908 30135 6920 30144
rect 2774 30064 2780 30116
rect 2832 30113 2838 30116
rect 2832 30067 2844 30113
rect 3504 30107 3562 30113
rect 3504 30073 3516 30107
rect 3550 30073 3562 30107
rect 3504 30067 3562 30073
rect 2832 30064 2838 30067
rect 1673 30039 1731 30045
rect 1673 30005 1685 30039
rect 1719 30036 1731 30039
rect 2958 30036 2964 30048
rect 1719 30008 2964 30036
rect 1719 30005 1731 30008
rect 1673 29999 1731 30005
rect 2958 29996 2964 30008
rect 3016 29996 3022 30048
rect 3418 29996 3424 30048
rect 3476 30036 3482 30048
rect 3528 30036 3556 30067
rect 4338 30064 4344 30116
rect 4396 30104 4402 30116
rect 5046 30107 5104 30113
rect 5046 30104 5058 30107
rect 4396 30076 5058 30104
rect 4396 30064 4402 30076
rect 5046 30073 5058 30076
rect 5092 30073 5104 30107
rect 5046 30067 5104 30073
rect 5810 30064 5816 30116
rect 5868 30104 5874 30116
rect 6564 30104 6592 30135
rect 6914 30132 6920 30135
rect 6972 30132 6978 30184
rect 8294 30132 8300 30184
rect 8352 30172 8358 30184
rect 8389 30175 8447 30181
rect 8389 30172 8401 30175
rect 8352 30144 8401 30172
rect 8352 30132 8358 30144
rect 8389 30141 8401 30144
rect 8435 30141 8447 30175
rect 8389 30135 8447 30141
rect 8573 30175 8631 30181
rect 8573 30141 8585 30175
rect 8619 30141 8631 30175
rect 8573 30135 8631 30141
rect 5868 30076 6592 30104
rect 8588 30104 8616 30135
rect 8846 30132 8852 30184
rect 8904 30132 8910 30184
rect 9122 30132 9128 30184
rect 9180 30132 9186 30184
rect 9217 30175 9275 30181
rect 9217 30141 9229 30175
rect 9263 30172 9275 30175
rect 9398 30172 9404 30184
rect 9263 30144 9404 30172
rect 9263 30141 9275 30144
rect 9217 30135 9275 30141
rect 9398 30132 9404 30144
rect 9456 30132 9462 30184
rect 9508 30172 9536 30203
rect 10980 30172 11008 30212
rect 11330 30200 11336 30212
rect 11388 30200 11394 30252
rect 20272 30240 20300 30271
rect 21542 30268 21548 30280
rect 21600 30268 21606 30320
rect 21913 30311 21971 30317
rect 21913 30277 21925 30311
rect 21959 30308 21971 30311
rect 21959 30280 22094 30308
rect 21959 30277 21971 30280
rect 21913 30271 21971 30277
rect 20438 30240 20444 30252
rect 20272 30212 20444 30240
rect 20438 30200 20444 30212
rect 20496 30200 20502 30252
rect 20901 30243 20959 30249
rect 20901 30209 20913 30243
rect 20947 30240 20959 30243
rect 21818 30240 21824 30252
rect 20947 30212 21824 30240
rect 20947 30209 20959 30212
rect 20901 30203 20959 30209
rect 21818 30200 21824 30212
rect 21876 30200 21882 30252
rect 9508 30144 11008 30172
rect 11054 30132 11060 30184
rect 11112 30132 11118 30184
rect 11238 30132 11244 30184
rect 11296 30132 11302 30184
rect 13081 30175 13139 30181
rect 13081 30141 13093 30175
rect 13127 30172 13139 30175
rect 13170 30172 13176 30184
rect 13127 30144 13176 30172
rect 13127 30141 13139 30144
rect 13081 30135 13139 30141
rect 13170 30132 13176 30144
rect 13228 30132 13234 30184
rect 13722 30132 13728 30184
rect 13780 30132 13786 30184
rect 15289 30175 15347 30181
rect 15289 30141 15301 30175
rect 15335 30141 15347 30175
rect 15289 30135 15347 30141
rect 9738 30107 9796 30113
rect 9738 30104 9750 30107
rect 8588 30076 9076 30104
rect 5868 30064 5874 30076
rect 3476 30008 3556 30036
rect 3476 29996 3482 30008
rect 6086 29996 6092 30048
rect 6144 30036 6150 30048
rect 6181 30039 6239 30045
rect 6181 30036 6193 30039
rect 6144 30008 6193 30036
rect 6144 29996 6150 30008
rect 6181 30005 6193 30008
rect 6227 30005 6239 30039
rect 6181 29999 6239 30005
rect 6362 29996 6368 30048
rect 6420 29996 6426 30048
rect 8570 29996 8576 30048
rect 8628 29996 8634 30048
rect 8662 29996 8668 30048
rect 8720 29996 8726 30048
rect 9048 30045 9076 30076
rect 9416 30076 9750 30104
rect 9033 30039 9091 30045
rect 9033 30005 9045 30039
rect 9079 30036 9091 30039
rect 9306 30036 9312 30048
rect 9079 30008 9312 30036
rect 9079 30005 9091 30008
rect 9033 29999 9091 30005
rect 9306 29996 9312 30008
rect 9364 29996 9370 30048
rect 9416 30045 9444 30076
rect 9738 30073 9750 30076
rect 9784 30073 9796 30107
rect 9738 30067 9796 30073
rect 11422 30064 11428 30116
rect 11480 30104 11486 30116
rect 11578 30107 11636 30113
rect 11578 30104 11590 30107
rect 11480 30076 11590 30104
rect 11480 30064 11486 30076
rect 11578 30073 11590 30076
rect 11624 30073 11636 30107
rect 13998 30104 14004 30116
rect 11578 30067 11636 30073
rect 13280 30076 14004 30104
rect 9401 30039 9459 30045
rect 9401 30005 9413 30039
rect 9447 30005 9459 30039
rect 9401 29999 9459 30005
rect 10594 29996 10600 30048
rect 10652 30036 10658 30048
rect 10870 30036 10876 30048
rect 10652 30008 10876 30036
rect 10652 29996 10658 30008
rect 10870 29996 10876 30008
rect 10928 29996 10934 30048
rect 13170 29996 13176 30048
rect 13228 30036 13234 30048
rect 13280 30045 13308 30076
rect 13998 30064 14004 30076
rect 14056 30064 14062 30116
rect 15044 30107 15102 30113
rect 15044 30073 15056 30107
rect 15090 30104 15102 30107
rect 15304 30104 15332 30135
rect 15378 30132 15384 30184
rect 15436 30172 15442 30184
rect 15565 30175 15623 30181
rect 15565 30172 15577 30175
rect 15436 30144 15577 30172
rect 15436 30132 15442 30144
rect 15565 30141 15577 30144
rect 15611 30141 15623 30175
rect 15565 30135 15623 30141
rect 15749 30175 15807 30181
rect 15749 30141 15761 30175
rect 15795 30172 15807 30175
rect 16114 30172 16120 30184
rect 15795 30144 16120 30172
rect 15795 30141 15807 30144
rect 15749 30135 15807 30141
rect 16114 30132 16120 30144
rect 16172 30132 16178 30184
rect 17405 30175 17463 30181
rect 17405 30172 17417 30175
rect 16868 30144 17417 30172
rect 16868 30116 16896 30144
rect 17405 30141 17417 30144
rect 17451 30141 17463 30175
rect 17405 30135 17463 30141
rect 18506 30132 18512 30184
rect 18564 30132 18570 30184
rect 18877 30175 18935 30181
rect 18877 30141 18889 30175
rect 18923 30172 18935 30175
rect 20533 30175 20591 30181
rect 18923 30144 19380 30172
rect 18923 30141 18935 30144
rect 18877 30135 18935 30141
rect 19352 30116 19380 30144
rect 20533 30141 20545 30175
rect 20579 30141 20591 30175
rect 20533 30135 20591 30141
rect 21453 30175 21511 30181
rect 21453 30141 21465 30175
rect 21499 30172 21511 30175
rect 22066 30172 22094 30280
rect 23658 30268 23664 30320
rect 23716 30308 23722 30320
rect 24121 30311 24179 30317
rect 24121 30308 24133 30311
rect 23716 30280 24133 30308
rect 23716 30268 23722 30280
rect 24121 30277 24133 30280
rect 24167 30277 24179 30311
rect 24121 30271 24179 30277
rect 24394 30240 24400 30252
rect 23768 30212 24400 30240
rect 21499 30144 22094 30172
rect 21499 30141 21511 30144
rect 21453 30135 21511 30141
rect 16850 30104 16856 30116
rect 15090 30076 15240 30104
rect 15304 30076 16856 30104
rect 15090 30073 15102 30076
rect 15044 30067 15102 30073
rect 13265 30039 13323 30045
rect 13265 30036 13277 30039
rect 13228 30008 13277 30036
rect 13228 29996 13234 30008
rect 13265 30005 13277 30008
rect 13311 30005 13323 30039
rect 13265 29999 13323 30005
rect 13538 29996 13544 30048
rect 13596 29996 13602 30048
rect 13909 30039 13967 30045
rect 13909 30005 13921 30039
rect 13955 30036 13967 30039
rect 14550 30036 14556 30048
rect 13955 30008 14556 30036
rect 13955 30005 13967 30008
rect 13909 29999 13967 30005
rect 14550 29996 14556 30008
rect 14608 29996 14614 30048
rect 15212 30036 15240 30076
rect 16850 30064 16856 30076
rect 16908 30064 16914 30116
rect 17138 30107 17196 30113
rect 17138 30104 17150 30107
rect 16960 30076 17150 30104
rect 15381 30039 15439 30045
rect 15381 30036 15393 30039
rect 15212 30008 15393 30036
rect 15381 30005 15393 30008
rect 15427 30005 15439 30039
rect 15381 29999 15439 30005
rect 15933 30039 15991 30045
rect 15933 30005 15945 30039
rect 15979 30036 15991 30039
rect 16960 30036 16988 30076
rect 17138 30073 17150 30076
rect 17184 30073 17196 30107
rect 17138 30067 17196 30073
rect 19144 30107 19202 30113
rect 19144 30073 19156 30107
rect 19190 30104 19202 30107
rect 19242 30104 19248 30116
rect 19190 30076 19248 30104
rect 19190 30073 19202 30076
rect 19144 30067 19202 30073
rect 19242 30064 19248 30076
rect 19300 30064 19306 30116
rect 19334 30064 19340 30116
rect 19392 30064 19398 30116
rect 20548 30104 20576 30135
rect 20548 30076 21496 30104
rect 21468 30048 21496 30076
rect 21542 30064 21548 30116
rect 21600 30064 21606 30116
rect 22066 30104 22094 30144
rect 22278 30132 22284 30184
rect 22336 30132 22342 30184
rect 22554 30181 22560 30184
rect 22548 30172 22560 30181
rect 22515 30144 22560 30172
rect 22548 30135 22560 30144
rect 22554 30132 22560 30135
rect 22612 30132 22618 30184
rect 23768 30104 23796 30212
rect 24394 30200 24400 30212
rect 24452 30200 24458 30252
rect 23845 30175 23903 30181
rect 23845 30141 23857 30175
rect 23891 30172 23903 30175
rect 24118 30172 24124 30184
rect 23891 30144 24124 30172
rect 23891 30141 23903 30144
rect 23845 30135 23903 30141
rect 24118 30132 24124 30144
rect 24176 30132 24182 30184
rect 25498 30132 25504 30184
rect 25556 30132 25562 30184
rect 25234 30107 25292 30113
rect 25234 30104 25246 30107
rect 22066 30076 23796 30104
rect 24044 30076 25246 30104
rect 15979 30008 16988 30036
rect 20993 30039 21051 30045
rect 15979 30005 15991 30008
rect 15933 29999 15991 30005
rect 20993 30005 21005 30039
rect 21039 30036 21051 30039
rect 21358 30036 21364 30048
rect 21039 30008 21364 30036
rect 21039 30005 21051 30008
rect 20993 29999 21051 30005
rect 21358 29996 21364 30008
rect 21416 29996 21422 30048
rect 21450 29996 21456 30048
rect 21508 29996 21514 30048
rect 22002 29996 22008 30048
rect 22060 29996 22066 30048
rect 23198 29996 23204 30048
rect 23256 30036 23262 30048
rect 24044 30045 24072 30076
rect 25234 30073 25246 30076
rect 25280 30073 25292 30107
rect 25234 30067 25292 30073
rect 23661 30039 23719 30045
rect 23661 30036 23673 30039
rect 23256 30008 23673 30036
rect 23256 29996 23262 30008
rect 23661 30005 23673 30008
rect 23707 30005 23719 30039
rect 23661 29999 23719 30005
rect 24029 30039 24087 30045
rect 24029 30005 24041 30039
rect 24075 30005 24087 30039
rect 24029 29999 24087 30005
rect 552 29946 27576 29968
rect 552 29894 7114 29946
rect 7166 29894 7178 29946
rect 7230 29894 7242 29946
rect 7294 29894 7306 29946
rect 7358 29894 7370 29946
rect 7422 29894 13830 29946
rect 13882 29894 13894 29946
rect 13946 29894 13958 29946
rect 14010 29894 14022 29946
rect 14074 29894 14086 29946
rect 14138 29894 20546 29946
rect 20598 29894 20610 29946
rect 20662 29894 20674 29946
rect 20726 29894 20738 29946
rect 20790 29894 20802 29946
rect 20854 29894 27262 29946
rect 27314 29894 27326 29946
rect 27378 29894 27390 29946
rect 27442 29894 27454 29946
rect 27506 29894 27518 29946
rect 27570 29894 27576 29946
rect 552 29872 27576 29894
rect 937 29835 995 29841
rect 937 29801 949 29835
rect 983 29832 995 29835
rect 1394 29832 1400 29844
rect 983 29804 1400 29832
rect 983 29801 995 29804
rect 937 29795 995 29801
rect 1394 29792 1400 29804
rect 1452 29792 1458 29844
rect 4338 29792 4344 29844
rect 4396 29792 4402 29844
rect 9122 29792 9128 29844
rect 9180 29832 9186 29844
rect 9401 29835 9459 29841
rect 9401 29832 9413 29835
rect 9180 29804 9413 29832
rect 9180 29792 9186 29804
rect 9401 29801 9413 29804
rect 9447 29801 9459 29835
rect 9401 29795 9459 29801
rect 10134 29792 10140 29844
rect 10192 29792 10198 29844
rect 10318 29792 10324 29844
rect 10376 29832 10382 29844
rect 10597 29835 10655 29841
rect 10597 29832 10609 29835
rect 10376 29804 10609 29832
rect 10376 29792 10382 29804
rect 10597 29801 10609 29804
rect 10643 29801 10655 29835
rect 10597 29795 10655 29801
rect 11054 29792 11060 29844
rect 11112 29832 11118 29844
rect 11885 29835 11943 29841
rect 11885 29832 11897 29835
rect 11112 29804 11897 29832
rect 11112 29792 11118 29804
rect 11885 29801 11897 29804
rect 11931 29801 11943 29835
rect 11885 29795 11943 29801
rect 11977 29835 12035 29841
rect 11977 29801 11989 29835
rect 12023 29832 12035 29835
rect 12710 29832 12716 29844
rect 12023 29804 12716 29832
rect 12023 29801 12035 29804
rect 11977 29795 12035 29801
rect 12710 29792 12716 29804
rect 12768 29792 12774 29844
rect 14550 29792 14556 29844
rect 14608 29832 14614 29844
rect 15102 29832 15108 29844
rect 14608 29804 15108 29832
rect 14608 29792 14614 29804
rect 15102 29792 15108 29804
rect 15160 29832 15166 29844
rect 15160 29804 15332 29832
rect 15160 29792 15166 29804
rect 3234 29724 3240 29776
rect 3292 29764 3298 29776
rect 3510 29764 3516 29776
rect 3292 29736 3516 29764
rect 3292 29724 3298 29736
rect 3510 29724 3516 29736
rect 3568 29764 3574 29776
rect 4617 29767 4675 29773
rect 4617 29764 4629 29767
rect 3568 29736 4629 29764
rect 3568 29724 3574 29736
rect 4617 29733 4629 29736
rect 4663 29764 4675 29767
rect 5534 29764 5540 29776
rect 4663 29736 5540 29764
rect 4663 29733 4675 29736
rect 4617 29727 4675 29733
rect 5534 29724 5540 29736
rect 5592 29724 5598 29776
rect 8938 29764 8944 29776
rect 5736 29736 8944 29764
rect 2061 29699 2119 29705
rect 2061 29665 2073 29699
rect 2107 29696 2119 29699
rect 2317 29699 2375 29705
rect 2107 29668 2268 29696
rect 2107 29665 2119 29668
rect 2061 29659 2119 29665
rect 2240 29628 2268 29668
rect 2317 29665 2329 29699
rect 2363 29696 2375 29699
rect 3252 29696 3280 29724
rect 2363 29668 3280 29696
rect 2363 29665 2375 29668
rect 2317 29659 2375 29665
rect 3326 29656 3332 29708
rect 3384 29696 3390 29708
rect 3789 29699 3847 29705
rect 3789 29696 3801 29699
rect 3384 29668 3801 29696
rect 3384 29656 3390 29668
rect 3789 29665 3801 29668
rect 3835 29665 3847 29699
rect 3789 29659 3847 29665
rect 3973 29699 4031 29705
rect 3973 29665 3985 29699
rect 4019 29665 4031 29699
rect 3973 29659 4031 29665
rect 3988 29628 4016 29659
rect 4154 29656 4160 29708
rect 4212 29656 4218 29708
rect 5353 29699 5411 29705
rect 5353 29665 5365 29699
rect 5399 29696 5411 29699
rect 5736 29696 5764 29736
rect 8938 29724 8944 29736
rect 8996 29724 9002 29776
rect 10336 29736 10640 29764
rect 5399 29668 5764 29696
rect 5399 29665 5411 29668
rect 5353 29659 5411 29665
rect 5994 29656 6000 29708
rect 6052 29656 6058 29708
rect 6270 29656 6276 29708
rect 6328 29656 6334 29708
rect 6546 29656 6552 29708
rect 6604 29656 6610 29708
rect 7006 29656 7012 29708
rect 7064 29656 7070 29708
rect 8288 29699 8346 29705
rect 8288 29665 8300 29699
rect 8334 29696 8346 29699
rect 8662 29696 8668 29708
rect 8334 29668 8668 29696
rect 8334 29665 8346 29668
rect 8288 29659 8346 29665
rect 8662 29656 8668 29668
rect 8720 29656 8726 29708
rect 10336 29705 10364 29736
rect 10612 29708 10640 29736
rect 11238 29724 11244 29776
rect 11296 29764 11302 29776
rect 11609 29767 11667 29773
rect 11609 29764 11621 29767
rect 11296 29736 11621 29764
rect 11296 29724 11302 29736
rect 11609 29733 11621 29736
rect 11655 29733 11667 29767
rect 11609 29727 11667 29733
rect 12980 29767 13038 29773
rect 12980 29733 12992 29767
rect 13026 29764 13038 29767
rect 13538 29764 13544 29776
rect 13026 29736 13544 29764
rect 13026 29733 13038 29736
rect 12980 29727 13038 29733
rect 13538 29724 13544 29736
rect 13596 29724 13602 29776
rect 14369 29767 14427 29773
rect 14369 29733 14381 29767
rect 14415 29764 14427 29767
rect 14415 29736 14688 29764
rect 14415 29733 14427 29736
rect 14369 29727 14427 29733
rect 10321 29699 10379 29705
rect 10321 29665 10333 29699
rect 10367 29665 10379 29699
rect 10321 29659 10379 29665
rect 10505 29699 10563 29705
rect 10505 29665 10517 29699
rect 10551 29665 10563 29699
rect 10505 29659 10563 29665
rect 5810 29628 5816 29640
rect 2240 29600 2544 29628
rect 3988 29600 5816 29628
rect 2516 29504 2544 29600
rect 5810 29588 5816 29600
rect 5868 29588 5874 29640
rect 6822 29588 6828 29640
rect 6880 29588 6886 29640
rect 8021 29631 8079 29637
rect 8021 29597 8033 29631
rect 8067 29597 8079 29631
rect 8021 29591 8079 29597
rect 2498 29452 2504 29504
rect 2556 29492 2562 29504
rect 2593 29495 2651 29501
rect 2593 29492 2605 29495
rect 2556 29464 2605 29492
rect 2556 29452 2562 29464
rect 2593 29461 2605 29464
rect 2639 29461 2651 29495
rect 2593 29455 2651 29461
rect 3602 29452 3608 29504
rect 3660 29492 3666 29504
rect 3881 29495 3939 29501
rect 3881 29492 3893 29495
rect 3660 29464 3893 29492
rect 3660 29452 3666 29464
rect 3881 29461 3893 29464
rect 3927 29461 3939 29495
rect 8036 29492 8064 29591
rect 10042 29588 10048 29640
rect 10100 29628 10106 29640
rect 10520 29628 10548 29659
rect 10594 29656 10600 29708
rect 10652 29656 10658 29708
rect 10781 29699 10839 29705
rect 10781 29665 10793 29699
rect 10827 29665 10839 29699
rect 10781 29659 10839 29665
rect 11333 29699 11391 29705
rect 11333 29665 11345 29699
rect 11379 29696 11391 29699
rect 12069 29699 12127 29705
rect 12069 29696 12081 29699
rect 11379 29668 12081 29696
rect 11379 29665 11391 29668
rect 11333 29659 11391 29665
rect 12069 29665 12081 29668
rect 12115 29696 12127 29699
rect 12115 29668 12434 29696
rect 12115 29665 12127 29668
rect 12069 29659 12127 29665
rect 10796 29628 10824 29659
rect 10100 29600 10824 29628
rect 12406 29628 12434 29668
rect 14550 29656 14556 29708
rect 14608 29656 14614 29708
rect 14660 29696 14688 29736
rect 15194 29724 15200 29776
rect 15252 29724 15258 29776
rect 15304 29764 15332 29804
rect 15378 29792 15384 29844
rect 15436 29792 15442 29844
rect 16114 29792 16120 29844
rect 16172 29792 16178 29844
rect 18506 29792 18512 29844
rect 18564 29832 18570 29844
rect 18693 29835 18751 29841
rect 18693 29832 18705 29835
rect 18564 29804 18705 29832
rect 18564 29792 18570 29804
rect 18693 29801 18705 29804
rect 18739 29832 18751 29835
rect 21542 29832 21548 29844
rect 18739 29804 21548 29832
rect 18739 29801 18751 29804
rect 18693 29795 18751 29801
rect 21542 29792 21548 29804
rect 21600 29792 21606 29844
rect 23658 29832 23664 29844
rect 22296 29804 23664 29832
rect 16301 29767 16359 29773
rect 15304 29736 15792 29764
rect 15764 29705 15792 29736
rect 16301 29733 16313 29767
rect 16347 29733 16359 29767
rect 16301 29727 16359 29733
rect 15657 29699 15715 29705
rect 15657 29696 15669 29699
rect 14660 29668 15669 29696
rect 15212 29640 15240 29668
rect 15657 29665 15669 29668
rect 15703 29665 15715 29699
rect 15657 29659 15715 29665
rect 15749 29699 15807 29705
rect 15749 29665 15761 29699
rect 15795 29665 15807 29699
rect 15749 29659 15807 29665
rect 12526 29628 12532 29640
rect 12406 29600 12532 29628
rect 10100 29588 10106 29600
rect 12526 29588 12532 29600
rect 12584 29588 12590 29640
rect 12618 29588 12624 29640
rect 12676 29628 12682 29640
rect 12713 29631 12771 29637
rect 12713 29628 12725 29631
rect 12676 29600 12725 29628
rect 12676 29588 12682 29600
rect 12713 29597 12725 29600
rect 12759 29597 12771 29631
rect 12713 29591 12771 29597
rect 15194 29588 15200 29640
rect 15252 29588 15258 29640
rect 15378 29588 15384 29640
rect 15436 29628 15442 29640
rect 16316 29628 16344 29727
rect 16758 29724 16764 29776
rect 16816 29764 16822 29776
rect 16853 29767 16911 29773
rect 16853 29764 16865 29767
rect 16816 29736 16865 29764
rect 16816 29724 16822 29736
rect 16853 29733 16865 29736
rect 16899 29733 16911 29767
rect 16853 29727 16911 29733
rect 17328 29736 18828 29764
rect 17328 29637 17356 29736
rect 17586 29705 17592 29708
rect 17580 29696 17592 29705
rect 17547 29668 17592 29696
rect 17580 29659 17592 29668
rect 17586 29656 17592 29659
rect 17644 29656 17650 29708
rect 18800 29705 18828 29736
rect 21358 29724 21364 29776
rect 21416 29764 21422 29776
rect 22296 29773 22324 29804
rect 23658 29792 23664 29804
rect 23716 29792 23722 29844
rect 24118 29792 24124 29844
rect 24176 29792 24182 29844
rect 22281 29767 22339 29773
rect 22281 29764 22293 29767
rect 21416 29736 21956 29764
rect 21416 29724 21422 29736
rect 18785 29699 18843 29705
rect 18785 29665 18797 29699
rect 18831 29665 18843 29699
rect 18785 29659 18843 29665
rect 18874 29656 18880 29708
rect 18932 29696 18938 29708
rect 19041 29699 19099 29705
rect 19041 29696 19053 29699
rect 18932 29668 19053 29696
rect 18932 29656 18938 29668
rect 19041 29665 19053 29668
rect 19087 29665 19099 29699
rect 19041 29659 19099 29665
rect 20438 29656 20444 29708
rect 20496 29696 20502 29708
rect 20496 29668 21404 29696
rect 20496 29656 20502 29668
rect 21376 29637 21404 29668
rect 21450 29656 21456 29708
rect 21508 29696 21514 29708
rect 21508 29668 21680 29696
rect 21508 29656 21514 29668
rect 17313 29631 17371 29637
rect 17313 29628 17325 29631
rect 15436 29600 16344 29628
rect 16868 29600 17325 29628
rect 15436 29588 15442 29600
rect 16868 29572 16896 29600
rect 17313 29597 17325 29600
rect 17359 29597 17371 29631
rect 20809 29631 20867 29637
rect 20809 29628 20821 29631
rect 17313 29591 17371 29597
rect 20180 29600 20821 29628
rect 14829 29563 14887 29569
rect 14829 29529 14841 29563
rect 14875 29560 14887 29563
rect 15286 29560 15292 29572
rect 14875 29532 15292 29560
rect 14875 29529 14887 29532
rect 14829 29523 14887 29529
rect 15286 29520 15292 29532
rect 15344 29560 15350 29572
rect 15473 29563 15531 29569
rect 15473 29560 15485 29563
rect 15344 29532 15485 29560
rect 15344 29520 15350 29532
rect 15473 29529 15485 29532
rect 15519 29529 15531 29563
rect 15473 29523 15531 29529
rect 16574 29520 16580 29572
rect 16632 29560 16638 29572
rect 16669 29563 16727 29569
rect 16669 29560 16681 29563
rect 16632 29532 16681 29560
rect 16632 29520 16638 29532
rect 16669 29529 16681 29532
rect 16715 29529 16727 29563
rect 16669 29523 16727 29529
rect 16850 29520 16856 29572
rect 16908 29520 16914 29572
rect 20070 29520 20076 29572
rect 20128 29560 20134 29572
rect 20180 29569 20208 29600
rect 20809 29597 20821 29600
rect 20855 29597 20867 29631
rect 20809 29591 20867 29597
rect 21361 29631 21419 29637
rect 21361 29597 21373 29631
rect 21407 29597 21419 29631
rect 21361 29591 21419 29597
rect 21545 29631 21603 29637
rect 21545 29597 21557 29631
rect 21591 29597 21603 29631
rect 21652 29628 21680 29668
rect 21818 29656 21824 29708
rect 21876 29656 21882 29708
rect 21928 29705 21956 29736
rect 22066 29736 22293 29764
rect 21913 29699 21971 29705
rect 21913 29665 21925 29699
rect 21959 29665 21971 29699
rect 21913 29659 21971 29665
rect 22066 29628 22094 29736
rect 22281 29733 22293 29736
rect 22327 29733 22339 29767
rect 22281 29727 22339 29733
rect 22462 29724 22468 29776
rect 22520 29724 22526 29776
rect 22557 29767 22615 29773
rect 22557 29733 22569 29767
rect 22603 29764 22615 29767
rect 22738 29764 22744 29776
rect 22603 29736 22744 29764
rect 22603 29733 22615 29736
rect 22557 29727 22615 29733
rect 22738 29724 22744 29736
rect 22796 29724 22802 29776
rect 23109 29767 23167 29773
rect 23109 29733 23121 29767
rect 23155 29764 23167 29767
rect 23937 29767 23995 29773
rect 23937 29764 23949 29767
rect 23155 29736 23949 29764
rect 23155 29733 23167 29736
rect 23109 29727 23167 29733
rect 23937 29733 23949 29736
rect 23983 29764 23995 29767
rect 25038 29764 25044 29776
rect 23983 29736 25044 29764
rect 23983 29733 23995 29736
rect 23937 29727 23995 29733
rect 25038 29724 25044 29736
rect 25096 29724 25102 29776
rect 22646 29656 22652 29708
rect 22704 29656 22710 29708
rect 22833 29699 22891 29705
rect 22833 29665 22845 29699
rect 22879 29696 22891 29699
rect 23474 29696 23480 29708
rect 22879 29668 23480 29696
rect 22879 29665 22891 29668
rect 22833 29659 22891 29665
rect 23474 29656 23480 29668
rect 23532 29696 23538 29708
rect 23569 29699 23627 29705
rect 23569 29696 23581 29699
rect 23532 29668 23581 29696
rect 23532 29656 23538 29668
rect 23569 29665 23581 29668
rect 23615 29665 23627 29699
rect 23569 29659 23627 29665
rect 24765 29699 24823 29705
rect 24765 29665 24777 29699
rect 24811 29696 24823 29699
rect 26421 29699 26479 29705
rect 26421 29696 26433 29699
rect 24811 29668 26433 29696
rect 24811 29665 24823 29668
rect 24765 29659 24823 29665
rect 26421 29665 26433 29668
rect 26467 29665 26479 29699
rect 26421 29659 26479 29665
rect 21652 29600 22094 29628
rect 21545 29591 21603 29597
rect 20165 29563 20223 29569
rect 20165 29560 20177 29563
rect 20128 29532 20177 29560
rect 20128 29520 20134 29532
rect 20165 29529 20177 29532
rect 20211 29529 20223 29563
rect 21560 29560 21588 29591
rect 24302 29588 24308 29640
rect 24360 29628 24366 29640
rect 24486 29628 24492 29640
rect 24360 29600 24492 29628
rect 24360 29588 24366 29600
rect 24486 29588 24492 29600
rect 24544 29628 24550 29640
rect 24673 29631 24731 29637
rect 24673 29628 24685 29631
rect 24544 29600 24685 29628
rect 24544 29588 24550 29600
rect 24673 29597 24685 29600
rect 24719 29597 24731 29631
rect 24673 29591 24731 29597
rect 26970 29588 26976 29640
rect 27028 29588 27034 29640
rect 21560 29532 22048 29560
rect 20165 29523 20223 29529
rect 22020 29504 22048 29532
rect 22554 29520 22560 29572
rect 22612 29560 22618 29572
rect 22612 29532 23244 29560
rect 22612 29520 22618 29532
rect 8386 29492 8392 29504
rect 8036 29464 8392 29492
rect 3881 29455 3939 29461
rect 8386 29452 8392 29464
rect 8444 29452 8450 29504
rect 12250 29452 12256 29504
rect 12308 29452 12314 29504
rect 13354 29452 13360 29504
rect 13412 29492 13418 29504
rect 14093 29495 14151 29501
rect 14093 29492 14105 29495
rect 13412 29464 14105 29492
rect 13412 29452 13418 29464
rect 14093 29461 14105 29464
rect 14139 29461 14151 29495
rect 14093 29455 14151 29461
rect 14737 29495 14795 29501
rect 14737 29461 14749 29495
rect 14783 29492 14795 29495
rect 15197 29495 15255 29501
rect 15197 29492 15209 29495
rect 14783 29464 15209 29492
rect 14783 29461 14795 29464
rect 14737 29455 14795 29461
rect 15197 29461 15209 29464
rect 15243 29461 15255 29495
rect 15197 29455 15255 29461
rect 15654 29452 15660 29504
rect 15712 29492 15718 29504
rect 16301 29495 16359 29501
rect 16301 29492 16313 29495
rect 15712 29464 16313 29492
rect 15712 29452 15718 29464
rect 16301 29461 16313 29464
rect 16347 29461 16359 29495
rect 16301 29455 16359 29461
rect 16942 29452 16948 29504
rect 17000 29452 17006 29504
rect 20254 29452 20260 29504
rect 20312 29452 20318 29504
rect 21450 29452 21456 29504
rect 21508 29492 21514 29504
rect 21729 29495 21787 29501
rect 21729 29492 21741 29495
rect 21508 29464 21741 29492
rect 21508 29452 21514 29464
rect 21729 29461 21741 29464
rect 21775 29461 21787 29495
rect 21729 29455 21787 29461
rect 22002 29452 22008 29504
rect 22060 29452 22066 29504
rect 22186 29452 22192 29504
rect 22244 29452 22250 29504
rect 22922 29452 22928 29504
rect 22980 29452 22986 29504
rect 23106 29452 23112 29504
rect 23164 29452 23170 29504
rect 23216 29492 23244 29532
rect 23382 29520 23388 29572
rect 23440 29560 23446 29572
rect 23477 29563 23535 29569
rect 23477 29560 23489 29563
rect 23440 29532 23489 29560
rect 23440 29520 23446 29532
rect 23477 29529 23489 29532
rect 23523 29529 23535 29563
rect 23477 29523 23535 29529
rect 25133 29563 25191 29569
rect 25133 29529 25145 29563
rect 25179 29560 25191 29563
rect 25406 29560 25412 29572
rect 25179 29532 25412 29560
rect 25179 29529 25191 29532
rect 25133 29523 25191 29529
rect 25406 29520 25412 29532
rect 25464 29520 25470 29572
rect 23566 29492 23572 29504
rect 23216 29464 23572 29492
rect 23566 29452 23572 29464
rect 23624 29452 23630 29504
rect 23750 29452 23756 29504
rect 23808 29492 23814 29504
rect 23937 29495 23995 29501
rect 23937 29492 23949 29495
rect 23808 29464 23949 29492
rect 23808 29452 23814 29464
rect 23937 29461 23949 29464
rect 23983 29461 23995 29495
rect 23937 29455 23995 29461
rect 552 29402 27416 29424
rect 552 29350 3756 29402
rect 3808 29350 3820 29402
rect 3872 29350 3884 29402
rect 3936 29350 3948 29402
rect 4000 29350 4012 29402
rect 4064 29350 10472 29402
rect 10524 29350 10536 29402
rect 10588 29350 10600 29402
rect 10652 29350 10664 29402
rect 10716 29350 10728 29402
rect 10780 29350 17188 29402
rect 17240 29350 17252 29402
rect 17304 29350 17316 29402
rect 17368 29350 17380 29402
rect 17432 29350 17444 29402
rect 17496 29350 23904 29402
rect 23956 29350 23968 29402
rect 24020 29350 24032 29402
rect 24084 29350 24096 29402
rect 24148 29350 24160 29402
rect 24212 29350 27416 29402
rect 552 29328 27416 29350
rect 5997 29291 6055 29297
rect 5997 29257 6009 29291
rect 6043 29288 6055 29291
rect 7006 29288 7012 29300
rect 6043 29260 7012 29288
rect 6043 29257 6055 29260
rect 5997 29251 6055 29257
rect 7006 29248 7012 29260
rect 7064 29248 7070 29300
rect 8570 29248 8576 29300
rect 8628 29248 8634 29300
rect 11422 29248 11428 29300
rect 11480 29248 11486 29300
rect 15654 29248 15660 29300
rect 15712 29248 15718 29300
rect 16301 29291 16359 29297
rect 16301 29257 16313 29291
rect 16347 29288 16359 29291
rect 16666 29288 16672 29300
rect 16347 29260 16672 29288
rect 16347 29257 16359 29260
rect 16301 29251 16359 29257
rect 16666 29248 16672 29260
rect 16724 29248 16730 29300
rect 18693 29291 18751 29297
rect 18693 29257 18705 29291
rect 18739 29288 18751 29291
rect 18874 29288 18880 29300
rect 18739 29260 18880 29288
rect 18739 29257 18751 29260
rect 18693 29251 18751 29257
rect 18874 29248 18880 29260
rect 18932 29248 18938 29300
rect 20346 29248 20352 29300
rect 20404 29248 20410 29300
rect 21450 29248 21456 29300
rect 21508 29248 21514 29300
rect 22557 29291 22615 29297
rect 22557 29257 22569 29291
rect 22603 29257 22615 29291
rect 22557 29251 22615 29257
rect 5718 29220 5724 29232
rect 5276 29192 5724 29220
rect 3510 29112 3516 29164
rect 3568 29112 3574 29164
rect 3602 29044 3608 29096
rect 3660 29084 3666 29096
rect 3769 29087 3827 29093
rect 3769 29084 3781 29087
rect 3660 29056 3781 29084
rect 3660 29044 3666 29056
rect 3769 29053 3781 29056
rect 3815 29053 3827 29087
rect 3769 29047 3827 29053
rect 5169 29087 5227 29093
rect 5169 29053 5181 29087
rect 5215 29084 5227 29087
rect 5276 29084 5304 29192
rect 5718 29180 5724 29192
rect 5776 29180 5782 29232
rect 5905 29223 5963 29229
rect 5905 29189 5917 29223
rect 5951 29220 5963 29223
rect 6362 29220 6368 29232
rect 5951 29192 6368 29220
rect 5951 29189 5963 29192
rect 5905 29183 5963 29189
rect 6362 29180 6368 29192
rect 6420 29180 6426 29232
rect 8389 29223 8447 29229
rect 8389 29189 8401 29223
rect 8435 29220 8447 29223
rect 8846 29220 8852 29232
rect 8435 29192 8852 29220
rect 8435 29189 8447 29192
rect 8389 29183 8447 29189
rect 8846 29180 8852 29192
rect 8904 29180 8910 29232
rect 8941 29223 8999 29229
rect 8941 29189 8953 29223
rect 8987 29220 8999 29223
rect 9033 29223 9091 29229
rect 9033 29220 9045 29223
rect 8987 29192 9045 29220
rect 8987 29189 8999 29192
rect 8941 29183 8999 29189
rect 9033 29189 9045 29192
rect 9079 29220 9091 29223
rect 10042 29220 10048 29232
rect 9079 29192 10048 29220
rect 9079 29189 9091 29192
rect 9033 29183 9091 29189
rect 10042 29180 10048 29192
rect 10100 29180 10106 29232
rect 12526 29180 12532 29232
rect 12584 29220 12590 29232
rect 17126 29220 17132 29232
rect 12584 29192 17132 29220
rect 12584 29180 12590 29192
rect 17126 29180 17132 29192
rect 17184 29220 17190 29232
rect 17184 29192 21496 29220
rect 17184 29180 17190 29192
rect 10318 29152 10324 29164
rect 5215 29056 5304 29084
rect 5368 29124 6224 29152
rect 5215 29053 5227 29056
rect 5169 29047 5227 29053
rect 5368 29028 5396 29124
rect 5445 29087 5503 29093
rect 5445 29053 5457 29087
rect 5491 29053 5503 29087
rect 5445 29047 5503 29053
rect 5537 29087 5595 29093
rect 5537 29053 5549 29087
rect 5583 29084 5595 29087
rect 5626 29084 5632 29096
rect 5583 29056 5632 29084
rect 5583 29053 5595 29056
rect 5537 29047 5595 29053
rect 5350 29016 5356 29028
rect 4908 28988 5356 29016
rect 4908 28957 4936 28988
rect 5350 28976 5356 28988
rect 5408 28976 5414 29028
rect 5460 29016 5488 29047
rect 5626 29044 5632 29056
rect 5684 29044 5690 29096
rect 5718 29044 5724 29096
rect 5776 29084 5782 29096
rect 6086 29084 6092 29096
rect 5776 29056 6092 29084
rect 5776 29044 5782 29056
rect 6086 29044 6092 29056
rect 6144 29044 6150 29096
rect 6196 29093 6224 29124
rect 10060 29124 10324 29152
rect 6181 29087 6239 29093
rect 6181 29053 6193 29087
rect 6227 29053 6239 29087
rect 6181 29047 6239 29053
rect 9033 29087 9091 29093
rect 9033 29053 9045 29087
rect 9079 29053 9091 29087
rect 9033 29047 9091 29053
rect 9217 29087 9275 29093
rect 9217 29053 9229 29087
rect 9263 29084 9275 29087
rect 9306 29084 9312 29096
rect 9263 29056 9312 29084
rect 9263 29053 9275 29056
rect 9217 29047 9275 29053
rect 6365 29019 6423 29025
rect 5460 28988 5580 29016
rect 5552 28960 5580 28988
rect 6365 28985 6377 29019
rect 6411 29016 6423 29019
rect 6638 29016 6644 29028
rect 6411 28988 6644 29016
rect 6411 28985 6423 28988
rect 6365 28979 6423 28985
rect 6638 28976 6644 28988
rect 6696 28976 6702 29028
rect 8294 28976 8300 29028
rect 8352 29016 8358 29028
rect 9048 29016 9076 29047
rect 9306 29044 9312 29056
rect 9364 29044 9370 29096
rect 9585 29087 9643 29093
rect 9585 29053 9597 29087
rect 9631 29084 9643 29087
rect 9950 29084 9956 29096
rect 9631 29056 9956 29084
rect 9631 29053 9643 29056
rect 9585 29047 9643 29053
rect 9950 29044 9956 29056
rect 10008 29044 10014 29096
rect 10060 29093 10088 29124
rect 10318 29112 10324 29124
rect 10376 29112 10382 29164
rect 12342 29152 12348 29164
rect 11624 29124 12348 29152
rect 10045 29087 10103 29093
rect 10045 29053 10057 29087
rect 10091 29053 10103 29087
rect 10045 29047 10103 29053
rect 10226 29044 10232 29096
rect 10284 29044 10290 29096
rect 11624 29093 11652 29124
rect 12342 29112 12348 29124
rect 12400 29152 12406 29164
rect 13630 29152 13636 29164
rect 12400 29124 13636 29152
rect 12400 29112 12406 29124
rect 13630 29112 13636 29124
rect 13688 29112 13694 29164
rect 14734 29112 14740 29164
rect 14792 29152 14798 29164
rect 18506 29152 18512 29164
rect 14792 29124 18512 29152
rect 14792 29112 14798 29124
rect 18506 29112 18512 29124
rect 18564 29112 18570 29164
rect 18966 29152 18972 29164
rect 18892 29124 18972 29152
rect 11609 29087 11667 29093
rect 11609 29053 11621 29087
rect 11655 29053 11667 29087
rect 11609 29047 11667 29053
rect 11698 29044 11704 29096
rect 11756 29044 11762 29096
rect 13173 29087 13231 29093
rect 13173 29053 13185 29087
rect 13219 29084 13231 29087
rect 13354 29084 13360 29096
rect 13219 29056 13360 29084
rect 13219 29053 13231 29056
rect 13173 29047 13231 29053
rect 13354 29044 13360 29056
rect 13412 29044 13418 29096
rect 15286 29044 15292 29096
rect 15344 29044 15350 29096
rect 15470 29044 15476 29096
rect 15528 29084 15534 29096
rect 16022 29084 16028 29096
rect 15528 29056 16028 29084
rect 15528 29044 15534 29056
rect 16022 29044 16028 29056
rect 16080 29044 16086 29096
rect 16574 29044 16580 29096
rect 16632 29044 16638 29096
rect 16758 29044 16764 29096
rect 16816 29044 16822 29096
rect 18892 29093 18920 29124
rect 18966 29112 18972 29124
rect 19024 29112 19030 29164
rect 20254 29152 20260 29164
rect 19260 29124 20260 29152
rect 16853 29087 16911 29093
rect 16853 29053 16865 29087
rect 16899 29053 16911 29087
rect 16853 29047 16911 29053
rect 18877 29087 18935 29093
rect 18877 29053 18889 29087
rect 18923 29053 18935 29087
rect 18877 29047 18935 29053
rect 19061 29087 19119 29093
rect 19061 29053 19073 29087
rect 19107 29084 19119 29087
rect 19150 29084 19156 29096
rect 19107 29056 19156 29084
rect 19107 29053 19119 29056
rect 19061 29047 19119 29053
rect 8352 28988 9076 29016
rect 8352 28976 8358 28988
rect 10962 28976 10968 29028
rect 11020 28976 11026 29028
rect 11146 28976 11152 29028
rect 11204 28976 11210 29028
rect 11425 29019 11483 29025
rect 11425 28985 11437 29019
rect 11471 29016 11483 29019
rect 12158 29016 12164 29028
rect 11471 28988 12164 29016
rect 11471 28985 11483 28988
rect 11425 28979 11483 28985
rect 12158 28976 12164 28988
rect 12216 28976 12222 29028
rect 12989 29019 13047 29025
rect 12989 28985 13001 29019
rect 13035 29016 13047 29019
rect 13078 29016 13084 29028
rect 13035 28988 13084 29016
rect 13035 28985 13047 28988
rect 12989 28979 13047 28985
rect 13078 28976 13084 28988
rect 13136 28976 13142 29028
rect 15838 28976 15844 29028
rect 15896 29016 15902 29028
rect 16117 29019 16175 29025
rect 16117 29016 16129 29019
rect 15896 28988 16129 29016
rect 15896 28976 15902 28988
rect 16117 28985 16129 28988
rect 16163 28985 16175 29019
rect 16117 28979 16175 28985
rect 16666 28976 16672 29028
rect 16724 28976 16730 29028
rect 16868 29016 16896 29047
rect 19150 29044 19156 29056
rect 19208 29044 19214 29096
rect 19260 29093 19288 29124
rect 20254 29112 20260 29124
rect 20312 29112 20318 29164
rect 20533 29155 20591 29161
rect 20533 29121 20545 29155
rect 20579 29152 20591 29155
rect 20898 29152 20904 29164
rect 20579 29124 20904 29152
rect 20579 29121 20591 29124
rect 20533 29115 20591 29121
rect 20898 29112 20904 29124
rect 20956 29112 20962 29164
rect 21358 29112 21364 29164
rect 21416 29112 21422 29164
rect 21468 29152 21496 29192
rect 21542 29180 21548 29232
rect 21600 29220 21606 29232
rect 21637 29223 21695 29229
rect 21637 29220 21649 29223
rect 21600 29192 21649 29220
rect 21600 29180 21606 29192
rect 21637 29189 21649 29192
rect 21683 29189 21695 29223
rect 22572 29220 22600 29251
rect 23106 29248 23112 29300
rect 23164 29248 23170 29300
rect 23566 29288 23572 29300
rect 23492 29260 23572 29288
rect 22738 29220 22744 29232
rect 22572 29192 22744 29220
rect 21637 29183 21695 29189
rect 22738 29180 22744 29192
rect 22796 29220 22802 29232
rect 23290 29220 23296 29232
rect 22796 29192 23296 29220
rect 22796 29180 22802 29192
rect 22554 29152 22560 29164
rect 21468 29124 22560 29152
rect 22554 29112 22560 29124
rect 22612 29112 22618 29164
rect 19245 29087 19303 29093
rect 19245 29053 19257 29087
rect 19291 29053 19303 29087
rect 19245 29047 19303 29053
rect 20070 29044 20076 29096
rect 20128 29044 20134 29096
rect 21266 29044 21272 29096
rect 21324 29044 21330 29096
rect 22462 29084 22468 29096
rect 22388 29056 22468 29084
rect 16776 28988 16896 29016
rect 18969 29019 19027 29025
rect 4893 28951 4951 28957
rect 4893 28917 4905 28951
rect 4939 28917 4951 28951
rect 4893 28911 4951 28917
rect 4982 28908 4988 28960
rect 5040 28908 5046 28960
rect 5534 28908 5540 28960
rect 5592 28908 5598 28960
rect 5626 28908 5632 28960
rect 5684 28948 5690 28960
rect 6089 28951 6147 28957
rect 6089 28948 6101 28951
rect 5684 28920 6101 28948
rect 5684 28908 5690 28920
rect 6089 28917 6101 28920
rect 6135 28917 6147 28951
rect 6089 28911 6147 28917
rect 8570 28908 8576 28960
rect 8628 28948 8634 28960
rect 8754 28948 8760 28960
rect 8628 28920 8760 28948
rect 8628 28908 8634 28920
rect 8754 28908 8760 28920
rect 8812 28908 8818 28960
rect 9398 28908 9404 28960
rect 9456 28908 9462 28960
rect 10134 28908 10140 28960
rect 10192 28908 10198 28960
rect 11330 28908 11336 28960
rect 11388 28908 11394 28960
rect 13262 28908 13268 28960
rect 13320 28948 13326 28960
rect 13357 28951 13415 28957
rect 13357 28948 13369 28951
rect 13320 28920 13369 28948
rect 13320 28908 13326 28920
rect 13357 28917 13369 28920
rect 13403 28917 13415 28951
rect 13357 28911 13415 28917
rect 16298 28908 16304 28960
rect 16356 28957 16362 28960
rect 16356 28951 16375 28957
rect 16363 28917 16375 28951
rect 16356 28911 16375 28917
rect 16485 28951 16543 28957
rect 16485 28917 16497 28951
rect 16531 28948 16543 28951
rect 16776 28948 16804 28988
rect 18969 28985 18981 29019
rect 19015 29016 19027 29019
rect 19426 29016 19432 29028
rect 19015 28988 19432 29016
rect 19015 28985 19027 28988
rect 18969 28979 19027 28985
rect 19426 28976 19432 28988
rect 19484 28976 19490 29028
rect 20346 28976 20352 29028
rect 20404 29016 20410 29028
rect 22388 29025 22416 29056
rect 22462 29044 22468 29056
rect 22520 29084 22526 29096
rect 22922 29084 22928 29096
rect 22520 29056 22928 29084
rect 22520 29044 22526 29056
rect 22922 29044 22928 29056
rect 22980 29044 22986 29096
rect 23017 29087 23075 29093
rect 23017 29053 23029 29087
rect 23063 29084 23075 29087
rect 23124 29084 23152 29192
rect 23290 29180 23296 29192
rect 23348 29180 23354 29232
rect 23063 29056 23152 29084
rect 23063 29053 23075 29056
rect 23017 29047 23075 29053
rect 23198 29044 23204 29096
rect 23256 29084 23262 29096
rect 23293 29087 23351 29093
rect 23293 29084 23305 29087
rect 23256 29056 23305 29084
rect 23256 29044 23262 29056
rect 23293 29053 23305 29056
rect 23339 29053 23351 29087
rect 23293 29047 23351 29053
rect 23492 29025 23520 29260
rect 23566 29248 23572 29260
rect 23624 29288 23630 29300
rect 26881 29291 26939 29297
rect 26881 29288 26893 29291
rect 23624 29260 26893 29288
rect 23624 29248 23630 29260
rect 26881 29257 26893 29260
rect 26927 29288 26939 29291
rect 26970 29288 26976 29300
rect 26927 29260 26976 29288
rect 26927 29257 26939 29260
rect 26881 29251 26939 29257
rect 26970 29248 26976 29260
rect 27028 29248 27034 29300
rect 24026 29112 24032 29164
rect 24084 29112 24090 29164
rect 23569 29087 23627 29093
rect 23569 29053 23581 29087
rect 23615 29084 23627 29087
rect 24118 29084 24124 29096
rect 23615 29056 24124 29084
rect 23615 29053 23627 29056
rect 23569 29047 23627 29053
rect 24118 29044 24124 29056
rect 24176 29044 24182 29096
rect 25498 29044 25504 29096
rect 25556 29084 25562 29096
rect 26142 29084 26148 29096
rect 25556 29056 26148 29084
rect 25556 29044 25562 29056
rect 26142 29044 26148 29056
rect 26200 29044 26206 29096
rect 24302 29025 24308 29028
rect 22373 29019 22431 29025
rect 22373 29016 22385 29019
rect 20404 28988 22385 29016
rect 20404 28976 20410 28988
rect 22373 28985 22385 28988
rect 22419 28985 22431 29019
rect 23477 29019 23535 29025
rect 22373 28979 22431 28985
rect 22756 28988 23428 29016
rect 16531 28920 16804 28948
rect 16531 28917 16543 28920
rect 16485 28911 16543 28917
rect 16356 28908 16362 28911
rect 17034 28908 17040 28960
rect 17092 28908 17098 28960
rect 22554 28908 22560 28960
rect 22612 28957 22618 28960
rect 22756 28957 22784 28988
rect 23400 28960 23428 28988
rect 23477 28985 23489 29019
rect 23523 28985 23535 29019
rect 23477 28979 23535 28985
rect 24296 28979 24308 29025
rect 24302 28976 24308 28979
rect 24360 28976 24366 29028
rect 24394 28976 24400 29028
rect 24452 29016 24458 29028
rect 24452 28988 25452 29016
rect 24452 28976 24458 28988
rect 22612 28951 22631 28957
rect 22619 28917 22631 28951
rect 22612 28911 22631 28917
rect 22741 28951 22799 28957
rect 22741 28917 22753 28951
rect 22787 28917 22799 28951
rect 22741 28911 22799 28917
rect 22612 28908 22618 28911
rect 22922 28908 22928 28960
rect 22980 28908 22986 28960
rect 23382 28908 23388 28960
rect 23440 28908 23446 28960
rect 25424 28957 25452 28988
rect 25590 28976 25596 29028
rect 25648 29016 25654 29028
rect 25746 29019 25804 29025
rect 25746 29016 25758 29019
rect 25648 28988 25758 29016
rect 25648 28976 25654 28988
rect 25746 28985 25758 28988
rect 25792 28985 25804 29019
rect 25746 28979 25804 28985
rect 25409 28951 25467 28957
rect 25409 28917 25421 28951
rect 25455 28917 25467 28951
rect 25409 28911 25467 28917
rect 552 28858 27576 28880
rect 552 28806 7114 28858
rect 7166 28806 7178 28858
rect 7230 28806 7242 28858
rect 7294 28806 7306 28858
rect 7358 28806 7370 28858
rect 7422 28806 13830 28858
rect 13882 28806 13894 28858
rect 13946 28806 13958 28858
rect 14010 28806 14022 28858
rect 14074 28806 14086 28858
rect 14138 28806 20546 28858
rect 20598 28806 20610 28858
rect 20662 28806 20674 28858
rect 20726 28806 20738 28858
rect 20790 28806 20802 28858
rect 20854 28806 27262 28858
rect 27314 28806 27326 28858
rect 27378 28806 27390 28858
rect 27442 28806 27454 28858
rect 27506 28806 27518 28858
rect 27570 28806 27576 28858
rect 552 28784 27576 28806
rect 3050 28704 3056 28756
rect 3108 28744 3114 28756
rect 3326 28744 3332 28756
rect 3108 28716 3332 28744
rect 3108 28704 3114 28716
rect 3326 28704 3332 28716
rect 3384 28744 3390 28756
rect 3384 28716 4016 28744
rect 3384 28704 3390 28716
rect 3510 28636 3516 28688
rect 3568 28676 3574 28688
rect 3988 28676 4016 28716
rect 4154 28704 4160 28756
rect 4212 28744 4218 28756
rect 4433 28747 4491 28753
rect 4433 28744 4445 28747
rect 4212 28716 4445 28744
rect 4212 28704 4218 28716
rect 4433 28713 4445 28716
rect 4479 28713 4491 28747
rect 4433 28707 4491 28713
rect 4601 28747 4659 28753
rect 4601 28713 4613 28747
rect 4647 28744 4659 28747
rect 4982 28744 4988 28756
rect 4647 28716 4988 28744
rect 4647 28713 4659 28716
rect 4601 28707 4659 28713
rect 4982 28704 4988 28716
rect 5040 28704 5046 28756
rect 5810 28704 5816 28756
rect 5868 28704 5874 28756
rect 6822 28704 6828 28756
rect 6880 28744 6886 28756
rect 6880 28716 8708 28744
rect 6880 28704 6886 28716
rect 8110 28685 8116 28688
rect 4801 28679 4859 28685
rect 4801 28676 4813 28679
rect 3568 28648 3924 28676
rect 3988 28648 4813 28676
rect 3568 28636 3574 28648
rect 3602 28568 3608 28620
rect 3660 28617 3666 28620
rect 3896 28617 3924 28648
rect 4801 28645 4813 28648
rect 4847 28645 4859 28679
rect 4801 28639 4859 28645
rect 8097 28679 8116 28685
rect 8097 28645 8109 28679
rect 8097 28639 8116 28645
rect 8110 28636 8116 28639
rect 8168 28636 8174 28688
rect 8297 28679 8355 28685
rect 8297 28645 8309 28679
rect 8343 28676 8355 28679
rect 8570 28676 8576 28688
rect 8343 28648 8576 28676
rect 8343 28645 8355 28648
rect 8297 28639 8355 28645
rect 8570 28636 8576 28648
rect 8628 28636 8634 28688
rect 3660 28571 3672 28617
rect 3881 28611 3939 28617
rect 3881 28577 3893 28611
rect 3927 28577 3939 28611
rect 3881 28571 3939 28577
rect 3660 28568 3666 28571
rect 5350 28568 5356 28620
rect 5408 28608 5414 28620
rect 6730 28617 6736 28620
rect 6181 28611 6239 28617
rect 6181 28608 6193 28611
rect 5408 28580 6193 28608
rect 5408 28568 5414 28580
rect 6181 28577 6193 28580
rect 6227 28577 6239 28611
rect 6181 28571 6239 28577
rect 6724 28571 6736 28617
rect 6730 28568 6736 28571
rect 6788 28568 6794 28620
rect 7834 28568 7840 28620
rect 7892 28608 7898 28620
rect 8680 28617 8708 28716
rect 10318 28704 10324 28756
rect 10376 28744 10382 28756
rect 13265 28747 13323 28753
rect 13265 28744 13277 28747
rect 10376 28716 10548 28744
rect 10376 28704 10382 28716
rect 9208 28679 9266 28685
rect 9208 28645 9220 28679
rect 9254 28676 9266 28679
rect 9398 28676 9404 28688
rect 9254 28648 9404 28676
rect 9254 28645 9266 28648
rect 9208 28639 9266 28645
rect 9398 28636 9404 28648
rect 9456 28636 9462 28688
rect 10520 28676 10548 28716
rect 12406 28716 13277 28744
rect 10520 28648 10652 28676
rect 8389 28611 8447 28617
rect 8389 28608 8401 28611
rect 7892 28580 8401 28608
rect 7892 28568 7898 28580
rect 8389 28577 8401 28580
rect 8435 28577 8447 28611
rect 8389 28571 8447 28577
rect 8481 28611 8539 28617
rect 8481 28577 8493 28611
rect 8527 28577 8539 28611
rect 8481 28571 8539 28577
rect 8665 28611 8723 28617
rect 8665 28577 8677 28611
rect 8711 28608 8723 28611
rect 9766 28608 9772 28620
rect 8711 28580 9772 28608
rect 8711 28577 8723 28580
rect 8665 28571 8723 28577
rect 6273 28543 6331 28549
rect 6273 28509 6285 28543
rect 6319 28509 6331 28543
rect 6273 28503 6331 28509
rect 2501 28407 2559 28413
rect 2501 28373 2513 28407
rect 2547 28404 2559 28407
rect 2866 28404 2872 28416
rect 2547 28376 2872 28404
rect 2547 28373 2559 28376
rect 2501 28367 2559 28373
rect 2866 28364 2872 28376
rect 2924 28364 2930 28416
rect 4617 28407 4675 28413
rect 4617 28373 4629 28407
rect 4663 28404 4675 28407
rect 5626 28404 5632 28416
rect 4663 28376 5632 28404
rect 4663 28373 4675 28376
rect 4617 28367 4675 28373
rect 5626 28364 5632 28376
rect 5684 28364 5690 28416
rect 6288 28404 6316 28503
rect 6454 28500 6460 28552
rect 6512 28500 6518 28552
rect 8018 28500 8024 28552
rect 8076 28540 8082 28552
rect 8496 28540 8524 28571
rect 9766 28568 9772 28580
rect 9824 28568 9830 28620
rect 10624 28617 10652 28648
rect 11514 28636 11520 28688
rect 11572 28676 11578 28688
rect 11609 28679 11667 28685
rect 11609 28676 11621 28679
rect 11572 28648 11621 28676
rect 11572 28636 11578 28648
rect 11609 28645 11621 28648
rect 11655 28676 11667 28679
rect 12406 28676 12434 28716
rect 13265 28713 13277 28716
rect 13311 28713 13323 28747
rect 13265 28707 13323 28713
rect 13449 28747 13507 28753
rect 13449 28713 13461 28747
rect 13495 28744 13507 28747
rect 13722 28744 13728 28756
rect 13495 28716 13728 28744
rect 13495 28713 13507 28716
rect 13449 28707 13507 28713
rect 11655 28648 12434 28676
rect 13280 28676 13308 28707
rect 13722 28704 13728 28716
rect 13780 28704 13786 28756
rect 14200 28716 15148 28744
rect 14200 28685 14228 28716
rect 14185 28679 14243 28685
rect 14185 28676 14197 28679
rect 13280 28648 14197 28676
rect 11655 28645 11667 28648
rect 11609 28639 11667 28645
rect 14185 28645 14197 28648
rect 14231 28645 14243 28679
rect 14185 28639 14243 28645
rect 15013 28679 15071 28685
rect 15013 28645 15025 28679
rect 15059 28645 15071 28679
rect 15120 28676 15148 28716
rect 15194 28704 15200 28756
rect 15252 28753 15258 28756
rect 15252 28747 15271 28753
rect 15259 28713 15271 28747
rect 15252 28707 15271 28713
rect 15381 28747 15439 28753
rect 15381 28713 15393 28747
rect 15427 28744 15439 28747
rect 15427 28716 16160 28744
rect 15427 28713 15439 28716
rect 15381 28707 15439 28713
rect 15252 28704 15258 28707
rect 15838 28676 15844 28688
rect 15120 28648 15844 28676
rect 15013 28639 15071 28645
rect 10401 28611 10459 28617
rect 10401 28577 10413 28611
rect 10447 28577 10459 28611
rect 10401 28571 10459 28577
rect 10597 28611 10655 28617
rect 10597 28577 10609 28611
rect 10643 28577 10655 28611
rect 10597 28571 10655 28577
rect 10965 28611 11023 28617
rect 10965 28577 10977 28611
rect 11011 28577 11023 28611
rect 10965 28571 11023 28577
rect 12897 28611 12955 28617
rect 12897 28577 12909 28611
rect 12943 28608 12955 28611
rect 12986 28608 12992 28620
rect 12943 28580 12992 28608
rect 12943 28577 12955 28580
rect 12897 28571 12955 28577
rect 8076 28512 8524 28540
rect 8941 28543 8999 28549
rect 8076 28500 8082 28512
rect 8941 28509 8953 28543
rect 8987 28509 8999 28543
rect 8941 28503 8999 28509
rect 7466 28432 7472 28484
rect 7524 28472 7530 28484
rect 7929 28475 7987 28481
rect 7929 28472 7941 28475
rect 7524 28444 7941 28472
rect 7524 28432 7530 28444
rect 7929 28441 7941 28444
rect 7975 28441 7987 28475
rect 7929 28435 7987 28441
rect 8294 28432 8300 28484
rect 8352 28472 8358 28484
rect 8389 28475 8447 28481
rect 8389 28472 8401 28475
rect 8352 28444 8401 28472
rect 8352 28432 8358 28444
rect 8389 28441 8401 28444
rect 8435 28441 8447 28475
rect 8389 28435 8447 28441
rect 8478 28432 8484 28484
rect 8536 28472 8542 28484
rect 8956 28472 8984 28503
rect 10226 28500 10232 28552
rect 10284 28540 10290 28552
rect 10419 28540 10447 28571
rect 10980 28540 11008 28571
rect 12986 28568 12992 28580
rect 13044 28608 13050 28620
rect 14461 28611 14519 28617
rect 14461 28608 14473 28611
rect 13044 28580 14473 28608
rect 13044 28568 13050 28580
rect 14461 28577 14473 28580
rect 14507 28577 14519 28611
rect 14461 28571 14519 28577
rect 14642 28568 14648 28620
rect 14700 28568 14706 28620
rect 15028 28608 15056 28639
rect 15838 28636 15844 28648
rect 15896 28636 15902 28688
rect 16132 28685 16160 28716
rect 16298 28704 16304 28756
rect 16356 28744 16362 28756
rect 16485 28747 16543 28753
rect 16485 28744 16497 28747
rect 16356 28716 16497 28744
rect 16356 28704 16362 28716
rect 16485 28713 16497 28716
rect 16531 28713 16543 28747
rect 16485 28707 16543 28713
rect 23750 28704 23756 28756
rect 23808 28704 23814 28756
rect 24213 28747 24271 28753
rect 24213 28713 24225 28747
rect 24259 28744 24271 28747
rect 24302 28744 24308 28756
rect 24259 28716 24308 28744
rect 24259 28713 24271 28716
rect 24213 28707 24271 28713
rect 24302 28704 24308 28716
rect 24360 28704 24366 28756
rect 25590 28704 25596 28756
rect 25648 28704 25654 28756
rect 16117 28679 16175 28685
rect 16117 28645 16129 28679
rect 16163 28676 16175 28679
rect 16574 28676 16580 28688
rect 16163 28648 16580 28676
rect 16163 28645 16175 28648
rect 16117 28639 16175 28645
rect 16574 28636 16580 28648
rect 16632 28636 16638 28688
rect 22189 28679 22247 28685
rect 16868 28648 18736 28676
rect 15470 28608 15476 28620
rect 15028 28580 15476 28608
rect 15470 28568 15476 28580
rect 15528 28568 15534 28620
rect 15565 28611 15623 28617
rect 15565 28577 15577 28611
rect 15611 28608 15623 28611
rect 15746 28608 15752 28620
rect 15611 28580 15752 28608
rect 15611 28577 15623 28580
rect 15565 28571 15623 28577
rect 10284 28512 10447 28540
rect 10520 28512 11008 28540
rect 13817 28543 13875 28549
rect 10284 28500 10290 28512
rect 8536 28444 8984 28472
rect 8536 28432 8542 28444
rect 10318 28432 10324 28484
rect 10376 28472 10382 28484
rect 10520 28472 10548 28512
rect 13817 28509 13829 28543
rect 13863 28540 13875 28543
rect 13906 28540 13912 28552
rect 13863 28512 13912 28540
rect 13863 28509 13875 28512
rect 13817 28503 13875 28509
rect 13906 28500 13912 28512
rect 13964 28540 13970 28552
rect 15194 28540 15200 28552
rect 13964 28512 15200 28540
rect 13964 28500 13970 28512
rect 15194 28500 15200 28512
rect 15252 28500 15258 28552
rect 15378 28500 15384 28552
rect 15436 28540 15442 28552
rect 15580 28540 15608 28571
rect 15746 28568 15752 28580
rect 15804 28568 15810 28620
rect 15436 28512 15608 28540
rect 15436 28500 15442 28512
rect 10376 28444 10548 28472
rect 10597 28475 10655 28481
rect 10376 28432 10382 28444
rect 10597 28441 10609 28475
rect 10643 28472 10655 28475
rect 10962 28472 10968 28484
rect 10643 28444 10968 28472
rect 10643 28441 10655 28444
rect 10597 28435 10655 28441
rect 10962 28432 10968 28444
rect 11020 28432 11026 28484
rect 11238 28432 11244 28484
rect 11296 28432 11302 28484
rect 14829 28475 14887 28481
rect 14829 28472 14841 28475
rect 14200 28444 14841 28472
rect 6638 28404 6644 28416
rect 6288 28376 6644 28404
rect 6638 28364 6644 28376
rect 6696 28364 6702 28416
rect 7834 28364 7840 28416
rect 7892 28364 7898 28416
rect 8113 28407 8171 28413
rect 8113 28373 8125 28407
rect 8159 28404 8171 28407
rect 8312 28404 8340 28432
rect 8159 28376 8340 28404
rect 8159 28373 8171 28376
rect 8113 28367 8171 28373
rect 10226 28364 10232 28416
rect 10284 28404 10290 28416
rect 11054 28404 11060 28416
rect 10284 28376 11060 28404
rect 10284 28364 10290 28376
rect 11054 28364 11060 28376
rect 11112 28364 11118 28416
rect 11330 28364 11336 28416
rect 11388 28404 11394 28416
rect 11609 28407 11667 28413
rect 11609 28404 11621 28407
rect 11388 28376 11621 28404
rect 11388 28364 11394 28376
rect 11609 28373 11621 28376
rect 11655 28373 11667 28407
rect 11609 28367 11667 28373
rect 11790 28364 11796 28416
rect 11848 28364 11854 28416
rect 13262 28364 13268 28416
rect 13320 28364 13326 28416
rect 14200 28413 14228 28444
rect 14829 28441 14841 28444
rect 14875 28441 14887 28475
rect 14829 28435 14887 28441
rect 15749 28475 15807 28481
rect 15749 28441 15761 28475
rect 15795 28472 15807 28475
rect 15856 28472 15884 28636
rect 16868 28620 16896 28648
rect 16301 28611 16359 28617
rect 16301 28577 16313 28611
rect 16347 28577 16359 28611
rect 16301 28571 16359 28577
rect 16761 28611 16819 28617
rect 16761 28577 16773 28611
rect 16807 28608 16819 28611
rect 16850 28608 16856 28620
rect 16807 28580 16856 28608
rect 16807 28577 16819 28580
rect 16761 28571 16819 28577
rect 15795 28444 15884 28472
rect 15795 28441 15807 28444
rect 15749 28435 15807 28441
rect 14185 28407 14243 28413
rect 14185 28373 14197 28407
rect 14231 28373 14243 28407
rect 14185 28367 14243 28373
rect 14274 28364 14280 28416
rect 14332 28404 14338 28416
rect 14369 28407 14427 28413
rect 14369 28404 14381 28407
rect 14332 28376 14381 28404
rect 14332 28364 14338 28376
rect 14369 28373 14381 28376
rect 14415 28373 14427 28407
rect 14369 28367 14427 28373
rect 15102 28364 15108 28416
rect 15160 28404 15166 28416
rect 15197 28407 15255 28413
rect 15197 28404 15209 28407
rect 15160 28376 15209 28404
rect 15160 28364 15166 28376
rect 15197 28373 15209 28376
rect 15243 28373 15255 28407
rect 16316 28404 16344 28571
rect 16850 28568 16856 28580
rect 16908 28568 16914 28620
rect 17034 28617 17040 28620
rect 17028 28608 17040 28617
rect 16995 28580 17040 28608
rect 17028 28571 17040 28580
rect 17034 28568 17040 28571
rect 17092 28568 17098 28620
rect 17586 28568 17592 28620
rect 17644 28608 17650 28620
rect 18325 28611 18383 28617
rect 18325 28608 18337 28611
rect 17644 28580 18337 28608
rect 17644 28568 17650 28580
rect 18325 28577 18337 28580
rect 18371 28577 18383 28611
rect 18325 28571 18383 28577
rect 18414 28568 18420 28620
rect 18472 28568 18478 28620
rect 18708 28617 18736 28648
rect 22189 28645 22201 28679
rect 22235 28676 22247 28679
rect 24854 28676 24860 28688
rect 22235 28648 24860 28676
rect 22235 28645 22247 28648
rect 22189 28639 22247 28645
rect 24854 28636 24860 28648
rect 24912 28636 24918 28688
rect 18693 28611 18751 28617
rect 18693 28577 18705 28611
rect 18739 28577 18751 28611
rect 18693 28571 18751 28577
rect 18782 28568 18788 28620
rect 18840 28608 18846 28620
rect 18949 28611 19007 28617
rect 18949 28608 18961 28611
rect 18840 28580 18961 28608
rect 18840 28568 18846 28580
rect 18949 28577 18961 28580
rect 18995 28577 19007 28611
rect 18949 28571 19007 28577
rect 19334 28568 19340 28620
rect 19392 28608 19398 28620
rect 21361 28611 21419 28617
rect 21361 28608 21373 28611
rect 19392 28580 21373 28608
rect 19392 28568 19398 28580
rect 21361 28577 21373 28580
rect 21407 28608 21419 28611
rect 22278 28608 22284 28620
rect 21407 28580 22284 28608
rect 21407 28577 21419 28580
rect 21361 28571 21419 28577
rect 22278 28568 22284 28580
rect 22336 28568 22342 28620
rect 22465 28611 22523 28617
rect 22465 28577 22477 28611
rect 22511 28577 22523 28611
rect 22465 28571 22523 28577
rect 22649 28611 22707 28617
rect 22649 28577 22661 28611
rect 22695 28608 22707 28611
rect 22922 28608 22928 28620
rect 22695 28580 22928 28608
rect 22695 28577 22707 28580
rect 22649 28571 22707 28577
rect 19702 28500 19708 28552
rect 19760 28540 19766 28552
rect 20165 28543 20223 28549
rect 20165 28540 20177 28543
rect 19760 28512 20177 28540
rect 19760 28500 19766 28512
rect 20165 28509 20177 28512
rect 20211 28509 20223 28543
rect 20165 28503 20223 28509
rect 20717 28543 20775 28549
rect 20717 28509 20729 28543
rect 20763 28540 20775 28543
rect 21634 28540 21640 28552
rect 20763 28512 21640 28540
rect 20763 28509 20775 28512
rect 20717 28503 20775 28509
rect 20073 28475 20131 28481
rect 20073 28441 20085 28475
rect 20119 28472 20131 28475
rect 20732 28472 20760 28503
rect 21634 28500 21640 28512
rect 21692 28540 21698 28552
rect 22480 28540 22508 28571
rect 22922 28568 22928 28580
rect 22980 28568 22986 28620
rect 23382 28568 23388 28620
rect 23440 28568 23446 28620
rect 23569 28611 23627 28617
rect 23569 28577 23581 28611
rect 23615 28608 23627 28611
rect 23658 28608 23664 28620
rect 23615 28580 23664 28608
rect 23615 28577 23627 28580
rect 23569 28571 23627 28577
rect 23658 28568 23664 28580
rect 23716 28568 23722 28620
rect 24029 28611 24087 28617
rect 24029 28577 24041 28611
rect 24075 28608 24087 28611
rect 24302 28608 24308 28620
rect 24075 28580 24308 28608
rect 24075 28577 24087 28580
rect 24029 28571 24087 28577
rect 24302 28568 24308 28580
rect 24360 28568 24366 28620
rect 25406 28568 25412 28620
rect 25464 28568 25470 28620
rect 25593 28611 25651 28617
rect 25593 28577 25605 28611
rect 25639 28577 25651 28611
rect 25593 28571 25651 28577
rect 21692 28512 22508 28540
rect 21692 28500 21698 28512
rect 25038 28500 25044 28552
rect 25096 28540 25102 28552
rect 25608 28540 25636 28571
rect 25096 28512 25636 28540
rect 25096 28500 25102 28512
rect 22370 28472 22376 28484
rect 20119 28444 20760 28472
rect 22066 28444 22376 28472
rect 20119 28441 20131 28444
rect 20073 28435 20131 28441
rect 16758 28404 16764 28416
rect 16316 28376 16764 28404
rect 15197 28367 15255 28373
rect 16758 28364 16764 28376
rect 16816 28404 16822 28416
rect 17862 28404 17868 28416
rect 16816 28376 17868 28404
rect 16816 28364 16822 28376
rect 17862 28364 17868 28376
rect 17920 28404 17926 28416
rect 18141 28407 18199 28413
rect 18141 28404 18153 28407
rect 17920 28376 18153 28404
rect 17920 28364 17926 28376
rect 18141 28373 18153 28376
rect 18187 28373 18199 28407
rect 18141 28367 18199 28373
rect 18966 28364 18972 28416
rect 19024 28404 19030 28416
rect 22066 28404 22094 28444
rect 22370 28432 22376 28444
rect 22428 28432 22434 28484
rect 19024 28376 22094 28404
rect 19024 28364 19030 28376
rect 22278 28364 22284 28416
rect 22336 28364 22342 28416
rect 552 28314 27416 28336
rect 552 28262 3756 28314
rect 3808 28262 3820 28314
rect 3872 28262 3884 28314
rect 3936 28262 3948 28314
rect 4000 28262 4012 28314
rect 4064 28262 10472 28314
rect 10524 28262 10536 28314
rect 10588 28262 10600 28314
rect 10652 28262 10664 28314
rect 10716 28262 10728 28314
rect 10780 28262 17188 28314
rect 17240 28262 17252 28314
rect 17304 28262 17316 28314
rect 17368 28262 17380 28314
rect 17432 28262 17444 28314
rect 17496 28262 23904 28314
rect 23956 28262 23968 28314
rect 24020 28262 24032 28314
rect 24084 28262 24096 28314
rect 24148 28262 24160 28314
rect 24212 28262 27416 28314
rect 552 28240 27416 28262
rect 3421 28203 3479 28209
rect 3421 28169 3433 28203
rect 3467 28200 3479 28203
rect 3602 28200 3608 28212
rect 3467 28172 3608 28200
rect 3467 28169 3479 28172
rect 3421 28163 3479 28169
rect 3602 28160 3608 28172
rect 3660 28160 3666 28212
rect 6086 28160 6092 28212
rect 6144 28160 6150 28212
rect 6730 28160 6736 28212
rect 6788 28200 6794 28212
rect 6917 28203 6975 28209
rect 6917 28200 6929 28203
rect 6788 28172 6929 28200
rect 6788 28160 6794 28172
rect 6917 28169 6929 28172
rect 6963 28169 6975 28203
rect 6917 28163 6975 28169
rect 8110 28160 8116 28212
rect 8168 28160 8174 28212
rect 9950 28160 9956 28212
rect 10008 28160 10014 28212
rect 10134 28160 10140 28212
rect 10192 28160 10198 28212
rect 12986 28160 12992 28212
rect 13044 28160 13050 28212
rect 13354 28160 13360 28212
rect 13412 28200 13418 28212
rect 13725 28203 13783 28209
rect 13725 28200 13737 28203
rect 13412 28172 13737 28200
rect 13412 28160 13418 28172
rect 13725 28169 13737 28172
rect 13771 28169 13783 28203
rect 13725 28163 13783 28169
rect 13906 28160 13912 28212
rect 13964 28160 13970 28212
rect 14001 28203 14059 28209
rect 14001 28169 14013 28203
rect 14047 28200 14059 28203
rect 14642 28200 14648 28212
rect 14047 28172 14648 28200
rect 14047 28169 14059 28172
rect 14001 28163 14059 28169
rect 10505 28135 10563 28141
rect 10505 28101 10517 28135
rect 10551 28132 10563 28135
rect 10962 28132 10968 28144
rect 10551 28104 10968 28132
rect 10551 28101 10563 28104
rect 10505 28095 10563 28101
rect 10962 28092 10968 28104
rect 11020 28092 11026 28144
rect 11146 28092 11152 28144
rect 11204 28092 11210 28144
rect 10318 28024 10324 28076
rect 10376 28064 10382 28076
rect 10376 28036 11008 28064
rect 10376 28024 10382 28036
rect 3234 27956 3240 28008
rect 3292 27956 3298 28008
rect 4065 27999 4123 28005
rect 4065 27965 4077 27999
rect 4111 27996 4123 27999
rect 4154 27996 4160 28008
rect 4111 27968 4160 27996
rect 4111 27965 4123 27968
rect 4065 27959 4123 27965
rect 4154 27956 4160 27968
rect 4212 27956 4218 28008
rect 5350 27956 5356 28008
rect 5408 27996 5414 28008
rect 5537 27999 5595 28005
rect 5537 27996 5549 27999
rect 5408 27968 5549 27996
rect 5408 27956 5414 27968
rect 5537 27965 5549 27968
rect 5583 27965 5595 27999
rect 5537 27959 5595 27965
rect 5718 27956 5724 28008
rect 5776 27996 5782 28008
rect 5813 27999 5871 28005
rect 5813 27996 5825 27999
rect 5776 27968 5825 27996
rect 5776 27956 5782 27968
rect 5813 27965 5825 27968
rect 5859 27965 5871 27999
rect 5813 27959 5871 27965
rect 6457 27999 6515 28005
rect 6457 27965 6469 27999
rect 6503 27996 6515 27999
rect 6822 27996 6828 28008
rect 6503 27968 6828 27996
rect 6503 27965 6515 27968
rect 6457 27959 6515 27965
rect 6822 27956 6828 27968
rect 6880 27956 6886 28008
rect 7101 27999 7159 28005
rect 7101 27965 7113 27999
rect 7147 27996 7159 27999
rect 7466 27996 7472 28008
rect 7147 27968 7472 27996
rect 7147 27965 7159 27968
rect 7101 27959 7159 27965
rect 7466 27956 7472 27968
rect 7524 27956 7530 28008
rect 7653 27999 7711 28005
rect 7653 27965 7665 27999
rect 7699 27965 7711 27999
rect 7653 27959 7711 27965
rect 2777 27931 2835 27937
rect 2777 27897 2789 27931
rect 2823 27897 2835 27931
rect 2777 27891 2835 27897
rect 2961 27931 3019 27937
rect 2961 27897 2973 27931
rect 3007 27928 3019 27931
rect 3142 27928 3148 27940
rect 3007 27900 3148 27928
rect 3007 27897 3019 27900
rect 2961 27891 3019 27897
rect 2593 27863 2651 27869
rect 2593 27829 2605 27863
rect 2639 27860 2651 27863
rect 2682 27860 2688 27872
rect 2639 27832 2688 27860
rect 2639 27829 2651 27832
rect 2593 27823 2651 27829
rect 2682 27820 2688 27832
rect 2740 27820 2746 27872
rect 2792 27860 2820 27891
rect 3142 27888 3148 27900
rect 3200 27888 3206 27940
rect 5629 27931 5687 27937
rect 5629 27897 5641 27931
rect 5675 27928 5687 27931
rect 6178 27928 6184 27940
rect 5675 27900 6184 27928
rect 5675 27897 5687 27900
rect 5629 27891 5687 27897
rect 6178 27888 6184 27900
rect 6236 27888 6242 27940
rect 6638 27888 6644 27940
rect 6696 27928 6702 27940
rect 7668 27928 7696 27959
rect 7834 27956 7840 28008
rect 7892 27996 7898 28008
rect 7929 27999 7987 28005
rect 7929 27996 7941 27999
rect 7892 27968 7941 27996
rect 7892 27956 7898 27968
rect 7929 27965 7941 27968
rect 7975 27996 7987 27999
rect 7975 27968 8340 27996
rect 7975 27965 7987 27968
rect 7929 27959 7987 27965
rect 6696 27900 7696 27928
rect 7745 27931 7803 27937
rect 6696 27888 6702 27900
rect 7745 27897 7757 27931
rect 7791 27928 7803 27931
rect 8018 27928 8024 27940
rect 7791 27900 8024 27928
rect 7791 27897 7803 27900
rect 7745 27891 7803 27897
rect 8018 27888 8024 27900
rect 8076 27888 8082 27940
rect 8312 27928 8340 27968
rect 8386 27956 8392 28008
rect 8444 27996 8450 28008
rect 9677 27999 9735 28005
rect 9677 27996 9689 27999
rect 8444 27968 9689 27996
rect 8444 27956 8450 27968
rect 9677 27965 9689 27968
rect 9723 27965 9735 27999
rect 9677 27959 9735 27965
rect 10042 27956 10048 28008
rect 10100 27996 10106 28008
rect 10781 27999 10839 28005
rect 10781 27996 10793 27999
rect 10100 27968 10793 27996
rect 10100 27956 10106 27968
rect 10781 27965 10793 27968
rect 10827 27965 10839 27999
rect 10781 27959 10839 27965
rect 10870 27956 10876 28008
rect 10928 27956 10934 28008
rect 10980 28005 11008 28036
rect 11330 28024 11336 28076
rect 11388 28024 11394 28076
rect 13372 28073 13400 28160
rect 13357 28067 13415 28073
rect 13357 28033 13369 28067
rect 13403 28033 13415 28067
rect 13357 28027 13415 28033
rect 10965 27999 11023 28005
rect 10965 27965 10977 27999
rect 11011 27965 11023 27999
rect 11238 27996 11244 28008
rect 10965 27959 11023 27965
rect 11072 27968 11244 27996
rect 8478 27928 8484 27940
rect 8312 27900 8484 27928
rect 8478 27888 8484 27900
rect 8536 27888 8542 27940
rect 8938 27888 8944 27940
rect 8996 27928 9002 27940
rect 10318 27928 10324 27940
rect 8996 27900 10324 27928
rect 8996 27888 9002 27900
rect 10318 27888 10324 27900
rect 10376 27888 10382 27940
rect 10597 27931 10655 27937
rect 10597 27897 10609 27931
rect 10643 27928 10655 27931
rect 11072 27928 11100 27968
rect 11238 27956 11244 27968
rect 11296 27996 11302 28008
rect 13078 27996 13084 28008
rect 11296 27968 13084 27996
rect 11296 27956 11302 27968
rect 13078 27956 13084 27968
rect 13136 27996 13142 28008
rect 13173 27999 13231 28005
rect 13173 27996 13185 27999
rect 13136 27968 13185 27996
rect 13136 27956 13142 27968
rect 13173 27965 13185 27968
rect 13219 27965 13231 27999
rect 13173 27959 13231 27965
rect 11606 27937 11612 27940
rect 10643 27900 11100 27928
rect 10643 27897 10655 27900
rect 10597 27891 10655 27897
rect 11600 27891 11612 27937
rect 11606 27888 11612 27891
rect 11664 27888 11670 27940
rect 2866 27860 2872 27872
rect 2792 27832 2872 27860
rect 2866 27820 2872 27832
rect 2924 27860 2930 27872
rect 3326 27860 3332 27872
rect 2924 27832 3332 27860
rect 2924 27820 2930 27832
rect 3326 27820 3332 27832
rect 3384 27820 3390 27872
rect 3878 27820 3884 27872
rect 3936 27820 3942 27872
rect 5902 27820 5908 27872
rect 5960 27860 5966 27872
rect 6273 27863 6331 27869
rect 6273 27860 6285 27863
rect 5960 27832 6285 27860
rect 5960 27820 5966 27832
rect 6273 27829 6285 27832
rect 6319 27829 6331 27863
rect 6273 27823 6331 27829
rect 6730 27820 6736 27872
rect 6788 27820 6794 27872
rect 8570 27820 8576 27872
rect 8628 27860 8634 27872
rect 10137 27863 10195 27869
rect 10137 27860 10149 27863
rect 8628 27832 10149 27860
rect 8628 27820 8634 27832
rect 10137 27829 10149 27832
rect 10183 27860 10195 27863
rect 11514 27860 11520 27872
rect 10183 27832 11520 27860
rect 10183 27829 10195 27832
rect 10137 27823 10195 27829
rect 11514 27820 11520 27832
rect 11572 27820 11578 27872
rect 12710 27820 12716 27872
rect 12768 27820 12774 27872
rect 13188 27860 13216 27959
rect 13541 27931 13599 27937
rect 13541 27897 13553 27931
rect 13587 27928 13599 27931
rect 13630 27928 13636 27940
rect 13587 27900 13636 27928
rect 13587 27897 13599 27900
rect 13541 27891 13599 27897
rect 13630 27888 13636 27900
rect 13688 27928 13694 27940
rect 14016 27928 14044 28163
rect 14642 28160 14648 28172
rect 14700 28160 14706 28212
rect 18414 28160 18420 28212
rect 18472 28160 18478 28212
rect 18693 28203 18751 28209
rect 18693 28169 18705 28203
rect 18739 28200 18751 28203
rect 18782 28200 18788 28212
rect 18739 28172 18788 28200
rect 18739 28169 18751 28172
rect 18693 28163 18751 28169
rect 18782 28160 18788 28172
rect 18840 28160 18846 28212
rect 20070 28160 20076 28212
rect 20128 28200 20134 28212
rect 20257 28203 20315 28209
rect 20257 28200 20269 28203
rect 20128 28172 20269 28200
rect 20128 28160 20134 28172
rect 20257 28169 20269 28172
rect 20303 28169 20315 28203
rect 20257 28163 20315 28169
rect 21085 28203 21143 28209
rect 21085 28169 21097 28203
rect 21131 28200 21143 28203
rect 21266 28200 21272 28212
rect 21131 28172 21272 28200
rect 21131 28169 21143 28172
rect 21085 28163 21143 28169
rect 21266 28160 21272 28172
rect 21324 28160 21330 28212
rect 21634 28160 21640 28212
rect 21692 28160 21698 28212
rect 22094 28160 22100 28212
rect 22152 28200 22158 28212
rect 22646 28200 22652 28212
rect 22152 28172 22652 28200
rect 22152 28160 22158 28172
rect 22646 28160 22652 28172
rect 22704 28160 22710 28212
rect 24029 28203 24087 28209
rect 24029 28169 24041 28203
rect 24075 28200 24087 28203
rect 24210 28200 24216 28212
rect 24075 28172 24216 28200
rect 24075 28169 24087 28172
rect 24029 28163 24087 28169
rect 24210 28160 24216 28172
rect 24268 28160 24274 28212
rect 24302 28160 24308 28212
rect 24360 28160 24366 28212
rect 24489 28203 24547 28209
rect 24489 28169 24501 28203
rect 24535 28169 24547 28203
rect 24489 28163 24547 28169
rect 17681 28135 17739 28141
rect 17681 28101 17693 28135
rect 17727 28101 17739 28135
rect 17681 28095 17739 28101
rect 15381 28067 15439 28073
rect 15381 28033 15393 28067
rect 15427 28064 15439 28067
rect 17696 28064 17724 28095
rect 20898 28092 20904 28144
rect 20956 28132 20962 28144
rect 22186 28132 22192 28144
rect 20956 28104 21496 28132
rect 20956 28092 20962 28104
rect 21468 28073 21496 28104
rect 21560 28104 22192 28132
rect 17773 28067 17831 28073
rect 17773 28064 17785 28067
rect 15427 28036 16344 28064
rect 17696 28036 17785 28064
rect 15427 28033 15439 28036
rect 15381 28027 15439 28033
rect 15654 27956 15660 28008
rect 15712 27956 15718 28008
rect 16316 28005 16344 28036
rect 17773 28033 17785 28036
rect 17819 28033 17831 28067
rect 17773 28027 17831 28033
rect 20625 28067 20683 28073
rect 20625 28033 20637 28067
rect 20671 28064 20683 28067
rect 21361 28067 21419 28073
rect 21361 28064 21373 28067
rect 20671 28036 21373 28064
rect 20671 28033 20683 28036
rect 20625 28027 20683 28033
rect 21361 28033 21373 28036
rect 21407 28033 21419 28067
rect 21361 28027 21419 28033
rect 21453 28067 21511 28073
rect 21453 28033 21465 28067
rect 21499 28033 21511 28067
rect 21453 28027 21511 28033
rect 16301 27999 16359 28005
rect 16301 27965 16313 27999
rect 16347 27996 16359 27999
rect 16850 27996 16856 28008
rect 16347 27968 16856 27996
rect 16347 27965 16359 27968
rect 16301 27959 16359 27965
rect 16850 27956 16856 27968
rect 16908 27996 16914 28008
rect 17034 27996 17040 28008
rect 16908 27968 17040 27996
rect 16908 27956 16914 27968
rect 17034 27956 17040 27968
rect 17092 27956 17098 28008
rect 18414 27956 18420 28008
rect 18472 27996 18478 28008
rect 18874 27996 18880 28008
rect 18472 27968 18880 27996
rect 18472 27956 18478 27968
rect 18874 27956 18880 27968
rect 18932 27956 18938 28008
rect 18966 27956 18972 28008
rect 19024 27956 19030 28008
rect 19061 27999 19119 28005
rect 19061 27965 19073 27999
rect 19107 27996 19119 27999
rect 19150 27996 19156 28008
rect 19107 27968 19156 27996
rect 19107 27965 19119 27968
rect 19061 27959 19119 27965
rect 13688 27900 14044 27928
rect 13688 27888 13694 27900
rect 14458 27888 14464 27940
rect 14516 27928 14522 27940
rect 15114 27931 15172 27937
rect 15114 27928 15126 27931
rect 14516 27900 15126 27928
rect 14516 27888 14522 27900
rect 15114 27897 15126 27900
rect 15160 27897 15172 27931
rect 15114 27891 15172 27897
rect 16209 27931 16267 27937
rect 16209 27897 16221 27931
rect 16255 27928 16267 27931
rect 16546 27931 16604 27937
rect 16546 27928 16558 27931
rect 16255 27900 16558 27928
rect 16255 27897 16267 27900
rect 16209 27891 16267 27897
rect 16546 27897 16558 27900
rect 16592 27897 16604 27931
rect 16546 27891 16604 27897
rect 18322 27888 18328 27940
rect 18380 27928 18386 27940
rect 19076 27928 19104 27959
rect 19150 27956 19156 27968
rect 19208 27956 19214 28008
rect 19245 27999 19303 28005
rect 19245 27965 19257 27999
rect 19291 27996 19303 27999
rect 19702 27996 19708 28008
rect 19291 27968 19708 27996
rect 19291 27965 19303 27968
rect 19245 27959 19303 27965
rect 19702 27956 19708 27968
rect 19760 27956 19766 28008
rect 20165 27999 20223 28005
rect 20165 27965 20177 27999
rect 20211 27996 20223 27999
rect 20346 27996 20352 28008
rect 20211 27968 20352 27996
rect 20211 27965 20223 27968
rect 20165 27959 20223 27965
rect 20346 27956 20352 27968
rect 20404 27956 20410 28008
rect 20809 27999 20867 28005
rect 20809 27965 20821 27999
rect 20855 27996 20867 27999
rect 20855 27968 21312 27996
rect 20855 27965 20867 27968
rect 20809 27959 20867 27965
rect 21284 27940 21312 27968
rect 18380 27900 19104 27928
rect 18380 27888 18386 27900
rect 20898 27888 20904 27940
rect 20956 27888 20962 27940
rect 21085 27931 21143 27937
rect 21085 27897 21097 27931
rect 21131 27897 21143 27931
rect 21085 27891 21143 27897
rect 13741 27863 13799 27869
rect 13741 27860 13753 27863
rect 13188 27832 13753 27860
rect 13741 27829 13753 27832
rect 13787 27829 13799 27863
rect 21100 27860 21128 27891
rect 21266 27888 21272 27940
rect 21324 27888 21330 27940
rect 21450 27860 21456 27872
rect 21100 27832 21456 27860
rect 13741 27823 13799 27829
rect 21450 27820 21456 27832
rect 21508 27860 21514 27872
rect 21560 27860 21588 28104
rect 22186 28092 22192 28104
rect 22244 28092 22250 28144
rect 23566 28092 23572 28144
rect 23624 28132 23630 28144
rect 24504 28132 24532 28163
rect 23624 28104 24532 28132
rect 23624 28092 23630 28104
rect 22922 28064 22928 28076
rect 22066 28036 22928 28064
rect 21729 27999 21787 28005
rect 21729 27965 21741 27999
rect 21775 27996 21787 27999
rect 22066 27996 22094 28036
rect 22922 28024 22928 28036
rect 22980 28024 22986 28076
rect 23109 28067 23167 28073
rect 23109 28033 23121 28067
rect 23155 28064 23167 28067
rect 24578 28064 24584 28076
rect 23155 28036 24584 28064
rect 23155 28033 23167 28036
rect 23109 28027 23167 28033
rect 24578 28024 24584 28036
rect 24636 28024 24642 28076
rect 21775 27968 22094 27996
rect 22189 27999 22247 28005
rect 21775 27965 21787 27968
rect 21729 27959 21787 27965
rect 22189 27965 22201 27999
rect 22235 27965 22247 27999
rect 22189 27959 22247 27965
rect 22373 27999 22431 28005
rect 22373 27965 22385 27999
rect 22419 27996 22431 27999
rect 22738 27996 22744 28008
rect 22419 27968 22744 27996
rect 22419 27965 22431 27968
rect 22373 27959 22431 27965
rect 22204 27928 22232 27959
rect 22738 27956 22744 27968
rect 22796 27956 22802 28008
rect 23014 27956 23020 28008
rect 23072 27956 23078 28008
rect 23201 27999 23259 28005
rect 23201 27965 23213 27999
rect 23247 27996 23259 27999
rect 23566 27996 23572 28008
rect 23247 27968 23572 27996
rect 23247 27965 23259 27968
rect 23201 27959 23259 27965
rect 23566 27956 23572 27968
rect 23624 27956 23630 28008
rect 23661 27999 23719 28005
rect 23661 27965 23673 27999
rect 23707 27996 23719 27999
rect 23707 27968 24348 27996
rect 23707 27965 23719 27968
rect 23661 27959 23719 27965
rect 22646 27928 22652 27940
rect 22204 27900 22652 27928
rect 22646 27888 22652 27900
rect 22704 27888 22710 27940
rect 23293 27931 23351 27937
rect 23293 27897 23305 27931
rect 23339 27928 23351 27931
rect 23382 27928 23388 27940
rect 23339 27900 23388 27928
rect 23339 27897 23351 27900
rect 23293 27891 23351 27897
rect 23382 27888 23388 27900
rect 23440 27888 23446 27940
rect 23477 27931 23535 27937
rect 23477 27897 23489 27931
rect 23523 27928 23535 27931
rect 23523 27900 23612 27928
rect 23523 27897 23535 27900
rect 23477 27891 23535 27897
rect 21508 27832 21588 27860
rect 21508 27820 21514 27832
rect 22186 27820 22192 27872
rect 22244 27860 22250 27872
rect 22281 27863 22339 27869
rect 22281 27860 22293 27863
rect 22244 27832 22293 27860
rect 22244 27820 22250 27832
rect 22281 27829 22293 27832
rect 22327 27829 22339 27863
rect 23584 27860 23612 27900
rect 23750 27888 23756 27940
rect 23808 27928 23814 27940
rect 23997 27931 24055 27937
rect 23997 27928 24009 27931
rect 23808 27900 24009 27928
rect 23808 27888 23814 27900
rect 23997 27897 24009 27900
rect 24043 27897 24055 27931
rect 23997 27891 24055 27897
rect 24210 27888 24216 27940
rect 24268 27888 24274 27940
rect 24320 27928 24348 27968
rect 25130 27956 25136 28008
rect 25188 27956 25194 28008
rect 24457 27931 24515 27937
rect 24457 27928 24469 27931
rect 24320 27900 24469 27928
rect 24457 27897 24469 27900
rect 24503 27897 24515 27931
rect 24457 27891 24515 27897
rect 24673 27931 24731 27937
rect 24673 27897 24685 27931
rect 24719 27928 24731 27931
rect 25038 27928 25044 27940
rect 24719 27900 25044 27928
rect 24719 27897 24731 27900
rect 24673 27891 24731 27897
rect 25038 27888 25044 27900
rect 25096 27888 25102 27940
rect 23658 27860 23664 27872
rect 23584 27832 23664 27860
rect 22281 27823 22339 27829
rect 23658 27820 23664 27832
rect 23716 27820 23722 27872
rect 23842 27820 23848 27872
rect 23900 27820 23906 27872
rect 25314 27820 25320 27872
rect 25372 27820 25378 27872
rect 552 27770 27576 27792
rect 552 27718 7114 27770
rect 7166 27718 7178 27770
rect 7230 27718 7242 27770
rect 7294 27718 7306 27770
rect 7358 27718 7370 27770
rect 7422 27718 13830 27770
rect 13882 27718 13894 27770
rect 13946 27718 13958 27770
rect 14010 27718 14022 27770
rect 14074 27718 14086 27770
rect 14138 27718 20546 27770
rect 20598 27718 20610 27770
rect 20662 27718 20674 27770
rect 20726 27718 20738 27770
rect 20790 27718 20802 27770
rect 20854 27718 27262 27770
rect 27314 27718 27326 27770
rect 27378 27718 27390 27770
rect 27442 27718 27454 27770
rect 27506 27718 27518 27770
rect 27570 27718 27576 27770
rect 552 27696 27576 27718
rect 2869 27659 2927 27665
rect 2869 27625 2881 27659
rect 2915 27656 2927 27659
rect 3234 27656 3240 27668
rect 2915 27628 3240 27656
rect 2915 27625 2927 27628
rect 2869 27619 2927 27625
rect 3234 27616 3240 27628
rect 3292 27616 3298 27668
rect 6086 27616 6092 27668
rect 6144 27656 6150 27668
rect 6365 27659 6423 27665
rect 6365 27656 6377 27659
rect 6144 27628 6377 27656
rect 6144 27616 6150 27628
rect 6365 27625 6377 27628
rect 6411 27656 6423 27659
rect 6914 27656 6920 27668
rect 6411 27628 6920 27656
rect 6411 27625 6423 27628
rect 6365 27619 6423 27625
rect 6914 27616 6920 27628
rect 6972 27616 6978 27668
rect 8018 27616 8024 27668
rect 8076 27656 8082 27668
rect 8076 27628 8616 27656
rect 8076 27616 8082 27628
rect 2685 27591 2743 27597
rect 2685 27557 2697 27591
rect 2731 27557 2743 27591
rect 2685 27551 2743 27557
rect 3780 27591 3838 27597
rect 3780 27557 3792 27591
rect 3826 27588 3838 27591
rect 3878 27588 3884 27600
rect 3826 27560 3884 27588
rect 3826 27557 3838 27560
rect 3780 27551 3838 27557
rect 1854 27480 1860 27532
rect 1912 27520 1918 27532
rect 2700 27520 2728 27551
rect 3878 27548 3884 27560
rect 3936 27548 3942 27600
rect 5261 27591 5319 27597
rect 5261 27557 5273 27591
rect 5307 27588 5319 27591
rect 5718 27588 5724 27600
rect 5307 27560 5724 27588
rect 5307 27557 5319 27560
rect 5261 27551 5319 27557
rect 5718 27548 5724 27560
rect 5776 27548 5782 27600
rect 6822 27588 6828 27600
rect 5828 27560 6828 27588
rect 1912 27492 2728 27520
rect 3145 27523 3203 27529
rect 1912 27480 1918 27492
rect 3145 27489 3157 27523
rect 3191 27520 3203 27523
rect 3234 27520 3240 27532
rect 3191 27492 3240 27520
rect 3191 27489 3203 27492
rect 3145 27483 3203 27489
rect 3234 27480 3240 27492
rect 3292 27480 3298 27532
rect 3513 27523 3571 27529
rect 3513 27489 3525 27523
rect 3559 27520 3571 27523
rect 3602 27520 3608 27532
rect 3559 27492 3608 27520
rect 3559 27489 3571 27492
rect 3513 27483 3571 27489
rect 3602 27480 3608 27492
rect 3660 27480 3666 27532
rect 5350 27480 5356 27532
rect 5408 27480 5414 27532
rect 5445 27523 5503 27529
rect 5445 27489 5457 27523
rect 5491 27520 5503 27523
rect 5828 27520 5856 27560
rect 6822 27548 6828 27560
rect 6880 27548 6886 27600
rect 8588 27597 8616 27628
rect 11606 27616 11612 27668
rect 11664 27616 11670 27668
rect 14458 27616 14464 27668
rect 14516 27616 14522 27668
rect 15654 27616 15660 27668
rect 15712 27656 15718 27668
rect 16393 27659 16451 27665
rect 16393 27656 16405 27659
rect 15712 27628 16405 27656
rect 15712 27616 15718 27628
rect 16393 27625 16405 27628
rect 16439 27625 16451 27659
rect 21358 27656 21364 27668
rect 16393 27619 16451 27625
rect 17696 27628 21364 27656
rect 8573 27591 8631 27597
rect 8573 27557 8585 27591
rect 8619 27557 8631 27591
rect 8573 27551 8631 27557
rect 11146 27548 11152 27600
rect 11204 27588 11210 27600
rect 12710 27588 12716 27600
rect 11204 27560 12716 27588
rect 11204 27548 11210 27560
rect 5491 27492 5856 27520
rect 5491 27489 5503 27492
rect 5445 27483 5503 27489
rect 5902 27480 5908 27532
rect 5960 27480 5966 27532
rect 6178 27480 6184 27532
rect 6236 27520 6242 27532
rect 6273 27523 6331 27529
rect 6273 27520 6285 27523
rect 6236 27492 6285 27520
rect 6236 27480 6242 27492
rect 6273 27489 6285 27492
rect 6319 27489 6331 27523
rect 6273 27483 6331 27489
rect 7006 27480 7012 27532
rect 7064 27520 7070 27532
rect 7478 27523 7536 27529
rect 7478 27520 7490 27523
rect 7064 27492 7490 27520
rect 7064 27480 7070 27492
rect 7478 27489 7490 27492
rect 7524 27489 7536 27523
rect 7478 27483 7536 27489
rect 10689 27523 10747 27529
rect 10689 27489 10701 27523
rect 10735 27520 10747 27523
rect 10870 27520 10876 27532
rect 10735 27492 10876 27520
rect 10735 27489 10747 27492
rect 10689 27483 10747 27489
rect 10870 27480 10876 27492
rect 10928 27480 10934 27532
rect 11790 27480 11796 27532
rect 11848 27480 11854 27532
rect 12084 27529 12112 27560
rect 12710 27548 12716 27560
rect 12768 27548 12774 27600
rect 16485 27591 16543 27597
rect 16485 27557 16497 27591
rect 16531 27588 16543 27591
rect 16758 27588 16764 27600
rect 16531 27560 16764 27588
rect 16531 27557 16543 27560
rect 16485 27551 16543 27557
rect 16758 27548 16764 27560
rect 16816 27588 16822 27600
rect 17586 27588 17592 27600
rect 16816 27560 17592 27588
rect 16816 27548 16822 27560
rect 17586 27548 17592 27560
rect 17644 27548 17650 27600
rect 12069 27523 12127 27529
rect 12069 27489 12081 27523
rect 12115 27489 12127 27523
rect 12069 27483 12127 27489
rect 13173 27523 13231 27529
rect 13173 27489 13185 27523
rect 13219 27520 13231 27523
rect 13354 27520 13360 27532
rect 13219 27492 13360 27520
rect 13219 27489 13231 27492
rect 13173 27483 13231 27489
rect 13354 27480 13360 27492
rect 13412 27480 13418 27532
rect 13630 27480 13636 27532
rect 13688 27520 13694 27532
rect 13725 27523 13783 27529
rect 13725 27520 13737 27523
rect 13688 27492 13737 27520
rect 13688 27480 13694 27492
rect 13725 27489 13737 27492
rect 13771 27489 13783 27523
rect 13725 27483 13783 27489
rect 14274 27480 14280 27532
rect 14332 27480 14338 27532
rect 14921 27523 14979 27529
rect 14921 27489 14933 27523
rect 14967 27520 14979 27523
rect 15102 27520 15108 27532
rect 14967 27492 15108 27520
rect 14967 27489 14979 27492
rect 14921 27483 14979 27489
rect 15102 27480 15108 27492
rect 15160 27480 15166 27532
rect 15470 27480 15476 27532
rect 15528 27520 15534 27532
rect 15657 27523 15715 27529
rect 15657 27520 15669 27523
rect 15528 27492 15669 27520
rect 15528 27480 15534 27492
rect 15657 27489 15669 27492
rect 15703 27489 15715 27523
rect 15657 27483 15715 27489
rect 15838 27480 15844 27532
rect 15896 27520 15902 27532
rect 16117 27523 16175 27529
rect 16117 27520 16129 27523
rect 15896 27492 16129 27520
rect 15896 27480 15902 27492
rect 16117 27489 16129 27492
rect 16163 27489 16175 27523
rect 16117 27483 16175 27489
rect 16577 27523 16635 27529
rect 16577 27489 16589 27523
rect 16623 27520 16635 27523
rect 16666 27520 16672 27532
rect 16623 27492 16672 27520
rect 16623 27489 16635 27492
rect 16577 27483 16635 27489
rect 16666 27480 16672 27492
rect 16724 27480 16730 27532
rect 17696 27520 17724 27628
rect 21358 27616 21364 27628
rect 21416 27616 21422 27668
rect 23477 27659 23535 27665
rect 21560 27628 21680 27656
rect 21453 27591 21511 27597
rect 21453 27588 21465 27591
rect 17880 27560 18736 27588
rect 16776 27492 17724 27520
rect 3050 27452 3056 27464
rect 2056 27424 3056 27452
rect 2056 27396 2084 27424
rect 3050 27412 3056 27424
rect 3108 27412 3114 27464
rect 3326 27412 3332 27464
rect 3384 27412 3390 27464
rect 5626 27412 5632 27464
rect 5684 27452 5690 27464
rect 5997 27455 6055 27461
rect 5997 27452 6009 27455
rect 5684 27424 6009 27452
rect 5684 27412 5690 27424
rect 5997 27421 6009 27424
rect 6043 27421 6055 27455
rect 5997 27415 6055 27421
rect 7745 27455 7803 27461
rect 7745 27421 7757 27455
rect 7791 27452 7803 27455
rect 8386 27452 8392 27464
rect 7791 27424 8392 27452
rect 7791 27421 7803 27424
rect 7745 27415 7803 27421
rect 8386 27412 8392 27424
rect 8444 27412 8450 27464
rect 8478 27412 8484 27464
rect 8536 27452 8542 27464
rect 9585 27455 9643 27461
rect 9585 27452 9597 27455
rect 8536 27424 9597 27452
rect 8536 27412 8542 27424
rect 9585 27421 9597 27424
rect 9631 27421 9643 27455
rect 9585 27415 9643 27421
rect 9766 27412 9772 27464
rect 9824 27452 9830 27464
rect 16776 27452 16804 27492
rect 17770 27480 17776 27532
rect 17828 27480 17834 27532
rect 17880 27529 17908 27560
rect 18708 27532 18736 27560
rect 21284 27560 21465 27588
rect 17865 27523 17923 27529
rect 17865 27489 17877 27523
rect 17911 27489 17923 27523
rect 17865 27483 17923 27489
rect 17954 27480 17960 27532
rect 18012 27520 18018 27532
rect 18121 27523 18179 27529
rect 18121 27520 18133 27523
rect 18012 27492 18133 27520
rect 18012 27480 18018 27492
rect 18121 27489 18133 27492
rect 18167 27489 18179 27523
rect 18121 27483 18179 27489
rect 18690 27480 18696 27532
rect 18748 27520 18754 27532
rect 19334 27520 19340 27532
rect 18748 27492 19340 27520
rect 18748 27480 18754 27492
rect 19334 27480 19340 27492
rect 19392 27480 19398 27532
rect 19426 27480 19432 27532
rect 19484 27520 19490 27532
rect 19593 27523 19651 27529
rect 19593 27520 19605 27523
rect 19484 27492 19605 27520
rect 19484 27480 19490 27492
rect 19593 27489 19605 27492
rect 19639 27489 19651 27523
rect 19593 27483 19651 27489
rect 9824 27424 16804 27452
rect 9824 27412 9830 27424
rect 17034 27412 17040 27464
rect 17092 27412 17098 27464
rect 21284 27452 21312 27560
rect 21453 27557 21465 27560
rect 21499 27557 21511 27591
rect 21453 27551 21511 27557
rect 21361 27523 21419 27529
rect 21361 27489 21373 27523
rect 21407 27520 21419 27523
rect 21560 27520 21588 27628
rect 21652 27588 21680 27628
rect 23477 27625 23489 27659
rect 23523 27656 23535 27659
rect 23566 27656 23572 27668
rect 23523 27628 23572 27656
rect 23523 27625 23535 27628
rect 23477 27619 23535 27625
rect 23566 27616 23572 27628
rect 23624 27616 23630 27668
rect 24210 27616 24216 27668
rect 24268 27656 24274 27668
rect 24857 27659 24915 27665
rect 24857 27656 24869 27659
rect 24268 27628 24869 27656
rect 24268 27616 24274 27628
rect 24857 27625 24869 27628
rect 24903 27625 24915 27659
rect 24857 27619 24915 27625
rect 22094 27588 22100 27600
rect 21652 27560 22100 27588
rect 22094 27548 22100 27560
rect 22152 27588 22158 27600
rect 22373 27591 22431 27597
rect 22373 27588 22385 27591
rect 22152 27560 22385 27588
rect 22152 27548 22158 27560
rect 22373 27557 22385 27560
rect 22419 27557 22431 27591
rect 23658 27588 23664 27600
rect 22373 27551 22431 27557
rect 23400 27560 23664 27588
rect 21407 27492 21588 27520
rect 21637 27523 21695 27529
rect 21407 27489 21419 27492
rect 21361 27483 21419 27489
rect 21637 27489 21649 27523
rect 21683 27489 21695 27523
rect 21637 27483 21695 27489
rect 21913 27523 21971 27529
rect 21913 27489 21925 27523
rect 21959 27520 21971 27523
rect 22186 27520 22192 27532
rect 21959 27492 22192 27520
rect 21959 27489 21971 27492
rect 21913 27483 21971 27489
rect 21542 27452 21548 27464
rect 21284 27424 21548 27452
rect 21542 27412 21548 27424
rect 21600 27412 21606 27464
rect 21652 27452 21680 27483
rect 22186 27480 22192 27492
rect 22244 27480 22250 27532
rect 22646 27480 22652 27532
rect 22704 27480 22710 27532
rect 22738 27480 22744 27532
rect 22796 27480 22802 27532
rect 22830 27480 22836 27532
rect 22888 27480 22894 27532
rect 23014 27480 23020 27532
rect 23072 27480 23078 27532
rect 23400 27529 23428 27560
rect 23658 27548 23664 27560
rect 23716 27588 23722 27600
rect 24118 27588 24124 27600
rect 23716 27560 24124 27588
rect 23716 27548 23722 27560
rect 24118 27548 24124 27560
rect 24176 27548 24182 27600
rect 23385 27523 23443 27529
rect 23385 27489 23397 27523
rect 23431 27489 23443 27523
rect 23385 27483 23443 27489
rect 23474 27480 23480 27532
rect 23532 27520 23538 27532
rect 23569 27523 23627 27529
rect 23569 27520 23581 27523
rect 23532 27492 23581 27520
rect 23532 27480 23538 27492
rect 23569 27489 23581 27492
rect 23615 27489 23627 27523
rect 23569 27483 23627 27489
rect 23845 27523 23903 27529
rect 23845 27489 23857 27523
rect 23891 27520 23903 27523
rect 24228 27520 24256 27616
rect 24581 27591 24639 27597
rect 24581 27557 24593 27591
rect 24627 27588 24639 27591
rect 25038 27588 25044 27600
rect 24627 27560 25044 27588
rect 24627 27557 24639 27560
rect 24581 27551 24639 27557
rect 25038 27548 25044 27560
rect 25096 27548 25102 27600
rect 25314 27548 25320 27600
rect 25372 27588 25378 27600
rect 25970 27591 26028 27597
rect 25970 27588 25982 27591
rect 25372 27560 25982 27588
rect 25372 27548 25378 27560
rect 25970 27557 25982 27560
rect 26016 27557 26028 27591
rect 25970 27551 26028 27557
rect 23891 27492 24256 27520
rect 23891 27489 23903 27492
rect 23845 27483 23903 27489
rect 26142 27480 26148 27532
rect 26200 27520 26206 27532
rect 26237 27523 26295 27529
rect 26237 27520 26249 27523
rect 26200 27492 26249 27520
rect 26200 27480 26206 27492
rect 26237 27489 26249 27492
rect 26283 27489 26295 27523
rect 26237 27483 26295 27489
rect 22005 27455 22063 27461
rect 22005 27452 22017 27455
rect 21652 27424 22017 27452
rect 22005 27421 22017 27424
rect 22051 27421 22063 27455
rect 23032 27452 23060 27480
rect 23753 27455 23811 27461
rect 23753 27452 23765 27455
rect 23032 27424 23765 27452
rect 22005 27415 22063 27421
rect 23753 27421 23765 27424
rect 23799 27421 23811 27455
rect 23753 27415 23811 27421
rect 2038 27344 2044 27396
rect 2096 27344 2102 27396
rect 2317 27387 2375 27393
rect 2317 27353 2329 27387
rect 2363 27384 2375 27387
rect 5077 27387 5135 27393
rect 2363 27356 3004 27384
rect 2363 27353 2375 27356
rect 2317 27347 2375 27353
rect 2682 27276 2688 27328
rect 2740 27276 2746 27328
rect 2976 27325 3004 27356
rect 5077 27353 5089 27387
rect 5123 27353 5135 27387
rect 5077 27347 5135 27353
rect 8941 27387 8999 27393
rect 8941 27353 8953 27387
rect 8987 27384 8999 27387
rect 8987 27356 9260 27384
rect 8987 27353 8999 27356
rect 8941 27347 8999 27353
rect 2961 27319 3019 27325
rect 2961 27285 2973 27319
rect 3007 27316 3019 27319
rect 3142 27316 3148 27328
rect 3007 27288 3148 27316
rect 3007 27285 3019 27288
rect 2961 27279 3019 27285
rect 3142 27276 3148 27288
rect 3200 27276 3206 27328
rect 4890 27276 4896 27328
rect 4948 27316 4954 27328
rect 5092 27316 5120 27347
rect 4948 27288 5120 27316
rect 4948 27276 4954 27288
rect 5166 27276 5172 27328
rect 5224 27316 5230 27328
rect 5629 27319 5687 27325
rect 5629 27316 5641 27319
rect 5224 27288 5641 27316
rect 5224 27276 5230 27288
rect 5629 27285 5641 27288
rect 5675 27285 5687 27319
rect 5629 27279 5687 27285
rect 5810 27276 5816 27328
rect 5868 27276 5874 27328
rect 6178 27276 6184 27328
rect 6236 27276 6242 27328
rect 9030 27276 9036 27328
rect 9088 27276 9094 27328
rect 9122 27276 9128 27328
rect 9180 27276 9186 27328
rect 9232 27316 9260 27356
rect 9306 27344 9312 27396
rect 9364 27344 9370 27396
rect 16850 27344 16856 27396
rect 16908 27384 16914 27396
rect 17126 27384 17132 27396
rect 16908 27356 17132 27384
rect 16908 27344 16914 27356
rect 17126 27344 17132 27356
rect 17184 27344 17190 27396
rect 21174 27344 21180 27396
rect 21232 27384 21238 27396
rect 21232 27356 21772 27384
rect 21232 27344 21238 27356
rect 9858 27316 9864 27328
rect 9232 27288 9864 27316
rect 9858 27276 9864 27288
rect 9916 27276 9922 27328
rect 10597 27319 10655 27325
rect 10597 27285 10609 27319
rect 10643 27316 10655 27319
rect 10870 27316 10876 27328
rect 10643 27288 10876 27316
rect 10643 27285 10655 27288
rect 10597 27279 10655 27285
rect 10870 27276 10876 27288
rect 10928 27276 10934 27328
rect 11974 27276 11980 27328
rect 12032 27276 12038 27328
rect 12986 27276 12992 27328
rect 13044 27316 13050 27328
rect 13081 27319 13139 27325
rect 13081 27316 13093 27319
rect 13044 27288 13093 27316
rect 13044 27276 13050 27288
rect 13081 27285 13093 27288
rect 13127 27285 13139 27319
rect 13081 27279 13139 27285
rect 13633 27319 13691 27325
rect 13633 27285 13645 27319
rect 13679 27316 13691 27319
rect 13814 27316 13820 27328
rect 13679 27288 13820 27316
rect 13679 27285 13691 27288
rect 13633 27279 13691 27285
rect 13814 27276 13820 27288
rect 13872 27276 13878 27328
rect 14829 27319 14887 27325
rect 14829 27285 14841 27319
rect 14875 27316 14887 27319
rect 14918 27316 14924 27328
rect 14875 27288 14924 27316
rect 14875 27285 14887 27288
rect 14829 27279 14887 27285
rect 14918 27276 14924 27288
rect 14976 27276 14982 27328
rect 15565 27319 15623 27325
rect 15565 27285 15577 27319
rect 15611 27316 15623 27319
rect 15654 27316 15660 27328
rect 15611 27288 15660 27316
rect 15611 27285 15623 27288
rect 15565 27279 15623 27285
rect 15654 27276 15660 27288
rect 15712 27276 15718 27328
rect 19242 27276 19248 27328
rect 19300 27276 19306 27328
rect 20714 27276 20720 27328
rect 20772 27276 20778 27328
rect 21542 27276 21548 27328
rect 21600 27316 21606 27328
rect 21744 27325 21772 27356
rect 21637 27319 21695 27325
rect 21637 27316 21649 27319
rect 21600 27288 21649 27316
rect 21600 27276 21606 27288
rect 21637 27285 21649 27288
rect 21683 27285 21695 27319
rect 21637 27279 21695 27285
rect 21729 27319 21787 27325
rect 21729 27285 21741 27319
rect 21775 27285 21787 27319
rect 22020 27316 22048 27415
rect 22465 27387 22523 27393
rect 22465 27384 22477 27387
rect 22204 27356 22477 27384
rect 22204 27316 22232 27356
rect 22465 27353 22477 27356
rect 22511 27353 22523 27387
rect 22465 27347 22523 27353
rect 23842 27344 23848 27396
rect 23900 27384 23906 27396
rect 24213 27387 24271 27393
rect 24213 27384 24225 27387
rect 23900 27356 24225 27384
rect 23900 27344 23906 27356
rect 24213 27353 24225 27356
rect 24259 27353 24271 27387
rect 24213 27347 24271 27353
rect 24765 27387 24823 27393
rect 24765 27353 24777 27387
rect 24811 27384 24823 27387
rect 25130 27384 25136 27396
rect 24811 27356 25136 27384
rect 24811 27353 24823 27356
rect 24765 27347 24823 27353
rect 25130 27344 25136 27356
rect 25188 27344 25194 27396
rect 22020 27288 22232 27316
rect 21729 27279 21787 27285
rect 22278 27276 22284 27328
rect 22336 27276 22342 27328
rect 24578 27276 24584 27328
rect 24636 27276 24642 27328
rect 552 27226 27416 27248
rect 552 27174 3756 27226
rect 3808 27174 3820 27226
rect 3872 27174 3884 27226
rect 3936 27174 3948 27226
rect 4000 27174 4012 27226
rect 4064 27174 10472 27226
rect 10524 27174 10536 27226
rect 10588 27174 10600 27226
rect 10652 27174 10664 27226
rect 10716 27174 10728 27226
rect 10780 27174 17188 27226
rect 17240 27174 17252 27226
rect 17304 27174 17316 27226
rect 17368 27174 17380 27226
rect 17432 27174 17444 27226
rect 17496 27174 23904 27226
rect 23956 27174 23968 27226
rect 24020 27174 24032 27226
rect 24084 27174 24096 27226
rect 24148 27174 24160 27226
rect 24212 27174 27416 27226
rect 552 27152 27416 27174
rect 2501 27115 2559 27121
rect 2501 27081 2513 27115
rect 2547 27112 2559 27115
rect 2774 27112 2780 27124
rect 2547 27084 2780 27112
rect 2547 27081 2559 27084
rect 2501 27075 2559 27081
rect 2774 27072 2780 27084
rect 2832 27072 2838 27124
rect 3973 27115 4031 27121
rect 3973 27081 3985 27115
rect 4019 27081 4031 27115
rect 3973 27075 4031 27081
rect 3988 27044 4016 27075
rect 4154 27072 4160 27124
rect 4212 27072 4218 27124
rect 5626 27072 5632 27124
rect 5684 27072 5690 27124
rect 5718 27072 5724 27124
rect 5776 27112 5782 27124
rect 5813 27115 5871 27121
rect 5813 27112 5825 27115
rect 5776 27084 5825 27112
rect 5776 27072 5782 27084
rect 5813 27081 5825 27084
rect 5859 27081 5871 27115
rect 7561 27115 7619 27121
rect 7561 27112 7573 27115
rect 5813 27075 5871 27081
rect 6656 27084 7573 27112
rect 4525 27047 4583 27053
rect 4525 27044 4537 27047
rect 3988 27016 4537 27044
rect 4525 27013 4537 27016
rect 4571 27013 4583 27047
rect 5166 27044 5172 27056
rect 4525 27007 4583 27013
rect 4632 27016 5172 27044
rect 3050 26936 3056 26988
rect 3108 26976 3114 26988
rect 3234 26976 3240 26988
rect 3108 26948 3240 26976
rect 3108 26936 3114 26948
rect 3234 26936 3240 26948
rect 3292 26976 3298 26988
rect 3605 26979 3663 26985
rect 3605 26976 3617 26979
rect 3292 26948 3617 26976
rect 3292 26936 3298 26948
rect 3605 26945 3617 26948
rect 3651 26976 3663 26979
rect 4632 26976 4660 27016
rect 5166 27004 5172 27016
rect 5224 27004 5230 27056
rect 3651 26948 4660 26976
rect 4801 26979 4859 26985
rect 3651 26945 3663 26948
rect 3605 26939 3663 26945
rect 4801 26945 4813 26979
rect 4847 26976 4859 26979
rect 5350 26976 5356 26988
rect 4847 26948 5356 26976
rect 4847 26945 4859 26948
rect 4801 26939 4859 26945
rect 5350 26936 5356 26948
rect 5408 26936 5414 26988
rect 842 26868 848 26920
rect 900 26868 906 26920
rect 2406 26868 2412 26920
rect 2464 26908 2470 26920
rect 2869 26911 2927 26917
rect 2869 26908 2881 26911
rect 2464 26880 2881 26908
rect 2464 26868 2470 26880
rect 2869 26877 2881 26880
rect 2915 26877 2927 26911
rect 2869 26871 2927 26877
rect 4709 26911 4767 26917
rect 4709 26877 4721 26911
rect 4755 26877 4767 26911
rect 4709 26871 4767 26877
rect 4893 26911 4951 26917
rect 4893 26877 4905 26911
rect 4939 26877 4951 26911
rect 4893 26871 4951 26877
rect 1118 26849 1124 26852
rect 1112 26803 1124 26849
rect 1118 26800 1124 26803
rect 1176 26800 1182 26852
rect 1486 26800 1492 26852
rect 1544 26840 1550 26852
rect 1854 26840 1860 26852
rect 1544 26812 1860 26840
rect 1544 26800 1550 26812
rect 1854 26800 1860 26812
rect 1912 26840 1918 26852
rect 2501 26843 2559 26849
rect 2501 26840 2513 26843
rect 1912 26812 2513 26840
rect 1912 26800 1918 26812
rect 2501 26809 2513 26812
rect 2547 26840 2559 26843
rect 3973 26843 4031 26849
rect 3973 26840 3985 26843
rect 2547 26812 3985 26840
rect 2547 26809 2559 26812
rect 2501 26803 2559 26809
rect 3973 26809 3985 26812
rect 4019 26809 4031 26843
rect 3973 26803 4031 26809
rect 2222 26732 2228 26784
rect 2280 26732 2286 26784
rect 2314 26732 2320 26784
rect 2372 26732 2378 26784
rect 4724 26772 4752 26871
rect 4908 26840 4936 26871
rect 4982 26868 4988 26920
rect 5040 26868 5046 26920
rect 5736 26908 5764 27072
rect 6656 27044 6684 27084
rect 7561 27081 7573 27084
rect 7607 27081 7619 27115
rect 7561 27075 7619 27081
rect 8757 27115 8815 27121
rect 8757 27081 8769 27115
rect 8803 27112 8815 27115
rect 9306 27112 9312 27124
rect 8803 27084 9312 27112
rect 8803 27081 8815 27084
rect 8757 27075 8815 27081
rect 9306 27072 9312 27084
rect 9364 27112 9370 27124
rect 10042 27112 10048 27124
rect 9364 27084 10048 27112
rect 9364 27072 9370 27084
rect 10042 27072 10048 27084
rect 10100 27072 10106 27124
rect 14553 27115 14611 27121
rect 14553 27081 14565 27115
rect 14599 27112 14611 27115
rect 16298 27112 16304 27124
rect 14599 27084 16304 27112
rect 14599 27081 14611 27084
rect 14553 27075 14611 27081
rect 16298 27072 16304 27084
rect 16356 27072 16362 27124
rect 17773 27115 17831 27121
rect 17773 27081 17785 27115
rect 17819 27112 17831 27115
rect 17954 27112 17960 27124
rect 17819 27084 17960 27112
rect 17819 27081 17831 27084
rect 17773 27075 17831 27081
rect 17954 27072 17960 27084
rect 18012 27072 18018 27124
rect 18509 27115 18567 27121
rect 18509 27081 18521 27115
rect 18555 27112 18567 27115
rect 19426 27112 19432 27124
rect 18555 27084 19432 27112
rect 18555 27081 18567 27084
rect 18509 27075 18567 27081
rect 19426 27072 19432 27084
rect 19484 27072 19490 27124
rect 21450 27072 21456 27124
rect 21508 27072 21514 27124
rect 21821 27115 21879 27121
rect 21821 27081 21833 27115
rect 21867 27112 21879 27115
rect 22094 27112 22100 27124
rect 21867 27084 22100 27112
rect 21867 27081 21879 27084
rect 21821 27075 21879 27081
rect 22094 27072 22100 27084
rect 22152 27072 22158 27124
rect 22738 27072 22744 27124
rect 22796 27112 22802 27124
rect 23201 27115 23259 27121
rect 23201 27112 23213 27115
rect 22796 27084 23213 27112
rect 22796 27072 22802 27084
rect 23201 27081 23213 27084
rect 23247 27081 23259 27115
rect 23201 27075 23259 27081
rect 24213 27115 24271 27121
rect 24213 27081 24225 27115
rect 24259 27112 24271 27115
rect 25133 27115 25191 27121
rect 25133 27112 25145 27115
rect 24259 27084 25145 27112
rect 24259 27081 24271 27084
rect 24213 27075 24271 27081
rect 25133 27081 25145 27084
rect 25179 27081 25191 27115
rect 25133 27075 25191 27081
rect 6288 27016 6684 27044
rect 6288 26976 6316 27016
rect 9122 27004 9128 27056
rect 9180 27004 9186 27056
rect 10321 27047 10379 27053
rect 10321 27013 10333 27047
rect 10367 27013 10379 27047
rect 10321 27007 10379 27013
rect 15105 27047 15163 27053
rect 15105 27013 15117 27047
rect 15151 27044 15163 27047
rect 15562 27044 15568 27056
rect 15151 27016 15568 27044
rect 15151 27013 15163 27016
rect 15105 27007 15163 27013
rect 6196 26948 6316 26976
rect 5092 26880 5764 26908
rect 5092 26840 5120 26880
rect 6086 26868 6092 26920
rect 6144 26868 6150 26920
rect 6196 26917 6224 26948
rect 6362 26936 6368 26988
rect 6420 26976 6426 26988
rect 6420 26948 6592 26976
rect 6420 26936 6426 26948
rect 6564 26917 6592 26948
rect 6914 26936 6920 26988
rect 6972 26936 6978 26988
rect 9140 26976 9168 27004
rect 9048 26948 9168 26976
rect 6181 26911 6239 26917
rect 6181 26877 6193 26911
rect 6227 26877 6239 26911
rect 6457 26911 6515 26917
rect 6457 26908 6469 26911
rect 6181 26871 6239 26877
rect 6288 26880 6469 26908
rect 4908 26812 5120 26840
rect 5718 26800 5724 26852
rect 5776 26840 5782 26852
rect 6288 26840 6316 26880
rect 6457 26877 6469 26880
rect 6503 26877 6515 26911
rect 6457 26871 6515 26877
rect 6549 26911 6607 26917
rect 6549 26877 6561 26911
rect 6595 26877 6607 26911
rect 6549 26871 6607 26877
rect 8110 26868 8116 26920
rect 8168 26868 8174 26920
rect 8478 26868 8484 26920
rect 8536 26868 8542 26920
rect 9048 26917 9076 26948
rect 9033 26911 9091 26917
rect 9033 26877 9045 26911
rect 9079 26877 9091 26911
rect 9033 26871 9091 26877
rect 9122 26868 9128 26920
rect 9180 26908 9186 26920
rect 9539 26911 9597 26917
rect 9180 26880 9225 26908
rect 9180 26868 9186 26880
rect 9539 26877 9551 26911
rect 9585 26908 9597 26911
rect 9585 26880 9720 26908
rect 9585 26877 9597 26880
rect 9539 26871 9597 26877
rect 5776 26812 6316 26840
rect 6365 26843 6423 26849
rect 5776 26800 5782 26812
rect 6365 26809 6377 26843
rect 6411 26840 6423 26843
rect 6914 26840 6920 26852
rect 6411 26812 6920 26840
rect 6411 26809 6423 26812
rect 6365 26803 6423 26809
rect 6914 26800 6920 26812
rect 6972 26800 6978 26852
rect 9309 26843 9367 26849
rect 9309 26809 9321 26843
rect 9355 26809 9367 26843
rect 9309 26803 9367 26809
rect 5534 26772 5540 26784
rect 4724 26744 5540 26772
rect 5534 26732 5540 26744
rect 5592 26772 5598 26784
rect 5902 26772 5908 26784
rect 5592 26744 5908 26772
rect 5592 26732 5598 26744
rect 5902 26732 5908 26744
rect 5960 26732 5966 26784
rect 6086 26732 6092 26784
rect 6144 26772 6150 26784
rect 6270 26772 6276 26784
rect 6144 26744 6276 26772
rect 6144 26732 6150 26744
rect 6270 26732 6276 26744
rect 6328 26732 6334 26784
rect 6733 26775 6791 26781
rect 6733 26741 6745 26775
rect 6779 26772 6791 26775
rect 6822 26772 6828 26784
rect 6779 26744 6828 26772
rect 6779 26741 6791 26744
rect 6733 26735 6791 26741
rect 6822 26732 6828 26744
rect 6880 26732 6886 26784
rect 7466 26732 7472 26784
rect 7524 26732 7530 26784
rect 8941 26775 8999 26781
rect 8941 26741 8953 26775
rect 8987 26772 8999 26775
rect 9324 26772 9352 26803
rect 9398 26800 9404 26852
rect 9456 26800 9462 26852
rect 9692 26840 9720 26880
rect 9766 26868 9772 26920
rect 9824 26868 9830 26920
rect 10045 26911 10103 26917
rect 10045 26877 10057 26911
rect 10091 26908 10103 26911
rect 10336 26908 10364 27007
rect 15562 27004 15568 27016
rect 15620 27004 15626 27056
rect 18322 27044 18328 27056
rect 17420 27016 18328 27044
rect 11701 26979 11759 26985
rect 11701 26945 11713 26979
rect 11747 26976 11759 26979
rect 12802 26976 12808 26988
rect 11747 26948 12808 26976
rect 11747 26945 11759 26948
rect 11701 26939 11759 26945
rect 10091 26880 10364 26908
rect 10091 26877 10103 26880
rect 10045 26871 10103 26877
rect 10502 26868 10508 26920
rect 10560 26868 10566 26920
rect 10597 26911 10655 26917
rect 10597 26877 10609 26911
rect 10643 26908 10655 26911
rect 10778 26908 10784 26920
rect 10643 26880 10784 26908
rect 10643 26877 10655 26880
rect 10597 26871 10655 26877
rect 10778 26868 10784 26880
rect 10836 26868 10842 26920
rect 10873 26911 10931 26917
rect 10873 26877 10885 26911
rect 10919 26908 10931 26911
rect 11054 26908 11060 26920
rect 10919 26880 11060 26908
rect 10919 26877 10931 26880
rect 10873 26871 10931 26877
rect 11054 26868 11060 26880
rect 11112 26868 11118 26920
rect 11146 26868 11152 26920
rect 11204 26908 11210 26920
rect 11425 26911 11483 26917
rect 11425 26908 11437 26911
rect 11204 26880 11437 26908
rect 11204 26868 11210 26880
rect 11425 26877 11437 26880
rect 11471 26877 11483 26911
rect 11425 26871 11483 26877
rect 11517 26911 11575 26917
rect 11517 26877 11529 26911
rect 11563 26877 11575 26911
rect 11517 26871 11575 26877
rect 11793 26911 11851 26917
rect 11793 26877 11805 26911
rect 11839 26908 11851 26911
rect 11974 26908 11980 26920
rect 11839 26880 11980 26908
rect 11839 26877 11851 26880
rect 11793 26871 11851 26877
rect 10134 26840 10140 26852
rect 9692 26812 10140 26840
rect 10134 26800 10140 26812
rect 10192 26800 10198 26852
rect 10689 26843 10747 26849
rect 10689 26809 10701 26843
rect 10735 26809 10747 26843
rect 11072 26840 11100 26868
rect 11532 26840 11560 26871
rect 11974 26868 11980 26880
rect 12032 26868 12038 26920
rect 12176 26917 12204 26948
rect 12802 26936 12808 26948
rect 12860 26936 12866 26988
rect 13173 26979 13231 26985
rect 13173 26945 13185 26979
rect 13219 26945 13231 26979
rect 13173 26939 13231 26945
rect 13280 26948 13860 26976
rect 12161 26911 12219 26917
rect 12161 26877 12173 26911
rect 12207 26877 12219 26911
rect 12161 26871 12219 26877
rect 12345 26911 12403 26917
rect 12345 26877 12357 26911
rect 12391 26908 12403 26911
rect 12894 26908 12900 26920
rect 12391 26880 12900 26908
rect 12391 26877 12403 26880
rect 12345 26871 12403 26877
rect 12894 26868 12900 26880
rect 12952 26868 12958 26920
rect 12986 26868 12992 26920
rect 13044 26868 13050 26920
rect 11072 26812 11560 26840
rect 12253 26843 12311 26849
rect 10689 26803 10747 26809
rect 12253 26809 12265 26843
rect 12299 26840 12311 26843
rect 13004 26840 13032 26868
rect 12299 26812 13032 26840
rect 13188 26840 13216 26939
rect 13280 26917 13308 26948
rect 13832 26920 13860 26948
rect 14108 26948 14964 26976
rect 13265 26911 13323 26917
rect 13265 26877 13277 26911
rect 13311 26877 13323 26911
rect 13265 26871 13323 26877
rect 13725 26911 13783 26917
rect 13725 26877 13737 26911
rect 13771 26877 13783 26911
rect 13725 26871 13783 26877
rect 13354 26840 13360 26852
rect 13188 26812 13360 26840
rect 12299 26809 12311 26812
rect 12253 26803 12311 26809
rect 8987 26744 9352 26772
rect 9677 26775 9735 26781
rect 8987 26741 8999 26744
rect 8941 26735 8999 26741
rect 9677 26741 9689 26775
rect 9723 26772 9735 26775
rect 9861 26775 9919 26781
rect 9861 26772 9873 26775
rect 9723 26744 9873 26772
rect 9723 26741 9735 26744
rect 9677 26735 9735 26741
rect 9861 26741 9873 26744
rect 9907 26741 9919 26775
rect 9861 26735 9919 26741
rect 10226 26732 10232 26784
rect 10284 26732 10290 26784
rect 10704 26772 10732 26803
rect 13354 26800 13360 26812
rect 13412 26840 13418 26852
rect 13740 26840 13768 26871
rect 13814 26868 13820 26920
rect 13872 26868 13878 26920
rect 14108 26917 14136 26948
rect 14936 26920 14964 26948
rect 15212 26948 15700 26976
rect 14093 26911 14151 26917
rect 14093 26877 14105 26911
rect 14139 26877 14151 26911
rect 14093 26871 14151 26877
rect 14274 26868 14280 26920
rect 14332 26868 14338 26920
rect 14826 26908 14832 26920
rect 14476 26880 14832 26908
rect 13412 26812 13768 26840
rect 13909 26843 13967 26849
rect 13412 26800 13418 26812
rect 13909 26809 13921 26843
rect 13955 26840 13967 26843
rect 14476 26840 14504 26880
rect 14826 26868 14832 26880
rect 14884 26868 14890 26920
rect 14918 26868 14924 26920
rect 14976 26868 14982 26920
rect 15212 26917 15240 26948
rect 15672 26920 15700 26948
rect 16942 26936 16948 26988
rect 17000 26976 17006 26988
rect 17000 26948 17356 26976
rect 17000 26936 17006 26948
rect 15197 26911 15255 26917
rect 15197 26877 15209 26911
rect 15243 26877 15255 26911
rect 15197 26871 15255 26877
rect 15562 26868 15568 26920
rect 15620 26868 15626 26920
rect 15654 26868 15660 26920
rect 15712 26868 15718 26920
rect 15838 26868 15844 26920
rect 15896 26868 15902 26920
rect 15933 26911 15991 26917
rect 15933 26877 15945 26911
rect 15979 26908 15991 26911
rect 17126 26908 17132 26920
rect 15979 26880 17132 26908
rect 15979 26877 15991 26880
rect 15933 26871 15991 26877
rect 17126 26868 17132 26880
rect 17184 26868 17190 26920
rect 17221 26911 17279 26917
rect 17221 26877 17233 26911
rect 17267 26877 17279 26911
rect 17221 26871 17279 26877
rect 13955 26812 14504 26840
rect 14553 26843 14611 26849
rect 13955 26809 13967 26812
rect 13909 26803 13967 26809
rect 14553 26809 14565 26843
rect 14599 26840 14611 26843
rect 15381 26843 15439 26849
rect 15381 26840 15393 26843
rect 14599 26812 15393 26840
rect 14599 26809 14611 26812
rect 14553 26803 14611 26809
rect 15381 26809 15393 26812
rect 15427 26809 15439 26843
rect 15381 26803 15439 26809
rect 11146 26772 11152 26784
rect 10704 26744 11152 26772
rect 11146 26732 11152 26744
rect 11204 26732 11210 26784
rect 11241 26775 11299 26781
rect 11241 26741 11253 26775
rect 11287 26772 11299 26775
rect 11422 26772 11428 26784
rect 11287 26744 11428 26772
rect 11287 26741 11299 26744
rect 11241 26735 11299 26741
rect 11422 26732 11428 26744
rect 11480 26732 11486 26784
rect 11606 26732 11612 26784
rect 11664 26772 11670 26784
rect 12529 26775 12587 26781
rect 12529 26772 12541 26775
rect 11664 26744 12541 26772
rect 11664 26732 11670 26744
rect 12529 26741 12541 26744
rect 12575 26741 12587 26775
rect 12529 26735 12587 26741
rect 12710 26732 12716 26784
rect 12768 26732 12774 26784
rect 12986 26732 12992 26784
rect 13044 26772 13050 26784
rect 13541 26775 13599 26781
rect 13541 26772 13553 26775
rect 13044 26744 13553 26772
rect 13044 26732 13050 26744
rect 13541 26741 13553 26744
rect 13587 26741 13599 26775
rect 13541 26735 13599 26741
rect 14369 26775 14427 26781
rect 14369 26741 14381 26775
rect 14415 26772 14427 26775
rect 14645 26775 14703 26781
rect 14645 26772 14657 26775
rect 14415 26744 14657 26772
rect 14415 26741 14427 26744
rect 14369 26735 14427 26741
rect 14645 26741 14657 26744
rect 14691 26741 14703 26775
rect 14645 26735 14703 26741
rect 15654 26732 15660 26784
rect 15712 26772 15718 26784
rect 16758 26772 16764 26784
rect 15712 26744 16764 26772
rect 15712 26732 15718 26744
rect 16758 26732 16764 26744
rect 16816 26732 16822 26784
rect 17236 26772 17264 26871
rect 17328 26840 17356 26948
rect 17420 26917 17448 27016
rect 18322 27004 18328 27016
rect 18380 27004 18386 27056
rect 21637 27047 21695 27053
rect 20180 27016 21588 27044
rect 19797 26979 19855 26985
rect 19797 26976 19809 26979
rect 17972 26948 19809 26976
rect 17405 26911 17463 26917
rect 17405 26877 17417 26911
rect 17451 26877 17463 26911
rect 17405 26871 17463 26877
rect 17589 26911 17647 26917
rect 17589 26877 17601 26911
rect 17635 26908 17647 26911
rect 17770 26908 17776 26920
rect 17635 26880 17776 26908
rect 17635 26877 17647 26880
rect 17589 26871 17647 26877
rect 17770 26868 17776 26880
rect 17828 26868 17834 26920
rect 17972 26917 18000 26948
rect 19797 26945 19809 26948
rect 19843 26945 19855 26979
rect 19797 26939 19855 26945
rect 17957 26911 18015 26917
rect 17957 26877 17969 26911
rect 18003 26877 18015 26911
rect 17957 26871 18015 26877
rect 18138 26868 18144 26920
rect 18196 26868 18202 26920
rect 18325 26911 18383 26917
rect 18325 26877 18337 26911
rect 18371 26908 18383 26911
rect 18414 26908 18420 26920
rect 18371 26880 18420 26908
rect 18371 26877 18383 26880
rect 18325 26871 18383 26877
rect 18414 26868 18420 26880
rect 18472 26868 18478 26920
rect 19242 26868 19248 26920
rect 19300 26908 19306 26920
rect 19337 26911 19395 26917
rect 19337 26908 19349 26911
rect 19300 26880 19349 26908
rect 19300 26868 19306 26880
rect 19337 26877 19349 26880
rect 19383 26908 19395 26911
rect 20180 26908 20208 27016
rect 21266 26936 21272 26988
rect 21324 26936 21330 26988
rect 19383 26880 20208 26908
rect 20441 26911 20499 26917
rect 19383 26877 19395 26880
rect 19337 26871 19395 26877
rect 20441 26877 20453 26911
rect 20487 26877 20499 26911
rect 20441 26871 20499 26877
rect 17494 26840 17500 26852
rect 17328 26812 17500 26840
rect 17494 26800 17500 26812
rect 17552 26800 17558 26852
rect 18230 26800 18236 26852
rect 18288 26800 18294 26852
rect 18693 26775 18751 26781
rect 18693 26772 18705 26775
rect 17236 26744 18705 26772
rect 18693 26741 18705 26744
rect 18739 26741 18751 26775
rect 20456 26772 20484 26871
rect 20898 26868 20904 26920
rect 20956 26868 20962 26920
rect 21082 26868 21088 26920
rect 21140 26868 21146 26920
rect 21174 26868 21180 26920
rect 21232 26868 21238 26920
rect 21453 26911 21511 26917
rect 21453 26877 21465 26911
rect 21499 26877 21511 26911
rect 21560 26908 21588 27016
rect 21637 27013 21649 27047
rect 21683 27044 21695 27047
rect 22462 27044 22468 27056
rect 21683 27016 22468 27044
rect 21683 27013 21695 27016
rect 21637 27007 21695 27013
rect 22462 27004 22468 27016
rect 22520 27004 22526 27056
rect 21910 26936 21916 26988
rect 21968 26976 21974 26988
rect 22646 26976 22652 26988
rect 21968 26948 22652 26976
rect 21968 26936 21974 26948
rect 22646 26936 22652 26948
rect 22704 26936 22710 26988
rect 23860 26948 24532 26976
rect 22005 26911 22063 26917
rect 21560 26880 21956 26908
rect 21453 26871 21511 26877
rect 20993 26843 21051 26849
rect 20993 26809 21005 26843
rect 21039 26840 21051 26843
rect 21468 26840 21496 26871
rect 21818 26840 21824 26852
rect 21039 26812 21824 26840
rect 21039 26809 21051 26812
rect 20993 26803 21051 26809
rect 21818 26800 21824 26812
rect 21876 26800 21882 26852
rect 21928 26840 21956 26880
rect 22005 26877 22017 26911
rect 22051 26908 22063 26911
rect 22094 26908 22100 26920
rect 22051 26880 22100 26908
rect 22051 26877 22063 26880
rect 22005 26871 22063 26877
rect 22094 26868 22100 26880
rect 22152 26868 22158 26920
rect 22189 26911 22247 26917
rect 22189 26877 22201 26911
rect 22235 26908 22247 26911
rect 22830 26908 22836 26920
rect 22235 26880 22836 26908
rect 22235 26877 22247 26880
rect 22189 26871 22247 26877
rect 22204 26840 22232 26871
rect 22830 26868 22836 26880
rect 22888 26868 22894 26920
rect 23293 26911 23351 26917
rect 23293 26877 23305 26911
rect 23339 26877 23351 26911
rect 23293 26871 23351 26877
rect 21928 26812 22232 26840
rect 23308 26840 23336 26871
rect 23750 26868 23756 26920
rect 23808 26908 23814 26920
rect 23860 26917 23888 26948
rect 24504 26917 24532 26948
rect 23845 26911 23903 26917
rect 23845 26908 23857 26911
rect 23808 26880 23857 26908
rect 23808 26868 23814 26880
rect 23845 26877 23857 26880
rect 23891 26877 23903 26911
rect 23845 26871 23903 26877
rect 24397 26911 24455 26917
rect 24397 26877 24409 26911
rect 24443 26877 24455 26911
rect 24397 26871 24455 26877
rect 24489 26911 24547 26917
rect 24489 26877 24501 26911
rect 24535 26877 24547 26911
rect 24489 26871 24547 26877
rect 24673 26911 24731 26917
rect 24673 26877 24685 26911
rect 24719 26908 24731 26911
rect 24765 26911 24823 26917
rect 24765 26908 24777 26911
rect 24719 26880 24777 26908
rect 24719 26877 24731 26880
rect 24673 26871 24731 26877
rect 24765 26877 24777 26880
rect 24811 26908 24823 26911
rect 25038 26908 25044 26920
rect 24811 26880 25044 26908
rect 24811 26877 24823 26880
rect 24765 26871 24823 26877
rect 24026 26840 24032 26852
rect 23308 26812 24032 26840
rect 24026 26800 24032 26812
rect 24084 26840 24090 26852
rect 24412 26840 24440 26871
rect 25038 26868 25044 26880
rect 25096 26868 25102 26920
rect 25314 26868 25320 26920
rect 25372 26908 25378 26920
rect 25593 26911 25651 26917
rect 25593 26908 25605 26911
rect 25372 26880 25605 26908
rect 25372 26868 25378 26880
rect 25593 26877 25605 26880
rect 25639 26908 25651 26911
rect 26142 26908 26148 26920
rect 25639 26880 26148 26908
rect 25639 26877 25651 26880
rect 25593 26871 25651 26877
rect 26142 26868 26148 26880
rect 26200 26868 26206 26920
rect 25866 26849 25872 26852
rect 24084 26812 25728 26840
rect 24084 26800 24090 26812
rect 20714 26772 20720 26784
rect 20456 26744 20720 26772
rect 18693 26735 18751 26741
rect 20714 26732 20720 26744
rect 20772 26772 20778 26784
rect 21910 26772 21916 26784
rect 20772 26744 21916 26772
rect 20772 26732 20778 26744
rect 21910 26732 21916 26744
rect 21968 26732 21974 26784
rect 22094 26732 22100 26784
rect 22152 26772 22158 26784
rect 23014 26772 23020 26784
rect 22152 26744 23020 26772
rect 22152 26732 22158 26744
rect 23014 26732 23020 26744
rect 23072 26732 23078 26784
rect 25130 26732 25136 26784
rect 25188 26732 25194 26784
rect 25317 26775 25375 26781
rect 25317 26741 25329 26775
rect 25363 26772 25375 26775
rect 25590 26772 25596 26784
rect 25363 26744 25596 26772
rect 25363 26741 25375 26744
rect 25317 26735 25375 26741
rect 25590 26732 25596 26744
rect 25648 26732 25654 26784
rect 25700 26772 25728 26812
rect 25860 26803 25872 26849
rect 25866 26800 25872 26803
rect 25924 26800 25930 26852
rect 26973 26775 27031 26781
rect 26973 26772 26985 26775
rect 25700 26744 26985 26772
rect 26973 26741 26985 26744
rect 27019 26741 27031 26775
rect 26973 26735 27031 26741
rect 552 26682 27576 26704
rect 552 26630 7114 26682
rect 7166 26630 7178 26682
rect 7230 26630 7242 26682
rect 7294 26630 7306 26682
rect 7358 26630 7370 26682
rect 7422 26630 13830 26682
rect 13882 26630 13894 26682
rect 13946 26630 13958 26682
rect 14010 26630 14022 26682
rect 14074 26630 14086 26682
rect 14138 26630 20546 26682
rect 20598 26630 20610 26682
rect 20662 26630 20674 26682
rect 20726 26630 20738 26682
rect 20790 26630 20802 26682
rect 20854 26630 27262 26682
rect 27314 26630 27326 26682
rect 27378 26630 27390 26682
rect 27442 26630 27454 26682
rect 27506 26630 27518 26682
rect 27570 26630 27576 26682
rect 552 26608 27576 26630
rect 1118 26528 1124 26580
rect 1176 26528 1182 26580
rect 2222 26528 2228 26580
rect 2280 26568 2286 26580
rect 2280 26540 2728 26568
rect 2280 26528 2286 26540
rect 2700 26509 2728 26540
rect 2774 26528 2780 26580
rect 2832 26528 2838 26580
rect 5537 26571 5595 26577
rect 5537 26537 5549 26571
rect 5583 26568 5595 26571
rect 5626 26568 5632 26580
rect 5583 26540 5632 26568
rect 5583 26537 5595 26540
rect 5537 26531 5595 26537
rect 5626 26528 5632 26540
rect 5684 26528 5690 26580
rect 6178 26528 6184 26580
rect 6236 26568 6242 26580
rect 8021 26571 8079 26577
rect 8021 26568 8033 26571
rect 6236 26540 8033 26568
rect 6236 26528 6242 26540
rect 8021 26537 8033 26540
rect 8067 26568 8079 26571
rect 8110 26568 8116 26580
rect 8067 26540 8116 26568
rect 8067 26537 8079 26540
rect 8021 26531 8079 26537
rect 8110 26528 8116 26540
rect 8168 26528 8174 26580
rect 9585 26571 9643 26577
rect 9585 26568 9597 26571
rect 8404 26540 9597 26568
rect 8404 26509 8432 26540
rect 9585 26537 9597 26540
rect 9631 26537 9643 26571
rect 9585 26531 9643 26537
rect 11422 26528 11428 26580
rect 11480 26528 11486 26580
rect 13173 26571 13231 26577
rect 13173 26537 13185 26571
rect 13219 26568 13231 26571
rect 14274 26568 14280 26580
rect 13219 26540 14280 26568
rect 13219 26537 13231 26540
rect 13173 26531 13231 26537
rect 14274 26528 14280 26540
rect 14332 26528 14338 26580
rect 16574 26568 16580 26580
rect 15764 26540 16580 26568
rect 2485 26503 2543 26509
rect 2485 26469 2497 26503
rect 2531 26500 2543 26503
rect 2685 26503 2743 26509
rect 2531 26472 2636 26500
rect 2531 26469 2543 26472
rect 2485 26463 2543 26469
rect 1305 26435 1363 26441
rect 1305 26401 1317 26435
rect 1351 26432 1363 26435
rect 2314 26432 2320 26444
rect 1351 26404 2320 26432
rect 1351 26401 1363 26404
rect 1305 26395 1363 26401
rect 2314 26392 2320 26404
rect 2372 26392 2378 26444
rect 2608 26432 2636 26472
rect 2685 26469 2697 26503
rect 2731 26500 2743 26503
rect 2961 26503 3019 26509
rect 2961 26500 2973 26503
rect 2731 26472 2973 26500
rect 2731 26469 2743 26472
rect 2685 26463 2743 26469
rect 2961 26469 2973 26472
rect 3007 26500 3019 26503
rect 8389 26503 8447 26509
rect 3007 26472 3280 26500
rect 3007 26469 3019 26472
rect 2961 26463 3019 26469
rect 3050 26432 3056 26444
rect 2608 26404 3056 26432
rect 3050 26392 3056 26404
rect 3108 26392 3114 26444
rect 3142 26392 3148 26444
rect 3200 26392 3206 26444
rect 3252 26441 3280 26472
rect 8389 26469 8401 26503
rect 8435 26469 8447 26503
rect 8605 26503 8663 26509
rect 8605 26500 8617 26503
rect 8389 26463 8447 26469
rect 8496 26472 8617 26500
rect 3237 26435 3295 26441
rect 3237 26401 3249 26435
rect 3283 26401 3295 26435
rect 3237 26395 3295 26401
rect 3329 26435 3387 26441
rect 3329 26401 3341 26435
rect 3375 26432 3387 26435
rect 4338 26432 4344 26444
rect 3375 26404 4344 26432
rect 3375 26401 3387 26404
rect 3329 26395 3387 26401
rect 4338 26392 4344 26404
rect 4396 26392 4402 26444
rect 5353 26435 5411 26441
rect 5353 26401 5365 26435
rect 5399 26432 5411 26435
rect 5442 26432 5448 26444
rect 5399 26404 5448 26432
rect 5399 26401 5411 26404
rect 5353 26395 5411 26401
rect 5442 26392 5448 26404
rect 5500 26392 5506 26444
rect 5629 26435 5687 26441
rect 5629 26401 5641 26435
rect 5675 26432 5687 26435
rect 5810 26432 5816 26444
rect 5675 26404 5816 26432
rect 5675 26401 5687 26404
rect 5629 26395 5687 26401
rect 5810 26392 5816 26404
rect 5868 26392 5874 26444
rect 5905 26435 5963 26441
rect 5905 26401 5917 26435
rect 5951 26401 5963 26435
rect 5905 26395 5963 26401
rect 3510 26324 3516 26376
rect 3568 26364 3574 26376
rect 3973 26367 4031 26373
rect 3973 26364 3985 26367
rect 3568 26336 3985 26364
rect 3568 26324 3574 26336
rect 3973 26333 3985 26336
rect 4019 26333 4031 26367
rect 5460 26364 5488 26392
rect 5920 26364 5948 26395
rect 6086 26392 6092 26444
rect 6144 26392 6150 26444
rect 6178 26392 6184 26444
rect 6236 26392 6242 26444
rect 6454 26392 6460 26444
rect 6512 26432 6518 26444
rect 6641 26435 6699 26441
rect 6641 26432 6653 26435
rect 6512 26404 6653 26432
rect 6512 26392 6518 26404
rect 6641 26401 6653 26404
rect 6687 26401 6699 26435
rect 6897 26435 6955 26441
rect 6897 26432 6909 26435
rect 6641 26395 6699 26401
rect 6748 26404 6909 26432
rect 6748 26364 6776 26404
rect 6897 26401 6909 26404
rect 6943 26401 6955 26435
rect 6897 26395 6955 26401
rect 8294 26392 8300 26444
rect 8352 26432 8358 26444
rect 8496 26432 8524 26472
rect 8605 26469 8617 26472
rect 8651 26500 8663 26503
rect 9950 26500 9956 26512
rect 8651 26472 9956 26500
rect 8651 26469 8663 26472
rect 8605 26463 8663 26469
rect 9950 26460 9956 26472
rect 10008 26500 10014 26512
rect 10565 26503 10623 26509
rect 10565 26500 10577 26503
rect 10008 26472 10577 26500
rect 10008 26460 10014 26472
rect 10565 26469 10577 26472
rect 10611 26469 10623 26503
rect 10565 26463 10623 26469
rect 10781 26503 10839 26509
rect 10781 26469 10793 26503
rect 10827 26500 10839 26503
rect 11698 26500 11704 26512
rect 10827 26472 11704 26500
rect 10827 26469 10839 26472
rect 10781 26463 10839 26469
rect 11698 26460 11704 26472
rect 11756 26460 11762 26512
rect 11793 26503 11851 26509
rect 11793 26469 11805 26503
rect 11839 26500 11851 26503
rect 12805 26503 12863 26509
rect 12805 26500 12817 26503
rect 11839 26472 12817 26500
rect 11839 26469 11851 26472
rect 11793 26463 11851 26469
rect 12805 26469 12817 26472
rect 12851 26469 12863 26503
rect 12805 26463 12863 26469
rect 9033 26435 9091 26441
rect 9033 26432 9045 26435
rect 8352 26404 8524 26432
rect 8772 26404 9045 26432
rect 8352 26392 8358 26404
rect 5460 26336 5948 26364
rect 6656 26336 6776 26364
rect 3973 26327 4031 26333
rect 2317 26299 2375 26305
rect 2317 26265 2329 26299
rect 2363 26296 2375 26299
rect 2406 26296 2412 26308
rect 2363 26268 2412 26296
rect 2363 26265 2375 26268
rect 2317 26259 2375 26265
rect 2406 26256 2412 26268
rect 2464 26256 2470 26308
rect 3326 26296 3332 26308
rect 2746 26268 3332 26296
rect 2501 26231 2559 26237
rect 2501 26197 2513 26231
rect 2547 26228 2559 26231
rect 2746 26228 2774 26268
rect 3326 26256 3332 26268
rect 3384 26296 3390 26308
rect 4154 26296 4160 26308
rect 3384 26268 4160 26296
rect 3384 26256 3390 26268
rect 4154 26256 4160 26268
rect 4212 26296 4218 26308
rect 4249 26299 4307 26305
rect 4249 26296 4261 26299
rect 4212 26268 4261 26296
rect 4212 26256 4218 26268
rect 4249 26265 4261 26268
rect 4295 26265 4307 26299
rect 4249 26259 4307 26265
rect 6362 26256 6368 26308
rect 6420 26256 6426 26308
rect 2547 26200 2774 26228
rect 4433 26231 4491 26237
rect 2547 26197 2559 26200
rect 2501 26191 2559 26197
rect 4433 26197 4445 26231
rect 4479 26228 4491 26231
rect 4614 26228 4620 26240
rect 4479 26200 4620 26228
rect 4479 26197 4491 26200
rect 4433 26191 4491 26197
rect 4614 26188 4620 26200
rect 4672 26188 4678 26240
rect 4982 26188 4988 26240
rect 5040 26228 5046 26240
rect 5169 26231 5227 26237
rect 5169 26228 5181 26231
rect 5040 26200 5181 26228
rect 5040 26188 5046 26200
rect 5169 26197 5181 26200
rect 5215 26197 5227 26231
rect 6656 26228 6684 26336
rect 8772 26305 8800 26404
rect 9033 26401 9045 26404
rect 9079 26401 9091 26435
rect 9033 26395 9091 26401
rect 9214 26392 9220 26444
rect 9272 26392 9278 26444
rect 9309 26435 9367 26441
rect 9309 26401 9321 26435
rect 9355 26432 9367 26435
rect 9582 26432 9588 26444
rect 9355 26404 9588 26432
rect 9355 26401 9367 26404
rect 9309 26395 9367 26401
rect 9582 26392 9588 26404
rect 9640 26392 9646 26444
rect 10042 26392 10048 26444
rect 10100 26432 10106 26444
rect 10137 26435 10195 26441
rect 10137 26432 10149 26435
rect 10100 26404 10149 26432
rect 10100 26392 10106 26404
rect 10137 26401 10149 26404
rect 10183 26401 10195 26435
rect 10137 26395 10195 26401
rect 10226 26392 10232 26444
rect 10284 26432 10290 26444
rect 11333 26435 11391 26441
rect 11333 26432 11345 26435
rect 10284 26404 11345 26432
rect 10284 26392 10290 26404
rect 11333 26401 11345 26404
rect 11379 26401 11391 26435
rect 11333 26395 11391 26401
rect 11606 26392 11612 26444
rect 11664 26392 11670 26444
rect 12066 26392 12072 26444
rect 12124 26392 12130 26444
rect 12253 26435 12311 26441
rect 12253 26401 12265 26435
rect 12299 26401 12311 26435
rect 12253 26395 12311 26401
rect 12345 26435 12403 26441
rect 12345 26401 12357 26435
rect 12391 26432 12403 26435
rect 12434 26432 12440 26444
rect 12391 26404 12440 26432
rect 12391 26401 12403 26404
rect 12345 26395 12403 26401
rect 11422 26324 11428 26376
rect 11480 26364 11486 26376
rect 12268 26364 12296 26395
rect 12434 26392 12440 26404
rect 12492 26392 12498 26444
rect 12710 26392 12716 26444
rect 12768 26392 12774 26444
rect 12986 26392 12992 26444
rect 13044 26392 13050 26444
rect 14734 26432 14740 26444
rect 13648 26404 14740 26432
rect 13648 26364 13676 26404
rect 14734 26392 14740 26404
rect 14792 26392 14798 26444
rect 15654 26392 15660 26444
rect 15712 26392 15718 26444
rect 15764 26441 15792 26540
rect 16574 26528 16580 26540
rect 16632 26528 16638 26580
rect 16666 26528 16672 26580
rect 16724 26568 16730 26580
rect 21634 26568 21640 26580
rect 16724 26540 21640 26568
rect 16724 26528 16730 26540
rect 21634 26528 21640 26540
rect 21692 26568 21698 26580
rect 22554 26568 22560 26580
rect 21692 26540 22560 26568
rect 21692 26528 21698 26540
rect 22554 26528 22560 26540
rect 22612 26528 22618 26580
rect 23750 26528 23756 26580
rect 23808 26568 23814 26580
rect 24003 26571 24061 26577
rect 24003 26568 24015 26571
rect 23808 26540 24015 26568
rect 23808 26528 23814 26540
rect 24003 26537 24015 26540
rect 24049 26537 24061 26571
rect 24003 26531 24061 26537
rect 25777 26571 25835 26577
rect 25777 26537 25789 26571
rect 25823 26568 25835 26571
rect 25866 26568 25872 26580
rect 25823 26540 25872 26568
rect 25823 26537 25835 26540
rect 25777 26531 25835 26537
rect 25866 26528 25872 26540
rect 25924 26528 25930 26580
rect 15933 26503 15991 26509
rect 15933 26469 15945 26503
rect 15979 26500 15991 26503
rect 19613 26503 19671 26509
rect 19613 26500 19625 26503
rect 15979 26472 16160 26500
rect 15979 26469 15991 26472
rect 15933 26463 15991 26469
rect 16132 26441 16160 26472
rect 18064 26472 19625 26500
rect 15749 26435 15807 26441
rect 15749 26401 15761 26435
rect 15795 26401 15807 26435
rect 15749 26395 15807 26401
rect 16117 26435 16175 26441
rect 16117 26401 16129 26435
rect 16163 26401 16175 26435
rect 16117 26395 16175 26401
rect 16298 26392 16304 26444
rect 16356 26392 16362 26444
rect 16666 26392 16672 26444
rect 16724 26392 16730 26444
rect 17313 26435 17371 26441
rect 17313 26401 17325 26435
rect 17359 26432 17371 26435
rect 17773 26435 17831 26441
rect 17773 26432 17785 26435
rect 17359 26404 17785 26432
rect 17359 26401 17371 26404
rect 17313 26395 17371 26401
rect 17773 26401 17785 26404
rect 17819 26432 17831 26435
rect 17862 26432 17868 26444
rect 17819 26404 17868 26432
rect 17819 26401 17831 26404
rect 17773 26395 17831 26401
rect 17862 26392 17868 26404
rect 17920 26392 17926 26444
rect 18064 26441 18092 26472
rect 19613 26469 19625 26472
rect 19659 26469 19671 26503
rect 19613 26463 19671 26469
rect 20441 26503 20499 26509
rect 20441 26469 20453 26503
rect 20487 26500 20499 26503
rect 21082 26500 21088 26512
rect 20487 26472 21088 26500
rect 20487 26469 20499 26472
rect 20441 26463 20499 26469
rect 21082 26460 21088 26472
rect 21140 26500 21146 26512
rect 21269 26503 21327 26509
rect 21269 26500 21281 26503
rect 21140 26472 21281 26500
rect 21140 26460 21146 26472
rect 21269 26469 21281 26472
rect 21315 26469 21327 26503
rect 24213 26503 24271 26509
rect 24213 26500 24225 26503
rect 21269 26463 21327 26469
rect 21376 26472 24225 26500
rect 18049 26435 18107 26441
rect 18049 26401 18061 26435
rect 18095 26401 18107 26435
rect 18049 26395 18107 26401
rect 18230 26392 18236 26444
rect 18288 26392 18294 26444
rect 18325 26435 18383 26441
rect 18325 26401 18337 26435
rect 18371 26401 18383 26435
rect 18325 26395 18383 26401
rect 11480 26336 13676 26364
rect 15933 26367 15991 26373
rect 11480 26324 11486 26336
rect 15933 26333 15945 26367
rect 15979 26364 15991 26367
rect 15979 26336 16804 26364
rect 15979 26333 15991 26336
rect 15933 26327 15991 26333
rect 8757 26299 8815 26305
rect 8757 26265 8769 26299
rect 8803 26265 8815 26299
rect 8757 26259 8815 26265
rect 10226 26256 10232 26308
rect 10284 26296 10290 26308
rect 10502 26296 10508 26308
rect 10284 26268 10508 26296
rect 10284 26256 10290 26268
rect 10502 26256 10508 26268
rect 10560 26256 10566 26308
rect 16022 26256 16028 26308
rect 16080 26296 16086 26308
rect 16776 26305 16804 26336
rect 16942 26324 16948 26376
rect 17000 26364 17006 26376
rect 17037 26367 17095 26373
rect 17037 26364 17049 26367
rect 17000 26336 17049 26364
rect 17000 26324 17006 26336
rect 17037 26333 17049 26336
rect 17083 26364 17095 26367
rect 17681 26367 17739 26373
rect 17681 26364 17693 26367
rect 17083 26336 17693 26364
rect 17083 26333 17095 26336
rect 17037 26327 17095 26333
rect 17681 26333 17693 26336
rect 17727 26333 17739 26367
rect 17681 26327 17739 26333
rect 17954 26324 17960 26376
rect 18012 26364 18018 26376
rect 18340 26364 18368 26395
rect 18414 26392 18420 26444
rect 18472 26392 18478 26444
rect 20622 26392 20628 26444
rect 20680 26392 20686 26444
rect 20717 26435 20775 26441
rect 20717 26401 20729 26435
rect 20763 26401 20775 26435
rect 20717 26395 20775 26401
rect 18012 26336 18828 26364
rect 18012 26324 18018 26336
rect 16301 26299 16359 26305
rect 16301 26296 16313 26299
rect 16080 26268 16313 26296
rect 16080 26256 16086 26268
rect 16301 26265 16313 26268
rect 16347 26265 16359 26299
rect 16301 26259 16359 26265
rect 16761 26299 16819 26305
rect 16761 26265 16773 26299
rect 16807 26265 16819 26299
rect 16761 26259 16819 26265
rect 17126 26256 17132 26308
rect 17184 26296 17190 26308
rect 17405 26299 17463 26305
rect 17405 26296 17417 26299
rect 17184 26268 17417 26296
rect 17184 26256 17190 26268
rect 17405 26265 17417 26268
rect 17451 26265 17463 26299
rect 17405 26259 17463 26265
rect 18230 26256 18236 26308
rect 18288 26296 18294 26308
rect 18693 26299 18751 26305
rect 18693 26296 18705 26299
rect 18288 26268 18705 26296
rect 18288 26256 18294 26268
rect 18693 26265 18705 26268
rect 18739 26265 18751 26299
rect 18800 26296 18828 26336
rect 19334 26324 19340 26376
rect 19392 26324 19398 26376
rect 20257 26367 20315 26373
rect 20257 26333 20269 26367
rect 20303 26364 20315 26367
rect 20346 26364 20352 26376
rect 20303 26336 20352 26364
rect 20303 26333 20315 26336
rect 20257 26327 20315 26333
rect 20346 26324 20352 26336
rect 20404 26324 20410 26376
rect 20732 26364 20760 26395
rect 20990 26392 20996 26444
rect 21048 26392 21054 26444
rect 21376 26364 21404 26472
rect 24213 26469 24225 26472
rect 24259 26500 24271 26503
rect 24857 26503 24915 26509
rect 24857 26500 24869 26503
rect 24259 26472 24869 26500
rect 24259 26469 24271 26472
rect 24213 26463 24271 26469
rect 24857 26469 24869 26472
rect 24903 26500 24915 26503
rect 24903 26472 24992 26500
rect 24903 26469 24915 26472
rect 24857 26463 24915 26469
rect 21542 26392 21548 26444
rect 21600 26392 21606 26444
rect 21818 26392 21824 26444
rect 21876 26392 21882 26444
rect 23109 26435 23167 26441
rect 23109 26401 23121 26435
rect 23155 26432 23167 26435
rect 23750 26432 23756 26444
rect 23155 26404 23756 26432
rect 23155 26401 23167 26404
rect 23109 26395 23167 26401
rect 23750 26392 23756 26404
rect 23808 26392 23814 26444
rect 20732 26336 21404 26364
rect 19702 26296 19708 26308
rect 18800 26268 19708 26296
rect 18693 26259 18751 26265
rect 19702 26256 19708 26268
rect 19760 26256 19766 26308
rect 6822 26228 6828 26240
rect 6656 26200 6828 26228
rect 5169 26191 5227 26197
rect 6822 26188 6828 26200
rect 6880 26188 6886 26240
rect 8570 26188 8576 26240
rect 8628 26188 8634 26240
rect 8662 26188 8668 26240
rect 8720 26228 8726 26240
rect 8849 26231 8907 26237
rect 8849 26228 8861 26231
rect 8720 26200 8861 26228
rect 8720 26188 8726 26200
rect 8849 26197 8861 26200
rect 8895 26197 8907 26231
rect 8849 26191 8907 26197
rect 9674 26188 9680 26240
rect 9732 26228 9738 26240
rect 10413 26231 10471 26237
rect 10413 26228 10425 26231
rect 9732 26200 10425 26228
rect 9732 26188 9738 26200
rect 10413 26197 10425 26200
rect 10459 26197 10471 26231
rect 10413 26191 10471 26197
rect 10597 26231 10655 26237
rect 10597 26197 10609 26231
rect 10643 26228 10655 26231
rect 10962 26228 10968 26240
rect 10643 26200 10968 26228
rect 10643 26197 10655 26200
rect 10597 26191 10655 26197
rect 10962 26188 10968 26200
rect 11020 26188 11026 26240
rect 11882 26188 11888 26240
rect 11940 26188 11946 26240
rect 16390 26188 16396 26240
rect 16448 26228 16454 26240
rect 16945 26231 17003 26237
rect 16945 26228 16957 26231
rect 16448 26200 16957 26228
rect 16448 26188 16454 26200
rect 16945 26197 16957 26200
rect 16991 26197 17003 26231
rect 16945 26191 17003 26197
rect 18598 26188 18604 26240
rect 18656 26188 18662 26240
rect 20162 26188 20168 26240
rect 20220 26228 20226 26240
rect 20732 26228 20760 26336
rect 21450 26324 21456 26376
rect 21508 26324 21514 26376
rect 22278 26364 22284 26376
rect 21560 26336 22284 26364
rect 21361 26299 21419 26305
rect 21361 26265 21373 26299
rect 21407 26296 21419 26299
rect 21560 26296 21588 26336
rect 22278 26324 22284 26336
rect 22336 26324 22342 26376
rect 24964 26364 24992 26472
rect 25038 26460 25044 26512
rect 25096 26460 25102 26512
rect 25590 26392 25596 26444
rect 25648 26392 25654 26444
rect 25038 26364 25044 26376
rect 24964 26336 25044 26364
rect 25038 26324 25044 26336
rect 25096 26324 25102 26376
rect 21407 26268 21588 26296
rect 21637 26299 21695 26305
rect 21407 26265 21419 26268
rect 21361 26259 21419 26265
rect 21637 26265 21649 26299
rect 21683 26296 21695 26299
rect 22186 26296 22192 26308
rect 21683 26268 22192 26296
rect 21683 26265 21695 26268
rect 21637 26259 21695 26265
rect 22186 26256 22192 26268
rect 22244 26256 22250 26308
rect 23845 26299 23903 26305
rect 23845 26265 23857 26299
rect 23891 26296 23903 26299
rect 24302 26296 24308 26308
rect 23891 26268 24308 26296
rect 23891 26265 23903 26268
rect 23845 26259 23903 26265
rect 24302 26256 24308 26268
rect 24360 26256 24366 26308
rect 20220 26200 20760 26228
rect 20220 26188 20226 26200
rect 20898 26188 20904 26240
rect 20956 26188 20962 26240
rect 23293 26231 23351 26237
rect 23293 26197 23305 26231
rect 23339 26228 23351 26231
rect 23382 26228 23388 26240
rect 23339 26200 23388 26228
rect 23339 26197 23351 26200
rect 23293 26191 23351 26197
rect 23382 26188 23388 26200
rect 23440 26188 23446 26240
rect 24026 26188 24032 26240
rect 24084 26188 24090 26240
rect 24670 26188 24676 26240
rect 24728 26188 24734 26240
rect 552 26138 27416 26160
rect 552 26086 3756 26138
rect 3808 26086 3820 26138
rect 3872 26086 3884 26138
rect 3936 26086 3948 26138
rect 4000 26086 4012 26138
rect 4064 26086 10472 26138
rect 10524 26086 10536 26138
rect 10588 26086 10600 26138
rect 10652 26086 10664 26138
rect 10716 26086 10728 26138
rect 10780 26086 17188 26138
rect 17240 26086 17252 26138
rect 17304 26086 17316 26138
rect 17368 26086 17380 26138
rect 17432 26086 17444 26138
rect 17496 26086 23904 26138
rect 23956 26086 23968 26138
rect 24020 26086 24032 26138
rect 24084 26086 24096 26138
rect 24148 26086 24160 26138
rect 24212 26086 27416 26138
rect 552 26064 27416 26086
rect 7006 25984 7012 26036
rect 7064 25984 7070 26036
rect 8021 26027 8079 26033
rect 8021 25993 8033 26027
rect 8067 26024 8079 26027
rect 8570 26024 8576 26036
rect 8067 25996 8576 26024
rect 8067 25993 8079 25996
rect 8021 25987 8079 25993
rect 8570 25984 8576 25996
rect 8628 26024 8634 26036
rect 8628 25996 9720 26024
rect 8628 25984 8634 25996
rect 2774 25956 2780 25968
rect 2332 25928 2780 25956
rect 2332 25829 2360 25928
rect 2774 25916 2780 25928
rect 2832 25916 2838 25968
rect 9692 25956 9720 25996
rect 9766 25984 9772 26036
rect 9824 26024 9830 26036
rect 9953 26027 10011 26033
rect 9953 26024 9965 26027
rect 9824 25996 9965 26024
rect 9824 25984 9830 25996
rect 9953 25993 9965 25996
rect 9999 25993 10011 26027
rect 9953 25987 10011 25993
rect 10226 25984 10232 26036
rect 10284 26024 10290 26036
rect 10413 26027 10471 26033
rect 10413 26024 10425 26027
rect 10284 25996 10425 26024
rect 10284 25984 10290 25996
rect 10413 25993 10425 25996
rect 10459 25993 10471 26027
rect 10413 25987 10471 25993
rect 11698 25984 11704 26036
rect 11756 26024 11762 26036
rect 11885 26027 11943 26033
rect 11885 26024 11897 26027
rect 11756 25996 11897 26024
rect 11756 25984 11762 25996
rect 11885 25993 11897 25996
rect 11931 25993 11943 26027
rect 11885 25987 11943 25993
rect 12406 25996 14780 26024
rect 10962 25956 10968 25968
rect 9692 25928 10968 25956
rect 10962 25916 10968 25928
rect 11020 25916 11026 25968
rect 11054 25916 11060 25968
rect 11112 25956 11118 25968
rect 12406 25956 12434 25996
rect 11112 25928 12434 25956
rect 14752 25956 14780 25996
rect 14826 25984 14832 26036
rect 14884 26024 14890 26036
rect 14921 26027 14979 26033
rect 14921 26024 14933 26027
rect 14884 25996 14933 26024
rect 14884 25984 14890 25996
rect 14921 25993 14933 25996
rect 14967 25993 14979 26027
rect 14921 25987 14979 25993
rect 15838 25984 15844 26036
rect 15896 26024 15902 26036
rect 16390 26024 16396 26036
rect 15896 25996 16396 26024
rect 15896 25984 15902 25996
rect 16390 25984 16396 25996
rect 16448 25984 16454 26036
rect 20441 26027 20499 26033
rect 20441 25993 20453 26027
rect 20487 26024 20499 26027
rect 20806 26024 20812 26036
rect 20487 25996 20812 26024
rect 20487 25993 20499 25996
rect 20441 25987 20499 25993
rect 20806 25984 20812 25996
rect 20864 25984 20870 26036
rect 20990 25984 20996 26036
rect 21048 26024 21054 26036
rect 22002 26024 22008 26036
rect 21048 25996 22008 26024
rect 21048 25984 21054 25996
rect 22002 25984 22008 25996
rect 22060 26024 22066 26036
rect 22281 26027 22339 26033
rect 22281 26024 22293 26027
rect 22060 25996 22293 26024
rect 22060 25984 22066 25996
rect 22281 25993 22293 25996
rect 22327 25993 22339 26027
rect 22281 25987 22339 25993
rect 23750 25984 23756 26036
rect 23808 26024 23814 26036
rect 23845 26027 23903 26033
rect 23845 26024 23857 26027
rect 23808 25996 23857 26024
rect 23808 25984 23814 25996
rect 23845 25993 23857 25996
rect 23891 25993 23903 26027
rect 23845 25987 23903 25993
rect 24026 25984 24032 26036
rect 24084 25984 24090 26036
rect 24670 25984 24676 26036
rect 24728 25984 24734 26036
rect 24949 26027 25007 26033
rect 24949 25993 24961 26027
rect 24995 26024 25007 26027
rect 25038 26024 25044 26036
rect 24995 25996 25044 26024
rect 24995 25993 25007 25996
rect 24949 25987 25007 25993
rect 25038 25984 25044 25996
rect 25096 25984 25102 26036
rect 16666 25956 16672 25968
rect 14752 25928 16672 25956
rect 11112 25916 11118 25928
rect 16666 25916 16672 25928
rect 16724 25916 16730 25968
rect 20717 25959 20775 25965
rect 20717 25925 20729 25959
rect 20763 25956 20775 25959
rect 21450 25956 21456 25968
rect 20763 25928 21456 25956
rect 20763 25925 20775 25928
rect 20717 25919 20775 25925
rect 2406 25848 2412 25900
rect 2464 25888 2470 25900
rect 2464 25860 2636 25888
rect 2464 25848 2470 25860
rect 2608 25829 2636 25860
rect 2682 25848 2688 25900
rect 2740 25848 2746 25900
rect 4982 25848 4988 25900
rect 5040 25848 5046 25900
rect 6914 25848 6920 25900
rect 6972 25888 6978 25900
rect 6972 25860 7420 25888
rect 6972 25848 6978 25860
rect 2317 25823 2375 25829
rect 2317 25789 2329 25823
rect 2363 25789 2375 25823
rect 2317 25783 2375 25789
rect 2501 25823 2559 25829
rect 2501 25789 2513 25823
rect 2547 25789 2559 25823
rect 2501 25783 2559 25789
rect 2593 25823 2651 25829
rect 2593 25789 2605 25823
rect 2639 25789 2651 25823
rect 2700 25820 2728 25848
rect 2777 25823 2835 25829
rect 2777 25820 2789 25823
rect 2700 25792 2789 25820
rect 2593 25783 2651 25789
rect 2777 25789 2789 25792
rect 2823 25789 2835 25823
rect 2777 25783 2835 25789
rect 2516 25752 2544 25783
rect 2866 25780 2872 25832
rect 2924 25780 2930 25832
rect 4430 25780 4436 25832
rect 4488 25820 4494 25832
rect 4893 25823 4951 25829
rect 4893 25820 4905 25823
rect 4488 25792 4905 25820
rect 4488 25780 4494 25792
rect 4893 25789 4905 25792
rect 4939 25789 4951 25823
rect 4893 25783 4951 25789
rect 5074 25780 5080 25832
rect 5132 25780 5138 25832
rect 5166 25780 5172 25832
rect 5224 25780 5230 25832
rect 6270 25780 6276 25832
rect 6328 25820 6334 25832
rect 7006 25820 7012 25832
rect 6328 25792 7012 25820
rect 6328 25780 6334 25792
rect 7006 25780 7012 25792
rect 7064 25820 7070 25832
rect 7392 25829 7420 25860
rect 9398 25848 9404 25900
rect 9456 25888 9462 25900
rect 10870 25888 10876 25900
rect 9456 25860 10272 25888
rect 9456 25848 9462 25860
rect 7193 25823 7251 25829
rect 7193 25820 7205 25823
rect 7064 25792 7205 25820
rect 7064 25780 7070 25792
rect 7193 25789 7205 25792
rect 7239 25789 7251 25823
rect 7193 25783 7251 25789
rect 7377 25823 7435 25829
rect 7377 25789 7389 25823
rect 7423 25789 7435 25823
rect 7377 25783 7435 25789
rect 7466 25780 7472 25832
rect 7524 25820 7530 25832
rect 7561 25823 7619 25829
rect 7561 25820 7573 25823
rect 7524 25792 7573 25820
rect 7524 25780 7530 25792
rect 7561 25789 7573 25792
rect 7607 25789 7619 25823
rect 8294 25820 8300 25832
rect 7561 25783 7619 25789
rect 8036 25792 8300 25820
rect 2685 25755 2743 25761
rect 2685 25752 2697 25755
rect 2516 25724 2697 25752
rect 2608 25696 2636 25724
rect 2685 25721 2697 25724
rect 2731 25721 2743 25755
rect 2685 25715 2743 25721
rect 3234 25712 3240 25764
rect 3292 25712 3298 25764
rect 3602 25712 3608 25764
rect 3660 25752 3666 25764
rect 3973 25755 4031 25761
rect 3973 25752 3985 25755
rect 3660 25724 3985 25752
rect 3660 25712 3666 25724
rect 3973 25721 3985 25724
rect 4019 25721 4031 25755
rect 3973 25715 4031 25721
rect 7285 25755 7343 25761
rect 7285 25721 7297 25755
rect 7331 25721 7343 25755
rect 7285 25715 7343 25721
rect 1854 25644 1860 25696
rect 1912 25684 1918 25696
rect 2317 25687 2375 25693
rect 2317 25684 2329 25687
rect 1912 25656 2329 25684
rect 1912 25644 1918 25656
rect 2317 25653 2329 25656
rect 2363 25653 2375 25687
rect 2317 25647 2375 25653
rect 2590 25644 2596 25696
rect 2648 25644 2654 25696
rect 3050 25644 3056 25696
rect 3108 25644 3114 25696
rect 4246 25644 4252 25696
rect 4304 25684 4310 25696
rect 4709 25687 4767 25693
rect 4709 25684 4721 25687
rect 4304 25656 4721 25684
rect 4304 25644 4310 25656
rect 4709 25653 4721 25656
rect 4755 25653 4767 25687
rect 7300 25684 7328 25715
rect 7834 25712 7840 25764
rect 7892 25712 7898 25764
rect 8036 25761 8064 25792
rect 8294 25780 8300 25792
rect 8352 25780 8358 25832
rect 8386 25780 8392 25832
rect 8444 25780 8450 25832
rect 8662 25829 8668 25832
rect 8656 25820 8668 25829
rect 8623 25792 8668 25820
rect 8656 25783 8668 25792
rect 8662 25780 8668 25783
rect 8720 25780 8726 25832
rect 10134 25780 10140 25832
rect 10192 25780 10198 25832
rect 10244 25829 10272 25860
rect 10520 25860 10876 25888
rect 10520 25829 10548 25860
rect 10870 25848 10876 25860
rect 10928 25848 10934 25900
rect 11146 25848 11152 25900
rect 11204 25888 11210 25900
rect 11701 25891 11759 25897
rect 11701 25888 11713 25891
rect 11204 25860 11713 25888
rect 11204 25848 11210 25860
rect 11701 25857 11713 25860
rect 11747 25888 11759 25891
rect 12618 25888 12624 25900
rect 11747 25860 12624 25888
rect 11747 25857 11759 25860
rect 11701 25851 11759 25857
rect 12618 25848 12624 25860
rect 12676 25888 12682 25900
rect 13541 25891 13599 25897
rect 13541 25888 13553 25891
rect 12676 25860 13553 25888
rect 12676 25848 12682 25860
rect 13541 25857 13553 25860
rect 13587 25857 13599 25891
rect 13541 25851 13599 25857
rect 14826 25848 14832 25900
rect 14884 25888 14890 25900
rect 15381 25891 15439 25897
rect 15381 25888 15393 25891
rect 14884 25860 15393 25888
rect 14884 25848 14890 25860
rect 15381 25857 15393 25860
rect 15427 25857 15439 25891
rect 15381 25851 15439 25857
rect 15746 25848 15752 25900
rect 15804 25888 15810 25900
rect 15841 25891 15899 25897
rect 15841 25888 15853 25891
rect 15804 25860 15853 25888
rect 15804 25848 15810 25860
rect 15841 25857 15853 25860
rect 15887 25857 15899 25891
rect 15841 25851 15899 25857
rect 16758 25848 16764 25900
rect 16816 25848 16822 25900
rect 18414 25888 18420 25900
rect 17880 25860 18420 25888
rect 17880 25832 17908 25860
rect 18414 25848 18420 25860
rect 18472 25848 18478 25900
rect 18690 25848 18696 25900
rect 18748 25848 18754 25900
rect 10229 25823 10287 25829
rect 10229 25789 10241 25823
rect 10275 25789 10287 25823
rect 10229 25783 10287 25789
rect 10505 25823 10563 25829
rect 10505 25789 10517 25823
rect 10551 25789 10563 25823
rect 10505 25783 10563 25789
rect 11238 25780 11244 25832
rect 11296 25820 11302 25832
rect 12437 25823 12495 25829
rect 12437 25820 12449 25823
rect 11296 25792 12449 25820
rect 11296 25780 11302 25792
rect 12437 25789 12449 25792
rect 12483 25789 12495 25823
rect 12437 25783 12495 25789
rect 12802 25780 12808 25832
rect 12860 25780 12866 25832
rect 15197 25823 15255 25829
rect 15197 25789 15209 25823
rect 15243 25820 15255 25823
rect 15470 25820 15476 25832
rect 15243 25792 15476 25820
rect 15243 25789 15255 25792
rect 15197 25783 15255 25789
rect 15470 25780 15476 25792
rect 15528 25780 15534 25832
rect 15657 25823 15715 25829
rect 15657 25789 15669 25823
rect 15703 25820 15715 25823
rect 16022 25820 16028 25832
rect 15703 25792 16028 25820
rect 15703 25789 15715 25792
rect 15657 25783 15715 25789
rect 16022 25780 16028 25792
rect 16080 25780 16086 25832
rect 16574 25780 16580 25832
rect 16632 25780 16638 25832
rect 17862 25780 17868 25832
rect 17920 25780 17926 25832
rect 18049 25823 18107 25829
rect 18049 25789 18061 25823
rect 18095 25820 18107 25823
rect 18138 25820 18144 25832
rect 18095 25792 18144 25820
rect 18095 25789 18107 25792
rect 18049 25783 18107 25789
rect 18138 25780 18144 25792
rect 18196 25780 18202 25832
rect 18230 25780 18236 25832
rect 18288 25780 18294 25832
rect 18598 25780 18604 25832
rect 18656 25820 18662 25832
rect 18949 25823 19007 25829
rect 18949 25820 18961 25823
rect 18656 25792 18961 25820
rect 18656 25780 18662 25792
rect 18949 25789 18961 25792
rect 18995 25789 19007 25823
rect 18949 25783 19007 25789
rect 20165 25823 20223 25829
rect 20165 25789 20177 25823
rect 20211 25820 20223 25823
rect 20254 25820 20260 25832
rect 20211 25792 20260 25820
rect 20211 25789 20223 25792
rect 20165 25783 20223 25789
rect 20254 25780 20260 25792
rect 20312 25820 20318 25832
rect 20622 25820 20628 25832
rect 20312 25792 20628 25820
rect 20312 25780 20318 25792
rect 20622 25780 20628 25792
rect 20680 25780 20686 25832
rect 8036 25755 8095 25761
rect 8036 25724 8049 25755
rect 8037 25721 8049 25724
rect 8083 25721 8095 25755
rect 9214 25752 9220 25764
rect 8037 25715 8095 25721
rect 8128 25724 9220 25752
rect 7926 25684 7932 25696
rect 7300 25656 7932 25684
rect 4709 25647 4767 25653
rect 7926 25644 7932 25656
rect 7984 25684 7990 25696
rect 8128 25684 8156 25724
rect 9214 25712 9220 25724
rect 9272 25712 9278 25764
rect 9858 25712 9864 25764
rect 9916 25752 9922 25764
rect 10318 25752 10324 25764
rect 9916 25724 10324 25752
rect 9916 25712 9922 25724
rect 10318 25712 10324 25724
rect 10376 25752 10382 25764
rect 10873 25755 10931 25761
rect 10873 25752 10885 25755
rect 10376 25724 10885 25752
rect 10376 25712 10382 25724
rect 10873 25721 10885 25724
rect 10919 25721 10931 25755
rect 10873 25715 10931 25721
rect 13630 25712 13636 25764
rect 13688 25752 13694 25764
rect 13786 25755 13844 25761
rect 13786 25752 13798 25755
rect 13688 25724 13798 25752
rect 13688 25712 13694 25724
rect 13786 25721 13798 25724
rect 13832 25721 13844 25755
rect 13786 25715 13844 25721
rect 17954 25712 17960 25764
rect 18012 25712 18018 25764
rect 20346 25752 20352 25764
rect 20088 25724 20352 25752
rect 7984 25656 8156 25684
rect 8205 25687 8263 25693
rect 7984 25644 7990 25656
rect 8205 25653 8217 25687
rect 8251 25684 8263 25687
rect 9398 25684 9404 25696
rect 8251 25656 9404 25684
rect 8251 25653 8263 25656
rect 8205 25647 8263 25653
rect 9398 25644 9404 25656
rect 9456 25644 9462 25696
rect 9769 25687 9827 25693
rect 9769 25653 9781 25687
rect 9815 25684 9827 25687
rect 10042 25684 10048 25696
rect 9815 25656 10048 25684
rect 9815 25653 9827 25656
rect 9769 25647 9827 25653
rect 10042 25644 10048 25656
rect 10100 25644 10106 25696
rect 12986 25644 12992 25696
rect 13044 25684 13050 25696
rect 13357 25687 13415 25693
rect 13357 25684 13369 25687
rect 13044 25656 13369 25684
rect 13044 25644 13050 25656
rect 13357 25653 13369 25656
rect 13403 25653 13415 25687
rect 13357 25647 13415 25653
rect 15010 25644 15016 25696
rect 15068 25644 15074 25696
rect 17678 25644 17684 25696
rect 17736 25644 17742 25696
rect 20088 25693 20116 25724
rect 20346 25712 20352 25724
rect 20404 25712 20410 25764
rect 20441 25755 20499 25761
rect 20441 25721 20453 25755
rect 20487 25752 20499 25755
rect 20732 25752 20760 25919
rect 21450 25916 21456 25928
rect 21508 25916 21514 25968
rect 24302 25916 24308 25968
rect 24360 25916 24366 25968
rect 21269 25891 21327 25897
rect 21269 25888 21281 25891
rect 20916 25860 21281 25888
rect 20916 25832 20944 25860
rect 21269 25857 21281 25860
rect 21315 25857 21327 25891
rect 21269 25851 21327 25857
rect 23661 25891 23719 25897
rect 23661 25857 23673 25891
rect 23707 25888 23719 25891
rect 25314 25888 25320 25900
rect 23707 25860 25320 25888
rect 23707 25857 23719 25860
rect 23661 25851 23719 25857
rect 25314 25848 25320 25860
rect 25372 25848 25378 25900
rect 20898 25780 20904 25832
rect 20956 25780 20962 25832
rect 20990 25780 20996 25832
rect 21048 25780 21054 25832
rect 21177 25823 21235 25829
rect 21177 25789 21189 25823
rect 21223 25789 21235 25823
rect 21177 25783 21235 25789
rect 20487 25724 20760 25752
rect 20487 25721 20499 25724
rect 20441 25715 20499 25721
rect 20073 25687 20131 25693
rect 20073 25653 20085 25687
rect 20119 25653 20131 25687
rect 20073 25647 20131 25653
rect 20162 25644 20168 25696
rect 20220 25684 20226 25696
rect 20257 25687 20315 25693
rect 20257 25684 20269 25687
rect 20220 25656 20269 25684
rect 20220 25644 20226 25656
rect 20257 25653 20269 25656
rect 20303 25653 20315 25687
rect 20364 25684 20392 25712
rect 21192 25684 21220 25783
rect 23382 25780 23388 25832
rect 23440 25829 23446 25832
rect 23440 25820 23452 25829
rect 25130 25820 25136 25832
rect 23440 25792 23485 25820
rect 24228 25792 25136 25820
rect 23440 25783 23452 25792
rect 23440 25780 23446 25783
rect 24228 25761 24256 25792
rect 25130 25780 25136 25792
rect 25188 25780 25194 25832
rect 25332 25820 25360 25848
rect 26329 25823 26387 25829
rect 26329 25820 26341 25823
rect 25332 25792 26341 25820
rect 26329 25789 26341 25792
rect 26375 25789 26387 25823
rect 26329 25783 26387 25789
rect 24213 25755 24271 25761
rect 24213 25721 24225 25755
rect 24259 25721 24271 25755
rect 25038 25752 25044 25764
rect 24213 25715 24271 25721
rect 24872 25724 25044 25752
rect 20364 25656 21220 25684
rect 20257 25647 20315 25653
rect 23382 25644 23388 25696
rect 23440 25684 23446 25696
rect 24003 25687 24061 25693
rect 24003 25684 24015 25687
rect 23440 25656 24015 25684
rect 23440 25644 23446 25656
rect 24003 25653 24015 25656
rect 24049 25653 24061 25687
rect 24003 25647 24061 25653
rect 24670 25644 24676 25696
rect 24728 25644 24734 25696
rect 24872 25693 24900 25724
rect 25038 25712 25044 25724
rect 25096 25712 25102 25764
rect 25222 25712 25228 25764
rect 25280 25752 25286 25764
rect 26062 25755 26120 25761
rect 26062 25752 26074 25755
rect 25280 25724 26074 25752
rect 25280 25712 25286 25724
rect 26062 25721 26074 25724
rect 26108 25721 26120 25755
rect 26062 25715 26120 25721
rect 24857 25687 24915 25693
rect 24857 25653 24869 25687
rect 24903 25653 24915 25687
rect 24857 25647 24915 25653
rect 552 25594 27576 25616
rect 552 25542 7114 25594
rect 7166 25542 7178 25594
rect 7230 25542 7242 25594
rect 7294 25542 7306 25594
rect 7358 25542 7370 25594
rect 7422 25542 13830 25594
rect 13882 25542 13894 25594
rect 13946 25542 13958 25594
rect 14010 25542 14022 25594
rect 14074 25542 14086 25594
rect 14138 25542 20546 25594
rect 20598 25542 20610 25594
rect 20662 25542 20674 25594
rect 20726 25542 20738 25594
rect 20790 25542 20802 25594
rect 20854 25542 27262 25594
rect 27314 25542 27326 25594
rect 27378 25542 27390 25594
rect 27442 25542 27454 25594
rect 27506 25542 27518 25594
rect 27570 25542 27576 25594
rect 552 25520 27576 25542
rect 2682 25480 2688 25492
rect 2608 25452 2688 25480
rect 1044 25384 1256 25412
rect 842 25304 848 25356
rect 900 25344 906 25356
rect 1044 25344 1072 25384
rect 1118 25353 1124 25356
rect 900 25316 1072 25344
rect 900 25304 906 25316
rect 1112 25307 1124 25353
rect 1118 25304 1124 25307
rect 1176 25304 1182 25356
rect 1228 25344 1256 25384
rect 2317 25347 2375 25353
rect 1228 25316 2084 25344
rect 2056 25208 2084 25316
rect 2317 25313 2329 25347
rect 2363 25344 2375 25347
rect 2406 25344 2412 25356
rect 2363 25316 2412 25344
rect 2363 25313 2375 25316
rect 2317 25307 2375 25313
rect 2406 25304 2412 25316
rect 2464 25304 2470 25356
rect 2501 25347 2559 25353
rect 2501 25313 2513 25347
rect 2547 25344 2559 25347
rect 2608 25344 2636 25452
rect 2682 25440 2688 25452
rect 2740 25480 2746 25492
rect 4157 25483 4215 25489
rect 4157 25480 4169 25483
rect 2740 25452 4169 25480
rect 2740 25440 2746 25452
rect 4157 25449 4169 25452
rect 4203 25449 4215 25483
rect 4157 25443 4215 25449
rect 4430 25440 4436 25492
rect 4488 25440 4494 25492
rect 5534 25440 5540 25492
rect 5592 25480 5598 25492
rect 5629 25483 5687 25489
rect 5629 25480 5641 25483
rect 5592 25452 5641 25480
rect 5592 25440 5598 25452
rect 5629 25449 5641 25452
rect 5675 25449 5687 25483
rect 5629 25443 5687 25449
rect 7834 25440 7840 25492
rect 7892 25480 7898 25492
rect 9953 25483 10011 25489
rect 9953 25480 9965 25483
rect 7892 25452 9965 25480
rect 7892 25440 7898 25452
rect 9953 25449 9965 25452
rect 9999 25449 10011 25483
rect 9953 25443 10011 25449
rect 10042 25440 10048 25492
rect 10100 25480 10106 25492
rect 10100 25452 12020 25480
rect 10100 25440 10106 25452
rect 3602 25412 3608 25424
rect 2792 25384 3608 25412
rect 2792 25353 2820 25384
rect 3602 25372 3608 25384
rect 3660 25372 3666 25424
rect 6914 25372 6920 25424
rect 6972 25412 6978 25424
rect 7929 25415 7987 25421
rect 7929 25412 7941 25415
rect 6972 25384 7941 25412
rect 6972 25372 6978 25384
rect 7929 25381 7941 25384
rect 7975 25381 7987 25415
rect 7929 25375 7987 25381
rect 8294 25372 8300 25424
rect 8352 25412 8358 25424
rect 9493 25415 9551 25421
rect 9493 25412 9505 25415
rect 8352 25384 9505 25412
rect 8352 25372 8358 25384
rect 9493 25381 9505 25384
rect 9539 25412 9551 25415
rect 11054 25412 11060 25424
rect 9539 25384 11060 25412
rect 9539 25381 9551 25384
rect 9493 25375 9551 25381
rect 11054 25372 11060 25384
rect 11112 25372 11118 25424
rect 11416 25415 11474 25421
rect 11416 25381 11428 25415
rect 11462 25412 11474 25415
rect 11882 25412 11888 25424
rect 11462 25384 11888 25412
rect 11462 25381 11474 25384
rect 11416 25375 11474 25381
rect 11882 25372 11888 25384
rect 11940 25372 11946 25424
rect 11992 25412 12020 25452
rect 12066 25440 12072 25492
rect 12124 25480 12130 25492
rect 12621 25483 12679 25489
rect 12621 25480 12633 25483
rect 12124 25452 12633 25480
rect 12124 25440 12130 25452
rect 12621 25449 12633 25452
rect 12667 25449 12679 25483
rect 12621 25443 12679 25449
rect 13630 25440 13636 25492
rect 13688 25480 13694 25492
rect 13909 25483 13967 25489
rect 13909 25480 13921 25483
rect 13688 25452 13921 25480
rect 13688 25440 13694 25452
rect 13909 25449 13921 25452
rect 13955 25449 13967 25483
rect 13909 25443 13967 25449
rect 14369 25483 14427 25489
rect 14369 25449 14381 25483
rect 14415 25449 14427 25483
rect 14369 25443 14427 25449
rect 14829 25483 14887 25489
rect 14829 25449 14841 25483
rect 14875 25480 14887 25483
rect 15010 25480 15016 25492
rect 14875 25452 15016 25480
rect 14875 25449 14887 25452
rect 14829 25443 14887 25449
rect 12773 25415 12831 25421
rect 12773 25412 12785 25415
rect 11992 25384 12785 25412
rect 12773 25381 12785 25384
rect 12819 25412 12831 25415
rect 12819 25384 12940 25412
rect 12819 25381 12831 25384
rect 12773 25375 12831 25381
rect 3050 25353 3056 25356
rect 2547 25316 2636 25344
rect 2777 25347 2835 25353
rect 2547 25313 2559 25316
rect 2501 25307 2559 25313
rect 2777 25313 2789 25347
rect 2823 25313 2835 25347
rect 3044 25344 3056 25353
rect 3011 25316 3056 25344
rect 2777 25307 2835 25313
rect 3044 25307 3056 25316
rect 2130 25236 2136 25288
rect 2188 25276 2194 25288
rect 2516 25276 2544 25307
rect 2188 25248 2544 25276
rect 2188 25236 2194 25248
rect 2792 25208 2820 25307
rect 3050 25304 3056 25307
rect 3108 25304 3114 25356
rect 4982 25304 4988 25356
rect 5040 25304 5046 25356
rect 5074 25304 5080 25356
rect 5132 25304 5138 25356
rect 7006 25304 7012 25356
rect 7064 25304 7070 25356
rect 7285 25347 7343 25353
rect 7285 25313 7297 25347
rect 7331 25344 7343 25347
rect 7650 25344 7656 25356
rect 7331 25316 7656 25344
rect 7331 25313 7343 25316
rect 7285 25307 7343 25313
rect 7650 25304 7656 25316
rect 7708 25304 7714 25356
rect 7745 25347 7803 25353
rect 7745 25313 7757 25347
rect 7791 25313 7803 25347
rect 7745 25307 7803 25313
rect 7837 25347 7895 25353
rect 7837 25313 7849 25347
rect 7883 25313 7895 25347
rect 7837 25307 7895 25313
rect 8113 25347 8171 25353
rect 8113 25313 8125 25347
rect 8159 25344 8171 25347
rect 8481 25347 8539 25353
rect 8481 25344 8493 25347
rect 8159 25316 8493 25344
rect 8159 25313 8171 25316
rect 8113 25307 8171 25313
rect 8481 25313 8493 25316
rect 8527 25313 8539 25347
rect 8481 25307 8539 25313
rect 9401 25347 9459 25353
rect 9401 25313 9413 25347
rect 9447 25344 9459 25347
rect 9582 25344 9588 25356
rect 9447 25316 9588 25344
rect 9447 25313 9459 25316
rect 9401 25307 9459 25313
rect 4709 25279 4767 25285
rect 4709 25245 4721 25279
rect 4755 25276 4767 25279
rect 4890 25276 4896 25288
rect 4755 25248 4896 25276
rect 4755 25245 4767 25248
rect 4709 25239 4767 25245
rect 4890 25236 4896 25248
rect 4948 25236 4954 25288
rect 5350 25236 5356 25288
rect 5408 25236 5414 25288
rect 6914 25236 6920 25288
rect 6972 25236 6978 25288
rect 7024 25276 7052 25304
rect 7760 25276 7788 25307
rect 7024 25248 7788 25276
rect 7852 25276 7880 25307
rect 9582 25304 9588 25316
rect 9640 25304 9646 25356
rect 9674 25304 9680 25356
rect 9732 25304 9738 25356
rect 10134 25304 10140 25356
rect 10192 25344 10198 25356
rect 10505 25347 10563 25353
rect 10505 25344 10517 25347
rect 10192 25316 10517 25344
rect 10192 25304 10198 25316
rect 10505 25313 10517 25316
rect 10551 25313 10563 25347
rect 10505 25307 10563 25313
rect 11146 25304 11152 25356
rect 11204 25304 11210 25356
rect 12912 25344 12940 25384
rect 12986 25372 12992 25424
rect 13044 25372 13050 25424
rect 13998 25344 14004 25356
rect 12912 25316 14004 25344
rect 13998 25304 14004 25316
rect 14056 25304 14062 25356
rect 14093 25347 14151 25353
rect 14093 25313 14105 25347
rect 14139 25344 14151 25347
rect 14384 25344 14412 25443
rect 15010 25440 15016 25452
rect 15068 25440 15074 25492
rect 19153 25483 19211 25489
rect 19153 25449 19165 25483
rect 19199 25480 19211 25483
rect 19334 25480 19340 25492
rect 19199 25452 19340 25480
rect 19199 25449 19211 25452
rect 19153 25443 19211 25449
rect 19334 25440 19340 25452
rect 19392 25440 19398 25492
rect 20254 25440 20260 25492
rect 20312 25440 20318 25492
rect 21358 25440 21364 25492
rect 21416 25480 21422 25492
rect 22094 25480 22100 25492
rect 21416 25452 22100 25480
rect 21416 25440 21422 25452
rect 22094 25440 22100 25452
rect 22152 25480 22158 25492
rect 22738 25480 22744 25492
rect 22152 25452 22744 25480
rect 22152 25440 22158 25452
rect 22738 25440 22744 25452
rect 22796 25440 22802 25492
rect 23382 25440 23388 25492
rect 23440 25440 23446 25492
rect 24302 25480 24308 25492
rect 23768 25452 24308 25480
rect 17678 25372 17684 25424
rect 17736 25412 17742 25424
rect 18018 25415 18076 25421
rect 18018 25412 18030 25415
rect 17736 25384 18030 25412
rect 17736 25372 17742 25384
rect 18018 25381 18030 25384
rect 18064 25381 18076 25415
rect 18018 25375 18076 25381
rect 14139 25316 14412 25344
rect 14737 25347 14795 25353
rect 14139 25313 14151 25316
rect 14093 25307 14151 25313
rect 14737 25313 14749 25347
rect 14783 25344 14795 25347
rect 14918 25344 14924 25356
rect 14783 25316 14924 25344
rect 14783 25313 14795 25316
rect 14737 25307 14795 25313
rect 14918 25304 14924 25316
rect 14976 25344 14982 25356
rect 18966 25344 18972 25356
rect 14976 25316 18972 25344
rect 14976 25304 14982 25316
rect 18966 25304 18972 25316
rect 19024 25304 19030 25356
rect 19352 25344 19380 25440
rect 22002 25372 22008 25424
rect 22060 25412 22066 25424
rect 23768 25421 23796 25452
rect 24302 25440 24308 25452
rect 24360 25440 24366 25492
rect 24765 25483 24823 25489
rect 24765 25449 24777 25483
rect 24811 25480 24823 25483
rect 25130 25480 25136 25492
rect 24811 25452 25136 25480
rect 24811 25449 24823 25452
rect 24765 25443 24823 25449
rect 25130 25440 25136 25452
rect 25188 25440 25194 25492
rect 25222 25440 25228 25492
rect 25280 25440 25286 25492
rect 23753 25415 23811 25421
rect 22060 25384 23060 25412
rect 22060 25372 22066 25384
rect 20165 25347 20223 25353
rect 20165 25344 20177 25347
rect 19352 25316 20177 25344
rect 20165 25313 20177 25316
rect 20211 25313 20223 25347
rect 20165 25307 20223 25313
rect 21266 25304 21272 25356
rect 21324 25344 21330 25356
rect 21821 25347 21879 25353
rect 21821 25344 21833 25347
rect 21324 25316 21833 25344
rect 21324 25304 21330 25316
rect 21821 25313 21833 25316
rect 21867 25313 21879 25347
rect 21821 25307 21879 25313
rect 22278 25304 22284 25356
rect 22336 25304 22342 25356
rect 22462 25304 22468 25356
rect 22520 25304 22526 25356
rect 22925 25347 22983 25353
rect 22925 25344 22937 25347
rect 22664 25316 22937 25344
rect 7852 25248 7972 25276
rect 2056 25180 2820 25208
rect 7944 25208 7972 25248
rect 8846 25236 8852 25288
rect 8904 25276 8910 25288
rect 9033 25279 9091 25285
rect 9033 25276 9045 25279
rect 8904 25248 9045 25276
rect 8904 25236 8910 25248
rect 9033 25245 9045 25248
rect 9079 25245 9091 25279
rect 9033 25239 9091 25245
rect 15010 25236 15016 25288
rect 15068 25236 15074 25288
rect 17034 25236 17040 25288
rect 17092 25276 17098 25288
rect 17770 25276 17776 25288
rect 17092 25248 17776 25276
rect 17092 25236 17098 25248
rect 17770 25236 17776 25248
rect 17828 25236 17834 25288
rect 21726 25236 21732 25288
rect 21784 25236 21790 25288
rect 22005 25279 22063 25285
rect 22005 25245 22017 25279
rect 22051 25276 22063 25279
rect 22189 25279 22247 25285
rect 22189 25276 22201 25279
rect 22051 25248 22201 25276
rect 22051 25245 22063 25248
rect 22005 25239 22063 25245
rect 22189 25245 22201 25248
rect 22235 25245 22247 25279
rect 22189 25239 22247 25245
rect 22370 25236 22376 25288
rect 22428 25236 22434 25288
rect 22664 25285 22692 25316
rect 22925 25313 22937 25316
rect 22971 25313 22983 25347
rect 23032 25344 23060 25384
rect 23753 25381 23765 25415
rect 23799 25381 23811 25415
rect 24670 25412 24676 25424
rect 23753 25375 23811 25381
rect 23952 25384 24676 25412
rect 23569 25347 23627 25353
rect 23569 25344 23581 25347
rect 23032 25316 23581 25344
rect 22925 25307 22983 25313
rect 23569 25313 23581 25316
rect 23615 25313 23627 25347
rect 23569 25307 23627 25313
rect 23845 25347 23903 25353
rect 23845 25313 23857 25347
rect 23891 25313 23903 25347
rect 23845 25307 23903 25313
rect 22649 25279 22707 25285
rect 22649 25245 22661 25279
rect 22695 25245 22707 25279
rect 22649 25239 22707 25245
rect 22741 25279 22799 25285
rect 22741 25245 22753 25279
rect 22787 25245 22799 25279
rect 22940 25276 22968 25307
rect 23106 25276 23112 25288
rect 22940 25248 23112 25276
rect 22741 25239 22799 25245
rect 9674 25208 9680 25220
rect 7944 25180 9680 25208
rect 9674 25168 9680 25180
rect 9732 25168 9738 25220
rect 9861 25211 9919 25217
rect 9861 25177 9873 25211
rect 9907 25208 9919 25211
rect 10318 25208 10324 25220
rect 9907 25180 10324 25208
rect 9907 25177 9919 25180
rect 9861 25171 9919 25177
rect 10318 25168 10324 25180
rect 10376 25168 10382 25220
rect 22756 25208 22784 25239
rect 23106 25236 23112 25248
rect 23164 25236 23170 25288
rect 23584 25276 23612 25307
rect 23750 25276 23756 25288
rect 23584 25248 23756 25276
rect 23750 25236 23756 25248
rect 23808 25276 23814 25288
rect 23860 25276 23888 25307
rect 23808 25248 23888 25276
rect 23808 25236 23814 25248
rect 23952 25208 23980 25384
rect 24670 25372 24676 25384
rect 24728 25372 24734 25424
rect 24854 25372 24860 25424
rect 24912 25412 24918 25424
rect 24912 25384 25360 25412
rect 24912 25372 24918 25384
rect 24029 25347 24087 25353
rect 24029 25313 24041 25347
rect 24075 25344 24087 25347
rect 24302 25344 24308 25356
rect 24075 25316 24308 25344
rect 24075 25313 24087 25316
rect 24029 25307 24087 25313
rect 24302 25304 24308 25316
rect 24360 25304 24366 25356
rect 25038 25304 25044 25356
rect 25096 25304 25102 25356
rect 25332 25353 25360 25384
rect 25317 25347 25375 25353
rect 25317 25313 25329 25347
rect 25363 25344 25375 25347
rect 25866 25344 25872 25356
rect 25363 25316 25872 25344
rect 25363 25313 25375 25316
rect 25317 25307 25375 25313
rect 25866 25304 25872 25316
rect 25924 25304 25930 25356
rect 25406 25236 25412 25288
rect 25464 25276 25470 25288
rect 26053 25279 26111 25285
rect 26053 25276 26065 25279
rect 25464 25248 26065 25276
rect 25464 25236 25470 25248
rect 26053 25245 26065 25248
rect 26099 25245 26111 25279
rect 26053 25239 26111 25245
rect 12406 25180 12848 25208
rect 2222 25100 2228 25152
rect 2280 25100 2286 25152
rect 2682 25100 2688 25152
rect 2740 25100 2746 25152
rect 4614 25100 4620 25152
rect 4672 25140 4678 25152
rect 5169 25143 5227 25149
rect 5169 25140 5181 25143
rect 4672 25112 5181 25140
rect 4672 25100 4678 25112
rect 5169 25109 5181 25112
rect 5215 25109 5227 25143
rect 5169 25103 5227 25109
rect 7558 25100 7564 25152
rect 7616 25100 7622 25152
rect 10962 25100 10968 25152
rect 11020 25140 11026 25152
rect 12406 25140 12434 25180
rect 11020 25112 12434 25140
rect 12529 25143 12587 25149
rect 11020 25100 11026 25112
rect 12529 25109 12541 25143
rect 12575 25140 12587 25143
rect 12710 25140 12716 25152
rect 12575 25112 12716 25140
rect 12575 25109 12587 25112
rect 12529 25103 12587 25109
rect 12710 25100 12716 25112
rect 12768 25100 12774 25152
rect 12820 25149 12848 25180
rect 22066 25180 22784 25208
rect 23124 25180 23980 25208
rect 12805 25143 12863 25149
rect 12805 25109 12817 25143
rect 12851 25109 12863 25143
rect 12805 25103 12863 25109
rect 17678 25100 17684 25152
rect 17736 25140 17742 25152
rect 22066 25140 22094 25180
rect 23124 25149 23152 25180
rect 17736 25112 22094 25140
rect 23109 25143 23167 25149
rect 17736 25100 17742 25112
rect 23109 25109 23121 25143
rect 23155 25109 23167 25143
rect 23109 25103 23167 25109
rect 23658 25100 23664 25152
rect 23716 25140 23722 25152
rect 23937 25143 23995 25149
rect 23937 25140 23949 25143
rect 23716 25112 23949 25140
rect 23716 25100 23722 25112
rect 23937 25109 23949 25112
rect 23983 25140 23995 25143
rect 24026 25140 24032 25152
rect 23983 25112 24032 25140
rect 23983 25109 23995 25112
rect 23937 25103 23995 25109
rect 24026 25100 24032 25112
rect 24084 25100 24090 25152
rect 552 25050 27416 25072
rect 552 24998 3756 25050
rect 3808 24998 3820 25050
rect 3872 24998 3884 25050
rect 3936 24998 3948 25050
rect 4000 24998 4012 25050
rect 4064 24998 10472 25050
rect 10524 24998 10536 25050
rect 10588 24998 10600 25050
rect 10652 24998 10664 25050
rect 10716 24998 10728 25050
rect 10780 24998 17188 25050
rect 17240 24998 17252 25050
rect 17304 24998 17316 25050
rect 17368 24998 17380 25050
rect 17432 24998 17444 25050
rect 17496 24998 23904 25050
rect 23956 24998 23968 25050
rect 24020 24998 24032 25050
rect 24084 24998 24096 25050
rect 24148 24998 24160 25050
rect 24212 24998 27416 25050
rect 552 24976 27416 24998
rect 1029 24939 1087 24945
rect 1029 24905 1041 24939
rect 1075 24936 1087 24939
rect 1118 24936 1124 24948
rect 1075 24908 1124 24936
rect 1075 24905 1087 24908
rect 1029 24899 1087 24905
rect 1118 24896 1124 24908
rect 1176 24896 1182 24948
rect 1857 24939 1915 24945
rect 1857 24905 1869 24939
rect 1903 24936 1915 24939
rect 1946 24936 1952 24948
rect 1903 24908 1952 24936
rect 1903 24905 1915 24908
rect 1857 24899 1915 24905
rect 1946 24896 1952 24908
rect 2004 24896 2010 24948
rect 2590 24896 2596 24948
rect 2648 24896 2654 24948
rect 2777 24939 2835 24945
rect 2777 24905 2789 24939
rect 2823 24936 2835 24939
rect 2866 24936 2872 24948
rect 2823 24908 2872 24936
rect 2823 24905 2835 24908
rect 2777 24899 2835 24905
rect 2866 24896 2872 24908
rect 2924 24896 2930 24948
rect 4154 24896 4160 24948
rect 4212 24896 4218 24948
rect 4525 24939 4583 24945
rect 4525 24905 4537 24939
rect 4571 24936 4583 24939
rect 5074 24936 5080 24948
rect 4571 24908 5080 24936
rect 4571 24905 4583 24908
rect 4525 24899 4583 24905
rect 5074 24896 5080 24908
rect 5132 24896 5138 24948
rect 5261 24939 5319 24945
rect 5261 24905 5273 24939
rect 5307 24936 5319 24939
rect 5350 24936 5356 24948
rect 5307 24908 5356 24936
rect 5307 24905 5319 24908
rect 5261 24899 5319 24905
rect 5350 24896 5356 24908
rect 5408 24896 5414 24948
rect 9582 24896 9588 24948
rect 9640 24896 9646 24948
rect 10045 24939 10103 24945
rect 10045 24905 10057 24939
rect 10091 24936 10103 24939
rect 10134 24936 10140 24948
rect 10091 24908 10140 24936
rect 10091 24905 10103 24908
rect 10045 24899 10103 24905
rect 10134 24896 10140 24908
rect 10192 24896 10198 24948
rect 11238 24896 11244 24948
rect 11296 24936 11302 24948
rect 11517 24939 11575 24945
rect 11517 24936 11529 24939
rect 11296 24908 11529 24936
rect 11296 24896 11302 24908
rect 11517 24905 11529 24908
rect 11563 24905 11575 24939
rect 11517 24899 11575 24905
rect 14550 24896 14556 24948
rect 14608 24896 14614 24948
rect 15470 24936 15476 24948
rect 15304 24908 15476 24936
rect 9600 24868 9628 24896
rect 9600 24840 10088 24868
rect 10060 24812 10088 24840
rect 2590 24760 2596 24812
rect 2648 24760 2654 24812
rect 2774 24760 2780 24812
rect 2832 24800 2838 24812
rect 2961 24803 3019 24809
rect 2961 24800 2973 24803
rect 2832 24772 2973 24800
rect 2832 24760 2838 24772
rect 2961 24769 2973 24772
rect 3007 24800 3019 24803
rect 3050 24800 3056 24812
rect 3007 24772 3056 24800
rect 3007 24769 3019 24772
rect 2961 24763 3019 24769
rect 3050 24760 3056 24772
rect 3108 24760 3114 24812
rect 4982 24760 4988 24812
rect 5040 24760 5046 24812
rect 8386 24800 8392 24812
rect 7484 24772 8392 24800
rect 1213 24735 1271 24741
rect 1213 24701 1225 24735
rect 1259 24732 1271 24735
rect 1259 24704 1716 24732
rect 1259 24701 1271 24704
rect 1213 24695 1271 24701
rect 1688 24605 1716 24704
rect 2222 24692 2228 24744
rect 2280 24732 2286 24744
rect 2608 24732 2636 24760
rect 2869 24735 2927 24741
rect 2869 24732 2881 24735
rect 2280 24704 2881 24732
rect 2280 24692 2286 24704
rect 2869 24701 2881 24704
rect 2915 24701 2927 24735
rect 2869 24695 2927 24701
rect 3510 24692 3516 24744
rect 3568 24732 3574 24744
rect 4065 24735 4123 24741
rect 4065 24732 4077 24735
rect 3568 24704 4077 24732
rect 3568 24692 3574 24704
rect 4065 24701 4077 24704
rect 4111 24701 4123 24735
rect 4065 24695 4123 24701
rect 1854 24673 1860 24676
rect 1841 24667 1860 24673
rect 1841 24633 1853 24667
rect 1841 24627 1860 24633
rect 1854 24624 1860 24627
rect 1912 24624 1918 24676
rect 2038 24624 2044 24676
rect 2096 24664 2102 24676
rect 2682 24673 2688 24676
rect 2409 24667 2467 24673
rect 2409 24664 2421 24667
rect 2096 24636 2421 24664
rect 2096 24624 2102 24636
rect 2409 24633 2421 24636
rect 2455 24633 2467 24667
rect 2409 24627 2467 24633
rect 2625 24667 2688 24673
rect 2625 24633 2637 24667
rect 2671 24633 2688 24667
rect 2625 24627 2688 24633
rect 2682 24624 2688 24627
rect 2740 24624 2746 24676
rect 4080 24664 4108 24695
rect 4890 24692 4896 24744
rect 4948 24692 4954 24744
rect 5000 24732 5028 24760
rect 7484 24744 7512 24772
rect 8386 24760 8392 24772
rect 8444 24760 8450 24812
rect 10042 24760 10048 24812
rect 10100 24760 10106 24812
rect 11146 24760 11152 24812
rect 11204 24800 11210 24812
rect 11977 24803 12035 24809
rect 11977 24800 11989 24803
rect 11204 24772 11989 24800
rect 11204 24760 11210 24772
rect 11977 24769 11989 24772
rect 12023 24769 12035 24803
rect 11977 24763 12035 24769
rect 13354 24760 13360 24812
rect 13412 24800 13418 24812
rect 13633 24803 13691 24809
rect 13633 24800 13645 24803
rect 13412 24772 13645 24800
rect 13412 24760 13418 24772
rect 13633 24769 13645 24772
rect 13679 24769 13691 24803
rect 13633 24763 13691 24769
rect 14277 24803 14335 24809
rect 14277 24769 14289 24803
rect 14323 24800 14335 24803
rect 14323 24772 15148 24800
rect 14323 24769 14335 24772
rect 14277 24763 14335 24769
rect 7101 24735 7159 24741
rect 5000 24704 6960 24732
rect 4080 24636 5764 24664
rect 5736 24605 5764 24636
rect 6178 24624 6184 24676
rect 6236 24664 6242 24676
rect 6834 24667 6892 24673
rect 6834 24664 6846 24667
rect 6236 24636 6846 24664
rect 6236 24624 6242 24636
rect 6834 24633 6846 24636
rect 6880 24633 6892 24667
rect 6932 24664 6960 24704
rect 7101 24701 7113 24735
rect 7147 24732 7159 24735
rect 7466 24732 7472 24744
rect 7147 24704 7472 24732
rect 7147 24701 7159 24704
rect 7101 24695 7159 24701
rect 7466 24692 7472 24704
rect 7524 24692 7530 24744
rect 7834 24692 7840 24744
rect 7892 24692 7898 24744
rect 8665 24735 8723 24741
rect 8665 24701 8677 24735
rect 8711 24732 8723 24735
rect 9490 24732 9496 24744
rect 8711 24704 9496 24732
rect 8711 24701 8723 24704
rect 8665 24695 8723 24701
rect 9490 24692 9496 24704
rect 9548 24732 9554 24744
rect 10137 24735 10195 24741
rect 10137 24732 10149 24735
rect 9548 24704 10149 24732
rect 9548 24692 9554 24704
rect 10137 24701 10149 24704
rect 10183 24732 10195 24735
rect 10404 24735 10462 24741
rect 10183 24704 10272 24732
rect 10183 24701 10195 24704
rect 10137 24695 10195 24701
rect 8754 24664 8760 24676
rect 6932 24636 8760 24664
rect 6834 24627 6892 24633
rect 8754 24624 8760 24636
rect 8812 24624 8818 24676
rect 8932 24667 8990 24673
rect 8932 24633 8944 24667
rect 8978 24664 8990 24667
rect 9306 24664 9312 24676
rect 8978 24636 9312 24664
rect 8978 24633 8990 24636
rect 8932 24627 8990 24633
rect 9306 24624 9312 24636
rect 9364 24624 9370 24676
rect 1673 24599 1731 24605
rect 1673 24565 1685 24599
rect 1719 24565 1731 24599
rect 1673 24559 1731 24565
rect 5721 24599 5779 24605
rect 5721 24565 5733 24599
rect 5767 24596 5779 24599
rect 6270 24596 6276 24608
rect 5767 24568 6276 24596
rect 5767 24565 5779 24568
rect 5721 24559 5779 24565
rect 6270 24556 6276 24568
rect 6328 24556 6334 24608
rect 6730 24556 6736 24608
rect 6788 24596 6794 24608
rect 7193 24599 7251 24605
rect 7193 24596 7205 24599
rect 6788 24568 7205 24596
rect 6788 24556 6794 24568
rect 7193 24565 7205 24568
rect 7239 24565 7251 24599
rect 10244 24596 10272 24704
rect 10404 24701 10416 24735
rect 10450 24701 10462 24735
rect 10404 24695 10462 24701
rect 10318 24624 10324 24676
rect 10376 24664 10382 24676
rect 10428 24664 10456 24695
rect 13998 24692 14004 24744
rect 14056 24732 14062 24744
rect 14458 24732 14464 24744
rect 14056 24704 14464 24732
rect 14056 24692 14062 24704
rect 14458 24692 14464 24704
rect 14516 24732 14522 24744
rect 14516 24701 14565 24732
rect 14516 24692 14519 24701
rect 10376 24636 10456 24664
rect 12244 24667 12302 24673
rect 10376 24624 10382 24636
rect 12244 24633 12256 24667
rect 12290 24664 12302 24667
rect 12618 24664 12624 24676
rect 12290 24636 12624 24664
rect 12290 24633 12302 24636
rect 12244 24627 12302 24633
rect 12618 24624 12624 24636
rect 12676 24624 12682 24676
rect 14507 24667 14519 24692
rect 14553 24667 14565 24701
rect 14642 24692 14648 24744
rect 14700 24732 14706 24744
rect 15013 24735 15071 24741
rect 15013 24732 15025 24735
rect 14700 24704 15025 24732
rect 14700 24692 14706 24704
rect 15013 24701 15025 24704
rect 15059 24701 15071 24735
rect 15013 24695 15071 24701
rect 14507 24661 14565 24667
rect 14737 24667 14795 24673
rect 14737 24633 14749 24667
rect 14783 24664 14795 24667
rect 15120 24664 15148 24772
rect 15304 24741 15332 24908
rect 15470 24896 15476 24908
rect 15528 24936 15534 24948
rect 15746 24936 15752 24948
rect 15528 24908 15752 24936
rect 15528 24896 15534 24908
rect 15746 24896 15752 24908
rect 15804 24936 15810 24948
rect 22097 24939 22155 24945
rect 15804 24908 17724 24936
rect 15804 24896 15810 24908
rect 17696 24880 17724 24908
rect 22097 24905 22109 24939
rect 22143 24936 22155 24939
rect 22370 24936 22376 24948
rect 22143 24908 22376 24936
rect 22143 24905 22155 24908
rect 22097 24899 22155 24905
rect 22370 24896 22376 24908
rect 22428 24896 22434 24948
rect 23109 24939 23167 24945
rect 23109 24905 23121 24939
rect 23155 24905 23167 24939
rect 23109 24899 23167 24905
rect 17678 24828 17684 24880
rect 17736 24828 17742 24880
rect 17770 24828 17776 24880
rect 17828 24828 17834 24880
rect 18049 24871 18107 24877
rect 18049 24837 18061 24871
rect 18095 24868 18107 24871
rect 18138 24868 18144 24880
rect 18095 24840 18144 24868
rect 18095 24837 18107 24840
rect 18049 24831 18107 24837
rect 18138 24828 18144 24840
rect 18196 24828 18202 24880
rect 22005 24871 22063 24877
rect 22005 24837 22017 24871
rect 22051 24868 22063 24871
rect 22186 24868 22192 24880
rect 22051 24840 22192 24868
rect 22051 24837 22063 24840
rect 22005 24831 22063 24837
rect 22186 24828 22192 24840
rect 22244 24828 22250 24880
rect 15473 24803 15531 24809
rect 15473 24769 15485 24803
rect 15519 24800 15531 24803
rect 15562 24800 15568 24812
rect 15519 24772 15568 24800
rect 15519 24769 15531 24772
rect 15473 24763 15531 24769
rect 15562 24760 15568 24772
rect 15620 24760 15626 24812
rect 17696 24800 17724 24828
rect 17604 24772 17724 24800
rect 17788 24800 17816 24828
rect 19337 24803 19395 24809
rect 19337 24800 19349 24803
rect 17788 24772 19349 24800
rect 15289 24735 15347 24741
rect 15289 24701 15301 24735
rect 15335 24701 15347 24735
rect 15289 24695 15347 24701
rect 15654 24692 15660 24744
rect 15712 24692 15718 24744
rect 15930 24692 15936 24744
rect 15988 24732 15994 24744
rect 17034 24732 17040 24744
rect 15988 24704 17040 24732
rect 15988 24692 15994 24704
rect 17034 24692 17040 24704
rect 17092 24692 17098 24744
rect 17604 24741 17632 24772
rect 19337 24769 19349 24772
rect 19383 24769 19395 24803
rect 23124 24800 23152 24899
rect 23750 24896 23756 24948
rect 23808 24936 23814 24948
rect 24029 24939 24087 24945
rect 24029 24936 24041 24939
rect 23808 24908 24041 24936
rect 23808 24896 23814 24908
rect 24029 24905 24041 24908
rect 24075 24905 24087 24939
rect 24029 24899 24087 24905
rect 24213 24871 24271 24877
rect 24213 24837 24225 24871
rect 24259 24837 24271 24871
rect 24213 24831 24271 24837
rect 19337 24763 19395 24769
rect 22066 24772 23152 24800
rect 23293 24803 23351 24809
rect 17589 24735 17647 24741
rect 17589 24701 17601 24735
rect 17635 24701 17647 24735
rect 17589 24695 17647 24701
rect 17681 24735 17739 24741
rect 17681 24701 17693 24735
rect 17727 24701 17739 24735
rect 17681 24695 17739 24701
rect 16178 24667 16236 24673
rect 16178 24664 16190 24667
rect 14783 24636 15148 24664
rect 15856 24636 16190 24664
rect 14783 24633 14795 24636
rect 14737 24627 14795 24633
rect 11146 24596 11152 24608
rect 10244 24568 11152 24596
rect 7193 24559 7251 24565
rect 11146 24556 11152 24568
rect 11204 24556 11210 24608
rect 13354 24556 13360 24608
rect 13412 24556 13418 24608
rect 13446 24556 13452 24608
rect 13504 24596 13510 24608
rect 14369 24599 14427 24605
rect 14369 24596 14381 24599
rect 13504 24568 14381 24596
rect 13504 24556 13510 24568
rect 14369 24565 14381 24568
rect 14415 24565 14427 24599
rect 14369 24559 14427 24565
rect 14826 24556 14832 24608
rect 14884 24556 14890 24608
rect 15102 24556 15108 24608
rect 15160 24556 15166 24608
rect 15856 24605 15884 24636
rect 16178 24633 16190 24636
rect 16224 24633 16236 24667
rect 17696 24664 17724 24695
rect 17954 24692 17960 24744
rect 18012 24732 18018 24744
rect 18049 24735 18107 24741
rect 18049 24732 18061 24735
rect 18012 24704 18061 24732
rect 18012 24692 18018 24704
rect 18049 24701 18061 24704
rect 18095 24701 18107 24735
rect 18049 24695 18107 24701
rect 18325 24735 18383 24741
rect 18325 24701 18337 24735
rect 18371 24701 18383 24735
rect 18325 24695 18383 24701
rect 16178 24627 16236 24633
rect 17328 24636 17724 24664
rect 18340 24664 18368 24695
rect 19058 24692 19064 24744
rect 19116 24692 19122 24744
rect 22066 24732 22094 24772
rect 23293 24769 23305 24803
rect 23339 24800 23351 24803
rect 24228 24800 24256 24831
rect 23339 24772 24256 24800
rect 23339 24769 23351 24772
rect 23293 24763 23351 24769
rect 19168 24704 22094 24732
rect 23017 24735 23075 24741
rect 18414 24664 18420 24676
rect 18340 24636 18420 24664
rect 15841 24599 15899 24605
rect 15841 24565 15853 24599
rect 15887 24565 15899 24599
rect 15841 24559 15899 24565
rect 16942 24556 16948 24608
rect 17000 24596 17006 24608
rect 17328 24605 17356 24636
rect 18414 24624 18420 24636
rect 18472 24664 18478 24676
rect 19168 24664 19196 24704
rect 23017 24701 23029 24735
rect 23063 24732 23075 24735
rect 23106 24732 23112 24744
rect 23063 24704 23112 24732
rect 23063 24701 23075 24704
rect 23017 24695 23075 24701
rect 23106 24692 23112 24704
rect 23164 24692 23170 24744
rect 19582 24667 19640 24673
rect 19582 24664 19594 24667
rect 18472 24636 19196 24664
rect 19260 24636 19594 24664
rect 18472 24624 18478 24636
rect 17313 24599 17371 24605
rect 17313 24596 17325 24599
rect 17000 24568 17325 24596
rect 17000 24556 17006 24568
rect 17313 24565 17325 24568
rect 17359 24565 17371 24599
rect 17313 24559 17371 24565
rect 17402 24556 17408 24608
rect 17460 24556 17466 24608
rect 19260 24605 19288 24636
rect 19582 24633 19594 24636
rect 19628 24633 19640 24667
rect 19582 24627 19640 24633
rect 21358 24624 21364 24676
rect 21416 24664 21422 24676
rect 21637 24667 21695 24673
rect 21637 24664 21649 24667
rect 21416 24636 21649 24664
rect 21416 24624 21422 24636
rect 21637 24633 21649 24636
rect 21683 24664 21695 24667
rect 21726 24664 21732 24676
rect 21683 24636 21732 24664
rect 21683 24633 21695 24636
rect 21637 24627 21695 24633
rect 21726 24624 21732 24636
rect 21784 24624 21790 24676
rect 23750 24624 23756 24676
rect 23808 24664 23814 24676
rect 23845 24667 23903 24673
rect 23845 24664 23857 24667
rect 23808 24636 23857 24664
rect 23808 24624 23814 24636
rect 23845 24633 23857 24636
rect 23891 24633 23903 24667
rect 23845 24627 23903 24633
rect 24026 24624 24032 24676
rect 24084 24673 24090 24676
rect 24084 24667 24103 24673
rect 24091 24633 24103 24667
rect 24228 24664 24256 24772
rect 24486 24760 24492 24812
rect 24544 24800 24550 24812
rect 24544 24772 25084 24800
rect 24544 24760 24550 24772
rect 24305 24735 24363 24741
rect 24305 24701 24317 24735
rect 24351 24732 24363 24735
rect 24394 24732 24400 24744
rect 24351 24704 24400 24732
rect 24351 24701 24363 24704
rect 24305 24695 24363 24701
rect 24394 24692 24400 24704
rect 24452 24692 24458 24744
rect 24581 24735 24639 24741
rect 24581 24701 24593 24735
rect 24627 24732 24639 24735
rect 24670 24732 24676 24744
rect 24627 24704 24676 24732
rect 24627 24701 24639 24704
rect 24581 24695 24639 24701
rect 24670 24692 24676 24704
rect 24728 24692 24734 24744
rect 24854 24741 24860 24744
rect 24847 24735 24860 24741
rect 24847 24732 24859 24735
rect 24780 24704 24859 24732
rect 24780 24664 24808 24704
rect 24847 24701 24859 24704
rect 24847 24695 24860 24701
rect 24854 24692 24860 24695
rect 24912 24692 24918 24744
rect 25056 24741 25084 24772
rect 25041 24735 25099 24741
rect 25041 24701 25053 24735
rect 25087 24701 25099 24735
rect 25041 24695 25099 24701
rect 25133 24735 25191 24741
rect 25133 24701 25145 24735
rect 25179 24701 25191 24735
rect 25133 24695 25191 24701
rect 24228 24636 24808 24664
rect 24084 24627 24103 24633
rect 24084 24624 24090 24627
rect 25148 24608 25176 24695
rect 25314 24692 25320 24744
rect 25372 24692 25378 24744
rect 25406 24692 25412 24744
rect 25464 24732 25470 24744
rect 25685 24735 25743 24741
rect 25685 24732 25697 24735
rect 25464 24704 25697 24732
rect 25464 24692 25470 24704
rect 25685 24701 25697 24704
rect 25731 24701 25743 24735
rect 25685 24695 25743 24701
rect 25952 24667 26010 24673
rect 25952 24633 25964 24667
rect 25998 24664 26010 24667
rect 26050 24664 26056 24676
rect 25998 24636 26056 24664
rect 25998 24633 26010 24636
rect 25952 24627 26010 24633
rect 26050 24624 26056 24636
rect 26108 24624 26114 24676
rect 19245 24599 19303 24605
rect 19245 24565 19257 24599
rect 19291 24565 19303 24599
rect 19245 24559 19303 24565
rect 20717 24599 20775 24605
rect 20717 24565 20729 24599
rect 20763 24596 20775 24599
rect 20898 24596 20904 24608
rect 20763 24568 20904 24596
rect 20763 24565 20775 24568
rect 20717 24559 20775 24565
rect 20898 24556 20904 24568
rect 20956 24556 20962 24608
rect 23382 24556 23388 24608
rect 23440 24596 23446 24608
rect 23569 24599 23627 24605
rect 23569 24596 23581 24599
rect 23440 24568 23581 24596
rect 23440 24556 23446 24568
rect 23569 24565 23581 24568
rect 23615 24565 23627 24599
rect 23569 24559 23627 24565
rect 24302 24556 24308 24608
rect 24360 24596 24366 24608
rect 24397 24599 24455 24605
rect 24397 24596 24409 24599
rect 24360 24568 24409 24596
rect 24360 24556 24366 24568
rect 24397 24565 24409 24568
rect 24443 24565 24455 24599
rect 24397 24559 24455 24565
rect 24762 24556 24768 24608
rect 24820 24556 24826 24608
rect 25041 24599 25099 24605
rect 25041 24565 25053 24599
rect 25087 24596 25099 24599
rect 25130 24596 25136 24608
rect 25087 24568 25136 24596
rect 25087 24565 25099 24568
rect 25041 24559 25099 24565
rect 25130 24556 25136 24568
rect 25188 24556 25194 24608
rect 25317 24599 25375 24605
rect 25317 24565 25329 24599
rect 25363 24596 25375 24599
rect 25774 24596 25780 24608
rect 25363 24568 25780 24596
rect 25363 24565 25375 24568
rect 25317 24559 25375 24565
rect 25774 24556 25780 24568
rect 25832 24556 25838 24608
rect 26878 24556 26884 24608
rect 26936 24596 26942 24608
rect 27065 24599 27123 24605
rect 27065 24596 27077 24599
rect 26936 24568 27077 24596
rect 26936 24556 26942 24568
rect 27065 24565 27077 24568
rect 27111 24565 27123 24599
rect 27065 24559 27123 24565
rect 552 24506 27576 24528
rect 552 24454 7114 24506
rect 7166 24454 7178 24506
rect 7230 24454 7242 24506
rect 7294 24454 7306 24506
rect 7358 24454 7370 24506
rect 7422 24454 13830 24506
rect 13882 24454 13894 24506
rect 13946 24454 13958 24506
rect 14010 24454 14022 24506
rect 14074 24454 14086 24506
rect 14138 24454 20546 24506
rect 20598 24454 20610 24506
rect 20662 24454 20674 24506
rect 20726 24454 20738 24506
rect 20790 24454 20802 24506
rect 20854 24454 27262 24506
rect 27314 24454 27326 24506
rect 27378 24454 27390 24506
rect 27442 24454 27454 24506
rect 27506 24454 27518 24506
rect 27570 24454 27576 24506
rect 552 24432 27576 24454
rect 6178 24352 6184 24404
rect 6236 24352 6242 24404
rect 6270 24352 6276 24404
rect 6328 24392 6334 24404
rect 7834 24392 7840 24404
rect 6328 24364 7840 24392
rect 6328 24352 6334 24364
rect 7834 24352 7840 24364
rect 7892 24352 7898 24404
rect 8846 24352 8852 24404
rect 8904 24352 8910 24404
rect 9306 24352 9312 24404
rect 9364 24352 9370 24404
rect 9950 24352 9956 24404
rect 10008 24392 10014 24404
rect 10318 24401 10324 24404
rect 10295 24395 10324 24401
rect 10295 24392 10307 24395
rect 10008 24364 10307 24392
rect 10008 24352 10014 24364
rect 10295 24361 10307 24364
rect 10295 24355 10324 24361
rect 10318 24352 10324 24355
rect 10376 24352 10382 24404
rect 12618 24352 12624 24404
rect 12676 24352 12682 24404
rect 12710 24352 12716 24404
rect 12768 24392 12774 24404
rect 12989 24395 13047 24401
rect 12989 24392 13001 24395
rect 12768 24364 13001 24392
rect 12768 24352 12774 24364
rect 12989 24361 13001 24364
rect 13035 24392 13047 24395
rect 14182 24392 14188 24404
rect 13035 24364 14188 24392
rect 13035 24361 13047 24364
rect 12989 24355 13047 24361
rect 14182 24352 14188 24364
rect 14240 24352 14246 24404
rect 15562 24352 15568 24404
rect 15620 24352 15626 24404
rect 15654 24352 15660 24404
rect 15712 24392 15718 24404
rect 16117 24395 16175 24401
rect 16117 24392 16129 24395
rect 15712 24364 16129 24392
rect 15712 24352 15718 24364
rect 16117 24361 16129 24364
rect 16163 24361 16175 24395
rect 16117 24355 16175 24361
rect 16577 24395 16635 24401
rect 16577 24361 16589 24395
rect 16623 24392 16635 24395
rect 17402 24392 17408 24404
rect 16623 24364 17408 24392
rect 16623 24361 16635 24364
rect 16577 24355 16635 24361
rect 17402 24352 17408 24364
rect 17460 24352 17466 24404
rect 19058 24352 19064 24404
rect 19116 24392 19122 24404
rect 19521 24395 19579 24401
rect 19521 24392 19533 24395
rect 19116 24364 19533 24392
rect 19116 24352 19122 24364
rect 19521 24361 19533 24364
rect 19567 24361 19579 24395
rect 19521 24355 19579 24361
rect 22097 24395 22155 24401
rect 22097 24361 22109 24395
rect 22143 24392 22155 24395
rect 22186 24392 22192 24404
rect 22143 24364 22192 24392
rect 22143 24361 22155 24364
rect 22097 24355 22155 24361
rect 22186 24352 22192 24364
rect 22244 24352 22250 24404
rect 23569 24395 23627 24401
rect 23569 24392 23581 24395
rect 23308 24364 23581 24392
rect 2590 24324 2596 24336
rect 1780 24296 2596 24324
rect 1780 24265 1808 24296
rect 2590 24284 2596 24296
rect 2648 24284 2654 24336
rect 6549 24327 6607 24333
rect 6549 24293 6561 24327
rect 6595 24324 6607 24327
rect 6914 24324 6920 24336
rect 6595 24296 6920 24324
rect 6595 24293 6607 24296
rect 6549 24287 6607 24293
rect 6914 24284 6920 24296
rect 6972 24324 6978 24336
rect 7009 24327 7067 24333
rect 7009 24324 7021 24327
rect 6972 24296 7021 24324
rect 6972 24284 6978 24296
rect 7009 24293 7021 24296
rect 7055 24293 7067 24327
rect 7009 24287 7067 24293
rect 7101 24327 7159 24333
rect 7101 24293 7113 24327
rect 7147 24324 7159 24327
rect 7147 24296 7512 24324
rect 7147 24293 7159 24296
rect 7101 24287 7159 24293
rect 1765 24259 1823 24265
rect 1765 24225 1777 24259
rect 1811 24225 1823 24259
rect 1765 24219 1823 24225
rect 1949 24259 2007 24265
rect 1949 24225 1961 24259
rect 1995 24256 2007 24259
rect 2225 24259 2283 24265
rect 1995 24228 2084 24256
rect 1995 24225 2007 24228
rect 1949 24219 2007 24225
rect 1854 24012 1860 24064
rect 1912 24012 1918 24064
rect 2056 24061 2084 24228
rect 2225 24225 2237 24259
rect 2271 24256 2283 24259
rect 2314 24256 2320 24268
rect 2271 24228 2320 24256
rect 2271 24225 2283 24228
rect 2225 24219 2283 24225
rect 2314 24216 2320 24228
rect 2372 24216 2378 24268
rect 2866 24216 2872 24268
rect 2924 24216 2930 24268
rect 4798 24216 4804 24268
rect 4856 24216 4862 24268
rect 6365 24259 6423 24265
rect 6365 24225 6377 24259
rect 6411 24225 6423 24259
rect 6365 24219 6423 24225
rect 6457 24259 6515 24265
rect 6457 24225 6469 24259
rect 6503 24225 6515 24259
rect 6457 24219 6515 24225
rect 2130 24148 2136 24200
rect 2188 24188 2194 24200
rect 2409 24191 2467 24197
rect 2409 24188 2421 24191
rect 2188 24160 2421 24188
rect 2188 24148 2194 24160
rect 2409 24157 2421 24160
rect 2455 24188 2467 24191
rect 4816 24188 4844 24216
rect 2455 24160 4844 24188
rect 2455 24157 2467 24160
rect 2409 24151 2467 24157
rect 3602 24080 3608 24132
rect 3660 24120 3666 24132
rect 5442 24120 5448 24132
rect 3660 24092 5448 24120
rect 3660 24080 3666 24092
rect 5442 24080 5448 24092
rect 5500 24080 5506 24132
rect 6380 24120 6408 24219
rect 6472 24188 6500 24219
rect 6730 24216 6736 24268
rect 6788 24216 6794 24268
rect 6822 24216 6828 24268
rect 6880 24216 6886 24268
rect 7190 24216 7196 24268
rect 7248 24216 7254 24268
rect 7484 24256 7512 24296
rect 7558 24284 7564 24336
rect 7616 24324 7622 24336
rect 7714 24327 7772 24333
rect 7714 24324 7726 24327
rect 7616 24296 7726 24324
rect 7616 24284 7622 24296
rect 7714 24293 7726 24296
rect 7760 24293 7772 24327
rect 7714 24287 7772 24293
rect 10505 24327 10563 24333
rect 10505 24293 10517 24327
rect 10551 24324 10563 24327
rect 10965 24327 11023 24333
rect 10965 24324 10977 24327
rect 10551 24296 10977 24324
rect 10551 24293 10563 24296
rect 10505 24287 10563 24293
rect 10965 24293 10977 24296
rect 11011 24293 11023 24327
rect 13446 24324 13452 24336
rect 10965 24287 11023 24293
rect 12820 24296 13452 24324
rect 8018 24256 8024 24268
rect 7484 24228 8024 24256
rect 8018 24216 8024 24228
rect 8076 24256 8082 24268
rect 8294 24256 8300 24268
rect 8076 24228 8300 24256
rect 8076 24216 8082 24228
rect 8294 24216 8300 24228
rect 8352 24216 8358 24268
rect 9398 24216 9404 24268
rect 9456 24256 9462 24268
rect 9493 24259 9551 24265
rect 9493 24256 9505 24259
rect 9456 24228 9505 24256
rect 9456 24216 9462 24228
rect 9493 24225 9505 24228
rect 9539 24225 9551 24259
rect 9493 24219 9551 24225
rect 9674 24216 9680 24268
rect 9732 24216 9738 24268
rect 9769 24259 9827 24265
rect 9769 24225 9781 24259
rect 9815 24256 9827 24259
rect 10042 24256 10048 24268
rect 9815 24228 10048 24256
rect 9815 24225 9827 24228
rect 9769 24219 9827 24225
rect 10042 24216 10048 24228
rect 10100 24216 10106 24268
rect 11146 24216 11152 24268
rect 11204 24256 11210 24268
rect 12820 24265 12848 24296
rect 13446 24284 13452 24296
rect 13504 24284 13510 24336
rect 15930 24324 15936 24336
rect 14200 24296 15936 24324
rect 11885 24259 11943 24265
rect 11885 24256 11897 24259
rect 11204 24228 11897 24256
rect 11204 24216 11210 24228
rect 11885 24225 11897 24228
rect 11931 24225 11943 24259
rect 11885 24219 11943 24225
rect 12805 24259 12863 24265
rect 12805 24225 12817 24259
rect 12851 24225 12863 24259
rect 12805 24219 12863 24225
rect 7374 24188 7380 24200
rect 6472 24160 7380 24188
rect 7374 24148 7380 24160
rect 7432 24148 7438 24200
rect 7466 24148 7472 24200
rect 7524 24148 7530 24200
rect 9692 24188 9720 24216
rect 9692 24160 9812 24188
rect 7006 24120 7012 24132
rect 6380 24092 7012 24120
rect 7006 24080 7012 24092
rect 7064 24120 7070 24132
rect 7190 24120 7196 24132
rect 7064 24092 7196 24120
rect 7064 24080 7070 24092
rect 7190 24080 7196 24092
rect 7248 24080 7254 24132
rect 9784 24120 9812 24160
rect 10226 24148 10232 24200
rect 10284 24188 10290 24200
rect 11517 24191 11575 24197
rect 11517 24188 11529 24191
rect 10284 24160 11529 24188
rect 10284 24148 10290 24160
rect 11517 24157 11529 24160
rect 11563 24157 11575 24191
rect 11517 24151 11575 24157
rect 10962 24120 10968 24132
rect 9784 24092 10968 24120
rect 10962 24080 10968 24092
rect 11020 24080 11026 24132
rect 11698 24080 11704 24132
rect 11756 24080 11762 24132
rect 11900 24120 11928 24219
rect 13078 24216 13084 24268
rect 13136 24216 13142 24268
rect 14200 24265 14228 24296
rect 15930 24284 15936 24296
rect 15988 24284 15994 24336
rect 21818 24324 21824 24336
rect 19076 24296 20576 24324
rect 14185 24259 14243 24265
rect 14185 24225 14197 24259
rect 14231 24225 14243 24259
rect 14185 24219 14243 24225
rect 14452 24259 14510 24265
rect 14452 24225 14464 24259
rect 14498 24256 14510 24259
rect 14826 24256 14832 24268
rect 14498 24228 14832 24256
rect 14498 24225 14510 24228
rect 14452 24219 14510 24225
rect 14826 24216 14832 24228
rect 14884 24216 14890 24268
rect 15010 24216 15016 24268
rect 15068 24256 15074 24268
rect 15068 24228 16068 24256
rect 15068 24216 15074 24228
rect 16040 24188 16068 24228
rect 16206 24216 16212 24268
rect 16264 24256 16270 24268
rect 19076 24265 19104 24296
rect 16485 24259 16543 24265
rect 16485 24256 16497 24259
rect 16264 24228 16497 24256
rect 16264 24216 16270 24228
rect 16485 24225 16497 24228
rect 16531 24225 16543 24259
rect 17773 24259 17831 24265
rect 17773 24256 17785 24259
rect 16485 24219 16543 24225
rect 17512 24228 17785 24256
rect 16390 24188 16396 24200
rect 16040 24160 16396 24188
rect 16390 24148 16396 24160
rect 16448 24188 16454 24200
rect 16669 24191 16727 24197
rect 16669 24188 16681 24191
rect 16448 24160 16681 24188
rect 16448 24148 16454 24160
rect 16669 24157 16681 24160
rect 16715 24157 16727 24191
rect 16669 24151 16727 24157
rect 11900 24092 14228 24120
rect 2041 24055 2099 24061
rect 2041 24021 2053 24055
rect 2087 24052 2099 24055
rect 2682 24052 2688 24064
rect 2087 24024 2688 24052
rect 2087 24021 2099 24024
rect 2041 24015 2099 24021
rect 2682 24012 2688 24024
rect 2740 24012 2746 24064
rect 2774 24012 2780 24064
rect 2832 24012 2838 24064
rect 4154 24012 4160 24064
rect 4212 24052 4218 24064
rect 4341 24055 4399 24061
rect 4341 24052 4353 24055
rect 4212 24024 4353 24052
rect 4212 24012 4218 24024
rect 4341 24021 4353 24024
rect 4387 24021 4399 24055
rect 4341 24015 4399 24021
rect 4709 24055 4767 24061
rect 4709 24021 4721 24055
rect 4755 24052 4767 24055
rect 4890 24052 4896 24064
rect 4755 24024 4896 24052
rect 4755 24021 4767 24024
rect 4709 24015 4767 24021
rect 4890 24012 4896 24024
rect 4948 24012 4954 24064
rect 7377 24055 7435 24061
rect 7377 24021 7389 24055
rect 7423 24052 7435 24055
rect 8754 24052 8760 24064
rect 7423 24024 8760 24052
rect 7423 24021 7435 24024
rect 7377 24015 7435 24021
rect 8754 24012 8760 24024
rect 8812 24012 8818 24064
rect 10134 24012 10140 24064
rect 10192 24012 10198 24064
rect 10321 24055 10379 24061
rect 10321 24021 10333 24055
rect 10367 24052 10379 24055
rect 10870 24052 10876 24064
rect 10367 24024 10876 24052
rect 10367 24021 10379 24024
rect 10321 24015 10379 24021
rect 10870 24012 10876 24024
rect 10928 24012 10934 24064
rect 11716 24052 11744 24080
rect 12986 24052 12992 24064
rect 11716 24024 12992 24052
rect 12986 24012 12992 24024
rect 13044 24052 13050 24064
rect 13722 24052 13728 24064
rect 13044 24024 13728 24052
rect 13044 24012 13050 24024
rect 13722 24012 13728 24024
rect 13780 24012 13786 24064
rect 14200 24052 14228 24092
rect 16482 24052 16488 24064
rect 14200 24024 16488 24052
rect 16482 24012 16488 24024
rect 16540 24052 16546 24064
rect 17512 24052 17540 24228
rect 17773 24225 17785 24228
rect 17819 24256 17831 24259
rect 19061 24259 19119 24265
rect 19061 24256 19073 24259
rect 17819 24228 19073 24256
rect 17819 24225 17831 24228
rect 17773 24219 17831 24225
rect 19061 24225 19073 24228
rect 19107 24225 19119 24259
rect 19889 24259 19947 24265
rect 19889 24256 19901 24259
rect 19061 24219 19119 24225
rect 19168 24228 19901 24256
rect 17957 24191 18015 24197
rect 17957 24157 17969 24191
rect 18003 24188 18015 24191
rect 18138 24188 18144 24200
rect 18003 24160 18144 24188
rect 18003 24157 18015 24160
rect 17957 24151 18015 24157
rect 18138 24148 18144 24160
rect 18196 24148 18202 24200
rect 18966 24148 18972 24200
rect 19024 24188 19030 24200
rect 19168 24188 19196 24228
rect 19889 24225 19901 24228
rect 19935 24225 19947 24259
rect 19889 24219 19947 24225
rect 19981 24259 20039 24265
rect 19981 24225 19993 24259
rect 20027 24256 20039 24259
rect 20349 24259 20407 24265
rect 20349 24256 20361 24259
rect 20027 24228 20361 24256
rect 20027 24225 20039 24228
rect 19981 24219 20039 24225
rect 20349 24225 20361 24228
rect 20395 24225 20407 24259
rect 20349 24219 20407 24225
rect 20438 24216 20444 24268
rect 20496 24256 20502 24268
rect 20548 24265 20576 24296
rect 20916 24296 21588 24324
rect 20916 24268 20944 24296
rect 20533 24259 20591 24265
rect 20533 24256 20545 24259
rect 20496 24228 20545 24256
rect 20496 24216 20502 24228
rect 20533 24225 20545 24228
rect 20579 24225 20591 24259
rect 20533 24219 20591 24225
rect 20717 24259 20775 24265
rect 20717 24225 20729 24259
rect 20763 24256 20775 24259
rect 20898 24256 20904 24268
rect 20763 24228 20904 24256
rect 20763 24225 20775 24228
rect 20717 24219 20775 24225
rect 20898 24216 20904 24228
rect 20956 24216 20962 24268
rect 20990 24216 20996 24268
rect 21048 24256 21054 24268
rect 21560 24265 21588 24296
rect 21652 24296 21824 24324
rect 21652 24265 21680 24296
rect 21818 24284 21824 24296
rect 21876 24324 21882 24336
rect 23308 24324 23336 24364
rect 23569 24361 23581 24364
rect 23615 24392 23627 24395
rect 24302 24392 24308 24404
rect 23615 24364 24308 24392
rect 23615 24361 23627 24364
rect 23569 24355 23627 24361
rect 24302 24352 24308 24364
rect 24360 24352 24366 24404
rect 24394 24352 24400 24404
rect 24452 24352 24458 24404
rect 25501 24395 25559 24401
rect 25501 24361 25513 24395
rect 25547 24392 25559 24395
rect 25793 24395 25851 24401
rect 25793 24392 25805 24395
rect 25547 24364 25805 24392
rect 25547 24361 25559 24364
rect 25501 24355 25559 24361
rect 25793 24361 25805 24364
rect 25839 24392 25851 24395
rect 25958 24392 25964 24404
rect 25839 24364 25964 24392
rect 25839 24361 25851 24364
rect 25793 24355 25851 24361
rect 25958 24352 25964 24364
rect 26016 24352 26022 24404
rect 26050 24352 26056 24404
rect 26108 24352 26114 24404
rect 21876 24296 23336 24324
rect 21876 24284 21882 24296
rect 23382 24284 23388 24336
rect 23440 24284 23446 24336
rect 24486 24284 24492 24336
rect 24544 24324 24550 24336
rect 24673 24327 24731 24333
rect 24673 24324 24685 24327
rect 24544 24296 24685 24324
rect 24544 24284 24550 24296
rect 24673 24293 24685 24296
rect 24719 24293 24731 24327
rect 24673 24287 24731 24293
rect 24854 24284 24860 24336
rect 24912 24284 24918 24336
rect 25222 24284 25228 24336
rect 25280 24324 25286 24336
rect 25590 24324 25596 24336
rect 25280 24296 25596 24324
rect 25280 24284 25286 24296
rect 25590 24284 25596 24296
rect 25648 24284 25654 24336
rect 26789 24327 26847 24333
rect 26789 24324 26801 24327
rect 25700 24296 26801 24324
rect 21361 24259 21419 24265
rect 21361 24256 21373 24259
rect 21048 24228 21373 24256
rect 21048 24216 21054 24228
rect 21361 24225 21373 24228
rect 21407 24225 21419 24259
rect 21361 24219 21419 24225
rect 21545 24259 21603 24265
rect 21545 24225 21557 24259
rect 21591 24225 21603 24259
rect 21545 24219 21603 24225
rect 21637 24259 21695 24265
rect 21637 24225 21649 24259
rect 21683 24225 21695 24259
rect 21637 24219 21695 24225
rect 21913 24259 21971 24265
rect 21913 24225 21925 24259
rect 21959 24256 21971 24259
rect 22186 24256 22192 24268
rect 21959 24228 22192 24256
rect 21959 24225 21971 24228
rect 21913 24219 21971 24225
rect 22186 24216 22192 24228
rect 22244 24216 22250 24268
rect 23658 24216 23664 24268
rect 23716 24216 23722 24268
rect 25130 24216 25136 24268
rect 25188 24216 25194 24268
rect 25314 24216 25320 24268
rect 25372 24256 25378 24268
rect 25700 24256 25728 24296
rect 26789 24293 26801 24296
rect 26835 24293 26847 24327
rect 26789 24287 26847 24293
rect 26237 24259 26295 24265
rect 26237 24256 26249 24259
rect 25372 24228 25728 24256
rect 25976 24228 26249 24256
rect 25372 24216 25378 24228
rect 19024 24160 19196 24188
rect 19245 24191 19303 24197
rect 19024 24148 19030 24160
rect 19245 24157 19257 24191
rect 19291 24188 19303 24191
rect 19794 24188 19800 24200
rect 19291 24160 19800 24188
rect 19291 24157 19303 24160
rect 19245 24151 19303 24157
rect 19794 24148 19800 24160
rect 19852 24148 19858 24200
rect 20070 24148 20076 24200
rect 20128 24148 20134 24200
rect 20806 24148 20812 24200
rect 20864 24188 20870 24200
rect 21729 24191 21787 24197
rect 21729 24188 21741 24191
rect 20864 24160 21741 24188
rect 20864 24148 20870 24160
rect 21729 24157 21741 24160
rect 21775 24188 21787 24191
rect 22094 24188 22100 24200
rect 21775 24160 22100 24188
rect 21775 24157 21787 24160
rect 21729 24151 21787 24157
rect 22094 24148 22100 24160
rect 22152 24148 22158 24200
rect 23293 24191 23351 24197
rect 23293 24157 23305 24191
rect 23339 24157 23351 24191
rect 23293 24151 23351 24157
rect 23308 24120 23336 24151
rect 23750 24148 23756 24200
rect 23808 24148 23814 24200
rect 25332 24188 25360 24216
rect 24421 24160 25360 24188
rect 23385 24123 23443 24129
rect 23385 24120 23397 24123
rect 23308 24092 23397 24120
rect 23385 24089 23397 24092
rect 23431 24089 23443 24123
rect 23385 24083 23443 24089
rect 16540 24024 17540 24052
rect 16540 24012 16546 24024
rect 17586 24012 17592 24064
rect 17644 24012 17650 24064
rect 18874 24012 18880 24064
rect 18932 24012 18938 24064
rect 22646 24012 22652 24064
rect 22704 24012 22710 24064
rect 23290 24012 23296 24064
rect 23348 24052 23354 24064
rect 24421 24052 24449 24160
rect 25976 24129 26004 24228
rect 26237 24225 26249 24228
rect 26283 24225 26295 24259
rect 26237 24219 26295 24225
rect 26878 24216 26884 24268
rect 26936 24216 26942 24268
rect 25961 24123 26019 24129
rect 25961 24089 25973 24123
rect 26007 24089 26019 24123
rect 25961 24083 26019 24089
rect 23348 24024 24449 24052
rect 23348 24012 23354 24024
rect 24486 24012 24492 24064
rect 24544 24012 24550 24064
rect 25774 24012 25780 24064
rect 25832 24012 25838 24064
rect 552 23962 27416 23984
rect 552 23910 3756 23962
rect 3808 23910 3820 23962
rect 3872 23910 3884 23962
rect 3936 23910 3948 23962
rect 4000 23910 4012 23962
rect 4064 23910 10472 23962
rect 10524 23910 10536 23962
rect 10588 23910 10600 23962
rect 10652 23910 10664 23962
rect 10716 23910 10728 23962
rect 10780 23910 17188 23962
rect 17240 23910 17252 23962
rect 17304 23910 17316 23962
rect 17368 23910 17380 23962
rect 17432 23910 17444 23962
rect 17496 23910 23904 23962
rect 23956 23910 23968 23962
rect 24020 23910 24032 23962
rect 24084 23910 24096 23962
rect 24148 23910 24160 23962
rect 24212 23910 27416 23962
rect 552 23888 27416 23910
rect 1213 23851 1271 23857
rect 1213 23817 1225 23851
rect 1259 23848 1271 23851
rect 1581 23851 1639 23857
rect 1581 23848 1593 23851
rect 1259 23820 1593 23848
rect 1259 23817 1271 23820
rect 1213 23811 1271 23817
rect 1581 23817 1593 23820
rect 1627 23817 1639 23851
rect 1581 23811 1639 23817
rect 2314 23808 2320 23860
rect 2372 23808 2378 23860
rect 2590 23808 2596 23860
rect 2648 23848 2654 23860
rect 2777 23851 2835 23857
rect 2777 23848 2789 23851
rect 2648 23820 2789 23848
rect 2648 23808 2654 23820
rect 2777 23817 2789 23820
rect 2823 23817 2835 23851
rect 4798 23848 4804 23860
rect 2777 23811 2835 23817
rect 3528 23820 4804 23848
rect 1397 23783 1455 23789
rect 1397 23780 1409 23783
rect 860 23752 1409 23780
rect 860 23653 888 23752
rect 1397 23749 1409 23752
rect 1443 23749 1455 23783
rect 1397 23743 1455 23749
rect 2038 23740 2044 23792
rect 2096 23780 2102 23792
rect 2501 23783 2559 23789
rect 2501 23780 2513 23783
rect 2096 23752 2513 23780
rect 2096 23740 2102 23752
rect 2501 23749 2513 23752
rect 2547 23749 2559 23783
rect 2501 23743 2559 23749
rect 2774 23712 2780 23724
rect 1320 23684 2780 23712
rect 1320 23653 1348 23684
rect 2774 23672 2780 23684
rect 2832 23672 2838 23724
rect 845 23647 903 23653
rect 845 23613 857 23647
rect 891 23613 903 23647
rect 845 23607 903 23613
rect 1121 23647 1179 23653
rect 1121 23613 1133 23647
rect 1167 23613 1179 23647
rect 1121 23607 1179 23613
rect 1305 23647 1363 23653
rect 1305 23613 1317 23647
rect 1351 23613 1363 23647
rect 1305 23607 1363 23613
rect 1949 23647 2007 23653
rect 1949 23613 1961 23647
rect 1995 23644 2007 23647
rect 3421 23647 3479 23653
rect 1995 23616 2636 23644
rect 1995 23613 2007 23616
rect 1949 23607 2007 23613
rect 1136 23576 1164 23607
rect 1854 23576 1860 23588
rect 1136 23548 1860 23576
rect 1854 23536 1860 23548
rect 1912 23536 1918 23588
rect 2130 23536 2136 23588
rect 2188 23536 2194 23588
rect 1029 23511 1087 23517
rect 1029 23477 1041 23511
rect 1075 23508 1087 23511
rect 1118 23508 1124 23520
rect 1075 23480 1124 23508
rect 1075 23477 1087 23480
rect 1029 23471 1087 23477
rect 1118 23468 1124 23480
rect 1176 23468 1182 23520
rect 1486 23468 1492 23520
rect 1544 23508 1550 23520
rect 1581 23511 1639 23517
rect 1581 23508 1593 23511
rect 1544 23480 1593 23508
rect 1544 23468 1550 23480
rect 1581 23477 1593 23480
rect 1627 23477 1639 23511
rect 1581 23471 1639 23477
rect 2314 23468 2320 23520
rect 2372 23517 2378 23520
rect 2372 23511 2391 23517
rect 2379 23477 2391 23511
rect 2372 23471 2391 23477
rect 2372 23468 2378 23471
rect 2498 23468 2504 23520
rect 2556 23508 2562 23520
rect 2608 23517 2636 23616
rect 3421 23613 3433 23647
rect 3467 23644 3479 23647
rect 3528 23644 3556 23820
rect 4798 23808 4804 23820
rect 4856 23808 4862 23860
rect 4893 23851 4951 23857
rect 4893 23817 4905 23851
rect 4939 23848 4951 23851
rect 4985 23851 5043 23857
rect 4985 23848 4997 23851
rect 4939 23820 4997 23848
rect 4939 23817 4951 23820
rect 4893 23811 4951 23817
rect 4985 23817 4997 23820
rect 5031 23817 5043 23851
rect 4985 23811 5043 23817
rect 4908 23780 4936 23811
rect 5166 23808 5172 23860
rect 5224 23848 5230 23860
rect 5350 23848 5356 23860
rect 5224 23820 5356 23848
rect 5224 23808 5230 23820
rect 5350 23808 5356 23820
rect 5408 23808 5414 23860
rect 6822 23808 6828 23860
rect 6880 23848 6886 23860
rect 8389 23851 8447 23857
rect 8389 23848 8401 23851
rect 6880 23820 8401 23848
rect 6880 23808 6886 23820
rect 8389 23817 8401 23820
rect 8435 23817 8447 23851
rect 8389 23811 8447 23817
rect 10226 23808 10232 23860
rect 10284 23848 10290 23860
rect 10873 23851 10931 23857
rect 10873 23848 10885 23851
rect 10284 23820 10885 23848
rect 10284 23808 10290 23820
rect 10873 23817 10885 23820
rect 10919 23817 10931 23851
rect 10873 23811 10931 23817
rect 12713 23851 12771 23857
rect 12713 23817 12725 23851
rect 12759 23848 12771 23851
rect 12894 23848 12900 23860
rect 12759 23820 12900 23848
rect 12759 23817 12771 23820
rect 12713 23811 12771 23817
rect 12894 23808 12900 23820
rect 12952 23848 12958 23860
rect 12952 23820 13676 23848
rect 12952 23808 12958 23820
rect 4080 23752 4936 23780
rect 3467 23616 3556 23644
rect 3467 23613 3479 23616
rect 3421 23607 3479 23613
rect 3786 23604 3792 23656
rect 3844 23604 3850 23656
rect 3878 23604 3884 23656
rect 3936 23604 3942 23656
rect 4080 23653 4108 23752
rect 7190 23740 7196 23792
rect 7248 23780 7254 23792
rect 7558 23780 7564 23792
rect 7248 23752 7564 23780
rect 7248 23740 7254 23752
rect 7558 23740 7564 23752
rect 7616 23740 7622 23792
rect 13648 23780 13676 23820
rect 13722 23808 13728 23860
rect 13780 23848 13786 23860
rect 14550 23848 14556 23860
rect 13780 23820 14556 23848
rect 13780 23808 13786 23820
rect 14550 23808 14556 23820
rect 14608 23808 14614 23860
rect 14642 23808 14648 23860
rect 14700 23808 14706 23860
rect 18138 23808 18144 23860
rect 18196 23848 18202 23860
rect 20806 23848 20812 23860
rect 18196 23820 20812 23848
rect 18196 23808 18202 23820
rect 20806 23808 20812 23820
rect 20864 23808 20870 23860
rect 23661 23851 23719 23857
rect 21192 23820 22232 23848
rect 14001 23783 14059 23789
rect 13648 23752 13952 23780
rect 4522 23672 4528 23724
rect 4580 23712 4586 23724
rect 4580 23684 5212 23712
rect 4580 23672 4586 23684
rect 3973 23647 4031 23653
rect 3973 23613 3985 23647
rect 4019 23613 4031 23647
rect 3973 23607 4031 23613
rect 4065 23647 4123 23653
rect 4065 23613 4077 23647
rect 4111 23613 4123 23647
rect 4065 23607 4123 23613
rect 2682 23536 2688 23588
rect 2740 23585 2746 23588
rect 2740 23579 2803 23585
rect 2740 23545 2757 23579
rect 2791 23576 2803 23579
rect 2791 23548 2833 23576
rect 2791 23545 2803 23548
rect 2740 23539 2803 23545
rect 2740 23536 2746 23539
rect 2866 23536 2872 23588
rect 2924 23576 2930 23588
rect 2961 23579 3019 23585
rect 2961 23576 2973 23579
rect 2924 23548 2973 23576
rect 2924 23536 2930 23548
rect 2961 23545 2973 23548
rect 3007 23545 3019 23579
rect 2961 23539 3019 23545
rect 3513 23579 3571 23585
rect 3513 23545 3525 23579
rect 3559 23545 3571 23579
rect 3513 23539 3571 23545
rect 2593 23511 2651 23517
rect 2593 23508 2605 23511
rect 2556 23480 2605 23508
rect 2556 23468 2562 23480
rect 2593 23477 2605 23480
rect 2639 23477 2651 23511
rect 3528 23508 3556 23539
rect 3694 23536 3700 23588
rect 3752 23576 3758 23588
rect 3988 23576 4016 23607
rect 4338 23604 4344 23656
rect 4396 23604 4402 23656
rect 4617 23647 4675 23653
rect 4617 23644 4629 23647
rect 4448 23616 4629 23644
rect 4448 23576 4476 23616
rect 4617 23613 4629 23616
rect 4663 23613 4675 23647
rect 4617 23607 4675 23613
rect 4709 23647 4767 23653
rect 4709 23613 4721 23647
rect 4755 23644 4767 23647
rect 4890 23644 4896 23656
rect 4755 23616 4896 23644
rect 4755 23613 4767 23616
rect 4709 23607 4767 23613
rect 3752 23548 4016 23576
rect 4080 23548 4476 23576
rect 3752 23536 3758 23548
rect 4080 23508 4108 23548
rect 4522 23536 4528 23588
rect 4580 23536 4586 23588
rect 3528 23480 4108 23508
rect 4249 23511 4307 23517
rect 2593 23471 2651 23477
rect 4249 23477 4261 23511
rect 4295 23508 4307 23511
rect 4614 23508 4620 23520
rect 4295 23480 4620 23508
rect 4295 23477 4307 23480
rect 4249 23471 4307 23477
rect 4614 23468 4620 23480
rect 4672 23468 4678 23520
rect 4816 23508 4844 23616
rect 4890 23604 4896 23616
rect 4948 23604 4954 23656
rect 4982 23604 4988 23656
rect 5040 23604 5046 23656
rect 5074 23604 5080 23656
rect 5132 23604 5138 23656
rect 5184 23644 5212 23684
rect 5442 23672 5448 23724
rect 5500 23672 5506 23724
rect 6472 23684 7880 23712
rect 6472 23644 6500 23684
rect 7852 23656 7880 23684
rect 9490 23672 9496 23724
rect 9548 23672 9554 23724
rect 10502 23672 10508 23724
rect 10560 23712 10566 23724
rect 10870 23712 10876 23724
rect 10560 23684 10876 23712
rect 10560 23672 10566 23684
rect 10870 23672 10876 23684
rect 10928 23712 10934 23724
rect 10965 23715 11023 23721
rect 10965 23712 10977 23715
rect 10928 23684 10977 23712
rect 10928 23672 10934 23684
rect 10965 23681 10977 23684
rect 11011 23681 11023 23715
rect 10965 23675 11023 23681
rect 5184 23616 6500 23644
rect 7745 23647 7803 23653
rect 7745 23613 7757 23647
rect 7791 23613 7803 23647
rect 7745 23607 7803 23613
rect 5712 23579 5770 23585
rect 5712 23545 5724 23579
rect 5758 23576 5770 23579
rect 6454 23576 6460 23588
rect 5758 23548 6460 23576
rect 5758 23545 5770 23548
rect 5712 23539 5770 23545
rect 6454 23536 6460 23548
rect 6512 23536 6518 23588
rect 7760 23576 7788 23607
rect 7834 23604 7840 23656
rect 7892 23644 7898 23656
rect 8941 23647 8999 23653
rect 8941 23644 8953 23647
rect 7892 23616 8953 23644
rect 7892 23604 7898 23616
rect 8941 23613 8953 23616
rect 8987 23613 8999 23647
rect 8941 23607 8999 23613
rect 11146 23604 11152 23656
rect 11204 23604 11210 23656
rect 11330 23604 11336 23656
rect 11388 23604 11394 23656
rect 12802 23604 12808 23656
rect 12860 23604 12866 23656
rect 13081 23647 13139 23653
rect 13081 23613 13093 23647
rect 13127 23644 13139 23647
rect 13354 23644 13360 23656
rect 13127 23616 13360 23644
rect 13127 23613 13139 23616
rect 13081 23607 13139 23613
rect 13354 23604 13360 23616
rect 13412 23604 13418 23656
rect 6840 23548 7788 23576
rect 9760 23579 9818 23585
rect 6840 23517 6868 23548
rect 9760 23545 9772 23579
rect 9806 23576 9818 23579
rect 9950 23576 9956 23588
rect 9806 23548 9956 23576
rect 9806 23545 9818 23548
rect 9760 23539 9818 23545
rect 9950 23536 9956 23548
rect 10008 23536 10014 23588
rect 11600 23579 11658 23585
rect 11600 23545 11612 23579
rect 11646 23576 11658 23579
rect 11790 23576 11796 23588
rect 11646 23548 11796 23576
rect 11646 23545 11658 23548
rect 11600 23539 11658 23545
rect 11790 23536 11796 23548
rect 11848 23536 11854 23588
rect 11882 23536 11888 23588
rect 11940 23576 11946 23588
rect 13924 23585 13952 23752
rect 14001 23749 14013 23783
rect 14047 23780 14059 23783
rect 14182 23780 14188 23792
rect 14047 23752 14188 23780
rect 14047 23749 14059 23752
rect 14001 23743 14059 23749
rect 14182 23740 14188 23752
rect 14240 23740 14246 23792
rect 15010 23740 15016 23792
rect 15068 23780 15074 23792
rect 15068 23752 15240 23780
rect 15068 23740 15074 23752
rect 15102 23672 15108 23724
rect 15160 23672 15166 23724
rect 15212 23721 15240 23752
rect 19794 23740 19800 23792
rect 19852 23780 19858 23792
rect 20073 23783 20131 23789
rect 20073 23780 20085 23783
rect 19852 23752 20085 23780
rect 19852 23740 19858 23752
rect 20073 23749 20085 23752
rect 20119 23780 20131 23783
rect 20346 23780 20352 23792
rect 20119 23752 20352 23780
rect 20119 23749 20131 23752
rect 20073 23743 20131 23749
rect 20346 23740 20352 23752
rect 20404 23740 20410 23792
rect 21192 23780 21220 23820
rect 20824 23752 21220 23780
rect 15197 23715 15255 23721
rect 15197 23681 15209 23715
rect 15243 23681 15255 23715
rect 15197 23675 15255 23681
rect 15286 23672 15292 23724
rect 15344 23712 15350 23724
rect 16761 23715 16819 23721
rect 16761 23712 16773 23715
rect 15344 23684 16773 23712
rect 15344 23672 15350 23684
rect 16761 23681 16773 23684
rect 16807 23681 16819 23715
rect 16761 23675 16819 23681
rect 17770 23672 17776 23724
rect 17828 23712 17834 23724
rect 18693 23715 18751 23721
rect 18693 23712 18705 23715
rect 17828 23684 18705 23712
rect 17828 23672 17834 23684
rect 18693 23681 18705 23684
rect 18739 23681 18751 23715
rect 20824 23712 20852 23752
rect 21266 23740 21272 23792
rect 21324 23740 21330 23792
rect 21358 23740 21364 23792
rect 21416 23740 21422 23792
rect 18693 23675 18751 23681
rect 20732 23684 20852 23712
rect 14185 23647 14243 23653
rect 14185 23613 14197 23647
rect 14231 23644 14243 23647
rect 14274 23644 14280 23656
rect 14231 23616 14280 23644
rect 14231 23613 14243 23616
rect 14185 23607 14243 23613
rect 14274 23604 14280 23616
rect 14332 23604 14338 23656
rect 16485 23647 16543 23653
rect 16485 23613 16497 23647
rect 16531 23644 16543 23647
rect 16850 23644 16856 23656
rect 16531 23616 16856 23644
rect 16531 23613 16543 23616
rect 16485 23607 16543 23613
rect 16850 23604 16856 23616
rect 16908 23604 16914 23656
rect 18322 23604 18328 23656
rect 18380 23604 18386 23656
rect 20349 23647 20407 23653
rect 20349 23613 20361 23647
rect 20395 23644 20407 23647
rect 20438 23644 20444 23656
rect 20395 23616 20444 23644
rect 20395 23613 20407 23616
rect 20349 23607 20407 23613
rect 20438 23604 20444 23616
rect 20496 23604 20502 23656
rect 20732 23653 20760 23684
rect 20898 23672 20904 23724
rect 20956 23712 20962 23724
rect 20956 23684 21772 23712
rect 20956 23672 20962 23684
rect 20533 23647 20591 23653
rect 20533 23613 20545 23647
rect 20579 23613 20591 23647
rect 20533 23607 20591 23613
rect 20717 23647 20775 23653
rect 20717 23613 20729 23647
rect 20763 23613 20775 23647
rect 20717 23607 20775 23613
rect 13909 23579 13967 23585
rect 11940 23548 13584 23576
rect 11940 23536 11946 23548
rect 6825 23511 6883 23517
rect 6825 23508 6837 23511
rect 4816 23480 6837 23508
rect 6825 23477 6837 23480
rect 6871 23477 6883 23511
rect 6825 23471 6883 23477
rect 7006 23468 7012 23520
rect 7064 23508 7070 23520
rect 7193 23511 7251 23517
rect 7193 23508 7205 23511
rect 7064 23480 7205 23508
rect 7064 23468 7070 23480
rect 7193 23477 7205 23480
rect 7239 23477 7251 23511
rect 7193 23471 7251 23477
rect 7374 23468 7380 23520
rect 7432 23508 7438 23520
rect 7742 23508 7748 23520
rect 7432 23480 7748 23508
rect 7432 23468 7438 23480
rect 7742 23468 7748 23480
rect 7800 23468 7806 23520
rect 10042 23468 10048 23520
rect 10100 23508 10106 23520
rect 12066 23508 12072 23520
rect 10100 23480 12072 23508
rect 10100 23468 10106 23480
rect 12066 23468 12072 23480
rect 12124 23508 12130 23520
rect 12434 23508 12440 23520
rect 12124 23480 12440 23508
rect 12124 23468 12130 23480
rect 12434 23468 12440 23480
rect 12492 23508 12498 23520
rect 12897 23511 12955 23517
rect 12897 23508 12909 23511
rect 12492 23480 12909 23508
rect 12492 23468 12498 23480
rect 12897 23477 12909 23480
rect 12943 23508 12955 23511
rect 13078 23508 13084 23520
rect 12943 23480 13084 23508
rect 12943 23477 12955 23480
rect 12897 23471 12955 23477
rect 13078 23468 13084 23480
rect 13136 23468 13142 23520
rect 13556 23517 13584 23548
rect 13909 23545 13921 23579
rect 13955 23545 13967 23579
rect 13909 23539 13967 23545
rect 15654 23536 15660 23588
rect 15712 23576 15718 23588
rect 16025 23579 16083 23585
rect 16025 23576 16037 23579
rect 15712 23548 16037 23576
rect 15712 23536 15718 23548
rect 16025 23545 16037 23548
rect 16071 23576 16083 23579
rect 16298 23576 16304 23588
rect 16071 23548 16304 23576
rect 16071 23545 16083 23548
rect 16025 23539 16083 23545
rect 16298 23536 16304 23548
rect 16356 23536 16362 23588
rect 17006 23579 17064 23585
rect 17006 23576 17018 23579
rect 16684 23548 17018 23576
rect 13541 23511 13599 23517
rect 13541 23477 13553 23511
rect 13587 23477 13599 23511
rect 13541 23471 13599 23477
rect 13709 23511 13767 23517
rect 13709 23477 13721 23511
rect 13755 23508 13767 23511
rect 14458 23508 14464 23520
rect 13755 23480 14464 23508
rect 13755 23477 13767 23480
rect 13709 23471 13767 23477
rect 14458 23468 14464 23480
rect 14516 23468 14522 23520
rect 15010 23468 15016 23520
rect 15068 23468 15074 23520
rect 15838 23468 15844 23520
rect 15896 23508 15902 23520
rect 16684 23517 16712 23548
rect 17006 23545 17018 23548
rect 17052 23545 17064 23579
rect 18938 23579 18996 23585
rect 18938 23576 18950 23579
rect 17006 23539 17064 23545
rect 18524 23548 18950 23576
rect 18524 23517 18552 23548
rect 18938 23545 18950 23548
rect 18984 23545 18996 23579
rect 20548 23576 20576 23607
rect 20990 23604 20996 23656
rect 21048 23604 21054 23656
rect 21082 23604 21088 23656
rect 21140 23604 21146 23656
rect 21744 23653 21772 23684
rect 21499 23647 21557 23653
rect 21499 23644 21511 23647
rect 21192 23616 21511 23644
rect 20898 23576 20904 23588
rect 20548 23548 20904 23576
rect 18938 23539 18996 23545
rect 20898 23536 20904 23548
rect 20956 23576 20962 23588
rect 21192 23576 21220 23616
rect 21499 23613 21511 23616
rect 21545 23613 21557 23647
rect 21499 23607 21557 23613
rect 21729 23647 21787 23653
rect 21729 23613 21741 23647
rect 21775 23613 21787 23647
rect 21729 23607 21787 23613
rect 21818 23604 21824 23656
rect 21876 23653 21882 23656
rect 21876 23647 21915 23653
rect 21903 23613 21915 23647
rect 21876 23607 21915 23613
rect 22005 23647 22063 23653
rect 22005 23613 22017 23647
rect 22051 23613 22063 23647
rect 22005 23607 22063 23613
rect 21876 23604 21882 23607
rect 20956 23548 21220 23576
rect 20956 23536 20962 23548
rect 21634 23536 21640 23588
rect 21692 23536 21698 23588
rect 16117 23511 16175 23517
rect 16117 23508 16129 23511
rect 15896 23480 16129 23508
rect 15896 23468 15902 23480
rect 16117 23477 16129 23480
rect 16163 23477 16175 23511
rect 16117 23471 16175 23477
rect 16669 23511 16727 23517
rect 16669 23477 16681 23511
rect 16715 23477 16727 23511
rect 16669 23471 16727 23477
rect 18509 23511 18567 23517
rect 18509 23477 18521 23511
rect 18555 23477 18567 23511
rect 18509 23471 18567 23477
rect 20162 23468 20168 23520
rect 20220 23468 20226 23520
rect 21082 23468 21088 23520
rect 21140 23508 21146 23520
rect 21910 23508 21916 23520
rect 21140 23480 21916 23508
rect 21140 23468 21146 23480
rect 21910 23468 21916 23480
rect 21968 23508 21974 23520
rect 22020 23508 22048 23607
rect 22204 23520 22232 23820
rect 23661 23817 23673 23851
rect 23707 23848 23719 23851
rect 23750 23848 23756 23860
rect 23707 23820 23756 23848
rect 23707 23817 23719 23820
rect 23661 23811 23719 23817
rect 23750 23808 23756 23820
rect 23808 23808 23814 23860
rect 23842 23808 23848 23860
rect 23900 23848 23906 23860
rect 24029 23851 24087 23857
rect 24029 23848 24041 23851
rect 23900 23820 24041 23848
rect 23900 23808 23906 23820
rect 24029 23817 24041 23820
rect 24075 23848 24087 23851
rect 24394 23848 24400 23860
rect 24075 23820 24400 23848
rect 24075 23817 24087 23820
rect 24029 23811 24087 23817
rect 24394 23808 24400 23820
rect 24452 23808 24458 23860
rect 25501 23715 25559 23721
rect 25501 23681 25513 23715
rect 25547 23712 25559 23715
rect 25590 23712 25596 23724
rect 25547 23684 25596 23712
rect 25547 23681 25559 23684
rect 25501 23675 25559 23681
rect 25590 23672 25596 23684
rect 25648 23672 25654 23724
rect 22281 23647 22339 23653
rect 22281 23613 22293 23647
rect 22327 23644 22339 23647
rect 25406 23644 25412 23656
rect 22327 23616 25412 23644
rect 22327 23613 22339 23616
rect 22281 23607 22339 23613
rect 25406 23604 25412 23616
rect 25464 23604 25470 23656
rect 25958 23604 25964 23656
rect 26016 23604 26022 23656
rect 26694 23604 26700 23656
rect 26752 23604 26758 23656
rect 22548 23579 22606 23585
rect 22548 23545 22560 23579
rect 22594 23576 22606 23579
rect 22646 23576 22652 23588
rect 22594 23548 22652 23576
rect 22594 23545 22606 23548
rect 22548 23539 22606 23545
rect 22646 23536 22652 23548
rect 22704 23536 22710 23588
rect 24762 23536 24768 23588
rect 24820 23576 24826 23588
rect 25142 23579 25200 23585
rect 25142 23576 25154 23579
rect 24820 23548 25154 23576
rect 24820 23536 24826 23548
rect 25142 23545 25154 23548
rect 25188 23545 25200 23579
rect 25869 23579 25927 23585
rect 25869 23576 25881 23579
rect 25142 23539 25200 23545
rect 25240 23548 25881 23576
rect 21968 23480 22048 23508
rect 21968 23468 21974 23480
rect 22186 23468 22192 23520
rect 22244 23508 22250 23520
rect 25240 23508 25268 23548
rect 25869 23545 25881 23548
rect 25915 23576 25927 23579
rect 26605 23579 26663 23585
rect 26605 23576 26617 23579
rect 25915 23548 26617 23576
rect 25915 23545 25927 23548
rect 25869 23539 25927 23545
rect 26605 23545 26617 23548
rect 26651 23545 26663 23579
rect 26605 23539 26663 23545
rect 22244 23480 25268 23508
rect 22244 23468 22250 23480
rect 25774 23468 25780 23520
rect 25832 23468 25838 23520
rect 552 23418 27576 23440
rect 552 23366 7114 23418
rect 7166 23366 7178 23418
rect 7230 23366 7242 23418
rect 7294 23366 7306 23418
rect 7358 23366 7370 23418
rect 7422 23366 13830 23418
rect 13882 23366 13894 23418
rect 13946 23366 13958 23418
rect 14010 23366 14022 23418
rect 14074 23366 14086 23418
rect 14138 23366 20546 23418
rect 20598 23366 20610 23418
rect 20662 23366 20674 23418
rect 20726 23366 20738 23418
rect 20790 23366 20802 23418
rect 20854 23366 27262 23418
rect 27314 23366 27326 23418
rect 27378 23366 27390 23418
rect 27442 23366 27454 23418
rect 27506 23366 27518 23418
rect 27570 23366 27576 23418
rect 552 23344 27576 23366
rect 2225 23307 2283 23313
rect 2225 23273 2237 23307
rect 2271 23304 2283 23307
rect 2866 23304 2872 23316
rect 2271 23276 2872 23304
rect 2271 23273 2283 23276
rect 2225 23267 2283 23273
rect 2866 23264 2872 23276
rect 2924 23264 2930 23316
rect 2961 23307 3019 23313
rect 2961 23273 2973 23307
rect 3007 23304 3019 23307
rect 3605 23307 3663 23313
rect 3007 23276 3556 23304
rect 3007 23273 3019 23276
rect 2961 23267 3019 23273
rect 2774 23196 2780 23248
rect 2832 23236 2838 23248
rect 3329 23239 3387 23245
rect 3329 23236 3341 23239
rect 2832 23208 3341 23236
rect 2832 23196 2838 23208
rect 3329 23205 3341 23208
rect 3375 23205 3387 23239
rect 3329 23199 3387 23205
rect 1118 23177 1124 23180
rect 1112 23168 1124 23177
rect 1079 23140 1124 23168
rect 1112 23131 1124 23140
rect 1118 23128 1124 23131
rect 1176 23128 1182 23180
rect 2501 23171 2559 23177
rect 2501 23137 2513 23171
rect 2547 23168 2559 23171
rect 2590 23168 2596 23180
rect 2547 23140 2596 23168
rect 2547 23137 2559 23140
rect 2501 23131 2559 23137
rect 2590 23128 2596 23140
rect 2648 23128 2654 23180
rect 3050 23128 3056 23180
rect 3108 23128 3114 23180
rect 3237 23171 3295 23177
rect 3237 23137 3249 23171
rect 3283 23137 3295 23171
rect 3237 23131 3295 23137
rect 3421 23171 3479 23177
rect 3421 23137 3433 23171
rect 3467 23137 3479 23171
rect 3528 23168 3556 23276
rect 3605 23273 3617 23307
rect 3651 23304 3663 23307
rect 3786 23304 3792 23316
rect 3651 23276 3792 23304
rect 3651 23273 3663 23276
rect 3605 23267 3663 23273
rect 3786 23264 3792 23276
rect 3844 23264 3850 23316
rect 4065 23307 4123 23313
rect 4065 23273 4077 23307
rect 4111 23304 4123 23307
rect 5074 23304 5080 23316
rect 4111 23276 5080 23304
rect 4111 23273 4123 23276
rect 4065 23267 4123 23273
rect 5074 23264 5080 23276
rect 5132 23264 5138 23316
rect 6454 23264 6460 23316
rect 6512 23264 6518 23316
rect 7558 23304 7564 23316
rect 6739 23276 7564 23304
rect 4154 23196 4160 23248
rect 4212 23236 4218 23248
rect 4212 23208 4292 23236
rect 4212 23196 4218 23208
rect 3694 23168 3700 23180
rect 3528 23140 3700 23168
rect 3421 23131 3479 23137
rect 842 23060 848 23112
rect 900 23060 906 23112
rect 3252 23032 3280 23131
rect 3326 23060 3332 23112
rect 3384 23100 3390 23112
rect 3436 23100 3464 23131
rect 3694 23128 3700 23140
rect 3752 23168 3758 23180
rect 4264 23177 4292 23208
rect 6086 23196 6092 23248
rect 6144 23236 6150 23248
rect 6739 23236 6767 23276
rect 7558 23264 7564 23276
rect 7616 23264 7622 23316
rect 7653 23307 7711 23313
rect 7653 23273 7665 23307
rect 7699 23304 7711 23307
rect 8570 23304 8576 23316
rect 7699 23276 8576 23304
rect 7699 23273 7711 23276
rect 7653 23267 7711 23273
rect 8570 23264 8576 23276
rect 8628 23264 8634 23316
rect 8680 23276 8984 23304
rect 6914 23236 6920 23248
rect 6144 23208 6767 23236
rect 6840 23208 6920 23236
rect 6144 23196 6150 23208
rect 4249 23171 4307 23177
rect 3752 23140 4200 23168
rect 3752 23128 3758 23140
rect 3384 23072 3464 23100
rect 3384 23060 3390 23072
rect 3602 23060 3608 23112
rect 3660 23100 3666 23112
rect 4172 23109 4200 23140
rect 4249 23137 4261 23171
rect 4295 23137 4307 23171
rect 4249 23131 4307 23137
rect 4338 23128 4344 23180
rect 4396 23168 4402 23180
rect 4525 23171 4583 23177
rect 4525 23168 4537 23171
rect 4396 23140 4537 23168
rect 4396 23128 4402 23140
rect 4525 23137 4537 23140
rect 4571 23137 4583 23171
rect 4525 23131 4583 23137
rect 4617 23171 4675 23177
rect 4617 23137 4629 23171
rect 4663 23137 4675 23171
rect 4617 23131 4675 23137
rect 4065 23103 4123 23109
rect 4065 23100 4077 23103
rect 3660 23072 4077 23100
rect 3660 23060 3666 23072
rect 4065 23069 4077 23072
rect 4111 23069 4123 23103
rect 4065 23063 4123 23069
rect 4157 23103 4215 23109
rect 4157 23069 4169 23103
rect 4203 23069 4215 23103
rect 4157 23063 4215 23069
rect 3510 23032 3516 23044
rect 2792 23004 3516 23032
rect 2792 22973 2820 23004
rect 3510 22992 3516 23004
rect 3568 22992 3574 23044
rect 4080 23032 4108 23063
rect 4430 23060 4436 23112
rect 4488 23060 4494 23112
rect 4632 23032 4660 23131
rect 4798 23128 4804 23180
rect 4856 23128 4862 23180
rect 5902 23128 5908 23180
rect 5960 23128 5966 23180
rect 6178 23128 6184 23180
rect 6236 23128 6242 23180
rect 6656 23177 6684 23208
rect 6641 23171 6699 23177
rect 6641 23137 6653 23171
rect 6687 23137 6699 23171
rect 6641 23131 6699 23137
rect 6730 23128 6736 23180
rect 6788 23128 6794 23180
rect 6840 23177 6868 23208
rect 6914 23196 6920 23208
rect 6972 23236 6978 23248
rect 7285 23239 7343 23245
rect 7285 23236 7297 23239
rect 6972 23208 7297 23236
rect 6972 23196 6978 23208
rect 7285 23205 7297 23208
rect 7331 23205 7343 23239
rect 7285 23199 7343 23205
rect 7377 23239 7435 23245
rect 7377 23205 7389 23239
rect 7423 23236 7435 23239
rect 8294 23236 8300 23248
rect 7423 23208 8300 23236
rect 7423 23205 7435 23208
rect 7377 23199 7435 23205
rect 8294 23196 8300 23208
rect 8352 23236 8358 23248
rect 8680 23236 8708 23276
rect 8352 23208 8708 23236
rect 8352 23196 8358 23208
rect 8754 23196 8760 23248
rect 8812 23236 8818 23248
rect 8858 23239 8916 23245
rect 8858 23236 8870 23239
rect 8812 23208 8870 23236
rect 8812 23196 8818 23208
rect 8858 23205 8870 23208
rect 8904 23205 8916 23239
rect 8956 23236 8984 23276
rect 9950 23264 9956 23316
rect 10008 23264 10014 23316
rect 12710 23304 12716 23316
rect 11440 23276 12716 23304
rect 11440 23236 11468 23276
rect 12710 23264 12716 23276
rect 12768 23264 12774 23316
rect 12805 23307 12863 23313
rect 12805 23273 12817 23307
rect 12851 23304 12863 23307
rect 13722 23304 13728 23316
rect 12851 23276 13728 23304
rect 12851 23273 12863 23276
rect 12805 23267 12863 23273
rect 13722 23264 13728 23276
rect 13780 23304 13786 23316
rect 14737 23307 14795 23313
rect 14737 23304 14749 23307
rect 13780 23276 14749 23304
rect 13780 23264 13786 23276
rect 14737 23273 14749 23276
rect 14783 23273 14795 23307
rect 14737 23267 14795 23273
rect 15010 23264 15016 23316
rect 15068 23304 15074 23316
rect 16666 23304 16672 23316
rect 15068 23276 16672 23304
rect 15068 23264 15074 23276
rect 16666 23264 16672 23276
rect 16724 23264 16730 23316
rect 16850 23264 16856 23316
rect 16908 23304 16914 23316
rect 17037 23307 17095 23313
rect 17037 23304 17049 23307
rect 16908 23276 17049 23304
rect 16908 23264 16914 23276
rect 17037 23273 17049 23276
rect 17083 23273 17095 23307
rect 17037 23267 17095 23273
rect 17497 23307 17555 23313
rect 17497 23273 17509 23307
rect 17543 23304 17555 23307
rect 17586 23304 17592 23316
rect 17543 23276 17592 23304
rect 17543 23273 17555 23276
rect 17497 23267 17555 23273
rect 17586 23264 17592 23276
rect 17644 23264 17650 23316
rect 18322 23264 18328 23316
rect 18380 23304 18386 23316
rect 18417 23307 18475 23313
rect 18417 23304 18429 23307
rect 18380 23276 18429 23304
rect 18380 23264 18386 23276
rect 18417 23273 18429 23276
rect 18463 23273 18475 23307
rect 18417 23267 18475 23273
rect 18874 23264 18880 23316
rect 18932 23264 18938 23316
rect 19613 23307 19671 23313
rect 19613 23273 19625 23307
rect 19659 23273 19671 23307
rect 19613 23267 19671 23273
rect 8956 23208 11468 23236
rect 8858 23199 8916 23205
rect 11790 23196 11796 23248
rect 11848 23196 11854 23248
rect 12161 23239 12219 23245
rect 12161 23205 12173 23239
rect 12207 23236 12219 23239
rect 12526 23236 12532 23248
rect 12207 23208 12532 23236
rect 12207 23205 12219 23208
rect 12161 23199 12219 23205
rect 12526 23196 12532 23208
rect 12584 23196 12590 23248
rect 13624 23239 13682 23245
rect 13624 23205 13636 23239
rect 13670 23236 13682 23239
rect 14182 23236 14188 23248
rect 13670 23208 14188 23236
rect 13670 23205 13682 23208
rect 13624 23199 13682 23205
rect 14182 23196 14188 23208
rect 14240 23196 14246 23248
rect 14550 23196 14556 23248
rect 14608 23236 14614 23248
rect 15028 23236 15056 23264
rect 16574 23236 16580 23248
rect 14608 23208 15056 23236
rect 15672 23208 16580 23236
rect 14608 23196 14614 23208
rect 6825 23171 6883 23177
rect 6825 23137 6837 23171
rect 6871 23137 6883 23171
rect 6825 23131 6883 23137
rect 6270 23060 6276 23112
rect 6328 23100 6334 23112
rect 6840 23100 6868 23131
rect 7006 23128 7012 23180
rect 7064 23128 7070 23180
rect 7098 23128 7104 23180
rect 7156 23128 7162 23180
rect 7469 23171 7527 23177
rect 7469 23137 7481 23171
rect 7515 23168 7527 23171
rect 7558 23168 7564 23180
rect 7515 23140 7564 23168
rect 7515 23137 7527 23140
rect 7469 23131 7527 23137
rect 7558 23128 7564 23140
rect 7616 23128 7622 23180
rect 9125 23171 9183 23177
rect 7668 23140 9076 23168
rect 6328 23072 6868 23100
rect 6328 23060 6334 23072
rect 4080 23004 4660 23032
rect 6638 22992 6644 23044
rect 6696 23032 6702 23044
rect 7668 23032 7696 23140
rect 9048 23100 9076 23140
rect 9125 23137 9137 23171
rect 9171 23168 9183 23171
rect 9490 23168 9496 23180
rect 9171 23140 9496 23168
rect 9171 23137 9183 23140
rect 9125 23131 9183 23137
rect 9490 23128 9496 23140
rect 9548 23128 9554 23180
rect 10134 23128 10140 23180
rect 10192 23128 10198 23180
rect 10318 23128 10324 23180
rect 10376 23128 10382 23180
rect 10413 23171 10471 23177
rect 10413 23137 10425 23171
rect 10459 23137 10471 23171
rect 10413 23131 10471 23137
rect 9048 23072 9628 23100
rect 6696 23004 7696 23032
rect 7745 23035 7803 23041
rect 6696 22992 6702 23004
rect 7745 23001 7757 23035
rect 7791 23032 7803 23035
rect 7834 23032 7840 23044
rect 7791 23004 7840 23032
rect 7791 23001 7803 23004
rect 7745 22995 7803 23001
rect 7834 22992 7840 23004
rect 7892 22992 7898 23044
rect 9600 23032 9628 23072
rect 9674 23060 9680 23112
rect 9732 23100 9738 23112
rect 10042 23100 10048 23112
rect 9732 23072 10048 23100
rect 9732 23060 9738 23072
rect 10042 23060 10048 23072
rect 10100 23100 10106 23112
rect 10428 23100 10456 23131
rect 11882 23128 11888 23180
rect 11940 23168 11946 23180
rect 11977 23171 12035 23177
rect 11977 23168 11989 23171
rect 11940 23140 11989 23168
rect 11940 23128 11946 23140
rect 11977 23137 11989 23140
rect 12023 23137 12035 23171
rect 11977 23131 12035 23137
rect 12066 23128 12072 23180
rect 12124 23168 12130 23180
rect 12253 23171 12311 23177
rect 12253 23168 12265 23171
rect 12124 23140 12265 23168
rect 12124 23128 12130 23140
rect 12253 23137 12265 23140
rect 12299 23137 12311 23171
rect 12253 23131 12311 23137
rect 12342 23128 12348 23180
rect 12400 23168 12406 23180
rect 12400 23128 12434 23168
rect 12894 23128 12900 23180
rect 12952 23128 12958 23180
rect 14366 23168 14372 23180
rect 13096 23140 14372 23168
rect 11422 23100 11428 23112
rect 10100 23072 10456 23100
rect 11265 23072 11428 23100
rect 10100 23060 10106 23072
rect 11265 23032 11293 23072
rect 11422 23060 11428 23072
rect 11480 23060 11486 23112
rect 11514 23060 11520 23112
rect 11572 23100 11578 23112
rect 12406 23100 12434 23128
rect 12713 23103 12771 23109
rect 12713 23100 12725 23103
rect 11572 23072 12725 23100
rect 11572 23060 11578 23072
rect 12713 23069 12725 23072
rect 12759 23100 12771 23103
rect 13096 23100 13124 23140
rect 14366 23128 14372 23140
rect 14424 23128 14430 23180
rect 15672 23177 15700 23208
rect 16574 23196 16580 23208
rect 16632 23196 16638 23248
rect 17405 23239 17463 23245
rect 17405 23205 17417 23239
rect 17451 23236 17463 23239
rect 17678 23236 17684 23248
rect 17451 23208 17684 23236
rect 17451 23205 17463 23208
rect 17405 23199 17463 23205
rect 15473 23171 15531 23177
rect 15473 23137 15485 23171
rect 15519 23137 15531 23171
rect 15473 23131 15531 23137
rect 15657 23171 15715 23177
rect 15657 23137 15669 23171
rect 15703 23137 15715 23171
rect 15657 23131 15715 23137
rect 12759 23072 13124 23100
rect 13357 23103 13415 23109
rect 12759 23069 12771 23072
rect 12713 23063 12771 23069
rect 13357 23069 13369 23103
rect 13403 23069 13415 23103
rect 13357 23063 13415 23069
rect 9600 23004 11293 23032
rect 11330 22992 11336 23044
rect 11388 23032 11394 23044
rect 12342 23032 12348 23044
rect 11388 23004 12348 23032
rect 11388 22992 11394 23004
rect 12342 22992 12348 23004
rect 12400 23032 12406 23044
rect 13372 23032 13400 23063
rect 12400 23004 13400 23032
rect 15488 23032 15516 23131
rect 15746 23128 15752 23180
rect 15804 23128 15810 23180
rect 16298 23128 16304 23180
rect 16356 23168 16362 23180
rect 16485 23171 16543 23177
rect 16485 23168 16497 23171
rect 16356 23140 16497 23168
rect 16356 23128 16362 23140
rect 16485 23137 16497 23140
rect 16531 23168 16543 23171
rect 17420 23168 17448 23199
rect 17678 23196 17684 23208
rect 17736 23196 17742 23248
rect 19628 23236 19656 23267
rect 20990 23264 20996 23316
rect 21048 23304 21054 23316
rect 21269 23307 21327 23313
rect 21269 23304 21281 23307
rect 21048 23276 21281 23304
rect 21048 23264 21054 23276
rect 21269 23273 21281 23276
rect 21315 23273 21327 23307
rect 21269 23267 21327 23273
rect 21910 23264 21916 23316
rect 21968 23264 21974 23316
rect 23290 23304 23296 23316
rect 22066 23276 23296 23304
rect 19950 23239 20008 23245
rect 19950 23236 19962 23239
rect 19628 23208 19962 23236
rect 19950 23205 19962 23208
rect 19996 23205 20008 23239
rect 22066 23236 22094 23276
rect 19950 23199 20008 23205
rect 21836 23208 22094 23236
rect 16531 23140 17448 23168
rect 16531 23137 16543 23140
rect 16485 23131 16543 23137
rect 18138 23128 18144 23180
rect 18196 23168 18202 23180
rect 18782 23168 18788 23180
rect 18196 23140 18788 23168
rect 18196 23128 18202 23140
rect 18782 23128 18788 23140
rect 18840 23128 18846 23180
rect 19429 23171 19487 23177
rect 19429 23137 19441 23171
rect 19475 23168 19487 23171
rect 19610 23168 19616 23180
rect 19475 23140 19616 23168
rect 19475 23137 19487 23140
rect 19429 23131 19487 23137
rect 19610 23128 19616 23140
rect 19668 23128 19674 23180
rect 21836 23177 21864 23208
rect 22186 23196 22192 23248
rect 22244 23196 22250 23248
rect 21453 23171 21511 23177
rect 21453 23168 21465 23171
rect 21100 23140 21465 23168
rect 15933 23103 15991 23109
rect 15933 23069 15945 23103
rect 15979 23100 15991 23103
rect 16577 23103 16635 23109
rect 16577 23100 16589 23103
rect 15979 23072 16589 23100
rect 15979 23069 15991 23072
rect 15933 23063 15991 23069
rect 16577 23069 16589 23072
rect 16623 23069 16635 23103
rect 16577 23063 16635 23069
rect 16669 23103 16727 23109
rect 16669 23069 16681 23103
rect 16715 23069 16727 23103
rect 16669 23063 16727 23069
rect 17681 23103 17739 23109
rect 17681 23069 17693 23103
rect 17727 23100 17739 23103
rect 19061 23103 19119 23109
rect 19061 23100 19073 23103
rect 17727 23072 19073 23100
rect 17727 23069 17739 23072
rect 17681 23063 17739 23069
rect 19061 23069 19073 23072
rect 19107 23100 19119 23103
rect 19334 23100 19340 23112
rect 19107 23072 19340 23100
rect 19107 23069 19119 23072
rect 19061 23063 19119 23069
rect 16117 23035 16175 23041
rect 16117 23032 16129 23035
rect 15488 23004 16129 23032
rect 12400 22992 12406 23004
rect 16117 23001 16129 23004
rect 16163 23001 16175 23035
rect 16117 22995 16175 23001
rect 16390 22992 16396 23044
rect 16448 23032 16454 23044
rect 16684 23032 16712 23063
rect 19334 23060 19340 23072
rect 19392 23060 19398 23112
rect 19705 23103 19763 23109
rect 19705 23069 19717 23103
rect 19751 23069 19763 23103
rect 19705 23063 19763 23069
rect 19720 23032 19748 23063
rect 16448 23004 16712 23032
rect 18892 23004 19748 23032
rect 16448 22992 16454 23004
rect 18892 22976 18920 23004
rect 20898 22992 20904 23044
rect 20956 23032 20962 23044
rect 21100 23041 21128 23140
rect 21453 23137 21465 23140
rect 21499 23137 21511 23171
rect 21453 23131 21511 23137
rect 21545 23171 21603 23177
rect 21545 23137 21557 23171
rect 21591 23137 21603 23171
rect 21545 23131 21603 23137
rect 21821 23171 21879 23177
rect 21821 23137 21833 23171
rect 21867 23137 21879 23171
rect 21821 23131 21879 23137
rect 21560 23100 21588 23131
rect 22094 23128 22100 23180
rect 22152 23128 22158 23180
rect 22278 23128 22284 23180
rect 22336 23128 22342 23180
rect 22480 23177 22508 23276
rect 23290 23264 23296 23276
rect 23348 23264 23354 23316
rect 24670 23264 24676 23316
rect 24728 23264 24734 23316
rect 26421 23307 26479 23313
rect 26421 23273 26433 23307
rect 26467 23304 26479 23307
rect 26694 23304 26700 23316
rect 26467 23276 26700 23304
rect 26467 23273 26479 23276
rect 26421 23267 26479 23273
rect 26694 23264 26700 23276
rect 26752 23264 26758 23316
rect 24305 23239 24363 23245
rect 24305 23205 24317 23239
rect 24351 23205 24363 23239
rect 24305 23199 24363 23205
rect 24521 23239 24579 23245
rect 24521 23205 24533 23239
rect 24567 23236 24579 23239
rect 25130 23236 25136 23248
rect 24567 23208 25136 23236
rect 24567 23205 24579 23208
rect 24521 23199 24579 23205
rect 22465 23171 22523 23177
rect 22465 23137 22477 23171
rect 22511 23137 22523 23171
rect 22465 23131 22523 23137
rect 23842 23128 23848 23180
rect 23900 23128 23906 23180
rect 24320 23168 24348 23199
rect 25130 23196 25136 23208
rect 25188 23196 25194 23248
rect 25590 23168 25596 23180
rect 24320 23140 25596 23168
rect 25590 23128 25596 23140
rect 25648 23128 25654 23180
rect 21634 23100 21640 23112
rect 21560 23072 21640 23100
rect 21634 23060 21640 23072
rect 21692 23100 21698 23112
rect 23753 23103 23811 23109
rect 23753 23100 23765 23103
rect 21692 23072 23765 23100
rect 21692 23060 21698 23072
rect 23753 23069 23765 23072
rect 23799 23069 23811 23103
rect 23753 23063 23811 23069
rect 24578 23060 24584 23112
rect 24636 23100 24642 23112
rect 25038 23100 25044 23112
rect 24636 23072 25044 23100
rect 24636 23060 24642 23072
rect 25038 23060 25044 23072
rect 25096 23060 25102 23112
rect 26878 23060 26884 23112
rect 26936 23100 26942 23112
rect 26973 23103 27031 23109
rect 26973 23100 26985 23103
rect 26936 23072 26985 23100
rect 26936 23060 26942 23072
rect 26973 23069 26985 23072
rect 27019 23069 27031 23103
rect 26973 23063 27031 23069
rect 21085 23035 21143 23041
rect 21085 23032 21097 23035
rect 20956 23004 21097 23032
rect 20956 22992 20962 23004
rect 21085 23001 21097 23004
rect 21131 23001 21143 23035
rect 21085 22995 21143 23001
rect 2777 22967 2835 22973
rect 2777 22933 2789 22967
rect 2823 22933 2835 22967
rect 2777 22927 2835 22933
rect 4522 22924 4528 22976
rect 4580 22964 4586 22976
rect 4709 22967 4767 22973
rect 4709 22964 4721 22967
rect 4580 22936 4721 22964
rect 4580 22924 4586 22936
rect 4709 22933 4721 22936
rect 4755 22933 4767 22967
rect 4709 22927 4767 22933
rect 9122 22924 9128 22976
rect 9180 22964 9186 22976
rect 11698 22964 11704 22976
rect 9180 22936 11704 22964
rect 9180 22924 9186 22936
rect 11698 22924 11704 22936
rect 11756 22924 11762 22976
rect 11790 22924 11796 22976
rect 11848 22964 11854 22976
rect 12986 22964 12992 22976
rect 11848 22936 12992 22964
rect 11848 22924 11854 22936
rect 12986 22924 12992 22936
rect 13044 22924 13050 22976
rect 13170 22924 13176 22976
rect 13228 22964 13234 22976
rect 13265 22967 13323 22973
rect 13265 22964 13277 22967
rect 13228 22936 13277 22964
rect 13228 22924 13234 22936
rect 13265 22933 13277 22936
rect 13311 22933 13323 22967
rect 13265 22927 13323 22933
rect 15289 22967 15347 22973
rect 15289 22933 15301 22967
rect 15335 22964 15347 22967
rect 15470 22964 15476 22976
rect 15335 22936 15476 22964
rect 15335 22933 15347 22936
rect 15289 22927 15347 22933
rect 15470 22924 15476 22936
rect 15528 22924 15534 22976
rect 18874 22924 18880 22976
rect 18932 22924 18938 22976
rect 20346 22924 20352 22976
rect 20404 22964 20410 22976
rect 21729 22967 21787 22973
rect 21729 22964 21741 22967
rect 20404 22936 21741 22964
rect 20404 22924 20410 22936
rect 21729 22933 21741 22936
rect 21775 22964 21787 22967
rect 22278 22964 22284 22976
rect 21775 22936 22284 22964
rect 21775 22933 21787 22936
rect 21729 22927 21787 22933
rect 22278 22924 22284 22936
rect 22336 22924 22342 22976
rect 24486 22924 24492 22976
rect 24544 22924 24550 22976
rect 552 22874 27416 22896
rect 552 22822 3756 22874
rect 3808 22822 3820 22874
rect 3872 22822 3884 22874
rect 3936 22822 3948 22874
rect 4000 22822 4012 22874
rect 4064 22822 10472 22874
rect 10524 22822 10536 22874
rect 10588 22822 10600 22874
rect 10652 22822 10664 22874
rect 10716 22822 10728 22874
rect 10780 22822 17188 22874
rect 17240 22822 17252 22874
rect 17304 22822 17316 22874
rect 17368 22822 17380 22874
rect 17432 22822 17444 22874
rect 17496 22822 23904 22874
rect 23956 22822 23968 22874
rect 24020 22822 24032 22874
rect 24084 22822 24096 22874
rect 24148 22822 24160 22874
rect 24212 22822 27416 22874
rect 552 22800 27416 22822
rect 2314 22720 2320 22772
rect 2372 22760 2378 22772
rect 2409 22763 2467 22769
rect 2409 22760 2421 22763
rect 2372 22732 2421 22760
rect 2372 22720 2378 22732
rect 2409 22729 2421 22732
rect 2455 22729 2467 22763
rect 2409 22723 2467 22729
rect 3326 22720 3332 22772
rect 3384 22760 3390 22772
rect 3513 22763 3571 22769
rect 3513 22760 3525 22763
rect 3384 22732 3525 22760
rect 3384 22720 3390 22732
rect 3513 22729 3525 22732
rect 3559 22729 3571 22763
rect 3513 22723 3571 22729
rect 3528 22692 3556 22723
rect 3602 22720 3608 22772
rect 3660 22760 3666 22772
rect 3697 22763 3755 22769
rect 3697 22760 3709 22763
rect 3660 22732 3709 22760
rect 3660 22720 3666 22732
rect 3697 22729 3709 22732
rect 3743 22729 3755 22763
rect 3697 22723 3755 22729
rect 5258 22720 5264 22772
rect 5316 22720 5322 22772
rect 7193 22763 7251 22769
rect 7193 22729 7205 22763
rect 7239 22760 7251 22763
rect 9122 22760 9128 22772
rect 7239 22732 9128 22760
rect 7239 22729 7251 22732
rect 7193 22723 7251 22729
rect 9122 22720 9128 22732
rect 9180 22720 9186 22772
rect 9766 22720 9772 22772
rect 9824 22760 9830 22772
rect 9861 22763 9919 22769
rect 9861 22760 9873 22763
rect 9824 22732 9873 22760
rect 9824 22720 9830 22732
rect 9861 22729 9873 22732
rect 9907 22729 9919 22763
rect 9861 22723 9919 22729
rect 11977 22763 12035 22769
rect 11977 22729 11989 22763
rect 12023 22729 12035 22763
rect 11977 22723 12035 22729
rect 13357 22763 13415 22769
rect 13357 22729 13369 22763
rect 13403 22760 13415 22763
rect 14274 22760 14280 22772
rect 13403 22732 14280 22760
rect 13403 22729 13415 22732
rect 13357 22723 13415 22729
rect 3528 22664 3648 22692
rect 3620 22624 3648 22664
rect 4614 22652 4620 22704
rect 4672 22692 4678 22704
rect 5077 22695 5135 22701
rect 5077 22692 5089 22695
rect 4672 22664 5089 22692
rect 4672 22652 4678 22664
rect 5077 22661 5089 22664
rect 5123 22661 5135 22695
rect 5077 22655 5135 22661
rect 7098 22652 7104 22704
rect 7156 22692 7162 22704
rect 7469 22695 7527 22701
rect 7469 22692 7481 22695
rect 7156 22664 7481 22692
rect 7156 22652 7162 22664
rect 7469 22661 7481 22664
rect 7515 22661 7527 22695
rect 7469 22655 7527 22661
rect 5166 22624 5172 22636
rect 3620 22596 5172 22624
rect 5166 22584 5172 22596
rect 5224 22584 5230 22636
rect 5350 22584 5356 22636
rect 5408 22584 5414 22636
rect 7558 22584 7564 22636
rect 7616 22624 7622 22636
rect 9876 22624 9904 22723
rect 11992 22692 12020 22723
rect 14274 22720 14280 22732
rect 14332 22720 14338 22772
rect 16574 22720 16580 22772
rect 16632 22720 16638 22772
rect 19610 22720 19616 22772
rect 19668 22720 19674 22772
rect 26878 22720 26884 22772
rect 26936 22720 26942 22772
rect 11348 22664 12020 22692
rect 11348 22636 11376 22664
rect 12986 22652 12992 22704
rect 13044 22692 13050 22704
rect 13817 22695 13875 22701
rect 13817 22692 13829 22695
rect 13044 22664 13829 22692
rect 13044 22652 13050 22664
rect 13817 22661 13829 22664
rect 13863 22661 13875 22695
rect 13817 22655 13875 22661
rect 14369 22695 14427 22701
rect 14369 22661 14381 22695
rect 14415 22692 14427 22695
rect 14458 22692 14464 22704
rect 14415 22664 14464 22692
rect 14415 22661 14427 22664
rect 14369 22655 14427 22661
rect 14458 22652 14464 22664
rect 14516 22652 14522 22704
rect 16390 22652 16396 22704
rect 16448 22692 16454 22704
rect 16669 22695 16727 22701
rect 16669 22692 16681 22695
rect 16448 22664 16681 22692
rect 16448 22652 16454 22664
rect 16669 22661 16681 22664
rect 16715 22661 16727 22695
rect 16669 22655 16727 22661
rect 17497 22695 17555 22701
rect 17497 22661 17509 22695
rect 17543 22692 17555 22695
rect 17543 22664 19380 22692
rect 17543 22661 17555 22664
rect 17497 22655 17555 22661
rect 19352 22636 19380 22664
rect 10689 22627 10747 22633
rect 10689 22624 10701 22627
rect 7616 22596 8140 22624
rect 9876 22596 10701 22624
rect 7616 22584 7622 22596
rect 2590 22516 2596 22568
rect 2648 22516 2654 22568
rect 2685 22559 2743 22565
rect 2685 22525 2697 22559
rect 2731 22556 2743 22559
rect 2866 22556 2872 22568
rect 2731 22528 2872 22556
rect 2731 22525 2743 22528
rect 2685 22519 2743 22525
rect 2866 22516 2872 22528
rect 2924 22556 2930 22568
rect 3237 22559 3295 22565
rect 3237 22556 3249 22559
rect 2924 22528 3249 22556
rect 2924 22516 2930 22528
rect 3237 22525 3249 22528
rect 3283 22525 3295 22559
rect 3237 22519 3295 22525
rect 4522 22516 4528 22568
rect 4580 22516 4586 22568
rect 4801 22559 4859 22565
rect 4801 22525 4813 22559
rect 4847 22556 4859 22559
rect 4982 22556 4988 22568
rect 4847 22528 4988 22556
rect 4847 22525 4859 22528
rect 4801 22519 4859 22525
rect 4982 22516 4988 22528
rect 5040 22556 5046 22568
rect 5258 22556 5264 22568
rect 5040 22528 5264 22556
rect 5040 22516 5046 22528
rect 5258 22516 5264 22528
rect 5316 22516 5322 22568
rect 5445 22559 5503 22565
rect 5445 22525 5457 22559
rect 5491 22525 5503 22559
rect 5445 22519 5503 22525
rect 5537 22559 5595 22565
rect 5537 22525 5549 22559
rect 5583 22556 5595 22559
rect 5626 22556 5632 22568
rect 5583 22528 5632 22556
rect 5583 22525 5595 22528
rect 5537 22519 5595 22525
rect 2961 22491 3019 22497
rect 2961 22457 2973 22491
rect 3007 22488 3019 22491
rect 3142 22488 3148 22500
rect 3007 22460 3148 22488
rect 3007 22457 3019 22460
rect 2961 22451 3019 22457
rect 3142 22448 3148 22460
rect 3200 22448 3206 22500
rect 5460 22488 5488 22519
rect 5626 22516 5632 22528
rect 5684 22516 5690 22568
rect 6362 22556 6368 22568
rect 5736 22528 6368 22556
rect 5736 22488 5764 22528
rect 6362 22516 6368 22528
rect 6420 22516 6426 22568
rect 7466 22516 7472 22568
rect 7524 22556 7530 22568
rect 8021 22559 8079 22565
rect 8021 22556 8033 22559
rect 7524 22528 8033 22556
rect 7524 22516 7530 22528
rect 8021 22525 8033 22528
rect 8067 22525 8079 22559
rect 8021 22519 8079 22525
rect 5460 22460 5764 22488
rect 5804 22491 5862 22497
rect 5804 22457 5816 22491
rect 5850 22488 5862 22491
rect 5902 22488 5908 22500
rect 5850 22460 5908 22488
rect 5850 22457 5862 22460
rect 5804 22451 5862 22457
rect 5902 22448 5908 22460
rect 5960 22448 5966 22500
rect 7377 22491 7435 22497
rect 7377 22457 7389 22491
rect 7423 22488 7435 22491
rect 7558 22488 7564 22500
rect 7423 22460 7564 22488
rect 7423 22457 7435 22460
rect 7377 22451 7435 22457
rect 7558 22448 7564 22460
rect 7616 22448 7622 22500
rect 8112 22488 8140 22596
rect 10689 22593 10701 22596
rect 10735 22593 10747 22627
rect 10689 22587 10747 22593
rect 11330 22584 11336 22636
rect 11388 22584 11394 22636
rect 11514 22584 11520 22636
rect 11572 22584 11578 22636
rect 12250 22584 12256 22636
rect 12308 22624 12314 22636
rect 12529 22627 12587 22633
rect 12529 22624 12541 22627
rect 12308 22596 12541 22624
rect 12308 22584 12314 22596
rect 12529 22593 12541 22596
rect 12575 22593 12587 22627
rect 12529 22587 12587 22593
rect 12894 22584 12900 22636
rect 12952 22624 12958 22636
rect 14918 22624 14924 22636
rect 12952 22596 14924 22624
rect 12952 22584 12958 22596
rect 14918 22584 14924 22596
rect 14976 22584 14982 22636
rect 17954 22584 17960 22636
rect 18012 22584 18018 22636
rect 19334 22584 19340 22636
rect 19392 22624 19398 22636
rect 20070 22624 20076 22636
rect 19392 22596 20076 22624
rect 19392 22584 19398 22596
rect 20070 22584 20076 22596
rect 20128 22624 20134 22636
rect 20165 22627 20223 22633
rect 20165 22624 20177 22627
rect 20128 22596 20177 22624
rect 20128 22584 20134 22596
rect 20165 22593 20177 22596
rect 20211 22593 20223 22627
rect 25038 22624 25044 22636
rect 20165 22587 20223 22593
rect 22066 22596 25044 22624
rect 8481 22559 8539 22565
rect 8481 22525 8493 22559
rect 8527 22556 8539 22559
rect 8527 22528 8892 22556
rect 8527 22525 8539 22528
rect 8481 22519 8539 22525
rect 8864 22500 8892 22528
rect 11882 22516 11888 22568
rect 11940 22556 11946 22568
rect 12161 22559 12219 22565
rect 12161 22556 12173 22559
rect 11940 22528 12173 22556
rect 11940 22516 11946 22528
rect 12161 22525 12173 22528
rect 12207 22525 12219 22559
rect 12161 22519 12219 22525
rect 12986 22516 12992 22568
rect 13044 22516 13050 22568
rect 13170 22516 13176 22568
rect 13228 22516 13234 22568
rect 13262 22516 13268 22568
rect 13320 22556 13326 22568
rect 13541 22559 13599 22565
rect 13541 22556 13553 22559
rect 13320 22528 13553 22556
rect 13320 22516 13326 22528
rect 13541 22525 13553 22528
rect 13587 22525 13599 22559
rect 13541 22519 13599 22525
rect 13725 22559 13783 22565
rect 13725 22525 13737 22559
rect 13771 22556 13783 22559
rect 14734 22556 14740 22568
rect 13771 22528 14740 22556
rect 13771 22525 13783 22528
rect 13725 22519 13783 22525
rect 14734 22516 14740 22528
rect 14792 22516 14798 22568
rect 15197 22559 15255 22565
rect 15197 22525 15209 22559
rect 15243 22556 15255 22559
rect 15286 22556 15292 22568
rect 15243 22528 15292 22556
rect 15243 22525 15255 22528
rect 15197 22519 15255 22525
rect 15286 22516 15292 22528
rect 15344 22516 15350 22568
rect 15470 22565 15476 22568
rect 15464 22556 15476 22565
rect 15431 22528 15476 22556
rect 15464 22519 15476 22528
rect 15470 22516 15476 22519
rect 15528 22516 15534 22568
rect 17129 22559 17187 22565
rect 17129 22556 17141 22559
rect 16868 22528 17141 22556
rect 8754 22497 8760 22500
rect 8112 22460 8600 22488
rect 2682 22380 2688 22432
rect 2740 22420 2746 22432
rect 2777 22423 2835 22429
rect 2777 22420 2789 22423
rect 2740 22392 2789 22420
rect 2740 22380 2746 22392
rect 2777 22389 2789 22392
rect 2823 22389 2835 22423
rect 2777 22383 2835 22389
rect 4246 22380 4252 22432
rect 4304 22420 4310 22432
rect 4617 22423 4675 22429
rect 4617 22420 4629 22423
rect 4304 22392 4629 22420
rect 4304 22380 4310 22392
rect 4617 22389 4629 22392
rect 4663 22389 4675 22423
rect 4617 22383 4675 22389
rect 4985 22423 5043 22429
rect 4985 22389 4997 22423
rect 5031 22420 5043 22423
rect 5718 22420 5724 22432
rect 5031 22392 5724 22420
rect 5031 22389 5043 22392
rect 4985 22383 5043 22389
rect 5718 22380 5724 22392
rect 5776 22380 5782 22432
rect 6914 22380 6920 22432
rect 6972 22380 6978 22432
rect 7006 22380 7012 22432
rect 7064 22380 7070 22432
rect 7177 22423 7235 22429
rect 7177 22389 7189 22423
rect 7223 22420 7235 22423
rect 8478 22420 8484 22432
rect 7223 22392 8484 22420
rect 7223 22389 7235 22392
rect 7177 22383 7235 22389
rect 8478 22380 8484 22392
rect 8536 22380 8542 22432
rect 8572 22420 8600 22460
rect 8748 22451 8760 22497
rect 8754 22448 8760 22451
rect 8812 22448 8818 22500
rect 8846 22448 8852 22500
rect 8904 22448 8910 22500
rect 11790 22488 11796 22500
rect 9646 22460 11796 22488
rect 9646 22420 9674 22460
rect 11790 22448 11796 22460
rect 11848 22448 11854 22500
rect 13354 22448 13360 22500
rect 13412 22488 13418 22500
rect 16868 22497 16896 22528
rect 17129 22525 17141 22528
rect 17175 22556 17187 22559
rect 17589 22559 17647 22565
rect 17589 22556 17601 22559
rect 17175 22528 17601 22556
rect 17175 22525 17187 22528
rect 17129 22519 17187 22525
rect 17589 22525 17601 22528
rect 17635 22525 17647 22559
rect 17589 22519 17647 22525
rect 17770 22516 17776 22568
rect 17828 22516 17834 22568
rect 22066 22556 22094 22596
rect 17880 22528 22094 22556
rect 14001 22491 14059 22497
rect 14001 22488 14013 22491
rect 13412 22460 14013 22488
rect 13412 22448 13418 22460
rect 14001 22457 14013 22460
rect 14047 22457 14059 22491
rect 14185 22491 14243 22497
rect 14185 22488 14197 22491
rect 14001 22451 14059 22457
rect 14108 22460 14197 22488
rect 8572 22392 9674 22420
rect 10134 22380 10140 22432
rect 10192 22380 10198 22432
rect 10410 22380 10416 22432
rect 10468 22420 10474 22432
rect 10873 22423 10931 22429
rect 10873 22420 10885 22423
rect 10468 22392 10885 22420
rect 10468 22380 10474 22392
rect 10873 22389 10885 22392
rect 10919 22389 10931 22423
rect 10873 22383 10931 22389
rect 11238 22380 11244 22432
rect 11296 22380 11302 22432
rect 12345 22423 12403 22429
rect 12345 22389 12357 22423
rect 12391 22420 12403 22423
rect 12802 22420 12808 22432
rect 12391 22392 12808 22420
rect 12391 22389 12403 22392
rect 12345 22383 12403 22389
rect 12802 22380 12808 22392
rect 12860 22420 12866 22432
rect 14108 22420 14136 22460
rect 14185 22457 14197 22460
rect 14231 22488 14243 22491
rect 16853 22491 16911 22497
rect 16853 22488 16865 22491
rect 14231 22460 16865 22488
rect 14231 22457 14243 22460
rect 14185 22451 14243 22457
rect 16853 22457 16865 22460
rect 16899 22457 16911 22491
rect 16853 22451 16911 22457
rect 16942 22448 16948 22500
rect 17000 22488 17006 22500
rect 17037 22491 17095 22497
rect 17037 22488 17049 22491
rect 17000 22460 17049 22488
rect 17000 22448 17006 22460
rect 17037 22457 17049 22460
rect 17083 22457 17095 22491
rect 17037 22451 17095 22457
rect 17218 22448 17224 22500
rect 17276 22488 17282 22500
rect 17313 22491 17371 22497
rect 17313 22488 17325 22491
rect 17276 22460 17325 22488
rect 17276 22448 17282 22460
rect 17313 22457 17325 22460
rect 17359 22457 17371 22491
rect 17313 22451 17371 22457
rect 12860 22392 14136 22420
rect 12860 22380 12866 22392
rect 15470 22380 15476 22432
rect 15528 22420 15534 22432
rect 17880 22420 17908 22528
rect 22370 22516 22376 22568
rect 22428 22516 22434 22568
rect 22554 22516 22560 22568
rect 22612 22516 22618 22568
rect 22664 22565 22692 22596
rect 25038 22584 25044 22596
rect 25096 22584 25102 22636
rect 25406 22584 25412 22636
rect 25464 22624 25470 22636
rect 25501 22627 25559 22633
rect 25501 22624 25513 22627
rect 25464 22596 25513 22624
rect 25464 22584 25470 22596
rect 25501 22593 25513 22596
rect 25547 22593 25559 22627
rect 25501 22587 25559 22593
rect 22649 22559 22707 22565
rect 22649 22525 22661 22559
rect 22695 22525 22707 22559
rect 22649 22519 22707 22525
rect 22922 22516 22928 22568
rect 22980 22516 22986 22568
rect 23198 22516 23204 22568
rect 23256 22516 23262 22568
rect 23474 22516 23480 22568
rect 23532 22556 23538 22568
rect 25774 22565 25780 22568
rect 23845 22559 23903 22565
rect 23845 22556 23857 22559
rect 23532 22528 23857 22556
rect 23532 22516 23538 22528
rect 23845 22525 23857 22528
rect 23891 22525 23903 22559
rect 25768 22556 25780 22565
rect 25735 22528 25780 22556
rect 23845 22519 23903 22525
rect 25768 22519 25780 22528
rect 25774 22516 25780 22519
rect 25832 22516 25838 22568
rect 19518 22448 19524 22500
rect 19576 22488 19582 22500
rect 19981 22491 20039 22497
rect 19981 22488 19993 22491
rect 19576 22460 19993 22488
rect 19576 22448 19582 22460
rect 19981 22457 19993 22460
rect 20027 22457 20039 22491
rect 19981 22451 20039 22457
rect 20073 22491 20131 22497
rect 20073 22457 20085 22491
rect 20119 22488 20131 22491
rect 20162 22488 20168 22500
rect 20119 22460 20168 22488
rect 20119 22457 20131 22460
rect 20073 22451 20131 22457
rect 20162 22448 20168 22460
rect 20220 22448 20226 22500
rect 15528 22392 17908 22420
rect 15528 22380 15534 22392
rect 22462 22380 22468 22432
rect 22520 22380 22526 22432
rect 22646 22380 22652 22432
rect 22704 22420 22710 22432
rect 22741 22423 22799 22429
rect 22741 22420 22753 22423
rect 22704 22392 22753 22420
rect 22704 22380 22710 22392
rect 22741 22389 22753 22392
rect 22787 22389 22799 22423
rect 22741 22383 22799 22389
rect 23014 22380 23020 22432
rect 23072 22420 23078 22432
rect 23109 22423 23167 22429
rect 23109 22420 23121 22423
rect 23072 22392 23121 22420
rect 23072 22380 23078 22392
rect 23109 22389 23121 22392
rect 23155 22389 23167 22423
rect 23109 22383 23167 22389
rect 23385 22423 23443 22429
rect 23385 22389 23397 22423
rect 23431 22420 23443 22423
rect 23934 22420 23940 22432
rect 23431 22392 23940 22420
rect 23431 22389 23443 22392
rect 23385 22383 23443 22389
rect 23934 22380 23940 22392
rect 23992 22380 23998 22432
rect 24029 22423 24087 22429
rect 24029 22389 24041 22423
rect 24075 22420 24087 22423
rect 24854 22420 24860 22432
rect 24075 22392 24860 22420
rect 24075 22389 24087 22392
rect 24029 22383 24087 22389
rect 24854 22380 24860 22392
rect 24912 22380 24918 22432
rect 552 22330 27576 22352
rect 552 22278 7114 22330
rect 7166 22278 7178 22330
rect 7230 22278 7242 22330
rect 7294 22278 7306 22330
rect 7358 22278 7370 22330
rect 7422 22278 13830 22330
rect 13882 22278 13894 22330
rect 13946 22278 13958 22330
rect 14010 22278 14022 22330
rect 14074 22278 14086 22330
rect 14138 22278 20546 22330
rect 20598 22278 20610 22330
rect 20662 22278 20674 22330
rect 20726 22278 20738 22330
rect 20790 22278 20802 22330
rect 20854 22278 27262 22330
rect 27314 22278 27326 22330
rect 27378 22278 27390 22330
rect 27442 22278 27454 22330
rect 27506 22278 27518 22330
rect 27570 22278 27576 22330
rect 552 22256 27576 22278
rect 3510 22176 3516 22228
rect 3568 22176 3574 22228
rect 4982 22176 4988 22228
rect 5040 22176 5046 22228
rect 5166 22176 5172 22228
rect 5224 22216 5230 22228
rect 7466 22216 7472 22228
rect 5224 22188 7472 22216
rect 5224 22176 5230 22188
rect 7466 22176 7472 22188
rect 7524 22176 7530 22228
rect 8754 22176 8760 22228
rect 8812 22216 8818 22228
rect 9033 22219 9091 22225
rect 9033 22216 9045 22219
rect 8812 22188 9045 22216
rect 8812 22176 8818 22188
rect 9033 22185 9045 22188
rect 9079 22185 9091 22219
rect 9033 22179 9091 22185
rect 9937 22219 9995 22225
rect 9937 22185 9949 22219
rect 9983 22216 9995 22219
rect 10226 22216 10232 22228
rect 9983 22188 10232 22216
rect 9983 22185 9995 22188
rect 9937 22179 9995 22185
rect 10226 22176 10232 22188
rect 10284 22176 10290 22228
rect 13354 22176 13360 22228
rect 13412 22216 13418 22228
rect 14458 22216 14464 22228
rect 13412 22188 14464 22216
rect 13412 22176 13418 22188
rect 14458 22176 14464 22188
rect 14516 22176 14522 22228
rect 16301 22219 16359 22225
rect 16301 22185 16313 22219
rect 16347 22185 16359 22219
rect 16301 22179 16359 22185
rect 1765 22151 1823 22157
rect 1765 22117 1777 22151
rect 1811 22148 1823 22151
rect 3528 22148 3556 22176
rect 1811 22120 2636 22148
rect 3528 22120 6868 22148
rect 1811 22117 1823 22120
rect 1765 22111 1823 22117
rect 2608 22092 2636 22120
rect 1949 22083 2007 22089
rect 1949 22049 1961 22083
rect 1995 22080 2007 22083
rect 2222 22080 2228 22092
rect 1995 22052 2228 22080
rect 1995 22049 2007 22052
rect 1949 22043 2007 22049
rect 2222 22040 2228 22052
rect 2280 22040 2286 22092
rect 2590 22040 2596 22092
rect 2648 22080 2654 22092
rect 3053 22083 3111 22089
rect 3053 22080 3065 22083
rect 2648 22052 3065 22080
rect 2648 22040 2654 22052
rect 3053 22049 3065 22052
rect 3099 22049 3111 22083
rect 3053 22043 3111 22049
rect 4798 22040 4804 22092
rect 4856 22080 4862 22092
rect 4893 22083 4951 22089
rect 4893 22080 4905 22083
rect 4856 22052 4905 22080
rect 4856 22040 4862 22052
rect 4893 22049 4905 22052
rect 4939 22049 4951 22083
rect 4893 22043 4951 22049
rect 5074 22040 5080 22092
rect 5132 22040 5138 22092
rect 5629 22083 5687 22089
rect 5629 22049 5641 22083
rect 5675 22080 5687 22083
rect 6273 22083 6331 22089
rect 6273 22080 6285 22083
rect 5675 22052 6285 22080
rect 5675 22049 5687 22052
rect 5629 22043 5687 22049
rect 6273 22049 6285 22052
rect 6319 22080 6331 22083
rect 6730 22080 6736 22092
rect 6319 22052 6736 22080
rect 6319 22049 6331 22052
rect 6273 22043 6331 22049
rect 6730 22040 6736 22052
rect 6788 22040 6794 22092
rect 6840 22080 6868 22120
rect 9416 22120 9628 22148
rect 9416 22092 9444 22120
rect 6914 22080 6920 22092
rect 6840 22052 6920 22080
rect 6914 22040 6920 22052
rect 6972 22040 6978 22092
rect 8570 22040 8576 22092
rect 8628 22089 8634 22092
rect 8628 22080 8640 22089
rect 9217 22083 9275 22089
rect 8628 22052 8673 22080
rect 8628 22043 8640 22052
rect 9217 22049 9229 22083
rect 9263 22049 9275 22083
rect 9398 22080 9404 22092
rect 9379 22052 9404 22080
rect 9217 22043 9275 22049
rect 8628 22040 8634 22043
rect 3142 21972 3148 22024
rect 3200 22012 3206 22024
rect 3326 22012 3332 22024
rect 3200 21984 3332 22012
rect 3200 21972 3206 21984
rect 3326 21972 3332 21984
rect 3384 21972 3390 22024
rect 5350 21972 5356 22024
rect 5408 21972 5414 22024
rect 6089 22015 6147 22021
rect 6089 21981 6101 22015
rect 6135 22012 6147 22015
rect 6178 22012 6184 22024
rect 6135 21984 6184 22012
rect 6135 21981 6147 21984
rect 6089 21975 6147 21981
rect 6178 21972 6184 21984
rect 6236 22012 6242 22024
rect 7650 22012 7656 22024
rect 6236 21984 7656 22012
rect 6236 21972 6242 21984
rect 7650 21972 7656 21984
rect 7708 21972 7714 22024
rect 8846 21972 8852 22024
rect 8904 21972 8910 22024
rect 9232 22012 9260 22043
rect 9398 22040 9404 22052
rect 9456 22040 9462 22092
rect 9490 22040 9496 22092
rect 9548 22040 9554 22092
rect 9600 22080 9628 22120
rect 10134 22108 10140 22160
rect 10192 22108 10198 22160
rect 12342 22108 12348 22160
rect 12400 22148 12406 22160
rect 13909 22151 13967 22157
rect 12400 22120 13400 22148
rect 12400 22108 12406 22120
rect 9600 22052 9904 22080
rect 9232 21984 9812 22012
rect 5534 21904 5540 21956
rect 5592 21944 5598 21956
rect 9784 21953 9812 21984
rect 9769 21947 9827 21953
rect 5592 21916 7972 21944
rect 5592 21904 5598 21916
rect 1394 21836 1400 21888
rect 1452 21876 1458 21888
rect 1581 21879 1639 21885
rect 1581 21876 1593 21879
rect 1452 21848 1593 21876
rect 1452 21836 1458 21848
rect 1581 21845 1593 21848
rect 1627 21845 1639 21879
rect 1581 21839 1639 21845
rect 3145 21879 3203 21885
rect 3145 21845 3157 21879
rect 3191 21876 3203 21879
rect 5442 21876 5448 21888
rect 3191 21848 5448 21876
rect 3191 21845 3203 21848
rect 3145 21839 3203 21845
rect 5442 21836 5448 21848
rect 5500 21836 5506 21888
rect 6365 21879 6423 21885
rect 6365 21845 6377 21879
rect 6411 21876 6423 21879
rect 6454 21876 6460 21888
rect 6411 21848 6460 21876
rect 6411 21845 6423 21848
rect 6365 21839 6423 21845
rect 6454 21836 6460 21848
rect 6512 21836 6518 21888
rect 7944 21876 7972 21916
rect 9769 21913 9781 21947
rect 9815 21913 9827 21947
rect 9876 21944 9904 22052
rect 10410 22040 10416 22092
rect 10468 22040 10474 22092
rect 10597 22083 10655 22089
rect 10597 22049 10609 22083
rect 10643 22080 10655 22083
rect 10965 22083 11023 22089
rect 10965 22080 10977 22083
rect 10643 22052 10977 22080
rect 10643 22049 10655 22052
rect 10597 22043 10655 22049
rect 10965 22049 10977 22052
rect 11011 22049 11023 22083
rect 10965 22043 11023 22049
rect 11330 22040 11336 22092
rect 11388 22080 11394 22092
rect 11790 22080 11796 22092
rect 11388 22052 11796 22080
rect 11388 22040 11394 22052
rect 11790 22040 11796 22052
rect 11848 22040 11854 22092
rect 12250 22040 12256 22092
rect 12308 22080 12314 22092
rect 12437 22083 12495 22089
rect 12437 22080 12449 22083
rect 12308 22052 12449 22080
rect 12308 22040 12314 22052
rect 12437 22049 12449 22052
rect 12483 22049 12495 22083
rect 12437 22043 12495 22049
rect 12621 22083 12679 22089
rect 12621 22049 12633 22083
rect 12667 22049 12679 22083
rect 12621 22043 12679 22049
rect 10134 21972 10140 22024
rect 10192 22012 10198 22024
rect 10229 22015 10287 22021
rect 10229 22012 10241 22015
rect 10192 21984 10241 22012
rect 10192 21972 10198 21984
rect 10229 21981 10241 21984
rect 10275 21981 10287 22015
rect 10229 21975 10287 21981
rect 12342 21972 12348 22024
rect 12400 22012 12406 22024
rect 12636 22012 12664 22043
rect 13372 22024 13400 22120
rect 13909 22117 13921 22151
rect 13955 22148 13967 22151
rect 14182 22148 14188 22160
rect 13955 22120 14188 22148
rect 13955 22117 13967 22120
rect 13909 22111 13967 22117
rect 14182 22108 14188 22120
rect 14240 22108 14246 22160
rect 15286 22148 15292 22160
rect 15212 22120 15292 22148
rect 13817 22083 13875 22089
rect 13817 22049 13829 22083
rect 13863 22080 13875 22083
rect 15013 22083 15071 22089
rect 15013 22080 15025 22083
rect 13863 22052 15025 22080
rect 13863 22049 13875 22052
rect 13817 22043 13875 22049
rect 15013 22049 15025 22052
rect 15059 22080 15071 22083
rect 15212 22080 15240 22120
rect 15286 22108 15292 22120
rect 15344 22148 15350 22160
rect 15749 22151 15807 22157
rect 15749 22148 15761 22151
rect 15344 22120 15761 22148
rect 15344 22108 15350 22120
rect 15749 22117 15761 22120
rect 15795 22117 15807 22151
rect 16316 22148 16344 22179
rect 16666 22176 16672 22228
rect 16724 22216 16730 22228
rect 19518 22216 19524 22228
rect 16724 22188 19524 22216
rect 16724 22176 16730 22188
rect 19518 22176 19524 22188
rect 19576 22176 19582 22228
rect 22097 22219 22155 22225
rect 22097 22185 22109 22219
rect 22143 22216 22155 22219
rect 22554 22216 22560 22228
rect 22143 22188 22560 22216
rect 22143 22185 22155 22188
rect 22097 22179 22155 22185
rect 22554 22176 22560 22188
rect 22612 22176 22618 22228
rect 22848 22188 23152 22216
rect 17034 22148 17040 22160
rect 16316 22120 17040 22148
rect 15749 22111 15807 22117
rect 17034 22108 17040 22120
rect 17092 22148 17098 22160
rect 17770 22148 17776 22160
rect 17092 22120 17776 22148
rect 17092 22108 17098 22120
rect 17770 22108 17776 22120
rect 17828 22108 17834 22160
rect 21726 22108 21732 22160
rect 21784 22148 21790 22160
rect 21821 22151 21879 22157
rect 21821 22148 21833 22151
rect 21784 22120 21833 22148
rect 21784 22108 21790 22120
rect 21821 22117 21833 22120
rect 21867 22148 21879 22151
rect 22005 22151 22063 22157
rect 21867 22120 21956 22148
rect 21867 22117 21879 22120
rect 21821 22111 21879 22117
rect 15059 22052 15240 22080
rect 15565 22083 15623 22089
rect 15059 22049 15071 22052
rect 15013 22043 15071 22049
rect 15565 22049 15577 22083
rect 15611 22049 15623 22083
rect 15565 22043 15623 22049
rect 15933 22083 15991 22089
rect 15933 22049 15945 22083
rect 15979 22080 15991 22083
rect 16117 22083 16175 22089
rect 16117 22080 16129 22083
rect 15979 22052 16129 22080
rect 15979 22049 15991 22052
rect 15933 22043 15991 22049
rect 16117 22049 16129 22052
rect 16163 22049 16175 22083
rect 16117 22043 16175 22049
rect 12400 21984 12664 22012
rect 12400 21972 12406 21984
rect 13354 21972 13360 22024
rect 13412 22012 13418 22024
rect 14737 22015 14795 22021
rect 14737 22012 14749 22015
rect 13412 21984 14749 22012
rect 13412 21972 13418 21984
rect 14737 21981 14749 21984
rect 14783 22012 14795 22015
rect 15194 22012 15200 22024
rect 14783 21984 15200 22012
rect 14783 21981 14795 21984
rect 14737 21975 14795 21981
rect 15194 21972 15200 21984
rect 15252 21972 15258 22024
rect 15289 22015 15347 22021
rect 15289 21981 15301 22015
rect 15335 22012 15347 22015
rect 15580 22012 15608 22043
rect 16758 22040 16764 22092
rect 16816 22080 16822 22092
rect 17129 22083 17187 22089
rect 17129 22080 17141 22083
rect 16816 22052 17141 22080
rect 16816 22040 16822 22052
rect 17129 22049 17141 22052
rect 17175 22080 17187 22083
rect 17865 22083 17923 22089
rect 17865 22080 17877 22083
rect 17175 22052 17877 22080
rect 17175 22049 17187 22052
rect 17129 22043 17187 22049
rect 17865 22049 17877 22052
rect 17911 22049 17923 22083
rect 17865 22043 17923 22049
rect 18785 22083 18843 22089
rect 18785 22049 18797 22083
rect 18831 22080 18843 22083
rect 18874 22080 18880 22092
rect 18831 22052 18880 22080
rect 18831 22049 18843 22052
rect 18785 22043 18843 22049
rect 18874 22040 18880 22052
rect 18932 22040 18938 22092
rect 19052 22083 19110 22089
rect 19052 22049 19064 22083
rect 19098 22080 19110 22083
rect 20162 22080 20168 22092
rect 19098 22052 20168 22080
rect 19098 22049 19110 22052
rect 19052 22043 19110 22049
rect 20162 22040 20168 22052
rect 20220 22040 20226 22092
rect 20349 22015 20407 22021
rect 20349 22012 20361 22015
rect 15335 21984 15608 22012
rect 20180 21984 20361 22012
rect 15335 21981 15347 21984
rect 15289 21975 15347 21981
rect 13446 21944 13452 21956
rect 9876 21916 13452 21944
rect 9769 21907 9827 21913
rect 13446 21904 13452 21916
rect 13504 21904 13510 21956
rect 15304 21944 15332 21975
rect 13740 21916 15332 21944
rect 13740 21888 13768 21916
rect 15746 21904 15752 21956
rect 15804 21944 15810 21956
rect 16114 21944 16120 21956
rect 15804 21916 16120 21944
rect 15804 21904 15810 21916
rect 16114 21904 16120 21916
rect 16172 21944 16178 21956
rect 17313 21947 17371 21953
rect 17313 21944 17325 21947
rect 16172 21916 17325 21944
rect 16172 21904 16178 21916
rect 17313 21913 17325 21916
rect 17359 21913 17371 21947
rect 17313 21907 17371 21913
rect 17770 21904 17776 21956
rect 17828 21904 17834 21956
rect 20180 21953 20208 21984
rect 20349 21981 20361 21984
rect 20395 22012 20407 22015
rect 21450 22012 21456 22024
rect 20395 21984 21456 22012
rect 20395 21981 20407 21984
rect 20349 21975 20407 21981
rect 21450 21972 21456 21984
rect 21508 21972 21514 22024
rect 21928 22012 21956 22120
rect 22005 22117 22017 22151
rect 22051 22148 22063 22151
rect 22465 22151 22523 22157
rect 22465 22148 22477 22151
rect 22051 22120 22477 22148
rect 22051 22117 22063 22120
rect 22005 22111 22063 22117
rect 22465 22117 22477 22120
rect 22511 22148 22523 22151
rect 22646 22148 22652 22160
rect 22511 22120 22652 22148
rect 22511 22117 22523 22120
rect 22465 22111 22523 22117
rect 22646 22108 22652 22120
rect 22704 22108 22710 22160
rect 22738 22108 22744 22160
rect 22796 22108 22802 22160
rect 22848 22157 22876 22188
rect 22833 22151 22891 22157
rect 22833 22117 22845 22151
rect 22879 22117 22891 22151
rect 22833 22111 22891 22117
rect 23014 22108 23020 22160
rect 23072 22157 23078 22160
rect 23072 22151 23091 22157
rect 23079 22117 23091 22151
rect 23124 22148 23152 22188
rect 23198 22176 23204 22228
rect 23256 22176 23262 22228
rect 23290 22148 23296 22160
rect 23124 22120 23296 22148
rect 23072 22111 23091 22117
rect 23072 22108 23078 22111
rect 23290 22108 23296 22120
rect 23348 22108 23354 22160
rect 22097 22083 22155 22089
rect 22097 22049 22109 22083
rect 22143 22080 22155 22083
rect 22278 22080 22284 22092
rect 22143 22052 22284 22080
rect 22143 22049 22155 22052
rect 22097 22043 22155 22049
rect 22278 22040 22284 22052
rect 22336 22080 22342 22092
rect 22373 22083 22431 22089
rect 22373 22080 22385 22083
rect 22336 22052 22385 22080
rect 22336 22040 22342 22052
rect 22373 22049 22385 22052
rect 22419 22049 22431 22083
rect 22373 22043 22431 22049
rect 22557 22083 22615 22089
rect 22557 22049 22569 22083
rect 22603 22080 22615 22083
rect 22756 22080 22784 22108
rect 22603 22052 22784 22080
rect 22603 22049 22615 22052
rect 22557 22043 22615 22049
rect 22388 22012 22416 22043
rect 23934 22040 23940 22092
rect 23992 22080 23998 22092
rect 24406 22083 24464 22089
rect 24406 22080 24418 22083
rect 23992 22052 24418 22080
rect 23992 22040 23998 22052
rect 24406 22049 24418 22052
rect 24452 22049 24464 22083
rect 24406 22043 24464 22049
rect 22922 22012 22928 22024
rect 21928 21984 22140 22012
rect 22388 21984 22928 22012
rect 22112 21956 22140 21984
rect 22922 21972 22928 21984
rect 22980 22012 22986 22024
rect 24673 22015 24731 22021
rect 22980 21984 23336 22012
rect 22980 21972 22986 21984
rect 20165 21947 20223 21953
rect 20165 21913 20177 21947
rect 20211 21913 20223 21947
rect 20165 21907 20223 21913
rect 22094 21904 22100 21956
rect 22152 21904 22158 21956
rect 22186 21904 22192 21956
rect 22244 21904 22250 21956
rect 22554 21904 22560 21956
rect 22612 21944 22618 21956
rect 23308 21953 23336 21984
rect 24673 21981 24685 22015
rect 24719 22012 24731 22015
rect 25590 22012 25596 22024
rect 24719 21984 25596 22012
rect 24719 21981 24731 21984
rect 24673 21975 24731 21981
rect 25590 21972 25596 21984
rect 25648 21972 25654 22024
rect 23293 21947 23351 21953
rect 22612 21916 23060 21944
rect 22612 21904 22618 21916
rect 9398 21876 9404 21888
rect 7944 21848 9404 21876
rect 9398 21836 9404 21848
rect 9456 21836 9462 21888
rect 9950 21836 9956 21888
rect 10008 21876 10014 21888
rect 10318 21876 10324 21888
rect 10008 21848 10324 21876
rect 10008 21836 10014 21848
rect 10318 21836 10324 21848
rect 10376 21836 10382 21888
rect 11149 21879 11207 21885
rect 11149 21845 11161 21879
rect 11195 21876 11207 21879
rect 11238 21876 11244 21888
rect 11195 21848 11244 21876
rect 11195 21845 11207 21848
rect 11149 21839 11207 21845
rect 11238 21836 11244 21848
rect 11296 21836 11302 21888
rect 12161 21879 12219 21885
rect 12161 21845 12173 21879
rect 12207 21876 12219 21879
rect 12250 21876 12256 21888
rect 12207 21848 12256 21876
rect 12207 21845 12219 21848
rect 12161 21839 12219 21845
rect 12250 21836 12256 21848
rect 12308 21876 12314 21888
rect 13262 21876 13268 21888
rect 12308 21848 13268 21876
rect 12308 21836 12314 21848
rect 13262 21836 13268 21848
rect 13320 21836 13326 21888
rect 13722 21836 13728 21888
rect 13780 21836 13786 21888
rect 15381 21879 15439 21885
rect 15381 21845 15393 21879
rect 15427 21876 15439 21879
rect 16482 21876 16488 21888
rect 15427 21848 16488 21876
rect 15427 21845 15439 21848
rect 15381 21839 15439 21845
rect 16482 21836 16488 21848
rect 16540 21876 16546 21888
rect 17218 21876 17224 21888
rect 16540 21848 17224 21876
rect 16540 21836 16546 21848
rect 17218 21836 17224 21848
rect 17276 21836 17282 21888
rect 20806 21836 20812 21888
rect 20864 21876 20870 21888
rect 20901 21879 20959 21885
rect 20901 21876 20913 21879
rect 20864 21848 20913 21876
rect 20864 21836 20870 21848
rect 20901 21845 20913 21848
rect 20947 21845 20959 21879
rect 20901 21839 20959 21845
rect 22738 21836 22744 21888
rect 22796 21836 22802 21888
rect 23032 21885 23060 21916
rect 23293 21913 23305 21947
rect 23339 21913 23351 21947
rect 23293 21907 23351 21913
rect 23017 21879 23075 21885
rect 23017 21845 23029 21879
rect 23063 21845 23075 21879
rect 23017 21839 23075 21845
rect 552 21786 27416 21808
rect 552 21734 3756 21786
rect 3808 21734 3820 21786
rect 3872 21734 3884 21786
rect 3936 21734 3948 21786
rect 4000 21734 4012 21786
rect 4064 21734 10472 21786
rect 10524 21734 10536 21786
rect 10588 21734 10600 21786
rect 10652 21734 10664 21786
rect 10716 21734 10728 21786
rect 10780 21734 17188 21786
rect 17240 21734 17252 21786
rect 17304 21734 17316 21786
rect 17368 21734 17380 21786
rect 17432 21734 17444 21786
rect 17496 21734 23904 21786
rect 23956 21734 23968 21786
rect 24020 21734 24032 21786
rect 24084 21734 24096 21786
rect 24148 21734 24160 21786
rect 24212 21734 27416 21786
rect 552 21712 27416 21734
rect 1578 21632 1584 21684
rect 1636 21672 1642 21684
rect 1946 21672 1952 21684
rect 1636 21644 1952 21672
rect 1636 21632 1642 21644
rect 1946 21632 1952 21644
rect 2004 21672 2010 21684
rect 2685 21675 2743 21681
rect 2685 21672 2697 21675
rect 2004 21644 2697 21672
rect 2004 21632 2010 21644
rect 2685 21641 2697 21644
rect 2731 21641 2743 21675
rect 2685 21635 2743 21641
rect 4246 21632 4252 21684
rect 4304 21672 4310 21684
rect 4893 21675 4951 21681
rect 4893 21672 4905 21675
rect 4304 21644 4905 21672
rect 4304 21632 4310 21644
rect 4893 21641 4905 21644
rect 4939 21641 4951 21675
rect 4893 21635 4951 21641
rect 5902 21632 5908 21684
rect 5960 21632 5966 21684
rect 7193 21675 7251 21681
rect 7193 21641 7205 21675
rect 7239 21672 7251 21675
rect 7558 21672 7564 21684
rect 7239 21644 7564 21672
rect 7239 21641 7251 21644
rect 7193 21635 7251 21641
rect 7558 21632 7564 21644
rect 7616 21632 7622 21684
rect 8573 21675 8631 21681
rect 8573 21641 8585 21675
rect 8619 21672 8631 21675
rect 8662 21672 8668 21684
rect 8619 21644 8668 21672
rect 8619 21641 8631 21644
rect 8573 21635 8631 21641
rect 8662 21632 8668 21644
rect 8720 21672 8726 21684
rect 9030 21672 9036 21684
rect 8720 21644 9036 21672
rect 8720 21632 8726 21644
rect 9030 21632 9036 21644
rect 9088 21632 9094 21684
rect 10137 21675 10195 21681
rect 10137 21641 10149 21675
rect 10183 21672 10195 21675
rect 11330 21672 11336 21684
rect 10183 21644 11336 21672
rect 10183 21641 10195 21644
rect 10137 21635 10195 21641
rect 11330 21632 11336 21644
rect 11388 21632 11394 21684
rect 13722 21632 13728 21684
rect 13780 21672 13786 21684
rect 13780 21644 14688 21672
rect 13780 21632 13786 21644
rect 2038 21564 2044 21616
rect 2096 21604 2102 21616
rect 2317 21607 2375 21613
rect 2317 21604 2329 21607
rect 2096 21576 2329 21604
rect 2096 21564 2102 21576
rect 2317 21573 2329 21576
rect 2363 21573 2375 21607
rect 5534 21604 5540 21616
rect 2317 21567 2375 21573
rect 5460 21576 5540 21604
rect 3237 21539 3295 21545
rect 3237 21536 3249 21539
rect 1872 21508 3249 21536
rect 842 21428 848 21480
rect 900 21468 906 21480
rect 1872 21468 1900 21508
rect 3237 21505 3249 21508
rect 3283 21505 3295 21539
rect 3237 21499 3295 21505
rect 900 21440 1900 21468
rect 900 21428 906 21440
rect 934 21360 940 21412
rect 992 21400 998 21412
rect 1090 21403 1148 21409
rect 1090 21400 1102 21403
rect 992 21372 1102 21400
rect 992 21360 998 21372
rect 1090 21369 1102 21372
rect 1136 21369 1148 21403
rect 1090 21363 1148 21369
rect 2958 21360 2964 21412
rect 3016 21400 3022 21412
rect 3482 21403 3540 21409
rect 3482 21400 3494 21403
rect 3016 21372 3494 21400
rect 3016 21360 3022 21372
rect 3482 21369 3494 21372
rect 3528 21369 3540 21403
rect 3482 21363 3540 21369
rect 4154 21360 4160 21412
rect 4212 21400 4218 21412
rect 5077 21403 5135 21409
rect 5077 21400 5089 21403
rect 4212 21372 5089 21400
rect 4212 21360 4218 21372
rect 5077 21369 5089 21372
rect 5123 21369 5135 21403
rect 5460 21400 5488 21576
rect 5534 21564 5540 21576
rect 5592 21564 5598 21616
rect 6730 21564 6736 21616
rect 6788 21604 6794 21616
rect 8938 21604 8944 21616
rect 6788 21576 8944 21604
rect 6788 21564 6794 21576
rect 8938 21564 8944 21576
rect 8996 21564 9002 21616
rect 11514 21564 11520 21616
rect 11572 21604 11578 21616
rect 14550 21604 14556 21616
rect 11572 21576 13860 21604
rect 11572 21564 11578 21576
rect 7006 21536 7012 21548
rect 5552 21508 7012 21536
rect 5552 21477 5580 21508
rect 7006 21496 7012 21508
rect 7064 21496 7070 21548
rect 7834 21536 7840 21548
rect 7208 21508 7840 21536
rect 5537 21471 5595 21477
rect 5537 21437 5549 21471
rect 5583 21437 5595 21471
rect 5537 21431 5595 21437
rect 5813 21471 5871 21477
rect 5813 21437 5825 21471
rect 5859 21437 5871 21471
rect 5813 21431 5871 21437
rect 5721 21403 5779 21409
rect 5721 21400 5733 21403
rect 5460 21372 5733 21400
rect 5077 21363 5135 21369
rect 5721 21369 5733 21372
rect 5767 21369 5779 21403
rect 5721 21363 5779 21369
rect 2225 21335 2283 21341
rect 2225 21301 2237 21335
rect 2271 21332 2283 21335
rect 2590 21332 2596 21344
rect 2271 21304 2596 21332
rect 2271 21301 2283 21304
rect 2225 21295 2283 21301
rect 2590 21292 2596 21304
rect 2648 21292 2654 21344
rect 2682 21292 2688 21344
rect 2740 21292 2746 21344
rect 2866 21292 2872 21344
rect 2924 21292 2930 21344
rect 3326 21292 3332 21344
rect 3384 21332 3390 21344
rect 4617 21335 4675 21341
rect 4617 21332 4629 21335
rect 3384 21304 4629 21332
rect 3384 21292 3390 21304
rect 4617 21301 4629 21304
rect 4663 21301 4675 21335
rect 4617 21295 4675 21301
rect 4706 21292 4712 21344
rect 4764 21292 4770 21344
rect 4890 21341 4896 21344
rect 4877 21335 4896 21341
rect 4877 21301 4889 21335
rect 4877 21295 4896 21301
rect 4890 21292 4896 21295
rect 4948 21292 4954 21344
rect 5353 21335 5411 21341
rect 5353 21301 5365 21335
rect 5399 21332 5411 21335
rect 5534 21332 5540 21344
rect 5399 21304 5540 21332
rect 5399 21301 5411 21304
rect 5353 21295 5411 21301
rect 5534 21292 5540 21304
rect 5592 21292 5598 21344
rect 5828 21332 5856 21431
rect 6086 21428 6092 21480
rect 6144 21428 6150 21480
rect 6270 21428 6276 21480
rect 6328 21428 6334 21480
rect 6454 21428 6460 21480
rect 6512 21428 6518 21480
rect 6641 21471 6699 21477
rect 6641 21437 6653 21471
rect 6687 21468 6699 21471
rect 6730 21468 6736 21480
rect 6687 21440 6736 21468
rect 6687 21437 6699 21440
rect 6641 21431 6699 21437
rect 6730 21428 6736 21440
rect 6788 21428 6794 21480
rect 7208 21468 7236 21508
rect 7834 21496 7840 21508
rect 7892 21536 7898 21548
rect 7892 21508 9674 21536
rect 7892 21496 7898 21508
rect 6932 21440 7236 21468
rect 7285 21471 7343 21477
rect 6181 21403 6239 21409
rect 6181 21369 6193 21403
rect 6227 21400 6239 21403
rect 6932 21400 6960 21440
rect 7285 21437 7297 21471
rect 7331 21437 7343 21471
rect 9646 21468 9674 21508
rect 11790 21496 11796 21548
rect 11848 21536 11854 21548
rect 12066 21536 12072 21548
rect 11848 21508 12072 21536
rect 11848 21496 11854 21508
rect 12066 21496 12072 21508
rect 12124 21536 12130 21548
rect 13081 21539 13139 21545
rect 12124 21508 12434 21536
rect 12124 21496 12130 21508
rect 9646 21440 11192 21468
rect 7285 21431 7343 21437
rect 6227 21372 6960 21400
rect 6227 21369 6239 21372
rect 6181 21363 6239 21369
rect 7006 21360 7012 21412
rect 7064 21400 7070 21412
rect 7300 21400 7328 21431
rect 7064 21372 7328 21400
rect 7929 21403 7987 21409
rect 7064 21360 7070 21372
rect 7929 21369 7941 21403
rect 7975 21400 7987 21403
rect 8757 21403 8815 21409
rect 8757 21400 8769 21403
rect 7975 21372 8769 21400
rect 7975 21369 7987 21372
rect 7929 21363 7987 21369
rect 8757 21369 8769 21372
rect 8803 21369 8815 21403
rect 8757 21363 8815 21369
rect 8938 21360 8944 21412
rect 8996 21400 9002 21412
rect 11054 21400 11060 21412
rect 8996 21372 11060 21400
rect 8996 21360 9002 21372
rect 11054 21360 11060 21372
rect 11112 21360 11118 21412
rect 7466 21332 7472 21344
rect 5828 21304 7472 21332
rect 7466 21292 7472 21304
rect 7524 21292 7530 21344
rect 8386 21292 8392 21344
rect 8444 21292 8450 21344
rect 8570 21341 8576 21344
rect 8557 21335 8576 21341
rect 8557 21301 8569 21335
rect 8557 21295 8576 21301
rect 8570 21292 8576 21295
rect 8628 21292 8634 21344
rect 11164 21332 11192 21440
rect 11238 21428 11244 21480
rect 11296 21477 11302 21480
rect 11296 21468 11308 21477
rect 11296 21440 11341 21468
rect 11296 21431 11308 21440
rect 11296 21428 11302 21431
rect 11422 21428 11428 21480
rect 11480 21468 11486 21480
rect 11517 21471 11575 21477
rect 11517 21468 11529 21471
rect 11480 21440 11529 21468
rect 11480 21428 11486 21440
rect 11517 21437 11529 21440
rect 11563 21437 11575 21471
rect 11517 21431 11575 21437
rect 12158 21428 12164 21480
rect 12216 21428 12222 21480
rect 12406 21468 12434 21508
rect 13081 21505 13093 21539
rect 13127 21536 13139 21539
rect 13722 21536 13728 21548
rect 13127 21508 13728 21536
rect 13127 21505 13139 21508
rect 13081 21499 13139 21505
rect 13722 21496 13728 21508
rect 13780 21496 13786 21548
rect 12529 21471 12587 21477
rect 12529 21468 12541 21471
rect 12406 21440 12541 21468
rect 12529 21437 12541 21440
rect 12575 21437 12587 21471
rect 12529 21431 12587 21437
rect 13265 21471 13323 21477
rect 13265 21437 13277 21471
rect 13311 21437 13323 21471
rect 13265 21431 13323 21437
rect 11882 21360 11888 21412
rect 11940 21400 11946 21412
rect 12342 21400 12348 21412
rect 11940 21372 12348 21400
rect 11940 21360 11946 21372
rect 12342 21360 12348 21372
rect 12400 21400 12406 21412
rect 13280 21400 13308 21431
rect 12400 21372 13308 21400
rect 12400 21360 12406 21372
rect 12526 21332 12532 21344
rect 11164 21304 12532 21332
rect 12526 21292 12532 21304
rect 12584 21292 12590 21344
rect 13078 21292 13084 21344
rect 13136 21332 13142 21344
rect 13541 21335 13599 21341
rect 13541 21332 13553 21335
rect 13136 21304 13553 21332
rect 13136 21292 13142 21304
rect 13541 21301 13553 21304
rect 13587 21301 13599 21335
rect 13832 21332 13860 21576
rect 13924 21576 14556 21604
rect 13924 21477 13952 21576
rect 14550 21564 14556 21576
rect 14608 21564 14614 21616
rect 14185 21539 14243 21545
rect 14185 21505 14197 21539
rect 14231 21536 14243 21539
rect 14366 21536 14372 21548
rect 14231 21508 14372 21536
rect 14231 21505 14243 21508
rect 14185 21499 14243 21505
rect 14366 21496 14372 21508
rect 14424 21496 14430 21548
rect 13909 21471 13967 21477
rect 13909 21437 13921 21471
rect 13955 21437 13967 21471
rect 13909 21431 13967 21437
rect 14001 21471 14059 21477
rect 14001 21437 14013 21471
rect 14047 21468 14059 21471
rect 14553 21471 14611 21477
rect 14553 21468 14565 21471
rect 14047 21440 14565 21468
rect 14047 21437 14059 21440
rect 14001 21431 14059 21437
rect 14553 21437 14565 21440
rect 14599 21437 14611 21471
rect 14660 21468 14688 21644
rect 20162 21632 20168 21684
rect 20220 21672 20226 21684
rect 20257 21675 20315 21681
rect 20257 21672 20269 21675
rect 20220 21644 20269 21672
rect 20220 21632 20226 21644
rect 20257 21641 20269 21644
rect 20303 21641 20315 21675
rect 22281 21675 22339 21681
rect 22281 21672 22293 21675
rect 20257 21635 20315 21641
rect 22066 21644 22293 21672
rect 14734 21564 14740 21616
rect 14792 21604 14798 21616
rect 16850 21604 16856 21616
rect 14792 21576 16856 21604
rect 14792 21564 14798 21576
rect 16850 21564 16856 21576
rect 16908 21564 16914 21616
rect 18509 21607 18567 21613
rect 18509 21573 18521 21607
rect 18555 21604 18567 21607
rect 18555 21576 19288 21604
rect 18555 21573 18567 21576
rect 18509 21567 18567 21573
rect 15194 21496 15200 21548
rect 15252 21536 15258 21548
rect 19260 21545 19288 21576
rect 21910 21564 21916 21616
rect 21968 21604 21974 21616
rect 22066 21604 22094 21644
rect 22281 21641 22293 21644
rect 22327 21672 22339 21675
rect 22370 21672 22376 21684
rect 22327 21644 22376 21672
rect 22327 21641 22339 21644
rect 22281 21635 22339 21641
rect 22370 21632 22376 21644
rect 22428 21632 22434 21684
rect 22462 21632 22468 21684
rect 22520 21672 22526 21684
rect 23109 21675 23167 21681
rect 23109 21672 23121 21675
rect 22520 21644 23121 21672
rect 22520 21632 22526 21644
rect 23109 21641 23121 21644
rect 23155 21641 23167 21675
rect 23109 21635 23167 21641
rect 23293 21675 23351 21681
rect 23293 21641 23305 21675
rect 23339 21672 23351 21675
rect 23474 21672 23480 21684
rect 23339 21644 23480 21672
rect 23339 21641 23351 21644
rect 23293 21635 23351 21641
rect 23474 21632 23480 21644
rect 23532 21632 23538 21684
rect 25590 21672 25596 21684
rect 25332 21644 25596 21672
rect 21968 21576 22094 21604
rect 21968 21564 21974 21576
rect 22186 21564 22192 21616
rect 22244 21604 22250 21616
rect 22244 21576 22324 21604
rect 22244 21564 22250 21576
rect 17129 21539 17187 21545
rect 17129 21536 17141 21539
rect 15252 21508 17141 21536
rect 15252 21496 15258 21508
rect 17129 21505 17141 21508
rect 17175 21505 17187 21539
rect 17129 21499 17187 21505
rect 19245 21539 19303 21545
rect 19245 21505 19257 21539
rect 19291 21536 19303 21539
rect 20346 21536 20352 21548
rect 19291 21508 20352 21536
rect 19291 21505 19303 21508
rect 19245 21499 19303 21505
rect 20346 21496 20352 21508
rect 20404 21496 20410 21548
rect 22296 21536 22324 21576
rect 22738 21564 22744 21616
rect 22796 21564 22802 21616
rect 23845 21607 23903 21613
rect 23845 21573 23857 21607
rect 23891 21573 23903 21607
rect 23845 21567 23903 21573
rect 23860 21536 23888 21567
rect 25332 21545 25360 21644
rect 25590 21632 25596 21644
rect 25648 21632 25654 21684
rect 22112 21508 23888 21536
rect 25225 21539 25283 21545
rect 14737 21471 14795 21477
rect 14737 21468 14749 21471
rect 14660 21440 14749 21468
rect 14553 21431 14611 21437
rect 14737 21437 14749 21440
rect 14783 21437 14795 21471
rect 15286 21468 15292 21480
rect 14737 21431 14795 21437
rect 14844 21440 15292 21468
rect 14568 21400 14596 21431
rect 14844 21400 14872 21440
rect 15286 21428 15292 21440
rect 15344 21428 15350 21480
rect 16114 21428 16120 21480
rect 16172 21428 16178 21480
rect 16206 21428 16212 21480
rect 16264 21468 16270 21480
rect 16264 21440 16896 21468
rect 16264 21428 16270 21440
rect 14568 21372 14872 21400
rect 15102 21360 15108 21412
rect 15160 21400 15166 21412
rect 16577 21403 16635 21409
rect 16577 21400 16589 21403
rect 15160 21372 16589 21400
rect 15160 21360 15166 21372
rect 16577 21369 16589 21372
rect 16623 21369 16635 21403
rect 16577 21363 16635 21369
rect 15654 21332 15660 21344
rect 13832 21304 15660 21332
rect 13541 21295 13599 21301
rect 15654 21292 15660 21304
rect 15712 21292 15718 21344
rect 15930 21292 15936 21344
rect 15988 21332 15994 21344
rect 16301 21335 16359 21341
rect 16301 21332 16313 21335
rect 15988 21304 16313 21332
rect 15988 21292 15994 21304
rect 16301 21301 16313 21304
rect 16347 21332 16359 21335
rect 16390 21332 16396 21344
rect 16347 21304 16396 21332
rect 16347 21301 16359 21304
rect 16301 21295 16359 21301
rect 16390 21292 16396 21304
rect 16448 21292 16454 21344
rect 16868 21341 16896 21440
rect 20162 21428 20168 21480
rect 20220 21428 20226 21480
rect 20438 21428 20444 21480
rect 20496 21428 20502 21480
rect 20806 21428 20812 21480
rect 20864 21428 20870 21480
rect 21082 21428 21088 21480
rect 21140 21428 21146 21480
rect 21266 21477 21272 21480
rect 21233 21471 21272 21477
rect 21233 21437 21245 21471
rect 21233 21431 21272 21437
rect 21266 21428 21272 21431
rect 21324 21428 21330 21480
rect 21591 21471 21649 21477
rect 21591 21437 21603 21471
rect 21637 21468 21649 21471
rect 22002 21468 22008 21480
rect 21637 21440 22008 21468
rect 21637 21437 21649 21440
rect 21591 21431 21649 21437
rect 22002 21428 22008 21440
rect 22060 21428 22066 21480
rect 22112 21468 22140 21508
rect 25225 21505 25237 21539
rect 25271 21536 25283 21539
rect 25317 21539 25375 21545
rect 25317 21536 25329 21539
rect 25271 21508 25329 21536
rect 25271 21505 25283 21508
rect 25225 21499 25283 21505
rect 25317 21505 25329 21508
rect 25363 21505 25375 21539
rect 25317 21499 25375 21505
rect 22181 21471 22239 21477
rect 22181 21468 22193 21471
rect 22112 21440 22193 21468
rect 22181 21437 22193 21440
rect 22227 21437 22239 21471
rect 22181 21431 22239 21437
rect 17402 21409 17408 21412
rect 17396 21363 17408 21409
rect 17402 21360 17408 21363
rect 17460 21360 17466 21412
rect 17954 21360 17960 21412
rect 18012 21400 18018 21412
rect 18693 21403 18751 21409
rect 18693 21400 18705 21403
rect 18012 21372 18705 21400
rect 18012 21360 18018 21372
rect 18693 21369 18705 21372
rect 18739 21369 18751 21403
rect 20533 21403 20591 21409
rect 20533 21400 20545 21403
rect 18693 21363 18751 21369
rect 18800 21372 20545 21400
rect 16853 21335 16911 21341
rect 16853 21301 16865 21335
rect 16899 21332 16911 21335
rect 18414 21332 18420 21344
rect 16899 21304 18420 21332
rect 16899 21301 16911 21304
rect 16853 21295 16911 21301
rect 18414 21292 18420 21304
rect 18472 21332 18478 21344
rect 18800 21332 18828 21372
rect 20533 21369 20545 21372
rect 20579 21369 20591 21403
rect 20533 21363 20591 21369
rect 20625 21403 20683 21409
rect 20625 21369 20637 21403
rect 20671 21369 20683 21403
rect 20625 21363 20683 21369
rect 18472 21304 18828 21332
rect 18472 21292 18478 21304
rect 18874 21292 18880 21344
rect 18932 21332 18938 21344
rect 19521 21335 19579 21341
rect 19521 21332 19533 21335
rect 18932 21304 19533 21332
rect 18932 21292 18938 21304
rect 19521 21301 19533 21304
rect 19567 21301 19579 21335
rect 19521 21295 19579 21301
rect 19794 21292 19800 21344
rect 19852 21332 19858 21344
rect 20640 21332 20668 21363
rect 20990 21360 20996 21412
rect 21048 21400 21054 21412
rect 21361 21403 21419 21409
rect 21361 21400 21373 21403
rect 21048 21372 21373 21400
rect 21048 21360 21054 21372
rect 21361 21369 21373 21372
rect 21407 21369 21419 21403
rect 21361 21363 21419 21369
rect 21453 21403 21511 21409
rect 21453 21369 21465 21403
rect 21499 21400 21511 21403
rect 21910 21400 21916 21412
rect 21499 21372 21916 21400
rect 21499 21369 21511 21372
rect 21453 21363 21511 21369
rect 21910 21360 21916 21372
rect 21968 21360 21974 21412
rect 22646 21360 22652 21412
rect 22704 21400 22710 21412
rect 22704 21372 24716 21400
rect 22704 21360 22710 21372
rect 19852 21304 20668 21332
rect 21729 21335 21787 21341
rect 19852 21292 19858 21304
rect 21729 21301 21741 21335
rect 21775 21332 21787 21335
rect 22370 21332 22376 21344
rect 21775 21304 22376 21332
rect 21775 21301 21787 21304
rect 21729 21295 21787 21301
rect 22370 21292 22376 21304
rect 22428 21292 22434 21344
rect 23109 21335 23167 21341
rect 23109 21301 23121 21335
rect 23155 21332 23167 21335
rect 23290 21332 23296 21344
rect 23155 21304 23296 21332
rect 23155 21301 23167 21304
rect 23109 21295 23167 21301
rect 23290 21292 23296 21304
rect 23348 21292 23354 21344
rect 24688 21332 24716 21372
rect 24854 21360 24860 21412
rect 24912 21400 24918 21412
rect 25590 21409 25596 21412
rect 24958 21403 25016 21409
rect 24958 21400 24970 21403
rect 24912 21372 24970 21400
rect 24912 21360 24918 21372
rect 24958 21369 24970 21372
rect 25004 21369 25016 21403
rect 24958 21363 25016 21369
rect 25584 21363 25596 21409
rect 25590 21360 25596 21363
rect 25648 21360 25654 21412
rect 26697 21335 26755 21341
rect 26697 21332 26709 21335
rect 24688 21304 26709 21332
rect 26697 21301 26709 21304
rect 26743 21332 26755 21335
rect 26970 21332 26976 21344
rect 26743 21304 26976 21332
rect 26743 21301 26755 21304
rect 26697 21295 26755 21301
rect 26970 21292 26976 21304
rect 27028 21292 27034 21344
rect 552 21242 27576 21264
rect 552 21190 7114 21242
rect 7166 21190 7178 21242
rect 7230 21190 7242 21242
rect 7294 21190 7306 21242
rect 7358 21190 7370 21242
rect 7422 21190 13830 21242
rect 13882 21190 13894 21242
rect 13946 21190 13958 21242
rect 14010 21190 14022 21242
rect 14074 21190 14086 21242
rect 14138 21190 20546 21242
rect 20598 21190 20610 21242
rect 20662 21190 20674 21242
rect 20726 21190 20738 21242
rect 20790 21190 20802 21242
rect 20854 21190 27262 21242
rect 27314 21190 27326 21242
rect 27378 21190 27390 21242
rect 27442 21190 27454 21242
rect 27506 21190 27518 21242
rect 27570 21190 27576 21242
rect 552 21168 27576 21190
rect 934 21088 940 21140
rect 992 21088 998 21140
rect 1394 21137 1400 21140
rect 1213 21131 1271 21137
rect 1213 21097 1225 21131
rect 1259 21097 1271 21131
rect 1213 21091 1271 21097
rect 1381 21131 1400 21137
rect 1381 21097 1393 21131
rect 1381 21091 1400 21097
rect 1121 20995 1179 21001
rect 1121 20961 1133 20995
rect 1167 20992 1179 20995
rect 1228 20992 1256 21091
rect 1394 21088 1400 21091
rect 1452 21088 1458 21140
rect 3234 21128 3240 21140
rect 2746 21100 3240 21128
rect 1578 21020 1584 21072
rect 1636 21020 1642 21072
rect 2593 21063 2651 21069
rect 2593 21029 2605 21063
rect 2639 21060 2651 21063
rect 2746 21060 2774 21100
rect 3234 21088 3240 21100
rect 3292 21128 3298 21140
rect 9766 21128 9772 21140
rect 3292 21100 9772 21128
rect 3292 21088 3298 21100
rect 2639 21032 2774 21060
rect 2639 21029 2651 21032
rect 2593 21023 2651 21029
rect 4798 21020 4804 21072
rect 4856 21020 4862 21072
rect 5169 21063 5227 21069
rect 5169 21060 5181 21063
rect 4908 21032 5181 21060
rect 1167 20964 1256 20992
rect 2685 20995 2743 21001
rect 1167 20961 1179 20964
rect 1121 20955 1179 20961
rect 2685 20961 2697 20995
rect 2731 20992 2743 20995
rect 2866 20992 2872 21004
rect 2731 20964 2872 20992
rect 2731 20961 2743 20964
rect 2685 20955 2743 20961
rect 2866 20952 2872 20964
rect 2924 20952 2930 21004
rect 3237 20995 3295 21001
rect 3237 20961 3249 20995
rect 3283 20992 3295 20995
rect 3326 20992 3332 21004
rect 3283 20964 3332 20992
rect 3283 20961 3295 20964
rect 3237 20955 3295 20961
rect 3326 20952 3332 20964
rect 3384 20992 3390 21004
rect 3697 20995 3755 21001
rect 3697 20992 3709 20995
rect 3384 20964 3709 20992
rect 3384 20952 3390 20964
rect 3697 20961 3709 20964
rect 3743 20961 3755 20995
rect 4908 20992 4936 21032
rect 5169 21029 5181 21032
rect 5215 21029 5227 21063
rect 5169 21023 5227 21029
rect 5258 21020 5264 21072
rect 5316 21060 5322 21072
rect 6730 21060 6736 21072
rect 5316 21032 6736 21060
rect 5316 21020 5322 21032
rect 6730 21020 6736 21032
rect 6788 21020 6794 21072
rect 6932 21069 6960 21100
rect 9766 21088 9772 21100
rect 9824 21088 9830 21140
rect 14737 21131 14795 21137
rect 14737 21097 14749 21131
rect 14783 21128 14795 21131
rect 15286 21128 15292 21140
rect 14783 21100 15292 21128
rect 14783 21097 14795 21100
rect 14737 21091 14795 21097
rect 15286 21088 15292 21100
rect 15344 21088 15350 21140
rect 15746 21088 15752 21140
rect 15804 21128 15810 21140
rect 15804 21100 16712 21128
rect 15804 21088 15810 21100
rect 6917 21063 6975 21069
rect 6917 21029 6929 21063
rect 6963 21029 6975 21063
rect 6917 21023 6975 21029
rect 8478 21020 8484 21072
rect 8536 21020 8542 21072
rect 9493 21063 9551 21069
rect 8711 21029 8769 21035
rect 3697 20955 3755 20961
rect 3804 20964 4936 20992
rect 5077 20995 5135 21001
rect 842 20884 848 20936
rect 900 20924 906 20936
rect 1765 20927 1823 20933
rect 1765 20924 1777 20927
rect 900 20896 1777 20924
rect 900 20884 906 20896
rect 1765 20893 1777 20896
rect 1811 20893 1823 20927
rect 1765 20887 1823 20893
rect 2774 20884 2780 20936
rect 2832 20924 2838 20936
rect 3145 20927 3203 20933
rect 3145 20924 3157 20927
rect 2832 20896 3157 20924
rect 2832 20884 2838 20896
rect 3145 20893 3157 20896
rect 3191 20924 3203 20927
rect 3804 20924 3832 20964
rect 5077 20961 5089 20995
rect 5123 20961 5135 20995
rect 5077 20955 5135 20961
rect 3191 20896 3832 20924
rect 3191 20893 3203 20896
rect 3145 20887 3203 20893
rect 4154 20884 4160 20936
rect 4212 20884 4218 20936
rect 4338 20884 4344 20936
rect 4396 20884 4402 20936
rect 4430 20884 4436 20936
rect 4488 20884 4494 20936
rect 4522 20884 4528 20936
rect 4580 20884 4586 20936
rect 4617 20927 4675 20933
rect 4617 20893 4629 20927
rect 4663 20924 4675 20927
rect 4663 20896 4936 20924
rect 4663 20893 4675 20896
rect 4617 20887 4675 20893
rect 4908 20868 4936 20896
rect 2869 20859 2927 20865
rect 2869 20825 2881 20859
rect 2915 20856 2927 20859
rect 2958 20856 2964 20868
rect 2915 20828 2964 20856
rect 2915 20825 2927 20828
rect 2869 20819 2927 20825
rect 2958 20816 2964 20828
rect 3016 20816 3022 20868
rect 4890 20816 4896 20868
rect 4948 20816 4954 20868
rect 5092 20856 5120 20955
rect 5442 20952 5448 21004
rect 5500 20952 5506 21004
rect 6178 20952 6184 21004
rect 6236 20992 6242 21004
rect 6822 20992 6828 21004
rect 6236 20964 6828 20992
rect 6236 20952 6242 20964
rect 6822 20952 6828 20964
rect 6880 20952 6886 21004
rect 8110 20952 8116 21004
rect 8168 21001 8174 21004
rect 8168 20955 8180 21001
rect 8168 20952 8174 20955
rect 8570 20952 8576 21004
rect 8628 20992 8634 21004
rect 8711 20995 8723 21029
rect 8757 21026 8769 21029
rect 9493 21029 9505 21063
rect 9539 21060 9551 21063
rect 9858 21060 9864 21072
rect 9539 21032 9864 21060
rect 9539 21029 9551 21032
rect 8757 21004 8791 21026
rect 9493 21023 9551 21029
rect 9858 21020 9864 21032
rect 9916 21020 9922 21072
rect 11882 21060 11888 21072
rect 11532 21032 11888 21060
rect 8757 20995 8760 21004
rect 8711 20992 8760 20995
rect 8628 20964 8760 20992
rect 8628 20952 8634 20964
rect 8754 20952 8760 20964
rect 8812 20992 8818 21004
rect 9309 20995 9367 21001
rect 9309 20992 9321 20995
rect 8812 20964 9321 20992
rect 8812 20952 8818 20964
rect 9309 20961 9321 20964
rect 9355 20961 9367 20995
rect 9309 20955 9367 20961
rect 9674 20952 9680 21004
rect 9732 20952 9738 21004
rect 10321 20995 10379 21001
rect 10321 20961 10333 20995
rect 10367 20961 10379 20995
rect 10321 20955 10379 20961
rect 10505 20995 10563 21001
rect 10505 20961 10517 20995
rect 10551 20992 10563 20995
rect 10781 20995 10839 21001
rect 10781 20992 10793 20995
rect 10551 20964 10793 20992
rect 10551 20961 10563 20964
rect 10505 20955 10563 20961
rect 10781 20961 10793 20964
rect 10827 20961 10839 20995
rect 10781 20955 10839 20961
rect 5718 20884 5724 20936
rect 5776 20924 5782 20936
rect 6089 20927 6147 20933
rect 6089 20924 6101 20927
rect 5776 20896 6101 20924
rect 5776 20884 5782 20896
rect 6089 20893 6101 20896
rect 6135 20893 6147 20927
rect 6089 20887 6147 20893
rect 8389 20927 8447 20933
rect 8389 20893 8401 20927
rect 8435 20924 8447 20927
rect 8846 20924 8852 20936
rect 8435 20896 8852 20924
rect 8435 20893 8447 20896
rect 8389 20887 8447 20893
rect 8846 20884 8852 20896
rect 8904 20924 8910 20936
rect 9582 20924 9588 20936
rect 8904 20896 9588 20924
rect 8904 20884 8910 20896
rect 9582 20884 9588 20896
rect 9640 20884 9646 20936
rect 10134 20884 10140 20936
rect 10192 20884 10198 20936
rect 10336 20924 10364 20955
rect 11422 20952 11428 21004
rect 11480 20952 11486 21004
rect 10336 20896 11100 20924
rect 7006 20856 7012 20868
rect 5092 20828 7012 20856
rect 1397 20791 1455 20797
rect 1397 20757 1409 20791
rect 1443 20788 1455 20791
rect 2406 20788 2412 20800
rect 1443 20760 2412 20788
rect 1443 20757 1455 20760
rect 1397 20751 1455 20757
rect 2406 20748 2412 20760
rect 2464 20748 2470 20800
rect 3973 20791 4031 20797
rect 3973 20757 3985 20791
rect 4019 20788 4031 20791
rect 5092 20788 5120 20828
rect 7006 20816 7012 20828
rect 7064 20816 7070 20868
rect 9674 20856 9680 20868
rect 8588 20828 9680 20856
rect 4019 20760 5120 20788
rect 4019 20757 4031 20760
rect 3973 20751 4031 20757
rect 5350 20748 5356 20800
rect 5408 20788 5414 20800
rect 8588 20788 8616 20828
rect 9674 20816 9680 20828
rect 9732 20816 9738 20868
rect 10152 20856 10180 20884
rect 11072 20865 11100 20896
rect 11330 20884 11336 20936
rect 11388 20924 11394 20936
rect 11532 20933 11560 21032
rect 11882 21020 11888 21032
rect 11940 21020 11946 21072
rect 12158 21060 12164 21072
rect 12100 21029 12164 21060
rect 12100 20998 12127 21029
rect 12115 20995 12127 20998
rect 12161 21020 12164 21029
rect 12216 21020 12222 21072
rect 12161 20995 12173 21020
rect 12115 20989 12173 20995
rect 12345 20995 12403 21001
rect 12345 20992 12357 20995
rect 12268 20964 12357 20992
rect 11517 20927 11575 20933
rect 11517 20924 11529 20927
rect 11388 20896 11529 20924
rect 11388 20884 11394 20896
rect 11517 20893 11529 20896
rect 11563 20893 11575 20927
rect 11517 20887 11575 20893
rect 11698 20884 11704 20936
rect 11756 20884 11762 20936
rect 12268 20865 12296 20964
rect 12345 20961 12357 20964
rect 12391 20961 12403 20995
rect 12345 20955 12403 20961
rect 12986 20952 12992 21004
rect 13044 20952 13050 21004
rect 13078 20952 13084 21004
rect 13136 20952 13142 21004
rect 13354 20952 13360 21004
rect 13412 20952 13418 21004
rect 13630 21001 13636 21004
rect 13624 20955 13636 21001
rect 13630 20952 13636 20955
rect 13688 20952 13694 21004
rect 15197 20995 15255 21001
rect 15197 20961 15209 20995
rect 15243 20992 15255 20995
rect 15286 20992 15292 21004
rect 15243 20964 15292 20992
rect 15243 20961 15255 20964
rect 15197 20955 15255 20961
rect 15286 20952 15292 20964
rect 15344 20952 15350 21004
rect 15378 20952 15384 21004
rect 15436 20952 15442 21004
rect 15470 20952 15476 21004
rect 15528 20952 15534 21004
rect 16206 20952 16212 21004
rect 16264 20952 16270 21004
rect 16393 20995 16451 21001
rect 16393 20961 16405 20995
rect 16439 20961 16451 20995
rect 16684 20992 16712 21100
rect 17402 21088 17408 21140
rect 17460 21088 17466 21140
rect 18969 21131 19027 21137
rect 18969 21097 18981 21131
rect 19015 21097 19027 21131
rect 18969 21091 19027 21097
rect 18874 21060 18880 21072
rect 18432 21032 18880 21060
rect 16945 20995 17003 21001
rect 16945 20992 16957 20995
rect 16684 20964 16957 20992
rect 16393 20955 16451 20961
rect 16945 20961 16957 20964
rect 16991 20961 17003 20995
rect 16945 20955 17003 20961
rect 13004 20924 13032 20952
rect 12340 20896 13032 20924
rect 11057 20859 11115 20865
rect 10152 20828 11008 20856
rect 5408 20760 8616 20788
rect 5408 20748 5414 20760
rect 8662 20748 8668 20800
rect 8720 20748 8726 20800
rect 8846 20748 8852 20800
rect 8904 20748 8910 20800
rect 10226 20748 10232 20800
rect 10284 20788 10290 20800
rect 10597 20791 10655 20797
rect 10597 20788 10609 20791
rect 10284 20760 10609 20788
rect 10284 20748 10290 20760
rect 10597 20757 10609 20760
rect 10643 20757 10655 20791
rect 10980 20788 11008 20828
rect 11057 20825 11069 20859
rect 11103 20825 11115 20859
rect 12253 20859 12311 20865
rect 11057 20819 11115 20825
rect 11992 20828 12204 20856
rect 11992 20788 12020 20828
rect 10980 20760 12020 20788
rect 10597 20751 10655 20757
rect 12066 20748 12072 20800
rect 12124 20748 12130 20800
rect 12176 20788 12204 20828
rect 12253 20825 12265 20859
rect 12299 20825 12311 20859
rect 12253 20819 12311 20825
rect 12340 20788 12368 20896
rect 15010 20884 15016 20936
rect 15068 20884 15074 20936
rect 15654 20884 15660 20936
rect 15712 20924 15718 20936
rect 16408 20924 16436 20955
rect 17034 20952 17040 21004
rect 17092 20992 17098 21004
rect 17129 20995 17187 21001
rect 17129 20992 17141 20995
rect 17092 20964 17141 20992
rect 17092 20952 17098 20964
rect 17129 20961 17141 20964
rect 17175 20961 17187 20995
rect 17129 20955 17187 20961
rect 17589 20995 17647 21001
rect 17589 20961 17601 20995
rect 17635 20961 17647 20995
rect 17589 20955 17647 20961
rect 15712 20896 16436 20924
rect 17313 20927 17371 20933
rect 15712 20884 15718 20896
rect 17313 20893 17325 20927
rect 17359 20924 17371 20927
rect 17604 20924 17632 20955
rect 17678 20952 17684 21004
rect 17736 20952 17742 21004
rect 17770 20952 17776 21004
rect 17828 20952 17834 21004
rect 17954 20952 17960 21004
rect 18012 20952 18018 21004
rect 18432 21001 18460 21032
rect 18874 21020 18880 21032
rect 18932 21020 18938 21072
rect 18984 21060 19012 21091
rect 20162 21088 20168 21140
rect 20220 21128 20226 21140
rect 20441 21131 20499 21137
rect 20441 21128 20453 21131
rect 20220 21100 20453 21128
rect 20220 21088 20226 21100
rect 20441 21097 20453 21100
rect 20487 21097 20499 21131
rect 20441 21091 20499 21097
rect 19306 21063 19364 21069
rect 19306 21060 19318 21063
rect 18984 21032 19318 21060
rect 19306 21029 19318 21032
rect 19352 21029 19364 21063
rect 20456 21060 20484 21091
rect 20990 21088 20996 21140
rect 21048 21088 21054 21140
rect 21082 21088 21088 21140
rect 21140 21128 21146 21140
rect 21269 21131 21327 21137
rect 21269 21128 21281 21131
rect 21140 21100 21281 21128
rect 21140 21088 21146 21100
rect 21269 21097 21281 21100
rect 21315 21097 21327 21131
rect 21269 21091 21327 21097
rect 21358 21088 21364 21140
rect 21416 21128 21422 21140
rect 21821 21131 21879 21137
rect 21821 21128 21833 21131
rect 21416 21100 21833 21128
rect 21416 21088 21422 21100
rect 21821 21097 21833 21100
rect 21867 21097 21879 21131
rect 21821 21091 21879 21097
rect 25590 21088 25596 21140
rect 25648 21088 25654 21140
rect 22002 21060 22008 21072
rect 20456 21032 22008 21060
rect 19306 21023 19364 21029
rect 22002 21020 22008 21032
rect 22060 21020 22066 21072
rect 22278 21020 22284 21072
rect 22336 21020 22342 21072
rect 23290 21020 23296 21072
rect 23348 21020 23354 21072
rect 23474 21020 23480 21072
rect 23532 21069 23538 21072
rect 23532 21063 23551 21069
rect 23539 21029 23551 21063
rect 26421 21063 26479 21069
rect 26421 21060 26433 21063
rect 23532 21023 23551 21029
rect 24872 21032 26433 21060
rect 23532 21020 23538 21023
rect 18417 20995 18475 21001
rect 18417 20961 18429 20995
rect 18463 20961 18475 20995
rect 18417 20955 18475 20961
rect 18601 20995 18659 21001
rect 18601 20961 18613 20995
rect 18647 20961 18659 20995
rect 18601 20955 18659 20961
rect 17862 20924 17868 20936
rect 17359 20896 17868 20924
rect 17359 20893 17371 20896
rect 17313 20887 17371 20893
rect 17862 20884 17868 20896
rect 17920 20884 17926 20936
rect 17770 20816 17776 20868
rect 17828 20856 17834 20868
rect 18616 20856 18644 20955
rect 18690 20952 18696 21004
rect 18748 20952 18754 21004
rect 18785 20995 18843 21001
rect 18785 20961 18797 20995
rect 18831 20992 18843 20995
rect 20438 20992 20444 21004
rect 18831 20964 20444 20992
rect 18831 20961 18843 20964
rect 18785 20955 18843 20961
rect 20438 20952 20444 20964
rect 20496 20952 20502 21004
rect 20533 20995 20591 21001
rect 20533 20961 20545 20995
rect 20579 20992 20591 20995
rect 21729 20995 21787 21001
rect 21729 20992 21741 20995
rect 20579 20964 21741 20992
rect 20579 20961 20591 20964
rect 20533 20955 20591 20961
rect 21729 20961 21741 20964
rect 21775 20992 21787 20995
rect 22296 20992 22324 21020
rect 21775 20964 22324 20992
rect 22557 20995 22615 21001
rect 21775 20961 21787 20964
rect 21729 20955 21787 20961
rect 22557 20961 22569 20995
rect 22603 20992 22615 20995
rect 23198 20992 23204 21004
rect 22603 20964 23204 20992
rect 22603 20961 22615 20964
rect 22557 20955 22615 20961
rect 23198 20952 23204 20964
rect 23256 20952 23262 21004
rect 24872 21001 24900 21032
rect 26421 21029 26433 21032
rect 26467 21029 26479 21063
rect 26421 21023 26479 21029
rect 24857 20995 24915 21001
rect 24857 20961 24869 20995
rect 24903 20961 24915 20995
rect 25409 20995 25467 21001
rect 25409 20992 25421 20995
rect 24857 20955 24915 20961
rect 25240 20964 25421 20992
rect 18966 20884 18972 20936
rect 19024 20924 19030 20936
rect 19061 20927 19119 20933
rect 19061 20924 19073 20927
rect 19024 20896 19073 20924
rect 19024 20884 19030 20896
rect 19061 20893 19073 20896
rect 19107 20893 19119 20927
rect 19061 20887 19119 20893
rect 22281 20927 22339 20933
rect 22281 20893 22293 20927
rect 22327 20924 22339 20927
rect 22646 20924 22652 20936
rect 22327 20896 22652 20924
rect 22327 20893 22339 20896
rect 22281 20887 22339 20893
rect 22646 20884 22652 20896
rect 22704 20884 22710 20936
rect 24949 20927 25007 20933
rect 24949 20893 24961 20927
rect 24995 20924 25007 20927
rect 25038 20924 25044 20936
rect 24995 20896 25044 20924
rect 24995 20893 25007 20896
rect 24949 20887 25007 20893
rect 25038 20884 25044 20896
rect 25096 20884 25102 20936
rect 17828 20828 18736 20856
rect 17828 20816 17834 20828
rect 12176 20760 12368 20788
rect 12434 20748 12440 20800
rect 12492 20748 12498 20800
rect 13265 20791 13323 20797
rect 13265 20757 13277 20791
rect 13311 20788 13323 20791
rect 13538 20788 13544 20800
rect 13311 20760 13544 20788
rect 13311 20757 13323 20760
rect 13265 20751 13323 20757
rect 13538 20748 13544 20760
rect 13596 20748 13602 20800
rect 13722 20748 13728 20800
rect 13780 20788 13786 20800
rect 15746 20788 15752 20800
rect 13780 20760 15752 20788
rect 13780 20748 13786 20760
rect 15746 20748 15752 20760
rect 15804 20748 15810 20800
rect 16298 20748 16304 20800
rect 16356 20748 16362 20800
rect 18708 20788 18736 20828
rect 20346 20816 20352 20868
rect 20404 20856 20410 20868
rect 21361 20859 21419 20865
rect 21361 20856 21373 20859
rect 20404 20828 21373 20856
rect 20404 20816 20410 20828
rect 19794 20788 19800 20800
rect 18708 20760 19800 20788
rect 19794 20748 19800 20760
rect 19852 20748 19858 20800
rect 20640 20797 20668 20828
rect 21361 20825 21373 20828
rect 21407 20825 21419 20859
rect 21361 20819 21419 20825
rect 21450 20816 21456 20868
rect 21508 20856 21514 20868
rect 21913 20859 21971 20865
rect 21913 20856 21925 20859
rect 21508 20828 21925 20856
rect 21508 20816 21514 20828
rect 21913 20825 21925 20828
rect 21959 20825 21971 20859
rect 21913 20819 21971 20825
rect 23290 20816 23296 20868
rect 23348 20856 23354 20868
rect 25240 20865 25268 20964
rect 25409 20961 25421 20964
rect 25455 20961 25467 20995
rect 25593 20995 25651 21001
rect 25593 20992 25605 20995
rect 25409 20955 25467 20961
rect 25516 20964 25605 20992
rect 25225 20859 25283 20865
rect 23348 20828 25176 20856
rect 23348 20816 23354 20828
rect 20625 20791 20683 20797
rect 20625 20757 20637 20791
rect 20671 20757 20683 20791
rect 20625 20751 20683 20757
rect 22462 20748 22468 20800
rect 22520 20748 22526 20800
rect 23477 20791 23535 20797
rect 23477 20757 23489 20791
rect 23523 20788 23535 20791
rect 23566 20788 23572 20800
rect 23523 20760 23572 20788
rect 23523 20757 23535 20760
rect 23477 20751 23535 20757
rect 23566 20748 23572 20760
rect 23624 20748 23630 20800
rect 23661 20791 23719 20797
rect 23661 20757 23673 20791
rect 23707 20788 23719 20791
rect 23750 20788 23756 20800
rect 23707 20760 23756 20788
rect 23707 20757 23719 20760
rect 23661 20751 23719 20757
rect 23750 20748 23756 20760
rect 23808 20748 23814 20800
rect 25148 20788 25176 20828
rect 25225 20825 25237 20859
rect 25271 20825 25283 20859
rect 25225 20819 25283 20825
rect 25516 20788 25544 20964
rect 25593 20961 25605 20964
rect 25639 20961 25651 20995
rect 25593 20955 25651 20961
rect 26970 20952 26976 21004
rect 27028 20952 27034 21004
rect 25148 20760 25544 20788
rect 552 20698 27416 20720
rect 552 20646 3756 20698
rect 3808 20646 3820 20698
rect 3872 20646 3884 20698
rect 3936 20646 3948 20698
rect 4000 20646 4012 20698
rect 4064 20646 10472 20698
rect 10524 20646 10536 20698
rect 10588 20646 10600 20698
rect 10652 20646 10664 20698
rect 10716 20646 10728 20698
rect 10780 20646 17188 20698
rect 17240 20646 17252 20698
rect 17304 20646 17316 20698
rect 17368 20646 17380 20698
rect 17432 20646 17444 20698
rect 17496 20646 23904 20698
rect 23956 20646 23968 20698
rect 24020 20646 24032 20698
rect 24084 20646 24096 20698
rect 24148 20646 24160 20698
rect 24212 20646 27416 20698
rect 552 20624 27416 20646
rect 1857 20587 1915 20593
rect 1857 20553 1869 20587
rect 1903 20584 1915 20587
rect 2314 20584 2320 20596
rect 1903 20556 2320 20584
rect 1903 20553 1915 20556
rect 1857 20547 1915 20553
rect 2314 20544 2320 20556
rect 2372 20544 2378 20596
rect 2501 20587 2559 20593
rect 2501 20553 2513 20587
rect 2547 20584 2559 20587
rect 2682 20584 2688 20596
rect 2547 20556 2688 20584
rect 2547 20553 2559 20556
rect 2501 20547 2559 20553
rect 2682 20544 2688 20556
rect 2740 20544 2746 20596
rect 3881 20587 3939 20593
rect 3881 20553 3893 20587
rect 3927 20584 3939 20587
rect 4433 20587 4491 20593
rect 3927 20556 4016 20584
rect 3927 20553 3939 20556
rect 3881 20547 3939 20553
rect 2038 20408 2044 20460
rect 2096 20448 2102 20460
rect 2777 20451 2835 20457
rect 2777 20448 2789 20451
rect 2096 20420 2360 20448
rect 2096 20408 2102 20420
rect 2133 20383 2191 20389
rect 2133 20349 2145 20383
rect 2179 20380 2191 20383
rect 2222 20380 2228 20392
rect 2179 20352 2228 20380
rect 2179 20349 2191 20352
rect 2133 20343 2191 20349
rect 2222 20340 2228 20352
rect 2280 20340 2286 20392
rect 2332 20389 2360 20420
rect 2424 20420 2789 20448
rect 2424 20392 2452 20420
rect 2777 20417 2789 20420
rect 2823 20417 2835 20451
rect 2777 20411 2835 20417
rect 2317 20383 2375 20389
rect 2317 20349 2329 20383
rect 2363 20349 2375 20383
rect 2317 20343 2375 20349
rect 2406 20340 2412 20392
rect 2464 20340 2470 20392
rect 2593 20383 2651 20389
rect 2593 20349 2605 20383
rect 2639 20349 2651 20383
rect 2593 20343 2651 20349
rect 1578 20272 1584 20324
rect 1636 20312 1642 20324
rect 2041 20315 2099 20321
rect 2041 20312 2053 20315
rect 1636 20284 2053 20312
rect 1636 20272 1642 20284
rect 2041 20281 2053 20284
rect 2087 20281 2099 20315
rect 2608 20312 2636 20343
rect 2682 20340 2688 20392
rect 2740 20340 2746 20392
rect 2869 20383 2927 20389
rect 2869 20349 2881 20383
rect 2915 20349 2927 20383
rect 2869 20343 2927 20349
rect 2774 20312 2780 20324
rect 2608 20284 2780 20312
rect 2041 20275 2099 20281
rect 2774 20272 2780 20284
rect 2832 20272 2838 20324
rect 1210 20204 1216 20256
rect 1268 20244 1274 20256
rect 1854 20253 1860 20256
rect 1673 20247 1731 20253
rect 1673 20244 1685 20247
rect 1268 20216 1685 20244
rect 1268 20204 1274 20216
rect 1673 20213 1685 20216
rect 1719 20213 1731 20247
rect 1673 20207 1731 20213
rect 1841 20247 1860 20253
rect 1841 20213 1853 20247
rect 1912 20244 1918 20256
rect 2133 20247 2191 20253
rect 2133 20244 2145 20247
rect 1912 20216 2145 20244
rect 1841 20207 1860 20213
rect 1854 20204 1860 20207
rect 1912 20204 1918 20216
rect 2133 20213 2145 20216
rect 2179 20213 2191 20247
rect 2133 20207 2191 20213
rect 2498 20204 2504 20256
rect 2556 20244 2562 20256
rect 2884 20244 2912 20343
rect 3326 20340 3332 20392
rect 3384 20380 3390 20392
rect 3605 20383 3663 20389
rect 3605 20380 3617 20383
rect 3384 20352 3617 20380
rect 3384 20340 3390 20352
rect 3605 20349 3617 20352
rect 3651 20349 3663 20383
rect 3605 20343 3663 20349
rect 2556 20216 2912 20244
rect 2556 20204 2562 20216
rect 3786 20204 3792 20256
rect 3844 20244 3850 20256
rect 3988 20244 4016 20556
rect 4433 20553 4445 20587
rect 4479 20584 4491 20587
rect 4522 20584 4528 20596
rect 4479 20556 4528 20584
rect 4479 20553 4491 20556
rect 4433 20547 4491 20553
rect 4522 20544 4528 20556
rect 4580 20544 4586 20596
rect 5077 20587 5135 20593
rect 5077 20553 5089 20587
rect 5123 20584 5135 20587
rect 5258 20584 5264 20596
rect 5123 20556 5264 20584
rect 5123 20553 5135 20556
rect 5077 20547 5135 20553
rect 5258 20544 5264 20556
rect 5316 20544 5322 20596
rect 6730 20544 6736 20596
rect 6788 20584 6794 20596
rect 7009 20587 7067 20593
rect 7009 20584 7021 20587
rect 6788 20556 7021 20584
rect 6788 20544 6794 20556
rect 7009 20553 7021 20556
rect 7055 20553 7067 20587
rect 7009 20547 7067 20553
rect 7929 20587 7987 20593
rect 7929 20553 7941 20587
rect 7975 20584 7987 20587
rect 8110 20584 8116 20596
rect 7975 20556 8116 20584
rect 7975 20553 7987 20556
rect 7929 20547 7987 20553
rect 8110 20544 8116 20556
rect 8168 20544 8174 20596
rect 8389 20587 8447 20593
rect 8389 20553 8401 20587
rect 8435 20584 8447 20587
rect 8478 20584 8484 20596
rect 8435 20556 8484 20584
rect 8435 20553 8447 20556
rect 8389 20547 8447 20553
rect 8478 20544 8484 20556
rect 8536 20544 8542 20596
rect 11330 20544 11336 20596
rect 11388 20544 11394 20596
rect 13630 20544 13636 20596
rect 13688 20584 13694 20596
rect 13725 20587 13783 20593
rect 13725 20584 13737 20587
rect 13688 20556 13737 20584
rect 13688 20544 13694 20556
rect 13725 20553 13737 20556
rect 13771 20553 13783 20587
rect 13725 20547 13783 20553
rect 15378 20544 15384 20596
rect 15436 20584 15442 20596
rect 15746 20584 15752 20596
rect 15436 20556 15752 20584
rect 15436 20544 15442 20556
rect 15746 20544 15752 20556
rect 15804 20584 15810 20596
rect 15933 20587 15991 20593
rect 15933 20584 15945 20587
rect 15804 20556 15945 20584
rect 15804 20544 15810 20556
rect 15933 20553 15945 20556
rect 15979 20553 15991 20587
rect 19886 20584 19892 20596
rect 15933 20547 15991 20553
rect 16408 20556 19892 20584
rect 4338 20476 4344 20528
rect 4396 20516 4402 20528
rect 4709 20519 4767 20525
rect 4709 20516 4721 20519
rect 4396 20488 4721 20516
rect 4396 20476 4402 20488
rect 4709 20485 4721 20488
rect 4755 20485 4767 20519
rect 4709 20479 4767 20485
rect 15838 20476 15844 20528
rect 15896 20516 15902 20528
rect 16408 20516 16436 20556
rect 19886 20544 19892 20556
rect 19944 20544 19950 20596
rect 22094 20584 22100 20596
rect 19996 20556 22100 20584
rect 15896 20488 16436 20516
rect 15896 20476 15902 20488
rect 17770 20476 17776 20528
rect 17828 20516 17834 20528
rect 17865 20519 17923 20525
rect 17865 20516 17877 20519
rect 17828 20488 17877 20516
rect 17828 20476 17834 20488
rect 17865 20485 17877 20488
rect 17911 20485 17923 20519
rect 17865 20479 17923 20485
rect 4065 20451 4123 20457
rect 4065 20417 4077 20451
rect 4111 20417 4123 20451
rect 4065 20411 4123 20417
rect 4080 20380 4108 20411
rect 4154 20408 4160 20460
rect 4212 20448 4218 20460
rect 5169 20451 5227 20457
rect 4212 20420 4568 20448
rect 4212 20408 4218 20420
rect 4246 20380 4252 20392
rect 4080 20352 4252 20380
rect 4246 20340 4252 20352
rect 4304 20380 4310 20392
rect 4540 20389 4568 20420
rect 5169 20417 5181 20451
rect 5215 20448 5227 20451
rect 5442 20448 5448 20460
rect 5215 20420 5448 20448
rect 5215 20417 5227 20420
rect 5169 20411 5227 20417
rect 5442 20408 5448 20420
rect 5500 20408 5506 20460
rect 13354 20408 13360 20460
rect 13412 20448 13418 20460
rect 14277 20451 14335 20457
rect 14277 20448 14289 20451
rect 13412 20420 14289 20448
rect 13412 20408 13418 20420
rect 14277 20417 14289 20420
rect 14323 20417 14335 20451
rect 14277 20411 14335 20417
rect 17313 20451 17371 20457
rect 17313 20417 17325 20451
rect 17359 20448 17371 20451
rect 17954 20448 17960 20460
rect 17359 20420 17960 20448
rect 17359 20417 17371 20420
rect 17313 20411 17371 20417
rect 17954 20408 17960 20420
rect 18012 20408 18018 20460
rect 18690 20408 18696 20460
rect 18748 20448 18754 20460
rect 19337 20451 19395 20457
rect 19337 20448 19349 20451
rect 18748 20420 19349 20448
rect 18748 20408 18754 20420
rect 19337 20417 19349 20420
rect 19383 20448 19395 20451
rect 19996 20448 20024 20556
rect 22094 20544 22100 20556
rect 22152 20544 22158 20596
rect 23385 20587 23443 20593
rect 23385 20553 23397 20587
rect 23431 20584 23443 20587
rect 23474 20584 23480 20596
rect 23431 20556 23480 20584
rect 23431 20553 23443 20556
rect 23385 20547 23443 20553
rect 23474 20544 23480 20556
rect 23532 20544 23538 20596
rect 24213 20519 24271 20525
rect 24213 20516 24225 20519
rect 20364 20488 21772 20516
rect 19383 20420 20024 20448
rect 19383 20417 19395 20420
rect 19337 20411 19395 20417
rect 20070 20408 20076 20460
rect 20128 20448 20134 20460
rect 20364 20457 20392 20488
rect 21744 20460 21772 20488
rect 23676 20488 24225 20516
rect 20349 20451 20407 20457
rect 20128 20420 20300 20448
rect 20128 20408 20134 20420
rect 4341 20383 4399 20389
rect 4341 20380 4353 20383
rect 4304 20352 4353 20380
rect 4304 20340 4310 20352
rect 4341 20349 4353 20352
rect 4387 20349 4399 20383
rect 4341 20343 4399 20349
rect 4525 20383 4583 20389
rect 4525 20349 4537 20383
rect 4571 20349 4583 20383
rect 4525 20343 4583 20349
rect 4890 20340 4896 20392
rect 4948 20340 4954 20392
rect 5629 20383 5687 20389
rect 5629 20349 5641 20383
rect 5675 20380 5687 20383
rect 5718 20380 5724 20392
rect 5675 20352 5724 20380
rect 5675 20349 5687 20352
rect 5629 20343 5687 20349
rect 5718 20340 5724 20352
rect 5776 20340 5782 20392
rect 7466 20340 7472 20392
rect 7524 20340 7530 20392
rect 7745 20383 7803 20389
rect 7745 20349 7757 20383
rect 7791 20380 7803 20383
rect 8386 20380 8392 20392
rect 7791 20352 8392 20380
rect 7791 20349 7803 20352
rect 7745 20343 7803 20349
rect 8386 20340 8392 20352
rect 8444 20340 8450 20392
rect 9674 20340 9680 20392
rect 9732 20380 9738 20392
rect 10226 20389 10232 20392
rect 9769 20383 9827 20389
rect 9769 20380 9781 20383
rect 9732 20352 9781 20380
rect 9732 20340 9738 20352
rect 9769 20349 9781 20352
rect 9815 20380 9827 20383
rect 9953 20383 10011 20389
rect 9953 20380 9965 20383
rect 9815 20352 9965 20380
rect 9815 20349 9827 20352
rect 9769 20343 9827 20349
rect 9953 20349 9965 20352
rect 9999 20349 10011 20383
rect 10220 20380 10232 20389
rect 10187 20352 10232 20380
rect 9953 20343 10011 20349
rect 10220 20343 10232 20352
rect 10226 20340 10232 20343
rect 10284 20340 10290 20392
rect 13538 20340 13544 20392
rect 13596 20340 13602 20392
rect 14001 20383 14059 20389
rect 14001 20349 14013 20383
rect 14047 20380 14059 20383
rect 14826 20380 14832 20392
rect 14047 20352 14832 20380
rect 14047 20349 14059 20352
rect 14001 20343 14059 20349
rect 14826 20340 14832 20352
rect 14884 20340 14890 20392
rect 16298 20340 16304 20392
rect 16356 20380 16362 20392
rect 17046 20383 17104 20389
rect 17046 20380 17058 20383
rect 16356 20352 17058 20380
rect 16356 20340 16362 20352
rect 17046 20349 17058 20352
rect 17092 20349 17104 20383
rect 17046 20343 17104 20349
rect 17681 20383 17739 20389
rect 17681 20349 17693 20383
rect 17727 20349 17739 20383
rect 17681 20343 17739 20349
rect 5534 20272 5540 20324
rect 5592 20312 5598 20324
rect 5874 20315 5932 20321
rect 5874 20312 5886 20315
rect 5592 20284 5886 20312
rect 5592 20272 5598 20284
rect 5874 20281 5886 20284
rect 5920 20281 5932 20315
rect 8478 20312 8484 20324
rect 5874 20275 5932 20281
rect 6012 20284 8484 20312
rect 6012 20244 6040 20284
rect 8478 20272 8484 20284
rect 8536 20272 8542 20324
rect 9030 20272 9036 20324
rect 9088 20312 9094 20324
rect 9502 20315 9560 20321
rect 9502 20312 9514 20315
rect 9088 20284 9514 20312
rect 9088 20272 9094 20284
rect 9502 20281 9514 20284
rect 9548 20281 9560 20315
rect 14522 20315 14580 20321
rect 14522 20312 14534 20315
rect 9502 20275 9560 20281
rect 14200 20284 14534 20312
rect 3844 20216 6040 20244
rect 7561 20247 7619 20253
rect 3844 20204 3850 20216
rect 7561 20213 7573 20247
rect 7607 20244 7619 20247
rect 7926 20244 7932 20256
rect 7607 20216 7932 20244
rect 7607 20213 7619 20216
rect 7561 20207 7619 20213
rect 7926 20204 7932 20216
rect 7984 20244 7990 20256
rect 12618 20244 12624 20256
rect 7984 20216 12624 20244
rect 7984 20204 7990 20216
rect 12618 20204 12624 20216
rect 12676 20204 12682 20256
rect 14200 20253 14228 20284
rect 14522 20281 14534 20284
rect 14568 20281 14580 20315
rect 17696 20312 17724 20343
rect 17862 20340 17868 20392
rect 17920 20380 17926 20392
rect 19613 20383 19671 20389
rect 19613 20380 19625 20383
rect 17920 20352 19625 20380
rect 17920 20340 17926 20352
rect 19613 20349 19625 20352
rect 19659 20349 19671 20383
rect 19613 20343 19671 20349
rect 18322 20312 18328 20324
rect 17696 20284 18328 20312
rect 14522 20275 14580 20281
rect 18322 20272 18328 20284
rect 18380 20312 18386 20324
rect 19242 20312 19248 20324
rect 18380 20284 19248 20312
rect 18380 20272 18386 20284
rect 19242 20272 19248 20284
rect 19300 20272 19306 20324
rect 19628 20312 19656 20343
rect 19702 20340 19708 20392
rect 19760 20340 19766 20392
rect 19981 20383 20039 20389
rect 19981 20349 19993 20383
rect 20027 20380 20039 20383
rect 20162 20380 20168 20392
rect 20027 20352 20168 20380
rect 20027 20349 20039 20352
rect 19981 20343 20039 20349
rect 20162 20340 20168 20352
rect 20220 20340 20226 20392
rect 20272 20380 20300 20420
rect 20349 20417 20361 20451
rect 20395 20417 20407 20451
rect 20349 20411 20407 20417
rect 20901 20451 20959 20457
rect 20901 20417 20913 20451
rect 20947 20448 20959 20451
rect 20947 20420 21588 20448
rect 20947 20417 20959 20420
rect 20901 20411 20959 20417
rect 21082 20380 21088 20392
rect 20272 20352 21088 20380
rect 21082 20340 21088 20352
rect 21140 20340 21146 20392
rect 21177 20383 21235 20389
rect 21177 20349 21189 20383
rect 21223 20380 21235 20383
rect 21450 20380 21456 20392
rect 21223 20352 21456 20380
rect 21223 20349 21235 20352
rect 21177 20343 21235 20349
rect 19628 20284 19748 20312
rect 14185 20247 14243 20253
rect 14185 20213 14197 20247
rect 14231 20213 14243 20247
rect 14185 20207 14243 20213
rect 15286 20204 15292 20256
rect 15344 20244 15350 20256
rect 15657 20247 15715 20253
rect 15657 20244 15669 20247
rect 15344 20216 15669 20244
rect 15344 20204 15350 20216
rect 15657 20213 15669 20216
rect 15703 20213 15715 20247
rect 15657 20207 15715 20213
rect 18046 20204 18052 20256
rect 18104 20244 18110 20256
rect 18693 20247 18751 20253
rect 18693 20244 18705 20247
rect 18104 20216 18705 20244
rect 18104 20204 18110 20216
rect 18693 20213 18705 20216
rect 18739 20213 18751 20247
rect 18693 20207 18751 20213
rect 19426 20204 19432 20256
rect 19484 20204 19490 20256
rect 19720 20244 19748 20284
rect 19794 20272 19800 20324
rect 19852 20272 19858 20324
rect 20438 20312 20444 20324
rect 19904 20284 20444 20312
rect 19904 20244 19932 20284
rect 20438 20272 20444 20284
rect 20496 20312 20502 20324
rect 21192 20312 21220 20343
rect 21450 20340 21456 20352
rect 21508 20340 21514 20392
rect 21560 20389 21588 20420
rect 21726 20408 21732 20460
rect 21784 20408 21790 20460
rect 22462 20448 22468 20460
rect 21836 20420 22468 20448
rect 21545 20383 21603 20389
rect 21545 20349 21557 20383
rect 21591 20349 21603 20383
rect 21545 20343 21603 20349
rect 21634 20340 21640 20392
rect 21692 20380 21698 20392
rect 21836 20380 21864 20420
rect 22462 20408 22468 20420
rect 22520 20408 22526 20460
rect 21692 20352 21864 20380
rect 21692 20340 21698 20352
rect 21910 20340 21916 20392
rect 21968 20340 21974 20392
rect 22002 20340 22008 20392
rect 22060 20340 22066 20392
rect 22189 20383 22247 20389
rect 22189 20349 22201 20383
rect 22235 20380 22247 20383
rect 22281 20383 22339 20389
rect 22281 20380 22293 20383
rect 22235 20352 22293 20380
rect 22235 20349 22247 20352
rect 22189 20343 22247 20349
rect 22281 20349 22293 20352
rect 22327 20349 22339 20383
rect 22281 20343 22339 20349
rect 22370 20340 22376 20392
rect 22428 20340 22434 20392
rect 22554 20340 22560 20392
rect 22612 20340 22618 20392
rect 22738 20340 22744 20392
rect 22796 20380 22802 20392
rect 23676 20389 23704 20488
rect 24213 20485 24225 20488
rect 24259 20485 24271 20519
rect 24213 20479 24271 20485
rect 23017 20383 23075 20389
rect 23017 20380 23029 20383
rect 22796 20352 23029 20380
rect 22796 20340 22802 20352
rect 23017 20349 23029 20352
rect 23063 20380 23075 20383
rect 23477 20383 23535 20389
rect 23477 20380 23489 20383
rect 23063 20352 23489 20380
rect 23063 20349 23075 20352
rect 23017 20343 23075 20349
rect 23477 20349 23489 20352
rect 23523 20349 23535 20383
rect 23477 20343 23535 20349
rect 23661 20383 23719 20389
rect 23661 20349 23673 20383
rect 23707 20349 23719 20383
rect 23661 20343 23719 20349
rect 20496 20284 21220 20312
rect 20496 20272 20502 20284
rect 21266 20272 21272 20324
rect 21324 20272 21330 20324
rect 21361 20315 21419 20321
rect 21361 20281 21373 20315
rect 21407 20312 21419 20315
rect 21407 20284 21588 20312
rect 21407 20281 21419 20284
rect 21361 20275 21419 20281
rect 21560 20256 21588 20284
rect 22830 20272 22836 20324
rect 22888 20312 22894 20324
rect 23198 20312 23204 20324
rect 22888 20284 23204 20312
rect 22888 20272 22894 20284
rect 23198 20272 23204 20284
rect 23256 20312 23262 20324
rect 23676 20312 23704 20343
rect 23750 20340 23756 20392
rect 23808 20380 23814 20392
rect 23937 20383 23995 20389
rect 23937 20380 23949 20383
rect 23808 20352 23949 20380
rect 23808 20340 23814 20352
rect 23937 20349 23949 20352
rect 23983 20349 23995 20383
rect 23937 20343 23995 20349
rect 25593 20383 25651 20389
rect 25593 20349 25605 20383
rect 25639 20349 25651 20383
rect 25593 20343 25651 20349
rect 25326 20315 25384 20321
rect 25326 20312 25338 20315
rect 23256 20284 23704 20312
rect 24136 20284 25338 20312
rect 23256 20272 23262 20284
rect 19720 20216 19932 20244
rect 20990 20204 20996 20256
rect 21048 20204 21054 20256
rect 21082 20204 21088 20256
rect 21140 20244 21146 20256
rect 21542 20244 21548 20256
rect 21140 20216 21548 20244
rect 21140 20204 21146 20216
rect 21542 20204 21548 20216
rect 21600 20204 21606 20256
rect 22738 20204 22744 20256
rect 22796 20204 22802 20256
rect 23566 20204 23572 20256
rect 23624 20204 23630 20256
rect 24136 20253 24164 20284
rect 25326 20281 25338 20284
rect 25372 20281 25384 20315
rect 25608 20312 25636 20343
rect 25866 20340 25872 20392
rect 25924 20380 25930 20392
rect 25961 20383 26019 20389
rect 25961 20380 25973 20383
rect 25924 20352 25973 20380
rect 25924 20340 25930 20352
rect 25961 20349 25973 20352
rect 26007 20349 26019 20383
rect 25961 20343 26019 20349
rect 26789 20315 26847 20321
rect 26789 20312 26801 20315
rect 25608 20284 26801 20312
rect 25326 20275 25384 20281
rect 26789 20281 26801 20284
rect 26835 20312 26847 20315
rect 27062 20312 27068 20324
rect 26835 20284 27068 20312
rect 26835 20281 26847 20284
rect 26789 20275 26847 20281
rect 27062 20272 27068 20284
rect 27120 20272 27126 20324
rect 24121 20247 24179 20253
rect 24121 20213 24133 20247
rect 24167 20213 24179 20247
rect 24121 20207 24179 20213
rect 552 20154 27576 20176
rect 552 20102 7114 20154
rect 7166 20102 7178 20154
rect 7230 20102 7242 20154
rect 7294 20102 7306 20154
rect 7358 20102 7370 20154
rect 7422 20102 13830 20154
rect 13882 20102 13894 20154
rect 13946 20102 13958 20154
rect 14010 20102 14022 20154
rect 14074 20102 14086 20154
rect 14138 20102 20546 20154
rect 20598 20102 20610 20154
rect 20662 20102 20674 20154
rect 20726 20102 20738 20154
rect 20790 20102 20802 20154
rect 20854 20102 27262 20154
rect 27314 20102 27326 20154
rect 27378 20102 27390 20154
rect 27442 20102 27454 20154
rect 27506 20102 27518 20154
rect 27570 20102 27576 20154
rect 552 20080 27576 20102
rect 2222 20000 2228 20052
rect 2280 20000 2286 20052
rect 2314 20000 2320 20052
rect 2372 20000 2378 20052
rect 4157 20043 4215 20049
rect 4157 20009 4169 20043
rect 4203 20040 4215 20043
rect 4430 20040 4436 20052
rect 4203 20012 4436 20040
rect 4203 20009 4215 20012
rect 4157 20003 4215 20009
rect 4430 20000 4436 20012
rect 4488 20000 4494 20052
rect 9030 20000 9036 20052
rect 9088 20000 9094 20052
rect 10962 20040 10968 20052
rect 9800 20012 10968 20040
rect 2240 19972 2268 20000
rect 2501 19975 2559 19981
rect 2501 19972 2513 19975
rect 2240 19944 2513 19972
rect 2501 19941 2513 19944
rect 2547 19972 2559 19975
rect 2547 19944 3372 19972
rect 2547 19941 2559 19944
rect 2501 19935 2559 19941
rect 3344 19916 3372 19944
rect 3694 19932 3700 19984
rect 3752 19972 3758 19984
rect 3881 19975 3939 19981
rect 3881 19972 3893 19975
rect 3752 19944 3893 19972
rect 3752 19932 3758 19944
rect 3881 19941 3893 19944
rect 3927 19941 3939 19975
rect 3881 19935 3939 19941
rect 1118 19913 1124 19916
rect 1112 19867 1124 19913
rect 1118 19864 1124 19867
rect 1176 19864 1182 19916
rect 2038 19864 2044 19916
rect 2096 19904 2102 19916
rect 2682 19904 2688 19916
rect 2096 19876 2688 19904
rect 2096 19864 2102 19876
rect 2682 19864 2688 19876
rect 2740 19864 2746 19916
rect 2774 19864 2780 19916
rect 2832 19864 2838 19916
rect 3326 19864 3332 19916
rect 3384 19864 3390 19916
rect 3421 19907 3479 19913
rect 3421 19873 3433 19907
rect 3467 19904 3479 19907
rect 3605 19907 3663 19913
rect 3605 19904 3617 19907
rect 3467 19876 3617 19904
rect 3467 19873 3479 19876
rect 3421 19867 3479 19873
rect 3605 19873 3617 19876
rect 3651 19873 3663 19907
rect 3605 19867 3663 19873
rect 3786 19864 3792 19916
rect 3844 19864 3850 19916
rect 3973 19907 4031 19913
rect 3973 19873 3985 19907
rect 4019 19904 4031 19907
rect 4448 19904 4476 20000
rect 8665 19975 8723 19981
rect 8665 19941 8677 19975
rect 8711 19972 8723 19975
rect 9800 19972 9828 20012
rect 10962 20000 10968 20012
rect 11020 20040 11026 20052
rect 12526 20040 12532 20052
rect 11020 20012 12532 20040
rect 11020 20000 11026 20012
rect 12526 20000 12532 20012
rect 12584 20000 12590 20052
rect 14826 20000 14832 20052
rect 14884 20000 14890 20052
rect 15013 20043 15071 20049
rect 15013 20009 15025 20043
rect 15059 20040 15071 20043
rect 15378 20040 15384 20052
rect 15059 20012 15384 20040
rect 15059 20009 15071 20012
rect 15013 20003 15071 20009
rect 15378 20000 15384 20012
rect 15436 20040 15442 20052
rect 15654 20040 15660 20052
rect 15436 20012 15660 20040
rect 15436 20000 15442 20012
rect 15654 20000 15660 20012
rect 15712 20000 15718 20052
rect 15765 20043 15823 20049
rect 15765 20040 15777 20043
rect 15764 20009 15777 20040
rect 15811 20009 15823 20043
rect 15764 20003 15823 20009
rect 12434 19972 12440 19984
rect 8711 19944 9828 19972
rect 9876 19944 12440 19972
rect 8711 19941 8723 19944
rect 8665 19935 8723 19941
rect 9876 19916 9904 19944
rect 4617 19907 4675 19913
rect 4617 19904 4629 19907
rect 4019 19876 4384 19904
rect 4448 19876 4629 19904
rect 4019 19873 4031 19876
rect 3973 19867 4031 19873
rect 842 19796 848 19848
rect 900 19796 906 19848
rect 4246 19728 4252 19780
rect 4304 19768 4310 19780
rect 4356 19768 4384 19876
rect 4617 19873 4629 19876
rect 4663 19873 4675 19907
rect 4617 19867 4675 19873
rect 4706 19864 4712 19916
rect 4764 19864 4770 19916
rect 4985 19907 5043 19913
rect 4985 19873 4997 19907
rect 5031 19904 5043 19907
rect 5074 19904 5080 19916
rect 5031 19876 5080 19904
rect 5031 19873 5043 19876
rect 4985 19867 5043 19873
rect 5074 19864 5080 19876
rect 5132 19864 5138 19916
rect 6172 19907 6230 19913
rect 6172 19873 6184 19907
rect 6218 19904 6230 19907
rect 6730 19904 6736 19916
rect 6218 19876 6736 19904
rect 6218 19873 6230 19876
rect 6172 19867 6230 19873
rect 6730 19864 6736 19876
rect 6788 19864 6794 19916
rect 7466 19864 7472 19916
rect 7524 19904 7530 19916
rect 8573 19907 8631 19913
rect 8573 19904 8585 19907
rect 7524 19876 8585 19904
rect 7524 19864 7530 19876
rect 8573 19873 8585 19876
rect 8619 19873 8631 19907
rect 8573 19867 8631 19873
rect 4430 19796 4436 19848
rect 4488 19836 4494 19848
rect 4890 19836 4896 19848
rect 4488 19808 4896 19836
rect 4488 19796 4494 19808
rect 4890 19796 4896 19808
rect 4948 19796 4954 19848
rect 5718 19796 5724 19848
rect 5776 19836 5782 19848
rect 5905 19839 5963 19845
rect 5905 19836 5917 19839
rect 5776 19808 5917 19836
rect 5776 19796 5782 19808
rect 5905 19805 5917 19808
rect 5951 19805 5963 19839
rect 7745 19839 7803 19845
rect 7745 19836 7757 19839
rect 5905 19799 5963 19805
rect 7300 19808 7757 19836
rect 7300 19777 7328 19808
rect 7745 19805 7757 19808
rect 7791 19805 7803 19839
rect 8588 19836 8616 19867
rect 8846 19864 8852 19916
rect 8904 19864 8910 19916
rect 9493 19907 9551 19913
rect 9493 19873 9505 19907
rect 9539 19873 9551 19907
rect 9493 19867 9551 19873
rect 9677 19907 9735 19913
rect 9677 19873 9689 19907
rect 9723 19904 9735 19907
rect 9858 19904 9864 19916
rect 9723 19876 9864 19904
rect 9723 19873 9735 19876
rect 9677 19867 9735 19873
rect 9309 19839 9367 19845
rect 9309 19836 9321 19839
rect 8588 19808 9321 19836
rect 7745 19799 7803 19805
rect 9309 19805 9321 19808
rect 9355 19805 9367 19839
rect 9508 19836 9536 19867
rect 9858 19864 9864 19876
rect 9916 19864 9922 19916
rect 11333 19907 11391 19913
rect 11333 19873 11345 19907
rect 11379 19904 11391 19907
rect 11422 19904 11428 19916
rect 11379 19876 11428 19904
rect 11379 19873 11391 19876
rect 11333 19867 11391 19873
rect 11422 19864 11428 19876
rect 11480 19864 11486 19916
rect 11808 19913 11836 19944
rect 12434 19932 12440 19944
rect 12492 19932 12498 19984
rect 12697 19975 12755 19981
rect 12697 19941 12709 19975
rect 12743 19972 12755 19975
rect 12802 19972 12808 19984
rect 12743 19944 12808 19972
rect 12743 19941 12755 19944
rect 12697 19935 12755 19941
rect 12802 19932 12808 19944
rect 12860 19932 12866 19984
rect 12897 19975 12955 19981
rect 12897 19941 12909 19975
rect 12943 19972 12955 19975
rect 12989 19975 13047 19981
rect 12989 19972 13001 19975
rect 12943 19944 13001 19972
rect 12943 19941 12955 19944
rect 12897 19935 12955 19941
rect 12989 19941 13001 19944
rect 13035 19941 13047 19975
rect 12989 19935 13047 19941
rect 15286 19932 15292 19984
rect 15344 19972 15350 19984
rect 15565 19975 15623 19981
rect 15565 19972 15577 19975
rect 15344 19944 15577 19972
rect 15344 19932 15350 19944
rect 15565 19941 15577 19944
rect 15611 19941 15623 19975
rect 15764 19972 15792 20003
rect 18690 20000 18696 20052
rect 18748 20000 18754 20052
rect 19794 20000 19800 20052
rect 19852 20040 19858 20052
rect 21082 20040 21088 20052
rect 19852 20012 21088 20040
rect 19852 20000 19858 20012
rect 21082 20000 21088 20012
rect 21140 20000 21146 20052
rect 21634 20040 21640 20052
rect 21284 20012 21640 20040
rect 17954 19972 17960 19984
rect 15565 19935 15623 19941
rect 15672 19944 15792 19972
rect 17328 19944 17960 19972
rect 15672 19916 15700 19944
rect 11793 19907 11851 19913
rect 11793 19873 11805 19907
rect 11839 19873 11851 19907
rect 11793 19867 11851 19873
rect 12069 19907 12127 19913
rect 12069 19873 12081 19907
rect 12115 19904 12127 19907
rect 12342 19904 12348 19916
rect 12115 19876 12348 19904
rect 12115 19873 12127 19876
rect 12069 19867 12127 19873
rect 12342 19864 12348 19876
rect 12400 19904 12406 19916
rect 13909 19907 13967 19913
rect 12400 19876 13768 19904
rect 12400 19864 12406 19876
rect 10042 19836 10048 19848
rect 9508 19808 10048 19836
rect 9309 19799 9367 19805
rect 10042 19796 10048 19808
rect 10100 19836 10106 19848
rect 10870 19836 10876 19848
rect 10100 19808 10876 19836
rect 10100 19796 10106 19808
rect 10870 19796 10876 19808
rect 10928 19796 10934 19848
rect 11149 19839 11207 19845
rect 11149 19805 11161 19839
rect 11195 19805 11207 19839
rect 11149 19799 11207 19805
rect 11241 19839 11299 19845
rect 11241 19805 11253 19839
rect 11287 19836 11299 19839
rect 12710 19836 12716 19848
rect 11287 19808 12716 19836
rect 11287 19805 11299 19808
rect 11241 19799 11299 19805
rect 7285 19771 7343 19777
rect 4304 19740 5764 19768
rect 4304 19728 4310 19740
rect 2958 19660 2964 19712
rect 3016 19660 3022 19712
rect 5077 19703 5135 19709
rect 5077 19669 5089 19703
rect 5123 19700 5135 19703
rect 5626 19700 5632 19712
rect 5123 19672 5632 19700
rect 5123 19669 5135 19672
rect 5077 19663 5135 19669
rect 5626 19660 5632 19672
rect 5684 19660 5690 19712
rect 5736 19700 5764 19740
rect 7285 19737 7297 19771
rect 7331 19737 7343 19771
rect 11164 19768 11192 19799
rect 12710 19796 12716 19808
rect 12768 19796 12774 19848
rect 12894 19796 12900 19848
rect 12952 19836 12958 19848
rect 13541 19839 13599 19845
rect 13541 19836 13553 19839
rect 12952 19808 13553 19836
rect 12952 19796 12958 19808
rect 13541 19805 13553 19808
rect 13587 19836 13599 19839
rect 13630 19836 13636 19848
rect 13587 19808 13636 19836
rect 13587 19805 13599 19808
rect 13541 19799 13599 19805
rect 13630 19796 13636 19808
rect 13688 19796 13694 19848
rect 12066 19768 12072 19780
rect 11164 19740 12072 19768
rect 7285 19731 7343 19737
rect 7300 19700 7328 19731
rect 12066 19728 12072 19740
rect 12124 19728 12130 19780
rect 13740 19768 13768 19876
rect 13909 19873 13921 19907
rect 13955 19904 13967 19907
rect 13955 19876 14688 19904
rect 13955 19873 13967 19876
rect 13909 19867 13967 19873
rect 14660 19848 14688 19876
rect 15654 19864 15660 19916
rect 15712 19864 15718 19916
rect 15746 19864 15752 19916
rect 15804 19904 15810 19916
rect 17328 19913 17356 19944
rect 17954 19932 17960 19944
rect 18012 19972 18018 19984
rect 19420 19975 19478 19981
rect 18012 19944 19012 19972
rect 18012 19932 18018 19944
rect 17586 19913 17592 19916
rect 16209 19907 16267 19913
rect 16209 19904 16221 19907
rect 15804 19876 16221 19904
rect 15804 19864 15810 19876
rect 16209 19873 16221 19876
rect 16255 19873 16267 19907
rect 16209 19867 16267 19873
rect 17313 19907 17371 19913
rect 17313 19873 17325 19907
rect 17359 19873 17371 19907
rect 17313 19867 17371 19873
rect 17580 19867 17592 19913
rect 17586 19864 17592 19867
rect 17644 19864 17650 19916
rect 18984 19848 19012 19944
rect 19420 19941 19432 19975
rect 19466 19972 19478 19975
rect 20990 19972 20996 19984
rect 19466 19944 20996 19972
rect 19466 19941 19478 19944
rect 19420 19935 19478 19941
rect 20990 19932 20996 19944
rect 21048 19932 21054 19984
rect 21284 19913 21312 20012
rect 21634 20000 21640 20012
rect 21692 20000 21698 20052
rect 21821 20043 21879 20049
rect 21821 20009 21833 20043
rect 21867 20040 21879 20043
rect 22554 20040 22560 20052
rect 21867 20012 22560 20040
rect 21867 20009 21879 20012
rect 21821 20003 21879 20009
rect 22554 20000 22560 20012
rect 22612 20000 22618 20052
rect 23198 20040 23204 20052
rect 22848 20012 23204 20040
rect 21453 19975 21511 19981
rect 21453 19941 21465 19975
rect 21499 19972 21511 19975
rect 21726 19972 21732 19984
rect 21499 19944 21732 19972
rect 21499 19941 21511 19944
rect 21453 19935 21511 19941
rect 21269 19907 21327 19913
rect 21269 19873 21281 19907
rect 21315 19873 21327 19907
rect 21269 19867 21327 19873
rect 14642 19796 14648 19848
rect 14700 19796 14706 19848
rect 16482 19836 16488 19848
rect 14752 19808 16488 19836
rect 14752 19768 14780 19808
rect 16482 19796 16488 19808
rect 16540 19796 16546 19848
rect 18966 19796 18972 19848
rect 19024 19836 19030 19848
rect 19153 19839 19211 19845
rect 19153 19836 19165 19839
rect 19024 19808 19165 19836
rect 19024 19796 19030 19808
rect 19153 19805 19165 19808
rect 19199 19805 19211 19839
rect 19153 19799 19211 19805
rect 13740 19740 14780 19768
rect 15381 19771 15439 19777
rect 15381 19737 15393 19771
rect 15427 19768 15439 19771
rect 20533 19771 20591 19777
rect 15427 19740 15884 19768
rect 15427 19737 15439 19740
rect 15381 19731 15439 19737
rect 15856 19712 15884 19740
rect 20533 19737 20545 19771
rect 20579 19768 20591 19771
rect 21468 19768 21496 19935
rect 21726 19932 21732 19944
rect 21784 19932 21790 19984
rect 22370 19972 22376 19984
rect 22296 19944 22376 19972
rect 21545 19907 21603 19913
rect 21545 19873 21557 19907
rect 21591 19873 21603 19907
rect 21545 19867 21603 19873
rect 21637 19907 21695 19913
rect 21637 19873 21649 19907
rect 21683 19904 21695 19907
rect 22094 19904 22100 19916
rect 21683 19876 22100 19904
rect 21683 19873 21695 19876
rect 21637 19867 21695 19873
rect 21560 19836 21588 19867
rect 22094 19864 22100 19876
rect 22152 19864 22158 19916
rect 22296 19913 22324 19944
rect 22370 19932 22376 19944
rect 22428 19972 22434 19984
rect 22428 19944 22600 19972
rect 22428 19932 22434 19944
rect 22281 19907 22339 19913
rect 22281 19873 22293 19907
rect 22327 19873 22339 19907
rect 22281 19867 22339 19873
rect 22465 19907 22523 19913
rect 22465 19873 22477 19907
rect 22511 19873 22523 19907
rect 22572 19904 22600 19944
rect 22646 19932 22652 19984
rect 22704 19981 22710 19984
rect 22704 19975 22767 19981
rect 22704 19941 22721 19975
rect 22755 19941 22767 19975
rect 22704 19935 22767 19941
rect 22704 19932 22710 19935
rect 22848 19904 22876 20012
rect 23198 20000 23204 20012
rect 23256 20000 23262 20052
rect 23569 20043 23627 20049
rect 23569 20009 23581 20043
rect 23615 20009 23627 20043
rect 23569 20003 23627 20009
rect 24121 20043 24179 20049
rect 24121 20009 24133 20043
rect 24167 20009 24179 20043
rect 24121 20003 24179 20009
rect 22925 19975 22983 19981
rect 22925 19941 22937 19975
rect 22971 19941 22983 19975
rect 22925 19935 22983 19941
rect 22572 19876 22876 19904
rect 22940 19904 22968 19935
rect 23382 19932 23388 19984
rect 23440 19932 23446 19984
rect 23584 19972 23612 20003
rect 24136 19972 24164 20003
rect 25326 19975 25384 19981
rect 25326 19972 25338 19975
rect 23584 19944 23980 19972
rect 24136 19944 25338 19972
rect 23952 19913 23980 19944
rect 25326 19941 25338 19944
rect 25372 19941 25384 19975
rect 25326 19935 25384 19941
rect 23845 19907 23903 19913
rect 23845 19904 23857 19907
rect 22940 19876 23857 19904
rect 22465 19867 22523 19873
rect 23845 19873 23857 19876
rect 23891 19873 23903 19907
rect 23845 19867 23903 19873
rect 23937 19907 23995 19913
rect 23937 19873 23949 19907
rect 23983 19873 23995 19907
rect 23937 19867 23995 19873
rect 22296 19836 22324 19867
rect 21560 19808 22324 19836
rect 22480 19836 22508 19867
rect 23566 19836 23572 19848
rect 22480 19808 23572 19836
rect 23566 19796 23572 19808
rect 23624 19796 23630 19848
rect 20579 19740 21496 19768
rect 22373 19771 22431 19777
rect 20579 19737 20591 19740
rect 20533 19731 20591 19737
rect 22373 19737 22385 19771
rect 22419 19768 22431 19771
rect 22419 19740 22968 19768
rect 22419 19737 22431 19740
rect 22373 19731 22431 19737
rect 5736 19672 7328 19700
rect 8386 19660 8392 19712
rect 8444 19660 8450 19712
rect 11698 19660 11704 19712
rect 11756 19660 11762 19712
rect 12434 19660 12440 19712
rect 12492 19700 12498 19712
rect 12529 19703 12587 19709
rect 12529 19700 12541 19703
rect 12492 19672 12541 19700
rect 12492 19660 12498 19672
rect 12529 19669 12541 19672
rect 12575 19669 12587 19703
rect 12529 19663 12587 19669
rect 12713 19703 12771 19709
rect 12713 19669 12725 19703
rect 12759 19700 12771 19703
rect 13170 19700 13176 19712
rect 12759 19672 13176 19700
rect 12759 19669 12771 19672
rect 12713 19663 12771 19669
rect 13170 19660 13176 19672
rect 13228 19660 13234 19712
rect 13814 19660 13820 19712
rect 13872 19660 13878 19712
rect 14001 19703 14059 19709
rect 14001 19669 14013 19703
rect 14047 19700 14059 19703
rect 14090 19700 14096 19712
rect 14047 19672 14096 19700
rect 14047 19669 14059 19672
rect 14001 19663 14059 19669
rect 14090 19660 14096 19672
rect 14148 19660 14154 19712
rect 15010 19660 15016 19712
rect 15068 19660 15074 19712
rect 15746 19660 15752 19712
rect 15804 19660 15810 19712
rect 15838 19660 15844 19712
rect 15896 19700 15902 19712
rect 15933 19703 15991 19709
rect 15933 19700 15945 19703
rect 15896 19672 15945 19700
rect 15896 19660 15902 19672
rect 15933 19669 15945 19672
rect 15979 19669 15991 19703
rect 15933 19663 15991 19669
rect 16850 19660 16856 19712
rect 16908 19660 16914 19712
rect 22557 19703 22615 19709
rect 22557 19669 22569 19703
rect 22603 19700 22615 19703
rect 22646 19700 22652 19712
rect 22603 19672 22652 19700
rect 22603 19669 22615 19672
rect 22557 19663 22615 19669
rect 22646 19660 22652 19672
rect 22704 19660 22710 19712
rect 22741 19703 22799 19709
rect 22741 19669 22753 19703
rect 22787 19700 22799 19703
rect 22830 19700 22836 19712
rect 22787 19672 22836 19700
rect 22787 19669 22799 19672
rect 22741 19663 22799 19669
rect 22830 19660 22836 19672
rect 22888 19660 22894 19712
rect 22940 19700 22968 19740
rect 23014 19728 23020 19780
rect 23072 19728 23078 19780
rect 23198 19728 23204 19780
rect 23256 19768 23262 19780
rect 23753 19771 23811 19777
rect 23753 19768 23765 19771
rect 23256 19740 23765 19768
rect 23256 19728 23262 19740
rect 23753 19737 23765 19740
rect 23799 19737 23811 19771
rect 23860 19768 23888 19867
rect 25593 19839 25651 19845
rect 25593 19805 25605 19839
rect 25639 19836 25651 19839
rect 27062 19836 27068 19848
rect 25639 19808 27068 19836
rect 25639 19805 25651 19808
rect 25593 19799 25651 19805
rect 27062 19796 27068 19808
rect 27120 19796 27126 19848
rect 24213 19771 24271 19777
rect 24213 19768 24225 19771
rect 23860 19740 24225 19768
rect 23753 19731 23811 19737
rect 24213 19737 24225 19740
rect 24259 19737 24271 19771
rect 24213 19731 24271 19737
rect 23385 19703 23443 19709
rect 23385 19700 23397 19703
rect 22940 19672 23397 19700
rect 23385 19669 23397 19672
rect 23431 19669 23443 19703
rect 23385 19663 23443 19669
rect 552 19610 27416 19632
rect 552 19558 3756 19610
rect 3808 19558 3820 19610
rect 3872 19558 3884 19610
rect 3936 19558 3948 19610
rect 4000 19558 4012 19610
rect 4064 19558 10472 19610
rect 10524 19558 10536 19610
rect 10588 19558 10600 19610
rect 10652 19558 10664 19610
rect 10716 19558 10728 19610
rect 10780 19558 17188 19610
rect 17240 19558 17252 19610
rect 17304 19558 17316 19610
rect 17368 19558 17380 19610
rect 17432 19558 17444 19610
rect 17496 19558 23904 19610
rect 23956 19558 23968 19610
rect 24020 19558 24032 19610
rect 24084 19558 24096 19610
rect 24148 19558 24160 19610
rect 24212 19558 27416 19610
rect 552 19536 27416 19558
rect 1029 19499 1087 19505
rect 1029 19465 1041 19499
rect 1075 19496 1087 19499
rect 1118 19496 1124 19508
rect 1075 19468 1124 19496
rect 1075 19465 1087 19468
rect 1029 19459 1087 19465
rect 1118 19456 1124 19468
rect 1176 19456 1182 19508
rect 1486 19456 1492 19508
rect 1544 19496 1550 19508
rect 2409 19499 2467 19505
rect 2409 19496 2421 19499
rect 1544 19468 2421 19496
rect 1544 19456 1550 19468
rect 2409 19465 2421 19468
rect 2455 19465 2467 19499
rect 2409 19459 2467 19465
rect 2593 19499 2651 19505
rect 2593 19465 2605 19499
rect 2639 19496 2651 19499
rect 2774 19496 2780 19508
rect 2639 19468 2780 19496
rect 2639 19465 2651 19468
rect 2593 19459 2651 19465
rect 2774 19456 2780 19468
rect 2832 19456 2838 19508
rect 2869 19499 2927 19505
rect 2869 19465 2881 19499
rect 2915 19496 2927 19499
rect 3326 19496 3332 19508
rect 2915 19468 3332 19496
rect 2915 19465 2927 19468
rect 2869 19459 2927 19465
rect 3326 19456 3332 19468
rect 3384 19456 3390 19508
rect 4246 19456 4252 19508
rect 4304 19456 4310 19508
rect 4430 19456 4436 19508
rect 4488 19456 4494 19508
rect 6730 19456 6736 19508
rect 6788 19456 6794 19508
rect 7469 19499 7527 19505
rect 7469 19465 7481 19499
rect 7515 19496 7527 19499
rect 7929 19499 7987 19505
rect 7929 19496 7941 19499
rect 7515 19468 7941 19496
rect 7515 19465 7527 19468
rect 7469 19459 7527 19465
rect 7929 19465 7941 19468
rect 7975 19496 7987 19499
rect 8110 19496 8116 19508
rect 7975 19468 8116 19496
rect 7975 19465 7987 19468
rect 7929 19459 7987 19465
rect 8110 19456 8116 19468
rect 8168 19496 8174 19508
rect 8757 19499 8815 19505
rect 8757 19496 8769 19499
rect 8168 19468 8769 19496
rect 8168 19456 8174 19468
rect 8757 19465 8769 19468
rect 8803 19465 8815 19499
rect 8757 19459 8815 19465
rect 12894 19456 12900 19508
rect 12952 19456 12958 19508
rect 13170 19456 13176 19508
rect 13228 19456 13234 19508
rect 13814 19456 13820 19508
rect 13872 19496 13878 19508
rect 15473 19499 15531 19505
rect 15473 19496 15485 19499
rect 13872 19468 15485 19496
rect 13872 19456 13878 19468
rect 15473 19465 15485 19468
rect 15519 19465 15531 19499
rect 15473 19459 15531 19465
rect 16206 19456 16212 19508
rect 16264 19456 16270 19508
rect 16945 19499 17003 19505
rect 16945 19465 16957 19499
rect 16991 19496 17003 19499
rect 17586 19496 17592 19508
rect 16991 19468 17592 19496
rect 16991 19465 17003 19468
rect 16945 19459 17003 19465
rect 17586 19456 17592 19468
rect 17644 19456 17650 19508
rect 20162 19456 20168 19508
rect 20220 19496 20226 19508
rect 20625 19499 20683 19505
rect 20625 19496 20637 19499
rect 20220 19468 20637 19496
rect 20220 19456 20226 19468
rect 20625 19465 20637 19468
rect 20671 19465 20683 19499
rect 20625 19459 20683 19465
rect 22646 19456 22652 19508
rect 22704 19496 22710 19508
rect 23014 19496 23020 19508
rect 22704 19468 23020 19496
rect 22704 19456 22710 19468
rect 23014 19456 23020 19468
rect 23072 19456 23078 19508
rect 2038 19388 2044 19440
rect 2096 19428 2102 19440
rect 2685 19431 2743 19437
rect 2685 19428 2697 19431
rect 2096 19400 2697 19428
rect 2096 19388 2102 19400
rect 2685 19397 2697 19400
rect 2731 19397 2743 19431
rect 5810 19428 5816 19440
rect 2685 19391 2743 19397
rect 5736 19400 5816 19428
rect 3329 19363 3387 19369
rect 3329 19360 3341 19363
rect 2746 19332 3341 19360
rect 1210 19252 1216 19304
rect 1268 19252 1274 19304
rect 1765 19295 1823 19301
rect 1765 19261 1777 19295
rect 1811 19292 1823 19295
rect 1854 19292 1860 19304
rect 1811 19264 1860 19292
rect 1811 19261 1823 19264
rect 1765 19255 1823 19261
rect 1854 19252 1860 19264
rect 1912 19252 1918 19304
rect 1949 19295 2007 19301
rect 1949 19261 1961 19295
rect 1995 19261 2007 19295
rect 2746 19292 2774 19332
rect 3329 19329 3341 19332
rect 3375 19360 3387 19363
rect 3602 19360 3608 19372
rect 3375 19332 3608 19360
rect 3375 19329 3387 19332
rect 3329 19323 3387 19329
rect 3602 19320 3608 19332
rect 3660 19320 3666 19372
rect 5626 19320 5632 19372
rect 5684 19320 5690 19372
rect 3421 19295 3479 19301
rect 3421 19292 3433 19295
rect 1949 19255 2007 19261
rect 2332 19264 2774 19292
rect 3068 19264 3433 19292
rect 1964 19224 1992 19255
rect 2332 19224 2360 19264
rect 1964 19196 2360 19224
rect 2498 19184 2504 19236
rect 2556 19224 2562 19236
rect 3068 19233 3096 19264
rect 3421 19261 3433 19264
rect 3467 19292 3479 19295
rect 3973 19295 4031 19301
rect 3973 19292 3985 19295
rect 3467 19264 3985 19292
rect 3467 19261 3479 19264
rect 3421 19255 3479 19261
rect 3973 19261 3985 19264
rect 4019 19261 4031 19295
rect 3973 19255 4031 19261
rect 4614 19252 4620 19304
rect 4672 19292 4678 19304
rect 4893 19295 4951 19301
rect 4893 19292 4905 19295
rect 4672 19264 4905 19292
rect 4672 19252 4678 19264
rect 4893 19261 4905 19264
rect 4939 19261 4951 19295
rect 4893 19255 4951 19261
rect 4985 19295 5043 19301
rect 4985 19261 4997 19295
rect 5031 19292 5043 19295
rect 5537 19295 5595 19301
rect 5031 19264 5488 19292
rect 5031 19261 5043 19264
rect 4985 19255 5043 19261
rect 5460 19233 5488 19264
rect 5537 19261 5549 19295
rect 5583 19292 5595 19295
rect 5736 19292 5764 19400
rect 5810 19388 5816 19400
rect 5868 19388 5874 19440
rect 7745 19431 7803 19437
rect 7745 19428 7757 19431
rect 7024 19400 7757 19428
rect 5583 19264 5764 19292
rect 5583 19261 5595 19264
rect 5537 19255 5595 19261
rect 5810 19252 5816 19304
rect 5868 19252 5874 19304
rect 5905 19295 5963 19301
rect 5905 19261 5917 19295
rect 5951 19261 5963 19295
rect 5905 19255 5963 19261
rect 6917 19295 6975 19301
rect 6917 19261 6929 19295
rect 6963 19292 6975 19295
rect 7024 19292 7052 19400
rect 7745 19397 7757 19400
rect 7791 19397 7803 19431
rect 7745 19391 7803 19397
rect 14642 19388 14648 19440
rect 14700 19428 14706 19440
rect 14921 19431 14979 19437
rect 14921 19428 14933 19431
rect 14700 19400 14933 19428
rect 14700 19388 14706 19400
rect 14921 19397 14933 19400
rect 14967 19397 14979 19431
rect 14921 19391 14979 19397
rect 17310 19388 17316 19440
rect 17368 19428 17374 19440
rect 17770 19428 17776 19440
rect 17368 19400 17776 19428
rect 17368 19388 17374 19400
rect 17770 19388 17776 19400
rect 17828 19388 17834 19440
rect 22094 19388 22100 19440
rect 22152 19428 22158 19440
rect 22152 19400 22508 19428
rect 22152 19388 22158 19400
rect 16393 19363 16451 19369
rect 7116 19332 7328 19360
rect 7116 19301 7144 19332
rect 6963 19264 7052 19292
rect 7101 19295 7159 19301
rect 6963 19261 6975 19264
rect 6917 19255 6975 19261
rect 7101 19261 7113 19295
rect 7147 19261 7159 19295
rect 7101 19255 7159 19261
rect 3053 19227 3111 19233
rect 3053 19224 3065 19227
rect 2556 19196 3065 19224
rect 2556 19184 2562 19196
rect 3053 19193 3065 19196
rect 3099 19193 3111 19227
rect 3053 19187 3111 19193
rect 5445 19227 5503 19233
rect 5445 19193 5457 19227
rect 5491 19193 5503 19227
rect 5445 19187 5503 19193
rect 5626 19184 5632 19236
rect 5684 19224 5690 19236
rect 5920 19224 5948 19255
rect 7190 19252 7196 19304
rect 7248 19252 7254 19304
rect 7300 19292 7328 19332
rect 16393 19329 16405 19363
rect 16439 19329 16451 19363
rect 17862 19360 17868 19372
rect 16393 19323 16451 19329
rect 17144 19332 17868 19360
rect 7742 19292 7748 19304
rect 7300 19264 7748 19292
rect 7742 19252 7748 19264
rect 7800 19252 7806 19304
rect 11514 19252 11520 19304
rect 11572 19252 11578 19304
rect 13354 19252 13360 19304
rect 13412 19292 13418 19304
rect 13541 19295 13599 19301
rect 13541 19292 13553 19295
rect 13412 19264 13553 19292
rect 13412 19252 13418 19264
rect 13541 19261 13553 19264
rect 13587 19261 13599 19295
rect 14090 19292 14096 19304
rect 13541 19255 13599 19261
rect 13648 19264 14096 19292
rect 7285 19227 7343 19233
rect 7285 19224 7297 19227
rect 5684 19196 5948 19224
rect 7116 19196 7297 19224
rect 5684 19184 5690 19196
rect 1949 19159 2007 19165
rect 1949 19125 1961 19159
rect 1995 19156 2007 19159
rect 2409 19159 2467 19165
rect 2409 19156 2421 19159
rect 1995 19128 2421 19156
rect 1995 19125 2007 19128
rect 1949 19119 2007 19125
rect 2409 19125 2421 19128
rect 2455 19125 2467 19159
rect 2409 19119 2467 19125
rect 2682 19116 2688 19168
rect 2740 19156 2746 19168
rect 2843 19159 2901 19165
rect 2843 19156 2855 19159
rect 2740 19128 2855 19156
rect 2740 19116 2746 19128
rect 2843 19125 2855 19128
rect 2889 19125 2901 19159
rect 2843 19119 2901 19125
rect 4614 19116 4620 19168
rect 4672 19156 4678 19168
rect 4709 19159 4767 19165
rect 4709 19156 4721 19159
rect 4672 19128 4721 19156
rect 4672 19116 4678 19128
rect 4709 19125 4721 19128
rect 4755 19125 4767 19159
rect 4709 19119 4767 19125
rect 5353 19159 5411 19165
rect 5353 19125 5365 19159
rect 5399 19156 5411 19159
rect 5902 19156 5908 19168
rect 5399 19128 5908 19156
rect 5399 19125 5411 19128
rect 5353 19119 5411 19125
rect 5902 19116 5908 19128
rect 5960 19116 5966 19168
rect 6454 19116 6460 19168
rect 6512 19156 6518 19168
rect 7116 19156 7144 19196
rect 7285 19193 7297 19196
rect 7331 19193 7343 19227
rect 7897 19227 7955 19233
rect 7897 19224 7909 19227
rect 7285 19187 7343 19193
rect 7500 19196 7909 19224
rect 7500 19168 7528 19196
rect 7897 19193 7909 19196
rect 7943 19224 7955 19227
rect 8113 19227 8171 19233
rect 7943 19193 7956 19224
rect 7897 19187 7956 19193
rect 8113 19193 8125 19227
rect 8159 19224 8171 19227
rect 8386 19224 8392 19236
rect 8159 19196 8392 19224
rect 8159 19193 8171 19196
rect 8113 19187 8171 19193
rect 6512 19128 7144 19156
rect 6512 19116 6518 19128
rect 7466 19116 7472 19168
rect 7524 19165 7530 19168
rect 7524 19159 7543 19165
rect 7531 19125 7543 19159
rect 7524 19119 7543 19125
rect 7524 19116 7530 19119
rect 7650 19116 7656 19168
rect 7708 19116 7714 19168
rect 7928 19156 7956 19187
rect 8386 19184 8392 19196
rect 8444 19184 8450 19236
rect 8570 19184 8576 19236
rect 8628 19184 8634 19236
rect 9490 19184 9496 19236
rect 9548 19224 9554 19236
rect 9766 19224 9772 19236
rect 9548 19196 9772 19224
rect 9548 19184 9554 19196
rect 9766 19184 9772 19196
rect 9824 19184 9830 19236
rect 11054 19184 11060 19236
rect 11112 19184 11118 19236
rect 11784 19227 11842 19233
rect 11784 19193 11796 19227
rect 11830 19224 11842 19227
rect 12250 19224 12256 19236
rect 11830 19196 12256 19224
rect 11830 19193 11842 19196
rect 11784 19187 11842 19193
rect 12250 19184 12256 19196
rect 12308 19184 12314 19236
rect 12989 19227 13047 19233
rect 12989 19193 13001 19227
rect 13035 19224 13047 19227
rect 13648 19224 13676 19264
rect 14090 19252 14096 19264
rect 14148 19252 14154 19304
rect 15194 19252 15200 19304
rect 15252 19252 15258 19304
rect 15286 19252 15292 19304
rect 15344 19252 15350 19304
rect 15565 19295 15623 19301
rect 15565 19261 15577 19295
rect 15611 19292 15623 19295
rect 15746 19292 15752 19304
rect 15611 19264 15752 19292
rect 15611 19261 15623 19264
rect 15565 19255 15623 19261
rect 15746 19252 15752 19264
rect 15804 19252 15810 19304
rect 15838 19252 15844 19304
rect 15896 19252 15902 19304
rect 16025 19295 16083 19301
rect 16025 19261 16037 19295
rect 16071 19292 16083 19295
rect 16114 19292 16120 19304
rect 16071 19264 16120 19292
rect 16071 19261 16083 19264
rect 16025 19255 16083 19261
rect 16114 19252 16120 19264
rect 16172 19252 16178 19304
rect 13035 19196 13676 19224
rect 13786 19227 13844 19233
rect 13035 19193 13047 19196
rect 12989 19187 13047 19193
rect 13786 19193 13798 19227
rect 13832 19224 13844 19227
rect 13832 19193 13860 19224
rect 13786 19187 13860 19193
rect 8754 19156 8760 19168
rect 8812 19165 8818 19168
rect 8812 19159 8831 19165
rect 7928 19128 8760 19156
rect 8754 19116 8760 19128
rect 8819 19125 8831 19159
rect 8812 19119 8831 19125
rect 8812 19116 8818 19119
rect 8938 19116 8944 19168
rect 8996 19116 9002 19168
rect 12802 19116 12808 19168
rect 12860 19156 12866 19168
rect 13189 19159 13247 19165
rect 13189 19156 13201 19159
rect 12860 19128 13201 19156
rect 12860 19116 12866 19128
rect 13189 19125 13201 19128
rect 13235 19125 13247 19159
rect 13189 19119 13247 19125
rect 13354 19116 13360 19168
rect 13412 19116 13418 19168
rect 13538 19116 13544 19168
rect 13596 19156 13602 19168
rect 13832 19156 13860 19187
rect 15470 19184 15476 19236
rect 15528 19224 15534 19236
rect 16408 19224 16436 19323
rect 16485 19295 16543 19301
rect 16485 19261 16497 19295
rect 16531 19292 16543 19295
rect 16850 19292 16856 19304
rect 16531 19264 16856 19292
rect 16531 19261 16543 19264
rect 16485 19255 16543 19261
rect 16850 19252 16856 19264
rect 16908 19252 16914 19304
rect 17144 19301 17172 19332
rect 17862 19320 17868 19332
rect 17920 19320 17926 19372
rect 22189 19363 22247 19369
rect 22189 19360 22201 19363
rect 22020 19332 22201 19360
rect 17129 19295 17187 19301
rect 17129 19261 17141 19295
rect 17175 19261 17187 19295
rect 17129 19255 17187 19261
rect 17310 19252 17316 19304
rect 17368 19252 17374 19304
rect 17497 19295 17555 19301
rect 17497 19261 17509 19295
rect 17543 19292 17555 19295
rect 18046 19292 18052 19304
rect 17543 19264 18052 19292
rect 17543 19261 17555 19264
rect 17497 19255 17555 19261
rect 18046 19252 18052 19264
rect 18104 19252 18110 19304
rect 18417 19295 18475 19301
rect 18417 19261 18429 19295
rect 18463 19292 18475 19295
rect 18966 19292 18972 19304
rect 18463 19264 18972 19292
rect 18463 19261 18475 19264
rect 18417 19255 18475 19261
rect 18966 19252 18972 19264
rect 19024 19292 19030 19304
rect 19153 19295 19211 19301
rect 19153 19292 19165 19295
rect 19024 19264 19165 19292
rect 19024 19252 19030 19264
rect 19153 19261 19165 19264
rect 19199 19261 19211 19295
rect 19153 19255 19211 19261
rect 21174 19252 21180 19304
rect 21232 19252 21238 19304
rect 21361 19295 21419 19301
rect 21361 19261 21373 19295
rect 21407 19292 21419 19295
rect 22020 19292 22048 19332
rect 22189 19329 22201 19332
rect 22235 19360 22247 19363
rect 22278 19360 22284 19372
rect 22235 19332 22284 19360
rect 22235 19329 22247 19332
rect 22189 19323 22247 19329
rect 22278 19320 22284 19332
rect 22336 19320 22342 19372
rect 21407 19264 22048 19292
rect 22097 19295 22155 19301
rect 21407 19261 21419 19264
rect 21361 19255 21419 19261
rect 22097 19261 22109 19295
rect 22143 19261 22155 19295
rect 22097 19255 22155 19261
rect 15528 19196 16436 19224
rect 15528 19184 15534 19196
rect 17218 19184 17224 19236
rect 17276 19184 17282 19236
rect 17586 19184 17592 19236
rect 17644 19184 17650 19236
rect 18506 19184 18512 19236
rect 18564 19224 18570 19236
rect 19058 19224 19064 19236
rect 18564 19196 19064 19224
rect 18564 19184 18570 19196
rect 19058 19184 19064 19196
rect 19116 19184 19122 19236
rect 19420 19227 19478 19233
rect 19420 19193 19432 19227
rect 19466 19224 19478 19227
rect 21082 19224 21088 19236
rect 19466 19196 21088 19224
rect 19466 19193 19478 19196
rect 19420 19187 19478 19193
rect 21082 19184 21088 19196
rect 21140 19184 21146 19236
rect 13596 19128 13860 19156
rect 13596 19116 13602 19128
rect 15010 19116 15016 19168
rect 15068 19116 15074 19168
rect 15657 19159 15715 19165
rect 15657 19125 15669 19159
rect 15703 19156 15715 19159
rect 15746 19156 15752 19168
rect 15703 19128 15752 19156
rect 15703 19125 15715 19128
rect 15657 19119 15715 19125
rect 15746 19116 15752 19128
rect 15804 19116 15810 19168
rect 17604 19156 17632 19184
rect 20438 19156 20444 19168
rect 17604 19128 20444 19156
rect 20438 19116 20444 19128
rect 20496 19116 20502 19168
rect 20533 19159 20591 19165
rect 20533 19125 20545 19159
rect 20579 19156 20591 19159
rect 21376 19156 21404 19255
rect 20579 19128 21404 19156
rect 20579 19125 20591 19128
rect 20533 19119 20591 19125
rect 21818 19116 21824 19168
rect 21876 19156 21882 19168
rect 22005 19159 22063 19165
rect 22005 19156 22017 19159
rect 21876 19128 22017 19156
rect 21876 19116 21882 19128
rect 22005 19125 22017 19128
rect 22051 19125 22063 19159
rect 22112 19156 22140 19255
rect 22370 19252 22376 19304
rect 22428 19252 22434 19304
rect 22480 19301 22508 19400
rect 22830 19320 22836 19372
rect 22888 19360 22894 19372
rect 22888 19332 23152 19360
rect 22888 19320 22894 19332
rect 22465 19295 22523 19301
rect 22465 19261 22477 19295
rect 22511 19261 22523 19295
rect 22465 19255 22523 19261
rect 22738 19252 22744 19304
rect 22796 19252 22802 19304
rect 23014 19252 23020 19304
rect 23072 19252 23078 19304
rect 23124 19292 23152 19332
rect 23290 19292 23296 19304
rect 23124 19264 23296 19292
rect 23290 19252 23296 19264
rect 23348 19292 23354 19304
rect 23569 19295 23627 19301
rect 23569 19292 23581 19295
rect 23348 19264 23581 19292
rect 23348 19252 23354 19264
rect 23569 19261 23581 19264
rect 23615 19292 23627 19295
rect 25130 19292 25136 19304
rect 23615 19264 25136 19292
rect 23615 19261 23627 19264
rect 23569 19255 23627 19261
rect 25130 19252 25136 19264
rect 25188 19252 25194 19304
rect 26973 19295 27031 19301
rect 26973 19261 26985 19295
rect 27019 19292 27031 19295
rect 27062 19292 27068 19304
rect 27019 19264 27068 19292
rect 27019 19261 27031 19264
rect 26973 19255 27031 19261
rect 27062 19252 27068 19264
rect 27120 19252 27126 19304
rect 22922 19184 22928 19236
rect 22980 19224 22986 19236
rect 23382 19224 23388 19236
rect 22980 19196 23388 19224
rect 22980 19184 22986 19196
rect 23382 19184 23388 19196
rect 23440 19184 23446 19236
rect 25774 19184 25780 19236
rect 25832 19224 25838 19236
rect 26706 19227 26764 19233
rect 26706 19224 26718 19227
rect 25832 19196 26718 19224
rect 25832 19184 25838 19196
rect 26706 19193 26718 19196
rect 26752 19193 26764 19227
rect 26706 19187 26764 19193
rect 22462 19156 22468 19168
rect 22112 19128 22468 19156
rect 22005 19119 22063 19125
rect 22462 19116 22468 19128
rect 22520 19116 22526 19168
rect 22649 19159 22707 19165
rect 22649 19125 22661 19159
rect 22695 19156 22707 19159
rect 22833 19159 22891 19165
rect 22833 19156 22845 19159
rect 22695 19128 22845 19156
rect 22695 19125 22707 19128
rect 22649 19119 22707 19125
rect 22833 19125 22845 19128
rect 22879 19125 22891 19159
rect 22833 19119 22891 19125
rect 23201 19159 23259 19165
rect 23201 19125 23213 19159
rect 23247 19156 23259 19159
rect 23290 19156 23296 19168
rect 23247 19128 23296 19156
rect 23247 19125 23259 19128
rect 23201 19119 23259 19125
rect 23290 19116 23296 19128
rect 23348 19116 23354 19168
rect 24762 19116 24768 19168
rect 24820 19156 24826 19168
rect 25593 19159 25651 19165
rect 25593 19156 25605 19159
rect 24820 19128 25605 19156
rect 24820 19116 24826 19128
rect 25593 19125 25605 19128
rect 25639 19125 25651 19159
rect 25593 19119 25651 19125
rect 552 19066 27576 19088
rect 552 19014 7114 19066
rect 7166 19014 7178 19066
rect 7230 19014 7242 19066
rect 7294 19014 7306 19066
rect 7358 19014 7370 19066
rect 7422 19014 13830 19066
rect 13882 19014 13894 19066
rect 13946 19014 13958 19066
rect 14010 19014 14022 19066
rect 14074 19014 14086 19066
rect 14138 19014 20546 19066
rect 20598 19014 20610 19066
rect 20662 19014 20674 19066
rect 20726 19014 20738 19066
rect 20790 19014 20802 19066
rect 20854 19014 27262 19066
rect 27314 19014 27326 19066
rect 27378 19014 27390 19066
rect 27442 19014 27454 19066
rect 27506 19014 27518 19066
rect 27570 19014 27576 19066
rect 552 18992 27576 19014
rect 2498 18912 2504 18964
rect 2556 18912 2562 18964
rect 5810 18912 5816 18964
rect 5868 18952 5874 18964
rect 6089 18955 6147 18961
rect 6089 18952 6101 18955
rect 5868 18924 6101 18952
rect 5868 18912 5874 18924
rect 6089 18921 6101 18924
rect 6135 18921 6147 18955
rect 6089 18915 6147 18921
rect 6362 18912 6368 18964
rect 6420 18952 6426 18964
rect 7929 18955 7987 18961
rect 7929 18952 7941 18955
rect 6420 18924 7941 18952
rect 6420 18912 6426 18924
rect 7929 18921 7941 18924
rect 7975 18952 7987 18955
rect 8570 18952 8576 18964
rect 7975 18924 8576 18952
rect 7975 18921 7987 18924
rect 7929 18915 7987 18921
rect 8570 18912 8576 18924
rect 8628 18912 8634 18964
rect 11054 18912 11060 18964
rect 11112 18952 11118 18964
rect 14369 18955 14427 18961
rect 14369 18952 14381 18955
rect 11112 18924 14381 18952
rect 11112 18912 11118 18924
rect 14369 18921 14381 18924
rect 14415 18952 14427 18955
rect 14415 18924 19288 18952
rect 14415 18921 14427 18924
rect 14369 18915 14427 18921
rect 2958 18844 2964 18896
rect 3016 18884 3022 18896
rect 3614 18887 3672 18893
rect 3614 18884 3626 18887
rect 3016 18856 3626 18884
rect 3016 18844 3022 18856
rect 3614 18853 3626 18856
rect 3660 18853 3672 18887
rect 6546 18884 6552 18896
rect 3614 18847 3672 18853
rect 5828 18856 6552 18884
rect 3881 18819 3939 18825
rect 3881 18785 3893 18819
rect 3927 18816 3939 18819
rect 5718 18816 5724 18828
rect 3927 18788 5724 18816
rect 3927 18785 3939 18788
rect 3881 18779 3939 18785
rect 5718 18776 5724 18788
rect 5776 18776 5782 18828
rect 5828 18825 5856 18856
rect 6546 18844 6552 18856
rect 6604 18844 6610 18896
rect 11514 18884 11520 18896
rect 7852 18856 11520 18884
rect 5813 18819 5871 18825
rect 5813 18785 5825 18819
rect 5859 18785 5871 18819
rect 5813 18779 5871 18785
rect 5994 18776 6000 18828
rect 6052 18776 6058 18828
rect 6086 18776 6092 18828
rect 6144 18776 6150 18828
rect 6273 18819 6331 18825
rect 6273 18785 6285 18819
rect 6319 18785 6331 18819
rect 6273 18779 6331 18785
rect 6288 18748 6316 18779
rect 7282 18776 7288 18828
rect 7340 18816 7346 18828
rect 7852 18825 7880 18856
rect 7570 18819 7628 18825
rect 7570 18816 7582 18819
rect 7340 18788 7582 18816
rect 7340 18776 7346 18788
rect 7570 18785 7582 18788
rect 7616 18785 7628 18819
rect 7570 18779 7628 18785
rect 7837 18819 7895 18825
rect 7837 18785 7849 18819
rect 7883 18785 7895 18819
rect 7837 18779 7895 18785
rect 8570 18776 8576 18828
rect 8628 18816 8634 18828
rect 9042 18819 9100 18825
rect 9042 18816 9054 18819
rect 8628 18788 9054 18816
rect 8628 18776 8634 18788
rect 9042 18785 9054 18788
rect 9088 18785 9100 18819
rect 9042 18779 9100 18785
rect 9324 18757 9352 18856
rect 10796 18825 10824 18856
rect 11514 18844 11520 18856
rect 11572 18844 11578 18896
rect 12250 18844 12256 18896
rect 12308 18844 12314 18896
rect 13173 18887 13231 18893
rect 13173 18853 13185 18887
rect 13219 18884 13231 18887
rect 13446 18884 13452 18896
rect 13219 18856 13452 18884
rect 13219 18853 13231 18856
rect 13173 18847 13231 18853
rect 13446 18844 13452 18856
rect 13504 18844 13510 18896
rect 13538 18844 13544 18896
rect 13596 18844 13602 18896
rect 13725 18887 13783 18893
rect 13725 18853 13737 18887
rect 13771 18884 13783 18887
rect 15194 18884 15200 18896
rect 13771 18856 15200 18884
rect 13771 18853 13783 18856
rect 13725 18847 13783 18853
rect 14384 18828 14412 18856
rect 15194 18844 15200 18856
rect 15252 18844 15258 18896
rect 19260 18893 19288 18924
rect 20438 18912 20444 18964
rect 20496 18952 20502 18964
rect 20533 18955 20591 18961
rect 20533 18952 20545 18955
rect 20496 18924 20545 18952
rect 20496 18912 20502 18924
rect 20533 18921 20545 18924
rect 20579 18952 20591 18955
rect 21266 18952 21272 18964
rect 20579 18924 21272 18952
rect 20579 18921 20591 18924
rect 20533 18915 20591 18921
rect 21266 18912 21272 18924
rect 21324 18912 21330 18964
rect 21358 18912 21364 18964
rect 21416 18952 21422 18964
rect 21913 18955 21971 18961
rect 21416 18924 21588 18952
rect 21416 18912 21422 18924
rect 21560 18893 21588 18924
rect 21913 18921 21925 18955
rect 21959 18952 21971 18955
rect 23014 18952 23020 18964
rect 21959 18924 23020 18952
rect 21959 18921 21971 18924
rect 21913 18915 21971 18921
rect 23014 18912 23020 18924
rect 23072 18912 23078 18964
rect 25774 18912 25780 18964
rect 25832 18912 25838 18964
rect 15657 18887 15715 18893
rect 15657 18853 15669 18887
rect 15703 18884 15715 18887
rect 19245 18887 19303 18893
rect 15703 18856 18920 18884
rect 15703 18853 15715 18856
rect 15657 18847 15715 18853
rect 10525 18819 10583 18825
rect 10525 18785 10537 18819
rect 10571 18816 10583 18819
rect 10781 18819 10839 18825
rect 10571 18788 10732 18816
rect 10571 18785 10583 18788
rect 10525 18779 10583 18785
rect 5920 18720 6316 18748
rect 9309 18751 9367 18757
rect 4982 18572 4988 18624
rect 5040 18612 5046 18624
rect 5920 18621 5948 18720
rect 9309 18717 9321 18751
rect 9355 18748 9367 18751
rect 9582 18748 9588 18760
rect 9355 18720 9588 18748
rect 9355 18717 9367 18720
rect 9309 18711 9367 18717
rect 9582 18708 9588 18720
rect 9640 18708 9646 18760
rect 10704 18748 10732 18788
rect 10781 18785 10793 18819
rect 10827 18785 10839 18819
rect 10781 18779 10839 18785
rect 11241 18819 11299 18825
rect 11241 18785 11253 18819
rect 11287 18785 11299 18819
rect 11241 18779 11299 18785
rect 10704 18720 10824 18748
rect 6454 18640 6460 18692
rect 6512 18640 6518 18692
rect 10796 18680 10824 18720
rect 11054 18708 11060 18760
rect 11112 18708 11118 18760
rect 11256 18748 11284 18779
rect 11422 18776 11428 18828
rect 11480 18776 11486 18828
rect 11698 18776 11704 18828
rect 11756 18776 11762 18828
rect 12434 18776 12440 18828
rect 12492 18776 12498 18828
rect 12618 18776 12624 18828
rect 12676 18776 12682 18828
rect 12713 18819 12771 18825
rect 12713 18785 12725 18819
rect 12759 18816 12771 18819
rect 13078 18816 13084 18828
rect 12759 18788 13084 18816
rect 12759 18785 12771 18788
rect 12713 18779 12771 18785
rect 13078 18776 13084 18788
rect 13136 18776 13142 18828
rect 13354 18776 13360 18828
rect 13412 18776 13418 18828
rect 13630 18776 13636 18828
rect 13688 18776 13694 18828
rect 14366 18776 14372 18828
rect 14424 18776 14430 18828
rect 16666 18776 16672 18828
rect 16724 18816 16730 18828
rect 17230 18819 17288 18825
rect 17230 18816 17242 18819
rect 16724 18788 17242 18816
rect 16724 18776 16730 18788
rect 17230 18785 17242 18788
rect 17276 18785 17288 18819
rect 17230 18779 17288 18785
rect 17678 18776 17684 18828
rect 17736 18816 17742 18828
rect 17845 18819 17903 18825
rect 17845 18816 17857 18819
rect 17736 18788 17857 18816
rect 17736 18776 17742 18788
rect 17845 18785 17857 18788
rect 17891 18785 17903 18819
rect 17845 18779 17903 18785
rect 12636 18748 12664 18776
rect 17497 18751 17555 18757
rect 11256 18720 11652 18748
rect 12636 18720 16068 18748
rect 11624 18692 11652 18720
rect 11517 18683 11575 18689
rect 11517 18680 11529 18683
rect 10796 18652 11529 18680
rect 11517 18649 11529 18652
rect 11563 18649 11575 18683
rect 11517 18643 11575 18649
rect 11606 18640 11612 18692
rect 11664 18680 11670 18692
rect 15930 18680 15936 18692
rect 11664 18652 15936 18680
rect 11664 18640 11670 18652
rect 15930 18640 15936 18652
rect 15988 18640 15994 18692
rect 5905 18615 5963 18621
rect 5905 18612 5917 18615
rect 5040 18584 5917 18612
rect 5040 18572 5046 18584
rect 5905 18581 5917 18584
rect 5951 18581 5963 18615
rect 5905 18575 5963 18581
rect 8386 18572 8392 18624
rect 8444 18612 8450 18624
rect 9401 18615 9459 18621
rect 9401 18612 9413 18615
rect 8444 18584 9413 18612
rect 8444 18572 8450 18584
rect 9401 18581 9413 18584
rect 9447 18612 9459 18615
rect 11054 18612 11060 18624
rect 9447 18584 11060 18612
rect 9447 18581 9459 18584
rect 9401 18575 9459 18581
rect 11054 18572 11060 18584
rect 11112 18572 11118 18624
rect 16040 18612 16068 18720
rect 17497 18717 17509 18751
rect 17543 18748 17555 18751
rect 17589 18751 17647 18757
rect 17589 18748 17601 18751
rect 17543 18720 17601 18748
rect 17543 18717 17555 18720
rect 17497 18711 17555 18717
rect 17589 18717 17601 18720
rect 17635 18717 17647 18751
rect 17589 18711 17647 18717
rect 16114 18640 16120 18692
rect 16172 18640 16178 18692
rect 17494 18612 17500 18624
rect 16040 18584 17500 18612
rect 17494 18572 17500 18584
rect 17552 18572 17558 18624
rect 17604 18612 17632 18711
rect 18892 18680 18920 18856
rect 19245 18853 19257 18887
rect 19291 18853 19303 18887
rect 19245 18847 19303 18853
rect 21545 18887 21603 18893
rect 21545 18853 21557 18887
rect 21591 18853 21603 18887
rect 21545 18847 21603 18853
rect 21726 18844 21732 18896
rect 21784 18884 21790 18896
rect 21784 18856 22232 18884
rect 21784 18844 21790 18856
rect 19058 18776 19064 18828
rect 19116 18816 19122 18828
rect 21358 18816 21364 18828
rect 19116 18788 21364 18816
rect 19116 18776 19122 18788
rect 21358 18776 21364 18788
rect 21416 18776 21422 18828
rect 21450 18776 21456 18828
rect 21508 18776 21514 18828
rect 21634 18776 21640 18828
rect 21692 18776 21698 18828
rect 21818 18776 21824 18828
rect 21876 18776 21882 18828
rect 22204 18825 22232 18856
rect 22278 18844 22284 18896
rect 22336 18844 22342 18896
rect 22388 18856 22876 18884
rect 22097 18819 22155 18825
rect 22097 18785 22109 18819
rect 22143 18785 22155 18819
rect 22097 18779 22155 18785
rect 22189 18819 22247 18825
rect 22189 18785 22201 18819
rect 22235 18816 22247 18819
rect 22388 18816 22416 18856
rect 22235 18788 22416 18816
rect 22235 18785 22247 18788
rect 22189 18779 22247 18785
rect 20898 18708 20904 18760
rect 20956 18748 20962 18760
rect 22112 18748 22140 18779
rect 22462 18776 22468 18828
rect 22520 18816 22526 18828
rect 22520 18788 22692 18816
rect 22520 18776 22526 18788
rect 20956 18720 22140 18748
rect 20956 18708 20962 18720
rect 22554 18708 22560 18760
rect 22612 18708 22618 18760
rect 22664 18748 22692 18788
rect 22738 18776 22744 18828
rect 22796 18776 22802 18828
rect 22848 18816 22876 18856
rect 22922 18844 22928 18896
rect 22980 18844 22986 18896
rect 23382 18884 23388 18896
rect 23032 18856 23388 18884
rect 23032 18816 23060 18856
rect 23382 18844 23388 18856
rect 23440 18844 23446 18896
rect 22848 18788 23060 18816
rect 23198 18776 23204 18828
rect 23256 18776 23262 18828
rect 25498 18776 25504 18828
rect 25556 18816 25562 18828
rect 25593 18819 25651 18825
rect 25593 18816 25605 18819
rect 25556 18788 25605 18816
rect 25556 18776 25562 18788
rect 25593 18785 25605 18788
rect 25639 18785 25651 18819
rect 25593 18779 25651 18785
rect 23109 18751 23167 18757
rect 23109 18748 23121 18751
rect 22664 18720 23121 18748
rect 23109 18717 23121 18720
rect 23155 18717 23167 18751
rect 23109 18711 23167 18717
rect 24946 18680 24952 18692
rect 18892 18652 24952 18680
rect 24946 18640 24952 18652
rect 25004 18640 25010 18692
rect 18874 18612 18880 18624
rect 17604 18584 18880 18612
rect 18874 18572 18880 18584
rect 18932 18572 18938 18624
rect 18969 18615 19027 18621
rect 18969 18581 18981 18615
rect 19015 18612 19027 18615
rect 19150 18612 19156 18624
rect 19015 18584 19156 18612
rect 19015 18581 19027 18584
rect 18969 18575 19027 18581
rect 19150 18572 19156 18584
rect 19208 18612 19214 18624
rect 20898 18612 20904 18624
rect 19208 18584 20904 18612
rect 19208 18572 19214 18584
rect 20898 18572 20904 18584
rect 20956 18572 20962 18624
rect 21082 18572 21088 18624
rect 21140 18612 21146 18624
rect 21269 18615 21327 18621
rect 21269 18612 21281 18615
rect 21140 18584 21281 18612
rect 21140 18572 21146 18584
rect 21269 18581 21281 18584
rect 21315 18581 21327 18615
rect 21269 18575 21327 18581
rect 22462 18572 22468 18624
rect 22520 18612 22526 18624
rect 22830 18612 22836 18624
rect 22520 18584 22836 18612
rect 22520 18572 22526 18584
rect 22830 18572 22836 18584
rect 22888 18572 22894 18624
rect 552 18522 27416 18544
rect 552 18470 3756 18522
rect 3808 18470 3820 18522
rect 3872 18470 3884 18522
rect 3936 18470 3948 18522
rect 4000 18470 4012 18522
rect 4064 18470 10472 18522
rect 10524 18470 10536 18522
rect 10588 18470 10600 18522
rect 10652 18470 10664 18522
rect 10716 18470 10728 18522
rect 10780 18470 17188 18522
rect 17240 18470 17252 18522
rect 17304 18470 17316 18522
rect 17368 18470 17380 18522
rect 17432 18470 17444 18522
rect 17496 18470 23904 18522
rect 23956 18470 23968 18522
rect 24020 18470 24032 18522
rect 24084 18470 24096 18522
rect 24148 18470 24160 18522
rect 24212 18470 27416 18522
rect 552 18448 27416 18470
rect 5074 18368 5080 18420
rect 5132 18408 5138 18420
rect 5261 18411 5319 18417
rect 5261 18408 5273 18411
rect 5132 18380 5273 18408
rect 5132 18368 5138 18380
rect 5261 18377 5273 18380
rect 5307 18377 5319 18411
rect 5261 18371 5319 18377
rect 6086 18368 6092 18420
rect 6144 18368 6150 18420
rect 7282 18368 7288 18420
rect 7340 18368 7346 18420
rect 8570 18368 8576 18420
rect 8628 18368 8634 18420
rect 13170 18368 13176 18420
rect 13228 18408 13234 18420
rect 13817 18411 13875 18417
rect 13817 18408 13829 18411
rect 13228 18380 13829 18408
rect 13228 18368 13234 18380
rect 13817 18377 13829 18380
rect 13863 18377 13875 18411
rect 13817 18371 13875 18377
rect 15749 18411 15807 18417
rect 15749 18377 15761 18411
rect 15795 18408 15807 18411
rect 16393 18411 16451 18417
rect 16393 18408 16405 18411
rect 15795 18380 16405 18408
rect 15795 18377 15807 18380
rect 15749 18371 15807 18377
rect 16393 18377 16405 18380
rect 16439 18377 16451 18411
rect 16393 18371 16451 18377
rect 16666 18368 16672 18420
rect 16724 18368 16730 18420
rect 17405 18411 17463 18417
rect 17405 18377 17417 18411
rect 17451 18408 17463 18411
rect 17678 18408 17684 18420
rect 17451 18380 17684 18408
rect 17451 18377 17463 18380
rect 17405 18371 17463 18377
rect 17678 18368 17684 18380
rect 17736 18368 17742 18420
rect 18417 18411 18475 18417
rect 18417 18377 18429 18411
rect 18463 18408 18475 18411
rect 18598 18408 18604 18420
rect 18463 18380 18604 18408
rect 18463 18377 18475 18380
rect 18417 18371 18475 18377
rect 18598 18368 18604 18380
rect 18656 18368 18662 18420
rect 20349 18411 20407 18417
rect 20349 18377 20361 18411
rect 20395 18408 20407 18411
rect 21174 18408 21180 18420
rect 20395 18380 21180 18408
rect 20395 18377 20407 18380
rect 20349 18371 20407 18377
rect 21174 18368 21180 18380
rect 21232 18408 21238 18420
rect 21542 18408 21548 18420
rect 21232 18380 21548 18408
rect 21232 18368 21238 18380
rect 21542 18368 21548 18380
rect 21600 18368 21606 18420
rect 21652 18380 22094 18408
rect 6454 18300 6460 18352
rect 6512 18300 6518 18352
rect 15933 18343 15991 18349
rect 12176 18312 15884 18340
rect 4617 18275 4675 18281
rect 4617 18241 4629 18275
rect 4663 18272 4675 18275
rect 5258 18272 5264 18284
rect 4663 18244 5264 18272
rect 4663 18241 4675 18244
rect 4617 18235 4675 18241
rect 5258 18232 5264 18244
rect 5316 18232 5322 18284
rect 5626 18232 5632 18284
rect 5684 18272 5690 18284
rect 6472 18272 6500 18300
rect 5684 18244 6500 18272
rect 5684 18232 5690 18244
rect 1302 18164 1308 18216
rect 1360 18164 1366 18216
rect 2038 18164 2044 18216
rect 2096 18164 2102 18216
rect 2222 18164 2228 18216
rect 2280 18204 2286 18216
rect 2501 18207 2559 18213
rect 2501 18204 2513 18207
rect 2280 18176 2513 18204
rect 2280 18164 2286 18176
rect 2501 18173 2513 18176
rect 2547 18173 2559 18207
rect 2501 18167 2559 18173
rect 4522 18164 4528 18216
rect 4580 18164 4586 18216
rect 4982 18164 4988 18216
rect 5040 18164 5046 18216
rect 5445 18207 5503 18213
rect 5445 18173 5457 18207
rect 5491 18173 5503 18207
rect 5445 18167 5503 18173
rect 2056 18136 2084 18164
rect 2682 18136 2688 18148
rect 2056 18108 2688 18136
rect 2682 18096 2688 18108
rect 2740 18096 2746 18148
rect 4798 18096 4804 18148
rect 4856 18136 4862 18148
rect 5460 18136 5488 18167
rect 5534 18164 5540 18216
rect 5592 18204 5598 18216
rect 5736 18213 5764 18244
rect 6546 18232 6552 18284
rect 6604 18232 6610 18284
rect 7558 18232 7564 18284
rect 7616 18272 7622 18284
rect 12176 18281 12204 18312
rect 12161 18275 12219 18281
rect 7616 18244 9076 18272
rect 7616 18232 7622 18244
rect 5721 18207 5779 18213
rect 5592 18176 5637 18204
rect 5592 18164 5598 18176
rect 5721 18173 5733 18207
rect 5767 18173 5779 18207
rect 5721 18167 5779 18173
rect 5951 18207 6009 18213
rect 5951 18173 5963 18207
rect 5997 18204 6009 18207
rect 6362 18204 6368 18216
rect 5997 18176 6368 18204
rect 5997 18173 6009 18176
rect 5951 18167 6009 18173
rect 6362 18164 6368 18176
rect 6420 18164 6426 18216
rect 6457 18207 6515 18213
rect 6457 18173 6469 18207
rect 6503 18204 6515 18207
rect 6564 18204 6592 18232
rect 6503 18176 6592 18204
rect 7469 18207 7527 18213
rect 6503 18173 6515 18176
rect 6457 18167 6515 18173
rect 7469 18173 7481 18207
rect 7515 18204 7527 18207
rect 7650 18204 7656 18216
rect 7515 18176 7656 18204
rect 7515 18173 7527 18176
rect 7469 18167 7527 18173
rect 7650 18164 7656 18176
rect 7708 18164 7714 18216
rect 7760 18213 7788 18244
rect 7745 18207 7803 18213
rect 7745 18173 7757 18207
rect 7791 18173 7803 18207
rect 7745 18167 7803 18173
rect 8757 18207 8815 18213
rect 8757 18173 8769 18207
rect 8803 18204 8815 18207
rect 8938 18204 8944 18216
rect 8803 18176 8944 18204
rect 8803 18173 8815 18176
rect 8757 18167 8815 18173
rect 8938 18164 8944 18176
rect 8996 18164 9002 18216
rect 9048 18213 9076 18244
rect 12161 18241 12173 18275
rect 12207 18241 12219 18275
rect 12161 18235 12219 18241
rect 12253 18275 12311 18281
rect 12253 18241 12265 18275
rect 12299 18241 12311 18275
rect 12253 18235 12311 18241
rect 13265 18275 13323 18281
rect 13265 18241 13277 18275
rect 13311 18272 13323 18275
rect 15381 18275 15439 18281
rect 13311 18244 14596 18272
rect 13311 18241 13323 18244
rect 13265 18235 13323 18241
rect 9033 18207 9091 18213
rect 9033 18173 9045 18207
rect 9079 18173 9091 18207
rect 10229 18207 10287 18213
rect 10229 18204 10241 18207
rect 9033 18167 9091 18173
rect 9968 18176 10241 18204
rect 4856 18108 5488 18136
rect 5813 18139 5871 18145
rect 4856 18096 4862 18108
rect 5813 18105 5825 18139
rect 5859 18136 5871 18139
rect 6549 18139 6607 18145
rect 6549 18136 6561 18139
rect 5859 18108 6561 18136
rect 5859 18105 5871 18108
rect 5813 18099 5871 18105
rect 6549 18105 6561 18108
rect 6595 18105 6607 18139
rect 6549 18099 6607 18105
rect 9217 18139 9275 18145
rect 9217 18105 9229 18139
rect 9263 18136 9275 18139
rect 9490 18136 9496 18148
rect 9263 18108 9496 18136
rect 9263 18105 9275 18108
rect 9217 18099 9275 18105
rect 9490 18096 9496 18108
rect 9548 18096 9554 18148
rect 9582 18096 9588 18148
rect 9640 18136 9646 18148
rect 9968 18145 9996 18176
rect 10229 18173 10241 18176
rect 10275 18173 10287 18207
rect 10229 18167 10287 18173
rect 11238 18164 11244 18216
rect 11296 18204 11302 18216
rect 12066 18204 12072 18216
rect 11296 18176 12072 18204
rect 11296 18164 11302 18176
rect 12066 18164 12072 18176
rect 12124 18204 12130 18216
rect 12268 18204 12296 18235
rect 12124 18176 12296 18204
rect 12124 18164 12130 18176
rect 13354 18164 13360 18216
rect 13412 18164 13418 18216
rect 14366 18213 14372 18216
rect 14364 18204 14372 18213
rect 14327 18176 14372 18204
rect 14364 18167 14372 18176
rect 14366 18164 14372 18167
rect 14424 18164 14430 18216
rect 14568 18213 14596 18244
rect 14751 18244 15148 18272
rect 14751 18213 14779 18244
rect 15120 18216 15148 18244
rect 15381 18241 15393 18275
rect 15427 18272 15439 18275
rect 15746 18272 15752 18284
rect 15427 18244 15752 18272
rect 15427 18241 15439 18244
rect 15381 18235 15439 18241
rect 15746 18232 15752 18244
rect 15804 18232 15810 18284
rect 15856 18272 15884 18312
rect 15933 18309 15945 18343
rect 15979 18340 15991 18343
rect 16298 18340 16304 18352
rect 15979 18312 16304 18340
rect 15979 18309 15991 18312
rect 15933 18303 15991 18309
rect 16298 18300 16304 18312
rect 16356 18300 16362 18352
rect 21361 18343 21419 18349
rect 21361 18309 21373 18343
rect 21407 18340 21419 18343
rect 21450 18340 21456 18352
rect 21407 18312 21456 18340
rect 21407 18309 21419 18312
rect 21361 18303 21419 18309
rect 21450 18300 21456 18312
rect 21508 18300 21514 18352
rect 16574 18272 16580 18284
rect 15856 18244 16580 18272
rect 16574 18232 16580 18244
rect 16632 18272 16638 18284
rect 17862 18272 17868 18284
rect 16632 18244 17264 18272
rect 16632 18232 16638 18244
rect 14553 18207 14611 18213
rect 14553 18173 14565 18207
rect 14599 18173 14611 18207
rect 14553 18167 14611 18173
rect 14736 18207 14794 18213
rect 14736 18173 14748 18207
rect 14782 18173 14794 18207
rect 14736 18167 14794 18173
rect 14829 18207 14887 18213
rect 14829 18173 14841 18207
rect 14875 18204 14887 18207
rect 15010 18204 15016 18216
rect 14875 18176 15016 18204
rect 14875 18173 14887 18176
rect 14829 18167 14887 18173
rect 9953 18139 10011 18145
rect 9953 18136 9965 18139
rect 9640 18108 9965 18136
rect 9640 18096 9646 18108
rect 9953 18105 9965 18108
rect 9999 18105 10011 18139
rect 9953 18099 10011 18105
rect 10496 18139 10554 18145
rect 10496 18105 10508 18139
rect 10542 18136 10554 18139
rect 10962 18136 10968 18148
rect 10542 18108 10968 18136
rect 10542 18105 10554 18108
rect 10496 18099 10554 18105
rect 10962 18096 10968 18108
rect 11020 18096 11026 18148
rect 11146 18096 11152 18148
rect 11204 18136 11210 18148
rect 11204 18108 11744 18136
rect 11204 18096 11210 18108
rect 1118 18028 1124 18080
rect 1176 18028 1182 18080
rect 1854 18028 1860 18080
rect 1912 18028 1918 18080
rect 1946 18028 1952 18080
rect 2004 18068 2010 18080
rect 2317 18071 2375 18077
rect 2317 18068 2329 18071
rect 2004 18040 2329 18068
rect 2004 18028 2010 18040
rect 2317 18037 2329 18040
rect 2363 18037 2375 18071
rect 2317 18031 2375 18037
rect 4893 18071 4951 18077
rect 4893 18037 4905 18071
rect 4939 18068 4951 18071
rect 5442 18068 5448 18080
rect 4939 18040 5448 18068
rect 4939 18037 4951 18040
rect 4893 18031 4951 18037
rect 5442 18028 5448 18040
rect 5500 18028 5506 18080
rect 5994 18028 6000 18080
rect 6052 18068 6058 18080
rect 6270 18068 6276 18080
rect 6052 18040 6276 18068
rect 6052 18028 6058 18040
rect 6270 18028 6276 18040
rect 6328 18028 6334 18080
rect 7653 18071 7711 18077
rect 7653 18037 7665 18071
rect 7699 18068 7711 18071
rect 7834 18068 7840 18080
rect 7699 18040 7840 18068
rect 7699 18037 7711 18040
rect 7653 18031 7711 18037
rect 7834 18028 7840 18040
rect 7892 18028 7898 18080
rect 8294 18028 8300 18080
rect 8352 18068 8358 18080
rect 8941 18071 8999 18077
rect 8941 18068 8953 18071
rect 8352 18040 8953 18068
rect 8352 18028 8358 18040
rect 8941 18037 8953 18040
rect 8987 18037 8999 18071
rect 8941 18031 8999 18037
rect 11422 18028 11428 18080
rect 11480 18068 11486 18080
rect 11716 18077 11744 18108
rect 12802 18096 12808 18148
rect 12860 18136 12866 18148
rect 13785 18139 13843 18145
rect 13785 18136 13797 18139
rect 12860 18108 13797 18136
rect 12860 18096 12866 18108
rect 13785 18105 13797 18108
rect 13831 18105 13843 18139
rect 13785 18099 13843 18105
rect 14001 18139 14059 18145
rect 14001 18105 14013 18139
rect 14047 18136 14059 18139
rect 14461 18139 14519 18145
rect 14047 18108 14320 18136
rect 14047 18105 14059 18108
rect 14001 18099 14059 18105
rect 14292 18080 14320 18108
rect 14461 18105 14473 18139
rect 14507 18105 14519 18139
rect 14568 18136 14596 18167
rect 15010 18164 15016 18176
rect 15068 18164 15074 18216
rect 15102 18164 15108 18216
rect 15160 18164 15166 18216
rect 16298 18164 16304 18216
rect 16356 18204 16362 18216
rect 17236 18213 17264 18244
rect 17604 18244 17868 18272
rect 17604 18213 17632 18244
rect 17862 18232 17868 18244
rect 17920 18232 17926 18284
rect 16485 18207 16543 18213
rect 16485 18204 16497 18207
rect 16356 18176 16497 18204
rect 16356 18164 16362 18176
rect 16485 18173 16497 18176
rect 16531 18173 16543 18207
rect 16485 18167 16543 18173
rect 17221 18207 17279 18213
rect 17221 18173 17233 18207
rect 17267 18173 17279 18207
rect 17221 18167 17279 18173
rect 17589 18207 17647 18213
rect 17589 18173 17601 18207
rect 17635 18173 17647 18207
rect 17589 18167 17647 18173
rect 17678 18164 17684 18216
rect 17736 18164 17742 18216
rect 17770 18164 17776 18216
rect 17828 18164 17834 18216
rect 17954 18164 17960 18216
rect 18012 18164 18018 18216
rect 18138 18164 18144 18216
rect 18196 18164 18202 18216
rect 18966 18164 18972 18216
rect 19024 18164 19030 18216
rect 20898 18164 20904 18216
rect 20956 18164 20962 18216
rect 20993 18207 21051 18213
rect 20993 18173 21005 18207
rect 21039 18173 21051 18207
rect 20993 18167 21051 18173
rect 14921 18139 14979 18145
rect 14921 18136 14933 18139
rect 14568 18108 14933 18136
rect 14461 18099 14519 18105
rect 14921 18105 14933 18108
rect 14967 18105 14979 18139
rect 14921 18099 14979 18105
rect 11609 18071 11667 18077
rect 11609 18068 11621 18071
rect 11480 18040 11621 18068
rect 11480 18028 11486 18040
rect 11609 18037 11621 18040
rect 11655 18037 11667 18071
rect 11609 18031 11667 18037
rect 11701 18071 11759 18077
rect 11701 18037 11713 18071
rect 11747 18037 11759 18071
rect 11701 18031 11759 18037
rect 12066 18028 12072 18080
rect 12124 18028 12130 18080
rect 13630 18028 13636 18080
rect 13688 18028 13694 18080
rect 14182 18028 14188 18080
rect 14240 18028 14246 18080
rect 14274 18028 14280 18080
rect 14332 18028 14338 18080
rect 14476 18068 14504 18099
rect 15838 18096 15844 18148
rect 15896 18136 15902 18148
rect 16025 18139 16083 18145
rect 16025 18136 16037 18139
rect 15896 18108 16037 18136
rect 15896 18096 15902 18108
rect 16025 18105 16037 18108
rect 16071 18105 16083 18139
rect 16025 18099 16083 18105
rect 16114 18096 16120 18148
rect 16172 18136 16178 18148
rect 16209 18139 16267 18145
rect 16209 18136 16221 18139
rect 16172 18108 16221 18136
rect 16172 18096 16178 18108
rect 16209 18105 16221 18108
rect 16255 18105 16267 18139
rect 16209 18099 16267 18105
rect 19236 18139 19294 18145
rect 19236 18105 19248 18139
rect 19282 18136 19294 18139
rect 19426 18136 19432 18148
rect 19282 18108 19432 18136
rect 19282 18105 19294 18108
rect 19236 18099 19294 18105
rect 19426 18096 19432 18108
rect 19484 18096 19490 18148
rect 21008 18136 21036 18167
rect 21174 18164 21180 18216
rect 21232 18213 21238 18216
rect 21232 18207 21281 18213
rect 21232 18173 21235 18207
rect 21269 18173 21281 18207
rect 21232 18167 21281 18173
rect 21232 18164 21238 18167
rect 21358 18164 21364 18216
rect 21416 18164 21422 18216
rect 21652 18213 21680 18380
rect 22066 18340 22094 18380
rect 22462 18368 22468 18420
rect 22520 18408 22526 18420
rect 22741 18411 22799 18417
rect 22741 18408 22753 18411
rect 22520 18380 22753 18408
rect 22520 18368 22526 18380
rect 22741 18377 22753 18380
rect 22787 18377 22799 18411
rect 23290 18408 23296 18420
rect 22741 18371 22799 18377
rect 22848 18380 23296 18408
rect 22848 18340 22876 18380
rect 23290 18368 23296 18380
rect 23348 18368 23354 18420
rect 23382 18368 23388 18420
rect 23440 18408 23446 18420
rect 24213 18411 24271 18417
rect 24213 18408 24225 18411
rect 23440 18380 24225 18408
rect 23440 18368 23446 18380
rect 24213 18377 24225 18380
rect 24259 18377 24271 18411
rect 24213 18371 24271 18377
rect 25041 18411 25099 18417
rect 25041 18377 25053 18411
rect 25087 18408 25099 18411
rect 25317 18411 25375 18417
rect 25317 18408 25329 18411
rect 25087 18380 25329 18408
rect 25087 18377 25099 18380
rect 25041 18371 25099 18377
rect 25317 18377 25329 18380
rect 25363 18377 25375 18411
rect 25317 18371 25375 18377
rect 25498 18368 25504 18420
rect 25556 18368 25562 18420
rect 22066 18312 22876 18340
rect 23109 18343 23167 18349
rect 23109 18309 23121 18343
rect 23155 18340 23167 18343
rect 23569 18343 23627 18349
rect 23569 18340 23581 18343
rect 23155 18312 23581 18340
rect 23155 18309 23167 18312
rect 23109 18303 23167 18309
rect 23569 18309 23581 18312
rect 23615 18340 23627 18343
rect 24394 18340 24400 18352
rect 23615 18312 24400 18340
rect 23615 18309 23627 18312
rect 23569 18303 23627 18309
rect 24394 18300 24400 18312
rect 24452 18300 24458 18352
rect 24854 18300 24860 18352
rect 24912 18340 24918 18352
rect 25685 18343 25743 18349
rect 25685 18340 25697 18343
rect 24912 18312 25697 18340
rect 24912 18300 24918 18312
rect 25685 18309 25697 18312
rect 25731 18309 25743 18343
rect 25685 18303 25743 18309
rect 21818 18232 21824 18284
rect 21876 18272 21882 18284
rect 22554 18272 22560 18284
rect 21876 18244 22560 18272
rect 21876 18232 21882 18244
rect 22554 18232 22560 18244
rect 22612 18232 22618 18284
rect 23198 18272 23204 18284
rect 22848 18244 23204 18272
rect 21637 18207 21695 18213
rect 21637 18173 21649 18207
rect 21683 18173 21695 18207
rect 21637 18167 21695 18173
rect 22005 18207 22063 18213
rect 22005 18173 22017 18207
rect 22051 18173 22063 18207
rect 22005 18167 22063 18173
rect 22281 18207 22339 18213
rect 22281 18173 22293 18207
rect 22327 18204 22339 18207
rect 22848 18204 22876 18244
rect 23198 18232 23204 18244
rect 23256 18232 23262 18284
rect 24320 18244 24624 18272
rect 24320 18213 24348 18244
rect 22327 18176 22876 18204
rect 23385 18207 23443 18213
rect 22327 18173 22339 18176
rect 22281 18167 22339 18173
rect 23385 18173 23397 18207
rect 23431 18173 23443 18207
rect 23845 18207 23903 18213
rect 23845 18204 23857 18207
rect 23385 18167 23443 18173
rect 23492 18176 23857 18204
rect 21726 18136 21732 18148
rect 21008 18108 21732 18136
rect 21726 18096 21732 18108
rect 21784 18096 21790 18148
rect 22020 18136 22048 18167
rect 22370 18136 22376 18148
rect 22020 18108 22376 18136
rect 22370 18096 22376 18108
rect 22428 18096 22434 18148
rect 22465 18139 22523 18145
rect 22465 18105 22477 18139
rect 22511 18136 22523 18139
rect 22741 18139 22799 18145
rect 22741 18136 22753 18139
rect 22511 18108 22753 18136
rect 22511 18105 22523 18108
rect 22465 18099 22523 18105
rect 22741 18105 22753 18108
rect 22787 18105 22799 18139
rect 22741 18099 22799 18105
rect 22830 18096 22836 18148
rect 22888 18136 22894 18148
rect 23400 18136 23428 18167
rect 22888 18108 23428 18136
rect 22888 18096 22894 18108
rect 15194 18068 15200 18080
rect 14476 18040 15200 18068
rect 15194 18028 15200 18040
rect 15252 18028 15258 18080
rect 15286 18028 15292 18080
rect 15344 18028 15350 18080
rect 15378 18028 15384 18080
rect 15436 18068 15442 18080
rect 15749 18071 15807 18077
rect 15749 18068 15761 18071
rect 15436 18040 15761 18068
rect 15436 18028 15442 18040
rect 15749 18037 15761 18040
rect 15795 18037 15807 18071
rect 15749 18031 15807 18037
rect 17129 18071 17187 18077
rect 17129 18037 17141 18071
rect 17175 18068 17187 18071
rect 17586 18068 17592 18080
rect 17175 18040 17592 18068
rect 17175 18037 17187 18040
rect 17129 18031 17187 18037
rect 17586 18028 17592 18040
rect 17644 18068 17650 18080
rect 17770 18068 17776 18080
rect 17644 18040 17776 18068
rect 17644 18028 17650 18040
rect 17770 18028 17776 18040
rect 17828 18028 17834 18080
rect 20717 18071 20775 18077
rect 20717 18037 20729 18071
rect 20763 18068 20775 18071
rect 21545 18071 21603 18077
rect 21545 18068 21557 18071
rect 20763 18040 21557 18068
rect 20763 18037 20775 18040
rect 20717 18031 20775 18037
rect 21545 18037 21557 18040
rect 21591 18037 21603 18071
rect 21545 18031 21603 18037
rect 22094 18028 22100 18080
rect 22152 18028 22158 18080
rect 22557 18071 22615 18077
rect 22557 18037 22569 18071
rect 22603 18068 22615 18071
rect 23492 18068 23520 18176
rect 23845 18173 23857 18176
rect 23891 18173 23903 18207
rect 23845 18167 23903 18173
rect 24305 18207 24363 18213
rect 24305 18173 24317 18207
rect 24351 18173 24363 18207
rect 24305 18167 24363 18173
rect 24394 18164 24400 18216
rect 24452 18204 24458 18216
rect 24596 18213 24624 18244
rect 24581 18207 24639 18213
rect 24452 18176 24532 18204
rect 24452 18164 24458 18176
rect 24504 18136 24532 18176
rect 24581 18173 24593 18207
rect 24627 18204 24639 18207
rect 24762 18204 24768 18216
rect 24627 18176 24768 18204
rect 24627 18173 24639 18176
rect 24581 18167 24639 18173
rect 24762 18164 24768 18176
rect 24820 18204 24826 18216
rect 24857 18207 24915 18213
rect 24857 18204 24869 18207
rect 24820 18176 24869 18204
rect 24820 18164 24826 18176
rect 24857 18173 24869 18176
rect 24903 18173 24915 18207
rect 24857 18167 24915 18173
rect 27062 18164 27068 18216
rect 27120 18164 27126 18216
rect 24673 18139 24731 18145
rect 24673 18136 24685 18139
rect 24504 18108 24685 18136
rect 24673 18105 24685 18108
rect 24719 18105 24731 18139
rect 24673 18099 24731 18105
rect 25130 18096 25136 18148
rect 25188 18136 25194 18148
rect 25498 18136 25504 18148
rect 25188 18108 25504 18136
rect 25188 18096 25194 18108
rect 25498 18096 25504 18108
rect 25556 18096 25562 18148
rect 26602 18096 26608 18148
rect 26660 18136 26666 18148
rect 26798 18139 26856 18145
rect 26798 18136 26810 18139
rect 26660 18108 26810 18136
rect 26660 18096 26666 18108
rect 26798 18105 26810 18108
rect 26844 18105 26856 18139
rect 26798 18099 26856 18105
rect 22603 18040 23520 18068
rect 22603 18037 22615 18040
rect 22557 18031 22615 18037
rect 23934 18028 23940 18080
rect 23992 18068 23998 18080
rect 24029 18071 24087 18077
rect 24029 18068 24041 18071
rect 23992 18040 24041 18068
rect 23992 18028 23998 18040
rect 24029 18037 24041 18040
rect 24075 18037 24087 18071
rect 24029 18031 24087 18037
rect 24581 18071 24639 18077
rect 24581 18037 24593 18071
rect 24627 18068 24639 18071
rect 25333 18071 25391 18077
rect 25333 18068 25345 18071
rect 24627 18040 25345 18068
rect 24627 18037 24639 18040
rect 24581 18031 24639 18037
rect 25333 18037 25345 18040
rect 25379 18068 25391 18071
rect 25774 18068 25780 18080
rect 25379 18040 25780 18068
rect 25379 18037 25391 18040
rect 25333 18031 25391 18037
rect 25774 18028 25780 18040
rect 25832 18068 25838 18080
rect 26142 18068 26148 18080
rect 25832 18040 26148 18068
rect 25832 18028 25838 18040
rect 26142 18028 26148 18040
rect 26200 18028 26206 18080
rect 552 17978 27576 18000
rect 552 17926 7114 17978
rect 7166 17926 7178 17978
rect 7230 17926 7242 17978
rect 7294 17926 7306 17978
rect 7358 17926 7370 17978
rect 7422 17926 13830 17978
rect 13882 17926 13894 17978
rect 13946 17926 13958 17978
rect 14010 17926 14022 17978
rect 14074 17926 14086 17978
rect 14138 17926 20546 17978
rect 20598 17926 20610 17978
rect 20662 17926 20674 17978
rect 20726 17926 20738 17978
rect 20790 17926 20802 17978
rect 20854 17926 27262 17978
rect 27314 17926 27326 17978
rect 27378 17926 27390 17978
rect 27442 17926 27454 17978
rect 27506 17926 27518 17978
rect 27570 17926 27576 17978
rect 552 17904 27576 17926
rect 2222 17824 2228 17876
rect 2280 17824 2286 17876
rect 4433 17867 4491 17873
rect 4433 17833 4445 17867
rect 4479 17864 4491 17867
rect 4522 17864 4528 17876
rect 4479 17836 4528 17864
rect 4479 17833 4491 17836
rect 4433 17827 4491 17833
rect 4522 17824 4528 17836
rect 4580 17824 4586 17876
rect 4798 17824 4804 17876
rect 4856 17864 4862 17876
rect 4893 17867 4951 17873
rect 4893 17864 4905 17867
rect 4856 17836 4905 17864
rect 4856 17824 4862 17836
rect 4893 17833 4905 17836
rect 4939 17833 4951 17867
rect 4893 17827 4951 17833
rect 6625 17867 6683 17873
rect 6625 17833 6637 17867
rect 6671 17864 6683 17867
rect 6671 17836 7061 17864
rect 6671 17833 6683 17836
rect 6625 17827 6683 17833
rect 1118 17805 1124 17808
rect 1112 17796 1124 17805
rect 1079 17768 1124 17796
rect 1112 17759 1124 17768
rect 1118 17756 1124 17759
rect 1176 17756 1182 17808
rect 842 17688 848 17740
rect 900 17688 906 17740
rect 2240 17728 2268 17824
rect 4709 17799 4767 17805
rect 2746 17768 4384 17796
rect 2593 17731 2651 17737
rect 2593 17728 2605 17731
rect 2240 17700 2605 17728
rect 2593 17697 2605 17700
rect 2639 17728 2651 17731
rect 2746 17728 2774 17768
rect 2639 17700 2774 17728
rect 2639 17697 2651 17700
rect 2593 17691 2651 17697
rect 3050 17688 3056 17740
rect 3108 17728 3114 17740
rect 4356 17737 4384 17768
rect 4709 17765 4721 17799
rect 4755 17796 4767 17799
rect 5534 17796 5540 17808
rect 4755 17768 5540 17796
rect 4755 17765 4767 17768
rect 4709 17759 4767 17765
rect 4065 17731 4123 17737
rect 4065 17728 4077 17731
rect 3108 17700 4077 17728
rect 3108 17688 3114 17700
rect 4065 17697 4077 17700
rect 4111 17697 4123 17731
rect 4065 17691 4123 17697
rect 4341 17731 4399 17737
rect 4341 17697 4353 17731
rect 4387 17728 4399 17731
rect 4522 17728 4528 17740
rect 4387 17700 4528 17728
rect 4387 17697 4399 17700
rect 4341 17691 4399 17697
rect 4522 17688 4528 17700
rect 4580 17688 4586 17740
rect 4617 17731 4675 17737
rect 4617 17697 4629 17731
rect 4663 17697 4675 17731
rect 4617 17691 4675 17697
rect 5077 17731 5135 17737
rect 5077 17697 5089 17731
rect 5123 17697 5135 17731
rect 5077 17691 5135 17697
rect 2409 17663 2467 17669
rect 2409 17629 2421 17663
rect 2455 17629 2467 17663
rect 2409 17623 2467 17629
rect 2424 17592 2452 17623
rect 2498 17620 2504 17672
rect 2556 17620 2562 17672
rect 2682 17620 2688 17672
rect 2740 17620 2746 17672
rect 3973 17663 4031 17669
rect 3973 17629 3985 17663
rect 4019 17660 4031 17663
rect 4154 17660 4160 17672
rect 4019 17632 4160 17660
rect 4019 17629 4031 17632
rect 3973 17623 4031 17629
rect 4154 17620 4160 17632
rect 4212 17620 4218 17672
rect 3234 17592 3240 17604
rect 2424 17564 3240 17592
rect 3234 17552 3240 17564
rect 3292 17592 3298 17604
rect 4632 17592 4660 17691
rect 5092 17660 5120 17691
rect 5166 17688 5172 17740
rect 5224 17688 5230 17740
rect 5460 17737 5488 17768
rect 5534 17756 5540 17768
rect 5592 17756 5598 17808
rect 6825 17799 6883 17805
rect 6825 17796 6837 17799
rect 6748 17768 6837 17796
rect 5445 17731 5503 17737
rect 5445 17697 5457 17731
rect 5491 17697 5503 17731
rect 5445 17691 5503 17697
rect 6273 17731 6331 17737
rect 6273 17697 6285 17731
rect 6319 17728 6331 17731
rect 6454 17728 6460 17740
rect 6319 17700 6460 17728
rect 6319 17697 6331 17700
rect 6273 17691 6331 17697
rect 6454 17688 6460 17700
rect 6512 17688 6518 17740
rect 6748 17728 6776 17768
rect 6825 17765 6837 17768
rect 6871 17765 6883 17799
rect 6825 17759 6883 17765
rect 6914 17756 6920 17808
rect 6972 17756 6978 17808
rect 7033 17796 7061 17836
rect 7282 17824 7288 17876
rect 7340 17864 7346 17876
rect 8113 17867 8171 17873
rect 8113 17864 8125 17867
rect 7340 17836 8125 17864
rect 7340 17824 7346 17836
rect 8113 17833 8125 17836
rect 8159 17833 8171 17867
rect 8113 17827 8171 17833
rect 10042 17824 10048 17876
rect 10100 17824 10106 17876
rect 10962 17824 10968 17876
rect 11020 17824 11026 17876
rect 11701 17867 11759 17873
rect 11701 17833 11713 17867
rect 11747 17864 11759 17867
rect 12066 17864 12072 17876
rect 11747 17836 12072 17864
rect 11747 17833 11759 17836
rect 11701 17827 11759 17833
rect 12066 17824 12072 17836
rect 12124 17824 12130 17876
rect 13354 17824 13360 17876
rect 13412 17864 13418 17876
rect 13541 17867 13599 17873
rect 13541 17864 13553 17867
rect 13412 17836 13553 17864
rect 13412 17824 13418 17836
rect 13541 17833 13553 17836
rect 13587 17833 13599 17867
rect 13541 17827 13599 17833
rect 7117 17799 7175 17805
rect 7117 17796 7129 17799
rect 7033 17768 7129 17796
rect 7117 17765 7129 17768
rect 7163 17796 7175 17799
rect 7466 17796 7472 17808
rect 7163 17768 7472 17796
rect 7163 17765 7175 17768
rect 7117 17759 7175 17765
rect 7466 17756 7472 17768
rect 7524 17756 7530 17808
rect 7377 17731 7435 17737
rect 7377 17728 7389 17731
rect 6748 17700 7389 17728
rect 7377 17697 7389 17700
rect 7423 17697 7435 17731
rect 7377 17691 7435 17697
rect 9401 17731 9459 17737
rect 9401 17697 9413 17731
rect 9447 17728 9459 17731
rect 9953 17731 10011 17737
rect 9447 17700 9628 17728
rect 9447 17697 9459 17700
rect 9401 17691 9459 17697
rect 7466 17660 7472 17672
rect 5092 17632 7472 17660
rect 7466 17620 7472 17632
rect 7524 17660 7530 17672
rect 7929 17663 7987 17669
rect 7929 17660 7941 17663
rect 7524 17632 7941 17660
rect 7524 17620 7530 17632
rect 7929 17629 7941 17632
rect 7975 17629 7987 17663
rect 7929 17623 7987 17629
rect 8662 17620 8668 17672
rect 8720 17620 8726 17672
rect 7285 17595 7343 17601
rect 3292 17564 6040 17592
rect 3292 17552 3298 17564
rect 2866 17484 2872 17536
rect 2924 17484 2930 17536
rect 3326 17484 3332 17536
rect 3384 17484 3390 17536
rect 4249 17527 4307 17533
rect 4249 17493 4261 17527
rect 4295 17524 4307 17527
rect 4338 17524 4344 17536
rect 4295 17496 4344 17524
rect 4295 17493 4307 17496
rect 4249 17487 4307 17493
rect 4338 17484 4344 17496
rect 4396 17484 4402 17536
rect 5353 17527 5411 17533
rect 5353 17493 5365 17527
rect 5399 17524 5411 17527
rect 5534 17524 5540 17536
rect 5399 17496 5540 17524
rect 5399 17493 5411 17496
rect 5353 17487 5411 17493
rect 5534 17484 5540 17496
rect 5592 17484 5598 17536
rect 5626 17484 5632 17536
rect 5684 17524 5690 17536
rect 6012 17533 6040 17564
rect 7285 17561 7297 17595
rect 7331 17592 7343 17595
rect 7834 17592 7840 17604
rect 7331 17564 7840 17592
rect 7331 17561 7343 17564
rect 7285 17555 7343 17561
rect 7834 17552 7840 17564
rect 7892 17552 7898 17604
rect 9600 17601 9628 17700
rect 9953 17697 9965 17731
rect 9999 17728 10011 17731
rect 10226 17728 10232 17740
rect 9999 17700 10232 17728
rect 9999 17697 10011 17700
rect 9953 17691 10011 17697
rect 10226 17688 10232 17700
rect 10284 17688 10290 17740
rect 11146 17688 11152 17740
rect 11204 17688 11210 17740
rect 11422 17688 11428 17740
rect 11480 17688 11486 17740
rect 11514 17688 11520 17740
rect 11572 17688 11578 17740
rect 12434 17737 12440 17740
rect 12428 17691 12440 17737
rect 12434 17688 12440 17691
rect 12492 17688 12498 17740
rect 13556 17728 13584 17827
rect 14274 17824 14280 17876
rect 14332 17864 14338 17876
rect 14461 17867 14519 17873
rect 14461 17864 14473 17867
rect 14332 17836 14473 17864
rect 14332 17824 14338 17836
rect 14461 17833 14473 17836
rect 14507 17833 14519 17867
rect 14461 17827 14519 17833
rect 15565 17867 15623 17873
rect 15565 17833 15577 17867
rect 15611 17864 15623 17867
rect 15654 17864 15660 17876
rect 15611 17836 15660 17864
rect 15611 17833 15623 17836
rect 15565 17827 15623 17833
rect 15654 17824 15660 17836
rect 15712 17824 15718 17876
rect 17954 17824 17960 17876
rect 18012 17864 18018 17876
rect 18509 17867 18567 17873
rect 18509 17864 18521 17867
rect 18012 17836 18521 17864
rect 18012 17824 18018 17836
rect 18509 17833 18521 17836
rect 18555 17833 18567 17867
rect 18509 17827 18567 17833
rect 21269 17867 21327 17873
rect 21269 17833 21281 17867
rect 21315 17864 21327 17867
rect 21358 17864 21364 17876
rect 21315 17836 21364 17864
rect 21315 17833 21327 17836
rect 21269 17827 21327 17833
rect 21358 17824 21364 17836
rect 21416 17824 21422 17876
rect 22833 17867 22891 17873
rect 22833 17833 22845 17867
rect 22879 17864 22891 17867
rect 23198 17864 23204 17876
rect 22879 17836 23204 17864
rect 22879 17833 22891 17836
rect 22833 17827 22891 17833
rect 23198 17824 23204 17836
rect 23256 17824 23262 17876
rect 24394 17824 24400 17876
rect 24452 17864 24458 17876
rect 24489 17867 24547 17873
rect 24489 17864 24501 17867
rect 24452 17836 24501 17864
rect 24452 17824 24458 17836
rect 24489 17833 24501 17836
rect 24535 17833 24547 17867
rect 24489 17827 24547 17833
rect 24673 17867 24731 17873
rect 24673 17833 24685 17867
rect 24719 17864 24731 17867
rect 24854 17864 24860 17876
rect 24719 17836 24860 17864
rect 24719 17833 24731 17836
rect 24673 17827 24731 17833
rect 24854 17824 24860 17836
rect 24912 17824 24918 17876
rect 25501 17867 25559 17873
rect 25501 17833 25513 17867
rect 25547 17864 25559 17867
rect 26053 17867 26111 17873
rect 26053 17864 26065 17867
rect 25547 17836 26065 17864
rect 25547 17833 25559 17836
rect 25501 17827 25559 17833
rect 26053 17833 26065 17836
rect 26099 17833 26111 17867
rect 26053 17827 26111 17833
rect 26602 17824 26608 17876
rect 26660 17824 26666 17876
rect 14737 17799 14795 17805
rect 14737 17765 14749 17799
rect 14783 17796 14795 17799
rect 15286 17796 15292 17808
rect 14783 17768 15292 17796
rect 14783 17765 14795 17768
rect 14737 17759 14795 17765
rect 15286 17756 15292 17768
rect 15344 17756 15350 17808
rect 15580 17768 16896 17796
rect 13817 17731 13875 17737
rect 13817 17728 13829 17731
rect 13556 17700 13829 17728
rect 13817 17697 13829 17700
rect 13863 17697 13875 17731
rect 13817 17691 13875 17697
rect 14182 17688 14188 17740
rect 14240 17728 14246 17740
rect 14553 17731 14611 17737
rect 14553 17728 14565 17731
rect 14240 17700 14565 17728
rect 14240 17688 14246 17700
rect 14553 17697 14565 17700
rect 14599 17697 14611 17731
rect 14553 17691 14611 17697
rect 14829 17731 14887 17737
rect 14829 17697 14841 17731
rect 14875 17697 14887 17731
rect 14829 17691 14887 17697
rect 14921 17731 14979 17737
rect 14921 17697 14933 17731
rect 14967 17728 14979 17731
rect 15102 17728 15108 17740
rect 14967 17700 15108 17728
rect 14967 17697 14979 17700
rect 14921 17691 14979 17697
rect 10137 17663 10195 17669
rect 10137 17629 10149 17663
rect 10183 17660 10195 17663
rect 10183 17632 11192 17660
rect 10183 17629 10195 17632
rect 10137 17623 10195 17629
rect 11164 17604 11192 17632
rect 11882 17620 11888 17672
rect 11940 17660 11946 17672
rect 12161 17663 12219 17669
rect 12161 17660 12173 17663
rect 11940 17632 12173 17660
rect 11940 17620 11946 17632
rect 12161 17629 12173 17632
rect 12207 17629 12219 17663
rect 12161 17623 12219 17629
rect 9585 17595 9643 17601
rect 9585 17561 9597 17595
rect 9631 17561 9643 17595
rect 9585 17555 9643 17561
rect 11146 17552 11152 17604
rect 11204 17552 11210 17604
rect 14844 17592 14872 17691
rect 15102 17688 15108 17700
rect 15160 17688 15166 17740
rect 15197 17663 15255 17669
rect 15197 17629 15209 17663
rect 15243 17660 15255 17663
rect 15378 17660 15384 17672
rect 15243 17632 15384 17660
rect 15243 17629 15255 17632
rect 15197 17623 15255 17629
rect 15378 17620 15384 17632
rect 15436 17620 15442 17672
rect 15286 17592 15292 17604
rect 14844 17564 15292 17592
rect 15286 17552 15292 17564
rect 15344 17592 15350 17604
rect 15580 17592 15608 17768
rect 15657 17731 15715 17737
rect 15657 17697 15669 17731
rect 15703 17697 15715 17731
rect 15657 17691 15715 17697
rect 15749 17731 15807 17737
rect 15749 17697 15761 17731
rect 15795 17728 15807 17731
rect 15838 17728 15844 17740
rect 15795 17700 15844 17728
rect 15795 17697 15807 17700
rect 15749 17691 15807 17697
rect 15672 17660 15700 17691
rect 15838 17688 15844 17700
rect 15896 17688 15902 17740
rect 16868 17737 16896 17768
rect 17862 17756 17868 17808
rect 17920 17796 17926 17808
rect 19797 17799 19855 17805
rect 19797 17796 19809 17799
rect 17920 17768 19809 17796
rect 17920 17756 17926 17768
rect 19797 17765 19809 17768
rect 19843 17765 19855 17799
rect 19797 17759 19855 17765
rect 21174 17756 21180 17808
rect 21232 17796 21238 17808
rect 24581 17799 24639 17805
rect 21232 17768 24440 17796
rect 21232 17756 21238 17768
rect 15933 17731 15991 17737
rect 15933 17697 15945 17731
rect 15979 17728 15991 17731
rect 16301 17731 16359 17737
rect 16301 17728 16313 17731
rect 15979 17700 16313 17728
rect 15979 17697 15991 17700
rect 15933 17691 15991 17697
rect 16301 17697 16313 17700
rect 16347 17697 16359 17731
rect 16301 17691 16359 17697
rect 16853 17731 16911 17737
rect 16853 17697 16865 17731
rect 16899 17697 16911 17731
rect 16853 17691 16911 17697
rect 16942 17688 16948 17740
rect 17000 17728 17006 17740
rect 17037 17731 17095 17737
rect 17037 17728 17049 17731
rect 17000 17700 17049 17728
rect 17000 17688 17006 17700
rect 17037 17697 17049 17700
rect 17083 17697 17095 17731
rect 17037 17691 17095 17697
rect 17773 17731 17831 17737
rect 17773 17697 17785 17731
rect 17819 17697 17831 17731
rect 17773 17691 17831 17697
rect 17957 17731 18015 17737
rect 17957 17697 17969 17731
rect 18003 17728 18015 17731
rect 18230 17728 18236 17740
rect 18003 17700 18236 17728
rect 18003 17697 18015 17700
rect 17957 17691 18015 17697
rect 17788 17660 17816 17691
rect 18230 17688 18236 17700
rect 18288 17688 18294 17740
rect 19150 17688 19156 17740
rect 19208 17688 19214 17740
rect 19613 17731 19671 17737
rect 19613 17697 19625 17731
rect 19659 17697 19671 17731
rect 19613 17691 19671 17697
rect 18322 17660 18328 17672
rect 15672 17632 15884 17660
rect 17788 17632 18328 17660
rect 15344 17564 15608 17592
rect 15344 17552 15350 17564
rect 5813 17527 5871 17533
rect 5813 17524 5825 17527
rect 5684 17496 5825 17524
rect 5684 17484 5690 17496
rect 5813 17493 5825 17496
rect 5859 17493 5871 17527
rect 5813 17487 5871 17493
rect 5997 17527 6055 17533
rect 5997 17493 6009 17527
rect 6043 17493 6055 17527
rect 5997 17487 6055 17493
rect 6454 17484 6460 17536
rect 6512 17484 6518 17536
rect 6641 17527 6699 17533
rect 6641 17493 6653 17527
rect 6687 17524 6699 17527
rect 7101 17527 7159 17533
rect 7101 17524 7113 17527
rect 6687 17496 7113 17524
rect 6687 17493 6699 17496
rect 6641 17487 6699 17493
rect 7101 17493 7113 17496
rect 7147 17524 7159 17527
rect 8110 17524 8116 17536
rect 7147 17496 8116 17524
rect 7147 17493 7159 17496
rect 7101 17487 7159 17493
rect 8110 17484 8116 17496
rect 8168 17484 8174 17536
rect 9030 17484 9036 17536
rect 9088 17524 9094 17536
rect 9217 17527 9275 17533
rect 9217 17524 9229 17527
rect 9088 17496 9229 17524
rect 9088 17484 9094 17496
rect 9217 17493 9229 17496
rect 9263 17493 9275 17527
rect 9217 17487 9275 17493
rect 14734 17484 14740 17536
rect 14792 17524 14798 17536
rect 15105 17527 15163 17533
rect 15105 17524 15117 17527
rect 14792 17496 15117 17524
rect 14792 17484 14798 17496
rect 15105 17493 15117 17496
rect 15151 17493 15163 17527
rect 15105 17487 15163 17493
rect 15381 17527 15439 17533
rect 15381 17493 15393 17527
rect 15427 17524 15439 17527
rect 15746 17524 15752 17536
rect 15427 17496 15752 17524
rect 15427 17493 15439 17496
rect 15381 17487 15439 17493
rect 15746 17484 15752 17496
rect 15804 17484 15810 17536
rect 15856 17533 15884 17632
rect 18322 17620 18328 17632
rect 18380 17660 18386 17672
rect 19628 17660 19656 17691
rect 19702 17688 19708 17740
rect 19760 17728 19766 17740
rect 19886 17728 19892 17740
rect 19760 17700 19892 17728
rect 19760 17688 19766 17700
rect 19886 17688 19892 17700
rect 19944 17688 19950 17740
rect 19981 17731 20039 17737
rect 19981 17697 19993 17731
rect 20027 17728 20039 17731
rect 20346 17728 20352 17740
rect 20027 17700 20352 17728
rect 20027 17697 20039 17700
rect 19981 17691 20039 17697
rect 20346 17688 20352 17700
rect 20404 17688 20410 17740
rect 20990 17688 20996 17740
rect 21048 17728 21054 17740
rect 21407 17731 21465 17737
rect 21407 17728 21419 17731
rect 21048 17700 21419 17728
rect 21048 17688 21054 17700
rect 21407 17697 21419 17700
rect 21453 17697 21465 17731
rect 21407 17691 21465 17697
rect 21542 17688 21548 17740
rect 21600 17688 21606 17740
rect 21634 17688 21640 17740
rect 21692 17688 21698 17740
rect 21775 17737 21803 17768
rect 21765 17731 21823 17737
rect 21765 17697 21777 17731
rect 21811 17697 21823 17731
rect 21765 17691 21823 17697
rect 21910 17688 21916 17740
rect 21968 17688 21974 17740
rect 22186 17737 22192 17740
rect 22005 17731 22063 17737
rect 22005 17697 22017 17731
rect 22051 17697 22063 17731
rect 22005 17691 22063 17697
rect 22159 17731 22192 17737
rect 22159 17697 22171 17731
rect 22159 17691 22192 17697
rect 18380 17632 19656 17660
rect 22020 17660 22048 17691
rect 22186 17688 22192 17691
rect 22244 17688 22250 17740
rect 23934 17688 23940 17740
rect 23992 17737 23998 17740
rect 23992 17728 24004 17737
rect 24412 17728 24440 17768
rect 24581 17765 24593 17799
rect 24627 17796 24639 17799
rect 24762 17796 24768 17808
rect 24627 17768 24768 17796
rect 24627 17765 24639 17768
rect 24581 17759 24639 17765
rect 24762 17756 24768 17768
rect 24820 17756 24826 17808
rect 27062 17796 27068 17808
rect 25884 17768 27068 17796
rect 24670 17728 24676 17740
rect 23992 17700 24037 17728
rect 24412 17700 24676 17728
rect 23992 17691 24004 17700
rect 23992 17688 23998 17691
rect 24670 17688 24676 17700
rect 24728 17728 24734 17740
rect 25682 17728 25688 17740
rect 24728 17700 25688 17728
rect 24728 17688 24734 17700
rect 25682 17688 25688 17700
rect 25740 17688 25746 17740
rect 25774 17688 25780 17740
rect 25832 17688 25838 17740
rect 24213 17663 24271 17669
rect 22020 17632 22094 17660
rect 18380 17620 18386 17632
rect 22066 17604 22094 17632
rect 24213 17629 24225 17663
rect 24259 17660 24271 17663
rect 25884 17660 25912 17768
rect 27062 17756 27068 17768
rect 27120 17756 27126 17808
rect 25958 17688 25964 17740
rect 26016 17728 26022 17740
rect 26053 17731 26111 17737
rect 26053 17728 26065 17731
rect 26016 17700 26065 17728
rect 26016 17688 26022 17700
rect 26053 17697 26065 17700
rect 26099 17697 26111 17731
rect 26053 17691 26111 17697
rect 26142 17688 26148 17740
rect 26200 17728 26206 17740
rect 26237 17731 26295 17737
rect 26237 17728 26249 17731
rect 26200 17700 26249 17728
rect 26200 17688 26206 17700
rect 26237 17697 26249 17700
rect 26283 17697 26295 17731
rect 26237 17691 26295 17697
rect 26418 17688 26424 17740
rect 26476 17688 26482 17740
rect 24259 17632 25912 17660
rect 24259 17629 24271 17632
rect 24213 17623 24271 17629
rect 16850 17552 16856 17604
rect 16908 17592 16914 17604
rect 19334 17592 19340 17604
rect 16908 17564 19340 17592
rect 16908 17552 16914 17564
rect 19334 17552 19340 17564
rect 19392 17552 19398 17604
rect 22066 17564 22100 17604
rect 22094 17552 22100 17564
rect 22152 17552 22158 17604
rect 22373 17595 22431 17601
rect 22373 17561 22385 17595
rect 22419 17592 22431 17595
rect 22462 17592 22468 17604
rect 22419 17564 22468 17592
rect 22419 17561 22431 17564
rect 22373 17555 22431 17561
rect 22462 17552 22468 17564
rect 22520 17592 22526 17604
rect 22922 17592 22928 17604
rect 22520 17564 22928 17592
rect 22520 17552 22526 17564
rect 22922 17552 22928 17564
rect 22980 17552 22986 17604
rect 24857 17595 24915 17601
rect 24857 17561 24869 17595
rect 24903 17592 24915 17595
rect 24946 17592 24952 17604
rect 24903 17564 24952 17592
rect 24903 17561 24915 17564
rect 24857 17555 24915 17561
rect 24946 17552 24952 17564
rect 25004 17552 25010 17604
rect 25038 17552 25044 17604
rect 25096 17592 25102 17604
rect 25133 17595 25191 17601
rect 25133 17592 25145 17595
rect 25096 17564 25145 17592
rect 25096 17552 25102 17564
rect 25133 17561 25145 17564
rect 25179 17592 25191 17595
rect 25777 17595 25835 17601
rect 25777 17592 25789 17595
rect 25179 17564 25789 17592
rect 25179 17561 25191 17564
rect 25133 17555 25191 17561
rect 25777 17561 25789 17564
rect 25823 17561 25835 17595
rect 25777 17555 25835 17561
rect 15841 17527 15899 17533
rect 15841 17493 15853 17527
rect 15887 17524 15899 17527
rect 16758 17524 16764 17536
rect 15887 17496 16764 17524
rect 15887 17493 15899 17496
rect 15841 17487 15899 17493
rect 16758 17484 16764 17496
rect 16816 17484 16822 17536
rect 17221 17527 17279 17533
rect 17221 17493 17233 17527
rect 17267 17524 17279 17527
rect 17586 17524 17592 17536
rect 17267 17496 17592 17524
rect 17267 17493 17279 17496
rect 17221 17487 17279 17493
rect 17586 17484 17592 17496
rect 17644 17484 17650 17536
rect 19429 17527 19487 17533
rect 19429 17493 19441 17527
rect 19475 17524 19487 17527
rect 19518 17524 19524 17536
rect 19475 17496 19524 17524
rect 19475 17493 19487 17496
rect 19429 17487 19487 17493
rect 19518 17484 19524 17496
rect 19576 17484 19582 17536
rect 24302 17484 24308 17536
rect 24360 17484 24366 17536
rect 25498 17484 25504 17536
rect 25556 17484 25562 17536
rect 25685 17527 25743 17533
rect 25685 17493 25697 17527
rect 25731 17524 25743 17527
rect 26418 17524 26424 17536
rect 25731 17496 26424 17524
rect 25731 17493 25743 17496
rect 25685 17487 25743 17493
rect 26418 17484 26424 17496
rect 26476 17484 26482 17536
rect 552 17434 27416 17456
rect 552 17382 3756 17434
rect 3808 17382 3820 17434
rect 3872 17382 3884 17434
rect 3936 17382 3948 17434
rect 4000 17382 4012 17434
rect 4064 17382 10472 17434
rect 10524 17382 10536 17434
rect 10588 17382 10600 17434
rect 10652 17382 10664 17434
rect 10716 17382 10728 17434
rect 10780 17382 17188 17434
rect 17240 17382 17252 17434
rect 17304 17382 17316 17434
rect 17368 17382 17380 17434
rect 17432 17382 17444 17434
rect 17496 17382 23904 17434
rect 23956 17382 23968 17434
rect 24020 17382 24032 17434
rect 24084 17382 24096 17434
rect 24148 17382 24160 17434
rect 24212 17382 27416 17434
rect 552 17360 27416 17382
rect 1302 17280 1308 17332
rect 1360 17280 1366 17332
rect 1486 17280 1492 17332
rect 1544 17280 1550 17332
rect 2222 17280 2228 17332
rect 2280 17280 2286 17332
rect 2869 17323 2927 17329
rect 2869 17320 2881 17323
rect 2746 17292 2881 17320
rect 1504 17184 1532 17280
rect 1854 17212 1860 17264
rect 1912 17212 1918 17264
rect 2409 17255 2467 17261
rect 2409 17221 2421 17255
rect 2455 17252 2467 17255
rect 2498 17252 2504 17264
rect 2455 17224 2504 17252
rect 2455 17221 2467 17224
rect 2409 17215 2467 17221
rect 2498 17212 2504 17224
rect 2556 17212 2562 17264
rect 2746 17196 2774 17292
rect 2869 17289 2881 17292
rect 2915 17289 2927 17323
rect 2869 17283 2927 17289
rect 3050 17280 3056 17332
rect 3108 17280 3114 17332
rect 3234 17280 3240 17332
rect 3292 17280 3298 17332
rect 4985 17323 5043 17329
rect 4985 17289 4997 17323
rect 5031 17320 5043 17323
rect 5166 17320 5172 17332
rect 5031 17292 5172 17320
rect 5031 17289 5043 17292
rect 4985 17283 5043 17289
rect 5166 17280 5172 17292
rect 5224 17280 5230 17332
rect 5258 17280 5264 17332
rect 5316 17320 5322 17332
rect 5813 17323 5871 17329
rect 5316 17292 5580 17320
rect 5316 17280 5322 17292
rect 2682 17184 2688 17196
rect 1504 17156 2688 17184
rect 2682 17144 2688 17156
rect 2740 17156 2774 17196
rect 2740 17144 2746 17156
rect 3252 17116 3280 17280
rect 5442 17252 5448 17264
rect 5184 17224 5448 17252
rect 5184 17193 5212 17224
rect 5442 17212 5448 17224
rect 5500 17212 5506 17264
rect 5552 17252 5580 17292
rect 5813 17289 5825 17323
rect 5859 17320 5871 17323
rect 6270 17320 6276 17332
rect 5859 17292 6276 17320
rect 5859 17289 5871 17292
rect 5813 17283 5871 17289
rect 6270 17280 6276 17292
rect 6328 17280 6334 17332
rect 6825 17323 6883 17329
rect 6825 17289 6837 17323
rect 6871 17320 6883 17323
rect 8662 17320 8668 17332
rect 6871 17292 8668 17320
rect 6871 17289 6883 17292
rect 6825 17283 6883 17289
rect 6840 17252 6868 17283
rect 8662 17280 8668 17292
rect 8720 17280 8726 17332
rect 12434 17280 12440 17332
rect 12492 17320 12498 17332
rect 12621 17323 12679 17329
rect 12621 17320 12633 17323
rect 12492 17292 12633 17320
rect 12492 17280 12498 17292
rect 12621 17289 12633 17292
rect 12667 17289 12679 17323
rect 12621 17283 12679 17289
rect 15378 17280 15384 17332
rect 15436 17320 15442 17332
rect 16666 17320 16672 17332
rect 15436 17292 16672 17320
rect 15436 17280 15442 17292
rect 16666 17280 16672 17292
rect 16724 17280 16730 17332
rect 18046 17280 18052 17332
rect 18104 17320 18110 17332
rect 20349 17323 20407 17329
rect 20349 17320 20361 17323
rect 18104 17292 20361 17320
rect 18104 17280 18110 17292
rect 20349 17289 20361 17292
rect 20395 17289 20407 17323
rect 20349 17283 20407 17289
rect 21729 17323 21787 17329
rect 21729 17289 21741 17323
rect 21775 17320 21787 17323
rect 22094 17320 22100 17332
rect 21775 17292 22100 17320
rect 21775 17289 21787 17292
rect 21729 17283 21787 17289
rect 22094 17280 22100 17292
rect 22152 17280 22158 17332
rect 5552 17224 6868 17252
rect 15105 17255 15163 17261
rect 15105 17221 15117 17255
rect 15151 17252 15163 17255
rect 15194 17252 15200 17264
rect 15151 17224 15200 17252
rect 15151 17221 15163 17224
rect 15105 17215 15163 17221
rect 15194 17212 15200 17224
rect 15252 17212 15258 17264
rect 15286 17212 15292 17264
rect 15344 17252 15350 17264
rect 16301 17255 16359 17261
rect 16301 17252 16313 17255
rect 15344 17224 16313 17252
rect 15344 17212 15350 17224
rect 16301 17221 16313 17224
rect 16347 17221 16359 17255
rect 17954 17252 17960 17264
rect 16301 17215 16359 17221
rect 17696 17224 17960 17252
rect 5169 17187 5227 17193
rect 5169 17153 5181 17187
rect 5215 17153 5227 17187
rect 5169 17147 5227 17153
rect 5350 17144 5356 17196
rect 5408 17184 5414 17196
rect 5905 17187 5963 17193
rect 5905 17184 5917 17187
rect 5408 17156 5917 17184
rect 5408 17144 5414 17156
rect 5905 17153 5917 17156
rect 5951 17184 5963 17187
rect 6546 17184 6552 17196
rect 5951 17156 6552 17184
rect 5951 17153 5963 17156
rect 5905 17147 5963 17153
rect 6546 17144 6552 17156
rect 6604 17144 6610 17196
rect 11149 17187 11207 17193
rect 11149 17153 11161 17187
rect 11195 17184 11207 17187
rect 11422 17184 11428 17196
rect 11195 17156 11428 17184
rect 11195 17153 11207 17156
rect 11149 17147 11207 17153
rect 11422 17144 11428 17156
rect 11480 17144 11486 17196
rect 13630 17184 13636 17196
rect 12820 17156 13636 17184
rect 2746 17088 3280 17116
rect 1489 17051 1547 17057
rect 1489 17017 1501 17051
rect 1535 17048 1547 17051
rect 1946 17048 1952 17060
rect 1535 17020 1952 17048
rect 1535 17017 1547 17020
rect 1489 17011 1547 17017
rect 1946 17008 1952 17020
rect 2004 17008 2010 17060
rect 2041 17051 2099 17057
rect 2041 17017 2053 17051
rect 2087 17048 2099 17051
rect 2746 17048 2774 17088
rect 4338 17076 4344 17128
rect 4396 17125 4402 17128
rect 4396 17116 4408 17125
rect 4617 17119 4675 17125
rect 4396 17088 4441 17116
rect 4396 17079 4408 17088
rect 4617 17085 4629 17119
rect 4663 17085 4675 17119
rect 4617 17079 4675 17085
rect 4396 17076 4402 17079
rect 2087 17020 2774 17048
rect 2087 17017 2099 17020
rect 2041 17011 2099 17017
rect 2866 17008 2872 17060
rect 2924 17008 2930 17060
rect 4632 17048 4660 17079
rect 4890 17076 4896 17128
rect 4948 17076 4954 17128
rect 4982 17076 4988 17128
rect 5040 17116 5046 17128
rect 5445 17119 5503 17125
rect 5445 17116 5457 17119
rect 5040 17088 5457 17116
rect 5040 17076 5046 17088
rect 5445 17085 5457 17088
rect 5491 17085 5503 17119
rect 5445 17079 5503 17085
rect 5626 17076 5632 17128
rect 5684 17076 5690 17128
rect 6454 17076 6460 17128
rect 6512 17076 6518 17128
rect 6638 17076 6644 17128
rect 6696 17076 6702 17128
rect 6733 17119 6791 17125
rect 6733 17085 6745 17119
rect 6779 17116 6791 17119
rect 7558 17116 7564 17128
rect 6779 17088 7564 17116
rect 6779 17085 6791 17088
rect 6733 17079 6791 17085
rect 7558 17076 7564 17088
rect 7616 17076 7622 17128
rect 8205 17119 8263 17125
rect 8205 17085 8217 17119
rect 8251 17116 8263 17119
rect 8386 17116 8392 17128
rect 8251 17088 8392 17116
rect 8251 17085 8263 17088
rect 8205 17079 8263 17085
rect 8386 17076 8392 17088
rect 8444 17116 8450 17128
rect 9030 17125 9036 17128
rect 8757 17119 8815 17125
rect 8757 17116 8769 17119
rect 8444 17088 8769 17116
rect 8444 17076 8450 17088
rect 8757 17085 8769 17088
rect 8803 17085 8815 17119
rect 9024 17116 9036 17125
rect 8991 17088 9036 17116
rect 8757 17079 8815 17085
rect 9024 17079 9036 17088
rect 9030 17076 9036 17079
rect 9088 17076 9094 17128
rect 10229 17119 10287 17125
rect 10229 17116 10241 17119
rect 10152 17088 10241 17116
rect 6086 17048 6092 17060
rect 4632 17020 6092 17048
rect 6086 17008 6092 17020
rect 6144 17008 6150 17060
rect 7650 17008 7656 17060
rect 7708 17048 7714 17060
rect 7938 17051 7996 17057
rect 7938 17048 7950 17051
rect 7708 17020 7950 17048
rect 7708 17008 7714 17020
rect 7938 17017 7950 17020
rect 7984 17017 7996 17051
rect 7938 17011 7996 17017
rect 10152 16992 10180 17088
rect 10229 17085 10241 17088
rect 10275 17085 10287 17119
rect 10229 17079 10287 17085
rect 11054 17076 11060 17128
rect 11112 17076 11118 17128
rect 12820 17125 12848 17156
rect 13630 17144 13636 17156
rect 13688 17144 13694 17196
rect 15746 17144 15752 17196
rect 15804 17144 15810 17196
rect 17696 17193 17724 17224
rect 17954 17212 17960 17224
rect 18012 17252 18018 17264
rect 18012 17224 18920 17252
rect 18012 17212 18018 17224
rect 17681 17187 17739 17193
rect 17681 17153 17693 17187
rect 17727 17153 17739 17187
rect 17681 17147 17739 17153
rect 12805 17119 12863 17125
rect 12805 17085 12817 17119
rect 12851 17085 12863 17119
rect 12805 17079 12863 17085
rect 13078 17076 13084 17128
rect 13136 17076 13142 17128
rect 13538 17076 13544 17128
rect 13596 17116 13602 17128
rect 13725 17119 13783 17125
rect 13725 17116 13737 17119
rect 13596 17088 13737 17116
rect 13596 17076 13602 17088
rect 13725 17085 13737 17088
rect 13771 17085 13783 17119
rect 16850 17116 16856 17128
rect 13725 17079 13783 17085
rect 13832 17088 16856 17116
rect 12710 17008 12716 17060
rect 12768 17048 12774 17060
rect 13832 17048 13860 17088
rect 16850 17076 16856 17088
rect 16908 17076 16914 17128
rect 17425 17119 17483 17125
rect 17425 17085 17437 17119
rect 17471 17116 17483 17119
rect 17586 17116 17592 17128
rect 17471 17088 17592 17116
rect 17471 17085 17483 17088
rect 17425 17079 17483 17085
rect 17586 17076 17592 17088
rect 17644 17076 17650 17128
rect 17957 17119 18015 17125
rect 17957 17085 17969 17119
rect 18003 17116 18015 17119
rect 18046 17116 18052 17128
rect 18003 17088 18052 17116
rect 18003 17085 18015 17088
rect 17957 17079 18015 17085
rect 18046 17076 18052 17088
rect 18104 17076 18110 17128
rect 18322 17076 18328 17128
rect 18380 17076 18386 17128
rect 18892 17125 18920 17224
rect 21542 17144 21548 17196
rect 21600 17184 21606 17196
rect 23937 17187 23995 17193
rect 23937 17184 23949 17187
rect 21600 17156 23949 17184
rect 21600 17144 21606 17156
rect 23937 17153 23949 17156
rect 23983 17153 23995 17187
rect 23937 17147 23995 17153
rect 18877 17119 18935 17125
rect 18877 17085 18889 17119
rect 18923 17116 18935 17119
rect 18966 17116 18972 17128
rect 18923 17088 18972 17116
rect 18923 17085 18935 17088
rect 18877 17079 18935 17085
rect 18966 17076 18972 17088
rect 19024 17116 19030 17128
rect 19024 17088 19288 17116
rect 19024 17076 19030 17088
rect 19260 17060 19288 17088
rect 20990 17076 20996 17128
rect 21048 17076 21054 17128
rect 21450 17076 21456 17128
rect 21508 17076 21514 17128
rect 22278 17076 22284 17128
rect 22336 17116 22342 17128
rect 22741 17119 22799 17125
rect 22741 17116 22753 17119
rect 22336 17088 22753 17116
rect 22336 17076 22342 17088
rect 22741 17085 22753 17088
rect 22787 17085 22799 17119
rect 22741 17079 22799 17085
rect 22922 17076 22928 17128
rect 22980 17116 22986 17128
rect 23109 17119 23167 17125
rect 23109 17116 23121 17119
rect 22980 17088 23121 17116
rect 22980 17076 22986 17088
rect 23109 17085 23121 17088
rect 23155 17085 23167 17119
rect 23109 17079 23167 17085
rect 23198 17076 23204 17128
rect 23256 17076 23262 17128
rect 24029 17119 24087 17125
rect 24029 17085 24041 17119
rect 24075 17085 24087 17119
rect 24029 17079 24087 17085
rect 12768 17020 13860 17048
rect 13992 17051 14050 17057
rect 12768 17008 12774 17020
rect 13992 17017 14004 17051
rect 14038 17048 14050 17051
rect 15197 17051 15255 17057
rect 15197 17048 15209 17051
rect 14038 17020 15209 17048
rect 14038 17017 14050 17020
rect 13992 17011 14050 17017
rect 15197 17017 15209 17020
rect 15243 17017 15255 17051
rect 15197 17011 15255 17017
rect 17862 17008 17868 17060
rect 17920 17048 17926 17060
rect 18141 17051 18199 17057
rect 18141 17048 18153 17051
rect 17920 17020 18153 17048
rect 17920 17008 17926 17020
rect 18141 17017 18153 17020
rect 18187 17017 18199 17051
rect 18141 17011 18199 17017
rect 18230 17008 18236 17060
rect 18288 17048 18294 17060
rect 18414 17048 18420 17060
rect 18288 17020 18420 17048
rect 18288 17008 18294 17020
rect 18414 17008 18420 17020
rect 18472 17008 18478 17060
rect 19122 17051 19180 17057
rect 19122 17048 19134 17051
rect 18524 17020 19134 17048
rect 1854 16940 1860 16992
rect 1912 16980 1918 16992
rect 2241 16983 2299 16989
rect 2241 16980 2253 16983
rect 1912 16952 2253 16980
rect 1912 16940 1918 16952
rect 2241 16949 2253 16952
rect 2287 16949 2299 16983
rect 2241 16943 2299 16949
rect 4154 16940 4160 16992
rect 4212 16980 4218 16992
rect 5350 16980 5356 16992
rect 4212 16952 5356 16980
rect 4212 16940 4218 16952
rect 5350 16940 5356 16952
rect 5408 16940 5414 16992
rect 5442 16940 5448 16992
rect 5500 16980 5506 16992
rect 5537 16983 5595 16989
rect 5537 16980 5549 16983
rect 5500 16952 5549 16980
rect 5500 16940 5506 16952
rect 5537 16949 5549 16952
rect 5583 16949 5595 16983
rect 5537 16943 5595 16949
rect 6273 16983 6331 16989
rect 6273 16949 6285 16983
rect 6319 16980 6331 16983
rect 6362 16980 6368 16992
rect 6319 16952 6368 16980
rect 6319 16949 6331 16952
rect 6273 16943 6331 16949
rect 6362 16940 6368 16952
rect 6420 16940 6426 16992
rect 10134 16940 10140 16992
rect 10192 16940 10198 16992
rect 10318 16940 10324 16992
rect 10376 16940 10382 16992
rect 10686 16940 10692 16992
rect 10744 16940 10750 16992
rect 12526 16940 12532 16992
rect 12584 16980 12590 16992
rect 12989 16983 13047 16989
rect 12989 16980 13001 16983
rect 12584 16952 13001 16980
rect 12584 16940 12590 16952
rect 12989 16949 13001 16952
rect 13035 16980 13047 16983
rect 13446 16980 13452 16992
rect 13035 16952 13452 16980
rect 13035 16949 13047 16952
rect 12989 16943 13047 16949
rect 13446 16940 13452 16952
rect 13504 16940 13510 16992
rect 13814 16940 13820 16992
rect 13872 16980 13878 16992
rect 16850 16980 16856 16992
rect 13872 16952 16856 16980
rect 13872 16940 13878 16952
rect 16850 16940 16856 16952
rect 16908 16980 16914 16992
rect 17218 16980 17224 16992
rect 16908 16952 17224 16980
rect 16908 16940 16914 16952
rect 17218 16940 17224 16952
rect 17276 16940 17282 16992
rect 18524 16989 18552 17020
rect 19122 17017 19134 17020
rect 19168 17017 19180 17051
rect 19122 17011 19180 17017
rect 19242 17008 19248 17060
rect 19300 17008 19306 17060
rect 21729 17051 21787 17057
rect 21729 17017 21741 17051
rect 21775 17048 21787 17051
rect 22002 17048 22008 17060
rect 21775 17020 22008 17048
rect 21775 17017 21787 17020
rect 21729 17011 21787 17017
rect 22002 17008 22008 17020
rect 22060 17008 22066 17060
rect 23566 17048 23572 17060
rect 23032 17020 23572 17048
rect 18509 16983 18567 16989
rect 18509 16949 18521 16983
rect 18555 16949 18567 16983
rect 18509 16943 18567 16949
rect 20257 16983 20315 16989
rect 20257 16949 20269 16983
rect 20303 16980 20315 16983
rect 20990 16980 20996 16992
rect 20303 16952 20996 16980
rect 20303 16949 20315 16952
rect 20257 16943 20315 16949
rect 20990 16940 20996 16952
rect 21048 16940 21054 16992
rect 21545 16983 21603 16989
rect 21545 16949 21557 16983
rect 21591 16980 21603 16983
rect 22370 16980 22376 16992
rect 21591 16952 22376 16980
rect 21591 16949 21603 16952
rect 21545 16943 21603 16949
rect 22370 16940 22376 16952
rect 22428 16940 22434 16992
rect 23032 16989 23060 17020
rect 23566 17008 23572 17020
rect 23624 17008 23630 17060
rect 24044 17048 24072 17079
rect 24118 17076 24124 17128
rect 24176 17116 24182 17128
rect 24213 17119 24271 17125
rect 24213 17116 24225 17119
rect 24176 17088 24225 17116
rect 24176 17076 24182 17088
rect 24213 17085 24225 17088
rect 24259 17085 24271 17119
rect 24213 17079 24271 17085
rect 25038 17076 25044 17128
rect 25096 17076 25102 17128
rect 25682 17076 25688 17128
rect 25740 17076 25746 17128
rect 24946 17048 24952 17060
rect 24044 17020 24952 17048
rect 24946 17008 24952 17020
rect 25004 17048 25010 17060
rect 25225 17051 25283 17057
rect 25225 17048 25237 17051
rect 25004 17020 25237 17048
rect 25004 17008 25010 17020
rect 25225 17017 25237 17020
rect 25271 17048 25283 17051
rect 25952 17051 26010 17057
rect 25271 17020 25544 17048
rect 25271 17017 25283 17020
rect 25225 17011 25283 17017
rect 23017 16983 23075 16989
rect 23017 16949 23029 16983
rect 23063 16949 23075 16983
rect 23017 16943 23075 16949
rect 24394 16940 24400 16992
rect 24452 16980 24458 16992
rect 24857 16983 24915 16989
rect 24857 16980 24869 16983
rect 24452 16952 24869 16980
rect 24452 16940 24458 16952
rect 24857 16949 24869 16952
rect 24903 16949 24915 16983
rect 24857 16943 24915 16949
rect 25314 16940 25320 16992
rect 25372 16980 25378 16992
rect 25409 16983 25467 16989
rect 25409 16980 25421 16983
rect 25372 16952 25421 16980
rect 25372 16940 25378 16952
rect 25409 16949 25421 16952
rect 25455 16949 25467 16983
rect 25516 16980 25544 17020
rect 25952 17017 25964 17051
rect 25998 17048 26010 17051
rect 26050 17048 26056 17060
rect 25998 17020 26056 17048
rect 25998 17017 26010 17020
rect 25952 17011 26010 17017
rect 26050 17008 26056 17020
rect 26108 17008 26114 17060
rect 27065 16983 27123 16989
rect 27065 16980 27077 16983
rect 25516 16952 27077 16980
rect 25409 16943 25467 16949
rect 27065 16949 27077 16952
rect 27111 16949 27123 16983
rect 27065 16943 27123 16949
rect 552 16890 27576 16912
rect 552 16838 7114 16890
rect 7166 16838 7178 16890
rect 7230 16838 7242 16890
rect 7294 16838 7306 16890
rect 7358 16838 7370 16890
rect 7422 16838 13830 16890
rect 13882 16838 13894 16890
rect 13946 16838 13958 16890
rect 14010 16838 14022 16890
rect 14074 16838 14086 16890
rect 14138 16838 20546 16890
rect 20598 16838 20610 16890
rect 20662 16838 20674 16890
rect 20726 16838 20738 16890
rect 20790 16838 20802 16890
rect 20854 16838 27262 16890
rect 27314 16838 27326 16890
rect 27378 16838 27390 16890
rect 27442 16838 27454 16890
rect 27506 16838 27518 16890
rect 27570 16838 27576 16890
rect 552 16816 27576 16838
rect 1578 16736 1584 16788
rect 1636 16776 1642 16788
rect 2406 16776 2412 16788
rect 1636 16748 2412 16776
rect 1636 16736 1642 16748
rect 2332 16649 2360 16748
rect 2406 16736 2412 16748
rect 2464 16736 2470 16788
rect 2682 16736 2688 16788
rect 2740 16776 2746 16788
rect 4338 16776 4344 16788
rect 2740 16748 4344 16776
rect 2740 16736 2746 16748
rect 4338 16736 4344 16748
rect 4396 16736 4402 16788
rect 4893 16779 4951 16785
rect 4893 16745 4905 16779
rect 4939 16776 4951 16779
rect 4982 16776 4988 16788
rect 4939 16748 4988 16776
rect 4939 16745 4951 16748
rect 4893 16739 4951 16745
rect 4982 16736 4988 16748
rect 5040 16736 5046 16788
rect 5442 16736 5448 16788
rect 5500 16736 5506 16788
rect 7466 16736 7472 16788
rect 7524 16736 7530 16788
rect 7650 16736 7656 16788
rect 7708 16736 7714 16788
rect 8018 16736 8024 16788
rect 8076 16736 8082 16788
rect 9677 16779 9735 16785
rect 9677 16745 9689 16779
rect 9723 16776 9735 16779
rect 10134 16776 10140 16788
rect 9723 16748 10140 16776
rect 9723 16745 9735 16748
rect 9677 16739 9735 16745
rect 10134 16736 10140 16748
rect 10192 16736 10198 16788
rect 10226 16736 10232 16788
rect 10284 16736 10290 16788
rect 11330 16736 11336 16788
rect 11388 16776 11394 16788
rect 11517 16779 11575 16785
rect 11517 16776 11529 16779
rect 11388 16748 11529 16776
rect 11388 16736 11394 16748
rect 11517 16745 11529 16748
rect 11563 16745 11575 16779
rect 11517 16739 11575 16745
rect 12802 16736 12808 16788
rect 12860 16776 12866 16788
rect 12963 16779 13021 16785
rect 12963 16776 12975 16779
rect 12860 16748 12975 16776
rect 12860 16736 12866 16748
rect 12963 16745 12975 16748
rect 13009 16776 13021 16779
rect 13722 16776 13728 16788
rect 13009 16748 13728 16776
rect 13009 16745 13021 16748
rect 12963 16739 13021 16745
rect 13722 16736 13728 16748
rect 13780 16776 13786 16788
rect 14001 16779 14059 16785
rect 14001 16776 14013 16779
rect 13780 16748 14013 16776
rect 13780 16736 13786 16748
rect 14001 16745 14013 16748
rect 14047 16745 14059 16779
rect 14458 16776 14464 16788
rect 14001 16739 14059 16745
rect 14200 16748 14464 16776
rect 2930 16711 2988 16717
rect 2930 16708 2942 16711
rect 2424 16680 2942 16708
rect 2317 16643 2375 16649
rect 2317 16609 2329 16643
rect 2363 16609 2375 16643
rect 2317 16603 2375 16609
rect 2133 16575 2191 16581
rect 2133 16541 2145 16575
rect 2179 16572 2191 16575
rect 2424 16572 2452 16680
rect 2930 16677 2942 16680
rect 2976 16677 2988 16711
rect 7484 16708 7512 16736
rect 14200 16720 14228 16748
rect 14458 16736 14464 16748
rect 14516 16736 14522 16788
rect 15286 16736 15292 16788
rect 15344 16776 15350 16788
rect 16485 16779 16543 16785
rect 15344 16748 16344 16776
rect 15344 16736 15350 16748
rect 2930 16671 2988 16677
rect 5000 16680 7512 16708
rect 2498 16600 2504 16652
rect 2556 16600 2562 16652
rect 2593 16643 2651 16649
rect 2593 16609 2605 16643
rect 2639 16640 2651 16643
rect 3326 16640 3332 16652
rect 2639 16612 3332 16640
rect 2639 16609 2651 16612
rect 2593 16603 2651 16609
rect 3326 16600 3332 16612
rect 3384 16600 3390 16652
rect 5000 16649 5028 16680
rect 7558 16668 7564 16720
rect 7616 16708 7622 16720
rect 9769 16711 9827 16717
rect 7616 16680 8156 16708
rect 7616 16668 7622 16680
rect 4433 16643 4491 16649
rect 4433 16609 4445 16643
rect 4479 16640 4491 16643
rect 4985 16643 5043 16649
rect 4479 16612 4936 16640
rect 4479 16609 4491 16612
rect 4433 16603 4491 16609
rect 2179 16544 2452 16572
rect 2685 16575 2743 16581
rect 2179 16541 2191 16544
rect 2133 16535 2191 16541
rect 2685 16541 2697 16575
rect 2731 16541 2743 16575
rect 4908 16572 4936 16612
rect 4985 16609 4997 16643
rect 5031 16609 5043 16643
rect 5258 16640 5264 16652
rect 4985 16603 5043 16609
rect 5092 16612 5264 16640
rect 5092 16572 5120 16612
rect 5258 16600 5264 16612
rect 5316 16600 5322 16652
rect 6086 16600 6092 16652
rect 6144 16600 6150 16652
rect 6362 16649 6368 16652
rect 6356 16640 6368 16649
rect 6323 16612 6368 16640
rect 6356 16603 6368 16612
rect 6362 16600 6368 16603
rect 6420 16600 6426 16652
rect 6638 16600 6644 16652
rect 6696 16640 6702 16652
rect 6822 16640 6828 16652
rect 6696 16612 6828 16640
rect 6696 16600 6702 16612
rect 6822 16600 6828 16612
rect 6880 16640 6886 16652
rect 6880 16612 7788 16640
rect 6880 16600 6886 16612
rect 4908 16544 5120 16572
rect 7760 16572 7788 16612
rect 7834 16600 7840 16652
rect 7892 16600 7898 16652
rect 8128 16649 8156 16680
rect 9769 16677 9781 16711
rect 9815 16708 9827 16711
rect 10686 16708 10692 16720
rect 9815 16680 10692 16708
rect 9815 16677 9827 16680
rect 9769 16671 9827 16677
rect 10686 16668 10692 16680
rect 10744 16668 10750 16720
rect 12710 16708 12716 16720
rect 10796 16680 12716 16708
rect 8113 16643 8171 16649
rect 8113 16609 8125 16643
rect 8159 16609 8171 16643
rect 10137 16643 10195 16649
rect 10137 16640 10149 16643
rect 8113 16603 8171 16609
rect 8220 16612 10149 16640
rect 8220 16572 8248 16612
rect 10137 16609 10149 16612
rect 10183 16640 10195 16643
rect 10183 16612 10272 16640
rect 10183 16609 10195 16612
rect 10137 16603 10195 16609
rect 7760 16544 8248 16572
rect 2685 16535 2743 16541
rect 2590 16464 2596 16516
rect 2648 16504 2654 16516
rect 2700 16504 2728 16535
rect 9122 16532 9128 16584
rect 9180 16572 9186 16584
rect 9861 16575 9919 16581
rect 9861 16572 9873 16575
rect 9180 16544 9873 16572
rect 9180 16532 9186 16544
rect 9861 16541 9873 16544
rect 9907 16541 9919 16575
rect 10244 16572 10272 16612
rect 10318 16600 10324 16652
rect 10376 16600 10382 16652
rect 10796 16640 10824 16680
rect 12710 16668 12716 16680
rect 12768 16668 12774 16720
rect 13173 16711 13231 16717
rect 13173 16677 13185 16711
rect 13219 16708 13231 16711
rect 13265 16711 13323 16717
rect 13265 16708 13277 16711
rect 13219 16680 13277 16708
rect 13219 16677 13231 16680
rect 13173 16671 13231 16677
rect 13265 16677 13277 16680
rect 13311 16677 13323 16711
rect 13265 16671 13323 16677
rect 14182 16668 14188 16720
rect 14240 16668 14246 16720
rect 14553 16711 14611 16717
rect 14553 16677 14565 16711
rect 14599 16708 14611 16711
rect 14599 16680 14964 16708
rect 14599 16677 14611 16680
rect 14553 16671 14611 16677
rect 10428 16612 10824 16640
rect 10428 16572 10456 16612
rect 11422 16600 11428 16652
rect 11480 16600 11486 16652
rect 13630 16600 13636 16652
rect 13688 16640 13694 16652
rect 14369 16643 14427 16649
rect 14369 16640 14381 16643
rect 13688 16612 14381 16640
rect 13688 16600 13694 16612
rect 14369 16609 14381 16612
rect 14415 16609 14427 16643
rect 14369 16603 14427 16609
rect 14458 16600 14464 16652
rect 14516 16600 14522 16652
rect 14734 16600 14740 16652
rect 14792 16600 14798 16652
rect 14936 16649 14964 16680
rect 15838 16668 15844 16720
rect 15896 16708 15902 16720
rect 16316 16717 16344 16748
rect 16485 16745 16497 16779
rect 16531 16776 16543 16779
rect 16777 16779 16835 16785
rect 16777 16776 16789 16779
rect 16531 16748 16789 16776
rect 16531 16745 16543 16748
rect 16485 16739 16543 16745
rect 16777 16745 16789 16748
rect 16823 16745 16835 16779
rect 16777 16739 16835 16745
rect 16942 16736 16948 16788
rect 17000 16736 17006 16788
rect 17129 16779 17187 16785
rect 17129 16745 17141 16779
rect 17175 16776 17187 16779
rect 17678 16776 17684 16788
rect 17175 16748 17684 16776
rect 17175 16745 17187 16748
rect 17129 16739 17187 16745
rect 17678 16736 17684 16748
rect 17736 16776 17742 16788
rect 18322 16776 18328 16788
rect 17736 16748 18328 16776
rect 17736 16736 17742 16748
rect 18322 16736 18328 16748
rect 18380 16736 18386 16788
rect 18693 16779 18751 16785
rect 18693 16745 18705 16779
rect 18739 16776 18751 16779
rect 18739 16748 19472 16776
rect 18739 16745 18751 16748
rect 18693 16739 18751 16745
rect 16117 16711 16175 16717
rect 16117 16708 16129 16711
rect 15896 16680 16129 16708
rect 15896 16668 15902 16680
rect 16117 16677 16129 16680
rect 16163 16677 16175 16711
rect 16117 16671 16175 16677
rect 16301 16711 16359 16717
rect 16301 16677 16313 16711
rect 16347 16677 16359 16711
rect 16301 16671 16359 16677
rect 16577 16711 16635 16717
rect 16577 16677 16589 16711
rect 16623 16708 16635 16711
rect 16666 16708 16672 16720
rect 16623 16680 16672 16708
rect 16623 16677 16635 16680
rect 16577 16671 16635 16677
rect 16666 16668 16672 16680
rect 16724 16668 16730 16720
rect 17954 16708 17960 16720
rect 17328 16680 17960 16708
rect 14921 16643 14979 16649
rect 14921 16609 14933 16643
rect 14967 16609 14979 16643
rect 14921 16603 14979 16609
rect 15013 16643 15071 16649
rect 15013 16609 15025 16643
rect 15059 16640 15071 16643
rect 15194 16640 15200 16652
rect 15059 16612 15200 16640
rect 15059 16609 15071 16612
rect 15013 16603 15071 16609
rect 15194 16600 15200 16612
rect 15252 16600 15258 16652
rect 15286 16600 15292 16652
rect 15344 16600 15350 16652
rect 15562 16600 15568 16652
rect 15620 16600 15626 16652
rect 15930 16640 15936 16652
rect 15856 16612 15936 16640
rect 10244 16544 10456 16572
rect 9861 16535 9919 16541
rect 11146 16532 11152 16584
rect 11204 16572 11210 16584
rect 11609 16575 11667 16581
rect 11609 16572 11621 16575
rect 11204 16544 11621 16572
rect 11204 16532 11210 16544
rect 11609 16541 11621 16544
rect 11655 16541 11667 16575
rect 11609 16535 11667 16541
rect 13814 16532 13820 16584
rect 13872 16532 13878 16584
rect 15102 16532 15108 16584
rect 15160 16532 15166 16584
rect 15856 16581 15884 16612
rect 15930 16600 15936 16612
rect 15988 16600 15994 16652
rect 16482 16600 16488 16652
rect 16540 16640 16546 16652
rect 17037 16643 17095 16649
rect 17037 16640 17049 16643
rect 16540 16612 17049 16640
rect 16540 16600 16546 16612
rect 17037 16609 17049 16612
rect 17083 16609 17095 16643
rect 17037 16603 17095 16609
rect 17218 16600 17224 16652
rect 17276 16600 17282 16652
rect 17328 16649 17356 16680
rect 17954 16668 17960 16680
rect 18012 16668 18018 16720
rect 17586 16649 17592 16652
rect 17313 16643 17371 16649
rect 17313 16609 17325 16643
rect 17359 16609 17371 16643
rect 17313 16603 17371 16609
rect 17580 16603 17592 16649
rect 17586 16600 17592 16603
rect 17644 16600 17650 16652
rect 19444 16649 19472 16748
rect 20346 16736 20352 16788
rect 20404 16736 20410 16788
rect 21910 16736 21916 16788
rect 21968 16736 21974 16788
rect 22002 16736 22008 16788
rect 22060 16736 22066 16788
rect 24118 16736 24124 16788
rect 24176 16736 24182 16788
rect 24670 16736 24676 16788
rect 24728 16776 24734 16788
rect 24765 16779 24823 16785
rect 24765 16776 24777 16779
rect 24728 16748 24777 16776
rect 24728 16736 24734 16748
rect 24765 16745 24777 16748
rect 24811 16745 24823 16779
rect 24765 16739 24823 16745
rect 25314 16736 25320 16788
rect 25372 16736 25378 16788
rect 25501 16779 25559 16785
rect 25501 16745 25513 16779
rect 25547 16745 25559 16779
rect 25501 16739 25559 16745
rect 20990 16668 20996 16720
rect 21048 16708 21054 16720
rect 21928 16708 21956 16736
rect 21048 16680 21772 16708
rect 21928 16680 22600 16708
rect 21048 16668 21054 16680
rect 19429 16643 19487 16649
rect 19429 16609 19441 16643
rect 19475 16640 19487 16643
rect 19794 16640 19800 16652
rect 19475 16612 19800 16640
rect 19475 16609 19487 16612
rect 19429 16603 19487 16609
rect 19794 16600 19800 16612
rect 19852 16600 19858 16652
rect 21542 16600 21548 16652
rect 21600 16640 21606 16652
rect 21744 16649 21772 16680
rect 21637 16643 21695 16649
rect 21637 16640 21649 16643
rect 21600 16612 21649 16640
rect 21600 16600 21606 16612
rect 21637 16609 21649 16612
rect 21683 16609 21695 16643
rect 21637 16603 21695 16609
rect 21729 16643 21787 16649
rect 21729 16609 21741 16643
rect 21775 16609 21787 16643
rect 21729 16603 21787 16609
rect 22189 16643 22247 16649
rect 22189 16609 22201 16643
rect 22235 16609 22247 16643
rect 22189 16603 22247 16609
rect 15841 16575 15899 16581
rect 15841 16541 15853 16575
rect 15887 16541 15899 16575
rect 15841 16535 15899 16541
rect 20254 16532 20260 16584
rect 20312 16532 20318 16584
rect 20993 16575 21051 16581
rect 20993 16541 21005 16575
rect 21039 16572 21051 16575
rect 21082 16572 21088 16584
rect 21039 16544 21088 16572
rect 21039 16541 21051 16544
rect 20993 16535 21051 16541
rect 21082 16532 21088 16544
rect 21140 16532 21146 16584
rect 21269 16575 21327 16581
rect 21269 16541 21281 16575
rect 21315 16541 21327 16575
rect 21269 16535 21327 16541
rect 21361 16575 21419 16581
rect 21361 16541 21373 16575
rect 21407 16572 21419 16575
rect 21450 16572 21456 16584
rect 21407 16544 21456 16572
rect 21407 16541 21419 16544
rect 21361 16535 21419 16541
rect 4890 16504 4896 16516
rect 2648 16476 2728 16504
rect 3988 16476 4896 16504
rect 2648 16464 2654 16476
rect 2498 16396 2504 16448
rect 2556 16436 2562 16448
rect 3988 16436 4016 16476
rect 4890 16464 4896 16476
rect 4948 16504 4954 16516
rect 21284 16504 21312 16535
rect 21450 16532 21456 16544
rect 21508 16532 21514 16584
rect 22204 16572 22232 16603
rect 22278 16600 22284 16652
rect 22336 16600 22342 16652
rect 22370 16600 22376 16652
rect 22428 16600 22434 16652
rect 22572 16649 22600 16680
rect 22922 16668 22928 16720
rect 22980 16708 22986 16720
rect 22980 16680 23244 16708
rect 22980 16668 22986 16680
rect 22557 16643 22615 16649
rect 22557 16609 22569 16643
rect 22603 16609 22615 16643
rect 22557 16603 22615 16609
rect 22741 16643 22799 16649
rect 22741 16609 22753 16643
rect 22787 16640 22799 16643
rect 22830 16640 22836 16652
rect 22787 16612 22836 16640
rect 22787 16609 22799 16612
rect 22741 16603 22799 16609
rect 22830 16600 22836 16612
rect 22888 16600 22894 16652
rect 23014 16649 23020 16652
rect 23008 16603 23020 16649
rect 23014 16600 23020 16603
rect 23072 16600 23078 16652
rect 23216 16640 23244 16680
rect 24302 16668 24308 16720
rect 24360 16708 24366 16720
rect 24578 16708 24584 16720
rect 24360 16680 24584 16708
rect 24360 16668 24366 16680
rect 24578 16668 24584 16680
rect 24636 16708 24642 16720
rect 24636 16680 24992 16708
rect 24636 16668 24642 16680
rect 23216 16612 24348 16640
rect 22646 16572 22652 16584
rect 22204 16544 22652 16572
rect 22646 16532 22652 16544
rect 22704 16532 22710 16584
rect 24320 16581 24348 16612
rect 24394 16600 24400 16652
rect 24452 16600 24458 16652
rect 24854 16600 24860 16652
rect 24912 16600 24918 16652
rect 24964 16649 24992 16680
rect 24949 16643 25007 16649
rect 24949 16609 24961 16643
rect 24995 16609 25007 16643
rect 25516 16640 25544 16739
rect 26050 16736 26056 16788
rect 26108 16736 26114 16788
rect 25869 16643 25927 16649
rect 25869 16640 25881 16643
rect 25516 16612 25881 16640
rect 24949 16603 25007 16609
rect 25869 16609 25881 16612
rect 25915 16609 25927 16643
rect 25869 16603 25927 16609
rect 24305 16575 24363 16581
rect 24305 16541 24317 16575
rect 24351 16541 24363 16575
rect 24305 16535 24363 16541
rect 21634 16504 21640 16516
rect 4948 16476 5120 16504
rect 21284 16476 21640 16504
rect 4948 16464 4954 16476
rect 2556 16408 4016 16436
rect 4065 16439 4123 16445
rect 2556 16396 2562 16408
rect 4065 16405 4077 16439
rect 4111 16436 4123 16439
rect 4154 16436 4160 16448
rect 4111 16408 4160 16436
rect 4111 16405 4123 16408
rect 4065 16399 4123 16405
rect 4154 16396 4160 16408
rect 4212 16396 4218 16448
rect 4522 16396 4528 16448
rect 4580 16396 4586 16448
rect 5092 16445 5120 16476
rect 21634 16464 21640 16476
rect 21692 16464 21698 16516
rect 5077 16439 5135 16445
rect 5077 16405 5089 16439
rect 5123 16405 5135 16439
rect 5077 16399 5135 16405
rect 9306 16396 9312 16448
rect 9364 16396 9370 16448
rect 11054 16396 11060 16448
rect 11112 16396 11118 16448
rect 12618 16396 12624 16448
rect 12676 16436 12682 16448
rect 12805 16439 12863 16445
rect 12805 16436 12817 16439
rect 12676 16408 12817 16436
rect 12676 16396 12682 16408
rect 12805 16405 12817 16408
rect 12851 16405 12863 16439
rect 12805 16399 12863 16405
rect 12989 16439 13047 16445
rect 12989 16405 13001 16439
rect 13035 16436 13047 16439
rect 13170 16436 13176 16448
rect 13035 16408 13176 16436
rect 13035 16405 13047 16408
rect 12989 16399 13047 16405
rect 13170 16396 13176 16408
rect 13228 16396 13234 16448
rect 15473 16439 15531 16445
rect 15473 16405 15485 16439
rect 15519 16436 15531 16439
rect 15657 16439 15715 16445
rect 15657 16436 15669 16439
rect 15519 16408 15669 16436
rect 15519 16405 15531 16408
rect 15473 16399 15531 16405
rect 15657 16405 15669 16408
rect 15703 16405 15715 16439
rect 15657 16399 15715 16405
rect 15746 16396 15752 16448
rect 15804 16396 15810 16448
rect 16758 16396 16764 16448
rect 16816 16396 16822 16448
rect 18782 16396 18788 16448
rect 18840 16396 18846 16448
rect 19334 16396 19340 16448
rect 19392 16436 19398 16448
rect 19613 16439 19671 16445
rect 19613 16436 19625 16439
rect 19392 16408 19625 16436
rect 19392 16396 19398 16408
rect 19613 16405 19625 16408
rect 19659 16405 19671 16439
rect 19613 16399 19671 16405
rect 24854 16396 24860 16448
rect 24912 16436 24918 16448
rect 25317 16439 25375 16445
rect 25317 16436 25329 16439
rect 24912 16408 25329 16436
rect 24912 16396 24918 16408
rect 25317 16405 25329 16408
rect 25363 16436 25375 16439
rect 25498 16436 25504 16448
rect 25363 16408 25504 16436
rect 25363 16405 25375 16408
rect 25317 16399 25375 16405
rect 25498 16396 25504 16408
rect 25556 16396 25562 16448
rect 552 16346 27416 16368
rect 552 16294 3756 16346
rect 3808 16294 3820 16346
rect 3872 16294 3884 16346
rect 3936 16294 3948 16346
rect 4000 16294 4012 16346
rect 4064 16294 10472 16346
rect 10524 16294 10536 16346
rect 10588 16294 10600 16346
rect 10652 16294 10664 16346
rect 10716 16294 10728 16346
rect 10780 16294 17188 16346
rect 17240 16294 17252 16346
rect 17304 16294 17316 16346
rect 17368 16294 17380 16346
rect 17432 16294 17444 16346
rect 17496 16294 23904 16346
rect 23956 16294 23968 16346
rect 24020 16294 24032 16346
rect 24084 16294 24096 16346
rect 24148 16294 24160 16346
rect 24212 16294 27416 16346
rect 552 16272 27416 16294
rect 1397 16235 1455 16241
rect 1397 16201 1409 16235
rect 1443 16232 1455 16235
rect 2041 16235 2099 16241
rect 2041 16232 2053 16235
rect 1443 16204 2053 16232
rect 1443 16201 1455 16204
rect 1397 16195 1455 16201
rect 2041 16201 2053 16204
rect 2087 16201 2099 16235
rect 2041 16195 2099 16201
rect 4338 16192 4344 16244
rect 4396 16192 4402 16244
rect 11054 16232 11060 16244
rect 10336 16204 11060 16232
rect 2222 16164 2228 16176
rect 1596 16136 2228 16164
rect 1596 16037 1624 16136
rect 2222 16124 2228 16136
rect 2280 16164 2286 16176
rect 2498 16164 2504 16176
rect 2280 16136 2504 16164
rect 2280 16124 2286 16136
rect 2498 16124 2504 16136
rect 2556 16124 2562 16176
rect 1854 16056 1860 16108
rect 1912 16096 1918 16108
rect 3237 16099 3295 16105
rect 3237 16096 3249 16099
rect 1912 16068 3249 16096
rect 1912 16056 1918 16068
rect 3237 16065 3249 16068
rect 3283 16065 3295 16099
rect 3237 16059 3295 16065
rect 4709 16099 4767 16105
rect 4709 16065 4721 16099
rect 4755 16096 4767 16099
rect 5810 16096 5816 16108
rect 4755 16068 5816 16096
rect 4755 16065 4767 16068
rect 4709 16059 4767 16065
rect 5810 16056 5816 16068
rect 5868 16056 5874 16108
rect 1581 16031 1639 16037
rect 1581 15997 1593 16031
rect 1627 15997 1639 16031
rect 1581 15991 1639 15997
rect 1765 16031 1823 16037
rect 1765 15997 1777 16031
rect 1811 16028 1823 16031
rect 1946 16028 1952 16040
rect 1811 16000 1952 16028
rect 1811 15997 1823 16000
rect 1765 15991 1823 15997
rect 1946 15988 1952 16000
rect 2004 16028 2010 16040
rect 2317 16031 2375 16037
rect 2317 16028 2329 16031
rect 2004 16000 2329 16028
rect 2004 15988 2010 16000
rect 2317 15997 2329 16000
rect 2363 15997 2375 16031
rect 2317 15991 2375 15997
rect 2406 15988 2412 16040
rect 2464 15988 2470 16040
rect 2498 15988 2504 16040
rect 2556 15988 2562 16040
rect 3326 15988 3332 16040
rect 3384 16028 3390 16040
rect 3789 16031 3847 16037
rect 3789 16028 3801 16031
rect 3384 16000 3801 16028
rect 3384 15988 3390 16000
rect 3789 15997 3801 16000
rect 3835 15997 3847 16031
rect 3789 15991 3847 15997
rect 4525 16031 4583 16037
rect 4525 15997 4537 16031
rect 4571 16028 4583 16031
rect 4614 16028 4620 16040
rect 4571 16000 4620 16028
rect 4571 15997 4583 16000
rect 4525 15991 4583 15997
rect 4614 15988 4620 16000
rect 4672 15988 4678 16040
rect 4798 15988 4804 16040
rect 4856 16028 4862 16040
rect 5353 16031 5411 16037
rect 5353 16028 5365 16031
rect 4856 16000 5365 16028
rect 4856 15988 4862 16000
rect 5353 15997 5365 16000
rect 5399 15997 5411 16031
rect 5353 15991 5411 15997
rect 6454 15988 6460 16040
rect 6512 16028 6518 16040
rect 7101 16031 7159 16037
rect 7101 16028 7113 16031
rect 6512 16000 7113 16028
rect 6512 15988 6518 16000
rect 7101 15997 7113 16000
rect 7147 15997 7159 16031
rect 7101 15991 7159 15997
rect 10137 16031 10195 16037
rect 10137 15997 10149 16031
rect 10183 16028 10195 16031
rect 10336 16028 10364 16204
rect 11054 16192 11060 16204
rect 11112 16192 11118 16244
rect 13170 16192 13176 16244
rect 13228 16232 13234 16244
rect 13725 16235 13783 16241
rect 13725 16232 13737 16235
rect 13228 16204 13737 16232
rect 13228 16192 13234 16204
rect 13725 16201 13737 16204
rect 13771 16201 13783 16235
rect 13725 16195 13783 16201
rect 14185 16235 14243 16241
rect 14185 16201 14197 16235
rect 14231 16232 14243 16235
rect 15102 16232 15108 16244
rect 14231 16204 15108 16232
rect 14231 16201 14243 16204
rect 14185 16195 14243 16201
rect 15102 16192 15108 16204
rect 15160 16192 15166 16244
rect 15473 16235 15531 16241
rect 15473 16201 15485 16235
rect 15519 16232 15531 16235
rect 15562 16232 15568 16244
rect 15519 16204 15568 16232
rect 15519 16201 15531 16204
rect 15473 16195 15531 16201
rect 15562 16192 15568 16204
rect 15620 16192 15626 16244
rect 17497 16235 17555 16241
rect 17497 16201 17509 16235
rect 17543 16232 17555 16235
rect 17586 16232 17592 16244
rect 17543 16204 17592 16232
rect 17543 16201 17555 16204
rect 17497 16195 17555 16201
rect 17586 16192 17592 16204
rect 17644 16192 17650 16244
rect 22189 16235 22247 16241
rect 22189 16201 22201 16235
rect 22235 16232 22247 16235
rect 22370 16232 22376 16244
rect 22235 16204 22376 16232
rect 22235 16201 22247 16204
rect 22189 16195 22247 16201
rect 22370 16192 22376 16204
rect 22428 16192 22434 16244
rect 23014 16192 23020 16244
rect 23072 16192 23078 16244
rect 22097 16167 22155 16173
rect 22097 16133 22109 16167
rect 22143 16164 22155 16167
rect 22281 16167 22339 16173
rect 22281 16164 22293 16167
rect 22143 16136 22293 16164
rect 22143 16133 22155 16136
rect 22097 16127 22155 16133
rect 22281 16133 22293 16136
rect 22327 16133 22339 16167
rect 22281 16127 22339 16133
rect 15289 16099 15347 16105
rect 15289 16065 15301 16099
rect 15335 16096 15347 16099
rect 20809 16099 20867 16105
rect 15335 16068 15700 16096
rect 15335 16065 15347 16068
rect 15289 16059 15347 16065
rect 15672 16040 15700 16068
rect 20809 16065 20821 16099
rect 20855 16096 20867 16099
rect 21450 16096 21456 16108
rect 20855 16068 21456 16096
rect 20855 16065 20867 16068
rect 20809 16059 20867 16065
rect 21450 16056 21456 16068
rect 21508 16096 21514 16108
rect 21508 16068 21588 16096
rect 21508 16056 21514 16068
rect 10183 16000 10364 16028
rect 10413 16031 10471 16037
rect 10183 15997 10195 16000
rect 10137 15991 10195 15997
rect 10413 15997 10425 16031
rect 10459 16028 10471 16031
rect 11882 16028 11888 16040
rect 10459 16000 11888 16028
rect 10459 15997 10471 16000
rect 10413 15991 10471 15997
rect 2225 15963 2283 15969
rect 2225 15929 2237 15963
rect 2271 15960 2283 15963
rect 2424 15960 2452 15988
rect 4154 15960 4160 15972
rect 2271 15932 4160 15960
rect 2271 15929 2283 15932
rect 2225 15923 2283 15929
rect 4154 15920 4160 15932
rect 4212 15920 4218 15972
rect 9674 15920 9680 15972
rect 9732 15960 9738 15972
rect 10428 15960 10456 15991
rect 11882 15988 11888 16000
rect 11940 15988 11946 16040
rect 13814 16028 13820 16040
rect 13280 16000 13820 16028
rect 10658 15963 10716 15969
rect 10658 15960 10670 15963
rect 9732 15932 10456 15960
rect 10520 15932 10670 15960
rect 9732 15920 9738 15932
rect 1486 15852 1492 15904
rect 1544 15892 1550 15904
rect 1857 15895 1915 15901
rect 1857 15892 1869 15895
rect 1544 15864 1869 15892
rect 1544 15852 1550 15864
rect 1857 15861 1869 15864
rect 1903 15861 1915 15895
rect 1857 15855 1915 15861
rect 2025 15895 2083 15901
rect 2025 15861 2037 15895
rect 2071 15892 2083 15895
rect 2409 15895 2467 15901
rect 2409 15892 2421 15895
rect 2071 15864 2421 15892
rect 2071 15861 2083 15864
rect 2025 15855 2083 15861
rect 2409 15861 2421 15864
rect 2455 15861 2467 15895
rect 2409 15855 2467 15861
rect 4614 15852 4620 15904
rect 4672 15892 4678 15904
rect 4801 15895 4859 15901
rect 4801 15892 4813 15895
rect 4672 15864 4813 15892
rect 4672 15852 4678 15864
rect 4801 15861 4813 15864
rect 4847 15861 4859 15895
rect 4801 15855 4859 15861
rect 6546 15852 6552 15904
rect 6604 15852 6610 15904
rect 10321 15895 10379 15901
rect 10321 15861 10333 15895
rect 10367 15892 10379 15895
rect 10520 15892 10548 15932
rect 10658 15929 10670 15932
rect 10704 15929 10716 15963
rect 10658 15923 10716 15929
rect 12152 15963 12210 15969
rect 12152 15929 12164 15963
rect 12198 15960 12210 15963
rect 12434 15960 12440 15972
rect 12198 15932 12440 15960
rect 12198 15929 12210 15932
rect 12152 15923 12210 15929
rect 12434 15920 12440 15932
rect 12492 15920 12498 15972
rect 10367 15864 10548 15892
rect 10367 15861 10379 15864
rect 10321 15855 10379 15861
rect 11238 15852 11244 15904
rect 11296 15892 11302 15904
rect 13280 15901 13308 16000
rect 13814 15988 13820 16000
rect 13872 16028 13878 16040
rect 14093 16031 14151 16037
rect 14093 16028 14105 16031
rect 13872 16000 14105 16028
rect 13872 15988 13878 16000
rect 14093 15997 14105 16000
rect 14139 15997 14151 16031
rect 14093 15991 14151 15997
rect 15194 15988 15200 16040
rect 15252 15988 15258 16040
rect 15473 16031 15531 16037
rect 15473 15997 15485 16031
rect 15519 15997 15531 16031
rect 15473 15991 15531 15997
rect 13722 15969 13728 15972
rect 13709 15963 13728 15969
rect 13709 15929 13721 15963
rect 13709 15923 13728 15929
rect 13722 15920 13728 15923
rect 13780 15920 13786 15972
rect 13909 15963 13967 15969
rect 13909 15929 13921 15963
rect 13955 15960 13967 15963
rect 14458 15960 14464 15972
rect 13955 15932 14464 15960
rect 13955 15929 13967 15932
rect 13909 15923 13967 15929
rect 14458 15920 14464 15932
rect 14516 15960 14522 15972
rect 15488 15960 15516 15991
rect 15654 15988 15660 16040
rect 15712 15988 15718 16040
rect 17678 15988 17684 16040
rect 17736 15988 17742 16040
rect 17862 15988 17868 16040
rect 17920 15988 17926 16040
rect 18049 16031 18107 16037
rect 18049 15997 18061 16031
rect 18095 16028 18107 16031
rect 18782 16028 18788 16040
rect 18095 16000 18788 16028
rect 18095 15997 18107 16000
rect 18049 15991 18107 15997
rect 18782 15988 18788 16000
rect 18840 15988 18846 16040
rect 19242 15988 19248 16040
rect 19300 15988 19306 16040
rect 19518 16037 19524 16040
rect 19512 16028 19524 16037
rect 19479 16000 19524 16028
rect 19512 15991 19524 16000
rect 19518 15988 19524 15991
rect 19576 15988 19582 16040
rect 19794 15988 19800 16040
rect 19852 16028 19858 16040
rect 20717 16031 20775 16037
rect 20717 16028 20729 16031
rect 19852 16000 20729 16028
rect 19852 15988 19858 16000
rect 20717 15997 20729 16000
rect 20763 15997 20775 16031
rect 20717 15991 20775 15997
rect 21082 15988 21088 16040
rect 21140 15988 21146 16040
rect 21174 15988 21180 16040
rect 21232 16028 21238 16040
rect 21560 16037 21588 16068
rect 21634 16056 21640 16108
rect 21692 16096 21698 16108
rect 21692 16068 22094 16096
rect 21692 16056 21698 16068
rect 21269 16031 21327 16037
rect 21269 16028 21281 16031
rect 21232 16000 21281 16028
rect 21232 15988 21238 16000
rect 21269 15997 21281 16000
rect 21315 15997 21327 16031
rect 21269 15991 21327 15997
rect 21361 16031 21419 16037
rect 21361 15997 21373 16031
rect 21407 15997 21419 16031
rect 21361 15991 21419 15997
rect 21545 16031 21603 16037
rect 21545 15997 21557 16031
rect 21591 15997 21603 16031
rect 21545 15991 21603 15997
rect 14516 15932 15516 15960
rect 14516 15920 14522 15932
rect 17770 15920 17776 15972
rect 17828 15920 17834 15972
rect 11793 15895 11851 15901
rect 11793 15892 11805 15895
rect 11296 15864 11805 15892
rect 11296 15852 11302 15864
rect 11793 15861 11805 15864
rect 11839 15861 11851 15895
rect 11793 15855 11851 15861
rect 13265 15895 13323 15901
rect 13265 15861 13277 15895
rect 13311 15861 13323 15895
rect 13265 15855 13323 15861
rect 13354 15852 13360 15904
rect 13412 15892 13418 15904
rect 13541 15895 13599 15901
rect 13541 15892 13553 15895
rect 13412 15864 13553 15892
rect 13412 15852 13418 15864
rect 13541 15861 13553 15864
rect 13587 15861 13599 15895
rect 13541 15855 13599 15861
rect 20625 15895 20683 15901
rect 20625 15861 20637 15895
rect 20671 15892 20683 15895
rect 21082 15892 21088 15904
rect 20671 15864 21088 15892
rect 20671 15861 20683 15864
rect 20625 15855 20683 15861
rect 21082 15852 21088 15864
rect 21140 15852 21146 15904
rect 21269 15895 21327 15901
rect 21269 15861 21281 15895
rect 21315 15892 21327 15895
rect 21376 15892 21404 15991
rect 21726 15988 21732 16040
rect 21784 15988 21790 16040
rect 21818 15988 21824 16040
rect 21876 16028 21882 16040
rect 21913 16031 21971 16037
rect 21913 16028 21925 16031
rect 21876 16000 21925 16028
rect 21876 15988 21882 16000
rect 21913 15997 21925 16000
rect 21959 15997 21971 16031
rect 22066 16028 22094 16068
rect 23566 16056 23572 16108
rect 23624 16056 23630 16108
rect 24854 16096 24860 16108
rect 24320 16068 24860 16096
rect 23845 16031 23903 16037
rect 23845 16028 23857 16031
rect 22066 16000 23857 16028
rect 21913 15991 21971 15997
rect 23845 15997 23857 16000
rect 23891 15997 23903 16031
rect 23845 15991 23903 15997
rect 24029 16031 24087 16037
rect 24029 15997 24041 16031
rect 24075 16028 24087 16031
rect 24210 16028 24216 16040
rect 24075 16000 24216 16028
rect 24075 15997 24087 16000
rect 24029 15991 24087 15997
rect 22278 15960 22284 15972
rect 22066 15932 22284 15960
rect 22066 15892 22094 15932
rect 22278 15920 22284 15932
rect 22336 15920 22342 15972
rect 22646 15920 22652 15972
rect 22704 15920 22710 15972
rect 23860 15960 23888 15991
rect 24210 15988 24216 16000
rect 24268 15988 24274 16040
rect 24320 16037 24348 16068
rect 24854 16056 24860 16068
rect 24912 16056 24918 16108
rect 24305 16031 24363 16037
rect 24305 15997 24317 16031
rect 24351 15997 24363 16031
rect 24305 15991 24363 15997
rect 24486 15988 24492 16040
rect 24544 15988 24550 16040
rect 24578 15988 24584 16040
rect 24636 15988 24642 16040
rect 24670 15988 24676 16040
rect 24728 15988 24734 16040
rect 25041 16031 25099 16037
rect 25041 15997 25053 16031
rect 25087 16028 25099 16031
rect 25682 16028 25688 16040
rect 25087 16000 25688 16028
rect 25087 15997 25099 16000
rect 25041 15991 25099 15997
rect 25682 15988 25688 16000
rect 25740 15988 25746 16040
rect 24949 15963 25007 15969
rect 23860 15932 24624 15960
rect 21315 15864 22094 15892
rect 24213 15895 24271 15901
rect 21315 15861 21327 15864
rect 21269 15855 21327 15861
rect 24213 15861 24225 15895
rect 24259 15892 24271 15895
rect 24394 15892 24400 15904
rect 24259 15864 24400 15892
rect 24259 15861 24271 15864
rect 24213 15855 24271 15861
rect 24394 15852 24400 15864
rect 24452 15852 24458 15904
rect 24596 15892 24624 15932
rect 24949 15929 24961 15963
rect 24995 15960 25007 15963
rect 25286 15963 25344 15969
rect 25286 15960 25298 15963
rect 24995 15932 25298 15960
rect 24995 15929 25007 15932
rect 24949 15923 25007 15929
rect 25286 15929 25298 15932
rect 25332 15929 25344 15963
rect 25286 15923 25344 15929
rect 26234 15892 26240 15904
rect 24596 15864 26240 15892
rect 26234 15852 26240 15864
rect 26292 15892 26298 15904
rect 26421 15895 26479 15901
rect 26421 15892 26433 15895
rect 26292 15864 26433 15892
rect 26292 15852 26298 15864
rect 26421 15861 26433 15864
rect 26467 15861 26479 15895
rect 26421 15855 26479 15861
rect 552 15802 27576 15824
rect 552 15750 7114 15802
rect 7166 15750 7178 15802
rect 7230 15750 7242 15802
rect 7294 15750 7306 15802
rect 7358 15750 7370 15802
rect 7422 15750 13830 15802
rect 13882 15750 13894 15802
rect 13946 15750 13958 15802
rect 14010 15750 14022 15802
rect 14074 15750 14086 15802
rect 14138 15750 20546 15802
rect 20598 15750 20610 15802
rect 20662 15750 20674 15802
rect 20726 15750 20738 15802
rect 20790 15750 20802 15802
rect 20854 15750 27262 15802
rect 27314 15750 27326 15802
rect 27378 15750 27390 15802
rect 27442 15750 27454 15802
rect 27506 15750 27518 15802
rect 27570 15750 27576 15802
rect 552 15728 27576 15750
rect 1765 15691 1823 15697
rect 1765 15657 1777 15691
rect 1811 15688 1823 15691
rect 1811 15660 2084 15688
rect 1811 15657 1823 15660
rect 1765 15651 1823 15657
rect 1397 15555 1455 15561
rect 1397 15521 1409 15555
rect 1443 15552 1455 15555
rect 1486 15552 1492 15564
rect 1443 15524 1492 15552
rect 1443 15521 1455 15524
rect 1397 15515 1455 15521
rect 1486 15512 1492 15524
rect 1544 15512 1550 15564
rect 1670 15512 1676 15564
rect 1728 15512 1734 15564
rect 1854 15512 1860 15564
rect 1912 15512 1918 15564
rect 2056 15552 2084 15660
rect 3326 15648 3332 15700
rect 3384 15648 3390 15700
rect 6454 15648 6460 15700
rect 6512 15648 6518 15700
rect 6549 15691 6607 15697
rect 6549 15657 6561 15691
rect 6595 15688 6607 15691
rect 7006 15688 7012 15700
rect 6595 15660 7012 15688
rect 6595 15657 6607 15660
rect 6549 15651 6607 15657
rect 7006 15648 7012 15660
rect 7064 15688 7070 15700
rect 9033 15691 9091 15697
rect 9033 15688 9045 15691
rect 7064 15660 7512 15688
rect 7064 15648 7070 15660
rect 3602 15580 3608 15632
rect 3660 15620 3666 15632
rect 3850 15623 3908 15629
rect 3850 15620 3862 15623
rect 3660 15592 3862 15620
rect 3660 15580 3666 15592
rect 3850 15589 3862 15592
rect 3896 15589 3908 15623
rect 3850 15583 3908 15589
rect 6178 15580 6184 15632
rect 6236 15620 6242 15632
rect 7484 15620 7512 15660
rect 8864 15660 9045 15688
rect 8757 15623 8815 15629
rect 8757 15620 8769 15623
rect 6236 15592 6684 15620
rect 7484 15592 8769 15620
rect 6236 15580 6242 15592
rect 2205 15555 2263 15561
rect 2205 15552 2217 15555
rect 2056 15524 2217 15552
rect 2205 15521 2217 15524
rect 2251 15521 2263 15555
rect 2205 15515 2263 15521
rect 2590 15512 2596 15564
rect 2648 15552 2654 15564
rect 2648 15524 3648 15552
rect 2648 15512 2654 15524
rect 3620 15493 3648 15524
rect 5074 15512 5080 15564
rect 5132 15552 5138 15564
rect 6656 15561 6684 15592
rect 8757 15589 8769 15592
rect 8803 15589 8815 15623
rect 8757 15583 8815 15589
rect 5261 15555 5319 15561
rect 5261 15552 5273 15555
rect 5132 15524 5273 15552
rect 5132 15512 5138 15524
rect 5261 15521 5273 15524
rect 5307 15521 5319 15555
rect 5261 15515 5319 15521
rect 6641 15555 6699 15561
rect 6641 15521 6653 15555
rect 6687 15521 6699 15555
rect 6641 15515 6699 15521
rect 6917 15555 6975 15561
rect 6917 15521 6929 15555
rect 6963 15521 6975 15555
rect 6917 15515 6975 15521
rect 7285 15555 7343 15561
rect 7285 15521 7297 15555
rect 7331 15552 7343 15555
rect 8202 15552 8208 15564
rect 7331 15524 8208 15552
rect 7331 15521 7343 15524
rect 7285 15515 7343 15521
rect 1949 15487 2007 15493
rect 1949 15484 1961 15487
rect 1412 15456 1961 15484
rect 1412 15428 1440 15456
rect 1949 15453 1961 15456
rect 1995 15453 2007 15487
rect 1949 15447 2007 15453
rect 3605 15487 3663 15493
rect 3605 15453 3617 15487
rect 3651 15453 3663 15487
rect 3605 15447 3663 15453
rect 6181 15487 6239 15493
rect 6181 15453 6193 15487
rect 6227 15484 6239 15487
rect 6270 15484 6276 15496
rect 6227 15456 6276 15484
rect 6227 15453 6239 15456
rect 6181 15447 6239 15453
rect 1394 15376 1400 15428
rect 1452 15376 1458 15428
rect 1210 15308 1216 15360
rect 1268 15308 1274 15360
rect 1964 15348 1992 15447
rect 2590 15348 2596 15360
rect 1964 15320 2596 15348
rect 2590 15308 2596 15320
rect 2648 15308 2654 15360
rect 3620 15348 3648 15447
rect 6270 15444 6276 15456
rect 6328 15444 6334 15496
rect 6825 15487 6883 15493
rect 6825 15453 6837 15487
rect 6871 15453 6883 15487
rect 6932 15484 6960 15515
rect 8202 15512 8208 15524
rect 8260 15512 8266 15564
rect 8297 15555 8355 15561
rect 8297 15521 8309 15555
rect 8343 15552 8355 15555
rect 8864 15552 8892 15660
rect 9033 15657 9045 15660
rect 9079 15657 9091 15691
rect 9033 15651 9091 15657
rect 9401 15691 9459 15697
rect 9401 15657 9413 15691
rect 9447 15688 9459 15691
rect 10318 15688 10324 15700
rect 9447 15660 10324 15688
rect 9447 15657 9459 15660
rect 9401 15651 9459 15657
rect 10318 15648 10324 15660
rect 10376 15648 10382 15700
rect 11422 15648 11428 15700
rect 11480 15688 11486 15700
rect 11609 15691 11667 15697
rect 11609 15688 11621 15691
rect 11480 15660 11621 15688
rect 11480 15648 11486 15660
rect 11609 15657 11621 15660
rect 11655 15657 11667 15691
rect 11609 15651 11667 15657
rect 12434 15648 12440 15700
rect 12492 15648 12498 15700
rect 13081 15691 13139 15697
rect 13081 15657 13093 15691
rect 13127 15688 13139 15691
rect 13127 15660 14412 15688
rect 13127 15657 13139 15660
rect 13081 15651 13139 15657
rect 8941 15623 8999 15629
rect 8941 15589 8953 15623
rect 8987 15620 8999 15623
rect 9306 15620 9312 15632
rect 8987 15592 9312 15620
rect 8987 15589 8999 15592
rect 8941 15583 8999 15589
rect 9306 15580 9312 15592
rect 9364 15580 9370 15632
rect 12805 15623 12863 15629
rect 12805 15620 12817 15623
rect 12452 15592 12817 15620
rect 12452 15564 12480 15592
rect 12805 15589 12817 15592
rect 12851 15589 12863 15623
rect 12805 15583 12863 15589
rect 13449 15623 13507 15629
rect 13449 15589 13461 15623
rect 13495 15620 13507 15623
rect 13786 15623 13844 15629
rect 13786 15620 13798 15623
rect 13495 15592 13798 15620
rect 13495 15589 13507 15592
rect 13449 15583 13507 15589
rect 13786 15589 13798 15592
rect 13832 15589 13844 15623
rect 14384 15620 14412 15660
rect 14458 15648 14464 15700
rect 14516 15688 14522 15700
rect 14921 15691 14979 15697
rect 14921 15688 14933 15691
rect 14516 15660 14933 15688
rect 14516 15648 14522 15660
rect 14921 15657 14933 15660
rect 14967 15657 14979 15691
rect 14921 15651 14979 15657
rect 17678 15648 17684 15700
rect 17736 15688 17742 15700
rect 19153 15691 19211 15697
rect 17736 15660 18920 15688
rect 17736 15648 17742 15660
rect 16574 15620 16580 15632
rect 14384 15592 16580 15620
rect 13786 15583 13844 15589
rect 16574 15580 16580 15592
rect 16632 15580 16638 15632
rect 17497 15623 17555 15629
rect 17497 15620 17509 15623
rect 16868 15592 17509 15620
rect 16868 15564 16896 15592
rect 17497 15589 17509 15592
rect 17543 15589 17555 15623
rect 17497 15583 17555 15589
rect 17862 15580 17868 15632
rect 17920 15620 17926 15632
rect 18785 15623 18843 15629
rect 18785 15620 18797 15623
rect 17920 15592 18797 15620
rect 17920 15580 17926 15592
rect 18785 15589 18797 15592
rect 18831 15589 18843 15623
rect 18892 15620 18920 15660
rect 19153 15657 19165 15691
rect 19199 15657 19211 15691
rect 19153 15651 19211 15657
rect 19168 15620 19196 15651
rect 20254 15648 20260 15700
rect 20312 15688 20318 15700
rect 20625 15691 20683 15697
rect 20625 15688 20637 15691
rect 20312 15660 20637 15688
rect 20312 15648 20318 15660
rect 20625 15657 20637 15660
rect 20671 15657 20683 15691
rect 20625 15651 20683 15657
rect 19490 15623 19548 15629
rect 19490 15620 19502 15623
rect 18892 15592 19012 15620
rect 19168 15592 19502 15620
rect 18785 15583 18843 15589
rect 11238 15552 11244 15564
rect 8343 15524 8892 15552
rect 9140 15524 11244 15552
rect 8343 15521 8355 15524
rect 8297 15515 8355 15521
rect 9140 15496 9168 15524
rect 11238 15512 11244 15524
rect 11296 15512 11302 15564
rect 11425 15555 11483 15561
rect 11425 15521 11437 15555
rect 11471 15521 11483 15555
rect 11425 15515 11483 15521
rect 9122 15484 9128 15496
rect 6932 15456 9128 15484
rect 6825 15447 6883 15453
rect 6840 15416 6868 15447
rect 9122 15444 9128 15456
rect 9180 15444 9186 15496
rect 9214 15444 9220 15496
rect 9272 15484 9278 15496
rect 9493 15487 9551 15493
rect 9493 15484 9505 15487
rect 9272 15456 9505 15484
rect 9272 15444 9278 15456
rect 9493 15453 9505 15456
rect 9539 15453 9551 15487
rect 9493 15447 9551 15453
rect 9585 15487 9643 15493
rect 9585 15453 9597 15487
rect 9631 15484 9643 15487
rect 11330 15484 11336 15496
rect 9631 15456 11336 15484
rect 9631 15453 9643 15456
rect 9585 15447 9643 15453
rect 9600 15416 9628 15447
rect 11330 15444 11336 15456
rect 11388 15444 11394 15496
rect 11440 15484 11468 15515
rect 12434 15512 12440 15564
rect 12492 15512 12498 15564
rect 12618 15512 12624 15564
rect 12676 15512 12682 15564
rect 12897 15555 12955 15561
rect 12897 15521 12909 15555
rect 12943 15552 12955 15555
rect 12986 15552 12992 15564
rect 12943 15524 12992 15552
rect 12943 15521 12955 15524
rect 12897 15515 12955 15521
rect 12986 15512 12992 15524
rect 13044 15512 13050 15564
rect 13265 15555 13323 15561
rect 13265 15521 13277 15555
rect 13311 15552 13323 15555
rect 13354 15552 13360 15564
rect 13311 15524 13360 15552
rect 13311 15521 13323 15524
rect 13265 15515 13323 15521
rect 13354 15512 13360 15524
rect 13412 15512 13418 15564
rect 13538 15512 13544 15564
rect 13596 15512 13602 15564
rect 13648 15524 15516 15552
rect 11514 15484 11520 15496
rect 11440 15456 11520 15484
rect 11514 15444 11520 15456
rect 11572 15484 11578 15496
rect 13648 15484 13676 15524
rect 11572 15456 13676 15484
rect 11572 15444 11578 15456
rect 15194 15444 15200 15496
rect 15252 15484 15258 15496
rect 15381 15487 15439 15493
rect 15381 15484 15393 15487
rect 15252 15456 15393 15484
rect 15252 15444 15258 15456
rect 15381 15453 15393 15456
rect 15427 15453 15439 15487
rect 15488 15484 15516 15524
rect 15562 15512 15568 15564
rect 15620 15512 15626 15564
rect 16850 15512 16856 15564
rect 16908 15512 16914 15564
rect 17034 15512 17040 15564
rect 17092 15552 17098 15564
rect 17129 15555 17187 15561
rect 17129 15552 17141 15555
rect 17092 15524 17141 15552
rect 17092 15512 17098 15524
rect 17129 15521 17141 15524
rect 17175 15552 17187 15555
rect 17313 15555 17371 15561
rect 17313 15552 17325 15555
rect 17175 15524 17325 15552
rect 17175 15521 17187 15524
rect 17129 15515 17187 15521
rect 17313 15521 17325 15524
rect 17359 15521 17371 15555
rect 17313 15515 17371 15521
rect 18601 15555 18659 15561
rect 18601 15521 18613 15555
rect 18647 15521 18659 15555
rect 18601 15515 18659 15521
rect 17954 15484 17960 15496
rect 15488 15456 17960 15484
rect 15381 15447 15439 15453
rect 17954 15444 17960 15456
rect 18012 15444 18018 15496
rect 18616 15484 18644 15515
rect 18690 15512 18696 15564
rect 18748 15552 18754 15564
rect 18984 15561 19012 15592
rect 19490 15589 19502 15592
rect 19536 15589 19548 15623
rect 20640 15620 20668 15651
rect 22002 15648 22008 15700
rect 22060 15688 22066 15700
rect 22646 15688 22652 15700
rect 22060 15660 22652 15688
rect 22060 15648 22066 15660
rect 22646 15648 22652 15660
rect 22704 15648 22710 15700
rect 23017 15691 23075 15697
rect 23017 15657 23029 15691
rect 23063 15688 23075 15691
rect 23198 15688 23204 15700
rect 23063 15660 23204 15688
rect 23063 15657 23075 15660
rect 23017 15651 23075 15657
rect 23198 15648 23204 15660
rect 23256 15688 23262 15700
rect 24213 15691 24271 15697
rect 24213 15688 24225 15691
rect 23256 15660 24225 15688
rect 23256 15648 23262 15660
rect 24213 15657 24225 15660
rect 24259 15657 24271 15691
rect 24213 15651 24271 15657
rect 24486 15648 24492 15700
rect 24544 15688 24550 15700
rect 24673 15691 24731 15697
rect 24673 15688 24685 15691
rect 24544 15660 24685 15688
rect 24544 15648 24550 15660
rect 24673 15657 24685 15660
rect 24719 15657 24731 15691
rect 24673 15651 24731 15657
rect 20640 15592 21680 15620
rect 19490 15583 19548 15589
rect 18877 15555 18935 15561
rect 18877 15552 18889 15555
rect 18748 15524 18889 15552
rect 18748 15512 18754 15524
rect 18877 15521 18889 15524
rect 18923 15521 18935 15555
rect 18877 15515 18935 15521
rect 18969 15555 19027 15561
rect 18969 15521 18981 15555
rect 19015 15521 19027 15555
rect 18969 15515 19027 15521
rect 19242 15512 19248 15564
rect 19300 15512 19306 15564
rect 19334 15512 19340 15564
rect 19392 15512 19398 15564
rect 21082 15512 21088 15564
rect 21140 15552 21146 15564
rect 21545 15555 21603 15561
rect 21545 15552 21557 15555
rect 21140 15524 21557 15552
rect 21140 15512 21146 15524
rect 21545 15521 21557 15524
rect 21591 15521 21603 15555
rect 21652 15552 21680 15592
rect 21818 15580 21824 15632
rect 21876 15580 21882 15632
rect 22094 15580 22100 15632
rect 22152 15580 22158 15632
rect 22738 15580 22744 15632
rect 22796 15620 22802 15632
rect 22925 15623 22983 15629
rect 22925 15620 22937 15623
rect 22796 15592 22937 15620
rect 22796 15580 22802 15592
rect 22925 15589 22937 15592
rect 22971 15589 22983 15623
rect 22925 15583 22983 15589
rect 22005 15555 22063 15561
rect 22005 15553 22017 15555
rect 21928 15552 22017 15553
rect 21652 15525 22017 15552
rect 21652 15524 21956 15525
rect 21545 15515 21603 15521
rect 22005 15521 22017 15525
rect 22051 15521 22063 15555
rect 22005 15515 22063 15521
rect 22462 15512 22468 15564
rect 22520 15552 22526 15564
rect 22833 15555 22891 15561
rect 22833 15552 22845 15555
rect 22520 15524 22845 15552
rect 22520 15512 22526 15524
rect 22833 15521 22845 15524
rect 22879 15521 22891 15555
rect 22833 15515 22891 15521
rect 23293 15555 23351 15561
rect 23293 15521 23305 15555
rect 23339 15552 23351 15555
rect 24121 15555 24179 15561
rect 24121 15552 24133 15555
rect 23339 15524 24133 15552
rect 23339 15521 23351 15524
rect 23293 15515 23351 15521
rect 24121 15521 24133 15524
rect 24167 15552 24179 15555
rect 24213 15555 24271 15561
rect 24213 15552 24225 15555
rect 24167 15524 24225 15552
rect 24167 15521 24179 15524
rect 24121 15515 24179 15521
rect 24213 15521 24225 15524
rect 24259 15521 24271 15555
rect 24213 15515 24271 15521
rect 24394 15512 24400 15564
rect 24452 15512 24458 15564
rect 24578 15512 24584 15564
rect 24636 15512 24642 15564
rect 24670 15512 24676 15564
rect 24728 15552 24734 15564
rect 24765 15555 24823 15561
rect 24765 15552 24777 15555
rect 24728 15524 24777 15552
rect 24728 15512 24734 15524
rect 24765 15521 24777 15524
rect 24811 15521 24823 15555
rect 24765 15515 24823 15521
rect 19352 15484 19380 15512
rect 18616 15456 19380 15484
rect 21174 15444 21180 15496
rect 21232 15484 21238 15496
rect 21453 15487 21511 15493
rect 21453 15484 21465 15487
rect 21232 15456 21465 15484
rect 21232 15444 21238 15456
rect 21453 15453 21465 15456
rect 21499 15453 21511 15487
rect 21453 15447 21511 15453
rect 5000 15388 6868 15416
rect 6932 15388 9628 15416
rect 17129 15419 17187 15425
rect 4522 15348 4528 15360
rect 3620 15320 4528 15348
rect 4522 15308 4528 15320
rect 4580 15308 4586 15360
rect 4798 15308 4804 15360
rect 4856 15348 4862 15360
rect 5000 15357 5028 15388
rect 4985 15351 5043 15357
rect 4985 15348 4997 15351
rect 4856 15320 4997 15348
rect 4856 15308 4862 15320
rect 4985 15317 4997 15320
rect 5031 15317 5043 15351
rect 4985 15311 5043 15317
rect 5077 15351 5135 15357
rect 5077 15317 5089 15351
rect 5123 15348 5135 15351
rect 5166 15348 5172 15360
rect 5123 15320 5172 15348
rect 5123 15317 5135 15320
rect 5077 15311 5135 15317
rect 5166 15308 5172 15320
rect 5224 15308 5230 15360
rect 5810 15308 5816 15360
rect 5868 15348 5874 15360
rect 6270 15348 6276 15360
rect 5868 15320 6276 15348
rect 5868 15308 5874 15320
rect 6270 15308 6276 15320
rect 6328 15348 6334 15360
rect 6932 15348 6960 15388
rect 17129 15385 17141 15419
rect 17175 15416 17187 15419
rect 17586 15416 17592 15428
rect 17175 15388 17592 15416
rect 17175 15385 17187 15388
rect 17129 15379 17187 15385
rect 17586 15376 17592 15388
rect 17644 15376 17650 15428
rect 21468 15416 21496 15447
rect 21726 15444 21732 15496
rect 21784 15484 21790 15496
rect 21913 15487 21971 15493
rect 21913 15484 21925 15487
rect 21784 15456 21925 15484
rect 21784 15444 21790 15456
rect 21913 15453 21925 15456
rect 21959 15453 21971 15487
rect 21913 15447 21971 15453
rect 23569 15487 23627 15493
rect 23569 15453 23581 15487
rect 23615 15484 23627 15487
rect 23658 15484 23664 15496
rect 23615 15456 23664 15484
rect 23615 15453 23627 15456
rect 23569 15447 23627 15453
rect 23658 15444 23664 15456
rect 23716 15444 23722 15496
rect 22922 15416 22928 15428
rect 21468 15388 22928 15416
rect 22922 15376 22928 15388
rect 22980 15376 22986 15428
rect 23201 15419 23259 15425
rect 23201 15385 23213 15419
rect 23247 15416 23259 15419
rect 24412 15416 24440 15512
rect 24780 15484 24808 15515
rect 24946 15512 24952 15564
rect 25004 15552 25010 15564
rect 25133 15555 25191 15561
rect 25133 15552 25145 15555
rect 25004 15524 25145 15552
rect 25004 15512 25010 15524
rect 25133 15521 25145 15524
rect 25179 15521 25191 15555
rect 25133 15515 25191 15521
rect 25317 15555 25375 15561
rect 25317 15521 25329 15555
rect 25363 15552 25375 15555
rect 26602 15552 26608 15564
rect 25363 15524 26608 15552
rect 25363 15521 25375 15524
rect 25317 15515 25375 15521
rect 26602 15512 26608 15524
rect 26660 15512 26666 15564
rect 25593 15487 25651 15493
rect 25593 15484 25605 15487
rect 24780 15456 25605 15484
rect 25593 15453 25605 15456
rect 25639 15453 25651 15487
rect 25593 15447 25651 15453
rect 26234 15444 26240 15496
rect 26292 15444 26298 15496
rect 26970 15444 26976 15496
rect 27028 15444 27034 15496
rect 23247 15388 24440 15416
rect 25501 15419 25559 15425
rect 23247 15385 23259 15388
rect 23201 15379 23259 15385
rect 25501 15385 25513 15419
rect 25547 15416 25559 15419
rect 26786 15416 26792 15428
rect 25547 15388 26792 15416
rect 25547 15385 25559 15388
rect 25501 15379 25559 15385
rect 26786 15376 26792 15388
rect 26844 15376 26850 15428
rect 6328 15320 6960 15348
rect 6328 15308 6334 15320
rect 7190 15308 7196 15360
rect 7248 15308 7254 15360
rect 7469 15351 7527 15357
rect 7469 15317 7481 15351
rect 7515 15348 7527 15351
rect 7742 15348 7748 15360
rect 7515 15320 7748 15348
rect 7515 15317 7527 15320
rect 7469 15311 7527 15317
rect 7742 15308 7748 15320
rect 7800 15308 7806 15360
rect 8478 15308 8484 15360
rect 8536 15308 8542 15360
rect 8573 15351 8631 15357
rect 8573 15317 8585 15351
rect 8619 15348 8631 15351
rect 8754 15348 8760 15360
rect 8619 15320 8760 15348
rect 8619 15317 8631 15320
rect 8573 15311 8631 15317
rect 8754 15308 8760 15320
rect 8812 15308 8818 15360
rect 15749 15351 15807 15357
rect 15749 15317 15761 15351
rect 15795 15348 15807 15351
rect 16666 15348 16672 15360
rect 15795 15320 16672 15348
rect 15795 15317 15807 15320
rect 15749 15311 15807 15317
rect 16666 15308 16672 15320
rect 16724 15348 16730 15360
rect 17034 15348 17040 15360
rect 16724 15320 17040 15348
rect 16724 15308 16730 15320
rect 17034 15308 17040 15320
rect 17092 15308 17098 15360
rect 17681 15351 17739 15357
rect 17681 15317 17693 15351
rect 17727 15348 17739 15351
rect 18874 15348 18880 15360
rect 17727 15320 18880 15348
rect 17727 15317 17739 15320
rect 17681 15311 17739 15317
rect 18874 15308 18880 15320
rect 18932 15308 18938 15360
rect 21269 15351 21327 15357
rect 21269 15317 21281 15351
rect 21315 15348 21327 15351
rect 22002 15348 22008 15360
rect 21315 15320 22008 15348
rect 21315 15317 21327 15320
rect 21269 15311 21327 15317
rect 22002 15308 22008 15320
rect 22060 15308 22066 15360
rect 22554 15308 22560 15360
rect 22612 15308 22618 15360
rect 26421 15351 26479 15357
rect 26421 15317 26433 15351
rect 26467 15348 26479 15351
rect 26694 15348 26700 15360
rect 26467 15320 26700 15348
rect 26467 15317 26479 15320
rect 26421 15311 26479 15317
rect 26694 15308 26700 15320
rect 26752 15308 26758 15360
rect 552 15258 27416 15280
rect 552 15206 3756 15258
rect 3808 15206 3820 15258
rect 3872 15206 3884 15258
rect 3936 15206 3948 15258
rect 4000 15206 4012 15258
rect 4064 15206 10472 15258
rect 10524 15206 10536 15258
rect 10588 15206 10600 15258
rect 10652 15206 10664 15258
rect 10716 15206 10728 15258
rect 10780 15206 17188 15258
rect 17240 15206 17252 15258
rect 17304 15206 17316 15258
rect 17368 15206 17380 15258
rect 17432 15206 17444 15258
rect 17496 15206 23904 15258
rect 23956 15206 23968 15258
rect 24020 15206 24032 15258
rect 24084 15206 24096 15258
rect 24148 15206 24160 15258
rect 24212 15206 27416 15258
rect 552 15184 27416 15206
rect 2225 15147 2283 15153
rect 2225 15113 2237 15147
rect 2271 15144 2283 15147
rect 2498 15144 2504 15156
rect 2271 15116 2504 15144
rect 2271 15113 2283 15116
rect 2225 15107 2283 15113
rect 2498 15104 2504 15116
rect 2556 15104 2562 15156
rect 3602 15104 3608 15156
rect 3660 15144 3666 15156
rect 4065 15147 4123 15153
rect 4065 15144 4077 15147
rect 3660 15116 4077 15144
rect 3660 15104 3666 15116
rect 4065 15113 4077 15116
rect 4111 15113 4123 15147
rect 4065 15107 4123 15113
rect 6181 15147 6239 15153
rect 6181 15113 6193 15147
rect 6227 15144 6239 15147
rect 6914 15144 6920 15156
rect 6227 15116 6920 15144
rect 6227 15113 6239 15116
rect 6181 15107 6239 15113
rect 6914 15104 6920 15116
rect 6972 15144 6978 15156
rect 7190 15144 7196 15156
rect 6972 15116 7196 15144
rect 6972 15104 6978 15116
rect 7190 15104 7196 15116
rect 7248 15104 7254 15156
rect 8110 15104 8116 15156
rect 8168 15144 8174 15156
rect 12897 15147 12955 15153
rect 8168 15116 12434 15144
rect 8168 15104 8174 15116
rect 11241 15079 11299 15085
rect 11241 15045 11253 15079
rect 11287 15076 11299 15079
rect 12406 15076 12434 15116
rect 12897 15113 12909 15147
rect 12943 15144 12955 15147
rect 12986 15144 12992 15156
rect 12943 15116 12992 15144
rect 12943 15113 12955 15116
rect 12897 15107 12955 15113
rect 12986 15104 12992 15116
rect 13044 15104 13050 15156
rect 21818 15104 21824 15156
rect 21876 15144 21882 15156
rect 23658 15144 23664 15156
rect 21876 15116 23664 15144
rect 21876 15104 21882 15116
rect 23658 15104 23664 15116
rect 23716 15104 23722 15156
rect 26326 15104 26332 15156
rect 26384 15144 26390 15156
rect 26970 15144 26976 15156
rect 26384 15116 26976 15144
rect 26384 15104 26390 15116
rect 26970 15104 26976 15116
rect 27028 15144 27034 15156
rect 27065 15147 27123 15153
rect 27065 15144 27077 15147
rect 27028 15116 27077 15144
rect 27028 15104 27034 15116
rect 27065 15113 27077 15116
rect 27111 15113 27123 15147
rect 27065 15107 27123 15113
rect 14826 15076 14832 15088
rect 11287 15048 11376 15076
rect 12406 15048 14832 15076
rect 11287 15045 11299 15048
rect 11241 15039 11299 15045
rect 4154 14968 4160 15020
rect 4212 15008 4218 15020
rect 4212 14980 4384 15008
rect 4212 14968 4218 14980
rect 845 14943 903 14949
rect 845 14909 857 14943
rect 891 14940 903 14943
rect 1394 14940 1400 14952
rect 891 14912 1400 14940
rect 891 14909 903 14912
rect 845 14903 903 14909
rect 1394 14900 1400 14912
rect 1452 14900 1458 14952
rect 4356 14949 4384 14980
rect 4614 14968 4620 15020
rect 4672 14968 4678 15020
rect 4706 14968 4712 15020
rect 4764 14968 4770 15020
rect 11348 15017 11376 15048
rect 14826 15036 14832 15048
rect 14884 15036 14890 15088
rect 11333 15011 11391 15017
rect 11333 14977 11345 15011
rect 11379 14977 11391 15011
rect 12342 15008 12348 15020
rect 11333 14971 11391 14977
rect 12268 14980 12348 15008
rect 4249 14943 4307 14949
rect 4249 14909 4261 14943
rect 4295 14909 4307 14943
rect 4249 14903 4307 14909
rect 4341 14943 4399 14949
rect 4341 14909 4353 14943
rect 4387 14909 4399 14943
rect 4341 14903 4399 14909
rect 1112 14875 1170 14881
rect 1112 14841 1124 14875
rect 1158 14872 1170 14875
rect 1210 14872 1216 14884
rect 1158 14844 1216 14872
rect 1158 14841 1170 14844
rect 1112 14835 1170 14841
rect 1210 14832 1216 14844
rect 1268 14832 1274 14884
rect 4264 14804 4292 14903
rect 4522 14900 4528 14952
rect 4580 14940 4586 14952
rect 4801 14943 4859 14949
rect 4801 14940 4813 14943
rect 4580 14912 4813 14940
rect 4580 14900 4586 14912
rect 4801 14909 4813 14912
rect 4847 14940 4859 14943
rect 6086 14940 6092 14952
rect 4847 14912 6092 14940
rect 4847 14909 4859 14912
rect 4801 14903 4859 14909
rect 6086 14900 6092 14912
rect 6144 14940 6150 14952
rect 6546 14949 6552 14952
rect 6273 14943 6331 14949
rect 6273 14940 6285 14943
rect 6144 14912 6285 14940
rect 6144 14900 6150 14912
rect 6273 14909 6285 14912
rect 6319 14909 6331 14943
rect 6540 14940 6552 14949
rect 6507 14912 6552 14940
rect 6273 14903 6331 14909
rect 6540 14903 6552 14912
rect 6546 14900 6552 14903
rect 6604 14900 6610 14952
rect 7742 14900 7748 14952
rect 7800 14900 7806 14952
rect 7926 14900 7932 14952
rect 7984 14900 7990 14952
rect 8386 14900 8392 14952
rect 8444 14940 8450 14952
rect 9582 14940 9588 14952
rect 8444 14912 9588 14940
rect 8444 14900 8450 14912
rect 9582 14900 9588 14912
rect 9640 14940 9646 14952
rect 9861 14943 9919 14949
rect 9861 14940 9873 14943
rect 9640 14912 9873 14940
rect 9640 14900 9646 14912
rect 9861 14909 9873 14912
rect 9907 14909 9919 14943
rect 9861 14903 9919 14909
rect 10128 14943 10186 14949
rect 10128 14909 10140 14943
rect 10174 14940 10186 14943
rect 11146 14940 11152 14952
rect 10174 14912 11152 14940
rect 10174 14909 10186 14912
rect 10128 14903 10186 14909
rect 11146 14900 11152 14912
rect 11204 14900 11210 14952
rect 12268 14949 12296 14980
rect 12342 14968 12348 14980
rect 12400 15008 12406 15020
rect 13630 15008 13636 15020
rect 12400 14980 12756 15008
rect 12400 14968 12406 14980
rect 12253 14943 12311 14949
rect 12253 14909 12265 14943
rect 12299 14909 12311 14943
rect 12253 14903 12311 14909
rect 12529 14943 12587 14949
rect 12529 14909 12541 14943
rect 12575 14909 12587 14943
rect 12529 14903 12587 14909
rect 5068 14875 5126 14881
rect 5068 14872 5080 14875
rect 4816 14844 5080 14872
rect 4816 14804 4844 14844
rect 5068 14841 5080 14844
rect 5114 14872 5126 14875
rect 5166 14872 5172 14884
rect 5114 14844 5172 14872
rect 5114 14841 5126 14844
rect 5068 14835 5126 14841
rect 5166 14832 5172 14844
rect 5224 14832 5230 14884
rect 6178 14832 6184 14884
rect 6236 14872 6242 14884
rect 7837 14875 7895 14881
rect 7837 14872 7849 14875
rect 6236 14844 7849 14872
rect 6236 14832 6242 14844
rect 7837 14841 7849 14844
rect 7883 14841 7895 14875
rect 7837 14835 7895 14841
rect 8478 14832 8484 14884
rect 8536 14872 8542 14884
rect 8634 14875 8692 14881
rect 8634 14872 8646 14875
rect 8536 14844 8646 14872
rect 8536 14832 8542 14844
rect 8634 14841 8646 14844
rect 8680 14841 8692 14875
rect 8634 14835 8692 14841
rect 12158 14832 12164 14884
rect 12216 14872 12222 14884
rect 12437 14875 12495 14881
rect 12437 14872 12449 14875
rect 12216 14844 12449 14872
rect 12216 14832 12222 14844
rect 12437 14841 12449 14844
rect 12483 14872 12495 14875
rect 12544 14872 12572 14903
rect 12618 14900 12624 14952
rect 12676 14900 12682 14952
rect 12728 14949 12756 14980
rect 12912 14980 13636 15008
rect 12912 14949 12940 14980
rect 13630 14968 13636 14980
rect 13688 14968 13694 15020
rect 21910 15008 21916 15020
rect 17144 14980 21916 15008
rect 12713 14943 12771 14949
rect 12713 14909 12725 14943
rect 12759 14909 12771 14943
rect 12713 14903 12771 14909
rect 12897 14943 12955 14949
rect 12897 14909 12909 14943
rect 12943 14909 12955 14943
rect 12897 14903 12955 14909
rect 13081 14943 13139 14949
rect 13081 14909 13093 14943
rect 13127 14940 13139 14943
rect 14182 14940 14188 14952
rect 13127 14912 14188 14940
rect 13127 14909 13139 14912
rect 13081 14903 13139 14909
rect 14182 14900 14188 14912
rect 14240 14900 14246 14952
rect 14274 14900 14280 14952
rect 14332 14940 14338 14952
rect 15657 14943 15715 14949
rect 15657 14940 15669 14943
rect 14332 14912 15669 14940
rect 14332 14900 14338 14912
rect 15657 14909 15669 14912
rect 15703 14909 15715 14943
rect 16206 14940 16212 14952
rect 15657 14903 15715 14909
rect 15856 14912 16212 14940
rect 12483 14844 12572 14872
rect 12636 14844 12940 14872
rect 12483 14841 12495 14844
rect 12437 14835 12495 14841
rect 4264 14776 4844 14804
rect 7653 14807 7711 14813
rect 7653 14773 7665 14807
rect 7699 14804 7711 14807
rect 7742 14804 7748 14816
rect 7699 14776 7748 14804
rect 7699 14773 7711 14776
rect 7653 14767 7711 14773
rect 7742 14764 7748 14776
rect 7800 14764 7806 14816
rect 9582 14764 9588 14816
rect 9640 14804 9646 14816
rect 9769 14807 9827 14813
rect 9769 14804 9781 14807
rect 9640 14776 9781 14804
rect 9640 14764 9646 14776
rect 9769 14773 9781 14776
rect 9815 14773 9827 14807
rect 9769 14767 9827 14773
rect 11698 14764 11704 14816
rect 11756 14804 11762 14816
rect 11977 14807 12035 14813
rect 11977 14804 11989 14807
rect 11756 14776 11989 14804
rect 11756 14764 11762 14776
rect 11977 14773 11989 14776
rect 12023 14773 12035 14807
rect 11977 14767 12035 14773
rect 12069 14807 12127 14813
rect 12069 14773 12081 14807
rect 12115 14804 12127 14807
rect 12636 14804 12664 14844
rect 12912 14816 12940 14844
rect 13538 14832 13544 14884
rect 13596 14872 13602 14884
rect 14292 14872 14320 14900
rect 13596 14844 14320 14872
rect 13596 14832 13602 14844
rect 14826 14832 14832 14884
rect 14884 14872 14890 14884
rect 15105 14875 15163 14881
rect 15105 14872 15117 14875
rect 14884 14844 15117 14872
rect 14884 14832 14890 14844
rect 15105 14841 15117 14844
rect 15151 14872 15163 14875
rect 15194 14872 15200 14884
rect 15151 14844 15200 14872
rect 15151 14841 15163 14844
rect 15105 14835 15163 14841
rect 15194 14832 15200 14844
rect 15252 14832 15258 14884
rect 15289 14875 15347 14881
rect 15289 14841 15301 14875
rect 15335 14872 15347 14875
rect 15856 14872 15884 14912
rect 16206 14900 16212 14912
rect 16264 14940 16270 14952
rect 17144 14940 17172 14980
rect 21910 14968 21916 14980
rect 21968 14968 21974 15020
rect 24857 15011 24915 15017
rect 24857 14977 24869 15011
rect 24903 15008 24915 15011
rect 25038 15008 25044 15020
rect 24903 14980 25044 15008
rect 24903 14977 24915 14980
rect 24857 14971 24915 14977
rect 25038 14968 25044 14980
rect 25096 14968 25102 15020
rect 25682 14968 25688 15020
rect 25740 14968 25746 15020
rect 16264 14912 17172 14940
rect 17221 14943 17279 14949
rect 16264 14900 16270 14912
rect 17221 14909 17233 14943
rect 17267 14940 17279 14943
rect 17865 14943 17923 14949
rect 17865 14940 17877 14943
rect 17267 14912 17877 14940
rect 17267 14909 17279 14912
rect 17221 14903 17279 14909
rect 17865 14909 17877 14912
rect 17911 14909 17923 14943
rect 17865 14903 17923 14909
rect 15335 14844 15884 14872
rect 15924 14875 15982 14881
rect 15335 14841 15347 14844
rect 15289 14835 15347 14841
rect 15924 14841 15936 14875
rect 15970 14872 15982 14875
rect 16850 14872 16856 14884
rect 15970 14844 16856 14872
rect 15970 14841 15982 14844
rect 15924 14835 15982 14841
rect 16850 14832 16856 14844
rect 16908 14832 16914 14884
rect 12115 14776 12664 14804
rect 12115 14773 12127 14776
rect 12069 14767 12127 14773
rect 12894 14764 12900 14816
rect 12952 14764 12958 14816
rect 17037 14807 17095 14813
rect 17037 14773 17049 14807
rect 17083 14804 17095 14807
rect 17236 14804 17264 14903
rect 17880 14872 17908 14903
rect 17954 14900 17960 14952
rect 18012 14940 18018 14952
rect 18049 14943 18107 14949
rect 18049 14940 18061 14943
rect 18012 14912 18061 14940
rect 18012 14900 18018 14912
rect 18049 14909 18061 14912
rect 18095 14909 18107 14943
rect 18049 14903 18107 14909
rect 18233 14943 18291 14949
rect 18233 14909 18245 14943
rect 18279 14940 18291 14943
rect 18325 14943 18383 14949
rect 18325 14940 18337 14943
rect 18279 14912 18337 14940
rect 18279 14909 18291 14912
rect 18233 14903 18291 14909
rect 18325 14909 18337 14912
rect 18371 14909 18383 14943
rect 18325 14903 18383 14909
rect 22094 14900 22100 14952
rect 22152 14940 22158 14952
rect 22281 14943 22339 14949
rect 22281 14940 22293 14943
rect 22152 14912 22293 14940
rect 22152 14900 22158 14912
rect 22281 14909 22293 14912
rect 22327 14940 22339 14943
rect 22830 14940 22836 14952
rect 22327 14912 22836 14940
rect 22327 14909 22339 14912
rect 22281 14903 22339 14909
rect 22830 14900 22836 14912
rect 22888 14900 22894 14952
rect 25133 14943 25191 14949
rect 25133 14940 25145 14943
rect 24872 14912 25145 14940
rect 21082 14872 21088 14884
rect 17880 14844 21088 14872
rect 21082 14832 21088 14844
rect 21140 14832 21146 14884
rect 22554 14881 22560 14884
rect 22548 14872 22560 14881
rect 22515 14844 22560 14872
rect 22548 14835 22560 14844
rect 22554 14832 22560 14835
rect 22612 14832 22618 14884
rect 23290 14832 23296 14884
rect 23348 14872 23354 14884
rect 24213 14875 24271 14881
rect 24213 14872 24225 14875
rect 23348 14844 24225 14872
rect 23348 14832 23354 14844
rect 24213 14841 24225 14844
rect 24259 14872 24271 14875
rect 24872 14872 24900 14912
rect 25133 14909 25145 14912
rect 25179 14909 25191 14943
rect 25133 14903 25191 14909
rect 24259 14844 24900 14872
rect 24259 14841 24271 14844
rect 24213 14835 24271 14841
rect 24946 14832 24952 14884
rect 25004 14832 25010 14884
rect 25952 14875 26010 14881
rect 25952 14841 25964 14875
rect 25998 14872 26010 14875
rect 26418 14872 26424 14884
rect 25998 14844 26424 14872
rect 25998 14841 26010 14844
rect 25952 14835 26010 14841
rect 26418 14832 26424 14844
rect 26476 14832 26482 14884
rect 17083 14776 17264 14804
rect 17083 14773 17095 14776
rect 17037 14767 17095 14773
rect 17494 14764 17500 14816
rect 17552 14804 17558 14816
rect 17773 14807 17831 14813
rect 17773 14804 17785 14807
rect 17552 14776 17785 14804
rect 17552 14764 17558 14776
rect 17773 14773 17785 14776
rect 17819 14773 17831 14807
rect 17773 14767 17831 14773
rect 17954 14764 17960 14816
rect 18012 14804 18018 14816
rect 18509 14807 18567 14813
rect 18509 14804 18521 14807
rect 18012 14776 18521 14804
rect 18012 14764 18018 14776
rect 18509 14773 18521 14776
rect 18555 14773 18567 14807
rect 18509 14767 18567 14773
rect 23382 14764 23388 14816
rect 23440 14804 23446 14816
rect 24964 14804 24992 14832
rect 23440 14776 24992 14804
rect 25317 14807 25375 14813
rect 23440 14764 23446 14776
rect 25317 14773 25329 14807
rect 25363 14804 25375 14807
rect 26878 14804 26884 14816
rect 25363 14776 26884 14804
rect 25363 14773 25375 14776
rect 25317 14767 25375 14773
rect 26878 14764 26884 14776
rect 26936 14764 26942 14816
rect 552 14714 27576 14736
rect 552 14662 7114 14714
rect 7166 14662 7178 14714
rect 7230 14662 7242 14714
rect 7294 14662 7306 14714
rect 7358 14662 7370 14714
rect 7422 14662 13830 14714
rect 13882 14662 13894 14714
rect 13946 14662 13958 14714
rect 14010 14662 14022 14714
rect 14074 14662 14086 14714
rect 14138 14662 20546 14714
rect 20598 14662 20610 14714
rect 20662 14662 20674 14714
rect 20726 14662 20738 14714
rect 20790 14662 20802 14714
rect 20854 14662 27262 14714
rect 27314 14662 27326 14714
rect 27378 14662 27390 14714
rect 27442 14662 27454 14714
rect 27506 14662 27518 14714
rect 27570 14662 27576 14714
rect 552 14640 27576 14662
rect 2038 14600 2044 14612
rect 1688 14572 2044 14600
rect 1688 14544 1716 14572
rect 2038 14560 2044 14572
rect 2096 14560 2102 14612
rect 3326 14600 3332 14612
rect 2700 14572 3332 14600
rect 1670 14492 1676 14544
rect 1728 14492 1734 14544
rect 2700 14541 2728 14572
rect 3326 14560 3332 14572
rect 3384 14560 3390 14612
rect 9490 14600 9496 14612
rect 3712 14572 9496 14600
rect 3712 14541 3740 14572
rect 9490 14560 9496 14572
rect 9548 14560 9554 14612
rect 16850 14560 16856 14612
rect 16908 14560 16914 14612
rect 22465 14603 22523 14609
rect 22465 14569 22477 14603
rect 22511 14569 22523 14603
rect 22465 14563 22523 14569
rect 23569 14603 23627 14609
rect 23569 14569 23581 14603
rect 23615 14569 23627 14603
rect 23569 14563 23627 14569
rect 1857 14535 1915 14541
rect 1857 14501 1869 14535
rect 1903 14532 1915 14535
rect 2685 14535 2743 14541
rect 2685 14532 2697 14535
rect 1903 14504 2697 14532
rect 1903 14501 1915 14504
rect 1857 14495 1915 14501
rect 2685 14501 2697 14504
rect 2731 14501 2743 14535
rect 2685 14495 2743 14501
rect 2901 14535 2959 14541
rect 2901 14501 2913 14535
rect 2947 14532 2959 14535
rect 3697 14535 3755 14541
rect 2947 14504 3188 14532
rect 2947 14501 2959 14504
rect 2901 14495 2959 14501
rect 3160 14476 3188 14504
rect 3697 14501 3709 14535
rect 3743 14501 3755 14535
rect 3697 14495 3755 14501
rect 5074 14492 5080 14544
rect 5132 14492 5138 14544
rect 6181 14535 6239 14541
rect 6181 14532 6193 14535
rect 5736 14504 6193 14532
rect 1949 14467 2007 14473
rect 1949 14433 1961 14467
rect 1995 14433 2007 14467
rect 1949 14427 2007 14433
rect 1578 14220 1584 14272
rect 1636 14260 1642 14272
rect 1673 14263 1731 14269
rect 1673 14260 1685 14263
rect 1636 14232 1685 14260
rect 1636 14220 1642 14232
rect 1673 14229 1685 14232
rect 1719 14229 1731 14263
rect 1964 14260 1992 14427
rect 3142 14424 3148 14476
rect 3200 14424 3206 14476
rect 3326 14424 3332 14476
rect 3384 14424 3390 14476
rect 4798 14424 4804 14476
rect 4856 14424 4862 14476
rect 4893 14467 4951 14473
rect 4893 14433 4905 14467
rect 4939 14464 4951 14467
rect 5442 14464 5448 14476
rect 4939 14436 5448 14464
rect 4939 14433 4951 14436
rect 4893 14427 4951 14433
rect 5442 14424 5448 14436
rect 5500 14424 5506 14476
rect 4522 14356 4528 14408
rect 4580 14356 4586 14408
rect 4816 14396 4844 14424
rect 5736 14396 5764 14504
rect 6181 14501 6193 14504
rect 6227 14532 6239 14535
rect 6457 14535 6515 14541
rect 6457 14532 6469 14535
rect 6227 14504 6469 14532
rect 6227 14501 6239 14504
rect 6181 14495 6239 14501
rect 6457 14501 6469 14504
rect 6503 14501 6515 14535
rect 6457 14495 6515 14501
rect 7926 14492 7932 14544
rect 7984 14532 7990 14544
rect 8389 14535 8447 14541
rect 8389 14532 8401 14535
rect 7984 14504 8401 14532
rect 7984 14492 7990 14504
rect 8389 14501 8401 14504
rect 8435 14501 8447 14535
rect 8389 14495 8447 14501
rect 11330 14492 11336 14544
rect 11388 14492 11394 14544
rect 15562 14492 15568 14544
rect 15620 14532 15626 14544
rect 17405 14535 17463 14541
rect 17405 14532 17417 14535
rect 15620 14504 17417 14532
rect 15620 14492 15626 14504
rect 17405 14501 17417 14504
rect 17451 14501 17463 14535
rect 17405 14495 17463 14501
rect 17494 14492 17500 14544
rect 17552 14492 17558 14544
rect 22094 14532 22100 14544
rect 17972 14504 18828 14532
rect 17972 14476 18000 14504
rect 6917 14467 6975 14473
rect 6917 14433 6929 14467
rect 6963 14464 6975 14467
rect 7650 14464 7656 14476
rect 6963 14436 7656 14464
rect 6963 14433 6975 14436
rect 6917 14427 6975 14433
rect 7650 14424 7656 14436
rect 7708 14424 7714 14476
rect 7742 14424 7748 14476
rect 7800 14424 7806 14476
rect 8202 14424 8208 14476
rect 8260 14464 8266 14476
rect 8849 14467 8907 14473
rect 8849 14464 8861 14467
rect 8260 14436 8861 14464
rect 8260 14424 8266 14436
rect 8849 14433 8861 14436
rect 8895 14433 8907 14467
rect 8849 14427 8907 14433
rect 4816 14368 5764 14396
rect 6825 14399 6883 14405
rect 6825 14365 6837 14399
rect 6871 14396 6883 14399
rect 7466 14396 7472 14408
rect 6871 14368 7472 14396
rect 6871 14365 6883 14368
rect 6825 14359 6883 14365
rect 7466 14356 7472 14368
rect 7524 14356 7530 14408
rect 8754 14356 8760 14408
rect 8812 14356 8818 14408
rect 8864 14396 8892 14427
rect 9582 14424 9588 14476
rect 9640 14424 9646 14476
rect 11238 14424 11244 14476
rect 11296 14464 11302 14476
rect 11425 14467 11483 14473
rect 11425 14464 11437 14467
rect 11296 14436 11437 14464
rect 11296 14424 11302 14436
rect 11425 14433 11437 14436
rect 11471 14433 11483 14467
rect 11425 14427 11483 14433
rect 11698 14424 11704 14476
rect 11756 14424 11762 14476
rect 11793 14467 11851 14473
rect 11793 14433 11805 14467
rect 11839 14464 11851 14467
rect 11882 14464 11888 14476
rect 11839 14436 11888 14464
rect 11839 14433 11851 14436
rect 11793 14427 11851 14433
rect 11882 14424 11888 14436
rect 11940 14424 11946 14476
rect 12066 14473 12072 14476
rect 12060 14427 12072 14473
rect 12066 14424 12072 14427
rect 12124 14424 12130 14476
rect 14550 14473 14556 14476
rect 14544 14427 14556 14473
rect 14550 14424 14556 14427
rect 14608 14424 14614 14476
rect 17034 14424 17040 14476
rect 17092 14424 17098 14476
rect 17129 14467 17187 14473
rect 17129 14433 17141 14467
rect 17175 14464 17187 14467
rect 17954 14464 17960 14476
rect 17175 14436 17960 14464
rect 17175 14433 17187 14436
rect 17129 14427 17187 14433
rect 17954 14424 17960 14436
rect 18012 14424 18018 14476
rect 18138 14424 18144 14476
rect 18196 14464 18202 14476
rect 18702 14467 18760 14473
rect 18702 14464 18714 14467
rect 18196 14436 18714 14464
rect 18196 14424 18202 14436
rect 18702 14433 18714 14436
rect 18748 14433 18760 14467
rect 18800 14464 18828 14504
rect 19076 14504 22100 14532
rect 19076 14473 19104 14504
rect 22094 14492 22100 14504
rect 22152 14492 22158 14544
rect 22480 14532 22508 14563
rect 23014 14532 23020 14544
rect 22480 14504 23020 14532
rect 23014 14492 23020 14504
rect 23072 14532 23078 14544
rect 23072 14504 23244 14532
rect 23072 14492 23078 14504
rect 18969 14467 19027 14473
rect 18800 14436 18920 14464
rect 18702 14427 18760 14433
rect 13817 14399 13875 14405
rect 13817 14396 13829 14399
rect 8864 14368 9444 14396
rect 5813 14331 5871 14337
rect 2884 14300 3188 14328
rect 2222 14260 2228 14272
rect 1964 14232 2228 14260
rect 1673 14223 1731 14229
rect 2222 14220 2228 14232
rect 2280 14260 2286 14272
rect 2884 14269 2912 14300
rect 2869 14263 2927 14269
rect 2869 14260 2881 14263
rect 2280 14232 2881 14260
rect 2280 14220 2286 14232
rect 2869 14229 2881 14232
rect 2915 14229 2927 14263
rect 2869 14223 2927 14229
rect 2958 14220 2964 14272
rect 3016 14260 3022 14272
rect 3160 14269 3188 14300
rect 5813 14297 5825 14331
rect 5859 14328 5871 14331
rect 5859 14300 6868 14328
rect 5859 14297 5871 14300
rect 5813 14291 5871 14297
rect 3053 14263 3111 14269
rect 3053 14260 3065 14263
rect 3016 14232 3065 14260
rect 3016 14220 3022 14232
rect 3053 14229 3065 14232
rect 3099 14229 3111 14263
rect 3053 14223 3111 14229
rect 3145 14263 3203 14269
rect 3145 14229 3157 14263
rect 3191 14229 3203 14263
rect 3145 14223 3203 14229
rect 3513 14263 3571 14269
rect 3513 14229 3525 14263
rect 3559 14260 3571 14263
rect 5902 14260 5908 14272
rect 3559 14232 5908 14260
rect 3559 14229 3571 14232
rect 3513 14223 3571 14229
rect 5902 14220 5908 14232
rect 5960 14220 5966 14272
rect 6178 14220 6184 14272
rect 6236 14220 6242 14272
rect 6270 14220 6276 14272
rect 6328 14260 6334 14272
rect 6840 14269 6868 14300
rect 7006 14288 7012 14340
rect 7064 14328 7070 14340
rect 7101 14331 7159 14337
rect 7101 14328 7113 14331
rect 7064 14300 7113 14328
rect 7064 14288 7070 14300
rect 7101 14297 7113 14300
rect 7147 14297 7159 14331
rect 7101 14291 7159 14297
rect 9214 14288 9220 14340
rect 9272 14288 9278 14340
rect 9416 14337 9444 14368
rect 13188 14368 13829 14396
rect 9401 14331 9459 14337
rect 9401 14297 9413 14331
rect 9447 14297 9459 14331
rect 9401 14291 9459 14297
rect 13188 14272 13216 14368
rect 13817 14365 13829 14368
rect 13863 14365 13875 14399
rect 13817 14359 13875 14365
rect 14274 14356 14280 14408
rect 14332 14356 14338 14408
rect 16298 14356 16304 14408
rect 16356 14396 16362 14408
rect 16669 14399 16727 14405
rect 16669 14396 16681 14399
rect 16356 14368 16681 14396
rect 16356 14356 16362 14368
rect 16669 14365 16681 14368
rect 16715 14365 16727 14399
rect 18892 14396 18920 14436
rect 18969 14433 18981 14467
rect 19015 14464 19027 14467
rect 19061 14467 19119 14473
rect 19061 14464 19073 14467
rect 19015 14436 19073 14464
rect 19015 14433 19027 14436
rect 18969 14427 19027 14433
rect 19061 14433 19073 14436
rect 19107 14433 19119 14467
rect 19317 14467 19375 14473
rect 19317 14464 19329 14467
rect 19061 14427 19119 14433
rect 19168 14436 19329 14464
rect 19168 14396 19196 14436
rect 19317 14433 19329 14436
rect 19363 14433 19375 14467
rect 19317 14427 19375 14433
rect 20625 14467 20683 14473
rect 20625 14433 20637 14467
rect 20671 14464 20683 14467
rect 21082 14464 21088 14476
rect 20671 14436 21088 14464
rect 20671 14433 20683 14436
rect 20625 14427 20683 14433
rect 21082 14424 21088 14436
rect 21140 14424 21146 14476
rect 21266 14424 21272 14476
rect 21324 14424 21330 14476
rect 22281 14467 22339 14473
rect 22281 14464 22293 14467
rect 22066 14436 22293 14464
rect 18892 14368 19196 14396
rect 16669 14359 16727 14365
rect 15657 14331 15715 14337
rect 15657 14297 15669 14331
rect 15703 14328 15715 14331
rect 16316 14328 16344 14356
rect 15703 14300 16344 14328
rect 21284 14328 21312 14424
rect 21726 14356 21732 14408
rect 21784 14396 21790 14408
rect 22066 14396 22094 14436
rect 22281 14433 22293 14436
rect 22327 14433 22339 14467
rect 22281 14427 22339 14433
rect 22646 14424 22652 14476
rect 22704 14464 22710 14476
rect 23216 14473 23244 14504
rect 22925 14467 22983 14473
rect 22925 14464 22937 14467
rect 22704 14436 22937 14464
rect 22704 14424 22710 14436
rect 22925 14433 22937 14436
rect 22971 14433 22983 14467
rect 22925 14427 22983 14433
rect 23109 14467 23167 14473
rect 23109 14433 23121 14467
rect 23155 14433 23167 14467
rect 23109 14427 23167 14433
rect 23201 14467 23259 14473
rect 23201 14433 23213 14467
rect 23247 14433 23259 14467
rect 23201 14427 23259 14433
rect 21784 14368 22094 14396
rect 23124 14396 23152 14427
rect 23290 14424 23296 14476
rect 23348 14424 23354 14476
rect 23584 14464 23612 14563
rect 23750 14560 23756 14612
rect 23808 14600 23814 14612
rect 23808 14572 23888 14600
rect 23808 14560 23814 14572
rect 23860 14532 23888 14572
rect 25038 14560 25044 14612
rect 25096 14560 25102 14612
rect 25317 14535 25375 14541
rect 25317 14532 25329 14535
rect 23860 14504 25329 14532
rect 25317 14501 25329 14504
rect 25363 14501 25375 14535
rect 25317 14495 25375 14501
rect 25682 14492 25688 14544
rect 25740 14532 25746 14544
rect 26053 14535 26111 14541
rect 26053 14532 26065 14535
rect 25740 14504 26065 14532
rect 25740 14492 25746 14504
rect 26053 14501 26065 14504
rect 26099 14501 26111 14535
rect 26053 14495 26111 14501
rect 23917 14467 23975 14473
rect 23917 14464 23929 14467
rect 23584 14436 23929 14464
rect 23917 14433 23929 14436
rect 23963 14433 23975 14467
rect 23917 14427 23975 14433
rect 26602 14424 26608 14476
rect 26660 14464 26666 14476
rect 26697 14467 26755 14473
rect 26697 14464 26709 14467
rect 26660 14436 26709 14464
rect 26660 14424 26666 14436
rect 26697 14433 26709 14436
rect 26743 14433 26755 14467
rect 26697 14427 26755 14433
rect 26789 14467 26847 14473
rect 26789 14433 26801 14467
rect 26835 14433 26847 14467
rect 26789 14427 26847 14433
rect 23474 14396 23480 14408
rect 23124 14368 23480 14396
rect 21784 14356 21790 14368
rect 23474 14356 23480 14368
rect 23532 14356 23538 14408
rect 23661 14399 23719 14405
rect 23661 14365 23673 14399
rect 23707 14365 23719 14399
rect 23661 14359 23719 14365
rect 22002 14328 22008 14340
rect 21284 14300 22008 14328
rect 15703 14297 15715 14300
rect 15657 14291 15715 14297
rect 22002 14288 22008 14300
rect 22060 14328 22066 14340
rect 23566 14328 23572 14340
rect 22060 14300 23572 14328
rect 22060 14288 22066 14300
rect 23566 14288 23572 14300
rect 23624 14288 23630 14340
rect 6365 14263 6423 14269
rect 6365 14260 6377 14263
rect 6328 14232 6377 14260
rect 6328 14220 6334 14232
rect 6365 14229 6377 14232
rect 6411 14229 6423 14263
rect 6365 14223 6423 14229
rect 6825 14263 6883 14269
rect 6825 14229 6837 14263
rect 6871 14260 6883 14263
rect 6914 14260 6920 14272
rect 6871 14232 6920 14260
rect 6871 14229 6883 14232
rect 6825 14223 6883 14229
rect 6914 14220 6920 14232
rect 6972 14220 6978 14272
rect 13170 14220 13176 14272
rect 13228 14220 13234 14272
rect 13262 14220 13268 14272
rect 13320 14220 13326 14272
rect 13446 14220 13452 14272
rect 13504 14260 13510 14272
rect 15010 14260 15016 14272
rect 13504 14232 15016 14260
rect 13504 14220 13510 14232
rect 15010 14220 15016 14232
rect 15068 14220 15074 14272
rect 16114 14220 16120 14272
rect 16172 14220 16178 14272
rect 17589 14263 17647 14269
rect 17589 14229 17601 14263
rect 17635 14260 17647 14263
rect 18690 14260 18696 14272
rect 17635 14232 18696 14260
rect 17635 14229 17647 14232
rect 17589 14223 17647 14229
rect 18690 14220 18696 14232
rect 18748 14220 18754 14272
rect 20441 14263 20499 14269
rect 20441 14229 20453 14263
rect 20487 14260 20499 14263
rect 20714 14260 20720 14272
rect 20487 14232 20720 14260
rect 20487 14229 20499 14232
rect 20441 14223 20499 14229
rect 20714 14220 20720 14232
rect 20772 14220 20778 14272
rect 21085 14263 21143 14269
rect 21085 14229 21097 14263
rect 21131 14260 21143 14263
rect 23382 14260 23388 14272
rect 21131 14232 23388 14260
rect 21131 14229 21143 14232
rect 21085 14223 21143 14229
rect 23382 14220 23388 14232
rect 23440 14220 23446 14272
rect 23676 14260 23704 14359
rect 24946 14356 24952 14408
rect 25004 14396 25010 14408
rect 26804 14396 26832 14427
rect 26878 14424 26884 14476
rect 26936 14424 26942 14476
rect 26970 14424 26976 14476
rect 27028 14464 27034 14476
rect 27065 14467 27123 14473
rect 27065 14464 27077 14467
rect 27028 14436 27077 14464
rect 27028 14424 27034 14436
rect 27065 14433 27077 14436
rect 27111 14433 27123 14467
rect 27065 14427 27123 14433
rect 25004 14368 26832 14396
rect 25004 14356 25010 14368
rect 25682 14328 25688 14340
rect 24596 14300 25688 14328
rect 24596 14260 24624 14300
rect 25682 14288 25688 14300
rect 25740 14288 25746 14340
rect 23676 14232 24624 14260
rect 25774 14220 25780 14272
rect 25832 14260 25838 14272
rect 26421 14263 26479 14269
rect 26421 14260 26433 14263
rect 25832 14232 26433 14260
rect 25832 14220 25838 14232
rect 26421 14229 26433 14232
rect 26467 14229 26479 14263
rect 26421 14223 26479 14229
rect 552 14170 27416 14192
rect 552 14118 3756 14170
rect 3808 14118 3820 14170
rect 3872 14118 3884 14170
rect 3936 14118 3948 14170
rect 4000 14118 4012 14170
rect 4064 14118 10472 14170
rect 10524 14118 10536 14170
rect 10588 14118 10600 14170
rect 10652 14118 10664 14170
rect 10716 14118 10728 14170
rect 10780 14118 17188 14170
rect 17240 14118 17252 14170
rect 17304 14118 17316 14170
rect 17368 14118 17380 14170
rect 17432 14118 17444 14170
rect 17496 14118 23904 14170
rect 23956 14118 23968 14170
rect 24020 14118 24032 14170
rect 24084 14118 24096 14170
rect 24148 14118 24160 14170
rect 24212 14118 27416 14170
rect 552 14096 27416 14118
rect 2222 14016 2228 14068
rect 2280 14056 2286 14068
rect 2280 14028 2774 14056
rect 2280 14016 2286 14028
rect 845 13855 903 13861
rect 845 13821 857 13855
rect 891 13852 903 13855
rect 1394 13852 1400 13864
rect 891 13824 1400 13852
rect 891 13821 903 13824
rect 845 13815 903 13821
rect 1394 13812 1400 13824
rect 1452 13812 1458 13864
rect 2746 13852 2774 14028
rect 3142 14016 3148 14068
rect 3200 14056 3206 14068
rect 3237 14059 3295 14065
rect 3237 14056 3249 14059
rect 3200 14028 3249 14056
rect 3200 14016 3206 14028
rect 3237 14025 3249 14028
rect 3283 14025 3295 14059
rect 3237 14019 3295 14025
rect 10870 14016 10876 14068
rect 10928 14056 10934 14068
rect 10928 14028 11376 14056
rect 10928 14016 10934 14028
rect 8478 13948 8484 14000
rect 8536 13988 8542 14000
rect 8573 13991 8631 13997
rect 8573 13988 8585 13991
rect 8536 13960 8585 13988
rect 8536 13948 8542 13960
rect 8573 13957 8585 13960
rect 8619 13988 8631 13991
rect 10042 13988 10048 14000
rect 8619 13960 10048 13988
rect 8619 13957 8631 13960
rect 8573 13951 8631 13957
rect 10042 13948 10048 13960
rect 10100 13948 10106 14000
rect 11149 13923 11207 13929
rect 11149 13920 11161 13923
rect 10980 13892 11161 13920
rect 10980 13864 11008 13892
rect 11149 13889 11161 13892
rect 11195 13889 11207 13923
rect 11149 13883 11207 13889
rect 2961 13855 3019 13861
rect 2961 13852 2973 13855
rect 2746 13824 2973 13852
rect 2961 13821 2973 13824
rect 3007 13852 3019 13855
rect 3418 13852 3424 13864
rect 3007 13824 3424 13852
rect 3007 13821 3019 13824
rect 2961 13815 3019 13821
rect 3418 13812 3424 13824
rect 3476 13812 3482 13864
rect 4522 13812 4528 13864
rect 4580 13852 4586 13864
rect 4617 13855 4675 13861
rect 4617 13852 4629 13855
rect 4580 13824 4629 13852
rect 4580 13812 4586 13824
rect 4617 13821 4629 13824
rect 4663 13821 4675 13855
rect 4617 13815 4675 13821
rect 5077 13855 5135 13861
rect 5077 13821 5089 13855
rect 5123 13852 5135 13855
rect 5166 13852 5172 13864
rect 5123 13824 5172 13852
rect 5123 13821 5135 13824
rect 5077 13815 5135 13821
rect 5166 13812 5172 13824
rect 5224 13812 5230 13864
rect 5261 13855 5319 13861
rect 5261 13821 5273 13855
rect 5307 13852 5319 13855
rect 5442 13852 5448 13864
rect 5307 13824 5448 13852
rect 5307 13821 5319 13824
rect 5261 13815 5319 13821
rect 5442 13812 5448 13824
rect 5500 13812 5506 13864
rect 6546 13812 6552 13864
rect 6604 13812 6610 13864
rect 6638 13812 6644 13864
rect 6696 13812 6702 13864
rect 6733 13855 6791 13861
rect 6733 13821 6745 13855
rect 6779 13852 6791 13855
rect 6822 13852 6828 13864
rect 6779 13824 6828 13852
rect 6779 13821 6791 13824
rect 6733 13815 6791 13821
rect 6822 13812 6828 13824
rect 6880 13812 6886 13864
rect 8110 13812 8116 13864
rect 8168 13852 8174 13864
rect 8205 13855 8263 13861
rect 8205 13852 8217 13855
rect 8168 13824 8217 13852
rect 8168 13812 8174 13824
rect 8205 13821 8217 13824
rect 8251 13852 8263 13855
rect 8389 13855 8447 13861
rect 8389 13852 8401 13855
rect 8251 13824 8401 13852
rect 8251 13821 8263 13824
rect 8205 13815 8263 13821
rect 8389 13821 8401 13824
rect 8435 13852 8447 13855
rect 8757 13855 8815 13861
rect 8757 13852 8769 13855
rect 8435 13824 8769 13852
rect 8435 13821 8447 13824
rect 8389 13815 8447 13821
rect 8757 13821 8769 13824
rect 8803 13821 8815 13855
rect 8757 13815 8815 13821
rect 10962 13812 10968 13864
rect 11020 13812 11026 13864
rect 11348 13861 11376 14028
rect 12066 14016 12072 14068
rect 12124 14056 12130 14068
rect 12161 14059 12219 14065
rect 12161 14056 12173 14059
rect 12124 14028 12173 14056
rect 12124 14016 12130 14028
rect 12161 14025 12173 14028
rect 12207 14025 12219 14059
rect 12161 14019 12219 14025
rect 12897 14059 12955 14065
rect 12897 14025 12909 14059
rect 12943 14056 12955 14059
rect 13262 14056 13268 14068
rect 12943 14028 13268 14056
rect 12943 14025 12955 14028
rect 12897 14019 12955 14025
rect 13262 14016 13268 14028
rect 13320 14016 13326 14068
rect 14458 14016 14464 14068
rect 14516 14016 14522 14068
rect 14550 14016 14556 14068
rect 14608 14056 14614 14068
rect 14737 14059 14795 14065
rect 14737 14056 14749 14059
rect 14608 14028 14749 14056
rect 14608 14016 14614 14028
rect 14737 14025 14749 14028
rect 14783 14025 14795 14059
rect 14737 14019 14795 14025
rect 15010 14016 15016 14068
rect 15068 14056 15074 14068
rect 15473 14059 15531 14065
rect 15068 14028 15424 14056
rect 15068 14016 15074 14028
rect 12713 13991 12771 13997
rect 12713 13988 12725 13991
rect 12406 13960 12725 13988
rect 12406 13920 12434 13960
rect 12713 13957 12725 13960
rect 12759 13957 12771 13991
rect 12713 13951 12771 13957
rect 13357 13991 13415 13997
rect 13357 13957 13369 13991
rect 13403 13988 13415 13991
rect 14476 13988 14504 14016
rect 15102 13988 15108 14000
rect 13403 13960 15108 13988
rect 13403 13957 13415 13960
rect 13357 13951 13415 13957
rect 15102 13948 15108 13960
rect 15160 13948 15166 14000
rect 15289 13991 15347 13997
rect 15289 13957 15301 13991
rect 15335 13957 15347 13991
rect 15396 13988 15424 14028
rect 15473 14025 15485 14059
rect 15519 14056 15531 14059
rect 16114 14056 16120 14068
rect 15519 14028 16120 14056
rect 15519 14025 15531 14028
rect 15473 14019 15531 14025
rect 16114 14016 16120 14028
rect 16172 14016 16178 14068
rect 18049 14059 18107 14065
rect 18049 14025 18061 14059
rect 18095 14056 18107 14059
rect 18138 14056 18144 14068
rect 18095 14028 18144 14056
rect 18095 14025 18107 14028
rect 18049 14019 18107 14025
rect 18138 14016 18144 14028
rect 18196 14016 18202 14068
rect 19337 14059 19395 14065
rect 19337 14025 19349 14059
rect 19383 14056 19395 14059
rect 19613 14059 19671 14065
rect 19613 14056 19625 14059
rect 19383 14028 19625 14056
rect 19383 14025 19395 14028
rect 19337 14019 19395 14025
rect 19613 14025 19625 14028
rect 19659 14025 19671 14059
rect 19613 14019 19671 14025
rect 20073 14059 20131 14065
rect 20073 14025 20085 14059
rect 20119 14025 20131 14059
rect 20073 14019 20131 14025
rect 20717 14059 20775 14065
rect 20717 14025 20729 14059
rect 20763 14056 20775 14059
rect 21358 14056 21364 14068
rect 20763 14028 21364 14056
rect 20763 14025 20775 14028
rect 20717 14019 20775 14025
rect 18598 13988 18604 14000
rect 15396 13960 18604 13988
rect 15289 13951 15347 13957
rect 14182 13920 14188 13932
rect 12360 13892 12434 13920
rect 12912 13892 13400 13920
rect 12360 13861 12388 13892
rect 11057 13855 11115 13861
rect 11057 13821 11069 13855
rect 11103 13821 11115 13855
rect 11057 13815 11115 13821
rect 11333 13855 11391 13861
rect 11333 13821 11345 13855
rect 11379 13821 11391 13855
rect 11333 13815 11391 13821
rect 12345 13855 12403 13861
rect 12345 13821 12357 13855
rect 12391 13821 12403 13855
rect 12345 13815 12403 13821
rect 1112 13787 1170 13793
rect 1112 13753 1124 13787
rect 1158 13784 1170 13787
rect 1302 13784 1308 13796
rect 1158 13756 1308 13784
rect 1158 13753 1170 13756
rect 1112 13747 1170 13753
rect 1302 13744 1308 13756
rect 1360 13744 1366 13796
rect 4154 13744 4160 13796
rect 4212 13784 4218 13796
rect 4350 13787 4408 13793
rect 4350 13784 4362 13787
rect 4212 13756 4362 13784
rect 4212 13744 4218 13756
rect 4350 13753 4362 13756
rect 4396 13753 4408 13787
rect 4350 13747 4408 13753
rect 4706 13744 4712 13796
rect 4764 13784 4770 13796
rect 6656 13784 6684 13812
rect 4764 13756 6684 13784
rect 4764 13744 4770 13756
rect 10318 13744 10324 13796
rect 10376 13784 10382 13796
rect 10790 13787 10848 13793
rect 10790 13784 10802 13787
rect 10376 13756 10802 13784
rect 10376 13744 10382 13756
rect 10790 13753 10802 13756
rect 10836 13753 10848 13787
rect 10790 13747 10848 13753
rect 1762 13676 1768 13728
rect 1820 13716 1826 13728
rect 2317 13719 2375 13725
rect 2317 13716 2329 13719
rect 1820 13688 2329 13716
rect 1820 13676 1826 13688
rect 2317 13685 2329 13688
rect 2363 13685 2375 13719
rect 2317 13679 2375 13685
rect 3878 13676 3884 13728
rect 3936 13716 3942 13728
rect 4614 13716 4620 13728
rect 3936 13688 4620 13716
rect 3936 13676 3942 13688
rect 4614 13676 4620 13688
rect 4672 13716 4678 13728
rect 4893 13719 4951 13725
rect 4893 13716 4905 13719
rect 4672 13688 4905 13716
rect 4672 13676 4678 13688
rect 4893 13685 4905 13688
rect 4939 13685 4951 13719
rect 4893 13679 4951 13685
rect 6641 13719 6699 13725
rect 6641 13685 6653 13719
rect 6687 13716 6699 13719
rect 6730 13716 6736 13728
rect 6687 13688 6736 13716
rect 6687 13685 6699 13688
rect 6641 13679 6699 13685
rect 6730 13676 6736 13688
rect 6788 13676 6794 13728
rect 7926 13676 7932 13728
rect 7984 13716 7990 13728
rect 8021 13719 8079 13725
rect 8021 13716 8033 13719
rect 7984 13688 8033 13716
rect 7984 13676 7990 13688
rect 8021 13685 8033 13688
rect 8067 13685 8079 13719
rect 8021 13679 8079 13685
rect 8938 13676 8944 13728
rect 8996 13676 9002 13728
rect 9677 13719 9735 13725
rect 9677 13685 9689 13719
rect 9723 13716 9735 13719
rect 9950 13716 9956 13728
rect 9723 13688 9956 13716
rect 9723 13685 9735 13688
rect 9677 13679 9735 13685
rect 9950 13676 9956 13688
rect 10008 13676 10014 13728
rect 11072 13716 11100 13815
rect 12618 13812 12624 13864
rect 12676 13812 12682 13864
rect 11514 13744 11520 13796
rect 11572 13784 11578 13796
rect 12158 13784 12164 13796
rect 11572 13756 12164 13784
rect 11572 13744 11578 13756
rect 12158 13744 12164 13756
rect 12216 13784 12222 13796
rect 12912 13784 12940 13892
rect 13372 13864 13400 13892
rect 13464 13892 14188 13920
rect 13173 13855 13231 13861
rect 13173 13821 13185 13855
rect 13219 13852 13231 13855
rect 13219 13824 13308 13852
rect 13219 13821 13231 13824
rect 13173 13815 13231 13821
rect 12216 13756 12940 13784
rect 12216 13744 12222 13756
rect 12986 13744 12992 13796
rect 13044 13784 13050 13796
rect 13081 13787 13139 13793
rect 13081 13784 13093 13787
rect 13044 13756 13093 13784
rect 13044 13744 13050 13756
rect 13081 13753 13093 13756
rect 13127 13753 13139 13787
rect 13280 13784 13308 13824
rect 13354 13812 13360 13864
rect 13412 13812 13418 13864
rect 13464 13784 13492 13892
rect 14182 13880 14188 13892
rect 14240 13880 14246 13932
rect 14274 13880 14280 13932
rect 14332 13920 14338 13932
rect 14553 13923 14611 13929
rect 14553 13920 14565 13923
rect 14332 13892 14565 13920
rect 14332 13880 14338 13892
rect 14553 13889 14565 13892
rect 14599 13920 14611 13923
rect 14642 13920 14648 13932
rect 14599 13892 14648 13920
rect 14599 13889 14611 13892
rect 14553 13883 14611 13889
rect 14642 13880 14648 13892
rect 14700 13880 14706 13932
rect 15304 13920 15332 13951
rect 14936 13892 15332 13920
rect 13722 13812 13728 13864
rect 13780 13812 13786 13864
rect 14936 13861 14964 13892
rect 14921 13855 14979 13861
rect 14921 13821 14933 13855
rect 14967 13821 14979 13855
rect 14921 13815 14979 13821
rect 15102 13812 15108 13864
rect 15160 13852 15166 13864
rect 15197 13855 15255 13861
rect 15197 13852 15209 13855
rect 15160 13824 15209 13852
rect 15160 13812 15166 13824
rect 15197 13821 15209 13824
rect 15243 13821 15255 13855
rect 15197 13815 15255 13821
rect 16758 13812 16764 13864
rect 16816 13812 16822 13864
rect 17328 13861 17356 13960
rect 18598 13948 18604 13960
rect 18656 13948 18662 14000
rect 19429 13991 19487 13997
rect 19429 13957 19441 13991
rect 19475 13957 19487 13991
rect 19429 13951 19487 13957
rect 19444 13920 19472 13951
rect 19518 13948 19524 14000
rect 19576 13988 19582 14000
rect 20088 13988 20116 14019
rect 21358 14016 21364 14028
rect 21416 14016 21422 14068
rect 21726 14016 21732 14068
rect 21784 14016 21790 14068
rect 22094 14056 22100 14068
rect 21836 14028 22100 14056
rect 19576 13960 20116 13988
rect 20533 13991 20591 13997
rect 19576 13948 19582 13960
rect 20533 13957 20545 13991
rect 20579 13988 20591 13991
rect 20990 13988 20996 14000
rect 20579 13960 20996 13988
rect 20579 13957 20591 13960
rect 20533 13951 20591 13957
rect 20990 13948 20996 13960
rect 21048 13948 21054 14000
rect 21082 13948 21088 14000
rect 21140 13988 21146 14000
rect 21545 13991 21603 13997
rect 21545 13988 21557 13991
rect 21140 13960 21557 13988
rect 21140 13948 21146 13960
rect 21545 13957 21557 13960
rect 21591 13957 21603 13991
rect 21545 13951 21603 13957
rect 18248 13892 19472 13920
rect 19996 13892 20668 13920
rect 17129 13855 17187 13861
rect 17129 13821 17141 13855
rect 17175 13852 17187 13855
rect 17313 13855 17371 13861
rect 17175 13824 17264 13852
rect 17175 13821 17187 13824
rect 17129 13815 17187 13821
rect 13280 13756 13492 13784
rect 13081 13747 13139 13753
rect 14550 13744 14556 13796
rect 14608 13784 14614 13796
rect 15657 13787 15715 13793
rect 15657 13784 15669 13787
rect 14608 13756 15669 13784
rect 14608 13744 14614 13756
rect 15657 13753 15669 13756
rect 15703 13753 15715 13787
rect 17236 13784 17264 13824
rect 17313 13821 17325 13855
rect 17359 13821 17371 13855
rect 17313 13815 17371 13821
rect 17405 13855 17463 13861
rect 17405 13821 17417 13855
rect 17451 13852 17463 13855
rect 17586 13852 17592 13864
rect 17451 13824 17592 13852
rect 17451 13821 17463 13824
rect 17405 13815 17463 13821
rect 17586 13812 17592 13824
rect 17644 13852 17650 13864
rect 18248 13861 18276 13892
rect 18233 13855 18291 13861
rect 17644 13824 18184 13852
rect 17644 13812 17650 13824
rect 18046 13784 18052 13796
rect 17236 13756 18052 13784
rect 15657 13747 15715 13753
rect 18046 13744 18052 13756
rect 18104 13744 18110 13796
rect 18156 13784 18184 13824
rect 18233 13821 18245 13855
rect 18279 13821 18291 13855
rect 18506 13852 18512 13864
rect 18233 13815 18291 13821
rect 18340 13824 18512 13852
rect 18340 13784 18368 13824
rect 18506 13812 18512 13824
rect 18564 13812 18570 13864
rect 18690 13812 18696 13864
rect 18748 13812 18754 13864
rect 18966 13852 18972 13864
rect 18800 13824 18972 13852
rect 18156 13756 18368 13784
rect 18417 13787 18475 13793
rect 18417 13753 18429 13787
rect 18463 13784 18475 13787
rect 18800 13784 18828 13824
rect 18966 13812 18972 13824
rect 19024 13812 19030 13864
rect 19996 13861 20024 13892
rect 19981 13855 20039 13861
rect 19981 13821 19993 13855
rect 20027 13821 20039 13855
rect 19981 13815 20039 13821
rect 20346 13812 20352 13864
rect 20404 13812 20410 13864
rect 20640 13852 20668 13892
rect 20714 13880 20720 13932
rect 20772 13920 20778 13932
rect 21836 13929 21864 14028
rect 22094 14016 22100 14028
rect 22152 14016 22158 14068
rect 24765 14059 24823 14065
rect 24765 14025 24777 14059
rect 24811 14025 24823 14059
rect 24765 14019 24823 14025
rect 23198 13948 23204 14000
rect 23256 13988 23262 14000
rect 24780 13988 24808 14019
rect 23256 13960 24808 13988
rect 23256 13948 23262 13960
rect 24412 13929 24440 13960
rect 21269 13923 21327 13929
rect 21269 13920 21281 13923
rect 20772 13892 21281 13920
rect 20772 13880 20778 13892
rect 21269 13889 21281 13892
rect 21315 13889 21327 13923
rect 21269 13883 21327 13889
rect 21821 13923 21879 13929
rect 21821 13889 21833 13923
rect 21867 13889 21879 13923
rect 21821 13883 21879 13889
rect 24397 13923 24455 13929
rect 24397 13889 24409 13923
rect 24443 13889 24455 13923
rect 24397 13883 24455 13889
rect 20901 13855 20959 13861
rect 20640 13824 20852 13852
rect 18463 13756 18828 13784
rect 18463 13753 18475 13756
rect 18417 13747 18475 13753
rect 19058 13744 19064 13796
rect 19116 13784 19122 13796
rect 19797 13787 19855 13793
rect 19797 13784 19809 13787
rect 19116 13756 19809 13784
rect 19116 13744 19122 13756
rect 19797 13753 19809 13756
rect 19843 13753 19855 13787
rect 20824 13784 20852 13824
rect 20901 13821 20913 13855
rect 20947 13852 20959 13855
rect 21910 13852 21916 13864
rect 20947 13824 21916 13852
rect 20947 13821 20959 13824
rect 20901 13815 20959 13821
rect 21910 13812 21916 13824
rect 21968 13812 21974 13864
rect 23382 13812 23388 13864
rect 23440 13812 23446 13864
rect 23477 13855 23535 13861
rect 23477 13821 23489 13855
rect 23523 13852 23535 13855
rect 23750 13852 23756 13864
rect 23523 13824 23756 13852
rect 23523 13821 23535 13824
rect 23477 13815 23535 13821
rect 23750 13812 23756 13824
rect 23808 13852 23814 13864
rect 24765 13855 24823 13861
rect 24765 13852 24777 13855
rect 23808 13824 24777 13852
rect 23808 13812 23814 13824
rect 24765 13821 24777 13824
rect 24811 13821 24823 13855
rect 24765 13815 24823 13821
rect 24854 13812 24860 13864
rect 24912 13812 24918 13864
rect 25038 13812 25044 13864
rect 25096 13812 25102 13864
rect 25501 13855 25559 13861
rect 25501 13821 25513 13855
rect 25547 13852 25559 13855
rect 25590 13852 25596 13864
rect 25547 13824 25596 13852
rect 25547 13821 25559 13824
rect 25501 13815 25559 13821
rect 25590 13812 25596 13824
rect 25648 13812 25654 13864
rect 25774 13861 25780 13864
rect 25768 13852 25780 13861
rect 25735 13824 25780 13852
rect 25768 13815 25780 13824
rect 25774 13812 25780 13815
rect 25832 13812 25838 13864
rect 21266 13784 21272 13796
rect 20824 13756 21272 13784
rect 19797 13747 19855 13753
rect 21266 13744 21272 13756
rect 21324 13744 21330 13796
rect 22088 13787 22146 13793
rect 22088 13753 22100 13787
rect 22134 13784 22146 13787
rect 22186 13784 22192 13796
rect 22134 13756 22192 13784
rect 22134 13753 22146 13756
rect 22088 13747 22146 13753
rect 22186 13744 22192 13756
rect 22244 13744 22250 13796
rect 23400 13784 23428 13812
rect 23661 13787 23719 13793
rect 23661 13784 23673 13787
rect 23400 13756 23673 13784
rect 23661 13753 23673 13756
rect 23707 13784 23719 13787
rect 24394 13784 24400 13796
rect 23707 13756 24400 13784
rect 23707 13753 23719 13756
rect 23661 13747 23719 13753
rect 24394 13744 24400 13756
rect 24452 13744 24458 13796
rect 11882 13716 11888 13728
rect 11072 13688 11888 13716
rect 11882 13676 11888 13688
rect 11940 13676 11946 13728
rect 12434 13676 12440 13728
rect 12492 13716 12498 13728
rect 12894 13725 12900 13728
rect 12529 13719 12587 13725
rect 12529 13716 12541 13719
rect 12492 13688 12541 13716
rect 12492 13676 12498 13688
rect 12529 13685 12541 13688
rect 12575 13685 12587 13719
rect 12529 13679 12587 13685
rect 12881 13719 12900 13725
rect 12881 13685 12893 13719
rect 12881 13679 12900 13685
rect 12894 13676 12900 13679
rect 12952 13676 12958 13728
rect 15010 13676 15016 13728
rect 15068 13716 15074 13728
rect 15105 13719 15163 13725
rect 15105 13716 15117 13719
rect 15068 13688 15117 13716
rect 15068 13676 15074 13688
rect 15105 13685 15117 13688
rect 15151 13685 15163 13719
rect 15105 13679 15163 13685
rect 15194 13676 15200 13728
rect 15252 13716 15258 13728
rect 15447 13719 15505 13725
rect 15447 13716 15459 13719
rect 15252 13688 15459 13716
rect 15252 13676 15258 13688
rect 15447 13685 15459 13688
rect 15493 13685 15505 13719
rect 15447 13679 15505 13685
rect 16206 13676 16212 13728
rect 16264 13676 16270 13728
rect 16942 13676 16948 13728
rect 17000 13676 17006 13728
rect 18874 13676 18880 13728
rect 18932 13716 18938 13728
rect 19587 13719 19645 13725
rect 19587 13716 19599 13719
rect 18932 13688 19599 13716
rect 18932 13676 18938 13688
rect 19587 13685 19599 13688
rect 19633 13685 19645 13719
rect 19587 13679 19645 13685
rect 23290 13676 23296 13728
rect 23348 13676 23354 13728
rect 23566 13676 23572 13728
rect 23624 13716 23630 13728
rect 23845 13719 23903 13725
rect 23845 13716 23857 13719
rect 23624 13688 23857 13716
rect 23624 13676 23630 13688
rect 23845 13685 23857 13688
rect 23891 13685 23903 13719
rect 23845 13679 23903 13685
rect 24578 13676 24584 13728
rect 24636 13676 24642 13728
rect 26878 13676 26884 13728
rect 26936 13676 26942 13728
rect 552 13626 27576 13648
rect 552 13574 7114 13626
rect 7166 13574 7178 13626
rect 7230 13574 7242 13626
rect 7294 13574 7306 13626
rect 7358 13574 7370 13626
rect 7422 13574 13830 13626
rect 13882 13574 13894 13626
rect 13946 13574 13958 13626
rect 14010 13574 14022 13626
rect 14074 13574 14086 13626
rect 14138 13574 20546 13626
rect 20598 13574 20610 13626
rect 20662 13574 20674 13626
rect 20726 13574 20738 13626
rect 20790 13574 20802 13626
rect 20854 13574 27262 13626
rect 27314 13574 27326 13626
rect 27378 13574 27390 13626
rect 27442 13574 27454 13626
rect 27506 13574 27518 13626
rect 27570 13574 27576 13626
rect 552 13552 27576 13574
rect 1302 13472 1308 13524
rect 1360 13472 1366 13524
rect 3326 13472 3332 13524
rect 3384 13472 3390 13524
rect 3697 13515 3755 13521
rect 3697 13481 3709 13515
rect 3743 13512 3755 13515
rect 4154 13512 4160 13524
rect 3743 13484 4160 13512
rect 3743 13481 3755 13484
rect 3697 13475 3755 13481
rect 4154 13472 4160 13484
rect 4212 13472 4218 13524
rect 6089 13515 6147 13521
rect 6089 13481 6101 13515
rect 6135 13512 6147 13515
rect 6546 13512 6552 13524
rect 6135 13484 6552 13512
rect 6135 13481 6147 13484
rect 6089 13475 6147 13481
rect 6546 13472 6552 13484
rect 6604 13472 6610 13524
rect 7837 13515 7895 13521
rect 7837 13481 7849 13515
rect 7883 13481 7895 13515
rect 12434 13512 12440 13524
rect 7837 13475 7895 13481
rect 2685 13447 2743 13453
rect 2685 13413 2697 13447
rect 2731 13444 2743 13447
rect 2961 13447 3019 13453
rect 2961 13444 2973 13447
rect 2731 13416 2973 13444
rect 2731 13413 2743 13416
rect 2685 13407 2743 13413
rect 2961 13413 2973 13416
rect 3007 13413 3019 13447
rect 2961 13407 3019 13413
rect 3973 13447 4031 13453
rect 3973 13413 3985 13447
rect 4019 13444 4031 13447
rect 4402 13447 4460 13453
rect 4402 13444 4414 13447
rect 4019 13416 4414 13444
rect 4019 13413 4031 13416
rect 3973 13407 4031 13413
rect 4402 13413 4414 13416
rect 4448 13413 4460 13447
rect 6914 13444 6920 13456
rect 4402 13407 4460 13413
rect 6380 13416 6920 13444
rect 6380 13388 6408 13416
rect 6914 13404 6920 13416
rect 6972 13444 6978 13456
rect 7852 13444 7880 13475
rect 12406 13472 12440 13512
rect 12492 13512 12498 13524
rect 13446 13512 13452 13524
rect 12492 13484 13452 13512
rect 12492 13472 12498 13484
rect 13446 13472 13452 13484
rect 13504 13472 13510 13524
rect 14366 13521 14372 13524
rect 14093 13515 14151 13521
rect 14093 13481 14105 13515
rect 14139 13512 14151 13515
rect 14353 13515 14372 13521
rect 14353 13512 14365 13515
rect 14139 13484 14365 13512
rect 14139 13481 14151 13484
rect 14093 13475 14151 13481
rect 14353 13481 14365 13484
rect 14424 13512 14430 13524
rect 15102 13512 15108 13524
rect 14424 13484 15108 13512
rect 14353 13475 14372 13481
rect 14366 13472 14372 13475
rect 14424 13472 14430 13484
rect 15102 13472 15108 13484
rect 15160 13472 15166 13524
rect 18046 13472 18052 13524
rect 18104 13512 18110 13524
rect 18874 13521 18880 13524
rect 18693 13515 18751 13521
rect 18693 13512 18705 13515
rect 18104 13484 18705 13512
rect 18104 13472 18110 13484
rect 18693 13481 18705 13484
rect 18739 13481 18751 13515
rect 18693 13475 18751 13481
rect 18861 13515 18880 13521
rect 18861 13481 18873 13515
rect 18861 13475 18880 13481
rect 18874 13472 18880 13475
rect 18932 13472 18938 13524
rect 20809 13515 20867 13521
rect 20809 13481 20821 13515
rect 20855 13481 20867 13515
rect 20809 13475 20867 13481
rect 8386 13444 8392 13456
rect 6972 13416 7880 13444
rect 7944 13416 8392 13444
rect 6972 13404 6978 13416
rect 3142 13336 3148 13388
rect 3200 13336 3206 13388
rect 3418 13336 3424 13388
rect 3476 13336 3482 13388
rect 3513 13379 3571 13385
rect 3513 13345 3525 13379
rect 3559 13345 3571 13379
rect 3513 13339 3571 13345
rect 1854 13268 1860 13320
rect 1912 13268 1918 13320
rect 3528 13308 3556 13339
rect 3878 13336 3884 13388
rect 3936 13336 3942 13388
rect 4065 13379 4123 13385
rect 4065 13345 4077 13379
rect 4111 13376 4123 13379
rect 6178 13376 6184 13388
rect 4111 13348 6184 13376
rect 4111 13345 4123 13348
rect 4065 13339 4123 13345
rect 6178 13336 6184 13348
rect 6236 13336 6242 13388
rect 6270 13336 6276 13388
rect 6328 13336 6334 13388
rect 6362 13336 6368 13388
rect 6420 13336 6426 13388
rect 6730 13385 6736 13388
rect 6724 13376 6736 13385
rect 6691 13348 6736 13376
rect 6724 13339 6736 13348
rect 6730 13336 6736 13339
rect 6788 13336 6794 13388
rect 7944 13385 7972 13416
rect 8386 13404 8392 13416
rect 8444 13404 8450 13456
rect 9769 13447 9827 13453
rect 9769 13413 9781 13447
rect 9815 13444 9827 13447
rect 12406 13444 12434 13472
rect 9815 13416 12434 13444
rect 9815 13413 9827 13416
rect 9769 13407 9827 13413
rect 13354 13404 13360 13456
rect 13412 13444 13418 13456
rect 13725 13447 13783 13453
rect 13725 13444 13737 13447
rect 13412 13416 13737 13444
rect 13412 13404 13418 13416
rect 13725 13413 13737 13416
rect 13771 13413 13783 13447
rect 13725 13407 13783 13413
rect 13909 13447 13967 13453
rect 13909 13413 13921 13447
rect 13955 13444 13967 13447
rect 14182 13444 14188 13456
rect 13955 13416 14188 13444
rect 13955 13413 13967 13416
rect 13909 13407 13967 13413
rect 14182 13404 14188 13416
rect 14240 13404 14246 13456
rect 14550 13404 14556 13456
rect 14608 13404 14614 13456
rect 15841 13447 15899 13453
rect 15841 13413 15853 13447
rect 15887 13444 15899 13447
rect 16206 13444 16212 13456
rect 15887 13416 16212 13444
rect 15887 13413 15899 13416
rect 15841 13407 15899 13413
rect 16206 13404 16212 13416
rect 16264 13404 16270 13456
rect 16660 13447 16718 13453
rect 16660 13413 16672 13447
rect 16706 13444 16718 13447
rect 16942 13444 16948 13456
rect 16706 13416 16948 13444
rect 16706 13413 16718 13416
rect 16660 13407 16718 13413
rect 16942 13404 16948 13416
rect 17000 13404 17006 13456
rect 19058 13404 19064 13456
rect 19116 13404 19122 13456
rect 20472 13447 20530 13453
rect 20472 13413 20484 13447
rect 20518 13444 20530 13447
rect 20824 13444 20852 13475
rect 21266 13472 21272 13524
rect 21324 13472 21330 13524
rect 22005 13515 22063 13521
rect 22005 13481 22017 13515
rect 22051 13512 22063 13515
rect 22186 13512 22192 13524
rect 22051 13484 22192 13512
rect 22051 13481 22063 13484
rect 22005 13475 22063 13481
rect 22186 13472 22192 13484
rect 22244 13472 22250 13524
rect 25406 13512 25412 13524
rect 22940 13484 25412 13512
rect 21729 13447 21787 13453
rect 20518 13416 20852 13444
rect 20916 13416 21312 13444
rect 20518 13413 20530 13416
rect 20472 13407 20530 13413
rect 7929 13379 7987 13385
rect 7929 13345 7941 13379
rect 7975 13345 7987 13379
rect 7929 13339 7987 13345
rect 8196 13379 8254 13385
rect 8196 13345 8208 13379
rect 8242 13376 8254 13379
rect 9401 13379 9459 13385
rect 9401 13376 9413 13379
rect 8242 13348 9413 13376
rect 8242 13345 8254 13348
rect 8196 13339 8254 13345
rect 9401 13345 9413 13348
rect 9447 13345 9459 13379
rect 9401 13339 9459 13345
rect 9582 13336 9588 13388
rect 9640 13336 9646 13388
rect 9858 13336 9864 13388
rect 9916 13336 9922 13388
rect 9950 13336 9956 13388
rect 10008 13336 10014 13388
rect 10870 13336 10876 13388
rect 10928 13376 10934 13388
rect 10965 13379 11023 13385
rect 10965 13376 10977 13379
rect 10928 13348 10977 13376
rect 10928 13336 10934 13348
rect 10965 13345 10977 13348
rect 11011 13345 11023 13379
rect 10965 13339 11023 13345
rect 11149 13379 11207 13385
rect 11149 13345 11161 13379
rect 11195 13376 11207 13379
rect 11514 13376 11520 13388
rect 11195 13348 11520 13376
rect 11195 13345 11207 13348
rect 11149 13339 11207 13345
rect 11514 13336 11520 13348
rect 11572 13336 11578 13388
rect 15654 13336 15660 13388
rect 15712 13336 15718 13388
rect 15933 13379 15991 13385
rect 15933 13345 15945 13379
rect 15979 13376 15991 13379
rect 16022 13376 16028 13388
rect 15979 13348 16028 13376
rect 15979 13345 15991 13348
rect 15933 13339 15991 13345
rect 16022 13336 16028 13348
rect 16080 13336 16086 13388
rect 20916 13376 20944 13416
rect 19352 13348 20944 13376
rect 2884 13280 3556 13308
rect 4157 13311 4215 13317
rect 2314 13200 2320 13252
rect 2372 13200 2378 13252
rect 2884 13249 2912 13280
rect 4157 13277 4169 13311
rect 4203 13277 4215 13311
rect 4157 13271 4215 13277
rect 2869 13243 2927 13249
rect 2869 13209 2881 13243
rect 2915 13209 2927 13243
rect 2869 13203 2927 13209
rect 2682 13132 2688 13184
rect 2740 13132 2746 13184
rect 4172 13172 4200 13271
rect 5810 13268 5816 13320
rect 5868 13308 5874 13320
rect 6086 13308 6092 13320
rect 5868 13280 6092 13308
rect 5868 13268 5874 13280
rect 6086 13268 6092 13280
rect 6144 13268 6150 13320
rect 6457 13311 6515 13317
rect 6457 13277 6469 13311
rect 6503 13277 6515 13311
rect 6457 13271 6515 13277
rect 5350 13200 5356 13252
rect 5408 13240 5414 13252
rect 6472 13240 6500 13271
rect 13078 13268 13084 13320
rect 13136 13308 13142 13320
rect 13265 13311 13323 13317
rect 13265 13308 13277 13311
rect 13136 13280 13277 13308
rect 13136 13268 13142 13280
rect 13265 13277 13277 13280
rect 13311 13277 13323 13311
rect 13265 13271 13323 13277
rect 15378 13268 15384 13320
rect 15436 13268 15442 13320
rect 16390 13268 16396 13320
rect 16448 13268 16454 13320
rect 17957 13311 18015 13317
rect 17957 13308 17969 13311
rect 17788 13280 17969 13308
rect 5408 13212 6500 13240
rect 5408 13200 5414 13212
rect 8938 13200 8944 13252
rect 8996 13240 9002 13252
rect 15562 13240 15568 13252
rect 8996 13212 15568 13240
rect 8996 13200 9002 13212
rect 15562 13200 15568 13212
rect 15620 13200 15626 13252
rect 17678 13200 17684 13252
rect 17736 13240 17742 13252
rect 17788 13249 17816 13280
rect 17957 13277 17969 13280
rect 18003 13277 18015 13311
rect 19352 13308 19380 13348
rect 20990 13336 20996 13388
rect 21048 13336 21054 13388
rect 21284 13385 21312 13416
rect 21468 13416 21680 13444
rect 21468 13388 21496 13416
rect 21269 13379 21327 13385
rect 21269 13345 21281 13379
rect 21315 13345 21327 13379
rect 21269 13339 21327 13345
rect 21450 13336 21456 13388
rect 21508 13336 21514 13388
rect 21542 13336 21548 13388
rect 21600 13336 21606 13388
rect 21652 13376 21680 13416
rect 21729 13413 21741 13447
rect 21775 13444 21787 13447
rect 22738 13444 22744 13456
rect 21775 13416 22744 13444
rect 21775 13413 21787 13416
rect 21729 13407 21787 13413
rect 22738 13404 22744 13416
rect 22796 13404 22802 13456
rect 22462 13376 22468 13388
rect 21652 13348 22468 13376
rect 22462 13336 22468 13348
rect 22520 13336 22526 13388
rect 17957 13271 18015 13277
rect 18524 13280 19380 13308
rect 17773 13243 17831 13249
rect 17773 13240 17785 13243
rect 17736 13212 17785 13240
rect 17736 13200 17742 13212
rect 17773 13209 17785 13212
rect 17819 13209 17831 13243
rect 17773 13203 17831 13209
rect 4522 13172 4528 13184
rect 4172 13144 4528 13172
rect 4522 13132 4528 13144
rect 4580 13172 4586 13184
rect 5368 13172 5396 13200
rect 4580 13144 5396 13172
rect 4580 13132 4586 13144
rect 5442 13132 5448 13184
rect 5500 13172 5506 13184
rect 5537 13175 5595 13181
rect 5537 13172 5549 13175
rect 5500 13144 5549 13172
rect 5500 13132 5506 13144
rect 5537 13141 5549 13144
rect 5583 13141 5595 13175
rect 5537 13135 5595 13141
rect 9306 13132 9312 13184
rect 9364 13132 9370 13184
rect 10597 13175 10655 13181
rect 10597 13141 10609 13175
rect 10643 13172 10655 13175
rect 10870 13172 10876 13184
rect 10643 13144 10876 13172
rect 10643 13141 10655 13144
rect 10597 13135 10655 13141
rect 10870 13132 10876 13144
rect 10928 13132 10934 13184
rect 11149 13175 11207 13181
rect 11149 13141 11161 13175
rect 11195 13172 11207 13175
rect 11330 13172 11336 13184
rect 11195 13144 11336 13172
rect 11195 13141 11207 13144
rect 11149 13135 11207 13141
rect 11330 13132 11336 13144
rect 11388 13132 11394 13184
rect 12713 13175 12771 13181
rect 12713 13141 12725 13175
rect 12759 13172 12771 13175
rect 12802 13172 12808 13184
rect 12759 13144 12808 13172
rect 12759 13141 12771 13144
rect 12713 13135 12771 13141
rect 12802 13132 12808 13144
rect 12860 13132 12866 13184
rect 14185 13175 14243 13181
rect 14185 13141 14197 13175
rect 14231 13172 14243 13175
rect 14274 13172 14280 13184
rect 14231 13144 14280 13172
rect 14231 13141 14243 13144
rect 14185 13135 14243 13141
rect 14274 13132 14280 13144
rect 14332 13132 14338 13184
rect 14369 13175 14427 13181
rect 14369 13141 14381 13175
rect 14415 13172 14427 13175
rect 14737 13175 14795 13181
rect 14737 13172 14749 13175
rect 14415 13144 14749 13172
rect 14415 13141 14427 13144
rect 14369 13135 14427 13141
rect 14737 13141 14749 13144
rect 14783 13141 14795 13175
rect 14737 13135 14795 13141
rect 15470 13132 15476 13184
rect 15528 13132 15534 13184
rect 17586 13132 17592 13184
rect 17644 13172 17650 13184
rect 18524 13172 18552 13280
rect 19352 13252 19380 13280
rect 20714 13268 20720 13320
rect 20772 13308 20778 13320
rect 22094 13308 22100 13320
rect 20772 13280 22100 13308
rect 20772 13268 20778 13280
rect 22094 13268 22100 13280
rect 22152 13268 22158 13320
rect 22649 13311 22707 13317
rect 22649 13277 22661 13311
rect 22695 13308 22707 13311
rect 22741 13311 22799 13317
rect 22741 13308 22753 13311
rect 22695 13280 22753 13308
rect 22695 13277 22707 13280
rect 22649 13271 22707 13277
rect 22741 13277 22753 13280
rect 22787 13277 22799 13311
rect 22741 13271 22799 13277
rect 18601 13243 18659 13249
rect 18601 13209 18613 13243
rect 18647 13240 18659 13243
rect 18647 13212 18920 13240
rect 18647 13209 18659 13212
rect 18601 13203 18659 13209
rect 18892 13181 18920 13212
rect 19334 13200 19340 13252
rect 19392 13200 19398 13252
rect 21913 13243 21971 13249
rect 21913 13209 21925 13243
rect 21959 13240 21971 13243
rect 22940 13240 22968 13484
rect 25406 13472 25412 13484
rect 25464 13472 25470 13524
rect 26421 13515 26479 13521
rect 26421 13481 26433 13515
rect 26467 13512 26479 13515
rect 26602 13512 26608 13524
rect 26467 13484 26608 13512
rect 26467 13481 26479 13484
rect 26421 13475 26479 13481
rect 26602 13472 26608 13484
rect 26660 13472 26666 13524
rect 23566 13444 23572 13456
rect 23032 13416 23572 13444
rect 23032 13385 23060 13416
rect 23566 13404 23572 13416
rect 23624 13404 23630 13456
rect 24946 13444 24952 13456
rect 23768 13416 24952 13444
rect 23017 13379 23075 13385
rect 23017 13345 23029 13379
rect 23063 13345 23075 13379
rect 23017 13339 23075 13345
rect 23109 13379 23167 13385
rect 23109 13345 23121 13379
rect 23155 13345 23167 13379
rect 23109 13339 23167 13345
rect 23201 13379 23259 13385
rect 23201 13345 23213 13379
rect 23247 13376 23259 13379
rect 23290 13376 23296 13388
rect 23247 13348 23296 13376
rect 23247 13345 23259 13348
rect 23201 13339 23259 13345
rect 21959 13212 22968 13240
rect 21959 13209 21971 13212
rect 21913 13203 21971 13209
rect 23014 13200 23020 13252
rect 23072 13240 23078 13252
rect 23124 13240 23152 13339
rect 23290 13336 23296 13348
rect 23348 13336 23354 13388
rect 23768 13385 23796 13416
rect 24946 13404 24952 13416
rect 25004 13444 25010 13456
rect 25682 13444 25688 13456
rect 25004 13416 25688 13444
rect 25004 13404 25010 13416
rect 25682 13404 25688 13416
rect 25740 13404 25746 13456
rect 25884 13416 26924 13444
rect 25884 13385 25912 13416
rect 26896 13388 26924 13416
rect 23385 13379 23443 13385
rect 23385 13345 23397 13379
rect 23431 13376 23443 13379
rect 23477 13379 23535 13385
rect 23477 13376 23489 13379
rect 23431 13348 23489 13376
rect 23431 13345 23443 13348
rect 23385 13339 23443 13345
rect 23477 13345 23489 13348
rect 23523 13345 23535 13379
rect 23477 13339 23535 13345
rect 23661 13379 23719 13385
rect 23661 13345 23673 13379
rect 23707 13345 23719 13379
rect 23661 13339 23719 13345
rect 23753 13379 23811 13385
rect 23753 13345 23765 13379
rect 23799 13345 23811 13379
rect 23753 13339 23811 13345
rect 23845 13379 23903 13385
rect 23845 13345 23857 13379
rect 23891 13376 23903 13379
rect 25869 13379 25927 13385
rect 23891 13348 24072 13376
rect 23891 13345 23903 13348
rect 23845 13339 23903 13345
rect 23400 13308 23428 13339
rect 23308 13280 23428 13308
rect 23308 13252 23336 13280
rect 23072 13212 23152 13240
rect 23072 13200 23078 13212
rect 17644 13144 18552 13172
rect 18877 13175 18935 13181
rect 17644 13132 17650 13144
rect 18877 13141 18889 13175
rect 18923 13141 18935 13175
rect 23124 13172 23152 13212
rect 23290 13200 23296 13252
rect 23348 13200 23354 13252
rect 23382 13200 23388 13252
rect 23440 13240 23446 13252
rect 23676 13240 23704 13339
rect 23440 13212 23704 13240
rect 23440 13200 23446 13212
rect 23768 13172 23796 13339
rect 23124 13144 23796 13172
rect 24044 13172 24072 13348
rect 25869 13345 25881 13379
rect 25915 13345 25927 13379
rect 25869 13339 25927 13345
rect 26145 13379 26203 13385
rect 26145 13345 26157 13379
rect 26191 13376 26203 13379
rect 26602 13376 26608 13388
rect 26191 13348 26608 13376
rect 26191 13345 26203 13348
rect 26145 13339 26203 13345
rect 26602 13336 26608 13348
rect 26660 13336 26666 13388
rect 26878 13336 26884 13388
rect 26936 13376 26942 13388
rect 26973 13379 27031 13385
rect 26973 13376 26985 13379
rect 26936 13348 26985 13376
rect 26936 13336 26942 13348
rect 26973 13345 26985 13348
rect 27019 13345 27031 13379
rect 26973 13339 27031 13345
rect 24854 13268 24860 13320
rect 24912 13268 24918 13320
rect 25501 13311 25559 13317
rect 25501 13277 25513 13311
rect 25547 13277 25559 13311
rect 25501 13271 25559 13277
rect 26053 13311 26111 13317
rect 26053 13277 26065 13311
rect 26099 13308 26111 13311
rect 27062 13308 27068 13320
rect 26099 13280 27068 13308
rect 26099 13277 26111 13280
rect 26053 13271 26111 13277
rect 24121 13243 24179 13249
rect 24121 13209 24133 13243
rect 24167 13240 24179 13243
rect 25516 13240 25544 13271
rect 27062 13268 27068 13280
rect 27120 13268 27126 13320
rect 24167 13212 25544 13240
rect 24167 13209 24179 13212
rect 24121 13203 24179 13209
rect 24213 13175 24271 13181
rect 24213 13172 24225 13175
rect 24044 13144 24225 13172
rect 18877 13135 18935 13141
rect 24213 13141 24225 13144
rect 24259 13172 24271 13175
rect 24302 13172 24308 13184
rect 24259 13144 24308 13172
rect 24259 13141 24271 13144
rect 24213 13135 24271 13141
rect 24302 13132 24308 13144
rect 24360 13132 24366 13184
rect 24946 13132 24952 13184
rect 25004 13132 25010 13184
rect 25038 13132 25044 13184
rect 25096 13172 25102 13184
rect 25685 13175 25743 13181
rect 25685 13172 25697 13175
rect 25096 13144 25697 13172
rect 25096 13132 25102 13144
rect 25685 13141 25697 13144
rect 25731 13141 25743 13175
rect 25685 13135 25743 13141
rect 26145 13175 26203 13181
rect 26145 13141 26157 13175
rect 26191 13172 26203 13175
rect 26234 13172 26240 13184
rect 26191 13144 26240 13172
rect 26191 13141 26203 13144
rect 26145 13135 26203 13141
rect 26234 13132 26240 13144
rect 26292 13132 26298 13184
rect 552 13082 27416 13104
rect 552 13030 3756 13082
rect 3808 13030 3820 13082
rect 3872 13030 3884 13082
rect 3936 13030 3948 13082
rect 4000 13030 4012 13082
rect 4064 13030 10472 13082
rect 10524 13030 10536 13082
rect 10588 13030 10600 13082
rect 10652 13030 10664 13082
rect 10716 13030 10728 13082
rect 10780 13030 17188 13082
rect 17240 13030 17252 13082
rect 17304 13030 17316 13082
rect 17368 13030 17380 13082
rect 17432 13030 17444 13082
rect 17496 13030 23904 13082
rect 23956 13030 23968 13082
rect 24020 13030 24032 13082
rect 24084 13030 24096 13082
rect 24148 13030 24160 13082
rect 24212 13030 27416 13082
rect 552 13008 27416 13030
rect 1397 12971 1455 12977
rect 1397 12937 1409 12971
rect 1443 12968 1455 12971
rect 1854 12968 1860 12980
rect 1443 12940 1860 12968
rect 1443 12937 1455 12940
rect 1397 12931 1455 12937
rect 1854 12928 1860 12940
rect 1912 12928 1918 12980
rect 4522 12928 4528 12980
rect 4580 12968 4586 12980
rect 4801 12971 4859 12977
rect 4801 12968 4813 12971
rect 4580 12940 4813 12968
rect 4580 12928 4586 12940
rect 4801 12937 4813 12940
rect 4847 12937 4859 12971
rect 4801 12931 4859 12937
rect 1670 12860 1676 12912
rect 1728 12900 1734 12912
rect 1949 12903 2007 12909
rect 1949 12900 1961 12903
rect 1728 12872 1961 12900
rect 1728 12860 1734 12872
rect 1949 12869 1961 12872
rect 1995 12869 2007 12903
rect 1949 12863 2007 12869
rect 2038 12860 2044 12912
rect 2096 12900 2102 12912
rect 2958 12900 2964 12912
rect 2096 12872 2964 12900
rect 2096 12860 2102 12872
rect 2958 12860 2964 12872
rect 3016 12860 3022 12912
rect 3694 12900 3700 12912
rect 3436 12872 3700 12900
rect 1762 12792 1768 12844
rect 1820 12792 1826 12844
rect 1854 12792 1860 12844
rect 1912 12792 1918 12844
rect 1578 12724 1584 12776
rect 1636 12724 1642 12776
rect 1949 12767 2007 12773
rect 1949 12733 1961 12767
rect 1995 12764 2007 12767
rect 2056 12764 2084 12860
rect 1995 12736 2084 12764
rect 2225 12767 2283 12773
rect 1995 12733 2007 12736
rect 1949 12727 2007 12733
rect 2225 12733 2237 12767
rect 2271 12764 2283 12767
rect 2314 12764 2320 12776
rect 2271 12736 2320 12764
rect 2271 12733 2283 12736
rect 2225 12727 2283 12733
rect 2314 12724 2320 12736
rect 2372 12724 2378 12776
rect 2774 12724 2780 12776
rect 2832 12724 2838 12776
rect 3436 12773 3464 12872
rect 3694 12860 3700 12872
rect 3752 12900 3758 12912
rect 4816 12900 4844 12931
rect 5166 12928 5172 12980
rect 5224 12968 5230 12980
rect 6733 12971 6791 12977
rect 5224 12940 5764 12968
rect 5224 12928 5230 12940
rect 5442 12900 5448 12912
rect 3752 12872 4660 12900
rect 4816 12872 5448 12900
rect 3752 12860 3758 12872
rect 4522 12792 4528 12844
rect 4580 12792 4586 12844
rect 4632 12832 4660 12872
rect 5442 12860 5448 12872
rect 5500 12900 5506 12912
rect 5736 12900 5764 12940
rect 6733 12937 6745 12971
rect 6779 12968 6791 12971
rect 6822 12968 6828 12980
rect 6779 12940 6828 12968
rect 6779 12937 6791 12940
rect 6733 12931 6791 12937
rect 6822 12928 6828 12940
rect 6880 12928 6886 12980
rect 8941 12971 8999 12977
rect 8941 12937 8953 12971
rect 8987 12968 8999 12971
rect 9217 12971 9275 12977
rect 9217 12968 9229 12971
rect 8987 12940 9229 12968
rect 8987 12937 8999 12940
rect 8941 12931 8999 12937
rect 9217 12937 9229 12940
rect 9263 12937 9275 12971
rect 9217 12931 9275 12937
rect 10318 12928 10324 12980
rect 10376 12968 10382 12980
rect 10413 12971 10471 12977
rect 10413 12968 10425 12971
rect 10376 12940 10425 12968
rect 10376 12928 10382 12940
rect 10413 12937 10425 12940
rect 10459 12937 10471 12971
rect 10413 12931 10471 12937
rect 10689 12971 10747 12977
rect 10689 12937 10701 12971
rect 10735 12968 10747 12971
rect 10870 12968 10876 12980
rect 10735 12940 10876 12968
rect 10735 12937 10747 12940
rect 10689 12931 10747 12937
rect 10870 12928 10876 12940
rect 10928 12928 10934 12980
rect 12158 12928 12164 12980
rect 12216 12968 12222 12980
rect 12618 12968 12624 12980
rect 12216 12940 12624 12968
rect 12216 12928 12222 12940
rect 12618 12928 12624 12940
rect 12676 12928 12682 12980
rect 12802 12928 12808 12980
rect 12860 12928 12866 12980
rect 15562 12928 15568 12980
rect 15620 12968 15626 12980
rect 16577 12971 16635 12977
rect 15620 12940 16160 12968
rect 15620 12928 15626 12940
rect 6917 12903 6975 12909
rect 6917 12900 6929 12903
rect 5500 12872 5580 12900
rect 5736 12872 6929 12900
rect 5500 12860 5506 12872
rect 5552 12841 5580 12872
rect 6917 12869 6929 12872
rect 6963 12869 6975 12903
rect 6917 12863 6975 12869
rect 9125 12903 9183 12909
rect 9125 12869 9137 12903
rect 9171 12900 9183 12903
rect 9582 12900 9588 12912
rect 9171 12872 9588 12900
rect 9171 12869 9183 12872
rect 9125 12863 9183 12869
rect 9582 12860 9588 12872
rect 9640 12860 9646 12912
rect 9674 12860 9680 12912
rect 9732 12900 9738 12912
rect 10042 12900 10048 12912
rect 9732 12872 10048 12900
rect 9732 12860 9738 12872
rect 10042 12860 10048 12872
rect 10100 12900 10106 12912
rect 10778 12900 10784 12912
rect 10100 12872 10784 12900
rect 10100 12860 10106 12872
rect 10778 12860 10784 12872
rect 10836 12860 10842 12912
rect 12529 12903 12587 12909
rect 12529 12869 12541 12903
rect 12575 12900 12587 12903
rect 13078 12900 13084 12912
rect 12575 12872 13084 12900
rect 12575 12869 12587 12872
rect 12529 12863 12587 12869
rect 13078 12860 13084 12872
rect 13136 12860 13142 12912
rect 16132 12900 16160 12940
rect 16577 12937 16589 12971
rect 16623 12968 16635 12971
rect 16758 12968 16764 12980
rect 16623 12940 16764 12968
rect 16623 12937 16635 12940
rect 16577 12931 16635 12937
rect 16758 12928 16764 12940
rect 16816 12968 16822 12980
rect 17034 12968 17040 12980
rect 16816 12940 17040 12968
rect 16816 12928 16822 12940
rect 17034 12928 17040 12940
rect 17092 12928 17098 12980
rect 17144 12940 19656 12968
rect 17144 12900 17172 12940
rect 16132 12872 17172 12900
rect 19628 12900 19656 12940
rect 20346 12928 20352 12980
rect 20404 12928 20410 12980
rect 20456 12940 21772 12968
rect 20456 12900 20484 12940
rect 19628 12872 20484 12900
rect 4893 12835 4951 12841
rect 4893 12832 4905 12835
rect 4632 12804 4905 12832
rect 4893 12801 4905 12804
rect 4939 12801 4951 12835
rect 4893 12795 4951 12801
rect 5537 12835 5595 12841
rect 5537 12801 5549 12835
rect 5583 12801 5595 12835
rect 5537 12795 5595 12801
rect 6181 12835 6239 12841
rect 6181 12801 6193 12835
rect 6227 12832 6239 12835
rect 7101 12835 7159 12841
rect 6227 12804 6868 12832
rect 6227 12801 6239 12804
rect 6181 12795 6239 12801
rect 3421 12767 3479 12773
rect 3421 12733 3433 12767
rect 3467 12733 3479 12767
rect 3697 12767 3755 12773
rect 3697 12764 3709 12767
rect 3421 12727 3479 12733
rect 3528 12736 3709 12764
rect 2332 12696 2360 12724
rect 2866 12696 2872 12708
rect 2332 12668 2872 12696
rect 2866 12656 2872 12668
rect 2924 12696 2930 12708
rect 3528 12696 3556 12736
rect 3697 12733 3709 12736
rect 3743 12733 3755 12767
rect 3697 12727 3755 12733
rect 4338 12724 4344 12776
rect 4396 12724 4402 12776
rect 4433 12767 4491 12773
rect 4433 12733 4445 12767
rect 4479 12733 4491 12767
rect 4433 12727 4491 12733
rect 4617 12767 4675 12773
rect 4617 12733 4629 12767
rect 4663 12764 4675 12767
rect 4706 12764 4712 12776
rect 4663 12736 4712 12764
rect 4663 12733 4675 12736
rect 4617 12727 4675 12733
rect 2924 12668 3556 12696
rect 2924 12656 2930 12668
rect 3602 12656 3608 12708
rect 3660 12696 3666 12708
rect 4448 12696 4476 12727
rect 4706 12724 4712 12736
rect 4764 12724 4770 12776
rect 5077 12767 5135 12773
rect 5077 12733 5089 12767
rect 5123 12733 5135 12767
rect 5077 12727 5135 12733
rect 4798 12696 4804 12708
rect 3660 12668 4384 12696
rect 4448 12668 4804 12696
rect 3660 12656 3666 12668
rect 2133 12631 2191 12637
rect 2133 12597 2145 12631
rect 2179 12628 2191 12631
rect 2222 12628 2228 12640
rect 2179 12600 2228 12628
rect 2179 12597 2191 12600
rect 2133 12591 2191 12597
rect 2222 12588 2228 12600
rect 2280 12588 2286 12640
rect 2590 12588 2596 12640
rect 2648 12588 2654 12640
rect 3234 12588 3240 12640
rect 3292 12588 3298 12640
rect 4157 12631 4215 12637
rect 4157 12597 4169 12631
rect 4203 12628 4215 12631
rect 4246 12628 4252 12640
rect 4203 12600 4252 12628
rect 4203 12597 4215 12600
rect 4157 12591 4215 12597
rect 4246 12588 4252 12600
rect 4304 12588 4310 12640
rect 4356 12628 4384 12668
rect 4798 12656 4804 12668
rect 4856 12656 4862 12708
rect 5092 12628 5120 12727
rect 6362 12724 6368 12776
rect 6420 12724 6426 12776
rect 6546 12724 6552 12776
rect 6604 12724 6610 12776
rect 6840 12773 6868 12804
rect 7101 12801 7113 12835
rect 7147 12832 7159 12835
rect 8938 12832 8944 12844
rect 7147 12804 8944 12832
rect 7147 12801 7159 12804
rect 7101 12795 7159 12801
rect 8938 12792 8944 12804
rect 8996 12792 9002 12844
rect 9306 12792 9312 12844
rect 9364 12832 9370 12844
rect 9490 12832 9496 12844
rect 9364 12804 9496 12832
rect 9364 12792 9370 12804
rect 9490 12792 9496 12804
rect 9548 12832 9554 12844
rect 9769 12835 9827 12841
rect 9769 12832 9781 12835
rect 9548 12804 9781 12832
rect 9548 12792 9554 12804
rect 9769 12801 9781 12804
rect 9815 12801 9827 12835
rect 9769 12795 9827 12801
rect 9858 12792 9864 12844
rect 9916 12832 9922 12844
rect 9916 12804 11008 12832
rect 9916 12792 9922 12804
rect 9968 12773 9996 12804
rect 6825 12767 6883 12773
rect 6825 12733 6837 12767
rect 6871 12733 6883 12767
rect 6825 12727 6883 12733
rect 9953 12767 10011 12773
rect 9953 12733 9965 12767
rect 9999 12764 10011 12767
rect 10229 12767 10287 12773
rect 9999 12736 10033 12764
rect 9999 12733 10011 12736
rect 9953 12727 10011 12733
rect 10229 12733 10241 12767
rect 10275 12764 10287 12767
rect 10275 12736 10548 12764
rect 10275 12733 10287 12736
rect 10229 12727 10287 12733
rect 8757 12699 8815 12705
rect 8757 12665 8769 12699
rect 8803 12696 8815 12699
rect 8846 12696 8852 12708
rect 8803 12668 8852 12696
rect 8803 12665 8815 12668
rect 8757 12659 8815 12665
rect 8846 12656 8852 12668
rect 8904 12696 8910 12708
rect 9674 12696 9680 12708
rect 8904 12668 9680 12696
rect 8904 12656 8910 12668
rect 9674 12656 9680 12668
rect 9732 12656 9738 12708
rect 4356 12600 5120 12628
rect 5261 12631 5319 12637
rect 5261 12597 5273 12631
rect 5307 12628 5319 12631
rect 5994 12628 6000 12640
rect 5307 12600 6000 12628
rect 5307 12597 5319 12600
rect 5261 12591 5319 12597
rect 5994 12588 6000 12600
rect 6052 12588 6058 12640
rect 6178 12588 6184 12640
rect 6236 12628 6242 12640
rect 7101 12631 7159 12637
rect 7101 12628 7113 12631
rect 6236 12600 7113 12628
rect 6236 12588 6242 12600
rect 7101 12597 7113 12600
rect 7147 12597 7159 12631
rect 7101 12591 7159 12597
rect 8967 12631 9025 12637
rect 8967 12597 8979 12631
rect 9013 12628 9025 12631
rect 9766 12628 9772 12640
rect 9013 12600 9772 12628
rect 9013 12597 9025 12600
rect 8967 12591 9025 12597
rect 9766 12588 9772 12600
rect 9824 12588 9830 12640
rect 10045 12631 10103 12637
rect 10045 12597 10057 12631
rect 10091 12628 10103 12631
rect 10318 12628 10324 12640
rect 10091 12600 10324 12628
rect 10091 12597 10103 12600
rect 10045 12591 10103 12597
rect 10318 12588 10324 12600
rect 10376 12588 10382 12640
rect 10520 12637 10548 12736
rect 10778 12656 10784 12708
rect 10836 12696 10842 12708
rect 10873 12699 10931 12705
rect 10873 12696 10885 12699
rect 10836 12668 10885 12696
rect 10836 12656 10842 12668
rect 10873 12665 10885 12668
rect 10919 12665 10931 12699
rect 10980 12696 11008 12804
rect 12167 12804 13584 12832
rect 11149 12767 11207 12773
rect 11149 12733 11161 12767
rect 11195 12764 11207 12767
rect 11882 12764 11888 12776
rect 11195 12736 11888 12764
rect 11195 12733 11207 12736
rect 11149 12727 11207 12733
rect 11882 12724 11888 12736
rect 11940 12764 11946 12776
rect 12167 12764 12195 12804
rect 11940 12736 12195 12764
rect 11940 12724 11946 12736
rect 13078 12724 13084 12776
rect 13136 12724 13142 12776
rect 13265 12767 13323 12773
rect 13265 12733 13277 12767
rect 13311 12764 13323 12767
rect 13446 12764 13452 12776
rect 13311 12736 13452 12764
rect 13311 12733 13323 12736
rect 13265 12727 13323 12733
rect 13446 12724 13452 12736
rect 13504 12724 13510 12776
rect 13556 12773 13584 12804
rect 16390 12792 16396 12844
rect 16448 12832 16454 12844
rect 18693 12835 18751 12841
rect 18693 12832 18705 12835
rect 16448 12804 18705 12832
rect 16448 12792 16454 12804
rect 18693 12801 18705 12804
rect 18739 12801 18751 12835
rect 18693 12795 18751 12801
rect 20714 12792 20720 12844
rect 20772 12792 20778 12844
rect 21744 12832 21772 12940
rect 22830 12928 22836 12980
rect 22888 12968 22894 12980
rect 23014 12968 23020 12980
rect 22888 12940 23020 12968
rect 22888 12928 22894 12940
rect 23014 12928 23020 12940
rect 23072 12928 23078 12980
rect 23845 12971 23903 12977
rect 23845 12937 23857 12971
rect 23891 12968 23903 12971
rect 24854 12968 24860 12980
rect 23891 12940 24860 12968
rect 23891 12937 23903 12940
rect 23845 12931 23903 12937
rect 24854 12928 24860 12940
rect 24912 12928 24918 12980
rect 27062 12928 27068 12980
rect 27120 12928 27126 12980
rect 22097 12903 22155 12909
rect 22097 12869 22109 12903
rect 22143 12900 22155 12903
rect 23750 12900 23756 12912
rect 22143 12872 23756 12900
rect 22143 12869 22155 12872
rect 22097 12863 22155 12869
rect 22646 12832 22652 12844
rect 21744 12804 22652 12832
rect 13541 12767 13599 12773
rect 13541 12733 13553 12767
rect 13587 12764 13599 12767
rect 14642 12764 14648 12776
rect 13587 12736 14648 12764
rect 13587 12733 13599 12736
rect 13541 12727 13599 12733
rect 14642 12724 14648 12736
rect 14700 12764 14706 12776
rect 15197 12767 15255 12773
rect 15197 12764 15209 12767
rect 14700 12736 15209 12764
rect 14700 12724 14706 12736
rect 15197 12733 15209 12736
rect 15243 12764 15255 12767
rect 16408 12764 16436 12792
rect 15243 12736 16436 12764
rect 15243 12733 15255 12736
rect 15197 12727 15255 12733
rect 17586 12724 17592 12776
rect 17644 12724 17650 12776
rect 17678 12724 17684 12776
rect 17736 12724 17742 12776
rect 18509 12767 18567 12773
rect 18509 12733 18521 12767
rect 18555 12764 18567 12767
rect 18598 12764 18604 12776
rect 18555 12736 18604 12764
rect 18555 12733 18567 12736
rect 18509 12727 18567 12733
rect 18598 12724 18604 12736
rect 18656 12724 18662 12776
rect 19334 12724 19340 12776
rect 19392 12764 19398 12776
rect 20165 12767 20223 12773
rect 20165 12764 20177 12767
rect 19392 12736 20177 12764
rect 19392 12724 19398 12736
rect 20165 12733 20177 12736
rect 20211 12733 20223 12767
rect 20165 12727 20223 12733
rect 20349 12767 20407 12773
rect 20349 12733 20361 12767
rect 20395 12764 20407 12767
rect 21450 12764 21456 12776
rect 20395 12736 21456 12764
rect 20395 12733 20407 12736
rect 20349 12727 20407 12733
rect 21450 12724 21456 12736
rect 21508 12724 21514 12776
rect 21818 12724 21824 12776
rect 21876 12764 21882 12776
rect 22480 12773 22508 12804
rect 22646 12792 22652 12804
rect 22704 12832 22710 12844
rect 23290 12832 23296 12844
rect 22704 12804 23296 12832
rect 22704 12792 22710 12804
rect 23290 12792 23296 12804
rect 23348 12792 23354 12844
rect 23584 12841 23612 12872
rect 23750 12860 23756 12872
rect 23808 12860 23814 12912
rect 23569 12835 23627 12841
rect 23569 12801 23581 12835
rect 23615 12801 23627 12835
rect 23569 12795 23627 12801
rect 25225 12835 25283 12841
rect 25225 12801 25237 12835
rect 25271 12832 25283 12835
rect 25590 12832 25596 12844
rect 25271 12804 25596 12832
rect 25271 12801 25283 12804
rect 25225 12795 25283 12801
rect 25590 12792 25596 12804
rect 25648 12832 25654 12844
rect 25685 12835 25743 12841
rect 25685 12832 25697 12835
rect 25648 12804 25697 12832
rect 25648 12792 25654 12804
rect 25685 12801 25697 12804
rect 25731 12801 25743 12835
rect 25685 12795 25743 12801
rect 22465 12767 22523 12773
rect 21876 12736 22324 12764
rect 21876 12724 21882 12736
rect 11416 12699 11474 12705
rect 10980 12668 11376 12696
rect 10873 12659 10931 12665
rect 11348 12640 11376 12668
rect 11416 12665 11428 12699
rect 11462 12696 11474 12699
rect 11514 12696 11520 12708
rect 11462 12668 11520 12696
rect 11462 12665 11474 12668
rect 11416 12659 11474 12665
rect 11514 12656 11520 12668
rect 11572 12656 11578 12708
rect 12434 12656 12440 12708
rect 12492 12696 12498 12708
rect 12773 12699 12831 12705
rect 12773 12696 12785 12699
rect 12492 12668 12785 12696
rect 12492 12656 12498 12668
rect 12773 12665 12785 12668
rect 12819 12696 12831 12699
rect 12894 12696 12900 12708
rect 12819 12668 12900 12696
rect 12819 12665 12831 12668
rect 12773 12659 12831 12665
rect 12894 12656 12900 12668
rect 12952 12656 12958 12708
rect 12986 12656 12992 12708
rect 13044 12656 13050 12708
rect 13808 12699 13866 12705
rect 13808 12665 13820 12699
rect 13854 12696 13866 12699
rect 14182 12696 14188 12708
rect 13854 12668 14188 12696
rect 13854 12665 13866 12668
rect 13808 12659 13866 12665
rect 14182 12656 14188 12668
rect 14240 12656 14246 12708
rect 15470 12705 15476 12708
rect 15464 12696 15476 12705
rect 15431 12668 15476 12696
rect 15464 12659 15476 12668
rect 15470 12656 15476 12659
rect 15528 12656 15534 12708
rect 16114 12696 16120 12708
rect 15580 12668 16120 12696
rect 10505 12631 10563 12637
rect 10505 12597 10517 12631
rect 10551 12597 10563 12631
rect 10505 12591 10563 12597
rect 10673 12631 10731 12637
rect 10673 12597 10685 12631
rect 10719 12628 10731 12631
rect 10962 12628 10968 12640
rect 10719 12600 10968 12628
rect 10719 12597 10731 12600
rect 10673 12591 10731 12597
rect 10962 12588 10968 12600
rect 11020 12588 11026 12640
rect 11330 12588 11336 12640
rect 11388 12588 11394 12640
rect 11698 12588 11704 12640
rect 11756 12628 11762 12640
rect 12621 12631 12679 12637
rect 12621 12628 12633 12631
rect 11756 12600 12633 12628
rect 11756 12588 11762 12600
rect 12621 12597 12633 12600
rect 12667 12597 12679 12631
rect 12621 12591 12679 12597
rect 13078 12588 13084 12640
rect 13136 12628 13142 12640
rect 13173 12631 13231 12637
rect 13173 12628 13185 12631
rect 13136 12600 13185 12628
rect 13136 12588 13142 12600
rect 13173 12597 13185 12600
rect 13219 12597 13231 12631
rect 13173 12591 13231 12597
rect 14921 12631 14979 12637
rect 14921 12597 14933 12631
rect 14967 12628 14979 12631
rect 15378 12628 15384 12640
rect 14967 12600 15384 12628
rect 14967 12597 14979 12600
rect 14921 12591 14979 12597
rect 15378 12588 15384 12600
rect 15436 12628 15442 12640
rect 15580 12628 15608 12668
rect 16114 12656 16120 12668
rect 16172 12656 16178 12708
rect 17954 12656 17960 12708
rect 18012 12656 18018 12708
rect 18049 12699 18107 12705
rect 18049 12665 18061 12699
rect 18095 12696 18107 12699
rect 18417 12699 18475 12705
rect 18417 12696 18429 12699
rect 18095 12668 18429 12696
rect 18095 12665 18107 12668
rect 18049 12659 18107 12665
rect 18417 12665 18429 12668
rect 18463 12665 18475 12699
rect 18417 12659 18475 12665
rect 18960 12699 19018 12705
rect 18960 12665 18972 12699
rect 19006 12696 19018 12699
rect 19242 12696 19248 12708
rect 19006 12668 19248 12696
rect 19006 12665 19018 12668
rect 18960 12659 19018 12665
rect 19242 12656 19248 12668
rect 19300 12656 19306 12708
rect 20984 12699 21042 12705
rect 20984 12665 20996 12699
rect 21030 12696 21042 12699
rect 22189 12699 22247 12705
rect 22189 12696 22201 12699
rect 21030 12668 22201 12696
rect 21030 12665 21042 12668
rect 20984 12659 21042 12665
rect 22189 12665 22201 12668
rect 22235 12665 22247 12699
rect 22296 12696 22324 12736
rect 22465 12733 22477 12767
rect 22511 12733 22523 12767
rect 22465 12727 22523 12733
rect 22925 12767 22983 12773
rect 22925 12733 22937 12767
rect 22971 12764 22983 12767
rect 23017 12767 23075 12773
rect 23017 12764 23029 12767
rect 22971 12736 23029 12764
rect 22971 12733 22983 12736
rect 22925 12727 22983 12733
rect 23017 12733 23029 12736
rect 23063 12733 23075 12767
rect 23017 12727 23075 12733
rect 24946 12724 24952 12776
rect 25004 12773 25010 12776
rect 25004 12764 25016 12773
rect 26234 12764 26240 12776
rect 25004 12736 25049 12764
rect 25148 12736 26240 12764
rect 25004 12727 25016 12736
rect 25004 12724 25010 12727
rect 22557 12699 22615 12705
rect 22557 12696 22569 12699
rect 22296 12668 22569 12696
rect 22189 12659 22247 12665
rect 22557 12665 22569 12668
rect 22603 12665 22615 12699
rect 22557 12659 22615 12665
rect 22738 12656 22744 12708
rect 22796 12696 22802 12708
rect 25148 12696 25176 12736
rect 26234 12724 26240 12736
rect 26292 12724 26298 12776
rect 22796 12668 25176 12696
rect 22796 12656 22802 12668
rect 25222 12656 25228 12708
rect 25280 12696 25286 12708
rect 25930 12699 25988 12705
rect 25930 12696 25942 12699
rect 25280 12668 25942 12696
rect 25280 12656 25286 12668
rect 25930 12665 25942 12668
rect 25976 12665 25988 12699
rect 25930 12659 25988 12665
rect 15436 12600 15608 12628
rect 15436 12588 15442 12600
rect 15838 12588 15844 12640
rect 15896 12628 15902 12640
rect 17405 12631 17463 12637
rect 17405 12628 17417 12631
rect 15896 12600 17417 12628
rect 15896 12588 15902 12600
rect 17405 12597 17417 12600
rect 17451 12597 17463 12631
rect 17405 12591 17463 12597
rect 20070 12588 20076 12640
rect 20128 12588 20134 12640
rect 22646 12588 22652 12640
rect 22704 12588 22710 12640
rect 23290 12588 23296 12640
rect 23348 12628 23354 12640
rect 26050 12628 26056 12640
rect 23348 12600 26056 12628
rect 23348 12588 23354 12600
rect 26050 12588 26056 12600
rect 26108 12588 26114 12640
rect 552 12538 27576 12560
rect 552 12486 7114 12538
rect 7166 12486 7178 12538
rect 7230 12486 7242 12538
rect 7294 12486 7306 12538
rect 7358 12486 7370 12538
rect 7422 12486 13830 12538
rect 13882 12486 13894 12538
rect 13946 12486 13958 12538
rect 14010 12486 14022 12538
rect 14074 12486 14086 12538
rect 14138 12486 20546 12538
rect 20598 12486 20610 12538
rect 20662 12486 20674 12538
rect 20726 12486 20738 12538
rect 20790 12486 20802 12538
rect 20854 12486 27262 12538
rect 27314 12486 27326 12538
rect 27378 12486 27390 12538
rect 27442 12486 27454 12538
rect 27506 12486 27518 12538
rect 27570 12486 27576 12538
rect 552 12464 27576 12486
rect 2130 12384 2136 12436
rect 2188 12424 2194 12436
rect 2188 12396 2728 12424
rect 2188 12384 2194 12396
rect 1394 12356 1400 12368
rect 860 12328 1400 12356
rect 860 12297 888 12328
rect 1394 12316 1400 12328
rect 1452 12356 1458 12368
rect 2590 12365 2596 12368
rect 2584 12356 2596 12365
rect 1452 12328 2360 12356
rect 2551 12328 2596 12356
rect 1452 12316 1458 12328
rect 1118 12297 1124 12300
rect 845 12291 903 12297
rect 845 12257 857 12291
rect 891 12257 903 12291
rect 845 12251 903 12257
rect 1112 12251 1124 12297
rect 1118 12248 1124 12251
rect 1176 12248 1182 12300
rect 2332 12297 2360 12328
rect 2584 12319 2596 12328
rect 2590 12316 2596 12319
rect 2648 12316 2654 12368
rect 2700 12356 2728 12396
rect 3694 12384 3700 12436
rect 3752 12384 3758 12436
rect 4338 12384 4344 12436
rect 4396 12424 4402 12436
rect 5166 12424 5172 12436
rect 4396 12396 5172 12424
rect 4396 12384 4402 12396
rect 5166 12384 5172 12396
rect 5224 12384 5230 12436
rect 10965 12427 11023 12433
rect 10965 12424 10977 12427
rect 9508 12396 10977 12424
rect 7742 12356 7748 12368
rect 2700 12328 7748 12356
rect 7742 12316 7748 12328
rect 7800 12316 7806 12368
rect 9248 12359 9306 12365
rect 9248 12325 9260 12359
rect 9294 12356 9306 12359
rect 9508 12356 9536 12396
rect 10965 12393 10977 12396
rect 11011 12393 11023 12427
rect 10965 12387 11023 12393
rect 11514 12384 11520 12436
rect 11572 12384 11578 12436
rect 11885 12427 11943 12433
rect 11885 12393 11897 12427
rect 11931 12424 11943 12427
rect 12250 12424 12256 12436
rect 11931 12396 12256 12424
rect 11931 12393 11943 12396
rect 11885 12387 11943 12393
rect 12250 12384 12256 12396
rect 12308 12384 12314 12436
rect 13446 12384 13452 12436
rect 13504 12384 13510 12436
rect 13817 12427 13875 12433
rect 13817 12393 13829 12427
rect 13863 12424 13875 12427
rect 14182 12424 14188 12436
rect 13863 12396 14188 12424
rect 13863 12393 13875 12396
rect 13817 12387 13875 12393
rect 14182 12384 14188 12396
rect 14240 12384 14246 12436
rect 14274 12384 14280 12436
rect 14332 12384 14338 12436
rect 15654 12384 15660 12436
rect 15712 12384 15718 12436
rect 19242 12384 19248 12436
rect 19300 12384 19306 12436
rect 21453 12427 21511 12433
rect 21453 12393 21465 12427
rect 21499 12424 21511 12427
rect 22465 12427 22523 12433
rect 21499 12396 21956 12424
rect 21499 12393 21511 12396
rect 21453 12387 21511 12393
rect 9294 12328 9536 12356
rect 9294 12325 9306 12328
rect 9248 12319 9306 12325
rect 9582 12316 9588 12368
rect 9640 12316 9646 12368
rect 9766 12316 9772 12368
rect 9824 12365 9830 12368
rect 9824 12359 9843 12365
rect 9831 12325 9843 12359
rect 9824 12319 9843 12325
rect 9824 12316 9830 12319
rect 9950 12316 9956 12368
rect 10008 12356 10014 12368
rect 14292 12356 14320 12384
rect 10008 12328 11192 12356
rect 10008 12316 10014 12328
rect 2317 12291 2375 12297
rect 2317 12257 2329 12291
rect 2363 12257 2375 12291
rect 2317 12251 2375 12257
rect 3418 12248 3424 12300
rect 3476 12288 3482 12300
rect 3602 12288 3608 12300
rect 3476 12260 3608 12288
rect 3476 12248 3482 12260
rect 3602 12248 3608 12260
rect 3660 12248 3666 12300
rect 4246 12248 4252 12300
rect 4304 12248 4310 12300
rect 4525 12291 4583 12297
rect 4525 12257 4537 12291
rect 4571 12288 4583 12291
rect 4614 12288 4620 12300
rect 4571 12260 4620 12288
rect 4571 12257 4583 12260
rect 4525 12251 4583 12257
rect 4614 12248 4620 12260
rect 4672 12248 4678 12300
rect 4709 12291 4767 12297
rect 4709 12257 4721 12291
rect 4755 12288 4767 12291
rect 4893 12291 4951 12297
rect 4893 12288 4905 12291
rect 4755 12260 4905 12288
rect 4755 12257 4767 12260
rect 4709 12251 4767 12257
rect 4893 12257 4905 12260
rect 4939 12257 4951 12291
rect 4893 12251 4951 12257
rect 5350 12248 5356 12300
rect 5408 12288 5414 12300
rect 5813 12291 5871 12297
rect 5813 12288 5825 12291
rect 5408 12260 5825 12288
rect 5408 12248 5414 12260
rect 5813 12257 5825 12260
rect 5859 12257 5871 12291
rect 5813 12251 5871 12257
rect 5902 12248 5908 12300
rect 5960 12288 5966 12300
rect 11164 12297 11192 12328
rect 14016 12328 14320 12356
rect 6069 12291 6127 12297
rect 6069 12288 6081 12291
rect 5960 12260 6081 12288
rect 5960 12248 5966 12260
rect 6069 12257 6081 12260
rect 6115 12257 6127 12291
rect 6069 12251 6127 12257
rect 9493 12291 9551 12297
rect 9493 12257 9505 12291
rect 9539 12288 9551 12291
rect 11149 12291 11207 12297
rect 9539 12260 11100 12288
rect 9539 12257 9551 12260
rect 9493 12251 9551 12257
rect 4798 12180 4804 12232
rect 4856 12220 4862 12232
rect 5445 12223 5503 12229
rect 5445 12220 5457 12223
rect 4856 12192 5457 12220
rect 4856 12180 4862 12192
rect 5445 12189 5457 12192
rect 5491 12189 5503 12223
rect 5445 12183 5503 12189
rect 7837 12223 7895 12229
rect 7837 12189 7849 12223
rect 7883 12189 7895 12223
rect 7837 12183 7895 12189
rect 7006 12112 7012 12164
rect 7064 12152 7070 12164
rect 7285 12155 7343 12161
rect 7285 12152 7297 12155
rect 7064 12124 7297 12152
rect 7064 12112 7070 12124
rect 7285 12121 7297 12124
rect 7331 12121 7343 12155
rect 7285 12115 7343 12121
rect 2222 12044 2228 12096
rect 2280 12044 2286 12096
rect 4065 12087 4123 12093
rect 4065 12053 4077 12087
rect 4111 12084 4123 12087
rect 4154 12084 4160 12096
rect 4111 12056 4160 12084
rect 4111 12053 4123 12056
rect 4065 12047 4123 12053
rect 4154 12044 4160 12056
rect 4212 12044 4218 12096
rect 7193 12087 7251 12093
rect 7193 12053 7205 12087
rect 7239 12084 7251 12087
rect 7558 12084 7564 12096
rect 7239 12056 7564 12084
rect 7239 12053 7251 12056
rect 7193 12047 7251 12053
rect 7558 12044 7564 12056
rect 7616 12084 7622 12096
rect 7852 12084 7880 12183
rect 9582 12180 9588 12232
rect 9640 12220 9646 12232
rect 10597 12223 10655 12229
rect 10597 12220 10609 12223
rect 9640 12192 10609 12220
rect 9640 12180 9646 12192
rect 10597 12189 10609 12192
rect 10643 12189 10655 12223
rect 11072 12220 11100 12260
rect 11149 12257 11161 12291
rect 11195 12257 11207 12291
rect 11149 12251 11207 12257
rect 11330 12248 11336 12300
rect 11388 12248 11394 12300
rect 11422 12248 11428 12300
rect 11480 12248 11486 12300
rect 11698 12248 11704 12300
rect 11756 12248 11762 12300
rect 11977 12291 12035 12297
rect 11977 12257 11989 12291
rect 12023 12288 12035 12291
rect 12158 12288 12164 12300
rect 12023 12260 12164 12288
rect 12023 12257 12035 12260
rect 11977 12251 12035 12257
rect 12158 12248 12164 12260
rect 12216 12248 12222 12300
rect 12336 12291 12394 12297
rect 12336 12257 12348 12291
rect 12382 12288 12394 12291
rect 12710 12288 12716 12300
rect 12382 12260 12716 12288
rect 12382 12257 12394 12260
rect 12336 12251 12394 12257
rect 12710 12248 12716 12260
rect 12768 12248 12774 12300
rect 14016 12297 14044 12328
rect 14826 12316 14832 12368
rect 14884 12316 14890 12368
rect 18877 12359 18935 12365
rect 18877 12356 18889 12359
rect 15488 12328 18889 12356
rect 14001 12291 14059 12297
rect 14001 12257 14013 12291
rect 14047 12257 14059 12291
rect 14001 12251 14059 12257
rect 14185 12291 14243 12297
rect 14185 12257 14197 12291
rect 14231 12257 14243 12291
rect 14185 12251 14243 12257
rect 11882 12220 11888 12232
rect 11072 12192 11888 12220
rect 10597 12183 10655 12189
rect 11882 12180 11888 12192
rect 11940 12220 11946 12232
rect 12069 12223 12127 12229
rect 11940 12212 12020 12220
rect 12069 12212 12081 12223
rect 11940 12192 12081 12212
rect 11940 12180 11946 12192
rect 11992 12189 12081 12192
rect 12115 12189 12127 12223
rect 14200 12220 14228 12251
rect 14274 12248 14280 12300
rect 14332 12288 14338 12300
rect 14458 12288 14464 12300
rect 14332 12260 14464 12288
rect 14332 12248 14338 12260
rect 14458 12248 14464 12260
rect 14516 12248 14522 12300
rect 15488 12220 15516 12328
rect 18877 12325 18889 12328
rect 18923 12356 18935 12359
rect 19702 12356 19708 12368
rect 18923 12328 19708 12356
rect 18923 12325 18935 12328
rect 18877 12319 18935 12325
rect 19702 12316 19708 12328
rect 19760 12316 19766 12368
rect 15933 12291 15991 12297
rect 15933 12257 15945 12291
rect 15979 12288 15991 12291
rect 16206 12288 16212 12300
rect 15979 12260 16212 12288
rect 15979 12257 15991 12260
rect 15933 12251 15991 12257
rect 16206 12248 16212 12260
rect 16264 12248 16270 12300
rect 18506 12248 18512 12300
rect 18564 12288 18570 12300
rect 18785 12291 18843 12297
rect 18785 12288 18797 12291
rect 18564 12260 18797 12288
rect 18564 12248 18570 12260
rect 18785 12257 18797 12260
rect 18831 12257 18843 12291
rect 18785 12251 18843 12257
rect 18966 12248 18972 12300
rect 19024 12288 19030 12300
rect 19061 12291 19119 12297
rect 19061 12288 19073 12291
rect 19024 12260 19073 12288
rect 19024 12248 19030 12260
rect 19061 12257 19073 12260
rect 19107 12257 19119 12291
rect 19061 12251 19119 12257
rect 21634 12248 21640 12300
rect 21692 12286 21698 12300
rect 21928 12297 21956 12396
rect 22465 12393 22477 12427
rect 22511 12424 22523 12427
rect 22646 12424 22652 12436
rect 22511 12396 22652 12424
rect 22511 12393 22523 12396
rect 22465 12387 22523 12393
rect 22646 12384 22652 12396
rect 22704 12384 22710 12436
rect 23124 12396 23336 12424
rect 23124 12356 23152 12396
rect 22020 12328 23152 12356
rect 21821 12291 21879 12297
rect 21821 12286 21833 12291
rect 21692 12258 21833 12286
rect 21692 12248 21698 12258
rect 21821 12257 21833 12258
rect 21867 12257 21879 12291
rect 21821 12251 21879 12257
rect 21913 12291 21971 12297
rect 21913 12257 21925 12291
rect 21959 12257 21971 12291
rect 21913 12251 21971 12257
rect 11992 12184 12127 12189
rect 12069 12183 12127 12184
rect 13372 12192 15516 12220
rect 10045 12155 10103 12161
rect 10045 12152 10057 12155
rect 9784 12124 10057 12152
rect 7616 12056 7880 12084
rect 8113 12087 8171 12093
rect 7616 12044 7622 12056
rect 8113 12053 8125 12087
rect 8159 12084 8171 12087
rect 9122 12084 9128 12096
rect 8159 12056 9128 12084
rect 8159 12053 8171 12056
rect 8113 12047 8171 12053
rect 9122 12044 9128 12056
rect 9180 12044 9186 12096
rect 9784 12093 9812 12124
rect 10045 12121 10057 12124
rect 10091 12121 10103 12155
rect 10045 12115 10103 12121
rect 9769 12087 9827 12093
rect 9769 12053 9781 12087
rect 9815 12053 9827 12087
rect 9769 12047 9827 12053
rect 9953 12087 10011 12093
rect 9953 12053 9965 12087
rect 9999 12084 10011 12087
rect 10226 12084 10232 12096
rect 9999 12056 10232 12084
rect 9999 12053 10011 12056
rect 9953 12047 10011 12053
rect 10226 12044 10232 12056
rect 10284 12044 10290 12096
rect 10318 12044 10324 12096
rect 10376 12084 10382 12096
rect 12250 12084 12256 12096
rect 10376 12056 12256 12084
rect 10376 12044 10382 12056
rect 12250 12044 12256 12056
rect 12308 12084 12314 12096
rect 13372 12084 13400 12192
rect 15562 12180 15568 12232
rect 15620 12220 15626 12232
rect 15657 12223 15715 12229
rect 15657 12220 15669 12223
rect 15620 12192 15669 12220
rect 15620 12180 15626 12192
rect 15657 12189 15669 12192
rect 15703 12189 15715 12223
rect 15657 12183 15715 12189
rect 15841 12223 15899 12229
rect 15841 12189 15853 12223
rect 15887 12220 15899 12223
rect 16022 12220 16028 12232
rect 15887 12192 16028 12220
rect 15887 12189 15899 12192
rect 15841 12183 15899 12189
rect 16022 12180 16028 12192
rect 16080 12180 16086 12232
rect 17862 12180 17868 12232
rect 17920 12220 17926 12232
rect 18049 12223 18107 12229
rect 18049 12220 18061 12223
rect 17920 12192 18061 12220
rect 17920 12180 17926 12192
rect 18049 12189 18061 12192
rect 18095 12189 18107 12223
rect 18049 12183 18107 12189
rect 19702 12180 19708 12232
rect 19760 12220 19766 12232
rect 20070 12220 20076 12232
rect 19760 12192 20076 12220
rect 19760 12180 19766 12192
rect 20070 12180 20076 12192
rect 20128 12220 20134 12232
rect 20257 12223 20315 12229
rect 20257 12220 20269 12223
rect 20128 12192 20269 12220
rect 20128 12180 20134 12192
rect 20257 12189 20269 12192
rect 20303 12189 20315 12223
rect 20257 12183 20315 12189
rect 21729 12223 21787 12229
rect 21729 12189 21741 12223
rect 21775 12220 21787 12223
rect 22020 12220 22048 12328
rect 23198 12316 23204 12368
rect 23256 12316 23262 12368
rect 23308 12356 23336 12396
rect 23382 12384 23388 12436
rect 23440 12384 23446 12436
rect 23474 12384 23480 12436
rect 23532 12424 23538 12436
rect 23845 12427 23903 12433
rect 23845 12424 23857 12427
rect 23532 12396 23857 12424
rect 23532 12384 23538 12396
rect 23845 12393 23857 12396
rect 23891 12393 23903 12427
rect 25038 12424 25044 12436
rect 23845 12387 23903 12393
rect 23952 12396 25044 12424
rect 23952 12356 23980 12396
rect 25038 12384 25044 12396
rect 25096 12384 25102 12436
rect 25222 12384 25228 12436
rect 25280 12384 25286 12436
rect 26418 12384 26424 12436
rect 26476 12384 26482 12436
rect 23308 12328 23980 12356
rect 24029 12359 24087 12365
rect 24029 12325 24041 12359
rect 24075 12356 24087 12359
rect 24302 12356 24308 12368
rect 24075 12328 24308 12356
rect 24075 12325 24087 12328
rect 24029 12319 24087 12325
rect 24302 12316 24308 12328
rect 24360 12316 24366 12368
rect 25406 12316 25412 12368
rect 25464 12356 25470 12368
rect 26970 12356 26976 12368
rect 25464 12328 25820 12356
rect 25464 12316 25470 12328
rect 22462 12248 22468 12300
rect 22520 12288 22526 12300
rect 22741 12291 22799 12297
rect 22741 12288 22753 12291
rect 22520 12260 22753 12288
rect 22520 12248 22526 12260
rect 22741 12257 22753 12260
rect 22787 12257 22799 12291
rect 22741 12251 22799 12257
rect 22925 12291 22983 12297
rect 22925 12257 22937 12291
rect 22971 12288 22983 12291
rect 23017 12291 23075 12297
rect 23017 12288 23029 12291
rect 22971 12260 23029 12288
rect 22971 12257 22983 12260
rect 22925 12251 22983 12257
rect 23017 12257 23029 12260
rect 23063 12288 23075 12291
rect 23569 12291 23627 12297
rect 23569 12288 23581 12291
rect 23063 12260 23581 12288
rect 23063 12257 23075 12260
rect 23017 12251 23075 12257
rect 23569 12257 23581 12260
rect 23615 12288 23627 12291
rect 24213 12291 24271 12297
rect 24213 12288 24225 12291
rect 23615 12260 24225 12288
rect 23615 12257 23627 12260
rect 23569 12251 23627 12257
rect 24213 12257 24225 12260
rect 24259 12288 24271 12291
rect 24394 12288 24400 12300
rect 24259 12260 24400 12288
rect 24259 12257 24271 12260
rect 24213 12251 24271 12257
rect 24394 12248 24400 12260
rect 24452 12248 24458 12300
rect 25593 12291 25651 12297
rect 25593 12257 25605 12291
rect 25639 12257 25651 12291
rect 25593 12251 25651 12257
rect 21775 12192 22048 12220
rect 21775 12189 21787 12192
rect 21729 12183 21787 12189
rect 22094 12180 22100 12232
rect 22152 12220 22158 12232
rect 22189 12223 22247 12229
rect 22189 12220 22201 12223
rect 22152 12192 22201 12220
rect 22152 12180 22158 12192
rect 22189 12189 22201 12192
rect 22235 12189 22247 12223
rect 22189 12183 22247 12189
rect 24673 12223 24731 12229
rect 24673 12189 24685 12223
rect 24719 12220 24731 12223
rect 25317 12223 25375 12229
rect 25317 12220 25329 12223
rect 24719 12192 25329 12220
rect 24719 12189 24731 12192
rect 24673 12183 24731 12189
rect 25317 12189 25329 12192
rect 25363 12189 25375 12223
rect 25608 12220 25636 12251
rect 25682 12248 25688 12300
rect 25740 12248 25746 12300
rect 25792 12297 25820 12328
rect 26068 12328 26976 12356
rect 26068 12300 26096 12328
rect 26970 12316 26976 12328
rect 27028 12316 27034 12368
rect 25777 12291 25835 12297
rect 25777 12257 25789 12291
rect 25823 12257 25835 12291
rect 25777 12251 25835 12257
rect 25961 12291 26019 12297
rect 25961 12257 25973 12291
rect 26007 12288 26019 12291
rect 26050 12288 26056 12300
rect 26007 12260 26056 12288
rect 26007 12257 26019 12260
rect 25961 12251 26019 12257
rect 26050 12248 26056 12260
rect 26108 12248 26114 12300
rect 26694 12248 26700 12300
rect 26752 12248 26758 12300
rect 26789 12291 26847 12297
rect 26789 12257 26801 12291
rect 26835 12257 26847 12291
rect 26789 12251 26847 12257
rect 26142 12220 26148 12232
rect 25608 12192 26148 12220
rect 25317 12183 25375 12189
rect 26142 12180 26148 12192
rect 26200 12180 26206 12232
rect 13630 12112 13636 12164
rect 13688 12152 13694 12164
rect 14645 12155 14703 12161
rect 14645 12152 14657 12155
rect 13688 12124 14657 12152
rect 13688 12112 13694 12124
rect 14645 12121 14657 12124
rect 14691 12121 14703 12155
rect 24578 12152 24584 12164
rect 14645 12115 14703 12121
rect 21836 12124 24584 12152
rect 12308 12056 13400 12084
rect 12308 12044 12314 12056
rect 18138 12044 18144 12096
rect 18196 12084 18202 12096
rect 18693 12087 18751 12093
rect 18693 12084 18705 12087
rect 18196 12056 18705 12084
rect 18196 12044 18202 12056
rect 18693 12053 18705 12056
rect 18739 12053 18751 12087
rect 18693 12047 18751 12053
rect 19150 12044 19156 12096
rect 19208 12084 19214 12096
rect 21836 12093 21864 12124
rect 24578 12112 24584 12124
rect 24636 12112 24642 12164
rect 25682 12112 25688 12164
rect 25740 12152 25746 12164
rect 26804 12152 26832 12251
rect 26878 12248 26884 12300
rect 26936 12248 26942 12300
rect 26988 12288 27016 12316
rect 27065 12291 27123 12297
rect 27065 12288 27077 12291
rect 26988 12260 27077 12288
rect 27065 12257 27077 12260
rect 27111 12257 27123 12291
rect 27065 12251 27123 12257
rect 25740 12124 26832 12152
rect 25740 12112 25746 12124
rect 19705 12087 19763 12093
rect 19705 12084 19717 12087
rect 19208 12056 19717 12084
rect 19208 12044 19214 12056
rect 19705 12053 19717 12056
rect 19751 12053 19763 12087
rect 19705 12047 19763 12053
rect 21821 12087 21879 12093
rect 21821 12053 21833 12087
rect 21867 12053 21879 12087
rect 21821 12047 21879 12053
rect 22281 12087 22339 12093
rect 22281 12053 22293 12087
rect 22327 12084 22339 12087
rect 22554 12084 22560 12096
rect 22327 12056 22560 12084
rect 22327 12053 22339 12056
rect 22281 12047 22339 12053
rect 22554 12044 22560 12056
rect 22612 12044 22618 12096
rect 23198 12044 23204 12096
rect 23256 12084 23262 12096
rect 23661 12087 23719 12093
rect 23661 12084 23673 12087
rect 23256 12056 23673 12084
rect 23256 12044 23262 12056
rect 23661 12053 23673 12056
rect 23707 12053 23719 12087
rect 23661 12047 23719 12053
rect 552 11994 27416 12016
rect 552 11942 3756 11994
rect 3808 11942 3820 11994
rect 3872 11942 3884 11994
rect 3936 11942 3948 11994
rect 4000 11942 4012 11994
rect 4064 11942 10472 11994
rect 10524 11942 10536 11994
rect 10588 11942 10600 11994
rect 10652 11942 10664 11994
rect 10716 11942 10728 11994
rect 10780 11942 17188 11994
rect 17240 11942 17252 11994
rect 17304 11942 17316 11994
rect 17368 11942 17380 11994
rect 17432 11942 17444 11994
rect 17496 11942 23904 11994
rect 23956 11942 23968 11994
rect 24020 11942 24032 11994
rect 24084 11942 24096 11994
rect 24148 11942 24160 11994
rect 24212 11942 27416 11994
rect 552 11920 27416 11942
rect 1118 11840 1124 11892
rect 1176 11880 1182 11892
rect 1305 11883 1363 11889
rect 1305 11880 1317 11883
rect 1176 11852 1317 11880
rect 1176 11840 1182 11852
rect 1305 11849 1317 11852
rect 1351 11849 1363 11883
rect 1305 11843 1363 11849
rect 3421 11883 3479 11889
rect 3421 11849 3433 11883
rect 3467 11880 3479 11883
rect 3602 11880 3608 11892
rect 3467 11852 3608 11880
rect 3467 11849 3479 11852
rect 3421 11843 3479 11849
rect 3602 11840 3608 11852
rect 3660 11840 3666 11892
rect 4338 11880 4344 11892
rect 3712 11852 4344 11880
rect 3237 11815 3295 11821
rect 3237 11781 3249 11815
rect 3283 11812 3295 11815
rect 3712 11812 3740 11852
rect 4338 11840 4344 11852
rect 4396 11840 4402 11892
rect 4798 11840 4804 11892
rect 4856 11880 4862 11892
rect 5077 11883 5135 11889
rect 5077 11880 5089 11883
rect 4856 11852 5089 11880
rect 4856 11840 4862 11852
rect 5077 11849 5089 11852
rect 5123 11849 5135 11883
rect 5077 11843 5135 11849
rect 5629 11883 5687 11889
rect 5629 11849 5641 11883
rect 5675 11880 5687 11883
rect 5902 11880 5908 11892
rect 5675 11852 5908 11880
rect 5675 11849 5687 11852
rect 5629 11843 5687 11849
rect 5902 11840 5908 11852
rect 5960 11840 5966 11892
rect 6914 11840 6920 11892
rect 6972 11880 6978 11892
rect 7193 11883 7251 11889
rect 7193 11880 7205 11883
rect 6972 11852 7205 11880
rect 6972 11840 6978 11852
rect 7193 11849 7205 11852
rect 7239 11849 7251 11883
rect 7193 11843 7251 11849
rect 3283 11784 3740 11812
rect 3283 11781 3295 11784
rect 3237 11775 3295 11781
rect 2222 11704 2228 11756
rect 2280 11744 2286 11756
rect 2593 11747 2651 11753
rect 2593 11744 2605 11747
rect 2280 11716 2605 11744
rect 2280 11704 2286 11716
rect 2593 11713 2605 11716
rect 2639 11744 2651 11747
rect 2639 11716 2774 11744
rect 2639 11713 2651 11716
rect 2593 11707 2651 11713
rect 1394 11636 1400 11688
rect 1452 11676 1458 11688
rect 1857 11679 1915 11685
rect 1857 11676 1869 11679
rect 1452 11648 1869 11676
rect 1452 11636 1458 11648
rect 1857 11645 1869 11648
rect 1903 11645 1915 11679
rect 2746 11676 2774 11716
rect 6638 11704 6644 11756
rect 6696 11744 6702 11756
rect 7208 11744 7236 11843
rect 7466 11840 7472 11892
rect 7524 11840 7530 11892
rect 9582 11840 9588 11892
rect 9640 11840 9646 11892
rect 12161 11883 12219 11889
rect 12161 11849 12173 11883
rect 12207 11880 12219 11883
rect 12710 11880 12716 11892
rect 12207 11852 12716 11880
rect 12207 11849 12219 11852
rect 12161 11843 12219 11849
rect 12710 11840 12716 11852
rect 12768 11840 12774 11892
rect 12897 11883 12955 11889
rect 12897 11849 12909 11883
rect 12943 11880 12955 11883
rect 13262 11880 13268 11892
rect 12943 11852 13268 11880
rect 12943 11849 12955 11852
rect 12897 11843 12955 11849
rect 13262 11840 13268 11852
rect 13320 11880 13326 11892
rect 13446 11880 13452 11892
rect 13320 11852 13452 11880
rect 13320 11840 13326 11852
rect 13446 11840 13452 11852
rect 13504 11840 13510 11892
rect 14461 11883 14519 11889
rect 14461 11849 14473 11883
rect 14507 11880 14519 11883
rect 15654 11880 15660 11892
rect 14507 11852 15660 11880
rect 14507 11849 14519 11852
rect 14461 11843 14519 11849
rect 15654 11840 15660 11852
rect 15712 11880 15718 11892
rect 16117 11883 16175 11889
rect 16117 11880 16129 11883
rect 15712 11852 16129 11880
rect 15712 11840 15718 11852
rect 16117 11849 16129 11852
rect 16163 11880 16175 11883
rect 16206 11880 16212 11892
rect 16163 11852 16212 11880
rect 16163 11849 16175 11852
rect 16117 11843 16175 11849
rect 16206 11840 16212 11852
rect 16264 11840 16270 11892
rect 17862 11840 17868 11892
rect 17920 11840 17926 11892
rect 18138 11840 18144 11892
rect 18196 11840 18202 11892
rect 18966 11840 18972 11892
rect 19024 11840 19030 11892
rect 19150 11840 19156 11892
rect 19208 11840 19214 11892
rect 21818 11840 21824 11892
rect 21876 11840 21882 11892
rect 22281 11883 22339 11889
rect 22281 11849 22293 11883
rect 22327 11880 22339 11883
rect 24762 11880 24768 11892
rect 22327 11852 24768 11880
rect 22327 11849 22339 11852
rect 22281 11843 22339 11849
rect 24762 11840 24768 11852
rect 24820 11840 24826 11892
rect 25682 11880 25688 11892
rect 24872 11852 25688 11880
rect 20901 11815 20959 11821
rect 20901 11781 20913 11815
rect 20947 11812 20959 11815
rect 20990 11812 20996 11824
rect 20947 11784 20996 11812
rect 20947 11781 20959 11784
rect 20901 11775 20959 11781
rect 20990 11772 20996 11784
rect 21048 11812 21054 11824
rect 23106 11812 23112 11824
rect 21048 11784 23112 11812
rect 21048 11772 21054 11784
rect 23106 11772 23112 11784
rect 23164 11772 23170 11824
rect 10965 11747 11023 11753
rect 6696 11716 6960 11744
rect 7208 11716 8708 11744
rect 6696 11704 6702 11716
rect 3418 11676 3424 11688
rect 2746 11648 3424 11676
rect 1857 11639 1915 11645
rect 3418 11636 3424 11648
rect 3476 11636 3482 11688
rect 3697 11679 3755 11685
rect 3697 11645 3709 11679
rect 3743 11676 3755 11679
rect 5350 11676 5356 11688
rect 3743 11648 5356 11676
rect 3743 11645 3755 11648
rect 3697 11639 3755 11645
rect 5350 11636 5356 11648
rect 5408 11636 5414 11688
rect 5445 11679 5503 11685
rect 5445 11645 5457 11679
rect 5491 11645 5503 11679
rect 5445 11639 5503 11645
rect 5629 11679 5687 11685
rect 5629 11645 5641 11679
rect 5675 11676 5687 11679
rect 6273 11679 6331 11685
rect 6273 11676 6285 11679
rect 5675 11648 6285 11676
rect 5675 11645 5687 11648
rect 5629 11639 5687 11645
rect 6273 11645 6285 11648
rect 6319 11645 6331 11679
rect 6273 11639 6331 11645
rect 3436 11608 3464 11636
rect 3605 11611 3663 11617
rect 3605 11608 3617 11611
rect 3436 11580 3617 11608
rect 3605 11577 3617 11580
rect 3651 11577 3663 11611
rect 3605 11571 3663 11577
rect 3964 11611 4022 11617
rect 3964 11577 3976 11611
rect 4010 11608 4022 11611
rect 4062 11608 4068 11620
rect 4010 11580 4068 11608
rect 4010 11577 4022 11580
rect 3964 11571 4022 11577
rect 4062 11568 4068 11580
rect 4120 11568 4126 11620
rect 1854 11500 1860 11552
rect 1912 11540 1918 11552
rect 3418 11549 3424 11552
rect 2041 11543 2099 11549
rect 2041 11540 2053 11543
rect 1912 11512 2053 11540
rect 1912 11500 1918 11512
rect 2041 11509 2053 11512
rect 2087 11509 2099 11543
rect 2041 11503 2099 11509
rect 3405 11543 3424 11549
rect 3405 11509 3417 11543
rect 3405 11503 3424 11509
rect 3418 11500 3424 11503
rect 3476 11500 3482 11552
rect 5460 11540 5488 11639
rect 6730 11636 6736 11688
rect 6788 11676 6794 11688
rect 6825 11679 6883 11685
rect 6825 11676 6837 11679
rect 6788 11648 6837 11676
rect 6788 11636 6794 11648
rect 6825 11645 6837 11648
rect 6871 11645 6883 11679
rect 6932 11676 6960 11716
rect 7469 11679 7527 11685
rect 7469 11676 7481 11679
rect 6932 11648 7481 11676
rect 6825 11639 6883 11645
rect 7469 11645 7481 11648
rect 7515 11645 7527 11679
rect 7469 11639 7527 11645
rect 7558 11636 7564 11688
rect 7616 11636 7622 11688
rect 7760 11685 7788 11716
rect 7745 11679 7803 11685
rect 7745 11645 7757 11679
rect 7791 11645 7803 11679
rect 7745 11639 7803 11645
rect 8202 11636 8208 11688
rect 8260 11676 8266 11688
rect 8680 11685 8708 11716
rect 10965 11713 10977 11747
rect 11011 11744 11023 11747
rect 11882 11744 11888 11756
rect 11011 11716 11888 11744
rect 11011 11713 11023 11716
rect 10965 11707 11023 11713
rect 11882 11704 11888 11716
rect 11940 11704 11946 11756
rect 14737 11747 14795 11753
rect 14737 11713 14749 11747
rect 14783 11713 14795 11747
rect 14737 11707 14795 11713
rect 8481 11679 8539 11685
rect 8481 11676 8493 11679
rect 8260 11648 8493 11676
rect 8260 11636 8266 11648
rect 8481 11645 8493 11648
rect 8527 11645 8539 11679
rect 8481 11639 8539 11645
rect 8665 11679 8723 11685
rect 8665 11645 8677 11679
rect 8711 11645 8723 11679
rect 8665 11639 8723 11645
rect 12345 11679 12403 11685
rect 12345 11645 12357 11679
rect 12391 11645 12403 11679
rect 12345 11639 12403 11645
rect 6546 11568 6552 11620
rect 6604 11608 6610 11620
rect 7161 11611 7219 11617
rect 7161 11608 7173 11611
rect 6604 11580 7173 11608
rect 6604 11568 6610 11580
rect 7161 11577 7173 11580
rect 7207 11577 7219 11611
rect 7161 11571 7219 11577
rect 7377 11611 7435 11617
rect 7377 11577 7389 11611
rect 7423 11608 7435 11611
rect 7576 11608 7604 11636
rect 7423 11580 7604 11608
rect 7423 11577 7435 11580
rect 7377 11571 7435 11577
rect 10410 11568 10416 11620
rect 10468 11608 10474 11620
rect 10698 11611 10756 11617
rect 10698 11608 10710 11611
rect 10468 11580 10710 11608
rect 10468 11568 10474 11580
rect 10698 11577 10710 11580
rect 10744 11577 10756 11611
rect 12360 11608 12388 11639
rect 12526 11636 12532 11688
rect 12584 11676 12590 11688
rect 12621 11679 12679 11685
rect 12621 11676 12633 11679
rect 12584 11648 12633 11676
rect 12584 11636 12590 11648
rect 12621 11645 12633 11648
rect 12667 11645 12679 11679
rect 12621 11639 12679 11645
rect 14550 11636 14556 11688
rect 14608 11636 14614 11688
rect 14752 11676 14780 11707
rect 16390 11704 16396 11756
rect 16448 11744 16454 11756
rect 16485 11747 16543 11753
rect 16485 11744 16497 11747
rect 16448 11716 16497 11744
rect 16448 11704 16454 11716
rect 16485 11713 16497 11716
rect 16531 11713 16543 11747
rect 16485 11707 16543 11713
rect 20717 11747 20775 11753
rect 20717 11713 20729 11747
rect 20763 11744 20775 11747
rect 21082 11744 21088 11756
rect 20763 11716 21088 11744
rect 20763 11713 20775 11716
rect 20717 11707 20775 11713
rect 21082 11704 21088 11716
rect 21140 11704 21146 11756
rect 22094 11744 22100 11756
rect 21744 11716 22100 11744
rect 16408 11676 16436 11704
rect 21744 11688 21772 11716
rect 22094 11704 22100 11716
rect 22152 11704 22158 11756
rect 22480 11716 24624 11744
rect 14752 11648 16436 11676
rect 19058 11636 19064 11688
rect 19116 11636 19122 11688
rect 19702 11636 19708 11688
rect 19760 11636 19766 11688
rect 19978 11636 19984 11688
rect 20036 11636 20042 11688
rect 20993 11679 21051 11685
rect 20993 11676 21005 11679
rect 20640 11648 21005 11676
rect 12894 11617 12900 11620
rect 12881 11611 12900 11617
rect 12360 11580 12756 11608
rect 10698 11571 10756 11577
rect 6914 11540 6920 11552
rect 5460 11512 6920 11540
rect 6914 11500 6920 11512
rect 6972 11540 6978 11552
rect 7009 11543 7067 11549
rect 7009 11540 7021 11543
rect 6972 11512 7021 11540
rect 6972 11500 6978 11512
rect 7009 11509 7021 11512
rect 7055 11509 7067 11543
rect 7009 11503 7067 11509
rect 9398 11500 9404 11552
rect 9456 11540 9462 11552
rect 9493 11543 9551 11549
rect 9493 11540 9505 11543
rect 9456 11512 9505 11540
rect 9456 11500 9462 11512
rect 9493 11509 9505 11512
rect 9539 11509 9551 11543
rect 9493 11503 9551 11509
rect 11330 11500 11336 11552
rect 11388 11540 11394 11552
rect 12526 11540 12532 11552
rect 11388 11512 12532 11540
rect 11388 11500 11394 11512
rect 12526 11500 12532 11512
rect 12584 11500 12590 11552
rect 12728 11549 12756 11580
rect 12881 11577 12893 11611
rect 12881 11571 12900 11577
rect 12894 11568 12900 11571
rect 12952 11568 12958 11620
rect 12986 11568 12992 11620
rect 13044 11608 13050 11620
rect 13081 11611 13139 11617
rect 13081 11608 13093 11611
rect 13044 11580 13093 11608
rect 13044 11568 13050 11580
rect 13081 11577 13093 11580
rect 13127 11608 13139 11611
rect 13630 11608 13636 11620
rect 13127 11580 13636 11608
rect 13127 11577 13139 11580
rect 13081 11571 13139 11577
rect 13630 11568 13636 11580
rect 13688 11568 13694 11620
rect 14277 11611 14335 11617
rect 14277 11577 14289 11611
rect 14323 11608 14335 11611
rect 14568 11608 14596 11636
rect 14734 11608 14740 11620
rect 14323 11580 14740 11608
rect 14323 11577 14335 11580
rect 14277 11571 14335 11577
rect 14734 11568 14740 11580
rect 14792 11568 14798 11620
rect 15004 11611 15062 11617
rect 15004 11577 15016 11611
rect 15050 11608 15062 11611
rect 15378 11608 15384 11620
rect 15050 11580 15384 11608
rect 15050 11577 15062 11580
rect 15004 11571 15062 11577
rect 15378 11568 15384 11580
rect 15436 11568 15442 11620
rect 16752 11611 16810 11617
rect 16752 11577 16764 11611
rect 16798 11608 16810 11611
rect 16942 11608 16948 11620
rect 16798 11580 16948 11608
rect 16798 11577 16810 11580
rect 16752 11571 16810 11577
rect 16942 11568 16948 11580
rect 17000 11568 17006 11620
rect 18322 11568 18328 11620
rect 18380 11608 18386 11620
rect 19076 11608 19104 11636
rect 19337 11611 19395 11617
rect 19337 11608 19349 11611
rect 18380 11580 19349 11608
rect 18380 11568 18386 11580
rect 19337 11577 19349 11580
rect 19383 11577 19395 11611
rect 19337 11571 19395 11577
rect 12713 11543 12771 11549
rect 12713 11509 12725 11543
rect 12759 11509 12771 11543
rect 12713 11503 12771 11509
rect 14366 11500 14372 11552
rect 14424 11540 14430 11552
rect 14477 11543 14535 11549
rect 14477 11540 14489 11543
rect 14424 11512 14489 11540
rect 14424 11500 14430 11512
rect 14477 11509 14489 11512
rect 14523 11509 14535 11543
rect 14477 11503 14535 11509
rect 14645 11543 14703 11549
rect 14645 11509 14657 11543
rect 14691 11540 14703 11543
rect 15562 11540 15568 11552
rect 14691 11512 15568 11540
rect 14691 11509 14703 11512
rect 14645 11503 14703 11509
rect 15562 11500 15568 11512
rect 15620 11500 15626 11552
rect 17126 11500 17132 11552
rect 17184 11540 17190 11552
rect 17957 11543 18015 11549
rect 17957 11540 17969 11543
rect 17184 11512 17969 11540
rect 17184 11500 17190 11512
rect 17957 11509 17969 11512
rect 18003 11509 18015 11543
rect 17957 11503 18015 11509
rect 18125 11543 18183 11549
rect 18125 11509 18137 11543
rect 18171 11540 18183 11543
rect 18874 11540 18880 11552
rect 18171 11512 18880 11540
rect 18171 11509 18183 11512
rect 18125 11503 18183 11509
rect 18874 11500 18880 11512
rect 18932 11540 18938 11552
rect 19127 11543 19185 11549
rect 19127 11540 19139 11543
rect 18932 11512 19139 11540
rect 18932 11500 18938 11512
rect 19127 11509 19139 11512
rect 19173 11509 19185 11543
rect 19127 11503 19185 11509
rect 19610 11500 19616 11552
rect 19668 11500 19674 11552
rect 20346 11500 20352 11552
rect 20404 11540 20410 11552
rect 20640 11549 20668 11648
rect 20993 11645 21005 11648
rect 21039 11645 21051 11679
rect 20993 11639 21051 11645
rect 21726 11636 21732 11688
rect 21784 11636 21790 11688
rect 21821 11679 21879 11685
rect 21821 11645 21833 11679
rect 21867 11676 21879 11679
rect 21867 11673 22140 11676
rect 22278 11673 22284 11688
rect 21867 11648 22284 11673
rect 21867 11645 21879 11648
rect 22112 11645 22284 11648
rect 21821 11639 21879 11645
rect 22278 11636 22284 11645
rect 22336 11636 22342 11688
rect 22370 11636 22376 11688
rect 22428 11636 22434 11688
rect 21545 11611 21603 11617
rect 21545 11577 21557 11611
rect 21591 11608 21603 11611
rect 21913 11611 21971 11617
rect 21591 11580 21772 11608
rect 21591 11577 21603 11580
rect 21545 11571 21603 11577
rect 20625 11543 20683 11549
rect 20625 11540 20637 11543
rect 20404 11512 20637 11540
rect 20404 11500 20410 11512
rect 20625 11509 20637 11512
rect 20671 11509 20683 11543
rect 20625 11503 20683 11509
rect 20717 11543 20775 11549
rect 20717 11509 20729 11543
rect 20763 11540 20775 11543
rect 20898 11540 20904 11552
rect 20763 11512 20904 11540
rect 20763 11509 20775 11512
rect 20717 11503 20775 11509
rect 20898 11500 20904 11512
rect 20956 11500 20962 11552
rect 21744 11540 21772 11580
rect 21913 11577 21925 11611
rect 21959 11608 21971 11611
rect 22002 11608 22008 11620
rect 21959 11580 22008 11608
rect 21959 11577 21971 11580
rect 21913 11571 21971 11577
rect 22002 11568 22008 11580
rect 22060 11568 22066 11620
rect 22097 11611 22155 11617
rect 22097 11577 22109 11611
rect 22143 11608 22155 11611
rect 22480 11608 22508 11716
rect 22554 11636 22560 11688
rect 22612 11636 22618 11688
rect 22649 11679 22707 11685
rect 22649 11645 22661 11679
rect 22695 11645 22707 11679
rect 22649 11639 22707 11645
rect 22741 11679 22799 11685
rect 22741 11645 22753 11679
rect 22787 11676 22799 11679
rect 23845 11679 23903 11685
rect 23845 11676 23857 11679
rect 22787 11648 23857 11676
rect 22787 11645 22799 11648
rect 22741 11639 22799 11645
rect 23845 11645 23857 11648
rect 23891 11645 23903 11679
rect 23845 11639 23903 11645
rect 24397 11679 24455 11685
rect 24397 11645 24409 11679
rect 24443 11645 24455 11679
rect 24397 11639 24455 11645
rect 22143 11580 22508 11608
rect 22664 11608 22692 11639
rect 22664 11580 23152 11608
rect 22143 11577 22155 11580
rect 22097 11571 22155 11577
rect 22830 11540 22836 11552
rect 21744 11512 22836 11540
rect 22830 11500 22836 11512
rect 22888 11500 22894 11552
rect 23014 11500 23020 11552
rect 23072 11500 23078 11552
rect 23124 11540 23152 11580
rect 23198 11568 23204 11620
rect 23256 11568 23262 11620
rect 23385 11611 23443 11617
rect 23385 11577 23397 11611
rect 23431 11608 23443 11611
rect 23658 11608 23664 11620
rect 23431 11580 23664 11608
rect 23431 11577 23443 11580
rect 23385 11571 23443 11577
rect 23658 11568 23664 11580
rect 23716 11608 23722 11620
rect 24412 11608 24440 11639
rect 23716 11580 24440 11608
rect 24596 11608 24624 11716
rect 24872 11685 24900 11852
rect 25682 11840 25688 11852
rect 25740 11840 25746 11892
rect 26602 11840 26608 11892
rect 26660 11880 26666 11892
rect 26970 11880 26976 11892
rect 26660 11852 26976 11880
rect 26660 11840 26666 11852
rect 26970 11840 26976 11852
rect 27028 11880 27034 11892
rect 27065 11883 27123 11889
rect 27065 11880 27077 11883
rect 27028 11852 27077 11880
rect 27028 11840 27034 11852
rect 27065 11849 27077 11852
rect 27111 11849 27123 11883
rect 27065 11843 27123 11849
rect 25056 11716 25360 11744
rect 24857 11679 24915 11685
rect 24857 11645 24869 11679
rect 24903 11645 24915 11679
rect 24857 11639 24915 11645
rect 24946 11636 24952 11688
rect 25004 11636 25010 11688
rect 25056 11608 25084 11716
rect 25130 11636 25136 11688
rect 25188 11636 25194 11688
rect 25332 11685 25360 11716
rect 25590 11704 25596 11756
rect 25648 11744 25654 11756
rect 25685 11747 25743 11753
rect 25685 11744 25697 11747
rect 25648 11716 25697 11744
rect 25648 11704 25654 11716
rect 25685 11713 25697 11716
rect 25731 11713 25743 11747
rect 25685 11707 25743 11713
rect 25225 11679 25283 11685
rect 25225 11645 25237 11679
rect 25271 11645 25283 11679
rect 25225 11639 25283 11645
rect 25317 11679 25375 11685
rect 25317 11645 25329 11679
rect 25363 11676 25375 11679
rect 26418 11676 26424 11688
rect 25363 11648 26424 11676
rect 25363 11645 25375 11648
rect 25317 11639 25375 11645
rect 24596 11580 25084 11608
rect 23716 11568 23722 11580
rect 23474 11540 23480 11552
rect 23124 11512 23480 11540
rect 23474 11500 23480 11512
rect 23532 11500 23538 11552
rect 23569 11543 23627 11549
rect 23569 11509 23581 11543
rect 23615 11540 23627 11543
rect 24486 11540 24492 11552
rect 23615 11512 24492 11540
rect 23615 11509 23627 11512
rect 23569 11503 23627 11509
rect 24486 11500 24492 11512
rect 24544 11500 24550 11552
rect 24578 11500 24584 11552
rect 24636 11540 24642 11552
rect 24673 11543 24731 11549
rect 24673 11540 24685 11543
rect 24636 11512 24685 11540
rect 24636 11500 24642 11512
rect 24673 11509 24685 11512
rect 24719 11540 24731 11543
rect 25240 11540 25268 11639
rect 26418 11636 26424 11648
rect 26476 11636 26482 11688
rect 25593 11611 25651 11617
rect 25593 11577 25605 11611
rect 25639 11608 25651 11611
rect 25930 11611 25988 11617
rect 25930 11608 25942 11611
rect 25639 11580 25942 11608
rect 25639 11577 25651 11580
rect 25593 11571 25651 11577
rect 25930 11577 25942 11580
rect 25976 11577 25988 11611
rect 25930 11571 25988 11577
rect 24719 11512 25268 11540
rect 24719 11509 24731 11512
rect 24673 11503 24731 11509
rect 552 11450 27576 11472
rect 552 11398 7114 11450
rect 7166 11398 7178 11450
rect 7230 11398 7242 11450
rect 7294 11398 7306 11450
rect 7358 11398 7370 11450
rect 7422 11398 13830 11450
rect 13882 11398 13894 11450
rect 13946 11398 13958 11450
rect 14010 11398 14022 11450
rect 14074 11398 14086 11450
rect 14138 11398 20546 11450
rect 20598 11398 20610 11450
rect 20662 11398 20674 11450
rect 20726 11398 20738 11450
rect 20790 11398 20802 11450
rect 20854 11398 27262 11450
rect 27314 11398 27326 11450
rect 27378 11398 27390 11450
rect 27442 11398 27454 11450
rect 27506 11398 27518 11450
rect 27570 11398 27576 11450
rect 552 11376 27576 11398
rect 1394 11296 1400 11348
rect 1452 11296 1458 11348
rect 2593 11339 2651 11345
rect 2593 11305 2605 11339
rect 2639 11336 2651 11339
rect 3234 11336 3240 11348
rect 2639 11308 3240 11336
rect 2639 11305 2651 11308
rect 2593 11299 2651 11305
rect 3234 11296 3240 11308
rect 3292 11296 3298 11348
rect 6730 11296 6736 11348
rect 6788 11296 6794 11348
rect 6914 11296 6920 11348
rect 6972 11296 6978 11348
rect 9122 11296 9128 11348
rect 9180 11336 9186 11348
rect 9401 11339 9459 11345
rect 9180 11308 9352 11336
rect 9180 11296 9186 11308
rect 6549 11271 6607 11277
rect 6549 11237 6561 11271
rect 6595 11268 6607 11271
rect 6932 11268 6960 11296
rect 6595 11240 6960 11268
rect 6595 11237 6607 11240
rect 6549 11231 6607 11237
rect 8846 11228 8852 11280
rect 8904 11268 8910 11280
rect 9033 11271 9091 11277
rect 9033 11268 9045 11271
rect 8904 11240 9045 11268
rect 8904 11228 8910 11240
rect 9033 11237 9045 11240
rect 9079 11237 9091 11271
rect 9233 11271 9291 11277
rect 9233 11268 9245 11271
rect 9033 11231 9091 11237
rect 9140 11240 9245 11268
rect 1581 11203 1639 11209
rect 1581 11169 1593 11203
rect 1627 11200 1639 11203
rect 1670 11200 1676 11212
rect 1627 11172 1676 11200
rect 1627 11169 1639 11172
rect 1581 11163 1639 11169
rect 1670 11160 1676 11172
rect 1728 11160 1734 11212
rect 1854 11160 1860 11212
rect 1912 11160 1918 11212
rect 2961 11203 3019 11209
rect 2961 11169 2973 11203
rect 3007 11200 3019 11203
rect 4338 11200 4344 11212
rect 3007 11172 4344 11200
rect 3007 11169 3019 11172
rect 2961 11163 3019 11169
rect 4338 11160 4344 11172
rect 4396 11160 4402 11212
rect 6365 11203 6423 11209
rect 6365 11169 6377 11203
rect 6411 11200 6423 11203
rect 6638 11200 6644 11212
rect 6411 11172 6644 11200
rect 6411 11169 6423 11172
rect 6365 11163 6423 11169
rect 6638 11160 6644 11172
rect 6696 11160 6702 11212
rect 6822 11160 6828 11212
rect 6880 11200 6886 11212
rect 6917 11203 6975 11209
rect 6917 11200 6929 11203
rect 6880 11172 6929 11200
rect 6880 11160 6886 11172
rect 6917 11169 6929 11172
rect 6963 11169 6975 11203
rect 6917 11163 6975 11169
rect 7006 11160 7012 11212
rect 7064 11160 7070 11212
rect 7285 11203 7343 11209
rect 7285 11169 7297 11203
rect 7331 11200 7343 11203
rect 7558 11200 7564 11212
rect 7331 11172 7564 11200
rect 7331 11169 7343 11172
rect 7285 11163 7343 11169
rect 7558 11160 7564 11172
rect 7616 11160 7622 11212
rect 1765 11135 1823 11141
rect 1765 11101 1777 11135
rect 1811 11132 1823 11135
rect 2314 11132 2320 11144
rect 1811 11104 2320 11132
rect 1811 11101 1823 11104
rect 1765 11095 1823 11101
rect 2314 11092 2320 11104
rect 2372 11132 2378 11144
rect 3418 11132 3424 11144
rect 2372 11104 3424 11132
rect 2372 11092 2378 11104
rect 3418 11092 3424 11104
rect 3476 11092 3482 11144
rect 6086 11092 6092 11144
rect 6144 11132 6150 11144
rect 6733 11135 6791 11141
rect 6733 11132 6745 11135
rect 6144 11104 6745 11132
rect 6144 11092 6150 11104
rect 6733 11101 6745 11104
rect 6779 11101 6791 11135
rect 6733 11095 6791 11101
rect 7193 11135 7251 11141
rect 7193 11101 7205 11135
rect 7239 11132 7251 11135
rect 8202 11132 8208 11144
rect 7239 11104 8208 11132
rect 7239 11101 7251 11104
rect 7193 11095 7251 11101
rect 2409 11067 2467 11073
rect 2409 11033 2421 11067
rect 2455 11064 2467 11067
rect 2774 11064 2780 11076
rect 2455 11036 2780 11064
rect 2455 11033 2467 11036
rect 2409 11027 2467 11033
rect 2774 11024 2780 11036
rect 2832 11024 2838 11076
rect 7006 11024 7012 11076
rect 7064 11064 7070 11076
rect 7208 11064 7236 11095
rect 8202 11092 8208 11104
rect 8260 11092 8266 11144
rect 7064 11036 7236 11064
rect 7653 11067 7711 11073
rect 7064 11024 7070 11036
rect 7653 11033 7665 11067
rect 7699 11064 7711 11067
rect 8938 11064 8944 11076
rect 7699 11036 8944 11064
rect 7699 11033 7711 11036
rect 7653 11027 7711 11033
rect 8938 11024 8944 11036
rect 8996 11024 9002 11076
rect 9140 11064 9168 11240
rect 9233 11237 9245 11240
rect 9279 11237 9291 11271
rect 9233 11231 9291 11237
rect 9324 11200 9352 11308
rect 9401 11305 9413 11339
rect 9447 11336 9459 11339
rect 9950 11336 9956 11348
rect 9447 11308 9956 11336
rect 9447 11305 9459 11308
rect 9401 11299 9459 11305
rect 9950 11296 9956 11308
rect 10008 11296 10014 11348
rect 10410 11296 10416 11348
rect 10468 11296 10474 11348
rect 11882 11336 11888 11348
rect 10980 11308 11888 11336
rect 9582 11228 9588 11280
rect 9640 11228 9646 11280
rect 10045 11271 10103 11277
rect 10045 11237 10057 11271
rect 10091 11268 10103 11271
rect 10980 11268 11008 11308
rect 11882 11296 11888 11308
rect 11940 11296 11946 11348
rect 12526 11296 12532 11348
rect 12584 11336 12590 11348
rect 14553 11339 14611 11345
rect 12584 11308 13768 11336
rect 12584 11296 12590 11308
rect 13630 11268 13636 11280
rect 10091 11240 11008 11268
rect 11072 11240 13636 11268
rect 10091 11237 10103 11240
rect 10045 11231 10103 11237
rect 9493 11203 9551 11209
rect 9493 11200 9505 11203
rect 9324 11172 9505 11200
rect 9493 11169 9505 11172
rect 9539 11169 9551 11203
rect 9600 11200 9628 11228
rect 9677 11203 9735 11209
rect 9677 11200 9689 11203
rect 9600 11172 9689 11200
rect 9493 11163 9551 11169
rect 9677 11169 9689 11172
rect 9723 11169 9735 11203
rect 9677 11163 9735 11169
rect 9858 11160 9864 11212
rect 9916 11200 9922 11212
rect 9953 11203 10011 11209
rect 9953 11200 9965 11203
rect 9916 11172 9965 11200
rect 9916 11160 9922 11172
rect 9953 11169 9965 11172
rect 9999 11169 10011 11203
rect 9953 11163 10011 11169
rect 10226 11160 10232 11212
rect 10284 11160 10290 11212
rect 11072 11209 11100 11240
rect 11057 11203 11115 11209
rect 11057 11169 11069 11203
rect 11103 11169 11115 11203
rect 11057 11163 11115 11169
rect 11324 11203 11382 11209
rect 11324 11169 11336 11203
rect 11370 11200 11382 11203
rect 11606 11200 11612 11212
rect 11370 11172 11612 11200
rect 11370 11169 11382 11172
rect 11324 11163 11382 11169
rect 11606 11160 11612 11172
rect 11664 11160 11670 11212
rect 13188 11209 13216 11240
rect 13630 11228 13636 11240
rect 13688 11228 13694 11280
rect 13446 11209 13452 11212
rect 13173 11203 13231 11209
rect 13173 11169 13185 11203
rect 13219 11169 13231 11203
rect 13173 11163 13231 11169
rect 13440 11163 13452 11209
rect 13446 11160 13452 11163
rect 13504 11160 13510 11212
rect 13740 11200 13768 11308
rect 14553 11305 14565 11339
rect 14599 11336 14611 11339
rect 15286 11336 15292 11348
rect 14599 11308 15292 11336
rect 14599 11305 14611 11308
rect 14553 11299 14611 11305
rect 15286 11296 15292 11308
rect 15344 11296 15350 11348
rect 15378 11296 15384 11348
rect 15436 11296 15442 11348
rect 15749 11339 15807 11345
rect 15749 11305 15761 11339
rect 15795 11336 15807 11339
rect 15795 11308 16620 11336
rect 15795 11305 15807 11308
rect 15749 11299 15807 11305
rect 14274 11228 14280 11280
rect 14332 11268 14338 11280
rect 14332 11240 15884 11268
rect 14332 11228 14338 11240
rect 13740 11172 15424 11200
rect 9214 11092 9220 11144
rect 9272 11132 9278 11144
rect 9585 11135 9643 11141
rect 9585 11132 9597 11135
rect 9272 11104 9597 11132
rect 9272 11092 9278 11104
rect 9585 11101 9597 11104
rect 9631 11101 9643 11135
rect 9585 11095 9643 11101
rect 15286 11092 15292 11144
rect 15344 11092 15350 11144
rect 15396 11132 15424 11172
rect 15562 11160 15568 11212
rect 15620 11160 15626 11212
rect 15856 11209 15884 11240
rect 15841 11203 15899 11209
rect 15841 11169 15853 11203
rect 15887 11169 15899 11203
rect 15841 11163 15899 11169
rect 15948 11132 15976 11308
rect 16592 11280 16620 11308
rect 16942 11296 16948 11348
rect 17000 11296 17006 11348
rect 19705 11339 19763 11345
rect 19705 11336 19717 11339
rect 19168 11308 19717 11336
rect 16574 11228 16580 11280
rect 16632 11268 16638 11280
rect 17313 11271 17371 11277
rect 17313 11268 17325 11271
rect 16632 11240 17325 11268
rect 16632 11228 16638 11240
rect 17313 11237 17325 11240
rect 17359 11237 17371 11271
rect 17313 11231 17371 11237
rect 16114 11160 16120 11212
rect 16172 11160 16178 11212
rect 16206 11160 16212 11212
rect 16264 11200 16270 11212
rect 16301 11203 16359 11209
rect 16301 11200 16313 11203
rect 16264 11172 16313 11200
rect 16264 11160 16270 11172
rect 16301 11169 16313 11172
rect 16347 11169 16359 11203
rect 16301 11163 16359 11169
rect 17126 11160 17132 11212
rect 17184 11160 17190 11212
rect 17405 11203 17463 11209
rect 17405 11169 17417 11203
rect 17451 11169 17463 11203
rect 17405 11163 17463 11169
rect 17681 11203 17739 11209
rect 17681 11169 17693 11203
rect 17727 11200 17739 11203
rect 17862 11200 17868 11212
rect 17727 11172 17868 11200
rect 17727 11169 17739 11172
rect 17681 11163 17739 11169
rect 15396 11104 15976 11132
rect 17420 11132 17448 11163
rect 17862 11160 17868 11172
rect 17920 11160 17926 11212
rect 19168 11209 19196 11308
rect 19705 11305 19717 11308
rect 19751 11336 19763 11339
rect 19978 11336 19984 11348
rect 19751 11308 19984 11336
rect 19751 11305 19763 11308
rect 19705 11299 19763 11305
rect 19978 11296 19984 11308
rect 20036 11296 20042 11348
rect 20438 11296 20444 11348
rect 20496 11336 20502 11348
rect 21726 11336 21732 11348
rect 20496 11308 21732 11336
rect 20496 11296 20502 11308
rect 21726 11296 21732 11308
rect 21784 11296 21790 11348
rect 22002 11296 22008 11348
rect 22060 11296 22066 11348
rect 22462 11296 22468 11348
rect 22520 11296 22526 11348
rect 23198 11336 23204 11348
rect 22756 11308 23204 11336
rect 19610 11228 19616 11280
rect 19668 11228 19674 11280
rect 20806 11268 20812 11280
rect 20864 11277 20870 11280
rect 20776 11240 20812 11268
rect 20806 11228 20812 11240
rect 20864 11231 20876 11277
rect 20864 11228 20870 11231
rect 21542 11228 21548 11280
rect 21600 11268 21606 11280
rect 22020 11268 22048 11296
rect 22756 11268 22784 11308
rect 23198 11296 23204 11308
rect 23256 11336 23262 11348
rect 23474 11336 23480 11348
rect 23256 11308 23480 11336
rect 23256 11296 23262 11308
rect 23474 11296 23480 11308
rect 23532 11296 23538 11348
rect 23566 11296 23572 11348
rect 23624 11336 23630 11348
rect 24578 11336 24584 11348
rect 23624 11308 24584 11336
rect 23624 11296 23630 11308
rect 24578 11296 24584 11308
rect 24636 11296 24642 11348
rect 26142 11296 26148 11348
rect 26200 11336 26206 11348
rect 26421 11339 26479 11345
rect 26421 11336 26433 11339
rect 26200 11308 26433 11336
rect 26200 11296 26206 11308
rect 26421 11305 26433 11308
rect 26467 11305 26479 11339
rect 26421 11299 26479 11305
rect 21600 11240 22784 11268
rect 22824 11271 22882 11277
rect 21600 11228 21606 11240
rect 22824 11237 22836 11271
rect 22870 11268 22882 11271
rect 23014 11268 23020 11280
rect 22870 11240 23020 11268
rect 22870 11237 22882 11240
rect 22824 11231 22882 11237
rect 23014 11228 23020 11240
rect 23072 11228 23078 11280
rect 25164 11271 25222 11277
rect 25164 11237 25176 11271
rect 25210 11268 25222 11271
rect 25501 11271 25559 11277
rect 25501 11268 25513 11271
rect 25210 11240 25513 11268
rect 25210 11237 25222 11240
rect 25164 11231 25222 11237
rect 25501 11237 25513 11240
rect 25547 11237 25559 11271
rect 25501 11231 25559 11237
rect 19133 11203 19196 11209
rect 19133 11169 19145 11203
rect 19179 11172 19196 11203
rect 19245 11203 19303 11209
rect 19179 11169 19191 11172
rect 19133 11163 19191 11169
rect 19245 11169 19257 11203
rect 19291 11200 19303 11203
rect 20070 11200 20076 11212
rect 19291 11172 20076 11200
rect 19291 11169 19303 11172
rect 19245 11163 19303 11169
rect 20070 11160 20076 11172
rect 20128 11160 20134 11212
rect 21085 11203 21143 11209
rect 21085 11169 21097 11203
rect 21131 11200 21143 11203
rect 22002 11200 22008 11212
rect 21131 11172 22008 11200
rect 21131 11169 21143 11172
rect 21085 11163 21143 11169
rect 22002 11160 22008 11172
rect 22060 11200 22066 11212
rect 22557 11203 22615 11209
rect 22557 11200 22569 11203
rect 22060 11172 22569 11200
rect 22060 11160 22066 11172
rect 22557 11169 22569 11172
rect 22603 11169 22615 11203
rect 22557 11163 22615 11169
rect 27062 11160 27068 11212
rect 27120 11160 27126 11212
rect 18414 11132 18420 11144
rect 17420 11104 18420 11132
rect 18414 11092 18420 11104
rect 18472 11092 18478 11144
rect 19521 11135 19579 11141
rect 19521 11132 19533 11135
rect 19444 11104 19533 11132
rect 9766 11064 9772 11076
rect 9140 11036 9772 11064
rect 9766 11024 9772 11036
rect 9824 11064 9830 11076
rect 10318 11064 10324 11076
rect 9824 11036 10324 11064
rect 9824 11024 9830 11036
rect 10318 11024 10324 11036
rect 10376 11064 10382 11076
rect 10962 11064 10968 11076
rect 10376 11036 10968 11064
rect 10376 11024 10382 11036
rect 10962 11024 10968 11036
rect 11020 11024 11026 11076
rect 18969 11067 19027 11073
rect 18969 11064 18981 11067
rect 12360 11036 13032 11064
rect 2498 10956 2504 11008
rect 2556 10996 2562 11008
rect 2593 10999 2651 11005
rect 2593 10996 2605 10999
rect 2556 10968 2605 10996
rect 2556 10956 2562 10968
rect 2593 10965 2605 10968
rect 2639 10996 2651 10999
rect 2682 10996 2688 11008
rect 2639 10968 2688 10996
rect 2639 10965 2651 10968
rect 2593 10959 2651 10965
rect 2682 10956 2688 10968
rect 2740 10956 2746 11008
rect 6178 10956 6184 11008
rect 6236 10956 6242 11008
rect 9122 10956 9128 11008
rect 9180 10996 9186 11008
rect 9217 10999 9275 11005
rect 9217 10996 9229 10999
rect 9180 10968 9229 10996
rect 9180 10956 9186 10968
rect 9217 10965 9229 10968
rect 9263 10965 9275 10999
rect 9217 10959 9275 10965
rect 9306 10956 9312 11008
rect 9364 10996 9370 11008
rect 12360 10996 12388 11036
rect 9364 10968 12388 10996
rect 12437 10999 12495 11005
rect 9364 10956 9370 10968
rect 12437 10965 12449 10999
rect 12483 10996 12495 10999
rect 12894 10996 12900 11008
rect 12483 10968 12900 10996
rect 12483 10965 12495 10968
rect 12437 10959 12495 10965
rect 12894 10956 12900 10968
rect 12952 10956 12958 11008
rect 13004 10996 13032 11036
rect 14476 11036 14780 11064
rect 14476 10996 14504 11036
rect 13004 10968 14504 10996
rect 14642 10956 14648 11008
rect 14700 10956 14706 11008
rect 14752 10996 14780 11036
rect 16040 11036 16252 11064
rect 16040 10996 16068 11036
rect 14752 10968 16068 10996
rect 16114 10956 16120 11008
rect 16172 10956 16178 11008
rect 16224 10996 16252 11036
rect 17512 11036 18981 11064
rect 17512 10996 17540 11036
rect 18969 11033 18981 11036
rect 19015 11033 19027 11067
rect 18969 11027 19027 11033
rect 16224 10968 17540 10996
rect 17589 10999 17647 11005
rect 17589 10965 17601 10999
rect 17635 10996 17647 10999
rect 17862 10996 17868 11008
rect 17635 10968 17868 10996
rect 17635 10965 17647 10968
rect 17589 10959 17647 10965
rect 17862 10956 17868 10968
rect 17920 10956 17926 11008
rect 17954 10956 17960 11008
rect 18012 10996 18018 11008
rect 19444 10996 19472 11104
rect 19521 11101 19533 11104
rect 19567 11101 19579 11135
rect 19521 11095 19579 11101
rect 21913 11135 21971 11141
rect 21913 11101 21925 11135
rect 21959 11132 21971 11135
rect 22370 11132 22376 11144
rect 21959 11104 22376 11132
rect 21959 11101 21971 11104
rect 21913 11095 21971 11101
rect 22370 11092 22376 11104
rect 22428 11092 22434 11144
rect 25409 11135 25467 11141
rect 25409 11101 25421 11135
rect 25455 11132 25467 11135
rect 25590 11132 25596 11144
rect 25455 11104 25596 11132
rect 25455 11101 25467 11104
rect 25409 11095 25467 11101
rect 25590 11092 25596 11104
rect 25648 11092 25654 11144
rect 26050 11092 26056 11144
rect 26108 11092 26114 11144
rect 23566 11024 23572 11076
rect 23624 11064 23630 11076
rect 24029 11067 24087 11073
rect 24029 11064 24041 11067
rect 23624 11036 24041 11064
rect 23624 11024 23630 11036
rect 24029 11033 24041 11036
rect 24075 11033 24087 11067
rect 24029 11027 24087 11033
rect 20438 10996 20444 11008
rect 18012 10968 20444 10996
rect 18012 10956 18018 10968
rect 20438 10956 20444 10968
rect 20496 10956 20502 11008
rect 21634 10956 21640 11008
rect 21692 10996 21698 11008
rect 22186 10996 22192 11008
rect 21692 10968 22192 10996
rect 21692 10956 21698 10968
rect 22186 10956 22192 10968
rect 22244 10956 22250 11008
rect 23658 10956 23664 11008
rect 23716 10996 23722 11008
rect 23937 10999 23995 11005
rect 23937 10996 23949 10999
rect 23716 10968 23949 10996
rect 23716 10956 23722 10968
rect 23937 10965 23949 10968
rect 23983 10965 23995 10999
rect 23937 10959 23995 10965
rect 25406 10956 25412 11008
rect 25464 10996 25470 11008
rect 27062 10996 27068 11008
rect 25464 10968 27068 10996
rect 25464 10956 25470 10968
rect 27062 10956 27068 10968
rect 27120 10956 27126 11008
rect 552 10906 27416 10928
rect 552 10854 3756 10906
rect 3808 10854 3820 10906
rect 3872 10854 3884 10906
rect 3936 10854 3948 10906
rect 4000 10854 4012 10906
rect 4064 10854 10472 10906
rect 10524 10854 10536 10906
rect 10588 10854 10600 10906
rect 10652 10854 10664 10906
rect 10716 10854 10728 10906
rect 10780 10854 17188 10906
rect 17240 10854 17252 10906
rect 17304 10854 17316 10906
rect 17368 10854 17380 10906
rect 17432 10854 17444 10906
rect 17496 10854 23904 10906
rect 23956 10854 23968 10906
rect 24020 10854 24032 10906
rect 24084 10854 24096 10906
rect 24148 10854 24160 10906
rect 24212 10854 27416 10906
rect 552 10832 27416 10854
rect 3510 10752 3516 10804
rect 3568 10752 3574 10804
rect 5353 10795 5411 10801
rect 5353 10761 5365 10795
rect 5399 10792 5411 10795
rect 6178 10792 6184 10804
rect 5399 10764 6184 10792
rect 5399 10761 5411 10764
rect 5353 10755 5411 10761
rect 6178 10752 6184 10764
rect 6236 10752 6242 10804
rect 11330 10752 11336 10804
rect 11388 10792 11394 10804
rect 12986 10792 12992 10804
rect 11388 10764 12992 10792
rect 11388 10752 11394 10764
rect 12986 10752 12992 10764
rect 13044 10752 13050 10804
rect 13446 10752 13452 10804
rect 13504 10792 13510 10804
rect 13633 10795 13691 10801
rect 13633 10792 13645 10795
rect 13504 10764 13645 10792
rect 13504 10752 13510 10764
rect 13633 10761 13645 10764
rect 13679 10761 13691 10795
rect 13633 10755 13691 10761
rect 14369 10795 14427 10801
rect 14369 10761 14381 10795
rect 14415 10792 14427 10795
rect 14642 10792 14648 10804
rect 14415 10764 14648 10792
rect 14415 10761 14427 10764
rect 14369 10755 14427 10761
rect 14642 10752 14648 10764
rect 14700 10752 14706 10804
rect 16209 10795 16267 10801
rect 16209 10761 16221 10795
rect 16255 10792 16267 10795
rect 16485 10795 16543 10801
rect 16485 10792 16497 10795
rect 16255 10764 16497 10792
rect 16255 10761 16267 10764
rect 16209 10755 16267 10761
rect 16485 10761 16497 10764
rect 16531 10761 16543 10795
rect 18874 10792 18880 10804
rect 16485 10755 16543 10761
rect 16960 10764 18880 10792
rect 5997 10727 6055 10733
rect 5997 10724 6009 10727
rect 5460 10696 6009 10724
rect 2958 10616 2964 10668
rect 3016 10656 3022 10668
rect 3016 10628 3372 10656
rect 3016 10616 3022 10628
rect 2501 10591 2559 10597
rect 2501 10557 2513 10591
rect 2547 10588 2559 10591
rect 2590 10588 2596 10600
rect 2547 10560 2596 10588
rect 2547 10557 2559 10560
rect 2501 10551 2559 10557
rect 2590 10548 2596 10560
rect 2648 10548 2654 10600
rect 2774 10548 2780 10600
rect 2832 10548 2838 10600
rect 3237 10591 3295 10597
rect 3237 10588 3249 10591
rect 2976 10560 3249 10588
rect 2976 10464 3004 10560
rect 3237 10557 3249 10560
rect 3283 10557 3295 10591
rect 3237 10551 3295 10557
rect 3344 10520 3372 10628
rect 3418 10548 3424 10600
rect 3476 10588 3482 10600
rect 3973 10591 4031 10597
rect 3973 10588 3985 10591
rect 3476 10560 3985 10588
rect 3476 10548 3482 10560
rect 3973 10557 3985 10560
rect 4019 10557 4031 10591
rect 3973 10551 4031 10557
rect 4157 10591 4215 10597
rect 4157 10557 4169 10591
rect 4203 10588 4215 10591
rect 4249 10591 4307 10597
rect 4249 10588 4261 10591
rect 4203 10560 4261 10588
rect 4203 10557 4215 10560
rect 4157 10551 4215 10557
rect 4249 10557 4261 10560
rect 4295 10557 4307 10591
rect 4249 10551 4307 10557
rect 4798 10548 4804 10600
rect 4856 10548 4862 10600
rect 3510 10520 3516 10532
rect 3344 10492 3516 10520
rect 3510 10480 3516 10492
rect 3568 10480 3574 10532
rect 5337 10523 5395 10529
rect 5337 10489 5349 10523
rect 5383 10520 5395 10523
rect 5460 10520 5488 10696
rect 5997 10693 6009 10696
rect 6043 10724 6055 10727
rect 6043 10696 6684 10724
rect 6043 10693 6055 10696
rect 5997 10687 6055 10693
rect 5629 10659 5687 10665
rect 5629 10625 5641 10659
rect 5675 10656 5687 10659
rect 6181 10659 6239 10665
rect 6181 10656 6193 10659
rect 5675 10628 6193 10656
rect 5675 10625 5687 10628
rect 5629 10619 5687 10625
rect 6181 10625 6193 10628
rect 6227 10625 6239 10659
rect 6181 10619 6239 10625
rect 6656 10600 6684 10696
rect 9766 10684 9772 10736
rect 9824 10724 9830 10736
rect 11238 10724 11244 10736
rect 9824 10696 11244 10724
rect 9824 10684 9830 10696
rect 11238 10684 11244 10696
rect 11296 10684 11302 10736
rect 11992 10696 12204 10724
rect 7006 10616 7012 10668
rect 7064 10616 7070 10668
rect 9140 10628 9444 10656
rect 9140 10600 9168 10628
rect 5813 10591 5871 10597
rect 5813 10588 5825 10591
rect 5552 10560 5825 10588
rect 5552 10529 5580 10560
rect 5813 10557 5825 10560
rect 5859 10588 5871 10591
rect 5994 10588 6000 10600
rect 5859 10560 6000 10588
rect 5859 10557 5871 10560
rect 5813 10551 5871 10557
rect 5994 10548 6000 10560
rect 6052 10548 6058 10600
rect 6089 10591 6147 10597
rect 6089 10557 6101 10591
rect 6135 10588 6147 10591
rect 6135 10560 6592 10588
rect 6135 10557 6147 10560
rect 6089 10551 6147 10557
rect 6564 10529 6592 10560
rect 6638 10548 6644 10600
rect 6696 10548 6702 10600
rect 6822 10548 6828 10600
rect 6880 10588 6886 10600
rect 7101 10591 7159 10597
rect 7101 10588 7113 10591
rect 6880 10560 7113 10588
rect 6880 10548 6886 10560
rect 7101 10557 7113 10560
rect 7147 10557 7159 10591
rect 7101 10551 7159 10557
rect 8938 10548 8944 10600
rect 8996 10548 9002 10600
rect 9033 10591 9091 10597
rect 9033 10557 9045 10591
rect 9079 10588 9091 10591
rect 9122 10588 9128 10600
rect 9079 10560 9128 10588
rect 9079 10557 9091 10560
rect 9033 10551 9091 10557
rect 9122 10548 9128 10560
rect 9180 10548 9186 10600
rect 9214 10548 9220 10600
rect 9272 10548 9278 10600
rect 9306 10548 9312 10600
rect 9364 10548 9370 10600
rect 9416 10597 9444 10628
rect 9858 10616 9864 10668
rect 9916 10656 9922 10668
rect 9916 10628 10640 10656
rect 9916 10616 9922 10628
rect 9401 10591 9459 10597
rect 9401 10557 9413 10591
rect 9447 10557 9459 10591
rect 9401 10551 9459 10557
rect 9490 10548 9496 10600
rect 9548 10588 9554 10600
rect 9585 10591 9643 10597
rect 9585 10588 9597 10591
rect 9548 10560 9597 10588
rect 9548 10548 9554 10560
rect 9585 10557 9597 10560
rect 9631 10557 9643 10591
rect 9585 10551 9643 10557
rect 10318 10548 10324 10600
rect 10376 10548 10382 10600
rect 10612 10597 10640 10628
rect 10597 10591 10655 10597
rect 10597 10557 10609 10591
rect 10643 10557 10655 10591
rect 10597 10551 10655 10557
rect 10870 10548 10876 10600
rect 10928 10548 10934 10600
rect 11238 10548 11244 10600
rect 11296 10588 11302 10600
rect 11992 10597 12020 10696
rect 12176 10656 12204 10696
rect 12250 10684 12256 10736
rect 12308 10724 12314 10736
rect 16960 10724 16988 10764
rect 18874 10752 18880 10764
rect 18932 10752 18938 10804
rect 20070 10752 20076 10804
rect 20128 10752 20134 10804
rect 20165 10795 20223 10801
rect 20165 10761 20177 10795
rect 20211 10792 20223 10795
rect 21082 10792 21088 10804
rect 20211 10764 21088 10792
rect 20211 10761 20223 10764
rect 20165 10755 20223 10761
rect 21082 10752 21088 10764
rect 21140 10752 21146 10804
rect 25406 10752 25412 10804
rect 25464 10752 25470 10804
rect 26878 10792 26884 10804
rect 25516 10764 26884 10792
rect 12308 10696 15608 10724
rect 12308 10684 12314 10696
rect 12802 10656 12808 10668
rect 12176 10628 12808 10656
rect 12802 10616 12808 10628
rect 12860 10616 12866 10668
rect 12894 10616 12900 10668
rect 12952 10616 12958 10668
rect 12986 10616 12992 10668
rect 13044 10656 13050 10668
rect 13044 10628 15516 10656
rect 13044 10616 13050 10628
rect 11701 10591 11759 10597
rect 11701 10588 11713 10591
rect 11296 10560 11713 10588
rect 11296 10548 11302 10560
rect 11701 10557 11713 10560
rect 11747 10557 11759 10591
rect 11701 10551 11759 10557
rect 11885 10591 11943 10597
rect 11885 10557 11897 10591
rect 11931 10557 11943 10591
rect 11885 10551 11943 10557
rect 11977 10591 12035 10597
rect 11977 10557 11989 10591
rect 12023 10557 12035 10591
rect 11977 10551 12035 10557
rect 5383 10492 5488 10520
rect 5537 10523 5595 10529
rect 5383 10489 5395 10492
rect 5337 10483 5395 10489
rect 5537 10489 5549 10523
rect 5583 10489 5595 10523
rect 5537 10483 5595 10489
rect 6549 10523 6607 10529
rect 6549 10489 6561 10523
rect 6595 10520 6607 10523
rect 7650 10520 7656 10532
rect 6595 10492 7656 10520
rect 6595 10489 6607 10492
rect 6549 10483 6607 10489
rect 7650 10480 7656 10492
rect 7708 10480 7714 10532
rect 8956 10520 8984 10548
rect 11900 10520 11928 10551
rect 12158 10548 12164 10600
rect 12216 10548 12222 10600
rect 12265 10591 12323 10597
rect 12265 10557 12277 10591
rect 12311 10588 12323 10591
rect 12912 10588 12940 10616
rect 13081 10591 13139 10597
rect 13081 10588 13093 10591
rect 12311 10560 12756 10588
rect 12912 10560 13093 10588
rect 12311 10557 12323 10560
rect 12265 10551 12323 10557
rect 12066 10520 12072 10532
rect 8956 10492 12072 10520
rect 12066 10480 12072 10492
rect 12124 10480 12130 10532
rect 12728 10520 12756 10560
rect 13081 10557 13093 10560
rect 13127 10557 13139 10591
rect 13081 10551 13139 10557
rect 13262 10548 13268 10600
rect 13320 10548 13326 10600
rect 13817 10591 13875 10597
rect 13817 10557 13829 10591
rect 13863 10557 13875 10591
rect 13817 10551 13875 10557
rect 13173 10523 13231 10529
rect 13173 10520 13185 10523
rect 12728 10492 13185 10520
rect 13173 10489 13185 10492
rect 13219 10489 13231 10523
rect 13832 10520 13860 10551
rect 13998 10548 14004 10600
rect 14056 10548 14062 10600
rect 14093 10591 14151 10597
rect 14093 10557 14105 10591
rect 14139 10588 14151 10591
rect 14274 10588 14280 10600
rect 14139 10560 14280 10588
rect 14139 10557 14151 10560
rect 14093 10551 14151 10557
rect 14274 10548 14280 10560
rect 14332 10548 14338 10600
rect 14734 10588 14740 10600
rect 14568 10560 14740 10588
rect 14568 10532 14596 10560
rect 14734 10548 14740 10560
rect 14792 10588 14798 10600
rect 15378 10588 15384 10600
rect 14792 10560 15384 10588
rect 14792 10548 14798 10560
rect 15378 10548 15384 10560
rect 15436 10548 15442 10600
rect 13832 10492 14228 10520
rect 13173 10483 13231 10489
rect 2314 10412 2320 10464
rect 2372 10452 2378 10464
rect 2593 10455 2651 10461
rect 2593 10452 2605 10455
rect 2372 10424 2605 10452
rect 2372 10412 2378 10424
rect 2593 10421 2605 10424
rect 2639 10421 2651 10455
rect 2593 10415 2651 10421
rect 2958 10412 2964 10464
rect 3016 10412 3022 10464
rect 3329 10455 3387 10461
rect 3329 10421 3341 10455
rect 3375 10452 3387 10455
rect 3602 10452 3608 10464
rect 3375 10424 3608 10452
rect 3375 10421 3387 10424
rect 3329 10415 3387 10421
rect 3602 10412 3608 10424
rect 3660 10452 3666 10464
rect 3973 10455 4031 10461
rect 3973 10452 3985 10455
rect 3660 10424 3985 10452
rect 3660 10412 3666 10424
rect 3973 10421 3985 10424
rect 4019 10421 4031 10455
rect 3973 10415 4031 10421
rect 5074 10412 5080 10464
rect 5132 10452 5138 10464
rect 5169 10455 5227 10461
rect 5169 10452 5181 10455
rect 5132 10424 5181 10452
rect 5132 10412 5138 10424
rect 5169 10421 5181 10424
rect 5215 10421 5227 10455
rect 5169 10415 5227 10421
rect 6270 10412 6276 10464
rect 6328 10452 6334 10464
rect 6457 10455 6515 10461
rect 6457 10452 6469 10455
rect 6328 10424 6469 10452
rect 6328 10412 6334 10424
rect 6457 10421 6469 10424
rect 6503 10421 6515 10455
rect 6457 10415 6515 10421
rect 7466 10412 7472 10464
rect 7524 10412 7530 10464
rect 8757 10455 8815 10461
rect 8757 10421 8769 10455
rect 8803 10452 8815 10455
rect 8846 10452 8852 10464
rect 8803 10424 8852 10452
rect 8803 10421 8815 10424
rect 8757 10415 8815 10421
rect 8846 10412 8852 10424
rect 8904 10412 8910 10464
rect 8938 10412 8944 10464
rect 8996 10452 9002 10464
rect 9493 10455 9551 10461
rect 9493 10452 9505 10455
rect 8996 10424 9505 10452
rect 8996 10412 9002 10424
rect 9493 10421 9505 10424
rect 9539 10421 9551 10455
rect 9493 10415 9551 10421
rect 10134 10412 10140 10464
rect 10192 10412 10198 10464
rect 10505 10455 10563 10461
rect 10505 10421 10517 10455
rect 10551 10452 10563 10455
rect 11054 10452 11060 10464
rect 10551 10424 11060 10452
rect 10551 10421 10563 10424
rect 10505 10415 10563 10421
rect 11054 10412 11060 10424
rect 11112 10412 11118 10464
rect 11146 10412 11152 10464
rect 11204 10452 11210 10464
rect 11517 10455 11575 10461
rect 11517 10452 11529 10455
rect 11204 10424 11529 10452
rect 11204 10412 11210 10424
rect 11517 10421 11529 10424
rect 11563 10421 11575 10455
rect 11517 10415 11575 10421
rect 12250 10412 12256 10464
rect 12308 10452 12314 10464
rect 14200 10461 14228 10492
rect 14550 10480 14556 10532
rect 14608 10480 14614 10532
rect 15488 10520 15516 10628
rect 15580 10597 15608 10696
rect 16316 10696 16988 10724
rect 15565 10591 15623 10597
rect 15565 10557 15577 10591
rect 15611 10557 15623 10591
rect 15565 10551 15623 10557
rect 15654 10548 15660 10600
rect 15712 10548 15718 10600
rect 15838 10548 15844 10600
rect 15896 10548 15902 10600
rect 15933 10591 15991 10597
rect 15933 10557 15945 10591
rect 15979 10588 15991 10591
rect 16206 10588 16212 10600
rect 15979 10560 16212 10588
rect 15979 10557 15991 10560
rect 15933 10551 15991 10557
rect 16206 10548 16212 10560
rect 16264 10548 16270 10600
rect 16022 10520 16028 10532
rect 15488 10492 16028 10520
rect 16022 10480 16028 10492
rect 16080 10480 16086 10532
rect 16316 10520 16344 10696
rect 17034 10684 17040 10736
rect 17092 10684 17098 10736
rect 17954 10724 17960 10736
rect 17696 10696 17960 10724
rect 17052 10656 17080 10684
rect 17405 10659 17463 10665
rect 17405 10656 17417 10659
rect 17052 10628 17417 10656
rect 17405 10625 17417 10628
rect 17451 10625 17463 10659
rect 17405 10619 17463 10625
rect 17034 10548 17040 10600
rect 17092 10588 17098 10600
rect 17497 10591 17555 10597
rect 17497 10588 17509 10591
rect 17092 10560 17509 10588
rect 17092 10548 17098 10560
rect 17497 10557 17509 10560
rect 17543 10557 17555 10591
rect 17696 10588 17724 10696
rect 17954 10684 17960 10696
rect 18012 10684 18018 10736
rect 20438 10684 20444 10736
rect 20496 10724 20502 10736
rect 20625 10727 20683 10733
rect 20625 10724 20637 10727
rect 20496 10696 20637 10724
rect 20496 10684 20502 10696
rect 20625 10693 20637 10696
rect 20671 10693 20683 10727
rect 25516 10724 25544 10764
rect 26878 10752 26884 10764
rect 26936 10752 26942 10804
rect 20625 10687 20683 10693
rect 25148 10696 25544 10724
rect 17770 10616 17776 10668
rect 17828 10656 17834 10668
rect 18693 10659 18751 10665
rect 18693 10656 18705 10659
rect 17828 10628 18705 10656
rect 17828 10616 17834 10628
rect 18693 10625 18705 10628
rect 18739 10625 18751 10659
rect 18693 10619 18751 10625
rect 22094 10616 22100 10668
rect 22152 10616 22158 10668
rect 22462 10616 22468 10668
rect 22520 10656 22526 10668
rect 22830 10656 22836 10668
rect 22520 10628 22836 10656
rect 22520 10616 22526 10628
rect 22830 10616 22836 10628
rect 22888 10656 22894 10668
rect 24302 10656 24308 10668
rect 22888 10628 24308 10656
rect 22888 10616 22894 10628
rect 17696 10560 17816 10588
rect 17497 10551 17555 10557
rect 17788 10529 17816 10560
rect 17862 10548 17868 10600
rect 17920 10548 17926 10600
rect 18141 10591 18199 10597
rect 18141 10557 18153 10591
rect 18187 10557 18199 10591
rect 18141 10551 18199 10557
rect 17773 10523 17831 10529
rect 16224 10492 16344 10520
rect 16408 10492 17724 10520
rect 14366 10461 14372 10464
rect 12345 10455 12403 10461
rect 12345 10452 12357 10455
rect 12308 10424 12357 10452
rect 12308 10412 12314 10424
rect 12345 10421 12357 10424
rect 12391 10421 12403 10455
rect 12345 10415 12403 10421
rect 14185 10455 14243 10461
rect 14185 10421 14197 10455
rect 14231 10421 14243 10455
rect 14185 10415 14243 10421
rect 14353 10455 14372 10461
rect 14353 10421 14365 10455
rect 14353 10415 14372 10421
rect 14366 10412 14372 10415
rect 14424 10412 14430 10464
rect 15378 10412 15384 10464
rect 15436 10412 15442 10464
rect 16224 10461 16252 10492
rect 16408 10461 16436 10492
rect 16224 10455 16283 10461
rect 16224 10424 16237 10455
rect 16225 10421 16237 10424
rect 16271 10421 16283 10455
rect 16225 10415 16283 10421
rect 16393 10455 16451 10461
rect 16393 10421 16405 10455
rect 16439 10421 16451 10455
rect 16393 10415 16451 10421
rect 17218 10412 17224 10464
rect 17276 10412 17282 10464
rect 17696 10452 17724 10492
rect 17773 10489 17785 10523
rect 17819 10489 17831 10523
rect 18156 10520 18184 10551
rect 18230 10548 18236 10600
rect 18288 10588 18294 10600
rect 18325 10591 18383 10597
rect 18325 10588 18337 10591
rect 18288 10560 18337 10588
rect 18288 10548 18294 10560
rect 18325 10557 18337 10560
rect 18371 10557 18383 10591
rect 18325 10551 18383 10557
rect 18414 10548 18420 10600
rect 18472 10548 18478 10600
rect 20346 10548 20352 10600
rect 20404 10548 20410 10600
rect 20441 10591 20499 10597
rect 20441 10557 20453 10591
rect 20487 10588 20499 10591
rect 20990 10588 20996 10600
rect 20487 10560 20996 10588
rect 20487 10557 20499 10560
rect 20441 10551 20499 10557
rect 20990 10548 20996 10560
rect 21048 10548 21054 10600
rect 22002 10548 22008 10600
rect 22060 10548 22066 10600
rect 22741 10591 22799 10597
rect 22741 10557 22753 10591
rect 22787 10588 22799 10591
rect 23109 10591 23167 10597
rect 23109 10588 23121 10591
rect 22787 10560 23121 10588
rect 22787 10557 22799 10560
rect 22741 10551 22799 10557
rect 23109 10557 23121 10560
rect 23155 10557 23167 10591
rect 23109 10551 23167 10557
rect 23201 10591 23259 10597
rect 23201 10557 23213 10591
rect 23247 10557 23259 10591
rect 23201 10551 23259 10557
rect 17773 10483 17831 10489
rect 17880 10492 18184 10520
rect 17880 10452 17908 10492
rect 18506 10480 18512 10532
rect 18564 10520 18570 10532
rect 18938 10523 18996 10529
rect 18938 10520 18950 10523
rect 18564 10492 18950 10520
rect 18564 10480 18570 10492
rect 18938 10489 18950 10492
rect 18984 10489 18996 10523
rect 18938 10483 18996 10489
rect 19886 10480 19892 10532
rect 19944 10520 19950 10532
rect 20165 10523 20223 10529
rect 20165 10520 20177 10523
rect 19944 10492 20177 10520
rect 19944 10480 19950 10492
rect 20165 10489 20177 10492
rect 20211 10489 20223 10523
rect 20165 10483 20223 10489
rect 21760 10523 21818 10529
rect 21760 10489 21772 10523
rect 21806 10520 21818 10523
rect 22833 10523 22891 10529
rect 22833 10520 22845 10523
rect 21806 10492 22845 10520
rect 21806 10489 21818 10492
rect 21760 10483 21818 10489
rect 22833 10489 22845 10492
rect 22879 10489 22891 10523
rect 23216 10520 23244 10551
rect 23290 10548 23296 10600
rect 23348 10548 23354 10600
rect 23492 10597 23520 10628
rect 24302 10616 24308 10628
rect 24360 10656 24366 10668
rect 24762 10656 24768 10668
rect 24360 10628 24768 10656
rect 24360 10616 24366 10628
rect 24762 10616 24768 10628
rect 24820 10616 24826 10668
rect 23477 10591 23535 10597
rect 23477 10557 23489 10591
rect 23523 10557 23535 10591
rect 23477 10551 23535 10557
rect 23566 10548 23572 10600
rect 23624 10588 23630 10600
rect 25148 10597 25176 10696
rect 24213 10591 24271 10597
rect 24213 10588 24225 10591
rect 23624 10560 24225 10588
rect 23624 10548 23630 10560
rect 24213 10557 24225 10560
rect 24259 10557 24271 10591
rect 24213 10551 24271 10557
rect 25133 10591 25191 10597
rect 25133 10557 25145 10591
rect 25179 10557 25191 10591
rect 25133 10551 25191 10557
rect 25225 10591 25283 10597
rect 25225 10557 25237 10591
rect 25271 10588 25283 10591
rect 25314 10588 25320 10600
rect 25271 10560 25320 10588
rect 25271 10557 25283 10560
rect 25225 10551 25283 10557
rect 25314 10548 25320 10560
rect 25372 10548 25378 10600
rect 25501 10591 25559 10597
rect 25501 10557 25513 10591
rect 25547 10588 25559 10591
rect 25590 10588 25596 10600
rect 25547 10560 25596 10588
rect 25547 10557 25559 10560
rect 25501 10551 25559 10557
rect 25590 10548 25596 10560
rect 25648 10548 25654 10600
rect 23842 10520 23848 10532
rect 23216 10492 23848 10520
rect 22833 10483 22891 10489
rect 23842 10480 23848 10492
rect 23900 10480 23906 10532
rect 24762 10480 24768 10532
rect 24820 10520 24826 10532
rect 25409 10523 25467 10529
rect 25409 10520 25421 10523
rect 24820 10492 25421 10520
rect 24820 10480 24826 10492
rect 25409 10489 25421 10492
rect 25455 10489 25467 10523
rect 25746 10523 25804 10529
rect 25746 10520 25758 10523
rect 25409 10483 25467 10489
rect 25516 10492 25758 10520
rect 25516 10464 25544 10492
rect 25746 10489 25758 10492
rect 25792 10489 25804 10523
rect 25746 10483 25804 10489
rect 17696 10424 17908 10452
rect 17954 10412 17960 10464
rect 18012 10412 18018 10464
rect 24854 10412 24860 10464
rect 24912 10412 24918 10464
rect 24946 10412 24952 10464
rect 25004 10412 25010 10464
rect 25498 10412 25504 10464
rect 25556 10412 25562 10464
rect 552 10362 27576 10384
rect 552 10310 7114 10362
rect 7166 10310 7178 10362
rect 7230 10310 7242 10362
rect 7294 10310 7306 10362
rect 7358 10310 7370 10362
rect 7422 10310 13830 10362
rect 13882 10310 13894 10362
rect 13946 10310 13958 10362
rect 14010 10310 14022 10362
rect 14074 10310 14086 10362
rect 14138 10310 20546 10362
rect 20598 10310 20610 10362
rect 20662 10310 20674 10362
rect 20726 10310 20738 10362
rect 20790 10310 20802 10362
rect 20854 10310 27262 10362
rect 27314 10310 27326 10362
rect 27378 10310 27390 10362
rect 27442 10310 27454 10362
rect 27506 10310 27518 10362
rect 27570 10310 27576 10362
rect 552 10288 27576 10310
rect 3326 10248 3332 10260
rect 3252 10220 3332 10248
rect 2866 10180 2872 10192
rect 2792 10152 2872 10180
rect 2409 10115 2467 10121
rect 2409 10081 2421 10115
rect 2455 10112 2467 10115
rect 2590 10112 2596 10124
rect 2455 10084 2596 10112
rect 2455 10081 2467 10084
rect 2409 10075 2467 10081
rect 2590 10072 2596 10084
rect 2648 10072 2654 10124
rect 2792 10121 2820 10152
rect 2866 10140 2872 10152
rect 2924 10140 2930 10192
rect 3044 10183 3102 10189
rect 3044 10149 3056 10183
rect 3090 10180 3102 10183
rect 3252 10180 3280 10220
rect 3326 10208 3332 10220
rect 3384 10208 3390 10260
rect 4157 10251 4215 10257
rect 4157 10217 4169 10251
rect 4203 10248 4215 10251
rect 4798 10248 4804 10260
rect 4203 10220 4804 10248
rect 4203 10217 4215 10220
rect 4157 10211 4215 10217
rect 4798 10208 4804 10220
rect 4856 10208 4862 10260
rect 6638 10208 6644 10260
rect 6696 10248 6702 10260
rect 7009 10251 7067 10257
rect 7009 10248 7021 10251
rect 6696 10220 7021 10248
rect 6696 10208 6702 10220
rect 7009 10217 7021 10220
rect 7055 10217 7067 10251
rect 7009 10211 7067 10217
rect 7466 10208 7472 10260
rect 7524 10248 7530 10260
rect 7524 10220 10272 10248
rect 7524 10208 7530 10220
rect 7285 10183 7343 10189
rect 3090 10152 3280 10180
rect 4448 10152 7236 10180
rect 3090 10149 3102 10152
rect 3044 10143 3102 10149
rect 2777 10115 2835 10121
rect 2777 10081 2789 10115
rect 2823 10081 2835 10115
rect 4448 10112 4476 10152
rect 2777 10075 2835 10081
rect 2884 10084 4476 10112
rect 4516 10115 4574 10121
rect 2225 10047 2283 10053
rect 2225 10013 2237 10047
rect 2271 10013 2283 10047
rect 2225 10007 2283 10013
rect 2240 9976 2268 10007
rect 2314 10004 2320 10056
rect 2372 10004 2378 10056
rect 2501 10047 2559 10053
rect 2501 10013 2513 10047
rect 2547 10044 2559 10047
rect 2682 10044 2688 10056
rect 2547 10016 2688 10044
rect 2547 10013 2559 10016
rect 2501 10007 2559 10013
rect 2682 10004 2688 10016
rect 2740 10004 2746 10056
rect 2884 10044 2912 10084
rect 4516 10081 4528 10115
rect 4562 10112 4574 10115
rect 4890 10112 4896 10124
rect 4562 10084 4896 10112
rect 4562 10081 4574 10084
rect 4516 10075 4574 10081
rect 4890 10072 4896 10084
rect 4948 10072 4954 10124
rect 6270 10072 6276 10124
rect 6328 10072 6334 10124
rect 6914 10072 6920 10124
rect 6972 10072 6978 10124
rect 7101 10115 7159 10121
rect 7101 10081 7113 10115
rect 7147 10081 7159 10115
rect 7101 10075 7159 10081
rect 2792 10016 2912 10044
rect 2792 9976 2820 10016
rect 4246 10004 4252 10056
rect 4304 10004 4310 10056
rect 6822 10044 6828 10056
rect 5644 10016 6828 10044
rect 5644 9985 5672 10016
rect 6822 10004 6828 10016
rect 6880 10044 6886 10056
rect 7116 10044 7144 10075
rect 6880 10016 7144 10044
rect 7208 10044 7236 10152
rect 7285 10149 7297 10183
rect 7331 10180 7343 10183
rect 7650 10180 7656 10192
rect 7331 10152 7656 10180
rect 7331 10149 7343 10152
rect 7285 10143 7343 10149
rect 7650 10140 7656 10152
rect 7708 10140 7714 10192
rect 8588 10121 8616 10220
rect 9668 10183 9726 10189
rect 8680 10152 9168 10180
rect 8680 10124 8708 10152
rect 9140 10124 9168 10152
rect 9668 10149 9680 10183
rect 9714 10180 9726 10183
rect 10134 10180 10140 10192
rect 9714 10152 10140 10180
rect 9714 10149 9726 10152
rect 9668 10143 9726 10149
rect 10134 10140 10140 10152
rect 10192 10140 10198 10192
rect 7377 10115 7435 10121
rect 7377 10081 7389 10115
rect 7423 10112 7435 10115
rect 7469 10115 7527 10121
rect 7469 10112 7481 10115
rect 7423 10084 7481 10112
rect 7423 10081 7435 10084
rect 7377 10075 7435 10081
rect 7469 10081 7481 10084
rect 7515 10081 7527 10115
rect 8573 10115 8631 10121
rect 7469 10075 7527 10081
rect 7944 10084 8524 10112
rect 7944 10044 7972 10084
rect 7208 10016 7972 10044
rect 6880 10004 6886 10016
rect 8018 10004 8024 10056
rect 8076 10004 8082 10056
rect 8496 10044 8524 10084
rect 8573 10081 8585 10115
rect 8619 10081 8631 10115
rect 8573 10075 8631 10081
rect 8662 10072 8668 10124
rect 8720 10072 8726 10124
rect 8849 10115 8907 10121
rect 8849 10081 8861 10115
rect 8895 10081 8907 10115
rect 8849 10075 8907 10081
rect 8496 10016 8708 10044
rect 2240 9948 2820 9976
rect 5629 9979 5687 9985
rect 5629 9945 5641 9979
rect 5675 9945 5687 9979
rect 8478 9976 8484 9988
rect 5629 9939 5687 9945
rect 5736 9948 8484 9976
rect 2682 9868 2688 9920
rect 2740 9868 2746 9920
rect 3510 9868 3516 9920
rect 3568 9908 3574 9920
rect 5736 9908 5764 9948
rect 8478 9936 8484 9948
rect 8536 9936 8542 9988
rect 8680 9976 8708 10016
rect 8754 10004 8760 10056
rect 8812 10044 8818 10056
rect 8864 10044 8892 10075
rect 8938 10072 8944 10124
rect 8996 10072 9002 10124
rect 9122 10072 9128 10124
rect 9180 10072 9186 10124
rect 9309 10115 9367 10121
rect 9309 10081 9321 10115
rect 9355 10112 9367 10115
rect 10042 10112 10048 10124
rect 9355 10084 10048 10112
rect 9355 10081 9367 10084
rect 9309 10075 9367 10081
rect 10042 10072 10048 10084
rect 10100 10072 10106 10124
rect 10244 10112 10272 10220
rect 10318 10208 10324 10260
rect 10376 10248 10382 10260
rect 10965 10251 11023 10257
rect 10965 10248 10977 10251
rect 10376 10220 10977 10248
rect 10376 10208 10382 10220
rect 10965 10217 10977 10220
rect 11011 10217 11023 10251
rect 10965 10211 11023 10217
rect 11517 10251 11575 10257
rect 11517 10217 11529 10251
rect 11563 10248 11575 10251
rect 11606 10248 11612 10260
rect 11563 10220 11612 10248
rect 11563 10217 11575 10220
rect 11517 10211 11575 10217
rect 11606 10208 11612 10220
rect 11664 10208 11670 10260
rect 11882 10208 11888 10260
rect 11940 10248 11946 10260
rect 14182 10248 14188 10260
rect 11940 10220 14188 10248
rect 11940 10208 11946 10220
rect 14182 10208 14188 10220
rect 14240 10208 14246 10260
rect 15838 10248 15844 10260
rect 14936 10220 15844 10248
rect 10410 10140 10416 10192
rect 10468 10180 10474 10192
rect 11117 10183 11175 10189
rect 11117 10180 11129 10183
rect 10468 10152 11129 10180
rect 10468 10140 10474 10152
rect 11117 10149 11129 10152
rect 11163 10149 11175 10183
rect 11117 10143 11175 10149
rect 11330 10140 11336 10192
rect 11388 10140 11394 10192
rect 12237 10183 12295 10189
rect 12237 10180 12249 10183
rect 11900 10152 12249 10180
rect 11900 10124 11928 10152
rect 12237 10149 12249 10152
rect 12283 10180 12295 10183
rect 12342 10180 12348 10192
rect 12283 10152 12348 10180
rect 12283 10149 12295 10152
rect 12237 10143 12295 10149
rect 12342 10140 12348 10152
rect 12400 10140 12406 10192
rect 12437 10183 12495 10189
rect 12437 10149 12449 10183
rect 12483 10149 12495 10183
rect 12437 10143 12495 10149
rect 11701 10115 11759 10121
rect 10244 10084 11284 10112
rect 9214 10044 9220 10056
rect 8812 10016 9220 10044
rect 8812 10004 8818 10016
rect 9214 10004 9220 10016
rect 9272 10004 9278 10056
rect 9398 10004 9404 10056
rect 9456 10004 9462 10056
rect 8680 9948 9444 9976
rect 3568 9880 5764 9908
rect 6825 9911 6883 9917
rect 3568 9868 3574 9880
rect 6825 9877 6837 9911
rect 6871 9908 6883 9911
rect 6914 9908 6920 9920
rect 6871 9880 6920 9908
rect 6871 9877 6883 9880
rect 6825 9871 6883 9877
rect 6914 9868 6920 9880
rect 6972 9868 6978 9920
rect 8386 9868 8392 9920
rect 8444 9868 8450 9920
rect 9030 9868 9036 9920
rect 9088 9908 9094 9920
rect 9309 9911 9367 9917
rect 9309 9908 9321 9911
rect 9088 9880 9321 9908
rect 9088 9868 9094 9880
rect 9309 9877 9321 9880
rect 9355 9877 9367 9911
rect 9416 9908 9444 9948
rect 9766 9908 9772 9920
rect 9416 9880 9772 9908
rect 9309 9871 9367 9877
rect 9766 9868 9772 9880
rect 9824 9868 9830 9920
rect 10318 9868 10324 9920
rect 10376 9908 10382 9920
rect 10781 9911 10839 9917
rect 10781 9908 10793 9911
rect 10376 9880 10793 9908
rect 10376 9868 10382 9880
rect 10781 9877 10793 9880
rect 10827 9908 10839 9911
rect 10870 9908 10876 9920
rect 10827 9880 10876 9908
rect 10827 9877 10839 9880
rect 10781 9871 10839 9877
rect 10870 9868 10876 9880
rect 10928 9868 10934 9920
rect 11146 9868 11152 9920
rect 11204 9868 11210 9920
rect 11256 9908 11284 10084
rect 11701 10081 11713 10115
rect 11747 10081 11759 10115
rect 11701 10075 11759 10081
rect 11716 10044 11744 10075
rect 11882 10072 11888 10124
rect 11940 10072 11946 10124
rect 11974 10072 11980 10124
rect 12032 10072 12038 10124
rect 12452 10044 12480 10143
rect 12802 10140 12808 10192
rect 12860 10180 12866 10192
rect 13262 10180 13268 10192
rect 12860 10152 13268 10180
rect 12860 10140 12866 10152
rect 13004 10124 13032 10152
rect 13262 10140 13268 10152
rect 13320 10140 13326 10192
rect 12986 10072 12992 10124
rect 13044 10072 13050 10124
rect 13170 10072 13176 10124
rect 13228 10072 13234 10124
rect 14642 10072 14648 10124
rect 14700 10072 14706 10124
rect 14936 10121 14964 10220
rect 15838 10208 15844 10220
rect 15896 10208 15902 10260
rect 16022 10208 16028 10260
rect 16080 10248 16086 10260
rect 16393 10251 16451 10257
rect 16080 10220 16252 10248
rect 16080 10208 16086 10220
rect 15286 10140 15292 10192
rect 15344 10180 15350 10192
rect 16224 10180 16252 10220
rect 16393 10217 16405 10251
rect 16439 10248 16451 10251
rect 17034 10248 17040 10260
rect 16439 10220 17040 10248
rect 16439 10217 16451 10220
rect 16393 10211 16451 10217
rect 17034 10208 17040 10220
rect 17092 10208 17098 10260
rect 18322 10248 18328 10260
rect 17420 10220 18328 10248
rect 17420 10180 17448 10220
rect 18322 10208 18328 10220
rect 18380 10248 18386 10260
rect 18769 10251 18827 10257
rect 18380 10220 18552 10248
rect 18380 10208 18386 10220
rect 15344 10152 16160 10180
rect 16224 10152 17448 10180
rect 17528 10183 17586 10189
rect 15344 10140 15350 10152
rect 14737 10115 14795 10121
rect 14737 10081 14749 10115
rect 14783 10081 14795 10115
rect 14737 10075 14795 10081
rect 14921 10115 14979 10121
rect 14921 10081 14933 10115
rect 14967 10081 14979 10115
rect 14921 10075 14979 10081
rect 15013 10115 15071 10121
rect 15013 10081 15025 10115
rect 15059 10112 15071 10115
rect 16022 10112 16028 10124
rect 15059 10084 16028 10112
rect 15059 10081 15071 10084
rect 15013 10075 15071 10081
rect 12526 10044 12532 10056
rect 11716 10016 12112 10044
rect 12452 10016 12532 10044
rect 12084 9985 12112 10016
rect 12526 10004 12532 10016
rect 12584 10044 12590 10056
rect 14550 10044 14556 10056
rect 12584 10016 14556 10044
rect 12584 10004 12590 10016
rect 14550 10004 14556 10016
rect 14608 10004 14614 10056
rect 14752 10044 14780 10075
rect 16022 10072 16028 10084
rect 16080 10072 16086 10124
rect 16132 10121 16160 10152
rect 17528 10149 17540 10183
rect 17574 10180 17586 10183
rect 17954 10180 17960 10192
rect 17574 10152 17960 10180
rect 17574 10149 17586 10152
rect 17528 10143 17586 10149
rect 17954 10140 17960 10152
rect 18012 10140 18018 10192
rect 18414 10180 18420 10192
rect 18064 10152 18420 10180
rect 16117 10115 16175 10121
rect 16117 10081 16129 10115
rect 16163 10081 16175 10115
rect 16117 10075 16175 10081
rect 16206 10072 16212 10124
rect 16264 10072 16270 10124
rect 18064 10121 18092 10152
rect 18414 10140 18420 10152
rect 18472 10140 18478 10192
rect 18524 10180 18552 10220
rect 18769 10217 18781 10251
rect 18815 10248 18827 10251
rect 18874 10248 18880 10260
rect 18815 10220 18880 10248
rect 18815 10217 18827 10220
rect 18769 10211 18827 10217
rect 18874 10208 18880 10220
rect 18932 10208 18938 10260
rect 22005 10251 22063 10257
rect 22005 10217 22017 10251
rect 22051 10248 22063 10251
rect 23290 10248 23296 10260
rect 22051 10220 23296 10248
rect 22051 10217 22063 10220
rect 22005 10211 22063 10217
rect 23290 10208 23296 10220
rect 23348 10208 23354 10260
rect 23474 10208 23480 10260
rect 23532 10248 23538 10260
rect 26142 10248 26148 10260
rect 23532 10220 24992 10248
rect 23532 10208 23538 10220
rect 18969 10183 19027 10189
rect 18969 10180 18981 10183
rect 18524 10152 18981 10180
rect 18969 10149 18981 10152
rect 19015 10149 19027 10183
rect 18969 10143 19027 10149
rect 21542 10140 21548 10192
rect 21600 10180 21606 10192
rect 21637 10183 21695 10189
rect 21637 10180 21649 10183
rect 21600 10152 21649 10180
rect 21600 10140 21606 10152
rect 21637 10149 21649 10152
rect 21683 10149 21695 10183
rect 21637 10143 21695 10149
rect 21821 10183 21879 10189
rect 21821 10149 21833 10183
rect 21867 10180 21879 10183
rect 24854 10180 24860 10192
rect 21867 10152 24860 10180
rect 21867 10149 21879 10152
rect 21821 10143 21879 10149
rect 16301 10115 16359 10121
rect 16301 10081 16313 10115
rect 16347 10081 16359 10115
rect 16301 10075 16359 10081
rect 18049 10115 18107 10121
rect 18049 10081 18061 10115
rect 18095 10081 18107 10115
rect 18049 10075 18107 10081
rect 15562 10044 15568 10056
rect 14752 10016 15568 10044
rect 15562 10004 15568 10016
rect 15620 10004 15626 10056
rect 15654 10004 15660 10056
rect 15712 10004 15718 10056
rect 12069 9979 12127 9985
rect 12069 9945 12081 9979
rect 12115 9945 12127 9979
rect 15580 9976 15608 10004
rect 16316 9976 16344 10075
rect 18138 10072 18144 10124
rect 18196 10072 18202 10124
rect 18325 10115 18383 10121
rect 18325 10081 18337 10115
rect 18371 10112 18383 10115
rect 18371 10084 18644 10112
rect 18371 10081 18383 10084
rect 18325 10075 18383 10081
rect 17770 10004 17776 10056
rect 17828 10004 17834 10056
rect 18506 10004 18512 10056
rect 18564 10004 18570 10056
rect 16390 9976 16396 9988
rect 12069 9939 12127 9945
rect 12176 9948 12388 9976
rect 15580 9948 16396 9976
rect 12176 9908 12204 9948
rect 11256 9880 12204 9908
rect 12250 9868 12256 9920
rect 12308 9868 12314 9920
rect 12360 9908 12388 9948
rect 16390 9936 16396 9948
rect 16448 9936 16454 9988
rect 12894 9908 12900 9920
rect 12360 9880 12900 9908
rect 12894 9868 12900 9880
rect 12952 9868 12958 9920
rect 12989 9911 13047 9917
rect 12989 9877 13001 9911
rect 13035 9908 13047 9911
rect 13262 9908 13268 9920
rect 13035 9880 13268 9908
rect 13035 9877 13047 9880
rect 12989 9871 13047 9877
rect 13262 9868 13268 9880
rect 13320 9868 13326 9920
rect 14461 9911 14519 9917
rect 14461 9877 14473 9911
rect 14507 9908 14519 9911
rect 14918 9908 14924 9920
rect 14507 9880 14924 9908
rect 14507 9877 14519 9880
rect 14461 9871 14519 9877
rect 14918 9868 14924 9880
rect 14976 9868 14982 9920
rect 15105 9911 15163 9917
rect 15105 9877 15117 9911
rect 15151 9908 15163 9911
rect 15194 9908 15200 9920
rect 15151 9880 15200 9908
rect 15151 9877 15163 9880
rect 15105 9871 15163 9877
rect 15194 9868 15200 9880
rect 15252 9868 15258 9920
rect 17034 9868 17040 9920
rect 17092 9908 17098 9920
rect 17788 9908 17816 10004
rect 18616 9985 18644 10084
rect 20070 10072 20076 10124
rect 20128 10072 20134 10124
rect 22278 10072 22284 10124
rect 22336 10112 22342 10124
rect 22373 10115 22431 10121
rect 22373 10112 22385 10115
rect 22336 10084 22385 10112
rect 22336 10072 22342 10084
rect 22373 10081 22385 10084
rect 22419 10081 22431 10115
rect 22373 10075 22431 10081
rect 22465 10115 22523 10121
rect 22465 10081 22477 10115
rect 22511 10081 22523 10115
rect 22465 10075 22523 10081
rect 22480 10044 22508 10075
rect 22554 10072 22560 10124
rect 22612 10072 22618 10124
rect 22741 10115 22799 10121
rect 22741 10081 22753 10115
rect 22787 10112 22799 10115
rect 22830 10112 22836 10124
rect 22787 10084 22836 10112
rect 22787 10081 22799 10084
rect 22741 10075 22799 10081
rect 22830 10072 22836 10084
rect 22888 10072 22894 10124
rect 23014 10072 23020 10124
rect 23072 10072 23078 10124
rect 23109 10115 23167 10121
rect 23109 10081 23121 10115
rect 23155 10081 23167 10115
rect 23109 10075 23167 10081
rect 23201 10115 23259 10121
rect 23201 10081 23213 10115
rect 23247 10112 23259 10115
rect 23382 10112 23388 10124
rect 23247 10084 23388 10112
rect 23247 10081 23259 10084
rect 23201 10075 23259 10081
rect 23124 10044 23152 10075
rect 23382 10072 23388 10084
rect 23440 10112 23446 10124
rect 23440 10084 23888 10112
rect 23440 10072 23446 10084
rect 22480 10016 23152 10044
rect 18601 9979 18659 9985
rect 18601 9945 18613 9979
rect 18647 9945 18659 9979
rect 23124 9976 23152 10016
rect 23477 10047 23535 10053
rect 23477 10013 23489 10047
rect 23523 10044 23535 10047
rect 23569 10047 23627 10053
rect 23569 10044 23581 10047
rect 23523 10016 23581 10044
rect 23523 10013 23535 10016
rect 23477 10007 23535 10013
rect 23569 10013 23581 10016
rect 23615 10013 23627 10047
rect 23860 10044 23888 10084
rect 24302 10072 24308 10124
rect 24360 10072 24366 10124
rect 24486 10072 24492 10124
rect 24544 10072 24550 10124
rect 24578 10072 24584 10124
rect 24636 10072 24642 10124
rect 24688 10121 24716 10152
rect 24854 10140 24860 10152
rect 24912 10140 24918 10192
rect 24673 10115 24731 10121
rect 24673 10081 24685 10115
rect 24719 10081 24731 10115
rect 24964 10112 24992 10220
rect 25976 10220 26148 10248
rect 25130 10140 25136 10192
rect 25188 10180 25194 10192
rect 25976 10189 26004 10220
rect 26142 10208 26148 10220
rect 26200 10208 26206 10260
rect 26418 10208 26424 10260
rect 26476 10208 26482 10260
rect 25777 10183 25835 10189
rect 25777 10180 25789 10183
rect 25188 10152 25789 10180
rect 25188 10140 25194 10152
rect 25777 10149 25789 10152
rect 25823 10149 25835 10183
rect 25777 10143 25835 10149
rect 25961 10183 26019 10189
rect 25961 10149 25973 10183
rect 26007 10149 26019 10183
rect 25961 10143 26019 10149
rect 26145 10115 26203 10121
rect 26145 10112 26157 10115
rect 24964 10084 26157 10112
rect 24673 10075 24731 10081
rect 26145 10081 26157 10084
rect 26191 10081 26203 10115
rect 26145 10075 26203 10081
rect 26970 10072 26976 10124
rect 27028 10072 27034 10124
rect 25041 10047 25099 10053
rect 25041 10044 25053 10047
rect 23860 10016 25053 10044
rect 23569 10007 23627 10013
rect 25041 10013 25053 10016
rect 25087 10013 25099 10047
rect 25041 10007 25099 10013
rect 25130 10004 25136 10056
rect 25188 10044 25194 10056
rect 25593 10047 25651 10053
rect 25593 10044 25605 10047
rect 25188 10016 25605 10044
rect 25188 10004 25194 10016
rect 25593 10013 25605 10016
rect 25639 10013 25651 10047
rect 25593 10007 25651 10013
rect 23842 9976 23848 9988
rect 23124 9948 23848 9976
rect 18601 9939 18659 9945
rect 23842 9936 23848 9948
rect 23900 9976 23906 9988
rect 24578 9976 24584 9988
rect 23900 9948 24584 9976
rect 23900 9936 23906 9948
rect 24578 9936 24584 9948
rect 24636 9936 24642 9988
rect 24949 9979 25007 9985
rect 24949 9945 24961 9979
rect 24995 9976 25007 9979
rect 26050 9976 26056 9988
rect 24995 9948 26056 9976
rect 24995 9945 25007 9948
rect 24949 9939 25007 9945
rect 26050 9936 26056 9948
rect 26108 9936 26114 9988
rect 17092 9880 17816 9908
rect 18785 9911 18843 9917
rect 17092 9868 17098 9880
rect 18785 9877 18797 9911
rect 18831 9908 18843 9911
rect 19429 9911 19487 9917
rect 19429 9908 19441 9911
rect 18831 9880 19441 9908
rect 18831 9877 18843 9880
rect 18785 9871 18843 9877
rect 19429 9877 19441 9880
rect 19475 9877 19487 9911
rect 19429 9871 19487 9877
rect 22094 9868 22100 9920
rect 22152 9868 22158 9920
rect 23750 9868 23756 9920
rect 23808 9908 23814 9920
rect 24213 9911 24271 9917
rect 24213 9908 24225 9911
rect 23808 9880 24225 9908
rect 23808 9868 23814 9880
rect 24213 9877 24225 9880
rect 24259 9877 24271 9911
rect 24213 9871 24271 9877
rect 552 9818 27416 9840
rect 552 9766 3756 9818
rect 3808 9766 3820 9818
rect 3872 9766 3884 9818
rect 3936 9766 3948 9818
rect 4000 9766 4012 9818
rect 4064 9766 10472 9818
rect 10524 9766 10536 9818
rect 10588 9766 10600 9818
rect 10652 9766 10664 9818
rect 10716 9766 10728 9818
rect 10780 9766 17188 9818
rect 17240 9766 17252 9818
rect 17304 9766 17316 9818
rect 17368 9766 17380 9818
rect 17432 9766 17444 9818
rect 17496 9766 23904 9818
rect 23956 9766 23968 9818
rect 24020 9766 24032 9818
rect 24084 9766 24096 9818
rect 24148 9766 24160 9818
rect 24212 9766 27416 9818
rect 552 9744 27416 9766
rect 3237 9707 3295 9713
rect 3237 9673 3249 9707
rect 3283 9704 3295 9707
rect 3326 9704 3332 9716
rect 3283 9676 3332 9704
rect 3283 9673 3295 9676
rect 3237 9667 3295 9673
rect 3326 9664 3332 9676
rect 3384 9664 3390 9716
rect 4890 9664 4896 9716
rect 4948 9664 4954 9716
rect 7558 9664 7564 9716
rect 7616 9704 7622 9716
rect 7653 9707 7711 9713
rect 7653 9704 7665 9707
rect 7616 9676 7665 9704
rect 7616 9664 7622 9676
rect 7653 9673 7665 9676
rect 7699 9673 7711 9707
rect 7653 9667 7711 9673
rect 12434 9664 12440 9716
rect 12492 9704 12498 9716
rect 13170 9704 13176 9716
rect 12492 9676 13176 9704
rect 12492 9664 12498 9676
rect 13170 9664 13176 9676
rect 13228 9664 13234 9716
rect 14642 9704 14648 9716
rect 13556 9676 14648 9704
rect 2958 9596 2964 9648
rect 3016 9596 3022 9648
rect 7742 9596 7748 9648
rect 7800 9636 7806 9648
rect 12066 9636 12072 9648
rect 7800 9608 12072 9636
rect 7800 9596 7806 9608
rect 12066 9596 12072 9608
rect 12124 9596 12130 9648
rect 12158 9596 12164 9648
rect 12216 9636 12222 9648
rect 13556 9636 13584 9676
rect 14642 9664 14648 9676
rect 14700 9664 14706 9716
rect 15194 9664 15200 9716
rect 15252 9664 15258 9716
rect 15378 9664 15384 9716
rect 15436 9704 15442 9716
rect 18230 9704 18236 9716
rect 15436 9676 18236 9704
rect 15436 9664 15442 9676
rect 18230 9664 18236 9676
rect 18288 9664 18294 9716
rect 22278 9664 22284 9716
rect 22336 9704 22342 9716
rect 22465 9707 22523 9713
rect 22465 9704 22477 9707
rect 22336 9676 22477 9704
rect 22336 9664 22342 9676
rect 22465 9673 22477 9676
rect 22511 9673 22523 9707
rect 22465 9667 22523 9673
rect 23658 9664 23664 9716
rect 23716 9664 23722 9716
rect 25130 9704 25136 9716
rect 24780 9676 25136 9704
rect 12216 9608 13584 9636
rect 14921 9639 14979 9645
rect 12216 9596 12222 9608
rect 14921 9605 14933 9639
rect 14967 9636 14979 9639
rect 15654 9636 15660 9648
rect 14967 9608 15660 9636
rect 14967 9605 14979 9608
rect 14921 9599 14979 9605
rect 15654 9596 15660 9608
rect 15712 9636 15718 9648
rect 15712 9608 16528 9636
rect 15712 9596 15718 9608
rect 2593 9571 2651 9577
rect 2593 9537 2605 9571
rect 2639 9568 2651 9571
rect 2682 9568 2688 9580
rect 2639 9540 2688 9568
rect 2639 9537 2651 9540
rect 2593 9531 2651 9537
rect 2682 9528 2688 9540
rect 2740 9528 2746 9580
rect 3053 9571 3111 9577
rect 3053 9537 3065 9571
rect 3099 9537 3111 9571
rect 3053 9531 3111 9537
rect 7285 9571 7343 9577
rect 7285 9537 7297 9571
rect 7331 9568 7343 9571
rect 9398 9568 9404 9580
rect 7331 9540 9404 9568
rect 7331 9537 7343 9540
rect 7285 9531 7343 9537
rect 2133 9503 2191 9509
rect 2133 9469 2145 9503
rect 2179 9500 2191 9503
rect 2314 9500 2320 9512
rect 2179 9472 2320 9500
rect 2179 9469 2191 9472
rect 2133 9463 2191 9469
rect 2314 9460 2320 9472
rect 2372 9460 2378 9512
rect 2498 9460 2504 9512
rect 2556 9500 2562 9512
rect 2866 9500 2872 9512
rect 2556 9472 2872 9500
rect 2556 9460 2562 9472
rect 2866 9460 2872 9472
rect 2924 9460 2930 9512
rect 3068 9500 3096 9531
rect 9398 9528 9404 9540
rect 9456 9528 9462 9580
rect 9508 9540 9720 9568
rect 3421 9503 3479 9509
rect 3421 9500 3433 9503
rect 3068 9472 3433 9500
rect 3421 9469 3433 9472
rect 3467 9469 3479 9503
rect 3421 9463 3479 9469
rect 3602 9460 3608 9512
rect 3660 9500 3666 9512
rect 3973 9503 4031 9509
rect 3973 9500 3985 9503
rect 3660 9472 3985 9500
rect 3660 9460 3666 9472
rect 3973 9469 3985 9472
rect 4019 9469 4031 9503
rect 3973 9463 4031 9469
rect 4157 9503 4215 9509
rect 4157 9469 4169 9503
rect 4203 9500 4215 9503
rect 4249 9503 4307 9509
rect 4249 9500 4261 9503
rect 4203 9472 4261 9500
rect 4203 9469 4215 9472
rect 4157 9463 4215 9469
rect 4249 9469 4261 9472
rect 4295 9469 4307 9503
rect 4249 9463 4307 9469
rect 4617 9503 4675 9509
rect 4617 9469 4629 9503
rect 4663 9500 4675 9503
rect 4798 9500 4804 9512
rect 4663 9472 4804 9500
rect 4663 9469 4675 9472
rect 4617 9463 4675 9469
rect 4798 9460 4804 9472
rect 4856 9460 4862 9512
rect 5074 9460 5080 9512
rect 5132 9460 5138 9512
rect 7834 9460 7840 9512
rect 7892 9460 7898 9512
rect 7929 9503 7987 9509
rect 7929 9469 7941 9503
rect 7975 9500 7987 9503
rect 8113 9503 8171 9509
rect 7975 9472 8064 9500
rect 7975 9469 7987 9472
rect 7929 9463 7987 9469
rect 1946 9392 1952 9444
rect 2004 9392 2010 9444
rect 2774 9392 2780 9444
rect 2832 9432 2838 9444
rect 4065 9435 4123 9441
rect 4065 9432 4077 9435
rect 2832 9404 4077 9432
rect 2832 9392 2838 9404
rect 4065 9401 4077 9404
rect 4111 9401 4123 9435
rect 4065 9395 4123 9401
rect 4433 9435 4491 9441
rect 4433 9401 4445 9435
rect 4479 9401 4491 9435
rect 4433 9395 4491 9401
rect 2317 9367 2375 9373
rect 2317 9333 2329 9367
rect 2363 9364 2375 9367
rect 2958 9364 2964 9376
rect 2363 9336 2964 9364
rect 2363 9333 2375 9336
rect 2317 9327 2375 9333
rect 2958 9324 2964 9336
rect 3016 9324 3022 9376
rect 3418 9324 3424 9376
rect 3476 9364 3482 9376
rect 4448 9364 4476 9395
rect 6914 9392 6920 9444
rect 6972 9432 6978 9444
rect 7018 9435 7076 9441
rect 7018 9432 7030 9435
rect 6972 9404 7030 9432
rect 6972 9392 6978 9404
rect 7018 9401 7030 9404
rect 7064 9401 7076 9435
rect 7018 9395 7076 9401
rect 3476 9336 4476 9364
rect 5905 9367 5963 9373
rect 3476 9324 3482 9336
rect 5905 9333 5917 9367
rect 5951 9364 5963 9367
rect 7466 9364 7472 9376
rect 5951 9336 7472 9364
rect 5951 9333 5963 9336
rect 5905 9327 5963 9333
rect 7466 9324 7472 9336
rect 7524 9324 7530 9376
rect 8036 9364 8064 9472
rect 8113 9469 8125 9503
rect 8159 9469 8171 9503
rect 8113 9463 8171 9469
rect 8205 9503 8263 9509
rect 8205 9469 8217 9503
rect 8251 9500 8263 9503
rect 8754 9500 8760 9512
rect 8251 9472 8760 9500
rect 8251 9469 8263 9472
rect 8205 9463 8263 9469
rect 8128 9432 8156 9463
rect 8754 9460 8760 9472
rect 8812 9460 8818 9512
rect 9033 9503 9091 9509
rect 9033 9469 9045 9503
rect 9079 9469 9091 9503
rect 9033 9463 9091 9469
rect 9048 9432 9076 9463
rect 9122 9460 9128 9512
rect 9180 9500 9186 9512
rect 9217 9503 9275 9509
rect 9217 9500 9229 9503
rect 9180 9472 9229 9500
rect 9180 9460 9186 9472
rect 9217 9469 9229 9472
rect 9263 9500 9275 9503
rect 9508 9500 9536 9540
rect 9263 9472 9536 9500
rect 9263 9469 9275 9472
rect 9217 9463 9275 9469
rect 9582 9460 9588 9512
rect 9640 9460 9646 9512
rect 9692 9509 9720 9540
rect 11054 9528 11060 9580
rect 11112 9568 11118 9580
rect 12342 9568 12348 9580
rect 11112 9540 12348 9568
rect 11112 9528 11118 9540
rect 9677 9503 9735 9509
rect 9677 9469 9689 9503
rect 9723 9469 9735 9503
rect 9677 9463 9735 9469
rect 9861 9503 9919 9509
rect 9861 9469 9873 9503
rect 9907 9500 9919 9503
rect 10318 9500 10324 9512
rect 9907 9472 10324 9500
rect 9907 9469 9919 9472
rect 9861 9463 9919 9469
rect 10318 9460 10324 9472
rect 10376 9460 10382 9512
rect 9769 9435 9827 9441
rect 9769 9432 9781 9435
rect 8128 9404 9781 9432
rect 9769 9401 9781 9404
rect 9815 9401 9827 9435
rect 9769 9395 9827 9401
rect 8662 9364 8668 9376
rect 8036 9336 8668 9364
rect 8662 9324 8668 9336
rect 8720 9324 8726 9376
rect 8849 9367 8907 9373
rect 8849 9333 8861 9367
rect 8895 9364 8907 9367
rect 8938 9364 8944 9376
rect 8895 9336 8944 9364
rect 8895 9333 8907 9336
rect 8849 9327 8907 9333
rect 8938 9324 8944 9336
rect 8996 9324 9002 9376
rect 11330 9324 11336 9376
rect 11388 9324 11394 9376
rect 11440 9364 11468 9540
rect 12342 9528 12348 9540
rect 12400 9528 12406 9580
rect 13078 9568 13084 9580
rect 12544 9540 13084 9568
rect 11517 9503 11575 9509
rect 11517 9469 11529 9503
rect 11563 9500 11575 9503
rect 11698 9500 11704 9512
rect 11563 9472 11704 9500
rect 11563 9469 11575 9472
rect 11517 9463 11575 9469
rect 11698 9460 11704 9472
rect 11756 9460 11762 9512
rect 11793 9503 11851 9509
rect 11793 9469 11805 9503
rect 11839 9500 11851 9503
rect 11974 9500 11980 9512
rect 11839 9472 11980 9500
rect 11839 9469 11851 9472
rect 11793 9463 11851 9469
rect 11974 9460 11980 9472
rect 12032 9460 12038 9512
rect 12158 9460 12164 9512
rect 12216 9460 12222 9512
rect 12253 9503 12311 9509
rect 12253 9469 12265 9503
rect 12299 9469 12311 9503
rect 12253 9463 12311 9469
rect 12268 9432 12296 9463
rect 12434 9460 12440 9512
rect 12492 9460 12498 9512
rect 12544 9509 12572 9540
rect 13078 9528 13084 9540
rect 13136 9528 13142 9580
rect 15562 9528 15568 9580
rect 15620 9568 15626 9580
rect 15620 9540 15884 9568
rect 15620 9528 15626 9540
rect 12529 9503 12587 9509
rect 12529 9469 12541 9503
rect 12575 9469 12587 9503
rect 12529 9463 12587 9469
rect 12894 9460 12900 9512
rect 12952 9460 12958 9512
rect 12986 9460 12992 9512
rect 13044 9460 13050 9512
rect 13170 9460 13176 9512
rect 13228 9460 13234 9512
rect 13262 9460 13268 9512
rect 13320 9460 13326 9512
rect 13541 9503 13599 9509
rect 13541 9469 13553 9503
rect 13587 9500 13599 9503
rect 13630 9500 13636 9512
rect 13587 9472 13636 9500
rect 13587 9469 13599 9472
rect 13541 9463 13599 9469
rect 13630 9460 13636 9472
rect 13688 9460 13694 9512
rect 15856 9509 15884 9540
rect 16298 9528 16304 9580
rect 16356 9528 16362 9580
rect 15749 9503 15807 9509
rect 15749 9500 15761 9503
rect 13740 9472 15761 9500
rect 12912 9432 12940 9460
rect 13740 9432 13768 9472
rect 15749 9469 15761 9472
rect 15795 9469 15807 9503
rect 15749 9463 15807 9469
rect 15841 9503 15899 9509
rect 15841 9469 15853 9503
rect 15887 9469 15899 9503
rect 15841 9463 15899 9469
rect 15930 9460 15936 9512
rect 15988 9500 15994 9512
rect 16025 9503 16083 9509
rect 16025 9500 16037 9503
rect 15988 9472 16037 9500
rect 15988 9460 15994 9472
rect 16025 9469 16037 9472
rect 16071 9469 16083 9503
rect 16025 9463 16083 9469
rect 16117 9503 16175 9509
rect 16117 9469 16129 9503
rect 16163 9469 16175 9503
rect 16117 9463 16175 9469
rect 16209 9503 16267 9509
rect 16209 9469 16221 9503
rect 16255 9500 16267 9503
rect 16316 9500 16344 9528
rect 16255 9472 16344 9500
rect 16255 9469 16267 9472
rect 16209 9463 16267 9469
rect 12268 9404 12848 9432
rect 12912 9404 13768 9432
rect 13808 9435 13866 9441
rect 12820 9376 12848 9404
rect 13808 9401 13820 9435
rect 13854 9401 13866 9435
rect 13808 9395 13866 9401
rect 11701 9367 11759 9373
rect 11701 9364 11713 9367
rect 11440 9336 11713 9364
rect 11701 9333 11713 9336
rect 11747 9333 11759 9367
rect 11701 9327 11759 9333
rect 11974 9324 11980 9376
rect 12032 9324 12038 9376
rect 12710 9324 12716 9376
rect 12768 9324 12774 9376
rect 12802 9324 12808 9376
rect 12860 9364 12866 9376
rect 12986 9364 12992 9376
rect 12860 9336 12992 9364
rect 12860 9324 12866 9336
rect 12986 9324 12992 9336
rect 13044 9324 13050 9376
rect 13538 9324 13544 9376
rect 13596 9364 13602 9376
rect 13823 9364 13851 9395
rect 14366 9392 14372 9444
rect 14424 9432 14430 9444
rect 15165 9435 15223 9441
rect 15165 9432 15177 9435
rect 14424 9404 15177 9432
rect 14424 9392 14430 9404
rect 15165 9401 15177 9404
rect 15211 9401 15223 9435
rect 15165 9395 15223 9401
rect 15378 9392 15384 9444
rect 15436 9392 15442 9444
rect 16132 9432 16160 9463
rect 16390 9460 16396 9512
rect 16448 9460 16454 9512
rect 16500 9509 16528 9608
rect 22370 9596 22376 9648
rect 22428 9636 22434 9648
rect 24780 9636 24808 9676
rect 25130 9664 25136 9676
rect 25188 9664 25194 9716
rect 25498 9664 25504 9716
rect 25556 9664 25562 9716
rect 22428 9608 23060 9636
rect 22428 9596 22434 9608
rect 23032 9577 23060 9608
rect 23400 9608 24808 9636
rect 23017 9571 23075 9577
rect 23017 9537 23029 9571
rect 23063 9537 23075 9571
rect 23017 9531 23075 9537
rect 16485 9503 16543 9509
rect 16485 9469 16497 9503
rect 16531 9469 16543 9503
rect 16485 9463 16543 9469
rect 16669 9503 16727 9509
rect 16669 9469 16681 9503
rect 16715 9469 16727 9503
rect 16669 9463 16727 9469
rect 16301 9435 16359 9441
rect 16301 9432 16313 9435
rect 16132 9404 16313 9432
rect 16301 9401 16313 9404
rect 16347 9401 16359 9435
rect 16408 9432 16436 9460
rect 16684 9432 16712 9463
rect 18690 9460 18696 9512
rect 18748 9460 18754 9512
rect 18877 9503 18935 9509
rect 18877 9469 18889 9503
rect 18923 9500 18935 9503
rect 19518 9500 19524 9512
rect 18923 9472 19524 9500
rect 18923 9469 18935 9472
rect 18877 9463 18935 9469
rect 19518 9460 19524 9472
rect 19576 9460 19582 9512
rect 20533 9503 20591 9509
rect 20533 9469 20545 9503
rect 20579 9500 20591 9503
rect 20990 9500 20996 9512
rect 20579 9472 20996 9500
rect 20579 9469 20591 9472
rect 20533 9463 20591 9469
rect 20990 9460 20996 9472
rect 21048 9460 21054 9512
rect 21260 9503 21318 9509
rect 21260 9469 21272 9503
rect 21306 9500 21318 9503
rect 22094 9500 22100 9512
rect 21306 9472 22100 9500
rect 21306 9469 21318 9472
rect 21260 9463 21318 9469
rect 22094 9460 22100 9472
rect 22152 9460 22158 9512
rect 22646 9460 22652 9512
rect 22704 9500 22710 9512
rect 23400 9509 23428 9608
rect 27062 9596 27068 9648
rect 27120 9596 27126 9648
rect 23566 9528 23572 9580
rect 23624 9528 23630 9580
rect 24118 9528 24124 9580
rect 24176 9568 24182 9580
rect 24302 9568 24308 9580
rect 24176 9540 24308 9568
rect 24176 9528 24182 9540
rect 24302 9528 24308 9540
rect 24360 9568 24366 9580
rect 24360 9540 25820 9568
rect 24360 9528 24366 9540
rect 23385 9503 23443 9509
rect 23385 9500 23397 9503
rect 22704 9472 23397 9500
rect 22704 9460 22710 9472
rect 23385 9469 23397 9472
rect 23431 9469 23443 9503
rect 23845 9503 23903 9509
rect 23845 9500 23857 9503
rect 23385 9463 23443 9469
rect 23584 9472 23857 9500
rect 16408 9404 16712 9432
rect 16301 9395 16359 9401
rect 16942 9392 16948 9444
rect 17000 9432 17006 9444
rect 17000 9404 19748 9432
rect 17000 9392 17006 9404
rect 13596 9336 13851 9364
rect 13596 9324 13602 9336
rect 15010 9324 15016 9376
rect 15068 9324 15074 9376
rect 15565 9367 15623 9373
rect 15565 9333 15577 9367
rect 15611 9364 15623 9367
rect 15746 9364 15752 9376
rect 15611 9336 15752 9364
rect 15611 9333 15623 9336
rect 15565 9327 15623 9333
rect 15746 9324 15752 9336
rect 15804 9324 15810 9376
rect 15930 9324 15936 9376
rect 15988 9364 15994 9376
rect 16577 9367 16635 9373
rect 16577 9364 16589 9367
rect 15988 9336 16589 9364
rect 15988 9324 15994 9336
rect 16577 9333 16589 9336
rect 16623 9333 16635 9367
rect 16577 9327 16635 9333
rect 18782 9324 18788 9376
rect 18840 9324 18846 9376
rect 19153 9367 19211 9373
rect 19153 9333 19165 9367
rect 19199 9364 19211 9367
rect 19610 9364 19616 9376
rect 19199 9336 19616 9364
rect 19199 9333 19211 9336
rect 19153 9327 19211 9333
rect 19610 9324 19616 9336
rect 19668 9324 19674 9376
rect 19720 9364 19748 9404
rect 19978 9392 19984 9444
rect 20036 9432 20042 9444
rect 20266 9435 20324 9441
rect 20266 9432 20278 9435
rect 20036 9404 20278 9432
rect 20036 9392 20042 9404
rect 20266 9401 20278 9404
rect 20312 9401 20324 9435
rect 20266 9395 20324 9401
rect 21910 9392 21916 9444
rect 21968 9432 21974 9444
rect 23584 9432 23612 9472
rect 23845 9469 23857 9472
rect 23891 9469 23903 9503
rect 23845 9463 23903 9469
rect 24581 9503 24639 9509
rect 24581 9469 24593 9503
rect 24627 9500 24639 9503
rect 24670 9500 24676 9512
rect 24627 9472 24676 9500
rect 24627 9469 24639 9472
rect 24581 9463 24639 9469
rect 24670 9460 24676 9472
rect 24728 9460 24734 9512
rect 24872 9509 24900 9540
rect 24857 9503 24915 9509
rect 24857 9469 24869 9503
rect 24903 9469 24915 9503
rect 24857 9463 24915 9469
rect 25038 9460 25044 9512
rect 25096 9460 25102 9512
rect 25130 9460 25136 9512
rect 25188 9460 25194 9512
rect 25222 9460 25228 9512
rect 25280 9460 25286 9512
rect 25590 9460 25596 9512
rect 25648 9500 25654 9512
rect 25685 9503 25743 9509
rect 25685 9500 25697 9503
rect 25648 9472 25697 9500
rect 25648 9460 25654 9472
rect 25685 9469 25697 9472
rect 25731 9469 25743 9503
rect 25792 9500 25820 9540
rect 26234 9500 26240 9512
rect 25792 9472 26240 9500
rect 25685 9463 25743 9469
rect 26234 9460 26240 9472
rect 26292 9460 26298 9512
rect 21968 9404 23612 9432
rect 23661 9435 23719 9441
rect 21968 9392 21974 9404
rect 23661 9401 23673 9435
rect 23707 9432 23719 9435
rect 24946 9432 24952 9444
rect 23707 9404 24952 9432
rect 23707 9401 23719 9404
rect 23661 9395 23719 9401
rect 24946 9392 24952 9404
rect 25004 9392 25010 9444
rect 25608 9432 25636 9460
rect 25056 9404 25636 9432
rect 21358 9364 21364 9376
rect 19720 9336 21364 9364
rect 21358 9324 21364 9336
rect 21416 9324 21422 9376
rect 22186 9324 22192 9376
rect 22244 9364 22250 9376
rect 23201 9367 23259 9373
rect 23201 9364 23213 9367
rect 22244 9336 23213 9364
rect 22244 9324 22250 9336
rect 23201 9333 23213 9336
rect 23247 9333 23259 9367
rect 23201 9327 23259 9333
rect 24670 9324 24676 9376
rect 24728 9364 24734 9376
rect 25056 9364 25084 9404
rect 25774 9392 25780 9444
rect 25832 9432 25838 9444
rect 25930 9435 25988 9441
rect 25930 9432 25942 9435
rect 25832 9404 25942 9432
rect 25832 9392 25838 9404
rect 25930 9401 25942 9404
rect 25976 9401 25988 9435
rect 25930 9395 25988 9401
rect 24728 9336 25084 9364
rect 24728 9324 24734 9336
rect 25130 9324 25136 9376
rect 25188 9364 25194 9376
rect 26050 9364 26056 9376
rect 25188 9336 26056 9364
rect 25188 9324 25194 9336
rect 26050 9324 26056 9336
rect 26108 9324 26114 9376
rect 552 9274 27576 9296
rect 552 9222 7114 9274
rect 7166 9222 7178 9274
rect 7230 9222 7242 9274
rect 7294 9222 7306 9274
rect 7358 9222 7370 9274
rect 7422 9222 13830 9274
rect 13882 9222 13894 9274
rect 13946 9222 13958 9274
rect 14010 9222 14022 9274
rect 14074 9222 14086 9274
rect 14138 9222 20546 9274
rect 20598 9222 20610 9274
rect 20662 9222 20674 9274
rect 20726 9222 20738 9274
rect 20790 9222 20802 9274
rect 20854 9222 27262 9274
rect 27314 9222 27326 9274
rect 27378 9222 27390 9274
rect 27442 9222 27454 9274
rect 27506 9222 27518 9274
rect 27570 9222 27576 9274
rect 552 9200 27576 9222
rect 1394 9160 1400 9172
rect 860 9132 1400 9160
rect 860 9033 888 9132
rect 1394 9120 1400 9132
rect 1452 9160 1458 9172
rect 4154 9160 4160 9172
rect 1452 9132 4160 9160
rect 1452 9120 1458 9132
rect 4154 9120 4160 9132
rect 4212 9120 4218 9172
rect 7653 9163 7711 9169
rect 7653 9129 7665 9163
rect 7699 9129 7711 9163
rect 12158 9160 12164 9172
rect 7653 9123 7711 9129
rect 8772 9132 12164 9160
rect 2682 9101 2688 9104
rect 2669 9095 2688 9101
rect 2669 9061 2681 9095
rect 2669 9055 2688 9061
rect 2682 9052 2688 9055
rect 2740 9052 2746 9104
rect 2866 9052 2872 9104
rect 2924 9052 2930 9104
rect 3513 9095 3571 9101
rect 3513 9092 3525 9095
rect 3252 9064 3525 9092
rect 1118 9033 1124 9036
rect 845 9027 903 9033
rect 845 8993 857 9027
rect 891 8993 903 9027
rect 845 8987 903 8993
rect 1112 8987 1124 9033
rect 1118 8984 1124 8987
rect 1176 8984 1182 9036
rect 2314 8984 2320 9036
rect 2372 9024 2378 9036
rect 2372 8996 3096 9024
rect 2372 8984 2378 8996
rect 1946 8916 1952 8968
rect 2004 8956 2010 8968
rect 2004 8928 2912 8956
rect 2004 8916 2010 8928
rect 2056 8820 2084 8928
rect 2130 8848 2136 8900
rect 2188 8888 2194 8900
rect 2774 8888 2780 8900
rect 2188 8860 2780 8888
rect 2188 8848 2194 8860
rect 2774 8848 2780 8860
rect 2832 8848 2838 8900
rect 2884 8888 2912 8928
rect 2958 8916 2964 8968
rect 3016 8916 3022 8968
rect 3068 8956 3096 8996
rect 3142 8984 3148 9036
rect 3200 9024 3206 9036
rect 3252 9024 3280 9064
rect 3513 9061 3525 9064
rect 3559 9061 3571 9095
rect 7668 9092 7696 9123
rect 8772 9092 8800 9132
rect 12158 9120 12164 9132
rect 12216 9120 12222 9172
rect 13538 9120 13544 9172
rect 13596 9160 13602 9172
rect 13909 9163 13967 9169
rect 13909 9160 13921 9163
rect 13596 9132 13921 9160
rect 13596 9120 13602 9132
rect 13909 9129 13921 9132
rect 13955 9129 13967 9163
rect 13909 9123 13967 9129
rect 14182 9120 14188 9172
rect 14240 9160 14246 9172
rect 19521 9163 19579 9169
rect 19521 9160 19533 9163
rect 14240 9132 19533 9160
rect 14240 9120 14246 9132
rect 19521 9129 19533 9132
rect 19567 9129 19579 9163
rect 19521 9123 19579 9129
rect 19978 9120 19984 9172
rect 20036 9120 20042 9172
rect 22646 9120 22652 9172
rect 22704 9120 22710 9172
rect 24578 9160 24584 9172
rect 24412 9132 24584 9160
rect 10870 9092 10876 9104
rect 7668 9064 8800 9092
rect 3513 9055 3571 9061
rect 3200 8996 3280 9024
rect 3421 9027 3479 9033
rect 3200 8984 3206 8996
rect 3421 8993 3433 9027
rect 3467 8993 3479 9027
rect 3421 8987 3479 8993
rect 3605 9027 3663 9033
rect 3605 8993 3617 9027
rect 3651 8993 3663 9027
rect 3605 8987 3663 8993
rect 7285 9027 7343 9033
rect 7285 8993 7297 9027
rect 7331 9024 7343 9027
rect 7466 9024 7472 9036
rect 7331 8996 7472 9024
rect 7331 8993 7343 8996
rect 7285 8987 7343 8993
rect 3436 8956 3464 8987
rect 3068 8928 3464 8956
rect 3620 8888 3648 8987
rect 7466 8984 7472 8996
rect 7524 9024 7530 9036
rect 8018 9024 8024 9036
rect 7524 8996 8024 9024
rect 7524 8984 7530 8996
rect 8018 8984 8024 8996
rect 8076 8984 8082 9036
rect 8772 9033 8800 9064
rect 10244 9064 10876 9092
rect 8757 9027 8815 9033
rect 8757 8993 8769 9027
rect 8803 8993 8815 9027
rect 8757 8987 8815 8993
rect 8849 9027 8907 9033
rect 8849 8993 8861 9027
rect 8895 8993 8907 9027
rect 8849 8987 8907 8993
rect 7006 8916 7012 8968
rect 7064 8956 7070 8968
rect 7193 8959 7251 8965
rect 7193 8956 7205 8959
rect 7064 8928 7205 8956
rect 7064 8916 7070 8928
rect 7193 8925 7205 8928
rect 7239 8925 7251 8959
rect 7193 8919 7251 8925
rect 8662 8916 8668 8968
rect 8720 8956 8726 8968
rect 8864 8956 8892 8987
rect 9030 8984 9036 9036
rect 9088 8984 9094 9036
rect 9125 9027 9183 9033
rect 9125 8993 9137 9027
rect 9171 9024 9183 9027
rect 9214 9024 9220 9036
rect 9171 8996 9220 9024
rect 9171 8993 9183 8996
rect 9125 8987 9183 8993
rect 9214 8984 9220 8996
rect 9272 8984 9278 9036
rect 10244 9033 10272 9064
rect 10870 9052 10876 9064
rect 10928 9052 10934 9104
rect 11232 9095 11290 9101
rect 11232 9061 11244 9095
rect 11278 9092 11290 9095
rect 11330 9092 11336 9104
rect 11278 9064 11336 9092
rect 11278 9061 11290 9064
rect 11232 9055 11290 9061
rect 11330 9052 11336 9064
rect 11388 9052 11394 9104
rect 15010 9092 15016 9104
rect 14108 9064 15016 9092
rect 10229 9027 10287 9033
rect 10229 8993 10241 9027
rect 10275 8993 10287 9027
rect 10229 8987 10287 8993
rect 10318 8984 10324 9036
rect 10376 9024 10382 9036
rect 10413 9027 10471 9033
rect 10413 9024 10425 9027
rect 10376 8996 10425 9024
rect 10376 8984 10382 8996
rect 10413 8993 10425 8996
rect 10459 8993 10471 9027
rect 10413 8987 10471 8993
rect 12713 9027 12771 9033
rect 12713 8993 12725 9027
rect 12759 8993 12771 9027
rect 12713 8987 12771 8993
rect 8720 8928 8892 8956
rect 8720 8916 8726 8928
rect 9306 8916 9312 8968
rect 9364 8956 9370 8968
rect 10965 8959 11023 8965
rect 10965 8956 10977 8959
rect 9364 8928 10977 8956
rect 9364 8916 9370 8928
rect 10965 8925 10977 8928
rect 11011 8925 11023 8959
rect 10965 8919 11023 8925
rect 2884 8860 3648 8888
rect 7834 8848 7840 8900
rect 7892 8888 7898 8900
rect 9582 8888 9588 8900
rect 7892 8860 9588 8888
rect 7892 8848 7898 8860
rect 9582 8848 9588 8860
rect 9640 8888 9646 8900
rect 12728 8888 12756 8987
rect 12802 8984 12808 9036
rect 12860 8984 12866 9036
rect 12989 9027 13047 9033
rect 12989 8993 13001 9027
rect 13035 8993 13047 9027
rect 12989 8987 13047 8993
rect 13004 8956 13032 8987
rect 13078 8984 13084 9036
rect 13136 8984 13142 9036
rect 14108 9033 14136 9064
rect 15010 9052 15016 9064
rect 15068 9052 15074 9104
rect 15378 9052 15384 9104
rect 15436 9092 15442 9104
rect 16298 9092 16304 9104
rect 15436 9064 16304 9092
rect 15436 9052 15442 9064
rect 16298 9052 16304 9064
rect 16356 9052 16362 9104
rect 18690 9052 18696 9104
rect 18748 9092 18754 9104
rect 18748 9064 19334 9092
rect 18748 9052 18754 9064
rect 14093 9027 14151 9033
rect 14093 8993 14105 9027
rect 14139 8993 14151 9027
rect 14093 8987 14151 8993
rect 14182 8984 14188 9036
rect 14240 9024 14246 9036
rect 14277 9027 14335 9033
rect 14277 9024 14289 9027
rect 14240 8996 14289 9024
rect 14240 8984 14246 8996
rect 14277 8993 14289 8996
rect 14323 8993 14335 9027
rect 14277 8987 14335 8993
rect 14366 8984 14372 9036
rect 14424 8984 14430 9036
rect 15565 9027 15623 9033
rect 15565 8993 15577 9027
rect 15611 8993 15623 9027
rect 15565 8987 15623 8993
rect 13170 8956 13176 8968
rect 13004 8928 13176 8956
rect 13170 8916 13176 8928
rect 13228 8916 13234 8968
rect 15580 8956 15608 8987
rect 15654 8984 15660 9036
rect 15712 8984 15718 9036
rect 15838 8984 15844 9036
rect 15896 8984 15902 9036
rect 15930 8984 15936 9036
rect 15988 8984 15994 9036
rect 17304 9027 17362 9033
rect 17304 8993 17316 9027
rect 17350 9024 17362 9027
rect 17586 9024 17592 9036
rect 17350 8996 17592 9024
rect 17350 8993 17362 8996
rect 17304 8987 17362 8993
rect 17586 8984 17592 8996
rect 17644 8984 17650 9036
rect 19306 9024 19334 9064
rect 19610 9052 19616 9104
rect 19668 9092 19674 9104
rect 19668 9064 20852 9092
rect 19668 9052 19674 9064
rect 19521 9027 19579 9033
rect 19521 9024 19533 9027
rect 19306 8996 19533 9024
rect 19521 8993 19533 8996
rect 19567 8993 19579 9027
rect 19521 8987 19579 8993
rect 20162 8984 20168 9036
rect 20220 8984 20226 9036
rect 20438 8984 20444 9036
rect 20496 8984 20502 9036
rect 20824 9033 20852 9064
rect 20990 9052 20996 9104
rect 21048 9092 21054 9104
rect 21266 9092 21272 9104
rect 21048 9064 21272 9092
rect 21048 9052 21054 9064
rect 21266 9052 21272 9064
rect 21324 9092 21330 9104
rect 22002 9092 22008 9104
rect 21324 9064 22008 9092
rect 21324 9052 21330 9064
rect 22002 9052 22008 9064
rect 22060 9092 22066 9104
rect 22060 9064 24072 9092
rect 22060 9052 22066 9064
rect 20809 9027 20867 9033
rect 20809 8993 20821 9027
rect 20855 8993 20867 9027
rect 20809 8987 20867 8993
rect 21358 8984 21364 9036
rect 21416 9024 21422 9036
rect 21729 9027 21787 9033
rect 21729 9024 21741 9027
rect 21416 8996 21741 9024
rect 21416 8984 21422 8996
rect 21729 8993 21741 8996
rect 21775 9024 21787 9027
rect 21818 9024 21824 9036
rect 21775 8996 21824 9024
rect 21775 8993 21787 8996
rect 21729 8987 21787 8993
rect 21818 8984 21824 8996
rect 21876 8984 21882 9036
rect 23750 8984 23756 9036
rect 23808 9033 23814 9036
rect 23808 9024 23820 9033
rect 23808 8996 23853 9024
rect 23808 8987 23820 8996
rect 23808 8984 23814 8987
rect 14476 8928 15608 8956
rect 9640 8860 10456 8888
rect 9640 8848 9646 8860
rect 2225 8823 2283 8829
rect 2225 8820 2237 8823
rect 2056 8792 2237 8820
rect 2225 8789 2237 8792
rect 2271 8789 2283 8823
rect 2225 8783 2283 8789
rect 2498 8780 2504 8832
rect 2556 8780 2562 8832
rect 2590 8780 2596 8832
rect 2648 8820 2654 8832
rect 2685 8823 2743 8829
rect 2685 8820 2697 8823
rect 2648 8792 2697 8820
rect 2648 8780 2654 8792
rect 2685 8789 2697 8792
rect 2731 8789 2743 8823
rect 2685 8783 2743 8789
rect 3050 8780 3056 8832
rect 3108 8820 3114 8832
rect 3329 8823 3387 8829
rect 3329 8820 3341 8823
rect 3108 8792 3341 8820
rect 3108 8780 3114 8792
rect 3329 8789 3341 8792
rect 3375 8789 3387 8823
rect 3329 8783 3387 8789
rect 8294 8780 8300 8832
rect 8352 8820 8358 8832
rect 8573 8823 8631 8829
rect 8573 8820 8585 8823
rect 8352 8792 8585 8820
rect 8352 8780 8358 8792
rect 8573 8789 8585 8792
rect 8619 8789 8631 8823
rect 8573 8783 8631 8789
rect 10226 8780 10232 8832
rect 10284 8820 10290 8832
rect 10321 8823 10379 8829
rect 10321 8820 10333 8823
rect 10284 8792 10333 8820
rect 10284 8780 10290 8792
rect 10321 8789 10333 8792
rect 10367 8789 10379 8823
rect 10428 8820 10456 8860
rect 11900 8860 12756 8888
rect 11900 8820 11928 8860
rect 10428 8792 11928 8820
rect 10321 8783 10379 8789
rect 12342 8780 12348 8832
rect 12400 8780 12406 8832
rect 12434 8780 12440 8832
rect 12492 8820 12498 8832
rect 12529 8823 12587 8829
rect 12529 8820 12541 8823
rect 12492 8792 12541 8820
rect 12492 8780 12498 8792
rect 12529 8789 12541 8792
rect 12575 8789 12587 8823
rect 12728 8820 12756 8860
rect 14476 8820 14504 8928
rect 15746 8916 15752 8968
rect 15804 8956 15810 8968
rect 16758 8956 16764 8968
rect 15804 8928 16764 8956
rect 15804 8916 15810 8928
rect 16758 8916 16764 8928
rect 16816 8916 16822 8968
rect 17034 8916 17040 8968
rect 17092 8916 17098 8968
rect 19058 8956 19064 8968
rect 18432 8928 19064 8956
rect 18432 8897 18460 8928
rect 19058 8916 19064 8928
rect 19116 8956 19122 8968
rect 19153 8959 19211 8965
rect 19153 8956 19165 8959
rect 19116 8928 19165 8956
rect 19116 8916 19122 8928
rect 19153 8925 19165 8928
rect 19199 8925 19211 8959
rect 19153 8919 19211 8925
rect 19242 8916 19248 8968
rect 19300 8956 19306 8968
rect 19337 8959 19395 8965
rect 19337 8956 19349 8959
rect 19300 8928 19349 8956
rect 19300 8916 19306 8928
rect 19337 8925 19349 8928
rect 19383 8925 19395 8959
rect 19337 8919 19395 8925
rect 19426 8916 19432 8968
rect 19484 8956 19490 8968
rect 19886 8956 19892 8968
rect 19484 8928 19892 8956
rect 19484 8916 19490 8928
rect 19886 8916 19892 8928
rect 19944 8916 19950 8968
rect 20070 8916 20076 8968
rect 20128 8956 20134 8968
rect 24044 8965 24072 9064
rect 24118 8984 24124 9036
rect 24176 8984 24182 9036
rect 24302 8984 24308 9036
rect 24360 8984 24366 9036
rect 24412 9033 24440 9132
rect 24578 9120 24584 9132
rect 24636 9160 24642 9172
rect 25130 9160 25136 9172
rect 24636 9132 25136 9160
rect 24636 9120 24642 9132
rect 25130 9120 25136 9132
rect 25188 9120 25194 9172
rect 25593 9163 25651 9169
rect 25593 9129 25605 9163
rect 25639 9160 25651 9163
rect 25774 9160 25780 9172
rect 25639 9132 25780 9160
rect 25639 9129 25651 9132
rect 25593 9123 25651 9129
rect 25774 9120 25780 9132
rect 25832 9120 25838 9172
rect 25958 9120 25964 9172
rect 26016 9120 26022 9172
rect 24854 9092 24860 9104
rect 24504 9064 24860 9092
rect 24504 9033 24532 9064
rect 24854 9052 24860 9064
rect 24912 9052 24918 9104
rect 25222 9052 25228 9104
rect 25280 9092 25286 9104
rect 25976 9092 26004 9120
rect 26421 9095 26479 9101
rect 26421 9092 26433 9095
rect 25280 9064 26433 9092
rect 25280 9052 25286 9064
rect 26421 9061 26433 9064
rect 26467 9061 26479 9095
rect 26421 9055 26479 9061
rect 24397 9027 24455 9033
rect 24397 8993 24409 9027
rect 24443 8993 24455 9027
rect 24397 8987 24455 8993
rect 24489 9027 24547 9033
rect 24489 8993 24501 9027
rect 24535 8993 24547 9027
rect 24489 8987 24547 8993
rect 25869 9027 25927 9033
rect 25869 8993 25881 9027
rect 25915 8993 25927 9027
rect 25869 8987 25927 8993
rect 25961 9027 26019 9033
rect 25961 8993 25973 9027
rect 26007 8993 26019 9027
rect 25961 8987 26019 8993
rect 26053 9027 26111 9033
rect 26053 8993 26065 9027
rect 26099 9024 26111 9027
rect 26142 9024 26148 9036
rect 26099 8996 26148 9024
rect 26099 8993 26111 8996
rect 26053 8987 26111 8993
rect 20257 8959 20315 8965
rect 20257 8956 20269 8959
rect 20128 8928 20269 8956
rect 20128 8916 20134 8928
rect 20257 8925 20269 8928
rect 20303 8956 20315 8959
rect 20625 8959 20683 8965
rect 20625 8956 20637 8959
rect 20303 8928 20637 8956
rect 20303 8925 20315 8928
rect 20257 8919 20315 8925
rect 20625 8925 20637 8928
rect 20671 8925 20683 8959
rect 20625 8919 20683 8925
rect 20993 8959 21051 8965
rect 20993 8925 21005 8959
rect 21039 8925 21051 8959
rect 20993 8919 21051 8925
rect 24029 8959 24087 8965
rect 24029 8925 24041 8959
rect 24075 8956 24087 8959
rect 24670 8956 24676 8968
rect 24075 8928 24676 8956
rect 24075 8925 24087 8928
rect 24029 8919 24087 8925
rect 18417 8891 18475 8897
rect 18417 8857 18429 8891
rect 18463 8857 18475 8891
rect 18417 8851 18475 8857
rect 20349 8891 20407 8897
rect 20349 8857 20361 8891
rect 20395 8888 20407 8891
rect 20806 8888 20812 8900
rect 20395 8860 20812 8888
rect 20395 8857 20407 8860
rect 20349 8851 20407 8857
rect 20806 8848 20812 8860
rect 20864 8848 20870 8900
rect 12728 8792 14504 8820
rect 15381 8823 15439 8829
rect 12529 8783 12587 8789
rect 15381 8789 15393 8823
rect 15427 8820 15439 8823
rect 16850 8820 16856 8832
rect 15427 8792 16856 8820
rect 15427 8789 15439 8792
rect 15381 8783 15439 8789
rect 16850 8780 16856 8792
rect 16908 8780 16914 8832
rect 18601 8823 18659 8829
rect 18601 8789 18613 8823
rect 18647 8820 18659 8823
rect 18874 8820 18880 8832
rect 18647 8792 18880 8820
rect 18647 8789 18659 8792
rect 18601 8783 18659 8789
rect 18874 8780 18880 8792
rect 18932 8780 18938 8832
rect 19886 8780 19892 8832
rect 19944 8820 19950 8832
rect 21008 8820 21036 8919
rect 24670 8916 24676 8928
rect 24728 8916 24734 8968
rect 24765 8959 24823 8965
rect 24765 8925 24777 8959
rect 24811 8956 24823 8959
rect 24857 8959 24915 8965
rect 24857 8956 24869 8959
rect 24811 8928 24869 8956
rect 24811 8925 24823 8928
rect 24765 8919 24823 8925
rect 24857 8925 24869 8928
rect 24903 8925 24915 8959
rect 25884 8956 25912 8987
rect 24857 8919 24915 8925
rect 25792 8928 25912 8956
rect 25976 8956 26004 8987
rect 26142 8984 26148 8996
rect 26200 8984 26206 9036
rect 26234 8984 26240 9036
rect 26292 8984 26298 9036
rect 26878 8984 26884 9036
rect 26936 9024 26942 9036
rect 26973 9027 27031 9033
rect 26973 9024 26985 9027
rect 26936 8996 26985 9024
rect 26936 8984 26942 8996
rect 26973 8993 26985 8996
rect 27019 8993 27031 9027
rect 26973 8987 27031 8993
rect 25976 8928 26096 8956
rect 19944 8792 21036 8820
rect 21913 8823 21971 8829
rect 19944 8780 19950 8792
rect 21913 8789 21925 8823
rect 21959 8820 21971 8823
rect 24118 8820 24124 8832
rect 21959 8792 24124 8820
rect 21959 8789 21971 8792
rect 21913 8783 21971 8789
rect 24118 8780 24124 8792
rect 24176 8780 24182 8832
rect 24946 8780 24952 8832
rect 25004 8820 25010 8832
rect 25501 8823 25559 8829
rect 25501 8820 25513 8823
rect 25004 8792 25513 8820
rect 25004 8780 25010 8792
rect 25501 8789 25513 8792
rect 25547 8789 25559 8823
rect 25792 8820 25820 8928
rect 26068 8900 26096 8928
rect 26050 8848 26056 8900
rect 26108 8848 26114 8900
rect 26418 8820 26424 8832
rect 25792 8792 26424 8820
rect 25501 8783 25559 8789
rect 26418 8780 26424 8792
rect 26476 8780 26482 8832
rect 552 8730 27416 8752
rect 552 8678 3756 8730
rect 3808 8678 3820 8730
rect 3872 8678 3884 8730
rect 3936 8678 3948 8730
rect 4000 8678 4012 8730
rect 4064 8678 10472 8730
rect 10524 8678 10536 8730
rect 10588 8678 10600 8730
rect 10652 8678 10664 8730
rect 10716 8678 10728 8730
rect 10780 8678 17188 8730
rect 17240 8678 17252 8730
rect 17304 8678 17316 8730
rect 17368 8678 17380 8730
rect 17432 8678 17444 8730
rect 17496 8678 23904 8730
rect 23956 8678 23968 8730
rect 24020 8678 24032 8730
rect 24084 8678 24096 8730
rect 24148 8678 24160 8730
rect 24212 8678 27416 8730
rect 552 8656 27416 8678
rect 1118 8576 1124 8628
rect 1176 8576 1182 8628
rect 2133 8619 2191 8625
rect 2133 8585 2145 8619
rect 2179 8616 2191 8619
rect 2590 8616 2596 8628
rect 2179 8588 2596 8616
rect 2179 8585 2191 8588
rect 2133 8579 2191 8585
rect 2590 8576 2596 8588
rect 2648 8576 2654 8628
rect 2774 8576 2780 8628
rect 2832 8576 2838 8628
rect 3234 8576 3240 8628
rect 3292 8616 3298 8628
rect 4801 8619 4859 8625
rect 3292 8588 4476 8616
rect 3292 8576 3298 8588
rect 2409 8551 2467 8557
rect 2409 8517 2421 8551
rect 2455 8548 2467 8551
rect 3050 8548 3056 8560
rect 2455 8520 3056 8548
rect 2455 8517 2467 8520
rect 2409 8511 2467 8517
rect 3050 8508 3056 8520
rect 3108 8508 3114 8560
rect 2498 8480 2504 8492
rect 1320 8452 2504 8480
rect 1320 8421 1348 8452
rect 2498 8440 2504 8452
rect 2556 8440 2562 8492
rect 4448 8480 4476 8588
rect 4801 8585 4813 8619
rect 4847 8616 4859 8619
rect 5074 8616 5080 8628
rect 4847 8588 5080 8616
rect 4847 8585 4859 8588
rect 4801 8579 4859 8585
rect 5074 8576 5080 8588
rect 5132 8576 5138 8628
rect 11146 8616 11152 8628
rect 10428 8588 11152 8616
rect 6273 8551 6331 8557
rect 6273 8517 6285 8551
rect 6319 8548 6331 8551
rect 6546 8548 6552 8560
rect 6319 8520 6552 8548
rect 6319 8517 6331 8520
rect 6273 8511 6331 8517
rect 6546 8508 6552 8520
rect 6604 8508 6610 8560
rect 8478 8508 8484 8560
rect 8536 8548 8542 8560
rect 10428 8548 10456 8588
rect 11146 8576 11152 8588
rect 11204 8576 11210 8628
rect 11698 8576 11704 8628
rect 11756 8576 11762 8628
rect 11885 8619 11943 8625
rect 11885 8585 11897 8619
rect 11931 8616 11943 8619
rect 12161 8619 12219 8625
rect 12161 8616 12173 8619
rect 11931 8588 12173 8616
rect 11931 8585 11943 8588
rect 11885 8579 11943 8585
rect 12161 8585 12173 8588
rect 12207 8585 12219 8619
rect 12161 8579 12219 8585
rect 12897 8619 12955 8625
rect 12897 8585 12909 8619
rect 12943 8616 12955 8619
rect 13078 8616 13084 8628
rect 12943 8588 13084 8616
rect 12943 8585 12955 8588
rect 12897 8579 12955 8585
rect 13078 8576 13084 8588
rect 13136 8576 13142 8628
rect 14182 8576 14188 8628
rect 14240 8576 14246 8628
rect 17497 8619 17555 8625
rect 15028 8588 17448 8616
rect 8536 8520 10456 8548
rect 8536 8508 8542 8520
rect 9140 8489 9168 8520
rect 10502 8508 10508 8560
rect 10560 8548 10566 8560
rect 13722 8548 13728 8560
rect 10560 8520 13728 8548
rect 10560 8508 10566 8520
rect 13722 8508 13728 8520
rect 13780 8508 13786 8560
rect 15028 8548 15056 8588
rect 13924 8520 15056 8548
rect 9125 8483 9183 8489
rect 4448 8452 5028 8480
rect 1305 8415 1363 8421
rect 1305 8381 1317 8415
rect 1351 8381 1363 8415
rect 1305 8375 1363 8381
rect 1949 8415 2007 8421
rect 1949 8381 1961 8415
rect 1995 8381 2007 8415
rect 1949 8375 2007 8381
rect 1964 8344 1992 8375
rect 2130 8372 2136 8424
rect 2188 8372 2194 8424
rect 2590 8412 2596 8424
rect 2240 8384 2596 8412
rect 2240 8344 2268 8384
rect 2590 8372 2596 8384
rect 2648 8412 2654 8424
rect 2777 8415 2835 8421
rect 2777 8412 2789 8415
rect 2648 8384 2789 8412
rect 2648 8372 2654 8384
rect 2777 8381 2789 8384
rect 2823 8381 2835 8415
rect 2777 8375 2835 8381
rect 3050 8372 3056 8424
rect 3108 8372 3114 8424
rect 3421 8415 3479 8421
rect 3421 8381 3433 8415
rect 3467 8412 3479 8415
rect 4154 8412 4160 8424
rect 3467 8384 4160 8412
rect 3467 8381 3479 8384
rect 3421 8375 3479 8381
rect 4154 8372 4160 8384
rect 4212 8412 4218 8424
rect 4890 8412 4896 8424
rect 4212 8384 4896 8412
rect 4212 8372 4218 8384
rect 4890 8372 4896 8384
rect 4948 8372 4954 8424
rect 5000 8412 5028 8452
rect 9125 8449 9137 8483
rect 9171 8449 9183 8483
rect 9125 8443 9183 8449
rect 9306 8440 9312 8492
rect 9364 8480 9370 8492
rect 11241 8483 11299 8489
rect 11241 8480 11253 8483
rect 9364 8452 11253 8480
rect 9364 8440 9370 8452
rect 11241 8449 11253 8452
rect 11287 8480 11299 8483
rect 13630 8480 13636 8492
rect 11287 8452 13636 8480
rect 11287 8449 11299 8452
rect 11241 8443 11299 8449
rect 13630 8440 13636 8452
rect 13688 8440 13694 8492
rect 5000 8384 5948 8412
rect 2682 8344 2688 8356
rect 1964 8316 2268 8344
rect 2516 8316 2688 8344
rect 2516 8285 2544 8316
rect 2682 8304 2688 8316
rect 2740 8304 2746 8356
rect 3688 8347 3746 8353
rect 3688 8313 3700 8347
rect 3734 8344 3746 8347
rect 4246 8344 4252 8356
rect 3734 8316 4252 8344
rect 3734 8313 3746 8316
rect 3688 8307 3746 8313
rect 4246 8304 4252 8316
rect 4304 8304 4310 8356
rect 5160 8347 5218 8353
rect 5160 8313 5172 8347
rect 5206 8344 5218 8347
rect 5810 8344 5816 8356
rect 5206 8316 5816 8344
rect 5206 8313 5218 8316
rect 5160 8307 5218 8313
rect 5810 8304 5816 8316
rect 5868 8304 5874 8356
rect 5920 8344 5948 8384
rect 6914 8372 6920 8424
rect 6972 8412 6978 8424
rect 7101 8415 7159 8421
rect 7101 8412 7113 8415
rect 6972 8384 7113 8412
rect 6972 8372 6978 8384
rect 7101 8381 7113 8384
rect 7147 8381 7159 8415
rect 7101 8375 7159 8381
rect 9493 8415 9551 8421
rect 9493 8381 9505 8415
rect 9539 8381 9551 8415
rect 9493 8375 9551 8381
rect 9217 8347 9275 8353
rect 9217 8344 9229 8347
rect 5920 8316 9229 8344
rect 9217 8313 9229 8316
rect 9263 8313 9275 8347
rect 9508 8344 9536 8375
rect 9582 8372 9588 8424
rect 9640 8412 9646 8424
rect 9677 8415 9735 8421
rect 9677 8412 9689 8415
rect 9640 8384 9689 8412
rect 9640 8372 9646 8384
rect 9677 8381 9689 8384
rect 9723 8381 9735 8415
rect 9677 8375 9735 8381
rect 9861 8415 9919 8421
rect 9861 8381 9873 8415
rect 9907 8412 9919 8415
rect 10594 8412 10600 8424
rect 9907 8384 10600 8412
rect 9907 8381 9919 8384
rect 9861 8375 9919 8381
rect 10594 8372 10600 8384
rect 10652 8372 10658 8424
rect 12250 8412 12256 8424
rect 11072 8384 12256 8412
rect 10226 8344 10232 8356
rect 9508 8316 10232 8344
rect 9217 8307 9275 8313
rect 10226 8304 10232 8316
rect 10284 8304 10290 8356
rect 10318 8304 10324 8356
rect 10376 8344 10382 8356
rect 10413 8347 10471 8353
rect 10413 8344 10425 8347
rect 10376 8316 10425 8344
rect 10376 8304 10382 8316
rect 10413 8313 10425 8316
rect 10459 8313 10471 8347
rect 10413 8307 10471 8313
rect 10502 8304 10508 8356
rect 10560 8304 10566 8356
rect 2501 8279 2559 8285
rect 2501 8245 2513 8279
rect 2547 8245 2559 8279
rect 2501 8239 2559 8245
rect 7006 8236 7012 8288
rect 7064 8276 7070 8288
rect 7285 8279 7343 8285
rect 7285 8276 7297 8279
rect 7064 8248 7297 8276
rect 7064 8236 7070 8248
rect 7285 8245 7297 8248
rect 7331 8245 7343 8279
rect 7285 8239 7343 8245
rect 8018 8236 8024 8288
rect 8076 8276 8082 8288
rect 11072 8276 11100 8384
rect 11146 8304 11152 8356
rect 11204 8344 11210 8356
rect 11882 8353 11888 8356
rect 11869 8347 11888 8353
rect 11204 8316 11836 8344
rect 11204 8304 11210 8316
rect 8076 8248 11100 8276
rect 11808 8276 11836 8316
rect 11869 8313 11881 8347
rect 11869 8307 11888 8313
rect 11882 8304 11888 8307
rect 11940 8304 11946 8356
rect 12084 8353 12112 8384
rect 12250 8372 12256 8384
rect 12308 8372 12314 8424
rect 12342 8372 12348 8424
rect 12400 8412 12406 8424
rect 12713 8415 12771 8421
rect 12713 8412 12725 8415
rect 12400 8384 12725 8412
rect 12400 8372 12406 8384
rect 12713 8381 12725 8384
rect 12759 8412 12771 8415
rect 12897 8415 12955 8421
rect 12897 8412 12909 8415
rect 12759 8384 12909 8412
rect 12759 8381 12771 8384
rect 12713 8375 12771 8381
rect 12897 8381 12909 8384
rect 12943 8381 12955 8415
rect 12897 8375 12955 8381
rect 12986 8372 12992 8424
rect 13044 8412 13050 8424
rect 13081 8415 13139 8421
rect 13081 8412 13093 8415
rect 13044 8384 13093 8412
rect 13044 8372 13050 8384
rect 13081 8381 13093 8384
rect 13127 8381 13139 8415
rect 13081 8375 13139 8381
rect 12069 8347 12127 8353
rect 12069 8313 12081 8347
rect 12115 8313 12127 8347
rect 13924 8344 13952 8520
rect 15102 8508 15108 8560
rect 15160 8548 15166 8560
rect 15473 8551 15531 8557
rect 15473 8548 15485 8551
rect 15160 8520 15485 8548
rect 15160 8508 15166 8520
rect 15473 8517 15485 8520
rect 15519 8517 15531 8551
rect 15473 8511 15531 8517
rect 14642 8480 14648 8492
rect 14108 8452 14648 8480
rect 12069 8307 12127 8313
rect 12176 8316 13952 8344
rect 14001 8347 14059 8353
rect 12176 8276 12204 8316
rect 14001 8313 14013 8347
rect 14047 8344 14059 8347
rect 14108 8344 14136 8452
rect 14642 8440 14648 8452
rect 14700 8480 14706 8492
rect 16942 8480 16948 8492
rect 14700 8452 16948 8480
rect 14700 8440 14706 8452
rect 16942 8440 16948 8452
rect 17000 8440 17006 8492
rect 14826 8372 14832 8424
rect 14884 8412 14890 8424
rect 14884 8384 15148 8412
rect 14884 8372 14890 8384
rect 14274 8353 14280 8356
rect 14047 8316 14136 8344
rect 14217 8347 14280 8353
rect 14047 8313 14059 8316
rect 14001 8307 14059 8313
rect 14217 8313 14229 8347
rect 14263 8313 14280 8347
rect 14217 8307 14280 8313
rect 14274 8304 14280 8307
rect 14332 8304 14338 8356
rect 15120 8353 15148 8384
rect 15286 8372 15292 8424
rect 15344 8372 15350 8424
rect 15378 8372 15384 8424
rect 15436 8414 15442 8424
rect 15436 8386 15479 8414
rect 15436 8372 15442 8386
rect 15562 8372 15568 8424
rect 15620 8372 15626 8424
rect 16482 8372 16488 8424
rect 16540 8372 16546 8424
rect 14921 8347 14979 8353
rect 14921 8313 14933 8347
rect 14967 8313 14979 8347
rect 14921 8307 14979 8313
rect 15105 8347 15163 8353
rect 15105 8313 15117 8347
rect 15151 8313 15163 8347
rect 17420 8344 17448 8588
rect 17497 8585 17509 8619
rect 17543 8616 17555 8619
rect 17586 8616 17592 8628
rect 17543 8588 17592 8616
rect 17543 8585 17555 8588
rect 17497 8579 17555 8585
rect 17586 8576 17592 8588
rect 17644 8576 17650 8628
rect 18690 8576 18696 8628
rect 18748 8616 18754 8628
rect 18785 8619 18843 8625
rect 18785 8616 18797 8619
rect 18748 8588 18797 8616
rect 18748 8576 18754 8588
rect 18785 8585 18797 8588
rect 18831 8585 18843 8619
rect 18785 8579 18843 8585
rect 19518 8576 19524 8628
rect 19576 8576 19582 8628
rect 20438 8576 20444 8628
rect 20496 8616 20502 8628
rect 20533 8619 20591 8625
rect 20533 8616 20545 8619
rect 20496 8588 20545 8616
rect 20496 8576 20502 8588
rect 20533 8585 20545 8588
rect 20579 8585 20591 8619
rect 20533 8579 20591 8585
rect 22554 8576 22560 8628
rect 22612 8616 22618 8628
rect 23201 8619 23259 8625
rect 23201 8616 23213 8619
rect 22612 8588 23213 8616
rect 22612 8576 22618 8588
rect 23201 8585 23213 8588
rect 23247 8585 23259 8619
rect 23201 8579 23259 8585
rect 17954 8508 17960 8560
rect 18012 8548 18018 8560
rect 18049 8551 18107 8557
rect 18049 8548 18061 8551
rect 18012 8520 18061 8548
rect 18012 8508 18018 8520
rect 18049 8517 18061 8520
rect 18095 8548 18107 8551
rect 19242 8548 19248 8560
rect 18095 8520 19248 8548
rect 18095 8517 18107 8520
rect 18049 8511 18107 8517
rect 19242 8508 19248 8520
rect 19300 8508 19306 8560
rect 17865 8483 17923 8489
rect 17865 8449 17877 8483
rect 17911 8449 17923 8483
rect 19426 8480 19432 8492
rect 17865 8443 17923 8449
rect 18248 8452 19432 8480
rect 17681 8415 17739 8421
rect 17681 8381 17693 8415
rect 17727 8412 17739 8415
rect 17880 8412 17908 8443
rect 17727 8384 17908 8412
rect 17727 8381 17739 8384
rect 17681 8375 17739 8381
rect 18248 8344 18276 8452
rect 19426 8440 19432 8452
rect 19484 8440 19490 8492
rect 19705 8483 19763 8489
rect 19705 8449 19717 8483
rect 19751 8480 19763 8483
rect 20162 8480 20168 8492
rect 19751 8452 20168 8480
rect 19751 8449 19763 8452
rect 19705 8443 19763 8449
rect 20162 8440 20168 8452
rect 20220 8480 20226 8492
rect 24026 8480 24032 8492
rect 20220 8452 20300 8480
rect 20220 8440 20226 8452
rect 18690 8372 18696 8424
rect 18748 8372 18754 8424
rect 18874 8372 18880 8424
rect 18932 8372 18938 8424
rect 19058 8372 19064 8424
rect 19116 8412 19122 8424
rect 19153 8415 19211 8421
rect 19153 8412 19165 8415
rect 19116 8384 19165 8412
rect 19116 8372 19122 8384
rect 19153 8381 19165 8384
rect 19199 8381 19211 8415
rect 19153 8375 19211 8381
rect 17420 8316 18276 8344
rect 15105 8307 15163 8313
rect 11808 8248 12204 8276
rect 8076 8236 8082 8248
rect 14366 8236 14372 8288
rect 14424 8236 14430 8288
rect 14734 8236 14740 8288
rect 14792 8276 14798 8288
rect 14936 8276 14964 8307
rect 18322 8304 18328 8356
rect 18380 8304 18386 8356
rect 18708 8344 18736 8372
rect 19337 8347 19395 8353
rect 19337 8344 19349 8347
rect 18708 8316 19349 8344
rect 19337 8313 19349 8316
rect 19383 8313 19395 8347
rect 19444 8344 19472 8440
rect 19610 8372 19616 8424
rect 19668 8372 19674 8424
rect 19797 8415 19855 8421
rect 19797 8381 19809 8415
rect 19843 8412 19855 8415
rect 19886 8412 19892 8424
rect 19843 8384 19892 8412
rect 19843 8381 19855 8384
rect 19797 8375 19855 8381
rect 19886 8372 19892 8384
rect 19944 8372 19950 8424
rect 20070 8372 20076 8424
rect 20128 8372 20134 8424
rect 20272 8421 20300 8452
rect 21468 8452 24032 8480
rect 20257 8415 20315 8421
rect 20257 8381 20269 8415
rect 20303 8381 20315 8415
rect 20257 8375 20315 8381
rect 20441 8415 20499 8421
rect 20441 8381 20453 8415
rect 20487 8412 20499 8415
rect 20717 8415 20775 8421
rect 20717 8412 20729 8415
rect 20487 8384 20729 8412
rect 20487 8381 20499 8384
rect 20441 8375 20499 8381
rect 20717 8381 20729 8384
rect 20763 8381 20775 8415
rect 20717 8375 20775 8381
rect 20806 8372 20812 8424
rect 20864 8372 20870 8424
rect 21468 8421 21496 8452
rect 24026 8440 24032 8452
rect 24084 8440 24090 8492
rect 21453 8415 21511 8421
rect 21453 8381 21465 8415
rect 21499 8381 21511 8415
rect 21453 8375 21511 8381
rect 21545 8415 21603 8421
rect 21545 8381 21557 8415
rect 21591 8412 21603 8415
rect 21634 8412 21640 8424
rect 21591 8384 21640 8412
rect 21591 8381 21603 8384
rect 21545 8375 21603 8381
rect 21634 8372 21640 8384
rect 21692 8372 21698 8424
rect 21726 8372 21732 8424
rect 21784 8372 21790 8424
rect 23382 8372 23388 8424
rect 23440 8372 23446 8424
rect 24394 8412 24400 8424
rect 23492 8384 24400 8412
rect 20533 8347 20591 8353
rect 20533 8344 20545 8347
rect 19444 8316 20545 8344
rect 19337 8307 19395 8313
rect 20533 8313 20545 8316
rect 20579 8313 20591 8347
rect 20533 8307 20591 8313
rect 21818 8304 21824 8356
rect 21876 8344 21882 8356
rect 23492 8344 23520 8384
rect 24394 8372 24400 8384
rect 24452 8372 24458 8424
rect 24946 8372 24952 8424
rect 25004 8421 25010 8424
rect 25004 8412 25016 8421
rect 25225 8415 25283 8421
rect 25004 8384 25049 8412
rect 25004 8375 25016 8384
rect 25225 8381 25237 8415
rect 25271 8412 25283 8415
rect 25590 8412 25596 8424
rect 25271 8384 25596 8412
rect 25271 8381 25283 8384
rect 25225 8375 25283 8381
rect 25004 8372 25010 8375
rect 21876 8316 23520 8344
rect 21876 8304 21882 8316
rect 23566 8304 23572 8356
rect 23624 8344 23630 8356
rect 24118 8344 24124 8356
rect 23624 8316 24124 8344
rect 23624 8304 23630 8316
rect 24118 8304 24124 8316
rect 24176 8304 24182 8356
rect 25038 8304 25044 8356
rect 25096 8344 25102 8356
rect 25240 8344 25268 8375
rect 25590 8372 25596 8384
rect 25648 8372 25654 8424
rect 25096 8316 25268 8344
rect 25096 8304 25102 8316
rect 25682 8304 25688 8356
rect 25740 8344 25746 8356
rect 25838 8347 25896 8353
rect 25838 8344 25850 8347
rect 25740 8316 25850 8344
rect 25740 8304 25746 8316
rect 25838 8313 25850 8316
rect 25884 8313 25896 8347
rect 25838 8307 25896 8313
rect 14792 8248 14964 8276
rect 16301 8279 16359 8285
rect 14792 8236 14798 8248
rect 16301 8245 16313 8279
rect 16347 8276 16359 8279
rect 16390 8276 16396 8288
rect 16347 8248 16396 8276
rect 16347 8245 16359 8248
rect 16301 8239 16359 8245
rect 16390 8236 16396 8248
rect 16448 8236 16454 8288
rect 21358 8236 21364 8288
rect 21416 8236 21422 8288
rect 21542 8236 21548 8288
rect 21600 8276 21606 8288
rect 21637 8279 21695 8285
rect 21637 8276 21649 8279
rect 21600 8248 21649 8276
rect 21600 8236 21606 8248
rect 21637 8245 21649 8248
rect 21683 8245 21695 8279
rect 21637 8239 21695 8245
rect 23474 8236 23480 8288
rect 23532 8276 23538 8288
rect 23845 8279 23903 8285
rect 23845 8276 23857 8279
rect 23532 8248 23857 8276
rect 23532 8236 23538 8248
rect 23845 8245 23857 8248
rect 23891 8276 23903 8279
rect 24762 8276 24768 8288
rect 23891 8248 24768 8276
rect 23891 8245 23903 8248
rect 23845 8239 23903 8245
rect 24762 8236 24768 8248
rect 24820 8236 24826 8288
rect 25314 8236 25320 8288
rect 25372 8276 25378 8288
rect 26878 8276 26884 8288
rect 25372 8248 26884 8276
rect 25372 8236 25378 8248
rect 26878 8236 26884 8248
rect 26936 8276 26942 8288
rect 26973 8279 27031 8285
rect 26973 8276 26985 8279
rect 26936 8248 26985 8276
rect 26936 8236 26942 8248
rect 26973 8245 26985 8248
rect 27019 8245 27031 8279
rect 26973 8239 27031 8245
rect 552 8186 27576 8208
rect 552 8134 7114 8186
rect 7166 8134 7178 8186
rect 7230 8134 7242 8186
rect 7294 8134 7306 8186
rect 7358 8134 7370 8186
rect 7422 8134 13830 8186
rect 13882 8134 13894 8186
rect 13946 8134 13958 8186
rect 14010 8134 14022 8186
rect 14074 8134 14086 8186
rect 14138 8134 20546 8186
rect 20598 8134 20610 8186
rect 20662 8134 20674 8186
rect 20726 8134 20738 8186
rect 20790 8134 20802 8186
rect 20854 8134 27262 8186
rect 27314 8134 27326 8186
rect 27378 8134 27390 8186
rect 27442 8134 27454 8186
rect 27506 8134 27518 8186
rect 27570 8134 27576 8186
rect 552 8112 27576 8134
rect 10502 8072 10508 8084
rect 4172 8044 10508 8072
rect 4172 8013 4200 8044
rect 10502 8032 10508 8044
rect 10560 8032 10566 8084
rect 10594 8032 10600 8084
rect 10652 8072 10658 8084
rect 10652 8044 11008 8072
rect 10652 8032 10658 8044
rect 4157 8007 4215 8013
rect 4157 7973 4169 8007
rect 4203 7973 4215 8007
rect 4890 8004 4896 8016
rect 4157 7967 4215 7973
rect 4264 7976 4896 8004
rect 2501 7939 2559 7945
rect 2501 7905 2513 7939
rect 2547 7905 2559 7939
rect 2501 7899 2559 7905
rect 2685 7939 2743 7945
rect 2685 7905 2697 7939
rect 2731 7936 2743 7939
rect 3142 7936 3148 7948
rect 2731 7908 3148 7936
rect 2731 7905 2743 7908
rect 2685 7899 2743 7905
rect 2516 7868 2544 7899
rect 3142 7896 3148 7908
rect 3200 7896 3206 7948
rect 3421 7939 3479 7945
rect 3421 7905 3433 7939
rect 3467 7936 3479 7939
rect 4264 7936 4292 7976
rect 4890 7964 4896 7976
rect 4948 8004 4954 8016
rect 4948 7976 6132 8004
rect 4948 7964 4954 7976
rect 3467 7908 4292 7936
rect 3467 7905 3479 7908
rect 3421 7899 3479 7905
rect 4430 7896 4436 7948
rect 4488 7896 4494 7948
rect 5994 7896 6000 7948
rect 6052 7896 6058 7948
rect 6104 7936 6132 7976
rect 6638 7964 6644 8016
rect 6696 7964 6702 8016
rect 7006 7964 7012 8016
rect 7064 8004 7070 8016
rect 10980 8013 11008 8044
rect 12728 8044 17816 8072
rect 7162 8007 7220 8013
rect 7162 8004 7174 8007
rect 7064 7976 7174 8004
rect 7064 7964 7070 7976
rect 7162 7973 7174 7976
rect 7208 7973 7220 8007
rect 9462 8007 9520 8013
rect 9462 8004 9474 8007
rect 7162 7967 7220 7973
rect 9048 7976 9474 8004
rect 6917 7939 6975 7945
rect 6917 7936 6929 7939
rect 6104 7908 6929 7936
rect 6917 7905 6929 7908
rect 6963 7905 6975 7939
rect 6917 7899 6975 7905
rect 8389 7939 8447 7945
rect 8389 7905 8401 7939
rect 8435 7936 8447 7939
rect 8435 7908 8708 7936
rect 8435 7905 8447 7908
rect 8389 7899 8447 7905
rect 3234 7868 3240 7880
rect 2516 7840 3240 7868
rect 3234 7828 3240 7840
rect 3292 7828 3298 7880
rect 8680 7877 8708 7908
rect 8665 7871 8723 7877
rect 8665 7837 8677 7871
rect 8711 7837 8723 7871
rect 8665 7831 8723 7837
rect 4246 7760 4252 7812
rect 4304 7760 4310 7812
rect 5810 7760 5816 7812
rect 5868 7760 5874 7812
rect 6270 7760 6276 7812
rect 6328 7760 6334 7812
rect 6825 7803 6883 7809
rect 6825 7769 6837 7803
rect 6871 7800 6883 7803
rect 6914 7800 6920 7812
rect 6871 7772 6920 7800
rect 6871 7769 6883 7772
rect 6825 7763 6883 7769
rect 6914 7760 6920 7772
rect 6972 7760 6978 7812
rect 8846 7760 8852 7812
rect 8904 7760 8910 7812
rect 1118 7692 1124 7744
rect 1176 7732 1182 7744
rect 2501 7735 2559 7741
rect 2501 7732 2513 7735
rect 1176 7704 2513 7732
rect 1176 7692 1182 7704
rect 2501 7701 2513 7704
rect 2547 7701 2559 7735
rect 2501 7695 2559 7701
rect 2866 7692 2872 7744
rect 2924 7732 2930 7744
rect 6641 7735 6699 7741
rect 6641 7732 6653 7735
rect 2924 7704 6653 7732
rect 2924 7692 2930 7704
rect 6641 7701 6653 7704
rect 6687 7732 6699 7735
rect 8110 7732 8116 7744
rect 6687 7704 8116 7732
rect 6687 7701 6699 7704
rect 6641 7695 6699 7701
rect 8110 7692 8116 7704
rect 8168 7692 8174 7744
rect 8202 7692 8208 7744
rect 8260 7732 8266 7744
rect 8297 7735 8355 7741
rect 8297 7732 8309 7735
rect 8260 7704 8309 7732
rect 8260 7692 8266 7704
rect 8297 7701 8309 7704
rect 8343 7701 8355 7735
rect 8297 7695 8355 7701
rect 8573 7735 8631 7741
rect 8573 7701 8585 7735
rect 8619 7732 8631 7735
rect 9048 7732 9076 7976
rect 9462 7973 9474 7976
rect 9508 7973 9520 8007
rect 9462 7967 9520 7973
rect 10965 8007 11023 8013
rect 10965 7973 10977 8007
rect 11011 7973 11023 8007
rect 12728 8004 12756 8044
rect 10965 7967 11023 7973
rect 11256 7976 12756 8004
rect 9217 7939 9275 7945
rect 9217 7905 9229 7939
rect 9263 7936 9275 7939
rect 9306 7936 9312 7948
rect 9263 7908 9312 7936
rect 9263 7905 9275 7908
rect 9217 7899 9275 7905
rect 9306 7896 9312 7908
rect 9364 7896 9370 7948
rect 9766 7896 9772 7948
rect 9824 7936 9830 7948
rect 9824 7908 10824 7936
rect 9824 7896 9830 7908
rect 9122 7828 9128 7880
rect 9180 7828 9186 7880
rect 10796 7868 10824 7908
rect 10870 7896 10876 7948
rect 10928 7936 10934 7948
rect 11149 7939 11207 7945
rect 11149 7936 11161 7939
rect 10928 7908 11161 7936
rect 10928 7896 10934 7908
rect 11149 7905 11161 7908
rect 11195 7905 11207 7939
rect 11149 7899 11207 7905
rect 11256 7868 11284 7976
rect 12161 7939 12219 7945
rect 12161 7905 12173 7939
rect 12207 7936 12219 7939
rect 12621 7939 12679 7945
rect 12207 7908 12296 7936
rect 12207 7905 12219 7908
rect 12161 7899 12219 7905
rect 10796 7840 11284 7868
rect 12268 7812 12296 7908
rect 12621 7905 12633 7939
rect 12667 7905 12679 7939
rect 12621 7899 12679 7905
rect 12342 7828 12348 7880
rect 12400 7828 12406 7880
rect 12250 7760 12256 7812
rect 12308 7800 12314 7812
rect 12437 7803 12495 7809
rect 12437 7800 12449 7803
rect 12308 7772 12449 7800
rect 12308 7760 12314 7772
rect 12437 7769 12449 7772
rect 12483 7769 12495 7803
rect 12636 7800 12664 7899
rect 12728 7868 12756 7976
rect 12805 8007 12863 8013
rect 12805 7973 12817 8007
rect 12851 8004 12863 8007
rect 13170 8004 13176 8016
rect 12851 7976 13176 8004
rect 12851 7973 12863 7976
rect 12805 7967 12863 7973
rect 13170 7964 13176 7976
rect 13228 7964 13234 8016
rect 14274 8004 14280 8016
rect 13280 7976 14280 8004
rect 13280 7945 13308 7976
rect 14274 7964 14280 7976
rect 14332 8004 14338 8016
rect 15197 8007 15255 8013
rect 15197 8004 15209 8007
rect 14332 7976 15209 8004
rect 14332 7964 14338 7976
rect 15197 7973 15209 7976
rect 15243 7973 15255 8007
rect 17034 8004 17040 8016
rect 15197 7967 15255 7973
rect 16132 7976 17040 8004
rect 12897 7939 12955 7945
rect 12897 7905 12909 7939
rect 12943 7936 12955 7939
rect 13265 7939 13323 7945
rect 13265 7936 13277 7939
rect 12943 7908 13277 7936
rect 12943 7905 12955 7908
rect 12897 7899 12955 7905
rect 13265 7905 13277 7908
rect 13311 7905 13323 7939
rect 13265 7899 13323 7905
rect 13630 7896 13636 7948
rect 13688 7896 13694 7948
rect 13906 7945 13912 7948
rect 13900 7899 13912 7945
rect 13906 7896 13912 7899
rect 13964 7896 13970 7948
rect 15102 7896 15108 7948
rect 15160 7896 15166 7948
rect 15286 7896 15292 7948
rect 15344 7896 15350 7948
rect 15562 7896 15568 7948
rect 15620 7896 15626 7948
rect 15654 7896 15660 7948
rect 15712 7936 15718 7948
rect 16132 7945 16160 7976
rect 17034 7964 17040 7976
rect 17092 8004 17098 8016
rect 17092 7976 17724 8004
rect 17092 7964 17098 7976
rect 16390 7945 16396 7948
rect 15841 7939 15899 7945
rect 15841 7936 15853 7939
rect 15712 7908 15853 7936
rect 15712 7896 15718 7908
rect 15841 7905 15853 7908
rect 15887 7905 15899 7939
rect 15841 7899 15899 7905
rect 16117 7939 16175 7945
rect 16117 7905 16129 7939
rect 16163 7905 16175 7939
rect 16384 7936 16396 7945
rect 16351 7908 16396 7936
rect 16117 7899 16175 7905
rect 16384 7899 16396 7908
rect 16390 7896 16396 7899
rect 16448 7896 16454 7948
rect 17696 7880 17724 7976
rect 17788 7936 17816 8044
rect 18322 8032 18328 8084
rect 18380 8072 18386 8084
rect 18601 8075 18659 8081
rect 18601 8072 18613 8075
rect 18380 8044 18613 8072
rect 18380 8032 18386 8044
rect 18601 8041 18613 8044
rect 18647 8041 18659 8075
rect 18601 8035 18659 8041
rect 20898 8032 20904 8084
rect 20956 8072 20962 8084
rect 20993 8075 21051 8081
rect 20993 8072 21005 8075
rect 20956 8044 21005 8072
rect 20956 8032 20962 8044
rect 20993 8041 21005 8044
rect 21039 8041 21051 8075
rect 20993 8035 21051 8041
rect 22649 8075 22707 8081
rect 22649 8041 22661 8075
rect 22695 8072 22707 8075
rect 22695 8044 22784 8072
rect 22695 8041 22707 8044
rect 22649 8035 22707 8041
rect 18509 8007 18567 8013
rect 18509 7973 18521 8007
rect 18555 8004 18567 8007
rect 21910 8004 21916 8016
rect 18555 7976 21916 8004
rect 18555 7973 18567 7976
rect 18509 7967 18567 7973
rect 21910 7964 21916 7976
rect 21968 7964 21974 8016
rect 19061 7939 19119 7945
rect 19061 7936 19073 7939
rect 17788 7908 19073 7936
rect 19061 7905 19073 7908
rect 19107 7905 19119 7939
rect 19061 7899 19119 7905
rect 19521 7939 19579 7945
rect 19521 7905 19533 7939
rect 19567 7905 19579 7939
rect 19521 7899 19579 7905
rect 13081 7871 13139 7877
rect 13081 7868 13093 7871
rect 12728 7840 13093 7868
rect 13081 7837 13093 7840
rect 13127 7837 13139 7871
rect 13081 7831 13139 7837
rect 13170 7828 13176 7880
rect 13228 7828 13234 7880
rect 13354 7828 13360 7880
rect 13412 7828 13418 7880
rect 17678 7828 17684 7880
rect 17736 7828 17742 7880
rect 18782 7828 18788 7880
rect 18840 7828 18846 7880
rect 18877 7871 18935 7877
rect 18877 7837 18889 7871
rect 18923 7837 18935 7871
rect 18877 7831 18935 7837
rect 18969 7871 19027 7877
rect 18969 7837 18981 7871
rect 19015 7868 19027 7871
rect 19536 7868 19564 7899
rect 19610 7896 19616 7948
rect 19668 7896 19674 7948
rect 19797 7939 19855 7945
rect 19797 7905 19809 7939
rect 19843 7905 19855 7939
rect 19797 7899 19855 7905
rect 19889 7939 19947 7945
rect 19889 7905 19901 7939
rect 19935 7936 19947 7939
rect 20070 7936 20076 7948
rect 19935 7908 20076 7936
rect 19935 7905 19947 7908
rect 19889 7899 19947 7905
rect 19702 7868 19708 7880
rect 19015 7840 19708 7868
rect 19015 7837 19027 7840
rect 18969 7831 19027 7837
rect 13372 7800 13400 7828
rect 12636 7772 13400 7800
rect 12437 7763 12495 7769
rect 14734 7760 14740 7812
rect 14792 7800 14798 7812
rect 15013 7803 15071 7809
rect 15013 7800 15025 7803
rect 14792 7772 15025 7800
rect 14792 7760 14798 7772
rect 15013 7769 15025 7772
rect 15059 7800 15071 7803
rect 15470 7800 15476 7812
rect 15059 7772 15476 7800
rect 15059 7769 15071 7772
rect 15013 7763 15071 7769
rect 15470 7760 15476 7772
rect 15528 7760 15534 7812
rect 17052 7772 17908 7800
rect 8619 7704 9076 7732
rect 8619 7701 8631 7704
rect 8573 7695 8631 7701
rect 11330 7692 11336 7744
rect 11388 7692 11394 7744
rect 11977 7735 12035 7741
rect 11977 7701 11989 7735
rect 12023 7732 12035 7735
rect 12066 7732 12072 7744
rect 12023 7704 12072 7732
rect 12023 7701 12035 7704
rect 11977 7695 12035 7701
rect 12066 7692 12072 7704
rect 12124 7692 12130 7744
rect 13541 7735 13599 7741
rect 13541 7701 13553 7735
rect 13587 7732 13599 7735
rect 13998 7732 14004 7744
rect 13587 7704 14004 7732
rect 13587 7701 13599 7704
rect 13541 7695 13599 7701
rect 13998 7692 14004 7704
rect 14056 7692 14062 7744
rect 14550 7692 14556 7744
rect 14608 7732 14614 7744
rect 17052 7732 17080 7772
rect 14608 7704 17080 7732
rect 17497 7735 17555 7741
rect 14608 7692 14614 7704
rect 17497 7701 17509 7735
rect 17543 7732 17555 7735
rect 17770 7732 17776 7744
rect 17543 7704 17776 7732
rect 17543 7701 17555 7704
rect 17497 7695 17555 7701
rect 17770 7692 17776 7704
rect 17828 7692 17834 7744
rect 17880 7732 17908 7772
rect 18138 7760 18144 7812
rect 18196 7800 18202 7812
rect 18892 7800 18920 7831
rect 19702 7828 19708 7840
rect 19760 7828 19766 7880
rect 19812 7868 19840 7899
rect 20070 7896 20076 7908
rect 20128 7896 20134 7948
rect 20254 7896 20260 7948
rect 20312 7936 20318 7948
rect 20349 7939 20407 7945
rect 20349 7936 20361 7939
rect 20312 7908 20361 7936
rect 20312 7896 20318 7908
rect 20349 7905 20361 7908
rect 20395 7905 20407 7939
rect 20349 7899 20407 7905
rect 20625 7939 20683 7945
rect 20625 7905 20637 7939
rect 20671 7936 20683 7939
rect 20809 7939 20867 7945
rect 20671 7908 20760 7936
rect 20671 7905 20683 7908
rect 20625 7899 20683 7905
rect 19978 7868 19984 7880
rect 19812 7840 19984 7868
rect 19978 7828 19984 7840
rect 20036 7868 20042 7880
rect 20165 7871 20223 7877
rect 20165 7868 20177 7871
rect 20036 7840 20177 7868
rect 20036 7828 20042 7840
rect 20165 7837 20177 7840
rect 20211 7837 20223 7871
rect 20165 7831 20223 7837
rect 19518 7800 19524 7812
rect 18196 7772 19524 7800
rect 18196 7760 18202 7772
rect 19518 7760 19524 7772
rect 19576 7760 19582 7812
rect 20732 7800 20760 7908
rect 20809 7905 20821 7939
rect 20855 7905 20867 7939
rect 20809 7899 20867 7905
rect 20824 7868 20852 7899
rect 20898 7896 20904 7948
rect 20956 7896 20962 7948
rect 21085 7939 21143 7945
rect 21085 7905 21097 7939
rect 21131 7936 21143 7939
rect 21358 7936 21364 7948
rect 21131 7908 21364 7936
rect 21131 7905 21143 7908
rect 21085 7899 21143 7905
rect 21100 7868 21128 7899
rect 21358 7896 21364 7908
rect 21416 7896 21422 7948
rect 21542 7945 21548 7948
rect 21536 7936 21548 7945
rect 21503 7908 21548 7936
rect 21536 7899 21548 7908
rect 21542 7896 21548 7899
rect 21600 7896 21606 7948
rect 22756 7945 22784 8044
rect 23014 8032 23020 8084
rect 23072 8072 23078 8084
rect 23293 8075 23351 8081
rect 23293 8072 23305 8075
rect 23072 8044 23305 8072
rect 23072 8032 23078 8044
rect 23293 8041 23305 8044
rect 23339 8041 23351 8075
rect 23293 8035 23351 8041
rect 24026 8032 24032 8084
rect 24084 8032 24090 8084
rect 24302 8032 24308 8084
rect 24360 8072 24366 8084
rect 24765 8075 24823 8081
rect 24765 8072 24777 8075
rect 24360 8044 24777 8072
rect 24360 8032 24366 8044
rect 24765 8041 24777 8044
rect 24811 8041 24823 8075
rect 24765 8035 24823 8041
rect 24854 8032 24860 8084
rect 24912 8032 24918 8084
rect 25593 8075 25651 8081
rect 25593 8041 25605 8075
rect 25639 8072 25651 8075
rect 25682 8072 25688 8084
rect 25639 8044 25688 8072
rect 25639 8041 25651 8044
rect 25593 8035 25651 8041
rect 25682 8032 25688 8044
rect 25740 8032 25746 8084
rect 26050 8072 26056 8084
rect 25976 8044 26056 8072
rect 23109 8007 23167 8013
rect 23109 7973 23121 8007
rect 23155 8004 23167 8007
rect 24044 8004 24072 8032
rect 23155 7976 23796 8004
rect 23155 7973 23167 7976
rect 23109 7967 23167 7973
rect 22741 7939 22799 7945
rect 22741 7905 22753 7939
rect 22787 7905 22799 7939
rect 22741 7899 22799 7905
rect 22925 7939 22983 7945
rect 22925 7905 22937 7939
rect 22971 7936 22983 7939
rect 23382 7936 23388 7948
rect 22971 7908 23388 7936
rect 22971 7905 22983 7908
rect 22925 7899 22983 7905
rect 20824 7840 21128 7868
rect 21266 7828 21272 7880
rect 21324 7828 21330 7880
rect 22756 7868 22784 7899
rect 23382 7896 23388 7908
rect 23440 7896 23446 7948
rect 23474 7896 23480 7948
rect 23532 7896 23538 7948
rect 23566 7896 23572 7948
rect 23624 7936 23630 7948
rect 23768 7945 23796 7976
rect 23952 7976 24072 8004
rect 23952 7945 23980 7976
rect 24118 7964 24124 8016
rect 24176 8004 24182 8016
rect 24397 8007 24455 8013
rect 24397 8004 24409 8007
rect 24176 7976 24409 8004
rect 24176 7964 24182 7976
rect 24397 7973 24409 7976
rect 24443 8004 24455 8007
rect 24486 8004 24492 8016
rect 24443 7976 24492 8004
rect 24443 7973 24455 7976
rect 24397 7967 24455 7973
rect 24486 7964 24492 7976
rect 24544 7964 24550 8016
rect 24581 8007 24639 8013
rect 24581 7973 24593 8007
rect 24627 8004 24639 8007
rect 25314 8004 25320 8016
rect 24627 7976 25320 8004
rect 24627 7973 24639 7976
rect 24581 7967 24639 7973
rect 25314 7964 25320 7976
rect 25372 7964 25378 8016
rect 23661 7939 23719 7945
rect 23661 7936 23673 7939
rect 23624 7908 23673 7936
rect 23624 7896 23630 7908
rect 23661 7905 23673 7908
rect 23707 7905 23719 7939
rect 23661 7899 23719 7905
rect 23753 7939 23811 7945
rect 23753 7905 23765 7939
rect 23799 7905 23811 7939
rect 23753 7899 23811 7905
rect 23937 7939 23995 7945
rect 23937 7905 23949 7939
rect 23983 7905 23995 7939
rect 23937 7899 23995 7905
rect 24026 7896 24032 7948
rect 24084 7896 24090 7948
rect 24213 7939 24271 7945
rect 24213 7905 24225 7939
rect 24259 7905 24271 7939
rect 24213 7899 24271 7905
rect 24228 7868 24256 7899
rect 24762 7896 24768 7948
rect 24820 7936 24826 7948
rect 25409 7939 25467 7945
rect 25409 7936 25421 7939
rect 24820 7908 25421 7936
rect 24820 7896 24826 7908
rect 25409 7905 25421 7908
rect 25455 7905 25467 7939
rect 25409 7899 25467 7905
rect 25866 7896 25872 7948
rect 25924 7896 25930 7948
rect 25976 7945 26004 8044
rect 26050 8032 26056 8044
rect 26108 8032 26114 8084
rect 26418 8032 26424 8084
rect 26476 8032 26482 8084
rect 25961 7939 26019 7945
rect 25961 7905 25973 7939
rect 26007 7905 26019 7939
rect 25961 7899 26019 7905
rect 26053 7939 26111 7945
rect 26053 7905 26065 7939
rect 26099 7905 26111 7939
rect 26053 7899 26111 7905
rect 22756 7840 24256 7868
rect 26068 7868 26096 7899
rect 26234 7896 26240 7948
rect 26292 7896 26298 7948
rect 27062 7896 27068 7948
rect 27120 7896 27126 7948
rect 26786 7868 26792 7880
rect 26068 7840 26792 7868
rect 26786 7828 26792 7840
rect 26844 7828 26850 7880
rect 20898 7800 20904 7812
rect 20732 7772 20904 7800
rect 20898 7760 20904 7772
rect 20956 7760 20962 7812
rect 23845 7803 23903 7809
rect 23845 7800 23857 7803
rect 22572 7772 23857 7800
rect 18414 7732 18420 7744
rect 17880 7704 18420 7732
rect 18414 7692 18420 7704
rect 18472 7692 18478 7744
rect 18874 7692 18880 7744
rect 18932 7732 18938 7744
rect 19337 7735 19395 7741
rect 19337 7732 19349 7735
rect 18932 7704 19349 7732
rect 18932 7692 18938 7704
rect 19337 7701 19349 7704
rect 19383 7701 19395 7735
rect 19337 7695 19395 7701
rect 21910 7692 21916 7744
rect 21968 7732 21974 7744
rect 22572 7732 22600 7772
rect 23845 7769 23857 7772
rect 23891 7769 23903 7803
rect 23845 7763 23903 7769
rect 21968 7704 22600 7732
rect 21968 7692 21974 7704
rect 552 7642 27416 7664
rect 552 7590 3756 7642
rect 3808 7590 3820 7642
rect 3872 7590 3884 7642
rect 3936 7590 3948 7642
rect 4000 7590 4012 7642
rect 4064 7590 10472 7642
rect 10524 7590 10536 7642
rect 10588 7590 10600 7642
rect 10652 7590 10664 7642
rect 10716 7590 10728 7642
rect 10780 7590 17188 7642
rect 17240 7590 17252 7642
rect 17304 7590 17316 7642
rect 17368 7590 17380 7642
rect 17432 7590 17444 7642
rect 17496 7590 23904 7642
rect 23956 7590 23968 7642
rect 24020 7590 24032 7642
rect 24084 7590 24096 7642
rect 24148 7590 24160 7642
rect 24212 7590 27416 7642
rect 552 7568 27416 7590
rect 2130 7488 2136 7540
rect 2188 7528 2194 7540
rect 2590 7528 2596 7540
rect 2188 7500 2596 7528
rect 2188 7488 2194 7500
rect 2590 7488 2596 7500
rect 2648 7488 2654 7540
rect 3234 7488 3240 7540
rect 3292 7488 3298 7540
rect 4249 7531 4307 7537
rect 4249 7497 4261 7531
rect 4295 7497 4307 7531
rect 4249 7491 4307 7497
rect 4264 7460 4292 7491
rect 4430 7488 4436 7540
rect 4488 7488 4494 7540
rect 5905 7531 5963 7537
rect 5905 7497 5917 7531
rect 5951 7497 5963 7531
rect 5905 7491 5963 7497
rect 4525 7463 4583 7469
rect 4525 7460 4537 7463
rect 4264 7432 4537 7460
rect 4525 7429 4537 7432
rect 4571 7429 4583 7463
rect 5920 7460 5948 7491
rect 5994 7488 6000 7540
rect 6052 7528 6058 7540
rect 6089 7531 6147 7537
rect 6089 7528 6101 7531
rect 6052 7500 6101 7528
rect 6052 7488 6058 7500
rect 6089 7497 6101 7500
rect 6135 7497 6147 7531
rect 6089 7491 6147 7497
rect 6638 7488 6644 7540
rect 6696 7528 6702 7540
rect 7285 7531 7343 7537
rect 7285 7528 7297 7531
rect 6696 7500 7297 7528
rect 6696 7488 6702 7500
rect 7285 7497 7297 7500
rect 7331 7497 7343 7531
rect 7285 7491 7343 7497
rect 9122 7488 9128 7540
rect 9180 7528 9186 7540
rect 9309 7531 9367 7537
rect 9309 7528 9321 7531
rect 9180 7500 9321 7528
rect 9180 7488 9186 7500
rect 9309 7497 9321 7500
rect 9355 7497 9367 7531
rect 9309 7491 9367 7497
rect 9582 7488 9588 7540
rect 9640 7528 9646 7540
rect 9953 7531 10011 7537
rect 9953 7528 9965 7531
rect 9640 7500 9965 7528
rect 9640 7488 9646 7500
rect 9953 7497 9965 7500
rect 9999 7497 10011 7531
rect 9953 7491 10011 7497
rect 10226 7488 10232 7540
rect 10284 7528 10290 7540
rect 10284 7500 10548 7528
rect 10284 7488 10290 7500
rect 8018 7460 8024 7472
rect 5920 7432 8024 7460
rect 4525 7423 4583 7429
rect 8018 7420 8024 7432
rect 8076 7420 8082 7472
rect 8846 7420 8852 7472
rect 8904 7460 8910 7472
rect 9600 7460 9628 7488
rect 8904 7432 9628 7460
rect 8904 7420 8910 7432
rect 2961 7395 3019 7401
rect 2961 7361 2973 7395
rect 3007 7392 3019 7395
rect 3326 7392 3332 7404
rect 3007 7364 3332 7392
rect 3007 7361 3019 7364
rect 2961 7355 3019 7361
rect 3326 7352 3332 7364
rect 3384 7392 3390 7404
rect 3421 7395 3479 7401
rect 3421 7392 3433 7395
rect 3384 7364 3433 7392
rect 3384 7352 3390 7364
rect 3421 7361 3433 7364
rect 3467 7361 3479 7395
rect 3421 7355 3479 7361
rect 4890 7352 4896 7404
rect 4948 7392 4954 7404
rect 5537 7395 5595 7401
rect 5537 7392 5549 7395
rect 4948 7364 5549 7392
rect 4948 7352 4954 7364
rect 845 7327 903 7333
rect 845 7293 857 7327
rect 891 7324 903 7327
rect 1394 7324 1400 7336
rect 891 7296 1400 7324
rect 891 7293 903 7296
rect 845 7287 903 7293
rect 1394 7284 1400 7296
rect 1452 7324 1458 7336
rect 1670 7324 1676 7336
rect 1452 7296 1676 7324
rect 1452 7284 1458 7296
rect 1670 7284 1676 7296
rect 1728 7284 1734 7336
rect 2501 7327 2559 7333
rect 2501 7293 2513 7327
rect 2547 7324 2559 7327
rect 2590 7324 2596 7336
rect 2547 7296 2596 7324
rect 2547 7293 2559 7296
rect 2501 7287 2559 7293
rect 2590 7284 2596 7296
rect 2648 7284 2654 7336
rect 3510 7284 3516 7336
rect 3568 7284 3574 7336
rect 3605 7327 3663 7333
rect 3605 7293 3617 7327
rect 3651 7293 3663 7327
rect 3605 7287 3663 7293
rect 3697 7327 3755 7333
rect 3697 7293 3709 7327
rect 3743 7324 3755 7327
rect 3743 7296 4568 7324
rect 3743 7293 3755 7296
rect 3697 7287 3755 7293
rect 1118 7265 1124 7268
rect 1112 7256 1124 7265
rect 1079 7228 1124 7256
rect 1112 7219 1124 7228
rect 1118 7216 1124 7219
rect 1176 7216 1182 7268
rect 3234 7216 3240 7268
rect 3292 7256 3298 7268
rect 3620 7256 3648 7287
rect 3292 7228 3648 7256
rect 3292 7216 3298 7228
rect 4062 7216 4068 7268
rect 4120 7216 4126 7268
rect 2222 7148 2228 7200
rect 2280 7148 2286 7200
rect 4246 7148 4252 7200
rect 4304 7197 4310 7200
rect 4304 7191 4323 7197
rect 4311 7157 4323 7191
rect 4540 7188 4568 7296
rect 4614 7284 4620 7336
rect 4672 7324 4678 7336
rect 4709 7327 4767 7333
rect 4709 7324 4721 7327
rect 4672 7296 4721 7324
rect 4672 7284 4678 7296
rect 4709 7293 4721 7296
rect 4755 7293 4767 7327
rect 4709 7287 4767 7293
rect 4798 7284 4804 7336
rect 4856 7284 4862 7336
rect 4982 7324 4988 7336
rect 4908 7296 4988 7324
rect 4908 7256 4936 7296
rect 4982 7284 4988 7296
rect 5040 7284 5046 7336
rect 5092 7333 5120 7364
rect 5537 7361 5549 7364
rect 5583 7392 5595 7395
rect 6181 7395 6239 7401
rect 6181 7392 6193 7395
rect 5583 7364 6193 7392
rect 5583 7361 5595 7364
rect 5537 7355 5595 7361
rect 6181 7361 6193 7364
rect 6227 7361 6239 7395
rect 6181 7355 6239 7361
rect 6270 7352 6276 7404
rect 6328 7392 6334 7404
rect 6914 7392 6920 7404
rect 6328 7364 6920 7392
rect 6328 7352 6334 7364
rect 5077 7327 5135 7333
rect 5077 7293 5089 7327
rect 5123 7293 5135 7327
rect 5077 7287 5135 7293
rect 5445 7327 5503 7333
rect 5445 7293 5457 7327
rect 5491 7324 5503 7327
rect 5994 7324 6000 7336
rect 5491 7296 6000 7324
rect 5491 7293 5503 7296
rect 5445 7287 5503 7293
rect 5994 7284 6000 7296
rect 6052 7284 6058 7336
rect 6454 7324 6460 7336
rect 6415 7296 6460 7324
rect 6454 7284 6460 7296
rect 6512 7284 6518 7336
rect 6564 7333 6592 7364
rect 6914 7352 6920 7364
rect 6972 7352 6978 7404
rect 7469 7395 7527 7401
rect 7469 7361 7481 7395
rect 7515 7392 7527 7395
rect 7650 7392 7656 7404
rect 7515 7364 7656 7392
rect 7515 7361 7527 7364
rect 7469 7355 7527 7361
rect 6549 7327 6607 7333
rect 6549 7293 6561 7327
rect 6595 7293 6607 7327
rect 6549 7287 6607 7293
rect 6641 7327 6699 7333
rect 6641 7293 6653 7327
rect 6687 7324 6699 7327
rect 6730 7324 6736 7336
rect 6687 7296 6736 7324
rect 6687 7293 6699 7296
rect 6641 7287 6699 7293
rect 6730 7284 6736 7296
rect 6788 7284 6794 7336
rect 6822 7284 6828 7336
rect 6880 7284 6886 7336
rect 7193 7327 7251 7333
rect 7193 7293 7205 7327
rect 7239 7324 7251 7327
rect 7484 7324 7512 7355
rect 7650 7352 7656 7364
rect 7708 7392 7714 7404
rect 8113 7395 8171 7401
rect 8113 7392 8125 7395
rect 7708 7364 8125 7392
rect 7708 7352 7714 7364
rect 8113 7361 8125 7364
rect 8159 7361 8171 7395
rect 8113 7355 8171 7361
rect 9398 7352 9404 7404
rect 9456 7392 9462 7404
rect 9585 7395 9643 7401
rect 9585 7392 9597 7395
rect 9456 7364 9597 7392
rect 9456 7352 9462 7364
rect 9585 7361 9597 7364
rect 9631 7392 9643 7395
rect 9631 7364 10364 7392
rect 9631 7361 9643 7364
rect 9585 7355 9643 7361
rect 7239 7296 7512 7324
rect 7561 7327 7619 7333
rect 7239 7293 7251 7296
rect 7193 7287 7251 7293
rect 7561 7293 7573 7327
rect 7607 7293 7619 7327
rect 7561 7287 7619 7293
rect 8021 7327 8079 7333
rect 8021 7293 8033 7327
rect 8067 7324 8079 7327
rect 8067 7296 8156 7324
rect 8067 7293 8079 7296
rect 8021 7287 8079 7293
rect 5353 7259 5411 7265
rect 5353 7256 5365 7259
rect 4908 7228 5365 7256
rect 5353 7225 5365 7228
rect 5399 7225 5411 7259
rect 6472 7256 6500 7284
rect 7101 7259 7159 7265
rect 7101 7256 7113 7259
rect 5353 7219 5411 7225
rect 5460 7228 6040 7256
rect 6472 7228 7113 7256
rect 4706 7188 4712 7200
rect 4540 7160 4712 7188
rect 4304 7151 4323 7157
rect 4304 7148 4310 7151
rect 4706 7148 4712 7160
rect 4764 7188 4770 7200
rect 5460 7188 5488 7228
rect 4764 7160 5488 7188
rect 4764 7148 4770 7160
rect 5902 7148 5908 7200
rect 5960 7148 5966 7200
rect 6012 7188 6040 7228
rect 7101 7225 7113 7228
rect 7147 7225 7159 7259
rect 7576 7256 7604 7287
rect 7742 7256 7748 7268
rect 7576 7228 7748 7256
rect 7101 7219 7159 7225
rect 7742 7216 7748 7228
rect 7800 7256 7806 7268
rect 8128 7256 8156 7296
rect 8202 7284 8208 7336
rect 8260 7324 8266 7336
rect 8389 7327 8447 7333
rect 8389 7324 8401 7327
rect 8260 7296 8401 7324
rect 8260 7284 8266 7296
rect 8389 7293 8401 7296
rect 8435 7293 8447 7327
rect 8389 7287 8447 7293
rect 9493 7327 9551 7333
rect 9493 7293 9505 7327
rect 9539 7293 9551 7327
rect 9493 7287 9551 7293
rect 8570 7256 8576 7268
rect 7800 7228 8064 7256
rect 8128 7228 8576 7256
rect 7800 7216 7806 7228
rect 7006 7188 7012 7200
rect 6012 7160 7012 7188
rect 7006 7148 7012 7160
rect 7064 7148 7070 7200
rect 7834 7148 7840 7200
rect 7892 7188 7898 7200
rect 7929 7191 7987 7197
rect 7929 7188 7941 7191
rect 7892 7160 7941 7188
rect 7892 7148 7898 7160
rect 7929 7157 7941 7160
rect 7975 7157 7987 7191
rect 8036 7188 8064 7228
rect 8570 7216 8576 7228
rect 8628 7216 8634 7268
rect 9508 7256 9536 7287
rect 9674 7284 9680 7336
rect 9732 7284 9738 7336
rect 9766 7284 9772 7336
rect 9824 7284 9830 7336
rect 10137 7327 10195 7333
rect 10137 7293 10149 7327
rect 10183 7321 10195 7327
rect 10336 7324 10364 7364
rect 10520 7333 10548 7500
rect 13170 7488 13176 7540
rect 13228 7528 13234 7540
rect 13228 7500 13768 7528
rect 13228 7488 13234 7500
rect 12250 7420 12256 7472
rect 12308 7460 12314 7472
rect 13633 7463 13691 7469
rect 13633 7460 13645 7463
rect 12308 7432 13645 7460
rect 12308 7420 12314 7432
rect 12636 7401 12664 7432
rect 13633 7429 13645 7432
rect 13679 7429 13691 7463
rect 13740 7460 13768 7500
rect 13906 7488 13912 7540
rect 13964 7528 13970 7540
rect 14093 7531 14151 7537
rect 14093 7528 14105 7531
rect 13964 7500 14105 7528
rect 13964 7488 13970 7500
rect 14093 7497 14105 7500
rect 14139 7497 14151 7531
rect 14093 7491 14151 7497
rect 14182 7488 14188 7540
rect 14240 7528 14246 7540
rect 14829 7531 14887 7537
rect 14829 7528 14841 7531
rect 14240 7500 14841 7528
rect 14240 7488 14246 7500
rect 14829 7497 14841 7500
rect 14875 7497 14887 7531
rect 14829 7491 14887 7497
rect 15654 7488 15660 7540
rect 15712 7488 15718 7540
rect 16209 7531 16267 7537
rect 16209 7497 16221 7531
rect 16255 7528 16267 7531
rect 16298 7528 16304 7540
rect 16255 7500 16304 7528
rect 16255 7497 16267 7500
rect 16209 7491 16267 7497
rect 16298 7488 16304 7500
rect 16356 7488 16362 7540
rect 16393 7531 16451 7537
rect 16393 7497 16405 7531
rect 16439 7528 16451 7531
rect 16482 7528 16488 7540
rect 16439 7500 16488 7528
rect 16439 7497 16451 7500
rect 16393 7491 16451 7497
rect 16482 7488 16488 7500
rect 16540 7488 16546 7540
rect 18325 7531 18383 7537
rect 18325 7528 18337 7531
rect 17328 7500 18337 7528
rect 15672 7460 15700 7488
rect 13740 7432 15056 7460
rect 13633 7423 13691 7429
rect 12345 7395 12403 7401
rect 12345 7392 12357 7395
rect 11808 7364 12357 7392
rect 10413 7327 10471 7333
rect 10413 7324 10425 7327
rect 10183 7293 10272 7321
rect 10336 7296 10425 7324
rect 10137 7287 10195 7293
rect 10244 7256 10272 7293
rect 10413 7293 10425 7296
rect 10459 7293 10471 7327
rect 10413 7287 10471 7293
rect 10505 7327 10563 7333
rect 10505 7293 10517 7327
rect 10551 7293 10563 7327
rect 10505 7287 10563 7293
rect 10689 7327 10747 7333
rect 10689 7293 10701 7327
rect 10735 7324 10747 7327
rect 11330 7324 11336 7336
rect 10735 7296 11336 7324
rect 10735 7293 10747 7296
rect 10689 7287 10747 7293
rect 11330 7284 11336 7296
rect 11388 7284 11394 7336
rect 11808 7333 11836 7364
rect 12345 7361 12357 7364
rect 12391 7361 12403 7395
rect 12345 7355 12403 7361
rect 12621 7395 12679 7401
rect 12621 7361 12633 7395
rect 12667 7361 12679 7395
rect 12621 7355 12679 7361
rect 13998 7352 14004 7404
rect 14056 7352 14062 7404
rect 14550 7392 14556 7404
rect 14200 7364 14556 7392
rect 11793 7327 11851 7333
rect 11793 7293 11805 7327
rect 11839 7293 11851 7327
rect 11793 7287 11851 7293
rect 12066 7284 12072 7336
rect 12124 7284 12130 7336
rect 12253 7327 12311 7333
rect 12253 7293 12265 7327
rect 12299 7324 12311 7327
rect 12526 7324 12532 7336
rect 12299 7296 12532 7324
rect 12299 7293 12311 7296
rect 12253 7287 12311 7293
rect 12526 7284 12532 7296
rect 12584 7284 12590 7336
rect 12713 7327 12771 7333
rect 12713 7293 12725 7327
rect 12759 7293 12771 7327
rect 12713 7287 12771 7293
rect 12805 7327 12863 7333
rect 12805 7293 12817 7327
rect 12851 7324 12863 7327
rect 14200 7324 14228 7364
rect 14550 7352 14556 7364
rect 14608 7352 14614 7404
rect 15028 7336 15056 7432
rect 15304 7432 15700 7460
rect 15841 7463 15899 7469
rect 12851 7296 14228 7324
rect 14277 7327 14335 7333
rect 12851 7293 12863 7296
rect 12805 7287 12863 7293
rect 14277 7293 14289 7327
rect 14323 7324 14335 7327
rect 14366 7324 14372 7336
rect 14323 7296 14372 7324
rect 14323 7293 14335 7296
rect 14277 7287 14335 7293
rect 10597 7259 10655 7265
rect 10597 7256 10609 7259
rect 9508 7228 10609 7256
rect 10597 7225 10609 7228
rect 10643 7225 10655 7259
rect 10597 7219 10655 7225
rect 12342 7216 12348 7268
rect 12400 7256 12406 7268
rect 12728 7256 12756 7287
rect 12400 7228 12756 7256
rect 12400 7216 12406 7228
rect 8757 7191 8815 7197
rect 8757 7188 8769 7191
rect 8036 7160 8769 7188
rect 7929 7151 7987 7157
rect 8757 7157 8769 7160
rect 8803 7157 8815 7191
rect 8757 7151 8815 7157
rect 9674 7148 9680 7200
rect 9732 7188 9738 7200
rect 10318 7188 10324 7200
rect 9732 7160 10324 7188
rect 9732 7148 9738 7160
rect 10318 7148 10324 7160
rect 10376 7148 10382 7200
rect 11330 7148 11336 7200
rect 11388 7188 11394 7200
rect 11609 7191 11667 7197
rect 11609 7188 11621 7191
rect 11388 7160 11621 7188
rect 11388 7148 11394 7160
rect 11609 7157 11621 7160
rect 11655 7157 11667 7191
rect 11609 7151 11667 7157
rect 11698 7148 11704 7200
rect 11756 7188 11762 7200
rect 12820 7188 12848 7287
rect 14366 7284 14372 7296
rect 14424 7284 14430 7336
rect 15010 7284 15016 7336
rect 15068 7284 15074 7336
rect 15105 7327 15163 7333
rect 15105 7293 15117 7327
rect 15151 7324 15163 7327
rect 15194 7324 15200 7336
rect 15151 7296 15200 7324
rect 15151 7293 15163 7296
rect 15105 7287 15163 7293
rect 15194 7284 15200 7296
rect 15252 7284 15258 7336
rect 15304 7333 15332 7432
rect 15841 7429 15853 7463
rect 15887 7460 15899 7463
rect 16669 7463 16727 7469
rect 16669 7460 16681 7463
rect 15887 7432 16681 7460
rect 15887 7429 15899 7432
rect 15841 7423 15899 7429
rect 16669 7429 16681 7432
rect 16715 7429 16727 7463
rect 16669 7423 16727 7429
rect 15856 7392 15884 7423
rect 15672 7364 15884 7392
rect 15289 7327 15347 7333
rect 15289 7293 15301 7327
rect 15335 7293 15347 7327
rect 15289 7287 15347 7293
rect 15381 7327 15439 7333
rect 15381 7293 15393 7327
rect 15427 7324 15439 7327
rect 15562 7324 15568 7336
rect 15427 7296 15568 7324
rect 15427 7293 15439 7296
rect 15381 7287 15439 7293
rect 15562 7284 15568 7296
rect 15620 7324 15626 7336
rect 15672 7324 15700 7364
rect 15620 7296 15700 7324
rect 15749 7327 15807 7333
rect 15620 7284 15626 7296
rect 15749 7293 15761 7327
rect 15795 7324 15807 7327
rect 15795 7296 16712 7324
rect 15795 7293 15807 7296
rect 15749 7287 15807 7293
rect 16684 7268 16712 7296
rect 16942 7284 16948 7336
rect 17000 7284 17006 7336
rect 17034 7284 17040 7336
rect 17092 7284 17098 7336
rect 17126 7284 17132 7336
rect 17184 7284 17190 7336
rect 17328 7333 17356 7500
rect 18325 7497 18337 7500
rect 18371 7497 18383 7531
rect 18325 7491 18383 7497
rect 18414 7488 18420 7540
rect 18472 7528 18478 7540
rect 18472 7500 18828 7528
rect 18472 7488 18478 7500
rect 17681 7463 17739 7469
rect 17681 7429 17693 7463
rect 17727 7460 17739 7463
rect 17862 7460 17868 7472
rect 17727 7432 17868 7460
rect 17727 7429 17739 7432
rect 17681 7423 17739 7429
rect 17862 7420 17868 7432
rect 17920 7420 17926 7472
rect 17954 7420 17960 7472
rect 18012 7460 18018 7472
rect 18693 7463 18751 7469
rect 18693 7460 18705 7463
rect 18012 7432 18705 7460
rect 18012 7420 18018 7432
rect 18693 7429 18705 7432
rect 18739 7429 18751 7463
rect 18800 7460 18828 7500
rect 18874 7488 18880 7540
rect 18932 7488 18938 7540
rect 19518 7488 19524 7540
rect 19576 7488 19582 7540
rect 20898 7488 20904 7540
rect 20956 7528 20962 7540
rect 21634 7528 21640 7540
rect 20956 7500 21640 7528
rect 20956 7488 20962 7500
rect 21634 7488 21640 7500
rect 21692 7488 21698 7540
rect 21726 7488 21732 7540
rect 21784 7488 21790 7540
rect 25866 7488 25872 7540
rect 25924 7528 25930 7540
rect 26329 7531 26387 7537
rect 26329 7528 26341 7531
rect 25924 7500 26341 7528
rect 25924 7488 25930 7500
rect 26329 7497 26341 7500
rect 26375 7497 26387 7531
rect 26329 7491 26387 7497
rect 19429 7463 19487 7469
rect 18800 7432 18920 7460
rect 18693 7423 18751 7429
rect 18782 7392 18788 7404
rect 17880 7364 18788 7392
rect 17880 7333 17908 7364
rect 18782 7352 18788 7364
rect 18840 7352 18846 7404
rect 18892 7392 18920 7432
rect 19429 7429 19441 7463
rect 19475 7460 19487 7463
rect 19610 7460 19616 7472
rect 19475 7432 19616 7460
rect 19475 7429 19487 7432
rect 19429 7423 19487 7429
rect 19610 7420 19616 7432
rect 19668 7420 19674 7472
rect 19720 7432 22094 7460
rect 19720 7392 19748 7432
rect 18892 7364 19748 7392
rect 21376 7364 21864 7392
rect 17313 7327 17371 7333
rect 17313 7293 17325 7327
rect 17359 7293 17371 7327
rect 17313 7287 17371 7293
rect 17865 7327 17923 7333
rect 17865 7293 17877 7327
rect 17911 7293 17923 7327
rect 17865 7287 17923 7293
rect 16666 7216 16672 7268
rect 16724 7256 16730 7268
rect 17328 7256 17356 7287
rect 18138 7284 18144 7336
rect 18196 7284 18202 7336
rect 18230 7284 18236 7336
rect 18288 7284 18294 7336
rect 18417 7327 18475 7333
rect 18417 7293 18429 7327
rect 18463 7293 18475 7327
rect 19702 7324 19708 7336
rect 18417 7287 18475 7293
rect 18984 7296 19708 7324
rect 16724 7228 17356 7256
rect 16724 7216 16730 7228
rect 17770 7216 17776 7268
rect 17828 7256 17834 7268
rect 18432 7256 18460 7287
rect 18984 7256 19012 7296
rect 19702 7284 19708 7296
rect 19760 7284 19766 7336
rect 19978 7284 19984 7336
rect 20036 7284 20042 7336
rect 20070 7284 20076 7336
rect 20128 7324 20134 7336
rect 21376 7333 21404 7364
rect 20165 7327 20223 7333
rect 20165 7324 20177 7327
rect 20128 7296 20177 7324
rect 20128 7284 20134 7296
rect 20165 7293 20177 7296
rect 20211 7293 20223 7327
rect 20165 7287 20223 7293
rect 21361 7327 21419 7333
rect 21361 7293 21373 7327
rect 21407 7293 21419 7327
rect 21361 7287 21419 7293
rect 21453 7327 21511 7333
rect 21453 7293 21465 7327
rect 21499 7324 21511 7327
rect 21836 7324 21864 7364
rect 21910 7352 21916 7404
rect 21968 7352 21974 7404
rect 22066 7392 22094 7432
rect 22189 7395 22247 7401
rect 22189 7392 22201 7395
rect 22066 7364 22201 7392
rect 22189 7361 22201 7364
rect 22235 7361 22247 7395
rect 22189 7355 22247 7361
rect 26878 7352 26884 7404
rect 26936 7352 26942 7404
rect 22002 7324 22008 7336
rect 21499 7296 21772 7324
rect 21836 7296 22008 7324
rect 21499 7293 21511 7296
rect 21453 7287 21511 7293
rect 17828 7228 18460 7256
rect 18800 7228 19012 7256
rect 17828 7216 17834 7228
rect 11756 7160 12848 7188
rect 11756 7148 11762 7160
rect 13078 7148 13084 7200
rect 13136 7188 13142 7200
rect 13541 7191 13599 7197
rect 13541 7188 13553 7191
rect 13136 7160 13553 7188
rect 13136 7148 13142 7160
rect 13541 7157 13553 7160
rect 13587 7157 13599 7191
rect 13541 7151 13599 7157
rect 16206 7148 16212 7200
rect 16264 7148 16270 7200
rect 18049 7191 18107 7197
rect 18049 7157 18061 7191
rect 18095 7188 18107 7191
rect 18800 7188 18828 7228
rect 19058 7216 19064 7268
rect 19116 7256 19122 7268
rect 21174 7256 21180 7268
rect 19116 7228 21180 7256
rect 19116 7216 19122 7228
rect 21174 7216 21180 7228
rect 21232 7216 21238 7268
rect 21637 7259 21695 7265
rect 21637 7225 21649 7259
rect 21683 7225 21695 7259
rect 21744 7256 21772 7296
rect 22002 7284 22008 7296
rect 22060 7284 22066 7336
rect 22097 7327 22155 7333
rect 22097 7293 22109 7327
rect 22143 7324 22155 7327
rect 23014 7324 23020 7336
rect 22143 7296 23020 7324
rect 22143 7293 22155 7296
rect 22097 7287 22155 7293
rect 22112 7256 22140 7287
rect 23014 7284 23020 7296
rect 23072 7324 23078 7336
rect 23201 7327 23259 7333
rect 23201 7324 23213 7327
rect 23072 7296 23213 7324
rect 23072 7284 23078 7296
rect 23201 7293 23213 7296
rect 23247 7293 23259 7327
rect 23201 7287 23259 7293
rect 23290 7284 23296 7336
rect 23348 7284 23354 7336
rect 23477 7327 23535 7333
rect 23477 7293 23489 7327
rect 23523 7293 23535 7327
rect 23477 7287 23535 7293
rect 21744 7228 22140 7256
rect 23492 7256 23520 7287
rect 23566 7284 23572 7336
rect 23624 7284 23630 7336
rect 24397 7327 24455 7333
rect 24397 7293 24409 7327
rect 24443 7324 24455 7327
rect 24578 7324 24584 7336
rect 24443 7296 24584 7324
rect 24443 7293 24455 7296
rect 24397 7287 24455 7293
rect 24578 7284 24584 7296
rect 24636 7284 24642 7336
rect 24673 7327 24731 7333
rect 24673 7293 24685 7327
rect 24719 7324 24731 7327
rect 24719 7296 25084 7324
rect 24719 7293 24731 7296
rect 24673 7287 24731 7293
rect 25056 7268 25084 7296
rect 23750 7256 23756 7268
rect 23492 7228 23756 7256
rect 21637 7219 21695 7225
rect 18095 7160 18828 7188
rect 18861 7191 18919 7197
rect 18095 7157 18107 7160
rect 18049 7151 18107 7157
rect 18861 7157 18873 7191
rect 18907 7188 18919 7191
rect 19518 7188 19524 7200
rect 18907 7160 19524 7188
rect 18907 7157 18919 7160
rect 18861 7151 18919 7157
rect 19518 7148 19524 7160
rect 19576 7148 19582 7200
rect 21652 7188 21680 7219
rect 23750 7216 23756 7228
rect 23808 7216 23814 7268
rect 24918 7259 24976 7265
rect 24918 7256 24930 7259
rect 24596 7228 24930 7256
rect 21910 7188 21916 7200
rect 21652 7160 21916 7188
rect 21910 7148 21916 7160
rect 21968 7148 21974 7200
rect 22554 7148 22560 7200
rect 22612 7188 22618 7200
rect 24596 7197 24624 7228
rect 24918 7225 24930 7228
rect 24964 7225 24976 7259
rect 24918 7219 24976 7225
rect 25038 7216 25044 7268
rect 25096 7216 25102 7268
rect 23017 7191 23075 7197
rect 23017 7188 23029 7191
rect 22612 7160 23029 7188
rect 22612 7148 22618 7160
rect 23017 7157 23029 7160
rect 23063 7157 23075 7191
rect 23017 7151 23075 7157
rect 24581 7191 24639 7197
rect 24581 7157 24593 7191
rect 24627 7157 24639 7191
rect 24581 7151 24639 7157
rect 26050 7148 26056 7200
rect 26108 7148 26114 7200
rect 552 7098 27576 7120
rect 552 7046 7114 7098
rect 7166 7046 7178 7098
rect 7230 7046 7242 7098
rect 7294 7046 7306 7098
rect 7358 7046 7370 7098
rect 7422 7046 13830 7098
rect 13882 7046 13894 7098
rect 13946 7046 13958 7098
rect 14010 7046 14022 7098
rect 14074 7046 14086 7098
rect 14138 7046 20546 7098
rect 20598 7046 20610 7098
rect 20662 7046 20674 7098
rect 20726 7046 20738 7098
rect 20790 7046 20802 7098
rect 20854 7046 27262 7098
rect 27314 7046 27326 7098
rect 27378 7046 27390 7098
rect 27442 7046 27454 7098
rect 27506 7046 27518 7098
rect 27570 7046 27576 7098
rect 552 7024 27576 7046
rect 2130 6944 2136 6996
rect 2188 6944 2194 6996
rect 5902 6944 5908 6996
rect 5960 6984 5966 6996
rect 5997 6987 6055 6993
rect 5997 6984 6009 6987
rect 5960 6956 6009 6984
rect 5960 6944 5966 6956
rect 5997 6953 6009 6956
rect 6043 6953 6055 6987
rect 6822 6984 6828 6996
rect 5997 6947 6055 6953
rect 6196 6956 6828 6984
rect 2409 6919 2467 6925
rect 2409 6885 2421 6919
rect 2455 6916 2467 6919
rect 2590 6916 2596 6928
rect 2455 6888 2596 6916
rect 2455 6885 2467 6888
rect 2409 6879 2467 6885
rect 2590 6876 2596 6888
rect 2648 6916 2654 6928
rect 2648 6888 3096 6916
rect 2648 6876 2654 6888
rect 2041 6851 2099 6857
rect 2041 6817 2053 6851
rect 2087 6848 2099 6851
rect 2130 6848 2136 6860
rect 2087 6820 2136 6848
rect 2087 6817 2099 6820
rect 2041 6811 2099 6817
rect 2130 6808 2136 6820
rect 2188 6808 2194 6860
rect 2222 6808 2228 6860
rect 2280 6848 2286 6860
rect 2317 6851 2375 6857
rect 2317 6848 2329 6851
rect 2280 6820 2329 6848
rect 2280 6808 2286 6820
rect 2317 6817 2329 6820
rect 2363 6817 2375 6851
rect 2317 6811 2375 6817
rect 2501 6851 2559 6857
rect 2501 6817 2513 6851
rect 2547 6817 2559 6851
rect 2501 6811 2559 6817
rect 2849 6851 2907 6857
rect 2849 6817 2861 6851
rect 2895 6848 2907 6851
rect 2895 6817 2912 6848
rect 2849 6811 2912 6817
rect 2148 6780 2176 6808
rect 2516 6780 2544 6811
rect 2148 6752 2544 6780
rect 2593 6783 2651 6789
rect 2593 6749 2605 6783
rect 2639 6780 2651 6783
rect 2682 6780 2688 6792
rect 2639 6752 2688 6780
rect 2639 6749 2651 6752
rect 2593 6743 2651 6749
rect 2682 6740 2688 6752
rect 2740 6740 2746 6792
rect 2884 6780 2912 6811
rect 2958 6808 2964 6860
rect 3016 6808 3022 6860
rect 3068 6857 3096 6888
rect 3326 6876 3332 6928
rect 3384 6876 3390 6928
rect 4525 6919 4583 6925
rect 4525 6885 4537 6919
rect 4571 6885 4583 6919
rect 4525 6879 4583 6885
rect 3053 6851 3111 6857
rect 3053 6817 3065 6851
rect 3099 6817 3111 6851
rect 3053 6811 3111 6817
rect 3234 6808 3240 6860
rect 3292 6848 3298 6860
rect 3513 6851 3571 6857
rect 3513 6848 3525 6851
rect 3292 6820 3525 6848
rect 3292 6808 3298 6820
rect 3513 6817 3525 6820
rect 3559 6817 3571 6851
rect 3513 6811 3571 6817
rect 3602 6808 3608 6860
rect 3660 6808 3666 6860
rect 4246 6808 4252 6860
rect 4304 6848 4310 6860
rect 4540 6848 4568 6879
rect 4304 6820 4568 6848
rect 4304 6808 4310 6820
rect 4890 6808 4896 6860
rect 4948 6808 4954 6860
rect 4982 6808 4988 6860
rect 5040 6808 5046 6860
rect 5074 6808 5080 6860
rect 5132 6808 5138 6860
rect 5258 6808 5264 6860
rect 5316 6808 5322 6860
rect 5994 6808 6000 6860
rect 6052 6848 6058 6860
rect 6196 6857 6224 6956
rect 6822 6944 6828 6956
rect 6880 6944 6886 6996
rect 6914 6944 6920 6996
rect 6972 6984 6978 6996
rect 7469 6987 7527 6993
rect 7469 6984 7481 6987
rect 6972 6956 7481 6984
rect 6972 6944 6978 6956
rect 7469 6953 7481 6956
rect 7515 6953 7527 6987
rect 7469 6947 7527 6953
rect 7650 6944 7656 6996
rect 7708 6944 7714 6996
rect 11698 6984 11704 6996
rect 7760 6956 11704 6984
rect 6932 6916 6960 6944
rect 6564 6888 6960 6916
rect 6181 6851 6239 6857
rect 6181 6848 6193 6851
rect 6052 6820 6193 6848
rect 6052 6808 6058 6820
rect 6181 6817 6193 6820
rect 6227 6817 6239 6851
rect 6181 6811 6239 6817
rect 6273 6851 6331 6857
rect 6273 6817 6285 6851
rect 6319 6817 6331 6851
rect 6273 6811 6331 6817
rect 4433 6783 4491 6789
rect 2884 6752 3556 6780
rect 3142 6672 3148 6724
rect 3200 6712 3206 6724
rect 3329 6715 3387 6721
rect 3329 6712 3341 6715
rect 3200 6684 3341 6712
rect 3200 6672 3206 6684
rect 3329 6681 3341 6684
rect 3375 6681 3387 6715
rect 3329 6675 3387 6681
rect 3528 6656 3556 6752
rect 4433 6749 4445 6783
rect 4479 6780 4491 6783
rect 4614 6780 4620 6792
rect 4479 6752 4620 6780
rect 4479 6749 4491 6752
rect 4433 6743 4491 6749
rect 4614 6740 4620 6752
rect 4672 6740 4678 6792
rect 4709 6783 4767 6789
rect 4709 6749 4721 6783
rect 4755 6780 4767 6783
rect 4798 6780 4804 6792
rect 4755 6752 4804 6780
rect 4755 6749 4767 6752
rect 4709 6743 4767 6749
rect 4798 6740 4804 6752
rect 4856 6780 4862 6792
rect 5445 6783 5503 6789
rect 5445 6780 5457 6783
rect 4856 6752 5457 6780
rect 4856 6740 4862 6752
rect 5445 6749 5457 6752
rect 5491 6749 5503 6783
rect 6288 6780 6316 6811
rect 6454 6808 6460 6860
rect 6512 6808 6518 6860
rect 6564 6857 6592 6888
rect 7006 6876 7012 6928
rect 7064 6916 7070 6928
rect 7760 6916 7788 6956
rect 11698 6944 11704 6956
rect 11756 6944 11762 6996
rect 12526 6944 12532 6996
rect 12584 6984 12590 6996
rect 12805 6987 12863 6993
rect 12805 6984 12817 6987
rect 12584 6956 12817 6984
rect 12584 6944 12590 6956
rect 12805 6953 12817 6956
rect 12851 6953 12863 6987
rect 12805 6947 12863 6953
rect 13354 6944 13360 6996
rect 13412 6984 13418 6996
rect 13633 6987 13691 6993
rect 13633 6984 13645 6987
rect 13412 6956 13645 6984
rect 13412 6944 13418 6956
rect 13633 6953 13645 6956
rect 13679 6953 13691 6987
rect 13633 6947 13691 6953
rect 16206 6944 16212 6996
rect 16264 6984 16270 6996
rect 16485 6987 16543 6993
rect 16485 6984 16497 6987
rect 16264 6956 16497 6984
rect 16264 6944 16270 6956
rect 16485 6953 16497 6956
rect 16531 6953 16543 6987
rect 19058 6984 19064 6996
rect 16485 6947 16543 6953
rect 16868 6956 19064 6984
rect 7064 6888 7788 6916
rect 7064 6876 7070 6888
rect 8662 6876 8668 6928
rect 8720 6916 8726 6928
rect 11232 6919 11290 6925
rect 8720 6888 11192 6916
rect 8720 6876 8726 6888
rect 6549 6851 6607 6857
rect 6549 6817 6561 6851
rect 6595 6817 6607 6851
rect 6549 6811 6607 6817
rect 6638 6808 6644 6860
rect 6696 6808 6702 6860
rect 6822 6808 6828 6860
rect 6880 6808 6886 6860
rect 9306 6808 9312 6860
rect 9364 6848 9370 6860
rect 10965 6851 11023 6857
rect 10965 6848 10977 6851
rect 9364 6820 10977 6848
rect 9364 6808 9370 6820
rect 10965 6817 10977 6820
rect 11011 6817 11023 6851
rect 11164 6848 11192 6888
rect 11232 6885 11244 6919
rect 11278 6916 11290 6919
rect 11330 6916 11336 6928
rect 11278 6888 11336 6916
rect 11278 6885 11290 6888
rect 11232 6879 11290 6885
rect 11330 6876 11336 6888
rect 11388 6876 11394 6928
rect 16868 6916 16896 6956
rect 19058 6944 19064 6956
rect 19116 6944 19122 6996
rect 19610 6944 19616 6996
rect 19668 6944 19674 6996
rect 19702 6944 19708 6996
rect 19760 6984 19766 6996
rect 20165 6987 20223 6993
rect 20165 6984 20177 6987
rect 19760 6956 20177 6984
rect 19760 6944 19766 6956
rect 20165 6953 20177 6956
rect 20211 6953 20223 6987
rect 20165 6947 20223 6953
rect 24486 6944 24492 6996
rect 24544 6984 24550 6996
rect 24544 6956 25636 6984
rect 24544 6944 24550 6956
rect 17221 6919 17279 6925
rect 17221 6916 17233 6919
rect 11440 6888 16896 6916
rect 16960 6888 17233 6916
rect 11440 6848 11468 6888
rect 16960 6860 16988 6888
rect 17221 6885 17233 6888
rect 17267 6885 17279 6919
rect 17221 6879 17279 6885
rect 17678 6876 17684 6928
rect 17736 6916 17742 6928
rect 17736 6888 18184 6916
rect 17736 6876 17742 6888
rect 11164 6820 11468 6848
rect 10965 6811 11023 6817
rect 11514 6808 11520 6860
rect 11572 6848 11578 6860
rect 12437 6851 12495 6857
rect 12437 6848 12449 6851
rect 11572 6820 12449 6848
rect 11572 6808 11578 6820
rect 12437 6817 12449 6820
rect 12483 6817 12495 6851
rect 12437 6811 12495 6817
rect 12526 6808 12532 6860
rect 12584 6848 12590 6860
rect 12621 6851 12679 6857
rect 12621 6848 12633 6851
rect 12584 6820 12633 6848
rect 12584 6808 12590 6820
rect 12621 6817 12633 6820
rect 12667 6817 12679 6851
rect 12621 6811 12679 6817
rect 13078 6808 13084 6860
rect 13136 6808 13142 6860
rect 13541 6851 13599 6857
rect 13541 6817 13553 6851
rect 13587 6817 13599 6851
rect 13541 6811 13599 6817
rect 13725 6851 13783 6857
rect 13725 6817 13737 6851
rect 13771 6848 13783 6851
rect 14182 6848 14188 6860
rect 13771 6820 14188 6848
rect 13771 6817 13783 6820
rect 13725 6811 13783 6817
rect 6730 6780 6736 6792
rect 6288 6752 6736 6780
rect 5445 6743 5503 6749
rect 6730 6740 6736 6752
rect 6788 6780 6794 6792
rect 7009 6783 7067 6789
rect 7009 6780 7021 6783
rect 6788 6752 7021 6780
rect 6788 6740 6794 6752
rect 7009 6749 7021 6752
rect 7055 6749 7067 6783
rect 7009 6743 7067 6749
rect 12158 6740 12164 6792
rect 12216 6780 12222 6792
rect 12342 6780 12348 6792
rect 12216 6752 12348 6780
rect 12216 6740 12222 6752
rect 12342 6740 12348 6752
rect 12400 6780 12406 6792
rect 13556 6780 13584 6811
rect 14182 6808 14188 6820
rect 14240 6808 14246 6860
rect 16666 6808 16672 6860
rect 16724 6808 16730 6860
rect 16761 6851 16819 6857
rect 16761 6817 16773 6851
rect 16807 6817 16819 6851
rect 16761 6811 16819 6817
rect 12400 6752 13584 6780
rect 16776 6780 16804 6811
rect 16942 6808 16948 6860
rect 17000 6808 17006 6860
rect 17034 6808 17040 6860
rect 17092 6808 17098 6860
rect 17313 6851 17371 6857
rect 17313 6817 17325 6851
rect 17359 6848 17371 6851
rect 17589 6851 17647 6857
rect 17359 6820 17540 6848
rect 17359 6817 17371 6820
rect 17313 6811 17371 6817
rect 17126 6780 17132 6792
rect 16776 6752 17132 6780
rect 12400 6740 12406 6752
rect 17126 6740 17132 6752
rect 17184 6780 17190 6792
rect 17405 6783 17463 6789
rect 17405 6780 17417 6783
rect 17184 6752 17417 6780
rect 17184 6740 17190 6752
rect 17405 6749 17417 6752
rect 17451 6749 17463 6783
rect 17512 6780 17540 6820
rect 17589 6817 17601 6851
rect 17635 6848 17647 6851
rect 17635 6820 17724 6848
rect 17635 6817 17647 6820
rect 17589 6811 17647 6817
rect 17696 6792 17724 6820
rect 17770 6808 17776 6860
rect 17828 6808 17834 6860
rect 17865 6851 17923 6857
rect 17865 6817 17877 6851
rect 17911 6848 17923 6851
rect 17954 6848 17960 6860
rect 17911 6820 17960 6848
rect 17911 6817 17923 6820
rect 17865 6811 17923 6817
rect 17954 6808 17960 6820
rect 18012 6808 18018 6860
rect 18156 6792 18184 6888
rect 19904 6888 20208 6916
rect 18414 6857 18420 6860
rect 18397 6851 18420 6857
rect 18397 6817 18409 6851
rect 18397 6811 18420 6817
rect 18414 6808 18420 6811
rect 18472 6808 18478 6860
rect 19797 6851 19855 6857
rect 19797 6817 19809 6851
rect 19843 6848 19855 6851
rect 19904 6848 19932 6888
rect 19843 6820 19932 6848
rect 19981 6851 20039 6857
rect 19843 6817 19855 6820
rect 19797 6811 19855 6817
rect 19981 6817 19993 6851
rect 20027 6848 20039 6851
rect 20073 6851 20131 6857
rect 20073 6848 20085 6851
rect 20027 6820 20085 6848
rect 20027 6817 20039 6820
rect 19981 6811 20039 6817
rect 20073 6817 20085 6820
rect 20119 6817 20131 6851
rect 20180 6848 20208 6888
rect 21174 6876 21180 6928
rect 21232 6916 21238 6928
rect 21361 6919 21419 6925
rect 21361 6916 21373 6919
rect 21232 6888 21373 6916
rect 21232 6876 21238 6888
rect 21361 6885 21373 6888
rect 21407 6916 21419 6919
rect 21450 6916 21456 6928
rect 21407 6888 21456 6916
rect 21407 6885 21419 6888
rect 21361 6879 21419 6885
rect 21450 6876 21456 6888
rect 21508 6876 21514 6928
rect 21577 6919 21635 6925
rect 21577 6885 21589 6919
rect 21623 6916 21635 6919
rect 22002 6916 22008 6928
rect 21623 6888 22008 6916
rect 21623 6885 21635 6888
rect 21577 6879 21635 6885
rect 22002 6876 22008 6888
rect 22060 6916 22066 6928
rect 25314 6916 25320 6928
rect 22060 6876 22094 6916
rect 20254 6848 20260 6860
rect 20180 6820 20260 6848
rect 20073 6811 20131 6817
rect 17512 6752 17632 6780
rect 17405 6743 17463 6749
rect 17604 6724 17632 6752
rect 17678 6740 17684 6792
rect 17736 6780 17742 6792
rect 18046 6780 18052 6792
rect 17736 6752 18052 6780
rect 17736 6740 17742 6752
rect 18046 6740 18052 6752
rect 18104 6740 18110 6792
rect 18138 6740 18144 6792
rect 18196 6740 18202 6792
rect 19996 6780 20024 6811
rect 20254 6808 20260 6820
rect 20312 6808 20318 6860
rect 22066 6848 22094 6876
rect 24596 6888 25320 6916
rect 23109 6851 23167 6857
rect 23109 6848 23121 6851
rect 22066 6820 23121 6848
rect 23109 6817 23121 6820
rect 23155 6817 23167 6851
rect 23109 6811 23167 6817
rect 23290 6808 23296 6860
rect 23348 6808 23354 6860
rect 23566 6808 23572 6860
rect 23624 6808 23630 6860
rect 23750 6808 23756 6860
rect 23808 6848 23814 6860
rect 24121 6851 24179 6857
rect 24121 6848 24133 6851
rect 23808 6820 24133 6848
rect 23808 6808 23814 6820
rect 24121 6817 24133 6820
rect 24167 6817 24179 6851
rect 24121 6811 24179 6817
rect 24213 6851 24271 6857
rect 24213 6817 24225 6851
rect 24259 6848 24271 6851
rect 24596 6848 24624 6888
rect 24259 6820 24624 6848
rect 24673 6851 24731 6857
rect 24259 6817 24271 6820
rect 24213 6811 24271 6817
rect 24673 6817 24685 6851
rect 24719 6817 24731 6851
rect 24673 6811 24731 6817
rect 19536 6752 20024 6780
rect 23584 6780 23612 6808
rect 24397 6783 24455 6789
rect 24397 6780 24409 6783
rect 23584 6752 24409 6780
rect 7834 6672 7840 6724
rect 7892 6712 7898 6724
rect 8021 6715 8079 6721
rect 8021 6712 8033 6715
rect 7892 6684 8033 6712
rect 7892 6672 7898 6684
rect 8021 6681 8033 6684
rect 8067 6681 8079 6715
rect 14642 6712 14648 6724
rect 8021 6675 8079 6681
rect 12268 6684 14648 6712
rect 3510 6604 3516 6656
rect 3568 6644 3574 6656
rect 4065 6647 4123 6653
rect 4065 6644 4077 6647
rect 3568 6616 4077 6644
rect 3568 6604 3574 6616
rect 4065 6613 4077 6616
rect 4111 6613 4123 6647
rect 4065 6607 4123 6613
rect 7653 6647 7711 6653
rect 7653 6613 7665 6647
rect 7699 6644 7711 6647
rect 7742 6644 7748 6656
rect 7699 6616 7748 6644
rect 7699 6613 7711 6616
rect 7653 6607 7711 6613
rect 7742 6604 7748 6616
rect 7800 6604 7806 6656
rect 9030 6604 9036 6656
rect 9088 6644 9094 6656
rect 12268 6644 12296 6684
rect 14642 6672 14648 6684
rect 14700 6672 14706 6724
rect 17586 6672 17592 6724
rect 17644 6672 17650 6724
rect 19536 6721 19564 6752
rect 24397 6749 24409 6752
rect 24443 6749 24455 6783
rect 24688 6780 24716 6811
rect 24762 6808 24768 6860
rect 24820 6808 24826 6860
rect 24857 6851 24915 6857
rect 24857 6817 24869 6851
rect 24903 6817 24915 6851
rect 24964 6848 24992 6888
rect 25314 6876 25320 6888
rect 25372 6916 25378 6928
rect 25372 6888 25544 6916
rect 25372 6876 25378 6888
rect 25041 6851 25099 6857
rect 25041 6848 25053 6851
rect 24964 6820 25053 6848
rect 24857 6811 24915 6817
rect 25041 6817 25053 6820
rect 25087 6817 25099 6851
rect 25041 6811 25099 6817
rect 24872 6780 24900 6811
rect 25130 6808 25136 6860
rect 25188 6808 25194 6860
rect 25222 6808 25228 6860
rect 25280 6808 25286 6860
rect 25406 6808 25412 6860
rect 25464 6808 25470 6860
rect 25516 6857 25544 6888
rect 25501 6851 25559 6857
rect 25501 6817 25513 6851
rect 25547 6817 25559 6851
rect 25608 6848 25636 6956
rect 26418 6944 26424 6996
rect 26476 6984 26482 6996
rect 26476 6956 26648 6984
rect 26476 6944 26482 6956
rect 26620 6925 26648 6956
rect 26605 6919 26663 6925
rect 26605 6885 26617 6919
rect 26651 6885 26663 6919
rect 26605 6879 26663 6885
rect 25777 6851 25835 6857
rect 25777 6848 25789 6851
rect 25608 6820 25789 6848
rect 25501 6811 25559 6817
rect 25777 6817 25789 6820
rect 25823 6817 25835 6851
rect 25777 6811 25835 6817
rect 25424 6780 25452 6808
rect 24688 6752 24808 6780
rect 24872 6752 25452 6780
rect 25792 6780 25820 6811
rect 25958 6808 25964 6860
rect 26016 6808 26022 6860
rect 26142 6808 26148 6860
rect 26200 6808 26206 6860
rect 26421 6851 26479 6857
rect 26421 6817 26433 6851
rect 26467 6817 26479 6851
rect 26421 6811 26479 6817
rect 26436 6780 26464 6811
rect 26786 6808 26792 6860
rect 26844 6808 26850 6860
rect 25792 6752 26464 6780
rect 24397 6743 24455 6749
rect 19521 6715 19579 6721
rect 19521 6681 19533 6715
rect 19567 6681 19579 6715
rect 22554 6712 22560 6724
rect 19521 6675 19579 6681
rect 21560 6684 22560 6712
rect 9088 6616 12296 6644
rect 9088 6604 9094 6616
rect 12342 6604 12348 6656
rect 12400 6604 12406 6656
rect 13262 6604 13268 6656
rect 13320 6604 13326 6656
rect 18049 6647 18107 6653
rect 18049 6613 18061 6647
rect 18095 6644 18107 6647
rect 18414 6644 18420 6656
rect 18095 6616 18420 6644
rect 18095 6613 18107 6616
rect 18049 6607 18107 6613
rect 18414 6604 18420 6616
rect 18472 6604 18478 6656
rect 21560 6653 21588 6684
rect 22554 6672 22560 6684
rect 22612 6672 22618 6724
rect 23014 6672 23020 6724
rect 23072 6672 23078 6724
rect 24780 6712 24808 6752
rect 25222 6712 25228 6724
rect 24780 6684 25228 6712
rect 25222 6672 25228 6684
rect 25280 6672 25286 6724
rect 21545 6647 21603 6653
rect 21545 6613 21557 6647
rect 21591 6613 21603 6647
rect 21545 6607 21603 6613
rect 21634 6604 21640 6656
rect 21692 6644 21698 6656
rect 21729 6647 21787 6653
rect 21729 6644 21741 6647
rect 21692 6616 21741 6644
rect 21692 6604 21698 6616
rect 21729 6613 21741 6616
rect 21775 6613 21787 6647
rect 21729 6607 21787 6613
rect 24762 6604 24768 6656
rect 24820 6644 24826 6656
rect 25130 6644 25136 6656
rect 24820 6616 25136 6644
rect 24820 6604 24826 6616
rect 25130 6604 25136 6616
rect 25188 6604 25194 6656
rect 25682 6604 25688 6656
rect 25740 6604 25746 6656
rect 552 6554 27416 6576
rect 552 6502 3756 6554
rect 3808 6502 3820 6554
rect 3872 6502 3884 6554
rect 3936 6502 3948 6554
rect 4000 6502 4012 6554
rect 4064 6502 10472 6554
rect 10524 6502 10536 6554
rect 10588 6502 10600 6554
rect 10652 6502 10664 6554
rect 10716 6502 10728 6554
rect 10780 6502 17188 6554
rect 17240 6502 17252 6554
rect 17304 6502 17316 6554
rect 17368 6502 17380 6554
rect 17432 6502 17444 6554
rect 17496 6502 23904 6554
rect 23956 6502 23968 6554
rect 24020 6502 24032 6554
rect 24084 6502 24096 6554
rect 24148 6502 24160 6554
rect 24212 6502 27416 6554
rect 552 6480 27416 6502
rect 2961 6443 3019 6449
rect 2961 6409 2973 6443
rect 3007 6440 3019 6443
rect 3881 6443 3939 6449
rect 3881 6440 3893 6443
rect 3007 6412 3893 6440
rect 3007 6409 3019 6412
rect 2961 6403 3019 6409
rect 3881 6409 3893 6412
rect 3927 6409 3939 6443
rect 3881 6403 3939 6409
rect 4614 6400 4620 6452
rect 4672 6440 4678 6452
rect 4709 6443 4767 6449
rect 4709 6440 4721 6443
rect 4672 6412 4721 6440
rect 4672 6400 4678 6412
rect 4709 6409 4721 6412
rect 4755 6409 4767 6443
rect 4709 6403 4767 6409
rect 5994 6400 6000 6452
rect 6052 6400 6058 6452
rect 7469 6443 7527 6449
rect 7469 6409 7481 6443
rect 7515 6440 7527 6443
rect 7745 6443 7803 6449
rect 7745 6440 7757 6443
rect 7515 6412 7757 6440
rect 7515 6409 7527 6412
rect 7469 6403 7527 6409
rect 7745 6409 7757 6412
rect 7791 6409 7803 6443
rect 7745 6403 7803 6409
rect 9125 6443 9183 6449
rect 9125 6409 9137 6443
rect 9171 6440 9183 6443
rect 9401 6443 9459 6449
rect 9401 6440 9413 6443
rect 9171 6412 9413 6440
rect 9171 6409 9183 6412
rect 9125 6403 9183 6409
rect 9401 6409 9413 6412
rect 9447 6409 9459 6443
rect 9401 6403 9459 6409
rect 9950 6400 9956 6452
rect 10008 6440 10014 6452
rect 11514 6440 11520 6452
rect 10008 6412 11520 6440
rect 10008 6400 10014 6412
rect 11514 6400 11520 6412
rect 11572 6400 11578 6452
rect 12084 6412 12388 6440
rect 3602 6332 3608 6384
rect 3660 6332 3666 6384
rect 5258 6372 5264 6384
rect 4724 6344 5264 6372
rect 2884 6276 3464 6304
rect 2884 6245 2912 6276
rect 3436 6245 3464 6276
rect 4724 6248 4752 6344
rect 5258 6332 5264 6344
rect 5316 6332 5322 6384
rect 9214 6332 9220 6384
rect 9272 6372 9278 6384
rect 9309 6375 9367 6381
rect 9309 6372 9321 6375
rect 9272 6344 9321 6372
rect 9272 6332 9278 6344
rect 9309 6341 9321 6344
rect 9355 6341 9367 6375
rect 10318 6372 10324 6384
rect 9309 6335 9367 6341
rect 9600 6344 10324 6372
rect 5074 6304 5080 6316
rect 4816 6276 5080 6304
rect 2869 6239 2927 6245
rect 2869 6205 2881 6239
rect 2915 6205 2927 6239
rect 3053 6239 3111 6245
rect 3053 6236 3065 6239
rect 2869 6199 2927 6205
rect 2976 6208 3065 6236
rect 2976 6180 3004 6208
rect 3053 6205 3065 6208
rect 3099 6236 3111 6239
rect 3237 6239 3295 6245
rect 3237 6236 3249 6239
rect 3099 6208 3249 6236
rect 3099 6205 3111 6208
rect 3053 6199 3111 6205
rect 3237 6205 3249 6208
rect 3283 6205 3295 6239
rect 3237 6199 3295 6205
rect 3421 6239 3479 6245
rect 3421 6205 3433 6239
rect 3467 6236 3479 6239
rect 3510 6236 3516 6248
rect 3467 6208 3516 6236
rect 3467 6205 3479 6208
rect 3421 6199 3479 6205
rect 3510 6196 3516 6208
rect 3568 6196 3574 6248
rect 4341 6239 4399 6245
rect 4341 6205 4353 6239
rect 4387 6236 4399 6239
rect 4522 6236 4528 6248
rect 4387 6208 4528 6236
rect 4387 6205 4399 6208
rect 4341 6199 4399 6205
rect 4522 6196 4528 6208
rect 4580 6196 4586 6248
rect 4617 6239 4675 6245
rect 4617 6205 4629 6239
rect 4663 6236 4675 6239
rect 4706 6236 4712 6248
rect 4663 6208 4712 6236
rect 4663 6205 4675 6208
rect 4617 6199 4675 6205
rect 4706 6196 4712 6208
rect 4764 6196 4770 6248
rect 4816 6245 4844 6276
rect 5074 6264 5080 6276
rect 5132 6264 5138 6316
rect 6822 6304 6828 6316
rect 5920 6276 6828 6304
rect 4801 6239 4859 6245
rect 4801 6205 4813 6239
rect 4847 6205 4859 6239
rect 4801 6199 4859 6205
rect 4890 6196 4896 6248
rect 4948 6196 4954 6248
rect 5626 6196 5632 6248
rect 5684 6236 5690 6248
rect 5920 6245 5948 6276
rect 6822 6264 6828 6276
rect 6880 6264 6886 6316
rect 5905 6239 5963 6245
rect 5905 6236 5917 6239
rect 5684 6208 5917 6236
rect 5684 6196 5690 6208
rect 5905 6205 5917 6208
rect 5951 6205 5963 6239
rect 5905 6199 5963 6205
rect 6089 6239 6147 6245
rect 6089 6205 6101 6239
rect 6135 6205 6147 6239
rect 6089 6199 6147 6205
rect 2958 6128 2964 6180
rect 3016 6128 3022 6180
rect 3602 6128 3608 6180
rect 3660 6168 3666 6180
rect 3849 6171 3907 6177
rect 3849 6168 3861 6171
rect 3660 6140 3861 6168
rect 3660 6128 3666 6140
rect 3849 6137 3861 6140
rect 3895 6137 3907 6171
rect 3849 6131 3907 6137
rect 4062 6128 4068 6180
rect 4120 6128 4126 6180
rect 6104 6168 6132 6199
rect 6178 6196 6184 6248
rect 6236 6236 6242 6248
rect 6365 6239 6423 6245
rect 6365 6236 6377 6239
rect 6236 6208 6377 6236
rect 6236 6196 6242 6208
rect 6365 6205 6377 6208
rect 6411 6205 6423 6239
rect 6365 6199 6423 6205
rect 7101 6239 7159 6245
rect 7101 6205 7113 6239
rect 7147 6236 7159 6239
rect 7466 6236 7472 6248
rect 7147 6208 7472 6236
rect 7147 6205 7159 6208
rect 7101 6199 7159 6205
rect 7466 6196 7472 6208
rect 7524 6196 7530 6248
rect 8110 6196 8116 6248
rect 8168 6236 8174 6248
rect 9030 6236 9036 6248
rect 8168 6208 9036 6236
rect 8168 6196 8174 6208
rect 6546 6168 6552 6180
rect 6104 6140 6552 6168
rect 6546 6128 6552 6140
rect 6604 6128 6610 6180
rect 7006 6128 7012 6180
rect 7064 6168 7070 6180
rect 7285 6171 7343 6177
rect 7285 6168 7297 6171
rect 7064 6140 7297 6168
rect 7064 6128 7070 6140
rect 7285 6137 7297 6140
rect 7331 6137 7343 6171
rect 7285 6131 7343 6137
rect 7561 6171 7619 6177
rect 7561 6137 7573 6171
rect 7607 6168 7619 6171
rect 8662 6168 8668 6180
rect 7607 6140 8668 6168
rect 7607 6137 7619 6140
rect 7561 6131 7619 6137
rect 3694 6060 3700 6112
rect 3752 6060 3758 6112
rect 4080 6100 4108 6128
rect 7576 6100 7604 6131
rect 8662 6128 8668 6140
rect 8720 6128 8726 6180
rect 8956 6177 8984 6208
rect 9030 6196 9036 6208
rect 9088 6196 9094 6248
rect 9600 6245 9628 6344
rect 10318 6332 10324 6344
rect 10376 6332 10382 6384
rect 11977 6375 12035 6381
rect 11977 6372 11989 6375
rect 10612 6344 11989 6372
rect 9692 6276 10088 6304
rect 9692 6245 9720 6276
rect 10060 6248 10088 6276
rect 9585 6239 9643 6245
rect 9585 6205 9597 6239
rect 9631 6205 9643 6239
rect 9585 6199 9643 6205
rect 9677 6239 9735 6245
rect 9677 6205 9689 6239
rect 9723 6205 9735 6239
rect 9677 6199 9735 6205
rect 9858 6196 9864 6248
rect 9916 6196 9922 6248
rect 9950 6196 9956 6248
rect 10008 6196 10014 6248
rect 10042 6196 10048 6248
rect 10100 6196 10106 6248
rect 10336 6245 10364 6332
rect 10321 6239 10379 6245
rect 10321 6205 10333 6239
rect 10367 6236 10379 6239
rect 10502 6236 10508 6248
rect 10367 6208 10508 6236
rect 10367 6205 10379 6208
rect 10321 6199 10379 6205
rect 10502 6196 10508 6208
rect 10560 6196 10566 6248
rect 10612 6245 10640 6344
rect 11977 6341 11989 6344
rect 12023 6341 12035 6375
rect 11977 6335 12035 6341
rect 12084 6304 12112 6412
rect 12360 6384 12388 6412
rect 12526 6400 12532 6452
rect 12584 6400 12590 6452
rect 16209 6443 16267 6449
rect 16209 6409 16221 6443
rect 16255 6440 16267 6443
rect 16298 6440 16304 6452
rect 16255 6412 16304 6440
rect 16255 6409 16267 6412
rect 16209 6403 16267 6409
rect 16298 6400 16304 6412
rect 16356 6400 16362 6452
rect 23290 6400 23296 6452
rect 23348 6440 23354 6452
rect 23569 6443 23627 6449
rect 23569 6440 23581 6443
rect 23348 6412 23581 6440
rect 23348 6400 23354 6412
rect 23569 6409 23581 6412
rect 23615 6409 23627 6443
rect 23569 6403 23627 6409
rect 24394 6400 24400 6452
rect 24452 6400 24458 6452
rect 24578 6400 24584 6452
rect 24636 6400 24642 6452
rect 25314 6400 25320 6452
rect 25372 6400 25378 6452
rect 25406 6400 25412 6452
rect 25464 6440 25470 6452
rect 25777 6443 25835 6449
rect 25777 6440 25789 6443
rect 25464 6412 25789 6440
rect 25464 6400 25470 6412
rect 25777 6409 25789 6412
rect 25823 6409 25835 6443
rect 25777 6403 25835 6409
rect 12342 6332 12348 6384
rect 12400 6372 12406 6384
rect 12544 6372 12572 6400
rect 12400 6332 12434 6372
rect 12544 6344 12664 6372
rect 11716 6276 12112 6304
rect 12406 6304 12434 6332
rect 12406 6276 12572 6304
rect 10597 6239 10655 6245
rect 10597 6205 10609 6239
rect 10643 6205 10655 6239
rect 10597 6199 10655 6205
rect 10873 6239 10931 6245
rect 10873 6205 10885 6239
rect 10919 6236 10931 6239
rect 11514 6236 11520 6248
rect 10919 6208 11520 6236
rect 10919 6205 10931 6208
rect 10873 6199 10931 6205
rect 8941 6171 8999 6177
rect 8941 6137 8953 6171
rect 8987 6137 8999 6171
rect 8941 6131 8999 6137
rect 9157 6171 9215 6177
rect 9157 6137 9169 6171
rect 9203 6168 9215 6171
rect 9398 6168 9404 6180
rect 9203 6140 9404 6168
rect 9203 6137 9215 6140
rect 9157 6131 9215 6137
rect 9398 6128 9404 6140
rect 9456 6168 9462 6180
rect 10137 6171 10195 6177
rect 10137 6168 10149 6171
rect 9456 6140 10149 6168
rect 9456 6128 9462 6140
rect 10137 6137 10149 6140
rect 10183 6137 10195 6171
rect 10137 6131 10195 6137
rect 4080 6072 7604 6100
rect 7742 6060 7748 6112
rect 7800 6109 7806 6112
rect 7800 6103 7819 6109
rect 7807 6069 7819 6103
rect 7800 6063 7819 6069
rect 7800 6060 7806 6063
rect 7926 6060 7932 6112
rect 7984 6060 7990 6112
rect 9858 6060 9864 6112
rect 9916 6100 9922 6112
rect 10612 6100 10640 6199
rect 11514 6196 11520 6208
rect 11572 6196 11578 6248
rect 11716 6245 11744 6276
rect 11701 6239 11759 6245
rect 11701 6205 11713 6239
rect 11747 6205 11759 6239
rect 11701 6199 11759 6205
rect 11790 6196 11796 6248
rect 11848 6196 11854 6248
rect 12250 6196 12256 6248
rect 12308 6196 12314 6248
rect 12342 6196 12348 6248
rect 12400 6196 12406 6248
rect 12544 6245 12572 6276
rect 12529 6239 12587 6245
rect 12529 6205 12541 6239
rect 12575 6205 12587 6239
rect 12529 6199 12587 6205
rect 11977 6171 12035 6177
rect 11977 6137 11989 6171
rect 12023 6168 12035 6171
rect 12636 6168 12664 6344
rect 15746 6332 15752 6384
rect 15804 6332 15810 6384
rect 13262 6264 13268 6316
rect 13320 6304 13326 6316
rect 14921 6307 14979 6313
rect 13320 6276 13952 6304
rect 13320 6264 13326 6276
rect 13170 6196 13176 6248
rect 13228 6196 13234 6248
rect 13357 6239 13415 6245
rect 13357 6205 13369 6239
rect 13403 6236 13415 6239
rect 13924 6236 13952 6276
rect 14921 6273 14933 6307
rect 14967 6304 14979 6307
rect 15764 6304 15792 6332
rect 14967 6276 15792 6304
rect 14967 6273 14979 6276
rect 14921 6267 14979 6273
rect 21266 6264 21272 6316
rect 21324 6304 21330 6316
rect 21729 6307 21787 6313
rect 21729 6304 21741 6307
rect 21324 6276 21741 6304
rect 21324 6264 21330 6276
rect 21729 6273 21741 6276
rect 21775 6273 21787 6307
rect 21729 6267 21787 6273
rect 23566 6264 23572 6316
rect 23624 6304 23630 6316
rect 24029 6307 24087 6313
rect 24029 6304 24041 6307
rect 23624 6276 24041 6304
rect 23624 6264 23630 6276
rect 24029 6273 24041 6276
rect 24075 6273 24087 6307
rect 25958 6304 25964 6316
rect 24029 6267 24087 6273
rect 25240 6276 25964 6304
rect 14654 6239 14712 6245
rect 14654 6236 14666 6239
rect 13403 6208 13584 6236
rect 13924 6208 14666 6236
rect 13403 6205 13415 6208
rect 13357 6199 13415 6205
rect 12023 6140 12664 6168
rect 12023 6137 12035 6140
rect 11977 6131 12035 6137
rect 13556 6112 13584 6208
rect 14654 6205 14666 6208
rect 14700 6205 14712 6239
rect 15565 6239 15623 6245
rect 15565 6236 15577 6239
rect 14654 6199 14712 6205
rect 15304 6208 15577 6236
rect 15304 6180 15332 6208
rect 15565 6205 15577 6208
rect 15611 6205 15623 6239
rect 15565 6199 15623 6205
rect 15749 6239 15807 6245
rect 15749 6205 15761 6239
rect 15795 6205 15807 6239
rect 15749 6199 15807 6205
rect 15286 6128 15292 6180
rect 15344 6128 15350 6180
rect 15470 6128 15476 6180
rect 15528 6168 15534 6180
rect 15764 6168 15792 6199
rect 16574 6196 16580 6248
rect 16632 6236 16638 6248
rect 17034 6236 17040 6248
rect 16632 6208 17040 6236
rect 16632 6196 16638 6208
rect 17034 6196 17040 6208
rect 17092 6196 17098 6248
rect 17126 6196 17132 6248
rect 17184 6236 17190 6248
rect 17221 6239 17279 6245
rect 17221 6236 17233 6239
rect 17184 6208 17233 6236
rect 17184 6196 17190 6208
rect 17221 6205 17233 6208
rect 17267 6205 17279 6239
rect 17221 6199 17279 6205
rect 17405 6239 17463 6245
rect 17405 6205 17417 6239
rect 17451 6236 17463 6239
rect 17862 6236 17868 6248
rect 17451 6208 17868 6236
rect 17451 6205 17463 6208
rect 17405 6199 17463 6205
rect 15528 6140 15792 6168
rect 17236 6168 17264 6199
rect 17862 6196 17868 6208
rect 17920 6196 17926 6248
rect 21453 6239 21511 6245
rect 21453 6205 21465 6239
rect 21499 6236 21511 6239
rect 21634 6236 21640 6248
rect 21499 6208 21640 6236
rect 21499 6205 21511 6208
rect 21453 6199 21511 6205
rect 21634 6196 21640 6208
rect 21692 6196 21698 6248
rect 22922 6196 22928 6248
rect 22980 6236 22986 6248
rect 23385 6239 23443 6245
rect 23385 6236 23397 6239
rect 22980 6208 23397 6236
rect 22980 6196 22986 6208
rect 23385 6205 23397 6208
rect 23431 6205 23443 6239
rect 23385 6199 23443 6205
rect 25130 6196 25136 6248
rect 25188 6236 25194 6248
rect 25240 6245 25268 6276
rect 25958 6264 25964 6276
rect 26016 6264 26022 6316
rect 25225 6239 25283 6245
rect 25225 6236 25237 6239
rect 25188 6208 25237 6236
rect 25188 6196 25194 6208
rect 25225 6205 25237 6208
rect 25271 6205 25283 6239
rect 25225 6199 25283 6205
rect 25409 6239 25467 6245
rect 25409 6205 25421 6239
rect 25455 6236 25467 6239
rect 26050 6236 26056 6248
rect 25455 6208 26056 6236
rect 25455 6205 25467 6208
rect 25409 6199 25467 6205
rect 26050 6196 26056 6208
rect 26108 6236 26114 6248
rect 26145 6239 26203 6245
rect 26145 6236 26157 6239
rect 26108 6208 26157 6236
rect 26108 6196 26114 6208
rect 26145 6205 26157 6208
rect 26191 6205 26203 6239
rect 26145 6199 26203 6205
rect 17770 6168 17776 6180
rect 17236 6140 17776 6168
rect 15528 6128 15534 6140
rect 17770 6128 17776 6140
rect 17828 6128 17834 6180
rect 21974 6171 22032 6177
rect 21974 6168 21986 6171
rect 21652 6140 21986 6168
rect 9916 6072 10640 6100
rect 9916 6060 9922 6072
rect 12158 6060 12164 6112
rect 12216 6100 12222 6112
rect 13173 6103 13231 6109
rect 13173 6100 13185 6103
rect 12216 6072 13185 6100
rect 12216 6060 12222 6072
rect 13173 6069 13185 6072
rect 13219 6069 13231 6103
rect 13173 6063 13231 6069
rect 13538 6060 13544 6112
rect 13596 6060 13602 6112
rect 15105 6103 15163 6109
rect 15105 6069 15117 6103
rect 15151 6100 15163 6103
rect 15194 6100 15200 6112
rect 15151 6072 15200 6100
rect 15151 6069 15163 6072
rect 15105 6063 15163 6069
rect 15194 6060 15200 6072
rect 15252 6060 15258 6112
rect 15562 6060 15568 6112
rect 15620 6060 15626 6112
rect 16022 6060 16028 6112
rect 16080 6060 16086 6112
rect 16209 6103 16267 6109
rect 16209 6069 16221 6103
rect 16255 6100 16267 6103
rect 16482 6100 16488 6112
rect 16255 6072 16488 6100
rect 16255 6069 16267 6072
rect 16209 6063 16267 6069
rect 16482 6060 16488 6072
rect 16540 6060 16546 6112
rect 17218 6060 17224 6112
rect 17276 6100 17282 6112
rect 17586 6100 17592 6112
rect 17276 6072 17592 6100
rect 17276 6060 17282 6072
rect 17586 6060 17592 6072
rect 17644 6060 17650 6112
rect 21652 6109 21680 6140
rect 21974 6137 21986 6140
rect 22020 6137 22032 6171
rect 21974 6131 22032 6137
rect 23201 6171 23259 6177
rect 23201 6137 23213 6171
rect 23247 6137 23259 6171
rect 23201 6131 23259 6137
rect 24397 6171 24455 6177
rect 24397 6137 24409 6171
rect 24443 6168 24455 6171
rect 25682 6168 25688 6180
rect 24443 6140 25688 6168
rect 24443 6137 24455 6140
rect 24397 6131 24455 6137
rect 21637 6103 21695 6109
rect 21637 6069 21649 6103
rect 21683 6069 21695 6103
rect 21637 6063 21695 6069
rect 23106 6060 23112 6112
rect 23164 6100 23170 6112
rect 23216 6100 23244 6131
rect 25682 6128 25688 6140
rect 25740 6128 25746 6180
rect 25958 6128 25964 6180
rect 26016 6128 26022 6180
rect 23164 6072 23244 6100
rect 23164 6060 23170 6072
rect 552 6010 27576 6032
rect 552 5958 7114 6010
rect 7166 5958 7178 6010
rect 7230 5958 7242 6010
rect 7294 5958 7306 6010
rect 7358 5958 7370 6010
rect 7422 5958 13830 6010
rect 13882 5958 13894 6010
rect 13946 5958 13958 6010
rect 14010 5958 14022 6010
rect 14074 5958 14086 6010
rect 14138 5958 20546 6010
rect 20598 5958 20610 6010
rect 20662 5958 20674 6010
rect 20726 5958 20738 6010
rect 20790 5958 20802 6010
rect 20854 5958 27262 6010
rect 27314 5958 27326 6010
rect 27378 5958 27390 6010
rect 27442 5958 27454 6010
rect 27506 5958 27518 6010
rect 27570 5958 27576 6010
rect 552 5936 27576 5958
rect 3418 5856 3424 5908
rect 3476 5896 3482 5908
rect 3513 5899 3571 5905
rect 3513 5896 3525 5899
rect 3476 5868 3525 5896
rect 3476 5856 3482 5868
rect 3513 5865 3525 5868
rect 3559 5865 3571 5899
rect 3513 5859 3571 5865
rect 4890 5856 4896 5908
rect 4948 5856 4954 5908
rect 5626 5856 5632 5908
rect 5684 5856 5690 5908
rect 9953 5899 10011 5905
rect 9953 5865 9965 5899
rect 9999 5865 10011 5899
rect 9953 5859 10011 5865
rect 3694 5828 3700 5840
rect 2608 5800 3700 5828
rect 2608 5769 2636 5800
rect 3694 5788 3700 5800
rect 3752 5788 3758 5840
rect 4908 5828 4936 5856
rect 9306 5828 9312 5840
rect 4632 5800 4936 5828
rect 8588 5800 9312 5828
rect 2593 5763 2651 5769
rect 2593 5729 2605 5763
rect 2639 5729 2651 5763
rect 2593 5723 2651 5729
rect 3050 5720 3056 5772
rect 3108 5720 3114 5772
rect 3237 5763 3295 5769
rect 3237 5729 3249 5763
rect 3283 5760 3295 5763
rect 4154 5760 4160 5772
rect 3283 5732 4160 5760
rect 3283 5729 3295 5732
rect 3237 5723 3295 5729
rect 4154 5720 4160 5732
rect 4212 5720 4218 5772
rect 4246 5720 4252 5772
rect 4304 5720 4310 5772
rect 4522 5720 4528 5772
rect 4580 5720 4586 5772
rect 4632 5769 4660 5800
rect 4617 5763 4675 5769
rect 4617 5729 4629 5763
rect 4663 5729 4675 5763
rect 4617 5723 4675 5729
rect 4890 5720 4896 5772
rect 4948 5720 4954 5772
rect 5997 5763 6055 5769
rect 5997 5729 6009 5763
rect 6043 5760 6055 5763
rect 6178 5760 6184 5772
rect 6043 5732 6184 5760
rect 6043 5729 6055 5732
rect 5997 5723 6055 5729
rect 6178 5720 6184 5732
rect 6236 5720 6242 5772
rect 6270 5720 6276 5772
rect 6328 5720 6334 5772
rect 8202 5720 8208 5772
rect 8260 5769 8266 5772
rect 8588 5769 8616 5800
rect 9306 5788 9312 5800
rect 9364 5788 9370 5840
rect 9968 5828 9996 5859
rect 10042 5856 10048 5908
rect 10100 5856 10106 5908
rect 10502 5856 10508 5908
rect 10560 5856 10566 5908
rect 11790 5856 11796 5908
rect 11848 5896 11854 5908
rect 12342 5896 12348 5908
rect 11848 5868 12348 5896
rect 11848 5856 11854 5868
rect 12342 5856 12348 5868
rect 12400 5856 12406 5908
rect 13170 5856 13176 5908
rect 13228 5896 13234 5908
rect 13228 5868 14044 5896
rect 13228 5856 13234 5868
rect 10413 5831 10471 5837
rect 10413 5828 10425 5831
rect 9968 5800 10425 5828
rect 10413 5797 10425 5800
rect 10459 5828 10471 5831
rect 10459 5800 10732 5828
rect 10459 5797 10471 5800
rect 10413 5791 10471 5797
rect 8846 5769 8852 5772
rect 8260 5723 8272 5769
rect 8481 5763 8539 5769
rect 8481 5729 8493 5763
rect 8527 5760 8539 5763
rect 8573 5763 8631 5769
rect 8573 5760 8585 5763
rect 8527 5732 8585 5760
rect 8527 5729 8539 5732
rect 8481 5723 8539 5729
rect 8573 5729 8585 5732
rect 8619 5729 8631 5763
rect 8573 5723 8631 5729
rect 8840 5723 8852 5769
rect 8260 5720 8266 5723
rect 8846 5720 8852 5723
rect 8904 5720 8910 5772
rect 10134 5720 10140 5772
rect 10192 5760 10198 5772
rect 10704 5769 10732 5800
rect 13538 5788 13544 5840
rect 13596 5828 13602 5840
rect 14016 5837 14044 5868
rect 14182 5856 14188 5908
rect 14240 5856 14246 5908
rect 14369 5899 14427 5905
rect 14369 5865 14381 5899
rect 14415 5896 14427 5899
rect 15470 5896 15476 5908
rect 14415 5868 15476 5896
rect 14415 5865 14427 5868
rect 14369 5859 14427 5865
rect 15470 5856 15476 5868
rect 15528 5856 15534 5908
rect 16482 5856 16488 5908
rect 16540 5856 16546 5908
rect 17129 5899 17187 5905
rect 17129 5896 17141 5899
rect 16592 5868 17141 5896
rect 13817 5831 13875 5837
rect 13817 5828 13829 5831
rect 13596 5800 13829 5828
rect 13596 5788 13602 5800
rect 13817 5797 13829 5800
rect 13863 5797 13875 5831
rect 13817 5791 13875 5797
rect 14001 5831 14059 5837
rect 14001 5797 14013 5831
rect 14047 5828 14059 5831
rect 14550 5828 14556 5840
rect 14047 5800 14556 5828
rect 14047 5797 14059 5800
rect 14001 5791 14059 5797
rect 14550 5788 14556 5800
rect 14608 5788 14614 5840
rect 15562 5788 15568 5840
rect 15620 5828 15626 5840
rect 16592 5828 16620 5868
rect 17129 5865 17141 5868
rect 17175 5896 17187 5899
rect 21269 5899 21327 5905
rect 17175 5868 17540 5896
rect 17175 5865 17187 5868
rect 17129 5859 17187 5865
rect 17218 5828 17224 5840
rect 15620 5800 16620 5828
rect 16684 5800 17224 5828
rect 15620 5788 15626 5800
rect 10229 5763 10287 5769
rect 10229 5760 10241 5763
rect 10192 5732 10241 5760
rect 10192 5720 10198 5732
rect 10229 5729 10241 5732
rect 10275 5760 10287 5763
rect 10505 5763 10563 5769
rect 10505 5760 10517 5763
rect 10275 5732 10517 5760
rect 10275 5729 10287 5732
rect 10229 5723 10287 5729
rect 10505 5729 10517 5732
rect 10551 5729 10563 5763
rect 10505 5723 10563 5729
rect 10689 5763 10747 5769
rect 10689 5729 10701 5763
rect 10735 5729 10747 5763
rect 10689 5723 10747 5729
rect 15470 5720 15476 5772
rect 15528 5769 15534 5772
rect 15528 5723 15540 5769
rect 15528 5720 15534 5723
rect 16022 5720 16028 5772
rect 16080 5760 16086 5772
rect 16684 5769 16712 5800
rect 17218 5788 17224 5800
rect 17276 5828 17282 5840
rect 17405 5831 17463 5837
rect 17405 5828 17417 5831
rect 17276 5800 17417 5828
rect 17276 5788 17282 5800
rect 17405 5797 17417 5800
rect 17451 5797 17463 5831
rect 17405 5791 17463 5797
rect 16209 5763 16267 5769
rect 16209 5760 16221 5763
rect 16080 5732 16221 5760
rect 16080 5720 16086 5732
rect 16209 5729 16221 5732
rect 16255 5729 16267 5763
rect 16209 5723 16267 5729
rect 16669 5763 16727 5769
rect 16669 5729 16681 5763
rect 16715 5729 16727 5763
rect 16669 5723 16727 5729
rect 15746 5652 15752 5704
rect 15804 5652 15810 5704
rect 16761 5695 16819 5701
rect 16761 5661 16773 5695
rect 16807 5661 16819 5695
rect 17512 5692 17540 5868
rect 21269 5865 21281 5899
rect 21315 5865 21327 5899
rect 21269 5859 21327 5865
rect 21437 5899 21495 5905
rect 21437 5865 21449 5899
rect 21483 5896 21495 5899
rect 21818 5896 21824 5908
rect 21483 5868 21824 5896
rect 21483 5865 21495 5868
rect 21437 5859 21495 5865
rect 17770 5788 17776 5840
rect 17828 5788 17834 5840
rect 17862 5788 17868 5840
rect 17920 5788 17926 5840
rect 17788 5760 17816 5788
rect 18049 5763 18107 5769
rect 18049 5760 18061 5763
rect 17788 5732 18061 5760
rect 18049 5729 18061 5732
rect 18095 5729 18107 5763
rect 18049 5723 18107 5729
rect 19978 5720 19984 5772
rect 20036 5720 20042 5772
rect 21085 5763 21143 5769
rect 21085 5729 21097 5763
rect 21131 5760 21143 5763
rect 21284 5760 21312 5859
rect 21818 5856 21824 5868
rect 21876 5856 21882 5908
rect 23014 5856 23020 5908
rect 23072 5856 23078 5908
rect 25041 5899 25099 5905
rect 25041 5865 25053 5899
rect 25087 5896 25099 5899
rect 25222 5896 25228 5908
rect 25087 5868 25228 5896
rect 25087 5865 25099 5868
rect 25041 5859 25099 5865
rect 25222 5856 25228 5868
rect 25280 5856 25286 5908
rect 21542 5788 21548 5840
rect 21600 5828 21606 5840
rect 21637 5831 21695 5837
rect 21637 5828 21649 5831
rect 21600 5800 21649 5828
rect 21600 5788 21606 5800
rect 21637 5797 21649 5800
rect 21683 5797 21695 5831
rect 21910 5828 21916 5840
rect 21637 5791 21695 5797
rect 21836 5800 21916 5828
rect 21131 5732 21312 5760
rect 21131 5729 21143 5732
rect 21085 5723 21143 5729
rect 21726 5720 21732 5772
rect 21784 5720 21790 5772
rect 17773 5695 17831 5701
rect 17773 5692 17785 5695
rect 17512 5664 17785 5692
rect 16761 5655 16819 5661
rect 17773 5661 17785 5664
rect 17819 5661 17831 5695
rect 17773 5655 17831 5661
rect 7006 5584 7012 5636
rect 7064 5624 7070 5636
rect 7190 5624 7196 5636
rect 7064 5596 7196 5624
rect 7064 5584 7070 5596
rect 7190 5584 7196 5596
rect 7248 5584 7254 5636
rect 16776 5624 16804 5655
rect 19702 5652 19708 5704
rect 19760 5652 19766 5704
rect 21836 5692 21864 5800
rect 21910 5788 21916 5800
rect 21968 5788 21974 5840
rect 24670 5788 24676 5840
rect 24728 5828 24734 5840
rect 24728 5800 25176 5828
rect 24728 5788 24734 5800
rect 22922 5720 22928 5772
rect 22980 5720 22986 5772
rect 23106 5720 23112 5772
rect 23164 5720 23170 5772
rect 25148 5769 25176 5800
rect 25133 5763 25191 5769
rect 25133 5729 25145 5763
rect 25179 5729 25191 5763
rect 25133 5723 25191 5729
rect 20732 5664 21864 5692
rect 25148 5692 25176 5723
rect 25222 5720 25228 5772
rect 25280 5720 25286 5772
rect 25406 5720 25412 5772
rect 25464 5760 25470 5772
rect 25501 5763 25559 5769
rect 25501 5760 25513 5763
rect 25464 5732 25513 5760
rect 25464 5720 25470 5732
rect 25501 5729 25513 5732
rect 25547 5729 25559 5763
rect 25501 5723 25559 5729
rect 25682 5720 25688 5772
rect 25740 5720 25746 5772
rect 25593 5695 25651 5701
rect 25593 5692 25605 5695
rect 25148 5664 25605 5692
rect 16776 5596 17448 5624
rect 1118 5516 1124 5568
rect 1176 5556 1182 5568
rect 1213 5559 1271 5565
rect 1213 5556 1225 5559
rect 1176 5528 1225 5556
rect 1176 5516 1182 5528
rect 1213 5525 1225 5528
rect 1259 5525 1271 5559
rect 1213 5519 1271 5525
rect 2406 5516 2412 5568
rect 2464 5516 2470 5568
rect 3142 5516 3148 5568
rect 3200 5516 3206 5568
rect 7101 5559 7159 5565
rect 7101 5525 7113 5559
rect 7147 5556 7159 5559
rect 7466 5556 7472 5568
rect 7147 5528 7472 5556
rect 7147 5525 7159 5528
rect 7101 5519 7159 5525
rect 7466 5516 7472 5528
rect 7524 5516 7530 5568
rect 12437 5559 12495 5565
rect 12437 5525 12449 5559
rect 12483 5556 12495 5559
rect 12526 5556 12532 5568
rect 12483 5528 12532 5556
rect 12483 5525 12495 5528
rect 12437 5519 12495 5525
rect 12526 5516 12532 5528
rect 12584 5516 12590 5568
rect 16298 5516 16304 5568
rect 16356 5556 16362 5568
rect 16393 5559 16451 5565
rect 16393 5556 16405 5559
rect 16356 5528 16405 5556
rect 16356 5516 16362 5528
rect 16393 5525 16405 5528
rect 16439 5525 16451 5559
rect 16393 5519 16451 5525
rect 16574 5516 16580 5568
rect 16632 5556 16638 5568
rect 17420 5565 17448 5596
rect 17954 5584 17960 5636
rect 18012 5624 18018 5636
rect 20732 5633 20760 5664
rect 25593 5661 25605 5664
rect 25639 5661 25651 5695
rect 25593 5655 25651 5661
rect 18325 5627 18383 5633
rect 18325 5624 18337 5627
rect 18012 5596 18337 5624
rect 18012 5584 18018 5596
rect 18325 5593 18337 5596
rect 18371 5593 18383 5627
rect 18325 5587 18383 5593
rect 20717 5627 20775 5633
rect 20717 5593 20729 5627
rect 20763 5593 20775 5627
rect 20717 5587 20775 5593
rect 24302 5584 24308 5636
rect 24360 5584 24366 5636
rect 17221 5559 17279 5565
rect 17221 5556 17233 5559
rect 16632 5528 17233 5556
rect 16632 5516 16638 5528
rect 17221 5525 17233 5528
rect 17267 5525 17279 5559
rect 17221 5519 17279 5525
rect 17405 5559 17463 5565
rect 17405 5525 17417 5559
rect 17451 5556 17463 5559
rect 18233 5559 18291 5565
rect 18233 5556 18245 5559
rect 17451 5528 18245 5556
rect 17451 5525 17463 5528
rect 17405 5519 17463 5525
rect 18233 5525 18245 5528
rect 18279 5525 18291 5559
rect 18233 5519 18291 5525
rect 18874 5516 18880 5568
rect 18932 5556 18938 5568
rect 18969 5559 19027 5565
rect 18969 5556 18981 5559
rect 18932 5528 18981 5556
rect 18932 5516 18938 5528
rect 18969 5525 18981 5528
rect 19015 5525 19027 5559
rect 18969 5519 19027 5525
rect 19334 5516 19340 5568
rect 19392 5516 19398 5568
rect 20898 5516 20904 5568
rect 20956 5516 20962 5568
rect 21453 5559 21511 5565
rect 21453 5525 21465 5559
rect 21499 5556 21511 5559
rect 22097 5559 22155 5565
rect 22097 5556 22109 5559
rect 21499 5528 22109 5556
rect 21499 5525 21511 5528
rect 21453 5519 21511 5525
rect 22097 5525 22109 5528
rect 22143 5525 22155 5559
rect 22097 5519 22155 5525
rect 22554 5516 22560 5568
rect 22612 5516 22618 5568
rect 24578 5516 24584 5568
rect 24636 5556 24642 5568
rect 24673 5559 24731 5565
rect 24673 5556 24685 5559
rect 24636 5528 24685 5556
rect 24636 5516 24642 5528
rect 24673 5525 24685 5528
rect 24719 5525 24731 5559
rect 24673 5519 24731 5525
rect 24762 5516 24768 5568
rect 24820 5556 24826 5568
rect 24857 5559 24915 5565
rect 24857 5556 24869 5559
rect 24820 5528 24869 5556
rect 24820 5516 24826 5528
rect 24857 5525 24869 5528
rect 24903 5525 24915 5559
rect 24857 5519 24915 5525
rect 25314 5516 25320 5568
rect 25372 5556 25378 5568
rect 25409 5559 25467 5565
rect 25409 5556 25421 5559
rect 25372 5528 25421 5556
rect 25372 5516 25378 5528
rect 25409 5525 25421 5528
rect 25455 5525 25467 5559
rect 25409 5519 25467 5525
rect 552 5466 27416 5488
rect 552 5414 3756 5466
rect 3808 5414 3820 5466
rect 3872 5414 3884 5466
rect 3936 5414 3948 5466
rect 4000 5414 4012 5466
rect 4064 5414 10472 5466
rect 10524 5414 10536 5466
rect 10588 5414 10600 5466
rect 10652 5414 10664 5466
rect 10716 5414 10728 5466
rect 10780 5414 17188 5466
rect 17240 5414 17252 5466
rect 17304 5414 17316 5466
rect 17368 5414 17380 5466
rect 17432 5414 17444 5466
rect 17496 5414 23904 5466
rect 23956 5414 23968 5466
rect 24020 5414 24032 5466
rect 24084 5414 24096 5466
rect 24148 5414 24160 5466
rect 24212 5414 27416 5466
rect 552 5392 27416 5414
rect 3050 5312 3056 5364
rect 3108 5312 3114 5364
rect 4246 5312 4252 5364
rect 4304 5352 4310 5364
rect 5445 5355 5503 5361
rect 5445 5352 5457 5355
rect 4304 5324 5457 5352
rect 4304 5312 4310 5324
rect 5445 5321 5457 5324
rect 5491 5321 5503 5355
rect 5445 5315 5503 5321
rect 6270 5312 6276 5364
rect 6328 5312 6334 5364
rect 6454 5312 6460 5364
rect 6512 5352 6518 5364
rect 7561 5355 7619 5361
rect 6512 5324 7144 5352
rect 6512 5312 6518 5324
rect 4798 5244 4804 5296
rect 4856 5284 4862 5296
rect 5169 5287 5227 5293
rect 5169 5284 5181 5287
rect 4856 5256 5181 5284
rect 4856 5244 4862 5256
rect 5169 5253 5181 5256
rect 5215 5253 5227 5287
rect 6914 5284 6920 5296
rect 5169 5247 5227 5253
rect 5276 5256 6920 5284
rect 1670 5176 1676 5228
rect 1728 5176 1734 5228
rect 5276 5160 5304 5256
rect 6086 5176 6092 5228
rect 6144 5216 6150 5228
rect 6656 5225 6684 5256
rect 6914 5244 6920 5256
rect 6972 5244 6978 5296
rect 7116 5284 7144 5324
rect 7561 5321 7573 5355
rect 7607 5352 7619 5355
rect 7742 5352 7748 5364
rect 7607 5324 7748 5352
rect 7607 5321 7619 5324
rect 7561 5315 7619 5321
rect 7742 5312 7748 5324
rect 7800 5312 7806 5364
rect 8021 5355 8079 5361
rect 8021 5321 8033 5355
rect 8067 5352 8079 5355
rect 8202 5352 8208 5364
rect 8067 5324 8208 5352
rect 8067 5321 8079 5324
rect 8021 5315 8079 5321
rect 8202 5312 8208 5324
rect 8260 5312 8266 5364
rect 8846 5312 8852 5364
rect 8904 5352 8910 5364
rect 9033 5355 9091 5361
rect 9033 5352 9045 5355
rect 8904 5324 9045 5352
rect 8904 5312 8910 5324
rect 9033 5321 9045 5324
rect 9079 5321 9091 5355
rect 9033 5315 9091 5321
rect 11609 5355 11667 5361
rect 11609 5321 11621 5355
rect 11655 5352 11667 5355
rect 11790 5352 11796 5364
rect 11655 5324 11796 5352
rect 11655 5321 11667 5324
rect 11609 5315 11667 5321
rect 11790 5312 11796 5324
rect 11848 5312 11854 5364
rect 14550 5312 14556 5364
rect 14608 5312 14614 5364
rect 15194 5312 15200 5364
rect 15252 5352 15258 5364
rect 15289 5355 15347 5361
rect 15289 5352 15301 5355
rect 15252 5324 15301 5352
rect 15252 5312 15258 5324
rect 15289 5321 15301 5324
rect 15335 5321 15347 5355
rect 15289 5315 15347 5321
rect 15470 5312 15476 5364
rect 15528 5352 15534 5364
rect 15565 5355 15623 5361
rect 15565 5352 15577 5355
rect 15528 5324 15577 5352
rect 15528 5312 15534 5324
rect 15565 5321 15577 5324
rect 15611 5321 15623 5355
rect 15565 5315 15623 5321
rect 15746 5312 15752 5364
rect 15804 5352 15810 5364
rect 18138 5352 18144 5364
rect 15804 5324 18144 5352
rect 15804 5312 15810 5324
rect 7834 5284 7840 5296
rect 7116 5256 7840 5284
rect 6457 5219 6515 5225
rect 6457 5216 6469 5219
rect 6144 5188 6469 5216
rect 6144 5176 6150 5188
rect 6457 5185 6469 5188
rect 6503 5185 6515 5219
rect 6457 5179 6515 5185
rect 6641 5219 6699 5225
rect 6641 5185 6653 5219
rect 6687 5185 6699 5219
rect 6641 5179 6699 5185
rect 6733 5219 6791 5225
rect 6733 5185 6745 5219
rect 6779 5216 6791 5219
rect 7009 5219 7067 5225
rect 7009 5216 7021 5219
rect 6779 5188 7021 5216
rect 6779 5185 6791 5188
rect 6733 5179 6791 5185
rect 7009 5185 7021 5188
rect 7055 5185 7067 5219
rect 7009 5179 7067 5185
rect 1581 5151 1639 5157
rect 1581 5117 1593 5151
rect 1627 5117 1639 5151
rect 1581 5111 1639 5117
rect 1940 5151 1998 5157
rect 1940 5117 1952 5151
rect 1986 5148 1998 5151
rect 2406 5148 2412 5160
rect 1986 5120 2412 5148
rect 1986 5117 1998 5120
rect 1940 5111 1998 5117
rect 1596 5080 1624 5111
rect 2406 5108 2412 5120
rect 2464 5108 2470 5160
rect 3050 5108 3056 5160
rect 3108 5148 3114 5160
rect 3237 5151 3295 5157
rect 3237 5148 3249 5151
rect 3108 5120 3249 5148
rect 3108 5108 3114 5120
rect 3237 5117 3249 5120
rect 3283 5117 3295 5151
rect 3237 5111 3295 5117
rect 4065 5151 4123 5157
rect 4065 5117 4077 5151
rect 4111 5148 4123 5151
rect 4157 5151 4215 5157
rect 4157 5148 4169 5151
rect 4111 5120 4169 5148
rect 4111 5117 4123 5120
rect 4065 5111 4123 5117
rect 4157 5117 4169 5120
rect 4203 5117 4215 5151
rect 4157 5111 4215 5117
rect 4433 5151 4491 5157
rect 4433 5117 4445 5151
rect 4479 5148 4491 5151
rect 4982 5148 4988 5160
rect 4479 5120 4988 5148
rect 4479 5117 4491 5120
rect 4433 5111 4491 5117
rect 4982 5108 4988 5120
rect 5040 5108 5046 5160
rect 5258 5108 5264 5160
rect 5316 5108 5322 5160
rect 5445 5151 5503 5157
rect 5445 5117 5457 5151
rect 5491 5117 5503 5151
rect 5445 5111 5503 5117
rect 3326 5080 3332 5092
rect 1596 5052 3332 5080
rect 3326 5040 3332 5052
rect 3384 5040 3390 5092
rect 3421 5083 3479 5089
rect 3421 5049 3433 5083
rect 3467 5080 3479 5083
rect 4246 5080 4252 5092
rect 3467 5052 4252 5080
rect 3467 5049 3479 5052
rect 3421 5043 3479 5049
rect 4246 5040 4252 5052
rect 4304 5040 4310 5092
rect 1394 4972 1400 5024
rect 1452 4972 1458 5024
rect 3602 4972 3608 5024
rect 3660 4972 3666 5024
rect 5460 5012 5488 5111
rect 5902 5108 5908 5160
rect 5960 5150 5966 5160
rect 5997 5153 6055 5159
rect 5997 5150 6009 5153
rect 5960 5122 6009 5150
rect 5960 5108 5966 5122
rect 5997 5119 6009 5122
rect 6043 5119 6055 5153
rect 5997 5113 6055 5119
rect 6178 5108 6184 5160
rect 6236 5108 6242 5160
rect 7116 5157 7144 5256
rect 7834 5244 7840 5256
rect 7892 5284 7898 5296
rect 8294 5284 8300 5296
rect 7892 5256 8300 5284
rect 7892 5244 7898 5256
rect 8294 5244 8300 5256
rect 8352 5244 8358 5296
rect 11882 5244 11888 5296
rect 11940 5284 11946 5296
rect 12342 5284 12348 5296
rect 11940 5256 12348 5284
rect 11940 5244 11946 5256
rect 12342 5244 12348 5256
rect 12400 5244 12406 5296
rect 7190 5176 7196 5228
rect 7248 5216 7254 5228
rect 15562 5216 15568 5228
rect 7248 5188 7696 5216
rect 7248 5176 7254 5188
rect 6549 5151 6607 5157
rect 6549 5117 6561 5151
rect 6595 5117 6607 5151
rect 6549 5111 6607 5117
rect 6917 5151 6975 5157
rect 6917 5117 6929 5151
rect 6963 5117 6975 5151
rect 6917 5111 6975 5117
rect 7101 5151 7159 5157
rect 7101 5117 7113 5151
rect 7147 5117 7159 5151
rect 7101 5111 7159 5117
rect 6564 5080 6592 5111
rect 6932 5080 6960 5111
rect 7466 5108 7472 5160
rect 7524 5108 7530 5160
rect 7668 5157 7696 5188
rect 15350 5188 15568 5216
rect 7653 5151 7711 5157
rect 7653 5117 7665 5151
rect 7699 5117 7711 5151
rect 7653 5111 7711 5117
rect 7837 5151 7895 5157
rect 7837 5117 7849 5151
rect 7883 5148 7895 5151
rect 7926 5148 7932 5160
rect 7883 5120 7932 5148
rect 7883 5117 7895 5120
rect 7837 5111 7895 5117
rect 7926 5108 7932 5120
rect 7984 5108 7990 5160
rect 9214 5108 9220 5160
rect 9272 5108 9278 5160
rect 10505 5151 10563 5157
rect 10505 5117 10517 5151
rect 10551 5148 10563 5151
rect 10597 5151 10655 5157
rect 10597 5148 10609 5151
rect 10551 5120 10609 5148
rect 10551 5117 10563 5120
rect 10505 5111 10563 5117
rect 10597 5117 10609 5120
rect 10643 5117 10655 5151
rect 10597 5111 10655 5117
rect 10778 5108 10784 5160
rect 10836 5148 10842 5160
rect 10873 5151 10931 5157
rect 10873 5148 10885 5151
rect 10836 5120 10885 5148
rect 10836 5108 10842 5120
rect 10873 5117 10885 5120
rect 10919 5117 10931 5151
rect 10873 5111 10931 5117
rect 11885 5151 11943 5157
rect 11885 5117 11897 5151
rect 11931 5148 11943 5151
rect 11974 5148 11980 5160
rect 11931 5120 11980 5148
rect 11931 5117 11943 5120
rect 11885 5111 11943 5117
rect 11974 5108 11980 5120
rect 12032 5108 12038 5160
rect 12345 5151 12403 5157
rect 12345 5117 12357 5151
rect 12391 5148 12403 5151
rect 12526 5148 12532 5160
rect 12391 5120 12532 5148
rect 12391 5117 12403 5120
rect 12345 5111 12403 5117
rect 12526 5108 12532 5120
rect 12584 5108 12590 5160
rect 12618 5108 12624 5160
rect 12676 5108 12682 5160
rect 12710 5108 12716 5160
rect 12768 5108 12774 5160
rect 13446 5108 13452 5160
rect 13504 5148 13510 5160
rect 13541 5151 13599 5157
rect 13541 5148 13553 5151
rect 13504 5120 13553 5148
rect 13504 5108 13510 5120
rect 13541 5117 13553 5120
rect 13587 5117 13599 5151
rect 13541 5111 13599 5117
rect 13722 5108 13728 5160
rect 13780 5148 13786 5160
rect 13817 5151 13875 5157
rect 13817 5148 13829 5151
rect 13780 5120 13829 5148
rect 13780 5108 13786 5120
rect 13817 5117 13829 5120
rect 13863 5117 13875 5151
rect 13817 5111 13875 5117
rect 7006 5080 7012 5092
rect 6564 5052 7012 5080
rect 7006 5040 7012 5052
rect 7064 5080 7070 5092
rect 7558 5080 7564 5092
rect 7064 5052 7564 5080
rect 7064 5040 7070 5052
rect 7558 5040 7564 5052
rect 7616 5040 7622 5092
rect 11330 5040 11336 5092
rect 11388 5080 11394 5092
rect 12069 5083 12127 5089
rect 12069 5080 12081 5083
rect 11388 5052 12081 5080
rect 11388 5040 11394 5052
rect 12069 5049 12081 5052
rect 12115 5080 12127 5083
rect 12728 5080 12756 5108
rect 12115 5052 12756 5080
rect 12115 5049 12127 5052
rect 12069 5043 12127 5049
rect 14642 5040 14648 5092
rect 14700 5080 14706 5092
rect 15350 5089 15378 5188
rect 15562 5176 15568 5188
rect 15620 5176 15626 5228
rect 16224 5225 16252 5324
rect 18138 5312 18144 5324
rect 18196 5352 18202 5364
rect 21637 5355 21695 5361
rect 18196 5324 20300 5352
rect 18196 5312 18202 5324
rect 17589 5287 17647 5293
rect 17589 5253 17601 5287
rect 17635 5284 17647 5287
rect 17862 5284 17868 5296
rect 17635 5256 17868 5284
rect 17635 5253 17647 5256
rect 17589 5247 17647 5253
rect 17862 5244 17868 5256
rect 17920 5244 17926 5296
rect 19702 5244 19708 5296
rect 19760 5284 19766 5296
rect 19981 5287 20039 5293
rect 19981 5284 19993 5287
rect 19760 5256 19993 5284
rect 19760 5244 19766 5256
rect 19981 5253 19993 5256
rect 20027 5253 20039 5287
rect 19981 5247 20039 5253
rect 16209 5219 16267 5225
rect 16209 5185 16221 5219
rect 16255 5185 16267 5219
rect 18322 5216 18328 5228
rect 16209 5179 16267 5185
rect 17972 5188 18328 5216
rect 15749 5151 15807 5157
rect 15749 5148 15761 5151
rect 15488 5120 15761 5148
rect 15105 5083 15163 5089
rect 15105 5080 15117 5083
rect 14700 5052 15117 5080
rect 14700 5040 14706 5052
rect 15105 5049 15117 5052
rect 15151 5049 15163 5083
rect 15105 5043 15163 5049
rect 15321 5083 15379 5089
rect 15321 5049 15333 5083
rect 15367 5049 15379 5083
rect 15321 5043 15379 5049
rect 6178 5012 6184 5024
rect 5460 4984 6184 5012
rect 6178 4972 6184 4984
rect 6236 4972 6242 5024
rect 12253 5015 12311 5021
rect 12253 4981 12265 5015
rect 12299 5012 12311 5015
rect 12710 5012 12716 5024
rect 12299 4984 12716 5012
rect 12299 4981 12311 4984
rect 12253 4975 12311 4981
rect 12710 4972 12716 4984
rect 12768 4972 12774 5024
rect 13357 5015 13415 5021
rect 13357 4981 13369 5015
rect 13403 5012 13415 5015
rect 15194 5012 15200 5024
rect 13403 4984 15200 5012
rect 13403 4981 13415 4984
rect 13357 4975 13415 4981
rect 15194 4972 15200 4984
rect 15252 4972 15258 5024
rect 15488 5021 15516 5120
rect 15749 5117 15761 5120
rect 15795 5117 15807 5151
rect 15749 5111 15807 5117
rect 16298 5108 16304 5160
rect 16356 5148 16362 5160
rect 17972 5157 18000 5188
rect 18322 5176 18328 5188
rect 18380 5176 18386 5228
rect 18874 5176 18880 5228
rect 18932 5176 18938 5228
rect 20272 5225 20300 5324
rect 21637 5321 21649 5355
rect 21683 5352 21695 5355
rect 21726 5352 21732 5364
rect 21683 5324 21732 5352
rect 21683 5321 21695 5324
rect 21637 5315 21695 5321
rect 21726 5312 21732 5324
rect 21784 5312 21790 5364
rect 21818 5312 21824 5364
rect 21876 5352 21882 5364
rect 24302 5352 24308 5364
rect 21876 5324 24308 5352
rect 21876 5312 21882 5324
rect 23569 5287 23627 5293
rect 23569 5253 23581 5287
rect 23615 5284 23627 5287
rect 23658 5284 23664 5296
rect 23615 5256 23664 5284
rect 23615 5253 23627 5256
rect 23569 5247 23627 5253
rect 23658 5244 23664 5256
rect 23716 5244 23722 5296
rect 20257 5219 20315 5225
rect 20257 5185 20269 5219
rect 20303 5185 20315 5219
rect 20257 5179 20315 5185
rect 22554 5176 22560 5228
rect 22612 5176 22618 5228
rect 24228 5225 24256 5324
rect 24302 5312 24308 5324
rect 24360 5312 24366 5364
rect 24213 5219 24271 5225
rect 24213 5185 24225 5219
rect 24259 5185 24271 5219
rect 24213 5179 24271 5185
rect 24670 5176 24676 5228
rect 24728 5176 24734 5228
rect 25038 5176 25044 5228
rect 25096 5176 25102 5228
rect 16465 5151 16523 5157
rect 16465 5148 16477 5151
rect 16356 5120 16477 5148
rect 16356 5108 16362 5120
rect 16465 5117 16477 5120
rect 16511 5117 16523 5151
rect 16465 5111 16523 5117
rect 17957 5151 18015 5157
rect 17957 5117 17969 5151
rect 18003 5117 18015 5151
rect 17957 5111 18015 5117
rect 18138 5108 18144 5160
rect 18196 5108 18202 5160
rect 19150 5108 19156 5160
rect 19208 5108 19214 5160
rect 20524 5151 20582 5157
rect 20524 5117 20536 5151
rect 20570 5148 20582 5151
rect 20898 5148 20904 5160
rect 20570 5120 20904 5148
rect 20570 5117 20582 5120
rect 20524 5111 20582 5117
rect 20898 5108 20904 5120
rect 20956 5108 20962 5160
rect 21726 5108 21732 5160
rect 21784 5108 21790 5160
rect 21910 5108 21916 5160
rect 21968 5108 21974 5160
rect 22094 5108 22100 5160
rect 22152 5148 22158 5160
rect 22189 5151 22247 5157
rect 22189 5148 22201 5151
rect 22152 5120 22201 5148
rect 22152 5108 22158 5120
rect 22189 5117 22201 5120
rect 22235 5117 22247 5151
rect 22189 5111 22247 5117
rect 22833 5151 22891 5157
rect 22833 5117 22845 5151
rect 22879 5148 22891 5151
rect 23198 5148 23204 5160
rect 22879 5120 23204 5148
rect 22879 5117 22891 5120
rect 22833 5111 22891 5117
rect 23198 5108 23204 5120
rect 23256 5108 23262 5160
rect 24578 5108 24584 5160
rect 24636 5108 24642 5160
rect 25314 5157 25320 5160
rect 25308 5148 25320 5157
rect 25275 5120 25320 5148
rect 25308 5111 25320 5120
rect 25314 5108 25320 5111
rect 25372 5108 25378 5160
rect 15473 5015 15531 5021
rect 15473 4981 15485 5015
rect 15519 4981 15531 5015
rect 15473 4975 15531 4981
rect 18046 4972 18052 5024
rect 18104 4972 18110 5024
rect 19886 4972 19892 5024
rect 19944 4972 19950 5024
rect 24394 4972 24400 5024
rect 24452 5012 24458 5024
rect 24857 5015 24915 5021
rect 24857 5012 24869 5015
rect 24452 4984 24869 5012
rect 24452 4972 24458 4984
rect 24857 4981 24869 4984
rect 24903 4981 24915 5015
rect 24857 4975 24915 4981
rect 25682 4972 25688 5024
rect 25740 5012 25746 5024
rect 26421 5015 26479 5021
rect 26421 5012 26433 5015
rect 25740 4984 26433 5012
rect 25740 4972 25746 4984
rect 26421 4981 26433 4984
rect 26467 4981 26479 5015
rect 26421 4975 26479 4981
rect 552 4922 27576 4944
rect 552 4870 7114 4922
rect 7166 4870 7178 4922
rect 7230 4870 7242 4922
rect 7294 4870 7306 4922
rect 7358 4870 7370 4922
rect 7422 4870 13830 4922
rect 13882 4870 13894 4922
rect 13946 4870 13958 4922
rect 14010 4870 14022 4922
rect 14074 4870 14086 4922
rect 14138 4870 20546 4922
rect 20598 4870 20610 4922
rect 20662 4870 20674 4922
rect 20726 4870 20738 4922
rect 20790 4870 20802 4922
rect 20854 4870 27262 4922
rect 27314 4870 27326 4922
rect 27378 4870 27390 4922
rect 27442 4870 27454 4922
rect 27506 4870 27518 4922
rect 27570 4870 27576 4922
rect 552 4848 27576 4870
rect 2130 4768 2136 4820
rect 2188 4768 2194 4820
rect 2958 4768 2964 4820
rect 3016 4768 3022 4820
rect 3326 4768 3332 4820
rect 3384 4808 3390 4820
rect 3384 4780 4292 4808
rect 3384 4768 3390 4780
rect 3602 4740 3608 4752
rect 2976 4712 3608 4740
rect 1118 4632 1124 4684
rect 1176 4632 1182 4684
rect 1394 4632 1400 4684
rect 1452 4632 1458 4684
rect 2976 4681 3004 4712
rect 3602 4700 3608 4712
rect 3660 4700 3666 4752
rect 4264 4740 4292 4780
rect 4890 4768 4896 4820
rect 4948 4768 4954 4820
rect 4982 4768 4988 4820
rect 5040 4768 5046 4820
rect 5813 4811 5871 4817
rect 5813 4777 5825 4811
rect 5859 4777 5871 4811
rect 5813 4771 5871 4777
rect 5828 4740 5856 4771
rect 5902 4768 5908 4820
rect 5960 4808 5966 4820
rect 7742 4808 7748 4820
rect 5960 4780 7748 4808
rect 5960 4768 5966 4780
rect 4264 4712 5856 4740
rect 5994 4700 6000 4752
rect 6052 4700 6058 4752
rect 6454 4740 6460 4752
rect 6380 4712 6460 4740
rect 2961 4675 3019 4681
rect 2961 4641 2973 4675
rect 3007 4641 3019 4675
rect 2961 4635 3019 4641
rect 3142 4632 3148 4684
rect 3200 4632 3206 4684
rect 4706 4632 4712 4684
rect 4764 4632 4770 4684
rect 5166 4632 5172 4684
rect 5224 4632 5230 4684
rect 6380 4681 6408 4712
rect 6454 4700 6460 4712
rect 6512 4700 6518 4752
rect 6656 4749 6684 4780
rect 7742 4768 7748 4780
rect 7800 4808 7806 4820
rect 8294 4808 8300 4820
rect 7800 4780 8300 4808
rect 7800 4768 7806 4780
rect 8294 4768 8300 4780
rect 8352 4768 8358 4820
rect 8389 4811 8447 4817
rect 8389 4777 8401 4811
rect 8435 4808 8447 4811
rect 8570 4808 8576 4820
rect 8435 4780 8576 4808
rect 8435 4777 8447 4780
rect 8389 4771 8447 4777
rect 8570 4768 8576 4780
rect 8628 4768 8634 4820
rect 10778 4768 10784 4820
rect 10836 4768 10842 4820
rect 12161 4811 12219 4817
rect 12161 4777 12173 4811
rect 12207 4808 12219 4811
rect 12618 4808 12624 4820
rect 12207 4780 12624 4808
rect 12207 4777 12219 4780
rect 12161 4771 12219 4777
rect 12618 4768 12624 4780
rect 12676 4768 12682 4820
rect 13357 4811 13415 4817
rect 13357 4777 13369 4811
rect 13403 4808 13415 4811
rect 13722 4808 13728 4820
rect 13403 4780 13728 4808
rect 13403 4777 13415 4780
rect 13357 4771 13415 4777
rect 13722 4768 13728 4780
rect 13780 4768 13786 4820
rect 14826 4768 14832 4820
rect 14884 4808 14890 4820
rect 15197 4811 15255 4817
rect 15197 4808 15209 4811
rect 14884 4780 15209 4808
rect 14884 4768 14890 4780
rect 15197 4777 15209 4780
rect 15243 4777 15255 4811
rect 15197 4771 15255 4777
rect 18690 4768 18696 4820
rect 18748 4808 18754 4820
rect 18785 4811 18843 4817
rect 18785 4808 18797 4811
rect 18748 4780 18797 4808
rect 18748 4768 18754 4780
rect 18785 4777 18797 4780
rect 18831 4777 18843 4811
rect 18785 4771 18843 4777
rect 19150 4768 19156 4820
rect 19208 4768 19214 4820
rect 20254 4768 20260 4820
rect 20312 4768 20318 4820
rect 22005 4811 22063 4817
rect 22005 4777 22017 4811
rect 22051 4777 22063 4811
rect 22005 4771 22063 4777
rect 6641 4743 6699 4749
rect 6641 4709 6653 4743
rect 6687 4709 6699 4743
rect 11882 4740 11888 4752
rect 6641 4703 6699 4709
rect 7392 4712 8524 4740
rect 7392 4681 7420 4712
rect 6365 4675 6423 4681
rect 6365 4641 6377 4675
rect 6411 4641 6423 4675
rect 6365 4635 6423 4641
rect 6825 4675 6883 4681
rect 6825 4641 6837 4675
rect 6871 4672 6883 4675
rect 7101 4675 7159 4681
rect 7101 4672 7113 4675
rect 6871 4644 7113 4672
rect 6871 4641 6883 4644
rect 6825 4635 6883 4641
rect 7101 4641 7113 4644
rect 7147 4641 7159 4675
rect 7101 4635 7159 4641
rect 7377 4675 7435 4681
rect 7377 4641 7389 4675
rect 7423 4641 7435 4675
rect 7377 4635 7435 4641
rect 7558 4632 7564 4684
rect 7616 4672 7622 4684
rect 8496 4681 8524 4712
rect 11348 4712 11888 4740
rect 7653 4675 7711 4681
rect 7653 4672 7665 4675
rect 7616 4644 7665 4672
rect 7616 4632 7622 4644
rect 7653 4641 7665 4644
rect 7699 4641 7711 4675
rect 7653 4635 7711 4641
rect 8481 4675 8539 4681
rect 8481 4641 8493 4675
rect 8527 4641 8539 4675
rect 8481 4635 8539 4641
rect 10597 4675 10655 4681
rect 10597 4641 10609 4675
rect 10643 4641 10655 4675
rect 10597 4635 10655 4641
rect 11057 4675 11115 4681
rect 11057 4641 11069 4675
rect 11103 4672 11115 4675
rect 11146 4672 11152 4684
rect 11103 4644 11152 4672
rect 11103 4641 11115 4644
rect 11057 4635 11115 4641
rect 6914 4496 6920 4548
rect 6972 4536 6978 4548
rect 7098 4536 7104 4548
rect 6972 4508 7104 4536
rect 6972 4496 6978 4508
rect 7098 4496 7104 4508
rect 7156 4496 7162 4548
rect 10612 4536 10640 4635
rect 11146 4632 11152 4644
rect 11204 4632 11210 4684
rect 11238 4632 11244 4684
rect 11296 4632 11302 4684
rect 11348 4681 11376 4712
rect 11882 4700 11888 4712
rect 11940 4700 11946 4752
rect 11974 4700 11980 4752
rect 12032 4740 12038 4752
rect 12345 4743 12403 4749
rect 12345 4740 12357 4743
rect 12032 4712 12357 4740
rect 12032 4700 12038 4712
rect 12345 4709 12357 4712
rect 12391 4709 12403 4743
rect 12345 4703 12403 4709
rect 12710 4700 12716 4752
rect 12768 4700 12774 4752
rect 19334 4700 19340 4752
rect 19392 4700 19398 4752
rect 22020 4740 22048 4771
rect 22922 4768 22928 4820
rect 22980 4808 22986 4820
rect 23109 4811 23167 4817
rect 23109 4808 23121 4811
rect 22980 4780 23121 4808
rect 22980 4768 22986 4780
rect 23109 4777 23121 4780
rect 23155 4777 23167 4811
rect 23109 4771 23167 4777
rect 23198 4768 23204 4820
rect 23256 4768 23262 4820
rect 24394 4768 24400 4820
rect 24452 4768 24458 4820
rect 24578 4768 24584 4820
rect 24636 4808 24642 4820
rect 25133 4811 25191 4817
rect 25133 4808 25145 4811
rect 24636 4780 25145 4808
rect 24636 4768 24642 4780
rect 25133 4777 25145 4780
rect 25179 4777 25191 4811
rect 25133 4771 25191 4777
rect 25317 4743 25375 4749
rect 22020 4712 22094 4740
rect 11333 4675 11391 4681
rect 11333 4641 11345 4675
rect 11379 4641 11391 4675
rect 11333 4635 11391 4641
rect 11514 4632 11520 4684
rect 11572 4672 11578 4684
rect 12529 4675 12587 4681
rect 12529 4672 12541 4675
rect 11572 4644 12541 4672
rect 11572 4632 11578 4644
rect 12529 4641 12541 4644
rect 12575 4641 12587 4675
rect 12529 4635 12587 4641
rect 13170 4632 13176 4684
rect 13228 4632 13234 4684
rect 13446 4632 13452 4684
rect 13504 4632 13510 4684
rect 14458 4632 14464 4684
rect 14516 4632 14522 4684
rect 17773 4675 17831 4681
rect 17773 4641 17785 4675
rect 17819 4672 17831 4675
rect 17954 4672 17960 4684
rect 17819 4644 17960 4672
rect 17819 4641 17831 4644
rect 17773 4635 17831 4641
rect 17954 4632 17960 4644
rect 18012 4632 18018 4684
rect 18046 4632 18052 4684
rect 18104 4632 18110 4684
rect 18966 4632 18972 4684
rect 19024 4632 19030 4684
rect 19245 4675 19303 4681
rect 19245 4641 19257 4675
rect 19291 4672 19303 4675
rect 19352 4672 19380 4700
rect 19291 4644 19380 4672
rect 19521 4675 19579 4681
rect 19291 4641 19303 4644
rect 19245 4635 19303 4641
rect 19521 4641 19533 4675
rect 19567 4672 19579 4675
rect 20714 4672 20720 4684
rect 19567 4644 20720 4672
rect 19567 4641 19579 4644
rect 19521 4635 19579 4641
rect 20714 4632 20720 4644
rect 20772 4632 20778 4684
rect 21818 4632 21824 4684
rect 21876 4632 21882 4684
rect 22066 4672 22094 4712
rect 25317 4709 25329 4743
rect 25363 4740 25375 4743
rect 25406 4740 25412 4752
rect 25363 4712 25412 4740
rect 25363 4709 25375 4712
rect 25317 4703 25375 4709
rect 25406 4700 25412 4712
rect 25464 4700 25470 4752
rect 25501 4743 25559 4749
rect 25501 4709 25513 4743
rect 25547 4740 25559 4743
rect 25682 4740 25688 4752
rect 25547 4712 25688 4740
rect 25547 4709 25559 4712
rect 25501 4703 25559 4709
rect 25682 4700 25688 4712
rect 25740 4700 25746 4752
rect 22373 4675 22431 4681
rect 22373 4672 22385 4675
rect 22066 4644 22385 4672
rect 22373 4641 22385 4644
rect 22419 4641 22431 4675
rect 22373 4635 22431 4641
rect 23382 4632 23388 4684
rect 23440 4632 23446 4684
rect 24029 4675 24087 4681
rect 24029 4641 24041 4675
rect 24075 4672 24087 4675
rect 24762 4672 24768 4684
rect 24075 4644 24768 4672
rect 24075 4641 24087 4644
rect 24029 4635 24087 4641
rect 24762 4632 24768 4644
rect 24820 4632 24826 4684
rect 11425 4607 11483 4613
rect 11425 4573 11437 4607
rect 11471 4604 11483 4607
rect 11701 4607 11759 4613
rect 11701 4604 11713 4607
rect 11471 4576 11713 4604
rect 11471 4573 11483 4576
rect 11425 4567 11483 4573
rect 11701 4573 11713 4576
rect 11747 4573 11759 4607
rect 11701 4567 11759 4573
rect 11790 4564 11796 4616
rect 11848 4564 11854 4616
rect 11882 4564 11888 4616
rect 11940 4564 11946 4616
rect 11977 4607 12035 4613
rect 11977 4573 11989 4607
rect 12023 4573 12035 4607
rect 11977 4567 12035 4573
rect 14093 4607 14151 4613
rect 14093 4573 14105 4607
rect 14139 4604 14151 4607
rect 14185 4607 14243 4613
rect 14185 4604 14197 4607
rect 14139 4576 14197 4604
rect 14139 4573 14151 4576
rect 14093 4567 14151 4573
rect 14185 4573 14197 4576
rect 14231 4573 14243 4607
rect 14185 4567 14243 4573
rect 11054 4536 11060 4548
rect 10612 4508 11060 4536
rect 11054 4496 11060 4508
rect 11112 4496 11118 4548
rect 11149 4539 11207 4545
rect 11149 4505 11161 4539
rect 11195 4536 11207 4539
rect 11238 4536 11244 4548
rect 11195 4508 11244 4536
rect 11195 4505 11207 4508
rect 11149 4499 11207 4505
rect 11238 4496 11244 4508
rect 11296 4536 11302 4548
rect 11992 4536 12020 4567
rect 22094 4564 22100 4616
rect 22152 4564 22158 4616
rect 11296 4508 12020 4536
rect 11296 4496 11302 4508
rect 12342 4496 12348 4548
rect 12400 4536 12406 4548
rect 12897 4539 12955 4545
rect 12897 4536 12909 4539
rect 12400 4508 12909 4536
rect 12400 4496 12406 4508
rect 12897 4505 12909 4508
rect 12943 4505 12955 4539
rect 12897 4499 12955 4505
rect 24581 4539 24639 4545
rect 24581 4505 24593 4539
rect 24627 4536 24639 4539
rect 25222 4536 25228 4548
rect 24627 4508 25228 4536
rect 24627 4505 24639 4508
rect 24581 4499 24639 4505
rect 25222 4496 25228 4508
rect 25280 4496 25286 4548
rect 2685 4471 2743 4477
rect 2685 4437 2697 4471
rect 2731 4468 2743 4471
rect 2958 4468 2964 4480
rect 2731 4440 2964 4468
rect 2731 4437 2743 4440
rect 2685 4431 2743 4437
rect 2958 4428 2964 4440
rect 3016 4428 3022 4480
rect 5997 4471 6055 4477
rect 5997 4437 6009 4471
rect 6043 4468 6055 4471
rect 6086 4468 6092 4480
rect 6043 4440 6092 4468
rect 6043 4437 6055 4440
rect 5997 4431 6055 4437
rect 6086 4428 6092 4440
rect 6144 4428 6150 4480
rect 9398 4428 9404 4480
rect 9456 4428 9462 4480
rect 9674 4428 9680 4480
rect 9732 4428 9738 4480
rect 16298 4428 16304 4480
rect 16356 4468 16362 4480
rect 16393 4471 16451 4477
rect 16393 4468 16405 4471
rect 16356 4440 16405 4468
rect 16356 4428 16362 4440
rect 16393 4437 16405 4440
rect 16439 4437 16451 4471
rect 16393 4431 16451 4437
rect 24397 4471 24455 4477
rect 24397 4437 24409 4471
rect 24443 4468 24455 4471
rect 24486 4468 24492 4480
rect 24443 4440 24492 4468
rect 24443 4437 24455 4440
rect 24397 4431 24455 4437
rect 24486 4428 24492 4440
rect 24544 4428 24550 4480
rect 552 4378 27416 4400
rect 552 4326 3756 4378
rect 3808 4326 3820 4378
rect 3872 4326 3884 4378
rect 3936 4326 3948 4378
rect 4000 4326 4012 4378
rect 4064 4326 10472 4378
rect 10524 4326 10536 4378
rect 10588 4326 10600 4378
rect 10652 4326 10664 4378
rect 10716 4326 10728 4378
rect 10780 4326 17188 4378
rect 17240 4326 17252 4378
rect 17304 4326 17316 4378
rect 17368 4326 17380 4378
rect 17432 4326 17444 4378
rect 17496 4326 23904 4378
rect 23956 4326 23968 4378
rect 24020 4326 24032 4378
rect 24084 4326 24096 4378
rect 24148 4326 24160 4378
rect 24212 4326 27416 4378
rect 552 4304 27416 4326
rect 4246 4224 4252 4276
rect 4304 4224 4310 4276
rect 7558 4224 7564 4276
rect 7616 4224 7622 4276
rect 11054 4224 11060 4276
rect 11112 4224 11118 4276
rect 11238 4224 11244 4276
rect 11296 4224 11302 4276
rect 13170 4224 13176 4276
rect 13228 4264 13234 4276
rect 13633 4267 13691 4273
rect 13633 4264 13645 4267
rect 13228 4236 13645 4264
rect 13228 4224 13234 4236
rect 13633 4233 13645 4236
rect 13679 4233 13691 4267
rect 13633 4227 13691 4233
rect 14001 4267 14059 4273
rect 14001 4233 14013 4267
rect 14047 4233 14059 4267
rect 14001 4227 14059 4233
rect 14277 4267 14335 4273
rect 14277 4233 14289 4267
rect 14323 4264 14335 4267
rect 14458 4264 14464 4276
rect 14323 4236 14464 4264
rect 14323 4233 14335 4236
rect 14277 4227 14335 4233
rect 4890 4196 4896 4208
rect 4448 4168 4896 4196
rect 2958 4088 2964 4140
rect 3016 4128 3022 4140
rect 3237 4131 3295 4137
rect 3237 4128 3249 4131
rect 3016 4100 3249 4128
rect 3016 4088 3022 4100
rect 3237 4097 3249 4100
rect 3283 4097 3295 4131
rect 3237 4091 3295 4097
rect 1489 4063 1547 4069
rect 1489 4029 1501 4063
rect 1535 4060 1547 4063
rect 1581 4063 1639 4069
rect 1581 4060 1593 4063
rect 1535 4032 1593 4060
rect 1535 4029 1547 4032
rect 1489 4023 1547 4029
rect 1581 4029 1593 4032
rect 1627 4029 1639 4063
rect 1581 4023 1639 4029
rect 1857 4063 1915 4069
rect 1857 4029 1869 4063
rect 1903 4029 1915 4063
rect 1857 4023 1915 4029
rect 1872 3992 1900 4023
rect 2866 4020 2872 4072
rect 2924 4020 2930 4072
rect 3418 4020 3424 4072
rect 3476 4060 3482 4072
rect 3513 4063 3571 4069
rect 3513 4060 3525 4063
rect 3476 4032 3525 4060
rect 3476 4020 3482 4032
rect 3513 4029 3525 4032
rect 3559 4029 3571 4063
rect 3513 4023 3571 4029
rect 4341 4063 4399 4069
rect 4341 4029 4353 4063
rect 4387 4060 4399 4063
rect 4448 4060 4476 4168
rect 4890 4156 4896 4168
rect 4948 4196 4954 4208
rect 5258 4196 5264 4208
rect 4948 4168 5264 4196
rect 4948 4156 4954 4168
rect 5258 4156 5264 4168
rect 5316 4156 5322 4208
rect 11514 4156 11520 4208
rect 11572 4196 11578 4208
rect 11609 4199 11667 4205
rect 11609 4196 11621 4199
rect 11572 4168 11621 4196
rect 11572 4156 11578 4168
rect 11609 4165 11621 4168
rect 11655 4196 11667 4199
rect 12066 4196 12072 4208
rect 11655 4168 12072 4196
rect 11655 4165 11667 4168
rect 11609 4159 11667 4165
rect 12066 4156 12072 4168
rect 12124 4156 12130 4208
rect 14016 4196 14044 4227
rect 14458 4224 14464 4236
rect 14516 4224 14522 4276
rect 15841 4267 15899 4273
rect 15841 4233 15853 4267
rect 15887 4233 15899 4267
rect 15841 4227 15899 4233
rect 18325 4267 18383 4273
rect 18325 4233 18337 4267
rect 18371 4233 18383 4267
rect 18325 4227 18383 4233
rect 18509 4267 18567 4273
rect 18509 4233 18521 4267
rect 18555 4264 18567 4267
rect 18966 4264 18972 4276
rect 18555 4236 18972 4264
rect 18555 4233 18567 4236
rect 18509 4227 18567 4233
rect 15197 4199 15255 4205
rect 15197 4196 15209 4199
rect 14016 4168 15209 4196
rect 15197 4165 15209 4168
rect 15243 4196 15255 4199
rect 15856 4196 15884 4227
rect 15243 4168 15884 4196
rect 18340 4196 18368 4227
rect 18966 4224 18972 4236
rect 19024 4224 19030 4276
rect 22370 4224 22376 4276
rect 22428 4224 22434 4276
rect 22557 4267 22615 4273
rect 22557 4233 22569 4267
rect 22603 4264 22615 4267
rect 23382 4264 23388 4276
rect 22603 4236 23388 4264
rect 22603 4233 22615 4236
rect 22557 4227 22615 4233
rect 23382 4224 23388 4236
rect 23440 4224 23446 4276
rect 25317 4267 25375 4273
rect 25317 4233 25329 4267
rect 25363 4264 25375 4267
rect 25406 4264 25412 4276
rect 25363 4236 25412 4264
rect 25363 4233 25375 4236
rect 25317 4227 25375 4233
rect 25406 4224 25412 4236
rect 25464 4224 25470 4276
rect 18785 4199 18843 4205
rect 18785 4196 18797 4199
rect 18340 4168 18797 4196
rect 15243 4165 15255 4168
rect 15197 4159 15255 4165
rect 18785 4165 18797 4168
rect 18831 4196 18843 4199
rect 18831 4168 19196 4196
rect 18831 4165 18843 4168
rect 18785 4159 18843 4165
rect 8941 4131 8999 4137
rect 8941 4128 8953 4131
rect 4540 4100 8953 4128
rect 4540 4069 4568 4100
rect 4387 4032 4476 4060
rect 4525 4063 4583 4069
rect 4387 4029 4399 4032
rect 4341 4023 4399 4029
rect 4525 4029 4537 4063
rect 4571 4029 4583 4063
rect 4525 4023 4583 4029
rect 6089 4063 6147 4069
rect 6089 4029 6101 4063
rect 6135 4060 6147 4063
rect 6178 4060 6184 4072
rect 6135 4032 6184 4060
rect 6135 4029 6147 4032
rect 6089 4023 6147 4029
rect 4154 3992 4160 4004
rect 1872 3964 4160 3992
rect 4154 3952 4160 3964
rect 4212 3992 4218 4004
rect 4433 3995 4491 4001
rect 4433 3992 4445 3995
rect 4212 3964 4445 3992
rect 4212 3952 4218 3964
rect 4433 3961 4445 3964
rect 4479 3961 4491 3995
rect 6104 3992 6132 4023
rect 6178 4020 6184 4032
rect 6236 4020 6242 4072
rect 6273 4063 6331 4069
rect 6273 4029 6285 4063
rect 6319 4060 6331 4063
rect 7006 4060 7012 4072
rect 6319 4032 7012 4060
rect 6319 4029 6331 4032
rect 6273 4023 6331 4029
rect 7006 4020 7012 4032
rect 7064 4060 7070 4072
rect 7285 4063 7343 4069
rect 7285 4060 7297 4063
rect 7064 4032 7297 4060
rect 7064 4020 7070 4032
rect 7285 4029 7297 4032
rect 7331 4029 7343 4063
rect 7285 4023 7343 4029
rect 7650 4020 7656 4072
rect 7708 4060 7714 4072
rect 7760 4069 7788 4100
rect 8941 4097 8953 4100
rect 8987 4097 8999 4131
rect 8941 4091 8999 4097
rect 9398 4088 9404 4140
rect 9456 4088 9462 4140
rect 11146 4128 11152 4140
rect 10520 4100 11152 4128
rect 7745 4063 7803 4069
rect 7745 4060 7757 4063
rect 7708 4032 7757 4060
rect 7708 4020 7714 4032
rect 7745 4029 7757 4032
rect 7791 4029 7803 4063
rect 7745 4023 7803 4029
rect 7834 4020 7840 4072
rect 7892 4020 7898 4072
rect 8018 4020 8024 4072
rect 8076 4020 8082 4072
rect 8110 4020 8116 4072
rect 8168 4020 8174 4072
rect 8754 4060 8760 4072
rect 8220 4032 8760 4060
rect 6104 3964 6316 3992
rect 4433 3955 4491 3961
rect 2314 3884 2320 3936
rect 2372 3924 2378 3936
rect 2593 3927 2651 3933
rect 2593 3924 2605 3927
rect 2372 3896 2605 3924
rect 2372 3884 2378 3896
rect 2593 3893 2605 3896
rect 2639 3893 2651 3927
rect 2593 3887 2651 3893
rect 3053 3927 3111 3933
rect 3053 3893 3065 3927
rect 3099 3924 3111 3927
rect 3234 3924 3240 3936
rect 3099 3896 3240 3924
rect 3099 3893 3111 3896
rect 3053 3887 3111 3893
rect 3234 3884 3240 3896
rect 3292 3884 3298 3936
rect 5994 3884 6000 3936
rect 6052 3924 6058 3936
rect 6181 3927 6239 3933
rect 6181 3924 6193 3927
rect 6052 3896 6193 3924
rect 6052 3884 6058 3896
rect 6181 3893 6193 3896
rect 6227 3893 6239 3927
rect 6288 3924 6316 3964
rect 6914 3952 6920 4004
rect 6972 3992 6978 4004
rect 7101 3995 7159 4001
rect 7101 3992 7113 3995
rect 6972 3964 7113 3992
rect 6972 3952 6978 3964
rect 7101 3961 7113 3964
rect 7147 3961 7159 3995
rect 7101 3955 7159 3961
rect 7469 3995 7527 4001
rect 7469 3961 7481 3995
rect 7515 3992 7527 3995
rect 8220 3992 8248 4032
rect 8754 4020 8760 4032
rect 8812 4060 8818 4072
rect 8849 4063 8907 4069
rect 8849 4060 8861 4063
rect 8812 4032 8861 4060
rect 8812 4020 8818 4032
rect 8849 4029 8861 4032
rect 8895 4029 8907 4063
rect 8849 4023 8907 4029
rect 9030 4020 9036 4072
rect 9088 4020 9094 4072
rect 10520 4069 10548 4100
rect 11146 4088 11152 4100
rect 11204 4088 11210 4140
rect 15289 4131 15347 4137
rect 15289 4128 15301 4131
rect 12636 4100 13216 4128
rect 9677 4063 9735 4069
rect 9677 4029 9689 4063
rect 9723 4029 9735 4063
rect 9677 4023 9735 4029
rect 10505 4063 10563 4069
rect 10505 4029 10517 4063
rect 10551 4029 10563 4063
rect 10505 4023 10563 4029
rect 10689 4063 10747 4069
rect 10689 4029 10701 4063
rect 10735 4060 10747 4063
rect 11238 4060 11244 4072
rect 10735 4032 11244 4060
rect 10735 4029 10747 4032
rect 10689 4023 10747 4029
rect 7515 3964 8248 3992
rect 7515 3961 7527 3964
rect 7469 3955 7527 3961
rect 7484 3924 7512 3955
rect 8570 3952 8576 4004
rect 8628 3992 8634 4004
rect 9048 3992 9076 4020
rect 8628 3964 9076 3992
rect 9692 3992 9720 4023
rect 11238 4020 11244 4032
rect 11296 4060 11302 4072
rect 11790 4060 11796 4072
rect 11296 4032 11796 4060
rect 11296 4020 11302 4032
rect 11790 4020 11796 4032
rect 11848 4060 11854 4072
rect 12342 4060 12348 4072
rect 11848 4032 12348 4060
rect 11848 4020 11854 4032
rect 12342 4020 12348 4032
rect 12400 4060 12406 4072
rect 12636 4069 12664 4100
rect 12621 4063 12679 4069
rect 12621 4060 12633 4063
rect 12400 4032 12633 4060
rect 12400 4020 12406 4032
rect 12621 4029 12633 4032
rect 12667 4029 12679 4063
rect 12621 4023 12679 4029
rect 12802 4020 12808 4072
rect 12860 4020 12866 4072
rect 13188 4069 13216 4100
rect 15028 4100 15301 4128
rect 13173 4063 13231 4069
rect 13173 4029 13185 4063
rect 13219 4029 13231 4063
rect 13173 4023 13231 4029
rect 13265 4063 13323 4069
rect 13265 4029 13277 4063
rect 13311 4060 13323 4063
rect 13817 4063 13875 4069
rect 13817 4060 13829 4063
rect 13311 4032 13829 4060
rect 13311 4029 13323 4032
rect 13265 4023 13323 4029
rect 13817 4029 13829 4032
rect 13863 4029 13875 4063
rect 13817 4023 13875 4029
rect 14001 4063 14059 4069
rect 14001 4029 14013 4063
rect 14047 4029 14059 4063
rect 14001 4023 14059 4029
rect 14093 4063 14151 4069
rect 14093 4029 14105 4063
rect 14139 4060 14151 4063
rect 14182 4060 14188 4072
rect 14139 4032 14188 4060
rect 14139 4029 14151 4032
rect 14093 4023 14151 4029
rect 10597 3995 10655 4001
rect 10597 3992 10609 3995
rect 9692 3964 10609 3992
rect 8628 3952 8634 3964
rect 10597 3961 10609 3964
rect 10643 3961 10655 3995
rect 10597 3955 10655 3961
rect 13722 3952 13728 4004
rect 13780 3992 13786 4004
rect 14016 3992 14044 4023
rect 14182 4020 14188 4032
rect 14240 4020 14246 4072
rect 14734 4020 14740 4072
rect 14792 4060 14798 4072
rect 15028 4069 15056 4100
rect 15289 4097 15301 4100
rect 15335 4097 15347 4131
rect 15289 4091 15347 4097
rect 16298 4088 16304 4140
rect 16356 4088 16362 4140
rect 18322 4088 18328 4140
rect 18380 4128 18386 4140
rect 19168 4137 19196 4168
rect 19242 4156 19248 4208
rect 19300 4196 19306 4208
rect 19300 4168 21579 4196
rect 19300 4156 19334 4168
rect 19306 4137 19334 4156
rect 19153 4131 19211 4137
rect 18380 4100 18920 4128
rect 18380 4088 18386 4100
rect 15013 4063 15071 4069
rect 15013 4060 15025 4063
rect 14792 4032 15025 4060
rect 14792 4020 14798 4032
rect 15013 4029 15025 4032
rect 15059 4029 15071 4063
rect 15197 4063 15255 4069
rect 15197 4060 15209 4063
rect 15013 4023 15071 4029
rect 15120 4032 15209 4060
rect 13780 3964 14044 3992
rect 13780 3952 13786 3964
rect 6288 3896 7512 3924
rect 6181 3887 6239 3893
rect 7558 3884 7564 3936
rect 7616 3924 7622 3936
rect 8389 3927 8447 3933
rect 8389 3924 8401 3927
rect 7616 3896 8401 3924
rect 7616 3884 7622 3896
rect 8389 3893 8401 3896
rect 8435 3893 8447 3927
rect 8389 3887 8447 3893
rect 10413 3927 10471 3933
rect 10413 3893 10425 3927
rect 10459 3924 10471 3927
rect 10870 3924 10876 3936
rect 10459 3896 10876 3924
rect 10459 3893 10471 3896
rect 10413 3887 10471 3893
rect 10870 3884 10876 3896
rect 10928 3884 10934 3936
rect 11146 3884 11152 3936
rect 11204 3924 11210 3936
rect 11241 3927 11299 3933
rect 11241 3924 11253 3927
rect 11204 3896 11253 3924
rect 11204 3884 11210 3896
rect 11241 3893 11253 3896
rect 11287 3893 11299 3927
rect 11241 3887 11299 3893
rect 12710 3884 12716 3936
rect 12768 3884 12774 3936
rect 12802 3884 12808 3936
rect 12860 3924 12866 3936
rect 15120 3924 15148 4032
rect 15197 4029 15209 4032
rect 15243 4060 15255 4063
rect 15470 4060 15476 4072
rect 15243 4032 15476 4060
rect 15243 4029 15255 4032
rect 15197 4023 15255 4029
rect 15470 4020 15476 4032
rect 15528 4020 15534 4072
rect 15657 4063 15715 4069
rect 15657 4029 15669 4063
rect 15703 4060 15715 4063
rect 15841 4063 15899 4069
rect 15841 4060 15853 4063
rect 15703 4032 15853 4060
rect 15703 4029 15715 4032
rect 15657 4023 15715 4029
rect 15841 4029 15853 4032
rect 15887 4029 15899 4063
rect 15841 4023 15899 4029
rect 15930 4020 15936 4072
rect 15988 4020 15994 4072
rect 16482 4020 16488 4072
rect 16540 4060 16546 4072
rect 16577 4063 16635 4069
rect 16577 4060 16589 4063
rect 16540 4032 16589 4060
rect 16540 4020 16546 4032
rect 16577 4029 16589 4032
rect 16623 4029 16635 4063
rect 16577 4023 16635 4029
rect 16758 4020 16764 4072
rect 16816 4060 16822 4072
rect 17589 4063 17647 4069
rect 17589 4060 17601 4063
rect 16816 4032 17601 4060
rect 16816 4020 16822 4032
rect 17589 4029 17601 4032
rect 17635 4029 17647 4063
rect 17589 4023 17647 4029
rect 17957 4063 18015 4069
rect 17957 4029 17969 4063
rect 18003 4060 18015 4063
rect 18230 4060 18236 4072
rect 18003 4032 18236 4060
rect 18003 4029 18015 4032
rect 17957 4023 18015 4029
rect 17402 3992 17408 4004
rect 16132 3964 17408 3992
rect 12860 3896 15148 3924
rect 12860 3884 12866 3896
rect 15194 3884 15200 3936
rect 15252 3924 15258 3936
rect 16132 3924 16160 3964
rect 17402 3952 17408 3964
rect 17460 3952 17466 4004
rect 17604 3992 17632 4023
rect 18230 4020 18236 4032
rect 18288 4020 18294 4072
rect 18690 4060 18696 4072
rect 18432 4056 18696 4060
rect 18340 4032 18696 4056
rect 18340 4028 18460 4032
rect 18340 3992 18368 4028
rect 18690 4020 18696 4032
rect 18748 4020 18754 4072
rect 18782 4020 18788 4072
rect 18840 4060 18846 4072
rect 18892 4069 18920 4100
rect 19153 4097 19165 4131
rect 19199 4097 19211 4131
rect 19306 4131 19386 4137
rect 19306 4100 19340 4131
rect 19153 4091 19211 4097
rect 19328 4097 19340 4100
rect 19374 4097 19386 4131
rect 19328 4091 19386 4097
rect 19422 4131 19480 4137
rect 19422 4097 19434 4131
rect 19468 4128 19480 4131
rect 19705 4131 19763 4137
rect 19705 4128 19717 4131
rect 19468 4100 19717 4128
rect 19468 4097 19480 4100
rect 19422 4091 19480 4097
rect 19705 4097 19717 4100
rect 19751 4097 19763 4131
rect 19705 4091 19763 4097
rect 18877 4063 18935 4069
rect 18877 4060 18889 4063
rect 18840 4032 18889 4060
rect 18840 4020 18846 4032
rect 18877 4029 18889 4032
rect 18923 4029 18935 4063
rect 18877 4023 18935 4029
rect 18966 4020 18972 4072
rect 19024 4060 19030 4072
rect 20640 4069 20668 4168
rect 20714 4088 20720 4140
rect 20772 4128 20778 4140
rect 21358 4128 21364 4140
rect 20772 4100 21364 4128
rect 20772 4088 20778 4100
rect 21358 4088 21364 4100
rect 21416 4088 21422 4140
rect 21551 4069 21579 4168
rect 21637 4131 21695 4137
rect 21637 4097 21649 4131
rect 21683 4128 21695 4131
rect 22281 4131 22339 4137
rect 22281 4128 22293 4131
rect 21683 4100 22293 4128
rect 21683 4097 21695 4100
rect 21637 4091 21695 4097
rect 22281 4097 22293 4100
rect 22327 4097 22339 4131
rect 22281 4091 22339 4097
rect 19245 4063 19303 4069
rect 19245 4060 19257 4063
rect 19024 4032 19257 4060
rect 19024 4020 19030 4032
rect 19245 4029 19257 4032
rect 19291 4060 19303 4063
rect 19613 4063 19671 4069
rect 19613 4060 19625 4063
rect 19291 4032 19625 4060
rect 19291 4029 19303 4032
rect 19245 4023 19303 4029
rect 19613 4029 19625 4032
rect 19659 4029 19671 4063
rect 19613 4023 19671 4029
rect 19797 4063 19855 4069
rect 19797 4029 19809 4063
rect 19843 4029 19855 4063
rect 19797 4023 19855 4029
rect 20625 4063 20683 4069
rect 20625 4029 20637 4063
rect 20671 4029 20683 4063
rect 20625 4023 20683 4029
rect 20809 4063 20867 4069
rect 20809 4029 20821 4063
rect 20855 4029 20867 4063
rect 20809 4023 20867 4029
rect 21545 4063 21603 4069
rect 21545 4029 21557 4063
rect 21591 4029 21603 4063
rect 21545 4023 21603 4029
rect 17604 3964 18368 3992
rect 18506 3952 18512 4004
rect 18564 3992 18570 4004
rect 19812 3992 19840 4023
rect 20162 3992 20168 4004
rect 18564 3964 20168 3992
rect 18564 3952 18570 3964
rect 20162 3952 20168 3964
rect 20220 3952 20226 4004
rect 20438 3952 20444 4004
rect 20496 3992 20502 4004
rect 20824 3992 20852 4023
rect 22186 4020 22192 4072
rect 22244 4020 22250 4072
rect 22922 4020 22928 4072
rect 22980 4060 22986 4072
rect 23017 4063 23075 4069
rect 23017 4060 23029 4063
rect 22980 4032 23029 4060
rect 22980 4020 22986 4032
rect 23017 4029 23029 4032
rect 23063 4029 23075 4063
rect 23198 4060 23204 4072
rect 23017 4023 23075 4029
rect 23124 4032 23204 4060
rect 23124 3992 23152 4032
rect 23198 4020 23204 4032
rect 23256 4020 23262 4072
rect 23477 4063 23535 4069
rect 23477 4029 23489 4063
rect 23523 4060 23535 4063
rect 23750 4060 23756 4072
rect 23523 4032 23756 4060
rect 23523 4029 23535 4032
rect 23477 4023 23535 4029
rect 23750 4020 23756 4032
rect 23808 4020 23814 4072
rect 24213 4063 24271 4069
rect 24213 4029 24225 4063
rect 24259 4060 24271 4063
rect 24305 4063 24363 4069
rect 24305 4060 24317 4063
rect 24259 4032 24317 4060
rect 24259 4029 24271 4032
rect 24213 4023 24271 4029
rect 24305 4029 24317 4032
rect 24351 4029 24363 4063
rect 24305 4023 24363 4029
rect 24581 4063 24639 4069
rect 24581 4029 24593 4063
rect 24627 4029 24639 4063
rect 24581 4023 24639 4029
rect 24596 3992 24624 4023
rect 20496 3964 20852 3992
rect 20496 3952 20502 3964
rect 15252 3896 16160 3924
rect 16209 3927 16267 3933
rect 15252 3884 15258 3896
rect 16209 3893 16221 3927
rect 16255 3924 16267 3927
rect 16298 3924 16304 3936
rect 16255 3896 16304 3924
rect 16255 3893 16267 3896
rect 16209 3887 16267 3893
rect 16298 3884 16304 3896
rect 16356 3884 16362 3936
rect 17034 3884 17040 3936
rect 17092 3924 17098 3936
rect 17313 3927 17371 3933
rect 17313 3924 17325 3927
rect 17092 3896 17325 3924
rect 17092 3884 17098 3896
rect 17313 3893 17325 3896
rect 17359 3893 17371 3927
rect 17313 3887 17371 3893
rect 17773 3927 17831 3933
rect 17773 3893 17785 3927
rect 17819 3924 17831 3927
rect 17862 3924 17868 3936
rect 17819 3896 17868 3924
rect 17819 3893 17831 3896
rect 17773 3887 17831 3893
rect 17862 3884 17868 3896
rect 17920 3884 17926 3936
rect 18322 3884 18328 3936
rect 18380 3884 18386 3936
rect 18969 3927 19027 3933
rect 18969 3893 18981 3927
rect 19015 3924 19027 3927
rect 19978 3924 19984 3936
rect 19015 3896 19984 3924
rect 19015 3893 19027 3896
rect 18969 3887 19027 3893
rect 19978 3884 19984 3896
rect 20036 3884 20042 3936
rect 20824 3924 20852 3964
rect 22296 3964 23152 3992
rect 23676 3964 24624 3992
rect 22296 3924 22324 3964
rect 20824 3896 22324 3924
rect 22370 3884 22376 3936
rect 22428 3924 22434 3936
rect 23109 3927 23167 3933
rect 23109 3924 23121 3927
rect 22428 3896 23121 3924
rect 22428 3884 22434 3896
rect 23109 3893 23121 3896
rect 23155 3924 23167 3927
rect 23382 3924 23388 3936
rect 23155 3896 23388 3924
rect 23155 3893 23167 3896
rect 23109 3887 23167 3893
rect 23382 3884 23388 3896
rect 23440 3884 23446 3936
rect 23676 3933 23704 3964
rect 23661 3927 23719 3933
rect 23661 3893 23673 3927
rect 23707 3893 23719 3927
rect 23661 3887 23719 3893
rect 552 3834 27576 3856
rect 552 3782 7114 3834
rect 7166 3782 7178 3834
rect 7230 3782 7242 3834
rect 7294 3782 7306 3834
rect 7358 3782 7370 3834
rect 7422 3782 13830 3834
rect 13882 3782 13894 3834
rect 13946 3782 13958 3834
rect 14010 3782 14022 3834
rect 14074 3782 14086 3834
rect 14138 3782 20546 3834
rect 20598 3782 20610 3834
rect 20662 3782 20674 3834
rect 20726 3782 20738 3834
rect 20790 3782 20802 3834
rect 20854 3782 27262 3834
rect 27314 3782 27326 3834
rect 27378 3782 27390 3834
rect 27442 3782 27454 3834
rect 27506 3782 27518 3834
rect 27570 3782 27576 3834
rect 552 3760 27576 3782
rect 2866 3680 2872 3732
rect 2924 3720 2930 3732
rect 4985 3723 5043 3729
rect 2924 3692 4752 3720
rect 2924 3680 2930 3692
rect 3697 3655 3755 3661
rect 3697 3621 3709 3655
rect 3743 3652 3755 3655
rect 3973 3655 4031 3661
rect 3973 3652 3985 3655
rect 3743 3624 3985 3652
rect 3743 3621 3755 3624
rect 3697 3615 3755 3621
rect 3973 3621 3985 3624
rect 4019 3652 4031 3655
rect 4246 3652 4252 3664
rect 4019 3624 4252 3652
rect 4019 3621 4031 3624
rect 3973 3615 4031 3621
rect 4246 3612 4252 3624
rect 4304 3612 4310 3664
rect 4724 3652 4752 3692
rect 4985 3689 4997 3723
rect 5031 3720 5043 3723
rect 5166 3720 5172 3732
rect 5031 3692 5172 3720
rect 5031 3689 5043 3692
rect 4985 3683 5043 3689
rect 5166 3680 5172 3692
rect 5224 3680 5230 3732
rect 6457 3723 6515 3729
rect 6457 3689 6469 3723
rect 6503 3689 6515 3723
rect 7561 3723 7619 3729
rect 7561 3720 7573 3723
rect 6457 3683 6515 3689
rect 7392 3692 7573 3720
rect 6472 3652 6500 3683
rect 4724 3624 6500 3652
rect 7006 3612 7012 3664
rect 7064 3612 7070 3664
rect 3602 3544 3608 3596
rect 3660 3544 3666 3596
rect 3881 3587 3939 3593
rect 3881 3553 3893 3587
rect 3927 3584 3939 3587
rect 4062 3584 4068 3596
rect 3927 3556 4068 3584
rect 3927 3553 3939 3556
rect 3881 3547 3939 3553
rect 4062 3544 4068 3556
rect 4120 3544 4126 3596
rect 4154 3544 4160 3596
rect 4212 3544 4218 3596
rect 4341 3587 4399 3593
rect 4341 3553 4353 3587
rect 4387 3584 4399 3587
rect 4617 3587 4675 3593
rect 4617 3584 4629 3587
rect 4387 3556 4629 3584
rect 4387 3553 4399 3556
rect 4341 3547 4399 3553
rect 4617 3553 4629 3556
rect 4663 3553 4675 3587
rect 4617 3547 4675 3553
rect 6086 3544 6092 3596
rect 6144 3544 6150 3596
rect 6270 3544 6276 3596
rect 6328 3544 6334 3596
rect 6822 3544 6828 3596
rect 6880 3544 6886 3596
rect 6917 3587 6975 3593
rect 6917 3553 6929 3587
rect 6963 3584 6975 3587
rect 7024 3584 7052 3612
rect 6963 3556 7052 3584
rect 6963 3553 6975 3556
rect 6917 3547 6975 3553
rect 4709 3519 4767 3525
rect 4709 3485 4721 3519
rect 4755 3516 4767 3519
rect 6181 3519 6239 3525
rect 6181 3516 6193 3519
rect 4755 3488 6193 3516
rect 4755 3485 4767 3488
rect 4709 3479 4767 3485
rect 6181 3485 6193 3488
rect 6227 3516 6239 3519
rect 6546 3516 6552 3528
rect 6227 3488 6552 3516
rect 6227 3485 6239 3488
rect 6181 3479 6239 3485
rect 6546 3476 6552 3488
rect 6604 3476 6610 3528
rect 6733 3519 6791 3525
rect 6733 3485 6745 3519
rect 6779 3516 6791 3519
rect 7009 3519 7067 3525
rect 7009 3516 7021 3519
rect 6779 3488 7021 3516
rect 6779 3485 6791 3488
rect 6733 3479 6791 3485
rect 7009 3485 7021 3488
rect 7055 3485 7067 3519
rect 7009 3479 7067 3485
rect 3510 3408 3516 3460
rect 3568 3448 3574 3460
rect 5350 3448 5356 3460
rect 3568 3420 5356 3448
rect 3568 3408 3574 3420
rect 5350 3408 5356 3420
rect 5408 3448 5414 3460
rect 7282 3448 7288 3460
rect 5408 3420 7288 3448
rect 5408 3408 5414 3420
rect 7282 3408 7288 3420
rect 7340 3408 7346 3460
rect 4798 3340 4804 3392
rect 4856 3340 4862 3392
rect 6825 3383 6883 3389
rect 6825 3349 6837 3383
rect 6871 3380 6883 3383
rect 7392 3380 7420 3692
rect 7561 3689 7573 3692
rect 7607 3720 7619 3723
rect 8018 3720 8024 3732
rect 7607 3692 8024 3720
rect 7607 3689 7619 3692
rect 7561 3683 7619 3689
rect 8018 3680 8024 3692
rect 8076 3680 8082 3732
rect 9674 3720 9680 3732
rect 9324 3692 9680 3720
rect 7834 3652 7840 3664
rect 7484 3624 7840 3652
rect 7484 3593 7512 3624
rect 7834 3612 7840 3624
rect 7892 3612 7898 3664
rect 8754 3652 8760 3664
rect 8220 3624 8760 3652
rect 7469 3587 7527 3593
rect 7469 3553 7481 3587
rect 7515 3553 7527 3587
rect 7469 3547 7527 3553
rect 7650 3544 7656 3596
rect 7708 3544 7714 3596
rect 8220 3593 8248 3624
rect 8754 3612 8760 3624
rect 8812 3612 8818 3664
rect 8205 3587 8263 3593
rect 8205 3553 8217 3587
rect 8251 3553 8263 3587
rect 8205 3547 8263 3553
rect 8389 3587 8447 3593
rect 8389 3553 8401 3587
rect 8435 3584 8447 3587
rect 8570 3584 8576 3596
rect 8435 3556 8576 3584
rect 8435 3553 8447 3556
rect 8389 3547 8447 3553
rect 8570 3544 8576 3556
rect 8628 3544 8634 3596
rect 9125 3587 9183 3593
rect 9125 3553 9137 3587
rect 9171 3584 9183 3587
rect 9324 3584 9352 3692
rect 9674 3680 9680 3692
rect 9732 3680 9738 3732
rect 10134 3680 10140 3732
rect 10192 3680 10198 3732
rect 12345 3723 12403 3729
rect 12345 3689 12357 3723
rect 12391 3720 12403 3723
rect 12802 3720 12808 3732
rect 12391 3692 12808 3720
rect 12391 3689 12403 3692
rect 12345 3683 12403 3689
rect 12802 3680 12808 3692
rect 12860 3680 12866 3732
rect 13909 3723 13967 3729
rect 13909 3689 13921 3723
rect 13955 3720 13967 3723
rect 14182 3720 14188 3732
rect 13955 3692 14188 3720
rect 13955 3689 13967 3692
rect 13909 3683 13967 3689
rect 14182 3680 14188 3692
rect 14240 3680 14246 3732
rect 15470 3680 15476 3732
rect 15528 3729 15534 3732
rect 15528 3723 15547 3729
rect 15535 3689 15547 3723
rect 15528 3683 15547 3689
rect 15528 3680 15534 3683
rect 15930 3680 15936 3732
rect 15988 3680 15994 3732
rect 16482 3680 16488 3732
rect 16540 3680 16546 3732
rect 17402 3680 17408 3732
rect 17460 3720 17466 3732
rect 17460 3692 18276 3720
rect 17460 3680 17466 3692
rect 12710 3652 12716 3664
rect 9416 3624 12716 3652
rect 9416 3593 9444 3624
rect 12710 3612 12716 3624
rect 12768 3652 12774 3664
rect 12768 3624 12940 3652
rect 12768 3612 12774 3624
rect 9171 3556 9352 3584
rect 9401 3587 9459 3593
rect 9171 3553 9183 3556
rect 9125 3547 9183 3553
rect 9401 3553 9413 3587
rect 9447 3553 9459 3587
rect 9401 3547 9459 3553
rect 10962 3544 10968 3596
rect 11020 3544 11026 3596
rect 11146 3544 11152 3596
rect 11204 3584 11210 3596
rect 11974 3584 11980 3596
rect 11204 3556 11980 3584
rect 11204 3544 11210 3556
rect 11974 3544 11980 3556
rect 12032 3584 12038 3596
rect 12437 3587 12495 3593
rect 12437 3584 12449 3587
rect 12032 3556 12449 3584
rect 12032 3544 12038 3556
rect 10980 3516 11008 3544
rect 11885 3519 11943 3525
rect 11885 3516 11897 3519
rect 10980 3488 11897 3516
rect 11885 3485 11897 3488
rect 11931 3485 11943 3519
rect 11885 3479 11943 3485
rect 6871 3352 7420 3380
rect 6871 3349 6883 3352
rect 6825 3343 6883 3349
rect 8018 3340 8024 3392
rect 8076 3380 8082 3392
rect 8297 3383 8355 3389
rect 8297 3380 8309 3383
rect 8076 3352 8309 3380
rect 8076 3340 8082 3352
rect 8297 3349 8309 3352
rect 8343 3349 8355 3383
rect 8297 3343 8355 3349
rect 11054 3340 11060 3392
rect 11112 3340 11118 3392
rect 11900 3380 11928 3479
rect 12176 3457 12204 3556
rect 12437 3553 12449 3556
rect 12483 3553 12495 3587
rect 12437 3547 12495 3553
rect 12621 3587 12679 3593
rect 12621 3553 12633 3587
rect 12667 3553 12679 3587
rect 12621 3547 12679 3553
rect 12161 3451 12219 3457
rect 12161 3417 12173 3451
rect 12207 3417 12219 3451
rect 12161 3411 12219 3417
rect 12636 3380 12664 3547
rect 12912 3516 12940 3624
rect 15102 3612 15108 3664
rect 15160 3652 15166 3664
rect 15289 3655 15347 3661
rect 15289 3652 15301 3655
rect 15160 3624 15301 3652
rect 15160 3612 15166 3624
rect 15289 3621 15301 3624
rect 15335 3621 15347 3655
rect 15948 3652 15976 3680
rect 17034 3652 17040 3664
rect 15948 3624 17040 3652
rect 15289 3615 15347 3621
rect 17034 3612 17040 3624
rect 17092 3612 17098 3664
rect 17862 3612 17868 3664
rect 17920 3612 17926 3664
rect 18248 3661 18276 3692
rect 18322 3680 18328 3732
rect 18380 3720 18386 3732
rect 18874 3720 18880 3732
rect 18380 3692 18880 3720
rect 18380 3680 18386 3692
rect 18874 3680 18880 3692
rect 18932 3680 18938 3732
rect 19981 3723 20039 3729
rect 19981 3689 19993 3723
rect 20027 3720 20039 3723
rect 20438 3720 20444 3732
rect 20027 3692 20444 3720
rect 20027 3689 20039 3692
rect 19981 3683 20039 3689
rect 20438 3680 20444 3692
rect 20496 3680 20502 3732
rect 21818 3680 21824 3732
rect 21876 3680 21882 3732
rect 25130 3680 25136 3732
rect 25188 3720 25194 3732
rect 25501 3723 25559 3729
rect 25501 3720 25513 3723
rect 25188 3692 25513 3720
rect 25188 3680 25194 3692
rect 25501 3689 25513 3692
rect 25547 3689 25559 3723
rect 25501 3683 25559 3689
rect 18233 3655 18291 3661
rect 18233 3621 18245 3655
rect 18279 3621 18291 3655
rect 18233 3615 18291 3621
rect 18690 3612 18696 3664
rect 18748 3652 18754 3664
rect 20809 3655 20867 3661
rect 18748 3624 20576 3652
rect 18748 3612 18754 3624
rect 13446 3544 13452 3596
rect 13504 3544 13510 3596
rect 13725 3587 13783 3593
rect 13725 3553 13737 3587
rect 13771 3584 13783 3587
rect 14182 3584 14188 3596
rect 13771 3556 14188 3584
rect 13771 3553 13783 3556
rect 13725 3547 13783 3553
rect 14182 3544 14188 3556
rect 14240 3544 14246 3596
rect 15378 3544 15384 3596
rect 15436 3584 15442 3596
rect 15749 3587 15807 3593
rect 15749 3584 15761 3587
rect 15436 3556 15761 3584
rect 15436 3544 15442 3556
rect 15749 3553 15761 3556
rect 15795 3553 15807 3587
rect 15749 3547 15807 3553
rect 16298 3544 16304 3596
rect 16356 3544 16362 3596
rect 18782 3544 18788 3596
rect 18840 3544 18846 3596
rect 18966 3544 18972 3596
rect 19024 3544 19030 3596
rect 19150 3544 19156 3596
rect 19208 3584 19214 3596
rect 19521 3587 19579 3593
rect 19521 3584 19533 3587
rect 19208 3556 19533 3584
rect 19208 3544 19214 3556
rect 19521 3553 19533 3556
rect 19567 3553 19579 3587
rect 19521 3547 19579 3553
rect 20162 3544 20168 3596
rect 20220 3544 20226 3596
rect 20548 3593 20576 3624
rect 20809 3621 20821 3655
rect 20855 3652 20867 3655
rect 21361 3655 21419 3661
rect 21361 3652 21373 3655
rect 20855 3624 21373 3652
rect 20855 3621 20867 3624
rect 20809 3615 20867 3621
rect 21361 3621 21373 3624
rect 21407 3621 21419 3655
rect 21361 3615 21419 3621
rect 23106 3612 23112 3664
rect 23164 3652 23170 3664
rect 23753 3655 23811 3661
rect 23753 3652 23765 3655
rect 23164 3624 23765 3652
rect 23164 3612 23170 3624
rect 23753 3621 23765 3624
rect 23799 3621 23811 3655
rect 23753 3615 23811 3621
rect 23983 3621 24041 3627
rect 23983 3618 23995 3621
rect 20533 3587 20591 3593
rect 20533 3553 20545 3587
rect 20579 3553 20591 3587
rect 20533 3547 20591 3553
rect 13633 3519 13691 3525
rect 12912 3488 13492 3516
rect 11900 3352 12664 3380
rect 12802 3340 12808 3392
rect 12860 3340 12866 3392
rect 13464 3389 13492 3488
rect 13633 3485 13645 3519
rect 13679 3516 13691 3519
rect 14274 3516 14280 3528
rect 13679 3488 14280 3516
rect 13679 3485 13691 3488
rect 13633 3479 13691 3485
rect 14274 3476 14280 3488
rect 14332 3476 14338 3528
rect 17954 3476 17960 3528
rect 18012 3516 18018 3528
rect 18049 3519 18107 3525
rect 18049 3516 18061 3519
rect 18012 3488 18061 3516
rect 18012 3476 18018 3488
rect 18049 3485 18061 3488
rect 18095 3516 18107 3519
rect 18138 3516 18144 3528
rect 18095 3488 18144 3516
rect 18095 3485 18107 3488
rect 18049 3479 18107 3485
rect 18138 3476 18144 3488
rect 18196 3516 18202 3528
rect 18598 3516 18604 3528
rect 18196 3488 18604 3516
rect 18196 3476 18202 3488
rect 18598 3476 18604 3488
rect 18656 3516 18662 3528
rect 19242 3516 19248 3528
rect 18656 3488 19248 3516
rect 18656 3476 18662 3488
rect 19242 3476 19248 3488
rect 19300 3476 19306 3528
rect 15657 3451 15715 3457
rect 15657 3417 15669 3451
rect 15703 3448 15715 3451
rect 16298 3448 16304 3460
rect 15703 3420 16304 3448
rect 15703 3417 15715 3420
rect 15657 3411 15715 3417
rect 16298 3408 16304 3420
rect 16356 3408 16362 3460
rect 18230 3408 18236 3460
rect 18288 3448 18294 3460
rect 18417 3451 18475 3457
rect 18417 3448 18429 3451
rect 18288 3420 18429 3448
rect 18288 3408 18294 3420
rect 18417 3417 18429 3420
rect 18463 3417 18475 3451
rect 18417 3411 18475 3417
rect 18966 3408 18972 3460
rect 19024 3448 19030 3460
rect 19797 3451 19855 3457
rect 19797 3448 19809 3451
rect 19024 3420 19809 3448
rect 19024 3408 19030 3420
rect 19797 3417 19809 3420
rect 19843 3417 19855 3451
rect 20548 3448 20576 3547
rect 20714 3544 20720 3596
rect 20772 3544 20778 3596
rect 20901 3587 20959 3593
rect 20901 3553 20913 3587
rect 20947 3553 20959 3587
rect 20901 3547 20959 3553
rect 21637 3587 21695 3593
rect 21637 3553 21649 3587
rect 21683 3584 21695 3587
rect 22554 3584 22560 3596
rect 21683 3556 22560 3584
rect 21683 3553 21695 3556
rect 21637 3547 21695 3553
rect 20622 3476 20628 3528
rect 20680 3516 20686 3528
rect 20916 3516 20944 3547
rect 22554 3544 22560 3556
rect 22612 3544 22618 3596
rect 23198 3544 23204 3596
rect 23256 3584 23262 3596
rect 23477 3587 23535 3593
rect 23477 3584 23489 3587
rect 23256 3556 23489 3584
rect 23256 3544 23262 3556
rect 23477 3553 23489 3556
rect 23523 3584 23535 3587
rect 23968 3587 23995 3618
rect 24029 3587 24041 3621
rect 23968 3584 24041 3587
rect 23523 3581 24041 3584
rect 23523 3556 23996 3581
rect 23523 3553 23535 3556
rect 23477 3547 23535 3553
rect 24762 3544 24768 3596
rect 24820 3544 24826 3596
rect 20680 3488 20944 3516
rect 21545 3519 21603 3525
rect 20680 3476 20686 3488
rect 21545 3485 21557 3519
rect 21591 3516 21603 3519
rect 22830 3516 22836 3528
rect 21591 3488 22836 3516
rect 21591 3485 21603 3488
rect 21545 3479 21603 3485
rect 22830 3476 22836 3488
rect 22888 3476 22894 3528
rect 23293 3519 23351 3525
rect 23293 3516 23305 3519
rect 22940 3488 23305 3516
rect 21634 3448 21640 3460
rect 20548 3420 21640 3448
rect 19797 3411 19855 3417
rect 21634 3408 21640 3420
rect 21692 3408 21698 3460
rect 22940 3392 22968 3488
rect 23293 3485 23305 3488
rect 23339 3485 23351 3519
rect 23293 3479 23351 3485
rect 24397 3519 24455 3525
rect 24397 3485 24409 3519
rect 24443 3516 24455 3519
rect 24489 3519 24547 3525
rect 24489 3516 24501 3519
rect 24443 3488 24501 3516
rect 24443 3485 24455 3488
rect 24397 3479 24455 3485
rect 24489 3485 24501 3488
rect 24535 3485 24547 3519
rect 24489 3479 24547 3485
rect 23308 3448 23336 3479
rect 23308 3420 23980 3448
rect 13449 3383 13507 3389
rect 13449 3349 13461 3383
rect 13495 3349 13507 3383
rect 13449 3343 13507 3349
rect 15470 3340 15476 3392
rect 15528 3340 15534 3392
rect 16390 3340 16396 3392
rect 16448 3380 16454 3392
rect 16577 3383 16635 3389
rect 16577 3380 16589 3383
rect 16448 3352 16589 3380
rect 16448 3340 16454 3352
rect 16577 3349 16589 3352
rect 16623 3349 16635 3383
rect 16577 3343 16635 3349
rect 20438 3340 20444 3392
rect 20496 3380 20502 3392
rect 20533 3383 20591 3389
rect 20533 3380 20545 3383
rect 20496 3352 20545 3380
rect 20496 3340 20502 3352
rect 20533 3349 20545 3352
rect 20579 3380 20591 3383
rect 20622 3380 20628 3392
rect 20579 3352 20628 3380
rect 20579 3349 20591 3352
rect 20533 3343 20591 3349
rect 20622 3340 20628 3352
rect 20680 3340 20686 3392
rect 21358 3340 21364 3392
rect 21416 3340 21422 3392
rect 22094 3340 22100 3392
rect 22152 3380 22158 3392
rect 22922 3380 22928 3392
rect 22152 3352 22928 3380
rect 22152 3340 22158 3352
rect 22922 3340 22928 3352
rect 22980 3340 22986 3392
rect 23658 3340 23664 3392
rect 23716 3340 23722 3392
rect 23952 3389 23980 3420
rect 23937 3383 23995 3389
rect 23937 3349 23949 3383
rect 23983 3349 23995 3383
rect 23937 3343 23995 3349
rect 24121 3383 24179 3389
rect 24121 3349 24133 3383
rect 24167 3380 24179 3383
rect 25038 3380 25044 3392
rect 24167 3352 25044 3380
rect 24167 3349 24179 3352
rect 24121 3343 24179 3349
rect 25038 3340 25044 3352
rect 25096 3340 25102 3392
rect 552 3290 27416 3312
rect 552 3238 3756 3290
rect 3808 3238 3820 3290
rect 3872 3238 3884 3290
rect 3936 3238 3948 3290
rect 4000 3238 4012 3290
rect 4064 3238 10472 3290
rect 10524 3238 10536 3290
rect 10588 3238 10600 3290
rect 10652 3238 10664 3290
rect 10716 3238 10728 3290
rect 10780 3238 17188 3290
rect 17240 3238 17252 3290
rect 17304 3238 17316 3290
rect 17368 3238 17380 3290
rect 17432 3238 17444 3290
rect 17496 3238 23904 3290
rect 23956 3238 23968 3290
rect 24020 3238 24032 3290
rect 24084 3238 24096 3290
rect 24148 3238 24160 3290
rect 24212 3238 27416 3290
rect 552 3216 27416 3238
rect 4246 3136 4252 3188
rect 4304 3136 4310 3188
rect 4433 3179 4491 3185
rect 4433 3145 4445 3179
rect 4479 3176 4491 3179
rect 4706 3176 4712 3188
rect 4479 3148 4712 3176
rect 4479 3145 4491 3148
rect 4433 3139 4491 3145
rect 4706 3136 4712 3148
rect 4764 3136 4770 3188
rect 4798 3136 4804 3188
rect 4856 3176 4862 3188
rect 5166 3176 5172 3188
rect 4856 3148 5172 3176
rect 4856 3136 4862 3148
rect 5166 3136 5172 3148
rect 5224 3136 5230 3188
rect 6733 3179 6791 3185
rect 6733 3145 6745 3179
rect 6779 3176 6791 3179
rect 6822 3176 6828 3188
rect 6779 3148 6828 3176
rect 6779 3145 6791 3148
rect 6733 3139 6791 3145
rect 6822 3136 6828 3148
rect 6880 3136 6886 3188
rect 9950 3136 9956 3188
rect 10008 3176 10014 3188
rect 10413 3179 10471 3185
rect 10413 3176 10425 3179
rect 10008 3148 10425 3176
rect 10008 3136 10014 3148
rect 10413 3145 10425 3148
rect 10459 3176 10471 3179
rect 10962 3176 10968 3188
rect 10459 3148 10968 3176
rect 10459 3145 10471 3148
rect 10413 3139 10471 3145
rect 10962 3136 10968 3148
rect 11020 3136 11026 3188
rect 12805 3179 12863 3185
rect 12805 3145 12817 3179
rect 12851 3176 12863 3179
rect 13446 3176 13452 3188
rect 12851 3148 13452 3176
rect 12851 3145 12863 3148
rect 12805 3139 12863 3145
rect 13446 3136 13452 3148
rect 13504 3136 13510 3188
rect 13722 3136 13728 3188
rect 13780 3136 13786 3188
rect 14274 3136 14280 3188
rect 14332 3176 14338 3188
rect 14826 3176 14832 3188
rect 14332 3148 14832 3176
rect 14332 3136 14338 3148
rect 14826 3136 14832 3148
rect 14884 3136 14890 3188
rect 15105 3179 15163 3185
rect 15105 3145 15117 3179
rect 15151 3145 15163 3179
rect 15105 3139 15163 3145
rect 15289 3179 15347 3185
rect 15289 3145 15301 3179
rect 15335 3176 15347 3179
rect 15378 3176 15384 3188
rect 15335 3148 15384 3176
rect 15335 3145 15347 3148
rect 15289 3139 15347 3145
rect 3602 3068 3608 3120
rect 3660 3108 3666 3120
rect 4614 3108 4620 3120
rect 3660 3080 4620 3108
rect 3660 3068 3666 3080
rect 4614 3068 4620 3080
rect 4672 3108 4678 3120
rect 5537 3111 5595 3117
rect 5537 3108 5549 3111
rect 4672 3080 5549 3108
rect 4672 3068 4678 3080
rect 5537 3077 5549 3080
rect 5583 3077 5595 3111
rect 5537 3071 5595 3077
rect 6086 3068 6092 3120
rect 6144 3108 6150 3120
rect 8018 3108 8024 3120
rect 6144 3080 8024 3108
rect 6144 3068 6150 3080
rect 8018 3068 8024 3080
rect 8076 3068 8082 3120
rect 9585 3111 9643 3117
rect 9585 3077 9597 3111
rect 9631 3108 9643 3111
rect 10226 3108 10232 3120
rect 9631 3080 10232 3108
rect 9631 3077 9643 3080
rect 9585 3071 9643 3077
rect 10226 3068 10232 3080
rect 10284 3068 10290 3120
rect 12066 3068 12072 3120
rect 12124 3108 12130 3120
rect 14734 3108 14740 3120
rect 12124 3080 14740 3108
rect 12124 3068 12130 3080
rect 4525 3043 4583 3049
rect 4525 3040 4537 3043
rect 4080 3012 4537 3040
rect 3142 2932 3148 2984
rect 3200 2972 3206 2984
rect 3329 2975 3387 2981
rect 3329 2972 3341 2975
rect 3200 2944 3341 2972
rect 3200 2932 3206 2944
rect 3329 2941 3341 2944
rect 3375 2941 3387 2975
rect 3329 2935 3387 2941
rect 3510 2932 3516 2984
rect 3568 2932 3574 2984
rect 4080 2981 4108 3012
rect 4525 3009 4537 3012
rect 4571 3009 4583 3043
rect 6270 3040 6276 3052
rect 4525 3003 4583 3009
rect 4724 3012 6276 3040
rect 4724 2981 4752 3012
rect 4065 2975 4123 2981
rect 4065 2941 4077 2975
rect 4111 2941 4123 2975
rect 4065 2935 4123 2941
rect 4157 2975 4215 2981
rect 4157 2941 4169 2975
rect 4203 2941 4215 2975
rect 4157 2935 4215 2941
rect 4709 2975 4767 2981
rect 4709 2941 4721 2975
rect 4755 2941 4767 2975
rect 4709 2935 4767 2941
rect 3421 2907 3479 2913
rect 3421 2904 3433 2907
rect 2746 2876 3433 2904
rect 1210 2796 1216 2848
rect 1268 2836 1274 2848
rect 2746 2836 2774 2876
rect 3421 2873 3433 2876
rect 3467 2904 3479 2907
rect 4172 2904 4200 2935
rect 4798 2932 4804 2984
rect 4856 2932 4862 2984
rect 4982 2932 4988 2984
rect 5040 2932 5046 2984
rect 5184 2981 5212 3012
rect 6270 3000 6276 3012
rect 6328 3040 6334 3052
rect 11146 3040 11152 3052
rect 6328 3012 6776 3040
rect 6328 3000 6334 3012
rect 5077 2975 5135 2981
rect 5077 2941 5089 2975
rect 5123 2941 5135 2975
rect 5077 2935 5135 2941
rect 5169 2975 5227 2981
rect 5169 2941 5181 2975
rect 5215 2972 5227 2975
rect 5258 2972 5264 2984
rect 5215 2944 5264 2972
rect 5215 2941 5227 2944
rect 5169 2935 5227 2941
rect 3467 2876 4200 2904
rect 5092 2904 5120 2935
rect 5258 2932 5264 2944
rect 5316 2932 5322 2984
rect 5350 2932 5356 2984
rect 5408 2932 5414 2984
rect 5629 2975 5687 2981
rect 5629 2941 5641 2975
rect 5675 2972 5687 2975
rect 5905 2975 5963 2981
rect 5675 2944 5856 2972
rect 5675 2941 5687 2944
rect 5629 2935 5687 2941
rect 5534 2904 5540 2916
rect 5092 2876 5540 2904
rect 3467 2873 3479 2876
rect 3421 2867 3479 2873
rect 5534 2864 5540 2876
rect 5592 2864 5598 2916
rect 1268 2808 2774 2836
rect 5828 2836 5856 2944
rect 5905 2941 5917 2975
rect 5951 2972 5963 2975
rect 6454 2972 6460 2984
rect 6512 2981 6518 2984
rect 6748 2981 6776 3012
rect 9784 3012 11152 3040
rect 6512 2975 6545 2981
rect 5951 2944 6460 2972
rect 5951 2941 5963 2944
rect 5905 2935 5963 2941
rect 6454 2932 6460 2944
rect 6533 2941 6545 2975
rect 6512 2935 6545 2941
rect 6641 2975 6699 2981
rect 6641 2941 6653 2975
rect 6687 2941 6699 2975
rect 6641 2935 6699 2941
rect 6733 2975 6791 2981
rect 6733 2941 6745 2975
rect 6779 2941 6791 2975
rect 6733 2935 6791 2941
rect 6512 2932 6518 2935
rect 6656 2904 6684 2935
rect 6914 2932 6920 2984
rect 6972 2932 6978 2984
rect 7742 2932 7748 2984
rect 7800 2972 7806 2984
rect 7837 2975 7895 2981
rect 7837 2972 7849 2975
rect 7800 2944 7849 2972
rect 7800 2932 7806 2944
rect 7837 2941 7849 2944
rect 7883 2941 7895 2975
rect 7837 2935 7895 2941
rect 7926 2932 7932 2984
rect 7984 2972 7990 2984
rect 8021 2975 8079 2981
rect 8021 2972 8033 2975
rect 7984 2944 8033 2972
rect 7984 2932 7990 2944
rect 8021 2941 8033 2944
rect 8067 2941 8079 2975
rect 8021 2935 8079 2941
rect 8294 2932 8300 2984
rect 8352 2972 8358 2984
rect 8389 2975 8447 2981
rect 8389 2972 8401 2975
rect 8352 2944 8401 2972
rect 8352 2932 8358 2944
rect 8389 2941 8401 2944
rect 8435 2941 8447 2975
rect 8389 2935 8447 2941
rect 7760 2904 7788 2932
rect 9784 2913 9812 3012
rect 10612 2981 10640 3012
rect 11146 3000 11152 3012
rect 11204 3000 11210 3052
rect 12713 3043 12771 3049
rect 12713 3040 12725 3043
rect 11808 3012 12725 3040
rect 10505 2975 10563 2981
rect 10505 2941 10517 2975
rect 10551 2972 10563 2975
rect 10597 2975 10655 2981
rect 10597 2972 10609 2975
rect 10551 2944 10609 2972
rect 10551 2941 10563 2944
rect 10505 2935 10563 2941
rect 10597 2941 10609 2944
rect 10643 2941 10655 2975
rect 10597 2935 10655 2941
rect 10751 2975 10809 2981
rect 10751 2941 10763 2975
rect 10797 2972 10809 2975
rect 10962 2972 10968 2984
rect 10797 2944 10968 2972
rect 10797 2941 10809 2944
rect 10751 2935 10809 2941
rect 10962 2932 10968 2944
rect 11020 2932 11026 2984
rect 11330 2932 11336 2984
rect 11388 2972 11394 2984
rect 11517 2975 11575 2981
rect 11517 2972 11529 2975
rect 11388 2944 11529 2972
rect 11388 2932 11394 2944
rect 11517 2941 11529 2944
rect 11563 2941 11575 2975
rect 11517 2935 11575 2941
rect 11808 2916 11836 3012
rect 12713 3009 12725 3012
rect 12759 3040 12771 3043
rect 12759 3012 13032 3040
rect 12759 3009 12771 3012
rect 12713 3003 12771 3009
rect 11977 2975 12035 2981
rect 11977 2941 11989 2975
rect 12023 2972 12035 2975
rect 12066 2972 12072 2984
rect 12023 2944 12072 2972
rect 12023 2941 12035 2944
rect 11977 2935 12035 2941
rect 12066 2932 12072 2944
rect 12124 2972 12130 2984
rect 12437 2975 12495 2981
rect 12437 2972 12449 2975
rect 12124 2944 12449 2972
rect 12124 2932 12130 2944
rect 12437 2941 12449 2944
rect 12483 2941 12495 2975
rect 12437 2935 12495 2941
rect 12529 2975 12587 2981
rect 12529 2941 12541 2975
rect 12575 2972 12587 2975
rect 12802 2972 12808 2984
rect 12575 2944 12808 2972
rect 12575 2941 12587 2944
rect 12529 2935 12587 2941
rect 12802 2932 12808 2944
rect 12860 2932 12866 2984
rect 13004 2981 13032 3012
rect 12989 2975 13047 2981
rect 12989 2941 13001 2975
rect 13035 2941 13047 2975
rect 12989 2935 13047 2941
rect 13173 2975 13231 2981
rect 13173 2941 13185 2975
rect 13219 2941 13231 2975
rect 13173 2935 13231 2941
rect 13357 2975 13415 2981
rect 13357 2941 13369 2975
rect 13403 2941 13415 2975
rect 13357 2935 13415 2941
rect 6656 2876 7788 2904
rect 9769 2907 9827 2913
rect 6656 2836 6684 2876
rect 9769 2873 9781 2907
rect 9815 2873 9827 2907
rect 9769 2867 9827 2873
rect 9950 2864 9956 2916
rect 10008 2864 10014 2916
rect 10060 2876 11652 2904
rect 5828 2808 6684 2836
rect 1268 2796 1274 2808
rect 7926 2796 7932 2848
rect 7984 2796 7990 2848
rect 9674 2796 9680 2848
rect 9732 2836 9738 2848
rect 10060 2845 10088 2876
rect 11624 2848 11652 2876
rect 11790 2864 11796 2916
rect 11848 2864 11854 2916
rect 13188 2904 13216 2935
rect 12406 2876 13216 2904
rect 13372 2904 13400 2935
rect 13538 2932 13544 2984
rect 13596 2932 13602 2984
rect 13725 2975 13783 2981
rect 13725 2941 13737 2975
rect 13771 2941 13783 2975
rect 13924 2972 13952 3080
rect 14734 3068 14740 3080
rect 14792 3108 14798 3120
rect 15120 3108 15148 3139
rect 15378 3136 15384 3148
rect 15436 3136 15442 3188
rect 15749 3179 15807 3185
rect 15749 3145 15761 3179
rect 15795 3145 15807 3179
rect 15749 3139 15807 3145
rect 17773 3179 17831 3185
rect 17773 3145 17785 3179
rect 17819 3176 17831 3179
rect 18414 3176 18420 3188
rect 17819 3148 18420 3176
rect 17819 3145 17831 3148
rect 17773 3139 17831 3145
rect 15470 3108 15476 3120
rect 14792 3080 15476 3108
rect 14792 3068 14798 3080
rect 15470 3068 15476 3080
rect 15528 3108 15534 3120
rect 15764 3108 15792 3139
rect 18414 3136 18420 3148
rect 18472 3176 18478 3188
rect 18782 3176 18788 3188
rect 18472 3148 18788 3176
rect 18472 3136 18478 3148
rect 18782 3136 18788 3148
rect 18840 3136 18846 3188
rect 20070 3136 20076 3188
rect 20128 3176 20134 3188
rect 21818 3176 21824 3188
rect 20128 3148 21824 3176
rect 20128 3136 20134 3148
rect 21818 3136 21824 3148
rect 21876 3136 21882 3188
rect 21910 3136 21916 3188
rect 21968 3176 21974 3188
rect 22094 3176 22100 3188
rect 21968 3148 22100 3176
rect 21968 3136 21974 3148
rect 22094 3136 22100 3148
rect 22152 3136 22158 3188
rect 22281 3179 22339 3185
rect 22281 3145 22293 3179
rect 22327 3176 22339 3179
rect 22554 3176 22560 3188
rect 22327 3148 22560 3176
rect 22327 3145 22339 3148
rect 22281 3139 22339 3145
rect 22554 3136 22560 3148
rect 22612 3136 22618 3188
rect 22922 3136 22928 3188
rect 22980 3176 22986 3188
rect 23017 3179 23075 3185
rect 23017 3176 23029 3179
rect 22980 3148 23029 3176
rect 22980 3136 22986 3148
rect 23017 3145 23029 3148
rect 23063 3145 23075 3179
rect 23017 3139 23075 3145
rect 23124 3148 23336 3176
rect 15528 3080 15792 3108
rect 17405 3111 17463 3117
rect 15528 3068 15534 3080
rect 17405 3077 17417 3111
rect 17451 3108 17463 3111
rect 17678 3108 17684 3120
rect 17451 3080 17684 3108
rect 17451 3077 17463 3080
rect 17405 3071 17463 3077
rect 17678 3068 17684 3080
rect 17736 3068 17742 3120
rect 19981 3111 20039 3117
rect 19981 3077 19993 3111
rect 20027 3108 20039 3111
rect 20622 3108 20628 3120
rect 20027 3080 20628 3108
rect 20027 3077 20039 3080
rect 19981 3071 20039 3077
rect 20622 3068 20628 3080
rect 20680 3068 20686 3120
rect 20717 3111 20775 3117
rect 20717 3077 20729 3111
rect 20763 3108 20775 3111
rect 23124 3108 23152 3148
rect 20763 3080 23152 3108
rect 23201 3111 23259 3117
rect 20763 3077 20775 3080
rect 20717 3071 20775 3077
rect 23201 3077 23213 3111
rect 23247 3077 23259 3111
rect 23308 3108 23336 3148
rect 23382 3136 23388 3188
rect 23440 3176 23446 3188
rect 23845 3179 23903 3185
rect 23845 3176 23857 3179
rect 23440 3148 23857 3176
rect 23440 3136 23446 3148
rect 23845 3145 23857 3148
rect 23891 3145 23903 3179
rect 23845 3139 23903 3145
rect 23934 3136 23940 3188
rect 23992 3176 23998 3188
rect 24213 3179 24271 3185
rect 24213 3176 24225 3179
rect 23992 3148 24225 3176
rect 23992 3136 23998 3148
rect 24213 3145 24225 3148
rect 24259 3145 24271 3179
rect 24213 3139 24271 3145
rect 24302 3136 24308 3188
rect 24360 3136 24366 3188
rect 24762 3136 24768 3188
rect 24820 3136 24826 3188
rect 23308 3080 24440 3108
rect 23201 3071 23259 3077
rect 15378 3000 15384 3052
rect 15436 3000 15442 3052
rect 16390 3000 16396 3052
rect 16448 3000 16454 3052
rect 17957 3043 18015 3049
rect 17957 3009 17969 3043
rect 18003 3040 18015 3043
rect 18138 3040 18144 3052
rect 18003 3012 18144 3040
rect 18003 3009 18015 3012
rect 17957 3003 18015 3009
rect 18138 3000 18144 3012
rect 18196 3000 18202 3052
rect 18966 3040 18972 3052
rect 18708 3012 18972 3040
rect 14047 2975 14105 2981
rect 14047 2972 14059 2975
rect 13924 2944 14059 2972
rect 13725 2935 13783 2941
rect 14047 2941 14059 2944
rect 14093 2941 14105 2975
rect 14047 2935 14105 2941
rect 14185 2975 14243 2981
rect 14185 2941 14197 2975
rect 14231 2941 14243 2975
rect 14185 2935 14243 2941
rect 13630 2904 13636 2916
rect 13372 2876 13636 2904
rect 10045 2839 10103 2845
rect 10045 2836 10057 2839
rect 9732 2808 10057 2836
rect 9732 2796 9738 2808
rect 10045 2805 10057 2808
rect 10091 2805 10103 2839
rect 10045 2799 10103 2805
rect 10134 2796 10140 2848
rect 10192 2836 10198 2848
rect 10962 2836 10968 2848
rect 10192 2808 10968 2836
rect 10192 2796 10198 2808
rect 10962 2796 10968 2808
rect 11020 2796 11026 2848
rect 11606 2796 11612 2848
rect 11664 2836 11670 2848
rect 12406 2836 12434 2876
rect 13630 2864 13636 2876
rect 13688 2904 13694 2916
rect 13740 2904 13768 2935
rect 13817 2907 13875 2913
rect 13817 2904 13829 2907
rect 13688 2876 13829 2904
rect 13688 2864 13694 2876
rect 13817 2873 13829 2876
rect 13863 2873 13875 2907
rect 13817 2867 13875 2873
rect 13906 2864 13912 2916
rect 13964 2904 13970 2916
rect 14200 2904 14228 2935
rect 14274 2932 14280 2984
rect 14332 2932 14338 2984
rect 14458 2932 14464 2984
rect 14516 2972 14522 2984
rect 14737 2975 14795 2981
rect 14737 2972 14749 2975
rect 14516 2944 14749 2972
rect 14516 2932 14522 2944
rect 14737 2941 14749 2944
rect 14783 2941 14795 2975
rect 14737 2935 14795 2941
rect 15930 2932 15936 2984
rect 15988 2972 15994 2984
rect 16117 2975 16175 2981
rect 16117 2972 16129 2975
rect 15988 2944 16129 2972
rect 15988 2932 15994 2944
rect 16117 2941 16129 2944
rect 16163 2941 16175 2975
rect 16117 2935 16175 2941
rect 16669 2975 16727 2981
rect 16669 2941 16681 2975
rect 16715 2941 16727 2975
rect 16669 2935 16727 2941
rect 13964 2876 14228 2904
rect 13964 2864 13970 2876
rect 15102 2864 15108 2916
rect 15160 2904 15166 2916
rect 15749 2907 15807 2913
rect 15749 2904 15761 2907
rect 15160 2876 15761 2904
rect 15160 2864 15166 2876
rect 15749 2873 15761 2876
rect 15795 2873 15807 2907
rect 16684 2904 16712 2935
rect 16850 2932 16856 2984
rect 16908 2972 16914 2984
rect 18708 2981 18736 3012
rect 18966 3000 18972 3012
rect 19024 3040 19030 3052
rect 19613 3043 19671 3049
rect 19613 3040 19625 3043
rect 19024 3012 19625 3040
rect 19024 3000 19030 3012
rect 19613 3009 19625 3012
rect 19659 3009 19671 3043
rect 19613 3003 19671 3009
rect 20438 3000 20444 3052
rect 20496 3040 20502 3052
rect 20809 3043 20867 3049
rect 20809 3040 20821 3043
rect 20496 3012 20821 3040
rect 20496 3000 20502 3012
rect 20809 3009 20821 3012
rect 20855 3009 20867 3043
rect 20809 3003 20867 3009
rect 21560 3012 21772 3040
rect 17497 2975 17555 2981
rect 17497 2972 17509 2975
rect 16908 2944 17509 2972
rect 16908 2932 16914 2944
rect 17497 2941 17509 2944
rect 17543 2972 17555 2975
rect 18233 2975 18291 2981
rect 18233 2972 18245 2975
rect 17543 2944 18245 2972
rect 17543 2941 17555 2944
rect 17497 2935 17555 2941
rect 18233 2941 18245 2944
rect 18279 2972 18291 2975
rect 18693 2975 18751 2981
rect 18693 2972 18705 2975
rect 18279 2944 18705 2972
rect 18279 2941 18291 2944
rect 18233 2935 18291 2941
rect 18693 2941 18705 2944
rect 18739 2941 18751 2975
rect 18693 2935 18751 2941
rect 18782 2932 18788 2984
rect 18840 2972 18846 2984
rect 19150 2972 19156 2984
rect 18840 2944 19156 2972
rect 18840 2932 18846 2944
rect 19150 2932 19156 2944
rect 19208 2972 19214 2984
rect 19797 2975 19855 2981
rect 19797 2972 19809 2975
rect 19208 2944 19809 2972
rect 19208 2932 19214 2944
rect 19797 2941 19809 2944
rect 19843 2941 19855 2975
rect 19797 2935 19855 2941
rect 20162 2932 20168 2984
rect 20220 2972 20226 2984
rect 20533 2975 20591 2981
rect 20533 2972 20545 2975
rect 20220 2944 20545 2972
rect 20220 2932 20226 2944
rect 20533 2941 20545 2944
rect 20579 2972 20591 2975
rect 21560 2972 21588 3012
rect 20579 2944 21588 2972
rect 20579 2941 20591 2944
rect 20533 2935 20591 2941
rect 21634 2932 21640 2984
rect 21692 2932 21698 2984
rect 21744 2981 21772 3012
rect 22002 3000 22008 3052
rect 22060 3040 22066 3052
rect 22465 3043 22523 3049
rect 22060 3012 22324 3040
rect 22060 3000 22066 3012
rect 21730 2975 21788 2981
rect 21730 2941 21742 2975
rect 21776 2941 21788 2975
rect 21730 2935 21788 2941
rect 15749 2867 15807 2873
rect 16316 2876 16712 2904
rect 11664 2808 12434 2836
rect 11664 2796 11670 2808
rect 12710 2796 12716 2848
rect 12768 2796 12774 2848
rect 13265 2839 13323 2845
rect 13265 2805 13277 2839
rect 13311 2836 13323 2839
rect 14182 2836 14188 2848
rect 13311 2808 14188 2836
rect 13311 2805 13323 2808
rect 13265 2799 13323 2805
rect 14182 2796 14188 2808
rect 14240 2796 14246 2848
rect 15933 2839 15991 2845
rect 15933 2805 15945 2839
rect 15979 2836 15991 2839
rect 16114 2836 16120 2848
rect 15979 2808 16120 2836
rect 15979 2805 15991 2808
rect 15933 2799 15991 2805
rect 16114 2796 16120 2808
rect 16172 2796 16178 2848
rect 16316 2845 16344 2876
rect 18414 2864 18420 2916
rect 18472 2864 18478 2916
rect 19061 2907 19119 2913
rect 19061 2873 19073 2907
rect 19107 2873 19119 2907
rect 21744 2904 21772 2935
rect 21818 2932 21824 2984
rect 21876 2972 21882 2984
rect 22296 2981 22324 3012
rect 22465 3009 22477 3043
rect 22511 3040 22523 3043
rect 22830 3040 22836 3052
rect 22511 3012 22836 3040
rect 22511 3009 22523 3012
rect 22465 3003 22523 3009
rect 22830 3000 22836 3012
rect 22888 3000 22894 3052
rect 22097 2975 22155 2981
rect 22097 2972 22109 2975
rect 21876 2944 22109 2972
rect 21876 2932 21882 2944
rect 22097 2941 22109 2944
rect 22143 2941 22155 2975
rect 22097 2935 22155 2941
rect 22281 2975 22339 2981
rect 22281 2941 22293 2975
rect 22327 2972 22339 2975
rect 22373 2975 22431 2981
rect 22373 2972 22385 2975
rect 22327 2944 22385 2972
rect 22327 2941 22339 2944
rect 22281 2935 22339 2941
rect 22373 2941 22385 2944
rect 22419 2941 22431 2975
rect 22557 2975 22615 2981
rect 22557 2972 22569 2975
rect 22373 2935 22431 2941
rect 22480 2944 22569 2972
rect 21910 2904 21916 2916
rect 21744 2876 21916 2904
rect 19061 2867 19119 2873
rect 16301 2839 16359 2845
rect 16301 2805 16313 2839
rect 16347 2805 16359 2839
rect 16301 2799 16359 2805
rect 18046 2796 18052 2848
rect 18104 2796 18110 2848
rect 18782 2796 18788 2848
rect 18840 2836 18846 2848
rect 19076 2836 19104 2867
rect 21910 2864 21916 2876
rect 21968 2864 21974 2916
rect 20346 2836 20352 2848
rect 18840 2808 20352 2836
rect 18840 2796 18846 2808
rect 20346 2796 20352 2808
rect 20404 2836 20410 2848
rect 22480 2836 22508 2944
rect 22557 2941 22569 2944
rect 22603 2972 22615 2975
rect 22649 2975 22707 2981
rect 22649 2972 22661 2975
rect 22603 2944 22661 2972
rect 22603 2941 22615 2944
rect 22557 2935 22615 2941
rect 22649 2941 22661 2944
rect 22695 2941 22707 2975
rect 23216 2972 23244 3071
rect 24412 3049 24440 3080
rect 24397 3043 24455 3049
rect 24397 3009 24409 3043
rect 24443 3009 24455 3043
rect 25314 3040 25320 3052
rect 24397 3003 24455 3009
rect 24504 3012 25320 3040
rect 23477 2975 23535 2981
rect 23477 2972 23489 2975
rect 23216 2944 23489 2972
rect 22649 2935 22707 2941
rect 23477 2941 23489 2944
rect 23523 2941 23535 2975
rect 23477 2935 23535 2941
rect 23658 2932 23664 2984
rect 23716 2972 23722 2984
rect 23845 2975 23903 2981
rect 23845 2972 23857 2975
rect 23716 2944 23857 2972
rect 23716 2932 23722 2944
rect 23845 2941 23857 2944
rect 23891 2941 23903 2975
rect 23845 2935 23903 2941
rect 24029 2975 24087 2981
rect 24029 2941 24041 2975
rect 24075 2941 24087 2975
rect 24029 2935 24087 2941
rect 23017 2907 23075 2913
rect 23017 2873 23029 2907
rect 23063 2904 23075 2907
rect 23106 2904 23112 2916
rect 23063 2876 23112 2904
rect 23063 2873 23075 2876
rect 23017 2867 23075 2873
rect 23106 2864 23112 2876
rect 23164 2864 23170 2916
rect 24044 2904 24072 2935
rect 24210 2932 24216 2984
rect 24268 2972 24274 2984
rect 24305 2975 24363 2981
rect 24305 2972 24317 2975
rect 24268 2944 24317 2972
rect 24268 2932 24274 2944
rect 24305 2941 24317 2944
rect 24351 2941 24363 2975
rect 24305 2935 24363 2941
rect 24504 2904 24532 3012
rect 25314 3000 25320 3012
rect 25372 3000 25378 3052
rect 24949 2975 25007 2981
rect 24949 2972 24961 2975
rect 23676 2876 24532 2904
rect 24688 2944 24961 2972
rect 23676 2845 23704 2876
rect 24688 2845 24716 2944
rect 24949 2941 24961 2944
rect 24995 2941 25007 2975
rect 24949 2935 25007 2941
rect 25038 2932 25044 2984
rect 25096 2932 25102 2984
rect 20404 2808 22508 2836
rect 23661 2839 23719 2845
rect 20404 2796 20410 2808
rect 23661 2805 23673 2839
rect 23707 2805 23719 2839
rect 23661 2799 23719 2805
rect 24673 2839 24731 2845
rect 24673 2805 24685 2839
rect 24719 2805 24731 2839
rect 24673 2799 24731 2805
rect 25130 2796 25136 2848
rect 25188 2836 25194 2848
rect 25225 2839 25283 2845
rect 25225 2836 25237 2839
rect 25188 2808 25237 2836
rect 25188 2796 25194 2808
rect 25225 2805 25237 2808
rect 25271 2805 25283 2839
rect 25225 2799 25283 2805
rect 552 2746 27576 2768
rect 552 2694 7114 2746
rect 7166 2694 7178 2746
rect 7230 2694 7242 2746
rect 7294 2694 7306 2746
rect 7358 2694 7370 2746
rect 7422 2694 13830 2746
rect 13882 2694 13894 2746
rect 13946 2694 13958 2746
rect 14010 2694 14022 2746
rect 14074 2694 14086 2746
rect 14138 2694 20546 2746
rect 20598 2694 20610 2746
rect 20662 2694 20674 2746
rect 20726 2694 20738 2746
rect 20790 2694 20802 2746
rect 20854 2694 27262 2746
rect 27314 2694 27326 2746
rect 27378 2694 27390 2746
rect 27442 2694 27454 2746
rect 27506 2694 27518 2746
rect 27570 2694 27576 2746
rect 552 2672 27576 2694
rect 4798 2592 4804 2644
rect 4856 2632 4862 2644
rect 4893 2635 4951 2641
rect 4893 2632 4905 2635
rect 4856 2604 4905 2632
rect 4856 2592 4862 2604
rect 4893 2601 4905 2604
rect 4939 2601 4951 2635
rect 7929 2635 7987 2641
rect 4893 2595 4951 2601
rect 5000 2604 6960 2632
rect 3605 2567 3663 2573
rect 3605 2564 3617 2567
rect 2746 2536 3617 2564
rect 2593 2499 2651 2505
rect 2593 2465 2605 2499
rect 2639 2496 2651 2499
rect 2746 2496 2774 2536
rect 3605 2533 3617 2536
rect 3651 2533 3663 2567
rect 3605 2527 3663 2533
rect 4540 2536 4844 2564
rect 4540 2508 4568 2536
rect 2639 2468 2774 2496
rect 2639 2465 2651 2468
rect 2593 2459 2651 2465
rect 3418 2456 3424 2508
rect 3476 2456 3482 2508
rect 3513 2499 3571 2505
rect 3513 2465 3525 2499
rect 3559 2465 3571 2499
rect 3513 2459 3571 2465
rect 3697 2499 3755 2505
rect 3697 2465 3709 2499
rect 3743 2496 3755 2499
rect 4062 2496 4068 2508
rect 3743 2468 4068 2496
rect 3743 2465 3755 2468
rect 3697 2459 3755 2465
rect 2225 2431 2283 2437
rect 2225 2397 2237 2431
rect 2271 2428 2283 2431
rect 2317 2431 2375 2437
rect 2317 2428 2329 2431
rect 2271 2400 2329 2428
rect 2271 2397 2283 2400
rect 2225 2391 2283 2397
rect 2317 2397 2329 2400
rect 2363 2397 2375 2431
rect 2317 2391 2375 2397
rect 3142 2388 3148 2440
rect 3200 2428 3206 2440
rect 3528 2428 3556 2459
rect 4062 2456 4068 2468
rect 4120 2456 4126 2508
rect 4522 2456 4528 2508
rect 4580 2456 4586 2508
rect 4706 2456 4712 2508
rect 4764 2456 4770 2508
rect 4724 2428 4752 2456
rect 3200 2400 4752 2428
rect 4816 2428 4844 2536
rect 4890 2456 4896 2508
rect 4948 2496 4954 2508
rect 5000 2505 5028 2604
rect 6932 2576 6960 2604
rect 7929 2601 7941 2635
rect 7975 2632 7987 2635
rect 8110 2632 8116 2644
rect 7975 2604 8116 2632
rect 7975 2601 7987 2604
rect 7929 2595 7987 2601
rect 8110 2592 8116 2604
rect 8168 2592 8174 2644
rect 12894 2632 12900 2644
rect 11164 2604 12900 2632
rect 6086 2564 6092 2576
rect 5184 2536 6092 2564
rect 4985 2499 5043 2505
rect 4985 2496 4997 2499
rect 4948 2468 4997 2496
rect 4948 2456 4954 2468
rect 4985 2465 4997 2468
rect 5031 2465 5043 2499
rect 4985 2459 5043 2465
rect 5184 2428 5212 2536
rect 6086 2524 6092 2536
rect 6144 2524 6150 2576
rect 6822 2524 6828 2576
rect 6880 2524 6886 2576
rect 6914 2524 6920 2576
rect 6972 2524 6978 2576
rect 8128 2564 8156 2592
rect 7484 2536 7788 2564
rect 8128 2536 8432 2564
rect 5258 2456 5264 2508
rect 5316 2496 5322 2508
rect 5445 2499 5503 2505
rect 5445 2496 5457 2499
rect 5316 2468 5457 2496
rect 5316 2456 5322 2468
rect 5445 2465 5457 2468
rect 5491 2465 5503 2499
rect 5445 2459 5503 2465
rect 5629 2499 5687 2505
rect 5629 2465 5641 2499
rect 5675 2465 5687 2499
rect 5629 2459 5687 2465
rect 5813 2499 5871 2505
rect 5813 2465 5825 2499
rect 5859 2496 5871 2499
rect 6178 2496 6184 2508
rect 5859 2468 6184 2496
rect 5859 2465 5871 2468
rect 5813 2459 5871 2465
rect 4816 2400 5212 2428
rect 5644 2428 5672 2459
rect 6178 2456 6184 2468
rect 6236 2456 6242 2508
rect 6641 2499 6699 2505
rect 6641 2465 6653 2499
rect 6687 2496 6699 2499
rect 6840 2496 6868 2524
rect 6687 2468 6868 2496
rect 6932 2496 6960 2524
rect 7484 2505 7512 2536
rect 7285 2499 7343 2505
rect 7285 2496 7297 2499
rect 6932 2468 7297 2496
rect 6687 2465 6699 2468
rect 6641 2459 6699 2465
rect 7285 2465 7297 2468
rect 7331 2465 7343 2499
rect 7285 2459 7343 2465
rect 7469 2499 7527 2505
rect 7469 2465 7481 2499
rect 7515 2465 7527 2499
rect 7469 2459 7527 2465
rect 7558 2456 7564 2508
rect 7616 2456 7622 2508
rect 7760 2505 7788 2536
rect 7745 2499 7803 2505
rect 7745 2465 7757 2499
rect 7791 2496 7803 2499
rect 7837 2499 7895 2505
rect 7837 2496 7849 2499
rect 7791 2468 7849 2496
rect 7791 2465 7803 2468
rect 7745 2459 7803 2465
rect 7837 2465 7849 2468
rect 7883 2496 7895 2499
rect 7926 2496 7932 2508
rect 7883 2468 7932 2496
rect 7883 2465 7895 2468
rect 7837 2459 7895 2465
rect 7926 2456 7932 2468
rect 7984 2456 7990 2508
rect 8018 2456 8024 2508
rect 8076 2456 8082 2508
rect 8113 2499 8171 2505
rect 8113 2465 8125 2499
rect 8159 2496 8171 2499
rect 8294 2496 8300 2508
rect 8159 2468 8300 2496
rect 8159 2465 8171 2468
rect 8113 2459 8171 2465
rect 8294 2456 8300 2468
rect 8352 2456 8358 2508
rect 8404 2505 8432 2536
rect 9968 2536 10456 2564
rect 8389 2499 8447 2505
rect 8389 2465 8401 2499
rect 8435 2465 8447 2499
rect 8389 2459 8447 2465
rect 9217 2499 9275 2505
rect 9217 2465 9229 2499
rect 9263 2496 9275 2499
rect 9490 2496 9496 2508
rect 9263 2468 9496 2496
rect 9263 2465 9275 2468
rect 9217 2459 9275 2465
rect 9490 2456 9496 2468
rect 9548 2456 9554 2508
rect 9674 2456 9680 2508
rect 9732 2456 9738 2508
rect 9968 2505 9996 2536
rect 9861 2499 9919 2505
rect 9861 2465 9873 2499
rect 9907 2496 9919 2499
rect 9953 2499 10011 2505
rect 9953 2496 9965 2499
rect 9907 2468 9965 2496
rect 9907 2465 9919 2468
rect 9861 2459 9919 2465
rect 9953 2465 9965 2468
rect 9999 2465 10011 2499
rect 9953 2459 10011 2465
rect 10134 2456 10140 2508
rect 10192 2456 10198 2508
rect 10226 2456 10232 2508
rect 10284 2456 10290 2508
rect 10428 2505 10456 2536
rect 10413 2499 10471 2505
rect 10413 2465 10425 2499
rect 10459 2496 10471 2499
rect 10965 2499 11023 2505
rect 10965 2496 10977 2499
rect 10459 2468 10977 2496
rect 10459 2465 10471 2468
rect 10413 2459 10471 2465
rect 10965 2465 10977 2468
rect 11011 2465 11023 2499
rect 10965 2459 11023 2465
rect 5994 2428 6000 2440
rect 5644 2400 6000 2428
rect 3200 2388 3206 2400
rect 4062 2320 4068 2372
rect 4120 2360 4126 2372
rect 5644 2360 5672 2400
rect 5994 2388 6000 2400
rect 6052 2388 6058 2440
rect 6914 2388 6920 2440
rect 6972 2388 6978 2440
rect 7006 2388 7012 2440
rect 7064 2428 7070 2440
rect 7377 2431 7435 2437
rect 7377 2428 7389 2431
rect 7064 2400 7389 2428
rect 7064 2388 7070 2400
rect 7377 2397 7389 2400
rect 7423 2397 7435 2431
rect 7377 2391 7435 2397
rect 4120 2332 5672 2360
rect 10244 2360 10272 2456
rect 10980 2428 11008 2459
rect 11054 2456 11060 2508
rect 11112 2496 11118 2508
rect 11164 2505 11192 2604
rect 12894 2592 12900 2604
rect 12952 2632 12958 2644
rect 12952 2604 13952 2632
rect 12952 2592 12958 2604
rect 11532 2536 11836 2564
rect 11532 2505 11560 2536
rect 11808 2508 11836 2536
rect 11149 2499 11207 2505
rect 11149 2496 11161 2499
rect 11112 2468 11161 2496
rect 11112 2456 11118 2468
rect 11149 2465 11161 2468
rect 11195 2465 11207 2499
rect 11149 2459 11207 2465
rect 11333 2499 11391 2505
rect 11333 2465 11345 2499
rect 11379 2465 11391 2499
rect 11333 2459 11391 2465
rect 11517 2499 11575 2505
rect 11517 2465 11529 2499
rect 11563 2465 11575 2499
rect 11517 2459 11575 2465
rect 11238 2428 11244 2440
rect 10980 2400 11244 2428
rect 11238 2388 11244 2400
rect 11296 2388 11302 2440
rect 11348 2428 11376 2459
rect 11606 2456 11612 2508
rect 11664 2456 11670 2508
rect 11790 2456 11796 2508
rect 11848 2456 11854 2508
rect 13924 2505 13952 2604
rect 15930 2592 15936 2644
rect 15988 2592 15994 2644
rect 18138 2592 18144 2644
rect 18196 2632 18202 2644
rect 20070 2632 20076 2644
rect 18196 2604 20076 2632
rect 18196 2592 18202 2604
rect 20070 2592 20076 2604
rect 20128 2592 20134 2644
rect 23017 2635 23075 2641
rect 23017 2601 23029 2635
rect 23063 2632 23075 2635
rect 23106 2632 23112 2644
rect 23063 2604 23112 2632
rect 23063 2601 23075 2604
rect 23017 2595 23075 2601
rect 23106 2592 23112 2604
rect 23164 2592 23170 2644
rect 23201 2635 23259 2641
rect 23201 2601 23213 2635
rect 23247 2601 23259 2635
rect 23201 2595 23259 2601
rect 23753 2635 23811 2641
rect 23753 2601 23765 2635
rect 23799 2632 23811 2635
rect 24302 2632 24308 2644
rect 23799 2604 24308 2632
rect 23799 2601 23811 2604
rect 23753 2595 23811 2601
rect 14001 2567 14059 2573
rect 14001 2533 14013 2567
rect 14047 2564 14059 2567
rect 18046 2564 18052 2576
rect 14047 2536 15608 2564
rect 14047 2533 14059 2536
rect 14001 2527 14059 2533
rect 13909 2499 13967 2505
rect 13909 2465 13921 2499
rect 13955 2465 13967 2499
rect 13909 2459 13967 2465
rect 14093 2499 14151 2505
rect 14093 2465 14105 2499
rect 14139 2496 14151 2499
rect 14274 2496 14280 2508
rect 14139 2468 14280 2496
rect 14139 2465 14151 2468
rect 14093 2459 14151 2465
rect 13538 2428 13544 2440
rect 11348 2400 13544 2428
rect 11348 2360 11376 2400
rect 13538 2388 13544 2400
rect 13596 2388 13602 2440
rect 13630 2388 13636 2440
rect 13688 2428 13694 2440
rect 14108 2428 14136 2459
rect 14274 2456 14280 2468
rect 14332 2456 14338 2508
rect 15470 2456 15476 2508
rect 15528 2496 15534 2508
rect 15580 2505 15608 2536
rect 17696 2536 18052 2564
rect 15565 2499 15623 2505
rect 15565 2496 15577 2499
rect 15528 2468 15577 2496
rect 15528 2456 15534 2468
rect 15565 2465 15577 2468
rect 15611 2465 15623 2499
rect 15565 2459 15623 2465
rect 16114 2456 16120 2508
rect 16172 2456 16178 2508
rect 16298 2456 16304 2508
rect 16356 2496 16362 2508
rect 17696 2505 17724 2536
rect 18046 2524 18052 2536
rect 18104 2524 18110 2576
rect 20438 2564 20444 2576
rect 19996 2536 20444 2564
rect 16393 2499 16451 2505
rect 16393 2496 16405 2499
rect 16356 2468 16405 2496
rect 16356 2456 16362 2468
rect 16393 2465 16405 2468
rect 16439 2465 16451 2499
rect 16393 2459 16451 2465
rect 17681 2499 17739 2505
rect 17681 2465 17693 2499
rect 17727 2465 17739 2499
rect 17681 2459 17739 2465
rect 17865 2499 17923 2505
rect 17865 2465 17877 2499
rect 17911 2496 17923 2499
rect 17954 2496 17960 2508
rect 17911 2468 17960 2496
rect 17911 2465 17923 2468
rect 17865 2459 17923 2465
rect 17954 2456 17960 2468
rect 18012 2456 18018 2508
rect 18138 2456 18144 2508
rect 18196 2456 18202 2508
rect 18598 2456 18604 2508
rect 18656 2456 18662 2508
rect 18782 2456 18788 2508
rect 18840 2456 18846 2508
rect 18877 2499 18935 2505
rect 18877 2465 18889 2499
rect 18923 2465 18935 2499
rect 18877 2459 18935 2465
rect 13688 2400 14136 2428
rect 15657 2431 15715 2437
rect 13688 2388 13694 2400
rect 15657 2397 15669 2431
rect 15703 2397 15715 2431
rect 18616 2428 18644 2456
rect 18892 2428 18920 2459
rect 18966 2456 18972 2508
rect 19024 2496 19030 2508
rect 19996 2505 20024 2536
rect 19061 2499 19119 2505
rect 19061 2496 19073 2499
rect 19024 2468 19073 2496
rect 19024 2456 19030 2468
rect 19061 2465 19073 2468
rect 19107 2465 19119 2499
rect 19061 2459 19119 2465
rect 19797 2499 19855 2505
rect 19797 2465 19809 2499
rect 19843 2465 19855 2499
rect 19797 2459 19855 2465
rect 19981 2499 20039 2505
rect 19981 2465 19993 2499
rect 20027 2465 20039 2499
rect 19981 2459 20039 2465
rect 18616 2400 18920 2428
rect 15657 2391 15715 2397
rect 10244 2332 11376 2360
rect 4120 2320 4126 2332
rect 12710 2320 12716 2372
rect 12768 2360 12774 2372
rect 15672 2360 15700 2391
rect 12768 2332 15700 2360
rect 12768 2320 12774 2332
rect 18046 2320 18052 2372
rect 18104 2360 18110 2372
rect 19812 2360 19840 2459
rect 20070 2456 20076 2508
rect 20128 2456 20134 2508
rect 20272 2505 20300 2536
rect 20438 2524 20444 2536
rect 20496 2564 20502 2576
rect 20496 2536 20760 2564
rect 20496 2524 20502 2536
rect 20732 2508 20760 2536
rect 22112 2536 22416 2564
rect 20257 2499 20315 2505
rect 20257 2465 20269 2499
rect 20303 2465 20315 2499
rect 20257 2459 20315 2465
rect 20346 2456 20352 2508
rect 20404 2496 20410 2508
rect 20625 2499 20683 2505
rect 20625 2496 20637 2499
rect 20404 2468 20637 2496
rect 20404 2456 20410 2468
rect 20625 2465 20637 2468
rect 20671 2465 20683 2499
rect 20625 2459 20683 2465
rect 20714 2456 20720 2508
rect 20772 2496 20778 2508
rect 20809 2499 20867 2505
rect 20809 2496 20821 2499
rect 20772 2468 20821 2496
rect 20772 2456 20778 2468
rect 20809 2465 20821 2468
rect 20855 2465 20867 2499
rect 20809 2459 20867 2465
rect 21913 2499 21971 2505
rect 21913 2465 21925 2499
rect 21959 2465 21971 2499
rect 21913 2459 21971 2465
rect 21928 2428 21956 2459
rect 22002 2456 22008 2508
rect 22060 2496 22066 2508
rect 22112 2505 22140 2536
rect 22097 2499 22155 2505
rect 22097 2496 22109 2499
rect 22060 2468 22109 2496
rect 22060 2456 22066 2468
rect 22097 2465 22109 2468
rect 22143 2465 22155 2499
rect 22097 2459 22155 2465
rect 22189 2499 22247 2505
rect 22189 2465 22201 2499
rect 22235 2496 22247 2499
rect 22278 2496 22284 2508
rect 22235 2468 22284 2496
rect 22235 2465 22247 2468
rect 22189 2459 22247 2465
rect 22278 2456 22284 2468
rect 22336 2456 22342 2508
rect 22388 2505 22416 2536
rect 22373 2499 22431 2505
rect 22373 2465 22385 2499
rect 22419 2465 22431 2499
rect 23216 2496 23244 2595
rect 24302 2592 24308 2604
rect 24360 2592 24366 2644
rect 23569 2499 23627 2505
rect 23569 2496 23581 2499
rect 23216 2468 23581 2496
rect 22373 2459 22431 2465
rect 23569 2465 23581 2468
rect 23615 2465 23627 2499
rect 23569 2459 23627 2465
rect 22649 2431 22707 2437
rect 22649 2428 22661 2431
rect 21928 2400 22661 2428
rect 21928 2360 21956 2400
rect 22649 2397 22661 2400
rect 22695 2397 22707 2431
rect 22649 2391 22707 2397
rect 18104 2332 21956 2360
rect 22097 2363 22155 2369
rect 18104 2320 18110 2332
rect 22097 2329 22109 2363
rect 22143 2360 22155 2363
rect 22186 2360 22192 2372
rect 22143 2332 22192 2360
rect 22143 2329 22155 2332
rect 22097 2323 22155 2329
rect 22186 2320 22192 2332
rect 22244 2320 22250 2372
rect 22373 2363 22431 2369
rect 22373 2329 22385 2363
rect 22419 2360 22431 2363
rect 23658 2360 23664 2372
rect 22419 2332 23664 2360
rect 22419 2329 22431 2332
rect 22373 2323 22431 2329
rect 23658 2320 23664 2332
rect 23716 2360 23722 2372
rect 24210 2360 24216 2372
rect 23716 2332 24216 2360
rect 23716 2320 23722 2332
rect 24210 2320 24216 2332
rect 24268 2320 24274 2372
rect 4154 2252 4160 2304
rect 4212 2292 4218 2304
rect 4525 2295 4583 2301
rect 4525 2292 4537 2295
rect 4212 2264 4537 2292
rect 4212 2252 4218 2264
rect 4525 2261 4537 2264
rect 4571 2292 4583 2295
rect 4982 2292 4988 2304
rect 4571 2264 4988 2292
rect 4571 2261 4583 2264
rect 4525 2255 4583 2261
rect 4982 2252 4988 2264
rect 5040 2252 5046 2304
rect 5534 2252 5540 2304
rect 5592 2292 5598 2304
rect 5629 2295 5687 2301
rect 5629 2292 5641 2295
rect 5592 2264 5641 2292
rect 5592 2252 5598 2264
rect 5629 2261 5641 2264
rect 5675 2292 5687 2295
rect 5902 2292 5908 2304
rect 5675 2264 5908 2292
rect 5675 2261 5687 2264
rect 5629 2255 5687 2261
rect 5902 2252 5908 2264
rect 5960 2252 5966 2304
rect 6270 2252 6276 2304
rect 6328 2292 6334 2304
rect 7009 2295 7067 2301
rect 7009 2292 7021 2295
rect 6328 2264 7021 2292
rect 6328 2252 6334 2264
rect 7009 2261 7021 2264
rect 7055 2261 7067 2295
rect 7009 2255 7067 2261
rect 7745 2295 7803 2301
rect 7745 2261 7757 2295
rect 7791 2292 7803 2295
rect 8202 2292 8208 2304
rect 7791 2264 8208 2292
rect 7791 2261 7803 2264
rect 7745 2255 7803 2261
rect 8202 2252 8208 2264
rect 8260 2252 8266 2304
rect 9674 2252 9680 2304
rect 9732 2252 9738 2304
rect 9950 2252 9956 2304
rect 10008 2292 10014 2304
rect 10137 2295 10195 2301
rect 10137 2292 10149 2295
rect 10008 2264 10149 2292
rect 10008 2252 10014 2264
rect 10137 2261 10149 2264
rect 10183 2261 10195 2295
rect 10137 2255 10195 2261
rect 10226 2252 10232 2304
rect 10284 2252 10290 2304
rect 11149 2295 11207 2301
rect 11149 2261 11161 2295
rect 11195 2292 11207 2295
rect 11238 2292 11244 2304
rect 11195 2264 11244 2292
rect 11195 2261 11207 2264
rect 11149 2255 11207 2261
rect 11238 2252 11244 2264
rect 11296 2252 11302 2304
rect 11330 2252 11336 2304
rect 11388 2292 11394 2304
rect 11517 2295 11575 2301
rect 11517 2292 11529 2295
rect 11388 2264 11529 2292
rect 11388 2252 11394 2264
rect 11517 2261 11529 2264
rect 11563 2261 11575 2295
rect 11517 2255 11575 2261
rect 11793 2295 11851 2301
rect 11793 2261 11805 2295
rect 11839 2292 11851 2295
rect 11882 2292 11888 2304
rect 11839 2264 11888 2292
rect 11839 2261 11851 2264
rect 11793 2255 11851 2261
rect 11882 2252 11888 2264
rect 11940 2252 11946 2304
rect 12250 2252 12256 2304
rect 12308 2292 12314 2304
rect 12345 2295 12403 2301
rect 12345 2292 12357 2295
rect 12308 2264 12357 2292
rect 12308 2252 12314 2264
rect 12345 2261 12357 2264
rect 12391 2261 12403 2295
rect 12345 2255 12403 2261
rect 15194 2252 15200 2304
rect 15252 2292 15258 2304
rect 15289 2295 15347 2301
rect 15289 2292 15301 2295
rect 15252 2264 15301 2292
rect 15252 2252 15258 2264
rect 15289 2261 15301 2264
rect 15335 2261 15347 2295
rect 15289 2255 15347 2261
rect 15749 2295 15807 2301
rect 15749 2261 15761 2295
rect 15795 2292 15807 2295
rect 16298 2292 16304 2304
rect 15795 2264 16304 2292
rect 15795 2261 15807 2264
rect 15749 2255 15807 2261
rect 16298 2252 16304 2264
rect 16356 2252 16362 2304
rect 16574 2252 16580 2304
rect 16632 2252 16638 2304
rect 17678 2252 17684 2304
rect 17736 2252 17742 2304
rect 18141 2295 18199 2301
rect 18141 2261 18153 2295
rect 18187 2292 18199 2295
rect 18506 2292 18512 2304
rect 18187 2264 18512 2292
rect 18187 2261 18199 2264
rect 18141 2255 18199 2261
rect 18506 2252 18512 2264
rect 18564 2252 18570 2304
rect 18785 2295 18843 2301
rect 18785 2261 18797 2295
rect 18831 2292 18843 2295
rect 18966 2292 18972 2304
rect 18831 2264 18972 2292
rect 18831 2261 18843 2264
rect 18785 2255 18843 2261
rect 18966 2252 18972 2264
rect 19024 2252 19030 2304
rect 19058 2252 19064 2304
rect 19116 2252 19122 2304
rect 19794 2252 19800 2304
rect 19852 2292 19858 2304
rect 19981 2295 20039 2301
rect 19981 2292 19993 2295
rect 19852 2264 19993 2292
rect 19852 2252 19858 2264
rect 19981 2261 19993 2264
rect 20027 2261 20039 2295
rect 19981 2255 20039 2261
rect 20254 2252 20260 2304
rect 20312 2252 20318 2304
rect 20809 2295 20867 2301
rect 20809 2261 20821 2295
rect 20855 2292 20867 2295
rect 21542 2292 21548 2304
rect 20855 2264 21548 2292
rect 20855 2261 20867 2264
rect 20809 2255 20867 2261
rect 21542 2252 21548 2264
rect 21600 2252 21606 2304
rect 23014 2252 23020 2304
rect 23072 2252 23078 2304
rect 552 2202 27416 2224
rect 552 2150 3756 2202
rect 3808 2150 3820 2202
rect 3872 2150 3884 2202
rect 3936 2150 3948 2202
rect 4000 2150 4012 2202
rect 4064 2150 10472 2202
rect 10524 2150 10536 2202
rect 10588 2150 10600 2202
rect 10652 2150 10664 2202
rect 10716 2150 10728 2202
rect 10780 2150 17188 2202
rect 17240 2150 17252 2202
rect 17304 2150 17316 2202
rect 17368 2150 17380 2202
rect 17432 2150 17444 2202
rect 17496 2150 23904 2202
rect 23956 2150 23968 2202
rect 24020 2150 24032 2202
rect 24084 2150 24096 2202
rect 24148 2150 24160 2202
rect 24212 2150 27416 2202
rect 552 2128 27416 2150
rect 5994 2088 6000 2100
rect 4816 2060 6000 2088
rect 4706 1952 4712 1964
rect 2792 1924 4712 1952
rect 934 1844 940 1896
rect 992 1844 998 1896
rect 1213 1887 1271 1893
rect 1213 1853 1225 1887
rect 1259 1853 1271 1887
rect 1213 1847 1271 1853
rect 1228 1816 1256 1847
rect 1762 1844 1768 1896
rect 1820 1884 1826 1896
rect 2041 1887 2099 1893
rect 2041 1884 2053 1887
rect 1820 1856 2053 1884
rect 1820 1844 1826 1856
rect 2041 1853 2053 1856
rect 2087 1853 2099 1887
rect 2041 1847 2099 1853
rect 2130 1844 2136 1896
rect 2188 1844 2194 1896
rect 2792 1893 2820 1924
rect 2777 1887 2835 1893
rect 2777 1853 2789 1887
rect 2823 1853 2835 1887
rect 2777 1847 2835 1853
rect 2961 1887 3019 1893
rect 2961 1853 2973 1887
rect 3007 1884 3019 1887
rect 3142 1884 3148 1896
rect 3007 1856 3148 1884
rect 3007 1853 3019 1856
rect 2961 1847 3019 1853
rect 3142 1844 3148 1856
rect 3200 1844 3206 1896
rect 3252 1893 3280 1924
rect 4706 1912 4712 1924
rect 4764 1912 4770 1964
rect 3237 1887 3295 1893
rect 3237 1853 3249 1887
rect 3283 1853 3295 1887
rect 3237 1847 3295 1853
rect 3421 1887 3479 1893
rect 3421 1853 3433 1887
rect 3467 1853 3479 1887
rect 3421 1847 3479 1853
rect 2869 1819 2927 1825
rect 2869 1816 2881 1819
rect 1228 1788 2881 1816
rect 2869 1785 2881 1788
rect 2915 1785 2927 1819
rect 3436 1816 3464 1847
rect 3510 1844 3516 1896
rect 3568 1844 3574 1896
rect 3697 1887 3755 1893
rect 3697 1853 3709 1887
rect 3743 1853 3755 1887
rect 3697 1847 3755 1853
rect 3712 1816 3740 1847
rect 4246 1844 4252 1896
rect 4304 1844 4310 1896
rect 4341 1887 4399 1893
rect 4341 1853 4353 1887
rect 4387 1853 4399 1887
rect 4341 1847 4399 1853
rect 4356 1816 4384 1847
rect 4522 1844 4528 1896
rect 4580 1844 4586 1896
rect 4614 1844 4620 1896
rect 4672 1844 4678 1896
rect 4816 1893 4844 2060
rect 5994 2048 6000 2060
rect 6052 2048 6058 2100
rect 10962 2048 10968 2100
rect 11020 2088 11026 2100
rect 11020 2060 12434 2088
rect 11020 2048 11026 2060
rect 6914 1980 6920 2032
rect 6972 2020 6978 2032
rect 7469 2023 7527 2029
rect 7469 2020 7481 2023
rect 6972 1992 7481 2020
rect 6972 1980 6978 1992
rect 7469 1989 7481 1992
rect 7515 1989 7527 2023
rect 7469 1983 7527 1989
rect 6270 1912 6276 1964
rect 6328 1912 6334 1964
rect 10226 1952 10232 1964
rect 9784 1924 10232 1952
rect 4801 1887 4859 1893
rect 4801 1853 4813 1887
rect 4847 1853 4859 1887
rect 4801 1847 4859 1853
rect 5077 1887 5135 1893
rect 5077 1853 5089 1887
rect 5123 1853 5135 1887
rect 5077 1847 5135 1853
rect 4632 1816 4660 1844
rect 3436 1788 4660 1816
rect 5092 1816 5120 1847
rect 5258 1844 5264 1896
rect 5316 1884 5322 1896
rect 5353 1887 5411 1893
rect 5353 1884 5365 1887
rect 5316 1856 5365 1884
rect 5316 1844 5322 1856
rect 5353 1853 5365 1856
rect 5399 1853 5411 1887
rect 5353 1847 5411 1853
rect 6181 1887 6239 1893
rect 6181 1853 6193 1887
rect 6227 1853 6239 1887
rect 6181 1847 6239 1853
rect 5442 1816 5448 1828
rect 5092 1788 5448 1816
rect 2869 1779 2927 1785
rect 5442 1776 5448 1788
rect 5500 1776 5506 1828
rect 6196 1816 6224 1847
rect 6546 1844 6552 1896
rect 6604 1844 6610 1896
rect 7377 1887 7435 1893
rect 7377 1853 7389 1887
rect 7423 1884 7435 1887
rect 7466 1884 7472 1896
rect 7423 1856 7472 1884
rect 7423 1853 7435 1856
rect 7377 1847 7435 1853
rect 7466 1844 7472 1856
rect 7524 1844 7530 1896
rect 9030 1844 9036 1896
rect 9088 1844 9094 1896
rect 9309 1887 9367 1893
rect 9309 1853 9321 1887
rect 9355 1884 9367 1887
rect 9784 1884 9812 1924
rect 10226 1912 10232 1924
rect 10284 1912 10290 1964
rect 12406 1952 12434 2060
rect 18874 2048 18880 2100
rect 18932 2088 18938 2100
rect 22278 2088 22284 2100
rect 18932 2060 22284 2088
rect 18932 2048 18938 2060
rect 20622 1980 20628 2032
rect 20680 2020 20686 2032
rect 20680 1992 20944 2020
rect 20680 1980 20686 1992
rect 14458 1952 14464 1964
rect 12406 1924 14464 1952
rect 9355 1856 9812 1884
rect 9355 1853 9367 1856
rect 9309 1847 9367 1853
rect 10042 1844 10048 1896
rect 10100 1884 10106 1896
rect 10137 1887 10195 1893
rect 10137 1884 10149 1887
rect 10100 1856 10149 1884
rect 10100 1844 10106 1856
rect 10137 1853 10149 1856
rect 10183 1853 10195 1887
rect 10137 1847 10195 1853
rect 10870 1844 10876 1896
rect 10928 1844 10934 1896
rect 11054 1844 11060 1896
rect 11112 1844 11118 1896
rect 11517 1887 11575 1893
rect 11517 1853 11529 1887
rect 11563 1884 11575 1887
rect 11609 1887 11667 1893
rect 11609 1884 11621 1887
rect 11563 1856 11621 1884
rect 11563 1853 11575 1856
rect 11517 1847 11575 1853
rect 11609 1853 11621 1856
rect 11655 1853 11667 1887
rect 11609 1847 11667 1853
rect 11882 1844 11888 1896
rect 11940 1844 11946 1896
rect 12710 1844 12716 1896
rect 12768 1844 12774 1896
rect 12805 1887 12863 1893
rect 12805 1853 12817 1887
rect 12851 1884 12863 1887
rect 12894 1884 12900 1896
rect 12851 1856 12900 1884
rect 12851 1853 12863 1856
rect 12805 1847 12863 1853
rect 12894 1844 12900 1856
rect 12952 1844 12958 1896
rect 13280 1893 13308 1924
rect 14458 1912 14464 1924
rect 14516 1912 14522 1964
rect 15194 1912 15200 1964
rect 15252 1912 15258 1964
rect 12989 1887 13047 1893
rect 12989 1853 13001 1887
rect 13035 1884 13047 1887
rect 13081 1887 13139 1893
rect 13081 1884 13093 1887
rect 13035 1856 13093 1884
rect 13035 1853 13047 1856
rect 12989 1847 13047 1853
rect 13081 1853 13093 1856
rect 13127 1853 13139 1887
rect 13081 1847 13139 1853
rect 13265 1887 13323 1893
rect 13265 1853 13277 1887
rect 13311 1853 13323 1887
rect 13265 1847 13323 1853
rect 6638 1816 6644 1828
rect 6196 1788 6644 1816
rect 6638 1776 6644 1788
rect 6696 1776 6702 1828
rect 11790 1776 11796 1828
rect 11848 1816 11854 1828
rect 13004 1816 13032 1847
rect 13538 1844 13544 1896
rect 13596 1844 13602 1896
rect 14093 1887 14151 1893
rect 14093 1853 14105 1887
rect 14139 1884 14151 1887
rect 14182 1884 14188 1896
rect 14139 1856 14188 1884
rect 14139 1853 14151 1856
rect 14093 1847 14151 1853
rect 14182 1844 14188 1856
rect 14240 1844 14246 1896
rect 14550 1844 14556 1896
rect 14608 1844 14614 1896
rect 15470 1844 15476 1896
rect 15528 1844 15534 1896
rect 16114 1844 16120 1896
rect 16172 1884 16178 1896
rect 16301 1887 16359 1893
rect 16301 1884 16313 1887
rect 16172 1856 16313 1884
rect 16172 1844 16178 1856
rect 16301 1853 16313 1856
rect 16347 1853 16359 1887
rect 16301 1847 16359 1853
rect 16390 1844 16396 1896
rect 16448 1844 16454 1896
rect 16853 1887 16911 1893
rect 16853 1853 16865 1887
rect 16899 1884 16911 1887
rect 17310 1884 17316 1896
rect 16899 1856 17316 1884
rect 16899 1853 16911 1856
rect 16853 1847 16911 1853
rect 17310 1844 17316 1856
rect 17368 1844 17374 1896
rect 17405 1887 17463 1893
rect 17405 1853 17417 1887
rect 17451 1884 17463 1887
rect 17586 1884 17592 1896
rect 17451 1856 17592 1884
rect 17451 1853 17463 1856
rect 17405 1847 17463 1853
rect 17586 1844 17592 1856
rect 17644 1844 17650 1896
rect 17862 1844 17868 1896
rect 17920 1844 17926 1896
rect 18690 1844 18696 1896
rect 18748 1844 18754 1896
rect 19153 1887 19211 1893
rect 19153 1853 19165 1887
rect 19199 1884 19211 1887
rect 19242 1884 19248 1896
rect 19199 1856 19248 1884
rect 19199 1853 19211 1856
rect 19153 1847 19211 1853
rect 19242 1844 19248 1856
rect 19300 1844 19306 1896
rect 19429 1887 19487 1893
rect 19429 1853 19441 1887
rect 19475 1884 19487 1887
rect 19521 1887 19579 1893
rect 19521 1884 19533 1887
rect 19475 1856 19533 1884
rect 19475 1853 19487 1856
rect 19429 1847 19487 1853
rect 19521 1853 19533 1856
rect 19567 1853 19579 1887
rect 19521 1847 19579 1853
rect 19794 1844 19800 1896
rect 19852 1844 19858 1896
rect 20438 1844 20444 1896
rect 20496 1884 20502 1896
rect 20916 1893 20944 1992
rect 20625 1887 20683 1893
rect 20625 1884 20637 1887
rect 20496 1856 20637 1884
rect 20496 1844 20502 1856
rect 20625 1853 20637 1856
rect 20671 1853 20683 1887
rect 20625 1847 20683 1853
rect 20901 1887 20959 1893
rect 20901 1853 20913 1887
rect 20947 1853 20959 1887
rect 21008 1884 21036 2060
rect 22278 2048 22284 2060
rect 22336 2048 22342 2100
rect 22370 1980 22376 2032
rect 22428 2020 22434 2032
rect 22649 2023 22707 2029
rect 22649 2020 22661 2023
rect 22428 1992 22661 2020
rect 22428 1980 22434 1992
rect 22649 1989 22661 1992
rect 22695 1989 22707 2023
rect 22649 1983 22707 1989
rect 23566 1912 23572 1964
rect 23624 1952 23630 1964
rect 23937 1955 23995 1961
rect 23937 1952 23949 1955
rect 23624 1924 23949 1952
rect 23624 1912 23630 1924
rect 23937 1921 23949 1924
rect 23983 1921 23995 1955
rect 23937 1915 23995 1921
rect 24854 1912 24860 1964
rect 24912 1952 24918 1964
rect 25133 1955 25191 1961
rect 25133 1952 25145 1955
rect 24912 1924 25145 1952
rect 24912 1912 24918 1924
rect 25133 1921 25145 1924
rect 25179 1921 25191 1955
rect 25133 1915 25191 1921
rect 21085 1887 21143 1893
rect 21085 1884 21097 1887
rect 21008 1856 21097 1884
rect 20901 1847 20959 1853
rect 21085 1853 21097 1856
rect 21131 1853 21143 1887
rect 21085 1847 21143 1853
rect 21177 1887 21235 1893
rect 21177 1853 21189 1887
rect 21223 1884 21235 1887
rect 21358 1884 21364 1896
rect 21223 1856 21364 1884
rect 21223 1853 21235 1856
rect 21177 1847 21235 1853
rect 21358 1844 21364 1856
rect 21416 1844 21422 1896
rect 21453 1887 21511 1893
rect 21453 1853 21465 1887
rect 21499 1853 21511 1887
rect 21453 1847 21511 1853
rect 11848 1788 13032 1816
rect 20993 1819 21051 1825
rect 11848 1776 11854 1788
rect 20993 1785 21005 1819
rect 21039 1816 21051 1819
rect 21468 1816 21496 1847
rect 22186 1844 22192 1896
rect 22244 1884 22250 1896
rect 22281 1887 22339 1893
rect 22281 1884 22293 1887
rect 22244 1856 22293 1884
rect 22244 1844 22250 1856
rect 22281 1853 22293 1856
rect 22327 1853 22339 1887
rect 22281 1847 22339 1853
rect 22373 1887 22431 1893
rect 22373 1853 22385 1887
rect 22419 1884 22431 1887
rect 22462 1884 22468 1896
rect 22419 1856 22468 1884
rect 22419 1853 22431 1856
rect 22373 1847 22431 1853
rect 22462 1844 22468 1856
rect 22520 1844 22526 1896
rect 23109 1887 23167 1893
rect 23109 1853 23121 1887
rect 23155 1884 23167 1887
rect 23382 1884 23388 1896
rect 23155 1856 23388 1884
rect 23155 1853 23167 1856
rect 23109 1847 23167 1853
rect 23382 1844 23388 1856
rect 23440 1844 23446 1896
rect 23661 1887 23719 1893
rect 23661 1853 23673 1887
rect 23707 1884 23719 1887
rect 23750 1884 23756 1896
rect 23707 1856 23756 1884
rect 23707 1853 23719 1856
rect 23661 1847 23719 1853
rect 23750 1844 23756 1856
rect 23808 1844 23814 1896
rect 24213 1887 24271 1893
rect 24213 1853 24225 1887
rect 24259 1884 24271 1887
rect 24302 1884 24308 1896
rect 24259 1856 24308 1884
rect 24259 1853 24271 1856
rect 24213 1847 24271 1853
rect 24302 1844 24308 1856
rect 24360 1844 24366 1896
rect 24946 1844 24952 1896
rect 25004 1884 25010 1896
rect 25041 1887 25099 1893
rect 25041 1884 25053 1887
rect 25004 1856 25053 1884
rect 25004 1844 25010 1856
rect 25041 1853 25053 1856
rect 25087 1853 25099 1887
rect 25041 1847 25099 1853
rect 25222 1844 25228 1896
rect 25280 1884 25286 1896
rect 25409 1887 25467 1893
rect 25409 1884 25421 1887
rect 25280 1856 25421 1884
rect 25280 1844 25286 1856
rect 25409 1853 25421 1856
rect 25455 1853 25467 1887
rect 25409 1847 25467 1853
rect 21039 1788 21496 1816
rect 21039 1785 21051 1788
rect 20993 1779 21051 1785
rect 2958 1708 2964 1760
rect 3016 1748 3022 1760
rect 3329 1751 3387 1757
rect 3329 1748 3341 1751
rect 3016 1720 3341 1748
rect 3016 1708 3022 1720
rect 3329 1717 3341 1720
rect 3375 1717 3387 1751
rect 3329 1711 3387 1717
rect 3602 1708 3608 1760
rect 3660 1708 3666 1760
rect 4433 1751 4491 1757
rect 4433 1717 4445 1751
rect 4479 1748 4491 1751
rect 4522 1748 4528 1760
rect 4479 1720 4528 1748
rect 4479 1717 4491 1720
rect 4433 1711 4491 1717
rect 4522 1708 4528 1720
rect 4580 1708 4586 1760
rect 4709 1751 4767 1757
rect 4709 1717 4721 1751
rect 4755 1748 4767 1751
rect 4798 1748 4804 1760
rect 4755 1720 4804 1748
rect 4755 1717 4767 1720
rect 4709 1711 4767 1717
rect 4798 1708 4804 1720
rect 4856 1708 4862 1760
rect 12897 1751 12955 1757
rect 12897 1717 12909 1751
rect 12943 1748 12955 1751
rect 12986 1748 12992 1760
rect 12943 1720 12992 1748
rect 12943 1717 12955 1720
rect 12897 1711 12955 1717
rect 12986 1708 12992 1720
rect 13044 1708 13050 1760
rect 13170 1708 13176 1760
rect 13228 1708 13234 1760
rect 552 1658 27576 1680
rect 552 1606 7114 1658
rect 7166 1606 7178 1658
rect 7230 1606 7242 1658
rect 7294 1606 7306 1658
rect 7358 1606 7370 1658
rect 7422 1606 13830 1658
rect 13882 1606 13894 1658
rect 13946 1606 13958 1658
rect 14010 1606 14022 1658
rect 14074 1606 14086 1658
rect 14138 1606 20546 1658
rect 20598 1606 20610 1658
rect 20662 1606 20674 1658
rect 20726 1606 20738 1658
rect 20790 1606 20802 1658
rect 20854 1606 27262 1658
rect 27314 1606 27326 1658
rect 27378 1606 27390 1658
rect 27442 1606 27454 1658
rect 27506 1606 27518 1658
rect 27570 1606 27576 1658
rect 552 1584 27576 1606
rect 8386 1544 8392 1556
rect 7668 1516 8392 1544
rect 2314 1476 2320 1488
rect 2056 1448 2320 1476
rect 1210 1368 1216 1420
rect 1268 1368 1274 1420
rect 2056 1417 2084 1448
rect 2314 1436 2320 1448
rect 2372 1436 2378 1488
rect 3510 1476 3516 1488
rect 2746 1448 3516 1476
rect 2041 1411 2099 1417
rect 2041 1377 2053 1411
rect 2087 1377 2099 1411
rect 2041 1371 2099 1377
rect 2133 1411 2191 1417
rect 2133 1377 2145 1411
rect 2179 1408 2191 1411
rect 2746 1408 2774 1448
rect 3510 1436 3516 1448
rect 3568 1436 3574 1488
rect 2179 1380 2774 1408
rect 2179 1377 2191 1380
rect 2133 1371 2191 1377
rect 2958 1368 2964 1420
rect 3016 1368 3022 1420
rect 3602 1368 3608 1420
rect 3660 1368 3666 1420
rect 4430 1368 4436 1420
rect 4488 1368 4494 1420
rect 4798 1368 4804 1420
rect 4856 1368 4862 1420
rect 5626 1368 5632 1420
rect 5684 1368 5690 1420
rect 6914 1408 6920 1420
rect 6748 1380 6920 1408
rect 937 1343 995 1349
rect 937 1309 949 1343
rect 983 1309 995 1343
rect 937 1303 995 1309
rect 952 1204 980 1303
rect 3234 1300 3240 1352
rect 3292 1300 3298 1352
rect 3326 1300 3332 1352
rect 3384 1300 3390 1352
rect 4525 1343 4583 1349
rect 4525 1309 4537 1343
rect 4571 1309 4583 1343
rect 4525 1303 4583 1309
rect 1302 1204 1308 1216
rect 952 1176 1308 1204
rect 1302 1164 1308 1176
rect 1360 1164 1366 1216
rect 4540 1204 4568 1303
rect 5442 1300 5448 1352
rect 5500 1340 5506 1352
rect 6748 1349 6776 1380
rect 6914 1368 6920 1380
rect 6972 1368 6978 1420
rect 7006 1368 7012 1420
rect 7064 1368 7070 1420
rect 7668 1408 7696 1516
rect 8386 1504 8392 1516
rect 8444 1504 8450 1556
rect 11146 1544 11152 1556
rect 10796 1516 11152 1544
rect 7837 1411 7895 1417
rect 7837 1408 7849 1411
rect 7668 1380 7849 1408
rect 7837 1377 7849 1380
rect 7883 1377 7895 1411
rect 7837 1371 7895 1377
rect 8202 1368 8208 1420
rect 8260 1368 8266 1420
rect 8938 1368 8944 1420
rect 8996 1408 9002 1420
rect 9033 1411 9091 1417
rect 9033 1408 9045 1411
rect 8996 1380 9045 1408
rect 8996 1368 9002 1380
rect 9033 1377 9045 1380
rect 9079 1377 9091 1411
rect 9033 1371 9091 1377
rect 9950 1368 9956 1420
rect 10008 1368 10014 1420
rect 10796 1417 10824 1516
rect 11146 1504 11152 1516
rect 11204 1504 11210 1556
rect 17770 1504 17776 1556
rect 17828 1544 17834 1556
rect 17828 1516 18460 1544
rect 17828 1504 17834 1516
rect 11054 1436 11060 1488
rect 11112 1436 11118 1488
rect 17034 1436 17040 1488
rect 17092 1476 17098 1488
rect 17092 1448 17632 1476
rect 17092 1436 17098 1448
rect 10781 1411 10839 1417
rect 10781 1377 10793 1411
rect 10827 1377 10839 1411
rect 11072 1408 11100 1436
rect 10781 1371 10839 1377
rect 10980 1380 11100 1408
rect 11241 1411 11299 1417
rect 6089 1343 6147 1349
rect 6089 1340 6101 1343
rect 5500 1312 6101 1340
rect 5500 1300 5506 1312
rect 6089 1309 6101 1312
rect 6135 1309 6147 1343
rect 6089 1303 6147 1309
rect 6733 1343 6791 1349
rect 6733 1309 6745 1343
rect 6779 1309 6791 1343
rect 6733 1303 6791 1309
rect 7926 1300 7932 1352
rect 7984 1300 7990 1352
rect 10980 1349 11008 1380
rect 11241 1377 11253 1411
rect 11287 1408 11299 1411
rect 11330 1408 11336 1420
rect 11287 1380 11336 1408
rect 11287 1377 11299 1380
rect 11241 1371 11299 1377
rect 11330 1368 11336 1380
rect 11388 1368 11394 1420
rect 12066 1368 12072 1420
rect 12124 1368 12130 1420
rect 12986 1368 12992 1420
rect 13044 1368 13050 1420
rect 13265 1411 13323 1417
rect 13265 1377 13277 1411
rect 13311 1408 13323 1411
rect 13538 1408 13544 1420
rect 13311 1380 13544 1408
rect 13311 1377 13323 1380
rect 13265 1371 13323 1377
rect 13538 1368 13544 1380
rect 13596 1368 13602 1420
rect 13633 1411 13691 1417
rect 13633 1377 13645 1411
rect 13679 1408 13691 1411
rect 13722 1408 13728 1420
rect 13679 1380 13728 1408
rect 13679 1377 13691 1380
rect 13633 1371 13691 1377
rect 13722 1368 13728 1380
rect 13780 1368 13786 1420
rect 14458 1368 14464 1420
rect 14516 1368 14522 1420
rect 14550 1368 14556 1420
rect 14608 1368 14614 1420
rect 14826 1368 14832 1420
rect 14884 1368 14890 1420
rect 15562 1368 15568 1420
rect 15620 1408 15626 1420
rect 15657 1411 15715 1417
rect 15657 1408 15669 1411
rect 15620 1380 15669 1408
rect 15620 1368 15626 1380
rect 15657 1377 15669 1380
rect 15703 1377 15715 1411
rect 15657 1371 15715 1377
rect 16298 1368 16304 1420
rect 16356 1408 16362 1420
rect 16393 1411 16451 1417
rect 16393 1408 16405 1411
rect 16356 1380 16405 1408
rect 16356 1368 16362 1380
rect 16393 1377 16405 1380
rect 16439 1377 16451 1411
rect 16393 1371 16451 1377
rect 16758 1368 16764 1420
rect 16816 1408 16822 1420
rect 17221 1411 17279 1417
rect 17221 1408 17233 1411
rect 16816 1380 17233 1408
rect 16816 1368 16822 1380
rect 17221 1377 17233 1380
rect 17267 1377 17279 1411
rect 17221 1371 17279 1377
rect 17310 1368 17316 1420
rect 17368 1368 17374 1420
rect 17604 1417 17632 1448
rect 17862 1436 17868 1488
rect 17920 1436 17926 1488
rect 17589 1411 17647 1417
rect 17589 1377 17601 1411
rect 17635 1377 17647 1411
rect 17880 1408 17908 1436
rect 18432 1417 18460 1516
rect 18506 1436 18512 1488
rect 18564 1436 18570 1488
rect 19058 1436 19064 1488
rect 19116 1476 19122 1488
rect 19116 1448 20024 1476
rect 19116 1436 19122 1448
rect 18417 1411 18475 1417
rect 17880 1380 18000 1408
rect 17589 1371 17647 1377
rect 9585 1343 9643 1349
rect 9585 1309 9597 1343
rect 9631 1340 9643 1343
rect 9677 1343 9735 1349
rect 9677 1340 9689 1343
rect 9631 1312 9689 1340
rect 9631 1309 9643 1312
rect 9585 1303 9643 1309
rect 9677 1309 9689 1312
rect 9723 1309 9735 1343
rect 9677 1303 9735 1309
rect 10965 1343 11023 1349
rect 10965 1309 10977 1343
rect 11011 1309 11023 1343
rect 10965 1303 11023 1309
rect 13354 1300 13360 1352
rect 13412 1300 13418 1352
rect 15933 1343 15991 1349
rect 15933 1309 15945 1343
rect 15979 1340 15991 1343
rect 16117 1343 16175 1349
rect 16117 1340 16129 1343
rect 15979 1312 16129 1340
rect 15979 1309 15991 1312
rect 15933 1303 15991 1309
rect 16117 1309 16129 1312
rect 16163 1309 16175 1343
rect 17972 1340 18000 1380
rect 18417 1377 18429 1411
rect 18463 1377 18475 1411
rect 18524 1408 18552 1436
rect 18785 1411 18843 1417
rect 18785 1408 18797 1411
rect 18524 1380 18797 1408
rect 18417 1371 18475 1377
rect 18785 1377 18797 1380
rect 18831 1377 18843 1411
rect 18785 1371 18843 1377
rect 18874 1368 18880 1420
rect 18932 1408 18938 1420
rect 19996 1417 20024 1448
rect 22278 1436 22284 1488
rect 22336 1476 22342 1488
rect 22336 1448 22784 1476
rect 22336 1436 22342 1448
rect 19613 1411 19671 1417
rect 19613 1408 19625 1411
rect 18932 1380 19625 1408
rect 18932 1368 18938 1380
rect 19613 1377 19625 1380
rect 19659 1377 19671 1411
rect 19613 1371 19671 1377
rect 19981 1411 20039 1417
rect 19981 1377 19993 1411
rect 20027 1377 20039 1411
rect 19981 1371 20039 1377
rect 20070 1368 20076 1420
rect 20128 1408 20134 1420
rect 20809 1411 20867 1417
rect 20809 1408 20821 1411
rect 20128 1380 20821 1408
rect 20128 1368 20134 1380
rect 20809 1377 20821 1380
rect 20855 1377 20867 1411
rect 20809 1371 20867 1377
rect 21542 1368 21548 1420
rect 21600 1368 21606 1420
rect 21634 1368 21640 1420
rect 21692 1408 21698 1420
rect 22373 1411 22431 1417
rect 22373 1408 22385 1411
rect 21692 1380 22385 1408
rect 21692 1368 21698 1380
rect 22373 1377 22385 1380
rect 22419 1377 22431 1411
rect 22373 1371 22431 1377
rect 22462 1368 22468 1420
rect 22520 1368 22526 1420
rect 22756 1417 22784 1448
rect 22922 1436 22928 1488
rect 22980 1476 22986 1488
rect 22980 1448 23980 1476
rect 22980 1436 22986 1448
rect 22741 1411 22799 1417
rect 22741 1377 22753 1411
rect 22787 1377 22799 1411
rect 22741 1371 22799 1377
rect 22830 1368 22836 1420
rect 22888 1408 22894 1420
rect 23952 1417 23980 1448
rect 23569 1411 23627 1417
rect 23569 1408 23581 1411
rect 22888 1380 23581 1408
rect 22888 1368 22894 1380
rect 23569 1377 23581 1380
rect 23615 1377 23627 1411
rect 23569 1371 23627 1377
rect 23937 1411 23995 1417
rect 23937 1377 23949 1411
rect 23983 1377 23995 1411
rect 23937 1371 23995 1377
rect 24302 1368 24308 1420
rect 24360 1408 24366 1420
rect 24765 1411 24823 1417
rect 24765 1408 24777 1411
rect 24360 1380 24777 1408
rect 24360 1368 24366 1380
rect 24765 1377 24777 1380
rect 24811 1377 24823 1411
rect 24765 1371 24823 1377
rect 24854 1368 24860 1420
rect 24912 1368 24918 1420
rect 25130 1368 25136 1420
rect 25188 1368 25194 1420
rect 25498 1368 25504 1420
rect 25556 1408 25562 1420
rect 25961 1411 26019 1417
rect 25961 1408 25973 1411
rect 25556 1380 25973 1408
rect 25556 1368 25562 1380
rect 25961 1377 25973 1380
rect 26007 1377 26019 1411
rect 25961 1371 26019 1377
rect 18509 1343 18567 1349
rect 18509 1340 18521 1343
rect 17972 1312 18521 1340
rect 16117 1303 16175 1309
rect 18509 1309 18521 1312
rect 18555 1309 18567 1343
rect 18509 1303 18567 1309
rect 19242 1300 19248 1352
rect 19300 1340 19306 1352
rect 19705 1343 19763 1349
rect 19705 1340 19717 1343
rect 19300 1312 19717 1340
rect 19300 1300 19306 1312
rect 19705 1309 19717 1312
rect 19751 1309 19763 1343
rect 19705 1303 19763 1309
rect 21266 1300 21272 1352
rect 21324 1300 21330 1352
rect 23382 1300 23388 1352
rect 23440 1340 23446 1352
rect 23661 1343 23719 1349
rect 23661 1340 23673 1343
rect 23440 1312 23673 1340
rect 23440 1300 23446 1312
rect 23661 1309 23673 1312
rect 23707 1309 23719 1343
rect 23661 1303 23719 1309
rect 5997 1275 6055 1281
rect 5997 1241 6009 1275
rect 6043 1272 6055 1275
rect 6043 1244 6868 1272
rect 6043 1241 6055 1244
rect 5997 1235 6055 1241
rect 6840 1216 6868 1244
rect 5442 1204 5448 1216
rect 4540 1176 5448 1204
rect 5442 1164 5448 1176
rect 5500 1164 5506 1216
rect 6641 1207 6699 1213
rect 6641 1173 6653 1207
rect 6687 1204 6699 1207
rect 6730 1204 6736 1216
rect 6687 1176 6736 1204
rect 6687 1173 6699 1176
rect 6641 1167 6699 1173
rect 6730 1164 6736 1176
rect 6788 1164 6794 1216
rect 6822 1164 6828 1216
rect 6880 1164 6886 1216
rect 9309 1207 9367 1213
rect 9309 1173 9321 1207
rect 9355 1204 9367 1207
rect 9398 1204 9404 1216
rect 9355 1176 9404 1204
rect 9355 1173 9367 1176
rect 9309 1167 9367 1173
rect 9398 1164 9404 1176
rect 9456 1164 9462 1216
rect 12243 1207 12301 1213
rect 12243 1173 12255 1207
rect 12289 1204 12301 1207
rect 13722 1204 13728 1216
rect 12289 1176 13728 1204
rect 12289 1173 12301 1176
rect 12243 1167 12301 1173
rect 13722 1164 13728 1176
rect 13780 1164 13786 1216
rect 19978 1164 19984 1216
rect 20036 1204 20042 1216
rect 20901 1207 20959 1213
rect 20901 1204 20913 1207
rect 20036 1176 20913 1204
rect 20036 1164 20042 1176
rect 20901 1173 20913 1176
rect 20947 1173 20959 1207
rect 20901 1167 20959 1173
rect 552 1114 27416 1136
rect 552 1062 3756 1114
rect 3808 1062 3820 1114
rect 3872 1062 3884 1114
rect 3936 1062 3948 1114
rect 4000 1062 4012 1114
rect 4064 1062 10472 1114
rect 10524 1062 10536 1114
rect 10588 1062 10600 1114
rect 10652 1062 10664 1114
rect 10716 1062 10728 1114
rect 10780 1062 17188 1114
rect 17240 1062 17252 1114
rect 17304 1062 17316 1114
rect 17368 1062 17380 1114
rect 17432 1062 17444 1114
rect 17496 1062 23904 1114
rect 23956 1062 23968 1114
rect 24020 1062 24032 1114
rect 24084 1062 24096 1114
rect 24148 1062 24160 1114
rect 24212 1062 27416 1114
rect 552 1040 27416 1062
rect 934 960 940 1012
rect 992 1000 998 1012
rect 1029 1003 1087 1009
rect 1029 1000 1041 1003
rect 992 972 1041 1000
rect 992 960 998 972
rect 1029 969 1041 972
rect 1075 969 1087 1003
rect 1029 963 1087 969
rect 1302 960 1308 1012
rect 1360 1000 1366 1012
rect 1397 1003 1455 1009
rect 1397 1000 1409 1003
rect 1360 972 1409 1000
rect 1360 960 1366 972
rect 1397 969 1409 972
rect 1443 969 1455 1003
rect 1397 963 1455 969
rect 3326 960 3332 1012
rect 3384 1000 3390 1012
rect 3421 1003 3479 1009
rect 3421 1000 3433 1003
rect 3384 972 3433 1000
rect 3384 960 3390 972
rect 3421 969 3433 972
rect 3467 969 3479 1003
rect 3421 963 3479 969
rect 5442 960 5448 1012
rect 5500 960 5506 1012
rect 7926 960 7932 1012
rect 7984 960 7990 1012
rect 9030 960 9036 1012
rect 9088 960 9094 1012
rect 13354 960 13360 1012
rect 13412 1000 13418 1012
rect 13633 1003 13691 1009
rect 13633 1000 13645 1003
rect 13412 972 13645 1000
rect 13412 960 13418 972
rect 13633 969 13645 972
rect 13679 969 13691 1003
rect 13633 963 13691 969
rect 21266 960 21272 1012
rect 21324 960 21330 1012
rect 21358 960 21364 1012
rect 21416 1000 21422 1012
rect 21545 1003 21603 1009
rect 21545 1000 21557 1003
rect 21416 972 21557 1000
rect 21416 960 21422 972
rect 21545 969 21557 972
rect 21591 969 21603 1003
rect 21545 963 21603 969
rect 23566 960 23572 1012
rect 23624 1000 23630 1012
rect 23661 1003 23719 1009
rect 23661 1000 23673 1003
rect 23624 972 23673 1000
rect 23624 960 23630 972
rect 23661 969 23673 972
rect 23707 969 23719 1003
rect 23661 963 23719 969
rect 3234 892 3240 944
rect 3292 932 3298 944
rect 3697 935 3755 941
rect 3697 932 3709 935
rect 3292 904 3709 932
rect 3292 892 3298 904
rect 3697 901 3709 904
rect 3743 901 3755 935
rect 3697 895 3755 901
rect 4154 864 4160 876
rect 2746 836 4160 864
rect 1949 799 2007 805
rect 1949 765 1961 799
rect 1995 796 2007 799
rect 2130 796 2136 808
rect 1995 768 2136 796
rect 1995 765 2007 768
rect 1949 759 2007 765
rect 2130 756 2136 768
rect 2188 756 2194 808
rect 2225 799 2283 805
rect 2225 765 2237 799
rect 2271 796 2283 799
rect 2746 796 2774 836
rect 4154 824 4160 836
rect 4212 824 4218 876
rect 4246 824 4252 876
rect 4304 824 4310 876
rect 6730 824 6736 876
rect 6788 824 6794 876
rect 9398 824 9404 876
rect 9456 824 9462 876
rect 10870 824 10876 876
rect 10928 864 10934 876
rect 10965 867 11023 873
rect 10965 864 10977 867
rect 10928 836 10977 864
rect 10928 824 10934 836
rect 10965 833 10977 836
rect 11011 833 11023 867
rect 10965 827 11023 833
rect 12250 824 12256 876
rect 12308 824 12314 876
rect 18690 824 18696 876
rect 18748 824 18754 876
rect 19978 824 19984 876
rect 20036 824 20042 876
rect 23750 824 23756 876
rect 23808 864 23814 876
rect 23845 867 23903 873
rect 23845 864 23857 867
rect 23808 836 23857 864
rect 23808 824 23814 836
rect 23845 833 23857 836
rect 23891 833 23903 867
rect 23845 827 23903 833
rect 2271 768 2774 796
rect 2271 765 2283 768
rect 2225 759 2283 765
rect 2866 756 2872 808
rect 2924 796 2930 808
rect 3053 799 3111 805
rect 3053 796 3065 799
rect 2924 768 3065 796
rect 2924 756 2930 768
rect 3053 765 3065 768
rect 3099 765 3111 799
rect 3053 759 3111 765
rect 4522 756 4528 808
rect 4580 756 4586 808
rect 5074 756 5080 808
rect 5132 796 5138 808
rect 5353 799 5411 805
rect 5353 796 5365 799
rect 5132 768 5365 796
rect 5132 756 5138 768
rect 5353 765 5365 768
rect 5399 765 5411 799
rect 5353 759 5411 765
rect 5902 756 5908 808
rect 5960 796 5966 808
rect 7009 799 7067 805
rect 7009 796 7021 799
rect 5960 768 7021 796
rect 5960 756 5966 768
rect 7009 765 7021 768
rect 7055 765 7067 799
rect 7009 759 7067 765
rect 7834 756 7840 808
rect 7892 756 7898 808
rect 9674 756 9680 808
rect 9732 756 9738 808
rect 10505 799 10563 805
rect 10505 765 10517 799
rect 10551 796 10563 799
rect 10594 796 10600 808
rect 10551 768 10600 796
rect 10551 765 10563 768
rect 10505 759 10563 765
rect 10594 756 10600 768
rect 10652 756 10658 808
rect 11238 756 11244 808
rect 11296 756 11302 808
rect 11698 756 11704 808
rect 11756 796 11762 808
rect 12069 799 12127 805
rect 12069 796 12081 799
rect 11756 768 12081 796
rect 11756 756 11762 768
rect 12069 765 12081 768
rect 12115 765 12127 799
rect 12069 759 12127 765
rect 12529 799 12587 805
rect 12529 765 12541 799
rect 12575 796 12587 799
rect 13170 796 13176 808
rect 12575 768 13176 796
rect 12575 765 12587 768
rect 12529 759 12587 765
rect 13170 756 13176 768
rect 13228 756 13234 808
rect 13354 756 13360 808
rect 13412 756 13418 808
rect 14001 799 14059 805
rect 14001 765 14013 799
rect 14047 796 14059 799
rect 14182 796 14188 808
rect 14047 768 14188 796
rect 14047 765 14059 768
rect 14001 759 14059 765
rect 14182 756 14188 768
rect 14240 756 14246 808
rect 14274 756 14280 808
rect 14332 756 14338 808
rect 15010 756 15016 808
rect 15068 796 15074 808
rect 15105 799 15163 805
rect 15105 796 15117 799
rect 15068 768 15117 796
rect 15068 756 15074 768
rect 15105 765 15117 768
rect 15151 765 15163 799
rect 15105 759 15163 765
rect 16209 799 16267 805
rect 16209 765 16221 799
rect 16255 796 16267 799
rect 16390 796 16396 808
rect 16255 768 16396 796
rect 16255 765 16267 768
rect 16209 759 16267 765
rect 16390 756 16396 768
rect 16448 756 16454 808
rect 16485 799 16543 805
rect 16485 765 16497 799
rect 16531 796 16543 799
rect 16574 796 16580 808
rect 16531 768 16580 796
rect 16531 765 16543 768
rect 16485 759 16543 765
rect 16574 756 16580 768
rect 16632 756 16638 808
rect 17218 756 17224 808
rect 17276 796 17282 808
rect 17313 799 17371 805
rect 17313 796 17325 799
rect 17276 768 17325 796
rect 17276 756 17282 768
rect 17313 765 17325 768
rect 17359 765 17371 799
rect 17313 759 17371 765
rect 17405 799 17463 805
rect 17405 765 17417 799
rect 17451 796 17463 799
rect 17586 796 17592 808
rect 17451 768 17592 796
rect 17451 765 17463 768
rect 17405 759 17463 765
rect 17586 756 17592 768
rect 17644 756 17650 808
rect 17678 756 17684 808
rect 17736 756 17742 808
rect 18322 756 18328 808
rect 18380 796 18386 808
rect 18509 799 18567 805
rect 18509 796 18521 799
rect 18380 768 18521 796
rect 18380 756 18386 768
rect 18509 765 18521 768
rect 18555 765 18567 799
rect 18509 759 18567 765
rect 18966 756 18972 808
rect 19024 756 19030 808
rect 19426 756 19432 808
rect 19484 796 19490 808
rect 19797 799 19855 805
rect 19797 796 19809 799
rect 19484 768 19809 796
rect 19484 756 19490 768
rect 19797 765 19809 768
rect 19843 765 19855 799
rect 19797 759 19855 765
rect 20254 756 20260 808
rect 20312 756 20318 808
rect 21082 756 21088 808
rect 21140 756 21146 808
rect 22189 799 22247 805
rect 22189 765 22201 799
rect 22235 796 22247 799
rect 22370 796 22376 808
rect 22235 768 22376 796
rect 22235 765 22247 768
rect 22189 759 22247 765
rect 22370 756 22376 768
rect 22428 756 22434 808
rect 22465 799 22523 805
rect 22465 765 22477 799
rect 22511 796 22523 799
rect 22554 796 22560 808
rect 22511 768 22560 796
rect 22511 765 22523 768
rect 22465 759 22523 765
rect 22554 756 22560 768
rect 22612 756 22618 808
rect 23290 756 23296 808
rect 23348 756 23354 808
rect 23658 756 23664 808
rect 23716 796 23722 808
rect 24121 799 24179 805
rect 24121 796 24133 799
rect 23716 768 24133 796
rect 23716 756 23722 768
rect 24121 765 24133 768
rect 24167 765 24179 799
rect 24121 759 24179 765
rect 24486 756 24492 808
rect 24544 796 24550 808
rect 24949 799 25007 805
rect 24949 796 24961 799
rect 24544 768 24961 796
rect 24544 756 24550 768
rect 24949 765 24961 768
rect 24995 765 25007 799
rect 24949 759 25007 765
rect 25041 799 25099 805
rect 25041 765 25053 799
rect 25087 796 25099 799
rect 25222 796 25228 808
rect 25087 768 25228 796
rect 25087 765 25099 768
rect 25041 759 25099 765
rect 25222 756 25228 768
rect 25280 756 25286 808
rect 25314 756 25320 808
rect 25372 756 25378 808
rect 26050 756 26056 808
rect 26108 796 26114 808
rect 26145 799 26203 805
rect 26145 796 26157 799
rect 26108 768 26157 796
rect 26108 756 26114 768
rect 26145 765 26157 768
rect 26191 765 26203 799
rect 26145 759 26203 765
rect 552 570 27576 592
rect 552 518 7114 570
rect 7166 518 7178 570
rect 7230 518 7242 570
rect 7294 518 7306 570
rect 7358 518 7370 570
rect 7422 518 13830 570
rect 13882 518 13894 570
rect 13946 518 13958 570
rect 14010 518 14022 570
rect 14074 518 14086 570
rect 14138 518 20546 570
rect 20598 518 20610 570
rect 20662 518 20674 570
rect 20726 518 20738 570
rect 20790 518 20802 570
rect 20854 518 27262 570
rect 27314 518 27326 570
rect 27378 518 27390 570
rect 27442 518 27454 570
rect 27506 518 27518 570
rect 27570 518 27576 570
rect 552 496 27576 518
rect 20438 416 20444 468
rect 20496 456 20502 468
rect 20622 456 20628 468
rect 20496 428 20628 456
rect 20496 416 20502 428
rect 20622 416 20628 428
rect 20680 416 20686 468
<< via1 >>
rect 16672 31084 16724 31136
rect 19432 31084 19484 31136
rect 7114 30982 7166 31034
rect 7178 30982 7230 31034
rect 7242 30982 7294 31034
rect 7306 30982 7358 31034
rect 7370 30982 7422 31034
rect 13830 30982 13882 31034
rect 13894 30982 13946 31034
rect 13958 30982 14010 31034
rect 14022 30982 14074 31034
rect 14086 30982 14138 31034
rect 20546 30982 20598 31034
rect 20610 30982 20662 31034
rect 20674 30982 20726 31034
rect 20738 30982 20790 31034
rect 20802 30982 20854 31034
rect 27262 30982 27314 31034
rect 27326 30982 27378 31034
rect 27390 30982 27442 31034
rect 27454 30982 27506 31034
rect 27518 30982 27570 31034
rect 10140 30855 10192 30864
rect 5632 30744 5684 30796
rect 10140 30821 10167 30855
rect 10167 30821 10192 30855
rect 10140 30812 10192 30821
rect 6368 30608 6420 30660
rect 7564 30744 7616 30796
rect 8760 30744 8812 30796
rect 10232 30744 10284 30796
rect 6920 30719 6972 30728
rect 6920 30685 6929 30719
rect 6929 30685 6963 30719
rect 6963 30685 6972 30719
rect 6920 30676 6972 30685
rect 8024 30719 8076 30728
rect 8024 30685 8033 30719
rect 8033 30685 8067 30719
rect 8067 30685 8076 30719
rect 8024 30676 8076 30685
rect 11704 30744 11756 30796
rect 12072 30744 12124 30796
rect 8760 30608 8812 30660
rect 11244 30608 11296 30660
rect 12716 30676 12768 30728
rect 16120 30812 16172 30864
rect 14188 30744 14240 30796
rect 14648 30744 14700 30796
rect 16672 30787 16724 30796
rect 16672 30753 16681 30787
rect 16681 30753 16715 30787
rect 16715 30753 16724 30787
rect 16672 30744 16724 30753
rect 17960 30812 18012 30864
rect 19432 30880 19484 30932
rect 19156 30812 19208 30864
rect 19340 30812 19392 30864
rect 20904 30812 20956 30864
rect 22100 30812 22152 30864
rect 17684 30787 17736 30796
rect 17684 30753 17693 30787
rect 17693 30753 17727 30787
rect 17727 30753 17736 30787
rect 17684 30744 17736 30753
rect 17776 30787 17828 30796
rect 17776 30753 17785 30787
rect 17785 30753 17819 30787
rect 17819 30753 17828 30787
rect 17776 30744 17828 30753
rect 18052 30787 18104 30796
rect 18052 30753 18061 30787
rect 18061 30753 18095 30787
rect 18095 30753 18104 30787
rect 18052 30744 18104 30753
rect 18788 30744 18840 30796
rect 19064 30787 19116 30796
rect 19064 30753 19073 30787
rect 19073 30753 19107 30787
rect 19107 30753 19116 30787
rect 19064 30744 19116 30753
rect 22928 30787 22980 30796
rect 22928 30753 22937 30787
rect 22937 30753 22971 30787
rect 22971 30753 22980 30787
rect 22928 30744 22980 30753
rect 23480 30744 23532 30796
rect 26424 30744 26476 30796
rect 6276 30583 6328 30592
rect 6276 30549 6285 30583
rect 6285 30549 6319 30583
rect 6319 30549 6328 30583
rect 6276 30540 6328 30549
rect 6920 30540 6972 30592
rect 9680 30540 9732 30592
rect 10324 30540 10376 30592
rect 11060 30540 11112 30592
rect 11704 30540 11756 30592
rect 13636 30583 13688 30592
rect 13636 30549 13645 30583
rect 13645 30549 13679 30583
rect 13679 30549 13688 30583
rect 13636 30540 13688 30549
rect 14004 30583 14056 30592
rect 14004 30549 14013 30583
rect 14013 30549 14047 30583
rect 14047 30549 14056 30583
rect 14004 30540 14056 30549
rect 14740 30540 14792 30592
rect 20444 30676 20496 30728
rect 23572 30676 23624 30728
rect 16764 30540 16816 30592
rect 17592 30540 17644 30592
rect 17776 30540 17828 30592
rect 18696 30540 18748 30592
rect 19248 30583 19300 30592
rect 19248 30549 19257 30583
rect 19257 30549 19291 30583
rect 19291 30549 19300 30583
rect 19248 30540 19300 30549
rect 19432 30608 19484 30660
rect 22376 30540 22428 30592
rect 22560 30540 22612 30592
rect 3756 30438 3808 30490
rect 3820 30438 3872 30490
rect 3884 30438 3936 30490
rect 3948 30438 4000 30490
rect 4012 30438 4064 30490
rect 10472 30438 10524 30490
rect 10536 30438 10588 30490
rect 10600 30438 10652 30490
rect 10664 30438 10716 30490
rect 10728 30438 10780 30490
rect 17188 30438 17240 30490
rect 17252 30438 17304 30490
rect 17316 30438 17368 30490
rect 17380 30438 17432 30490
rect 17444 30438 17496 30490
rect 23904 30438 23956 30490
rect 23968 30438 24020 30490
rect 24032 30438 24084 30490
rect 24096 30438 24148 30490
rect 24160 30438 24212 30490
rect 8024 30379 8076 30388
rect 8024 30345 8033 30379
rect 8033 30345 8067 30379
rect 8067 30345 8076 30379
rect 8024 30336 8076 30345
rect 12072 30336 12124 30388
rect 12716 30379 12768 30388
rect 12716 30345 12725 30379
rect 12725 30345 12759 30379
rect 12759 30345 12768 30379
rect 12716 30336 12768 30345
rect 4344 30268 4396 30320
rect 16028 30311 16080 30320
rect 16028 30277 16037 30311
rect 16037 30277 16071 30311
rect 16071 30277 16080 30311
rect 16028 30268 16080 30277
rect 18052 30268 18104 30320
rect 6460 30200 6512 30252
rect 8484 30200 8536 30252
rect 11336 30243 11388 30252
rect 3240 30175 3292 30184
rect 3240 30141 3249 30175
rect 3249 30141 3283 30175
rect 3283 30141 3292 30175
rect 3240 30132 3292 30141
rect 5540 30132 5592 30184
rect 6920 30175 6972 30184
rect 6920 30141 6954 30175
rect 6954 30141 6972 30175
rect 2780 30107 2832 30116
rect 2780 30073 2798 30107
rect 2798 30073 2832 30107
rect 2780 30064 2832 30073
rect 2964 29996 3016 30048
rect 3424 29996 3476 30048
rect 4344 30064 4396 30116
rect 5816 30064 5868 30116
rect 6920 30132 6972 30141
rect 8300 30132 8352 30184
rect 8852 30175 8904 30184
rect 8852 30141 8861 30175
rect 8861 30141 8895 30175
rect 8895 30141 8904 30175
rect 8852 30132 8904 30141
rect 9128 30175 9180 30184
rect 9128 30141 9137 30175
rect 9137 30141 9171 30175
rect 9171 30141 9180 30175
rect 9128 30132 9180 30141
rect 9404 30132 9456 30184
rect 11336 30209 11345 30243
rect 11345 30209 11379 30243
rect 11379 30209 11388 30243
rect 11336 30200 11388 30209
rect 21548 30268 21600 30320
rect 20444 30243 20496 30252
rect 20444 30209 20453 30243
rect 20453 30209 20487 30243
rect 20487 30209 20496 30243
rect 20444 30200 20496 30209
rect 21824 30200 21876 30252
rect 11060 30175 11112 30184
rect 11060 30141 11069 30175
rect 11069 30141 11103 30175
rect 11103 30141 11112 30175
rect 11060 30132 11112 30141
rect 11244 30175 11296 30184
rect 11244 30141 11253 30175
rect 11253 30141 11287 30175
rect 11287 30141 11296 30175
rect 11244 30132 11296 30141
rect 13176 30132 13228 30184
rect 13728 30175 13780 30184
rect 13728 30141 13737 30175
rect 13737 30141 13771 30175
rect 13771 30141 13780 30175
rect 13728 30132 13780 30141
rect 6092 29996 6144 30048
rect 6368 30039 6420 30048
rect 6368 30005 6377 30039
rect 6377 30005 6411 30039
rect 6411 30005 6420 30039
rect 6368 29996 6420 30005
rect 8576 30039 8628 30048
rect 8576 30005 8585 30039
rect 8585 30005 8619 30039
rect 8619 30005 8628 30039
rect 8576 29996 8628 30005
rect 8668 30039 8720 30048
rect 8668 30005 8677 30039
rect 8677 30005 8711 30039
rect 8711 30005 8720 30039
rect 8668 29996 8720 30005
rect 9312 29996 9364 30048
rect 11428 30064 11480 30116
rect 10600 29996 10652 30048
rect 10876 30039 10928 30048
rect 10876 30005 10885 30039
rect 10885 30005 10919 30039
rect 10919 30005 10928 30039
rect 10876 29996 10928 30005
rect 13176 29996 13228 30048
rect 14004 30064 14056 30116
rect 15384 30132 15436 30184
rect 16120 30132 16172 30184
rect 18512 30175 18564 30184
rect 18512 30141 18521 30175
rect 18521 30141 18555 30175
rect 18555 30141 18564 30175
rect 18512 30132 18564 30141
rect 23664 30268 23716 30320
rect 13544 30039 13596 30048
rect 13544 30005 13553 30039
rect 13553 30005 13587 30039
rect 13587 30005 13596 30039
rect 13544 29996 13596 30005
rect 14556 29996 14608 30048
rect 16856 30064 16908 30116
rect 19248 30064 19300 30116
rect 19340 30064 19392 30116
rect 21548 30107 21600 30116
rect 21548 30073 21557 30107
rect 21557 30073 21591 30107
rect 21591 30073 21600 30107
rect 21548 30064 21600 30073
rect 22284 30175 22336 30184
rect 22284 30141 22293 30175
rect 22293 30141 22327 30175
rect 22327 30141 22336 30175
rect 22284 30132 22336 30141
rect 22560 30175 22612 30184
rect 22560 30141 22594 30175
rect 22594 30141 22612 30175
rect 22560 30132 22612 30141
rect 24400 30200 24452 30252
rect 24124 30132 24176 30184
rect 25504 30175 25556 30184
rect 25504 30141 25513 30175
rect 25513 30141 25547 30175
rect 25547 30141 25556 30175
rect 25504 30132 25556 30141
rect 21364 29996 21416 30048
rect 21456 29996 21508 30048
rect 22008 30039 22060 30048
rect 22008 30005 22017 30039
rect 22017 30005 22051 30039
rect 22051 30005 22060 30039
rect 22008 29996 22060 30005
rect 23204 29996 23256 30048
rect 7114 29894 7166 29946
rect 7178 29894 7230 29946
rect 7242 29894 7294 29946
rect 7306 29894 7358 29946
rect 7370 29894 7422 29946
rect 13830 29894 13882 29946
rect 13894 29894 13946 29946
rect 13958 29894 14010 29946
rect 14022 29894 14074 29946
rect 14086 29894 14138 29946
rect 20546 29894 20598 29946
rect 20610 29894 20662 29946
rect 20674 29894 20726 29946
rect 20738 29894 20790 29946
rect 20802 29894 20854 29946
rect 27262 29894 27314 29946
rect 27326 29894 27378 29946
rect 27390 29894 27442 29946
rect 27454 29894 27506 29946
rect 27518 29894 27570 29946
rect 1400 29792 1452 29844
rect 4344 29835 4396 29844
rect 4344 29801 4353 29835
rect 4353 29801 4387 29835
rect 4387 29801 4396 29835
rect 4344 29792 4396 29801
rect 9128 29792 9180 29844
rect 10140 29835 10192 29844
rect 10140 29801 10149 29835
rect 10149 29801 10183 29835
rect 10183 29801 10192 29835
rect 10140 29792 10192 29801
rect 10324 29792 10376 29844
rect 11060 29792 11112 29844
rect 12716 29792 12768 29844
rect 14556 29792 14608 29844
rect 15108 29792 15160 29844
rect 3240 29724 3292 29776
rect 3516 29724 3568 29776
rect 5540 29724 5592 29776
rect 3332 29656 3384 29708
rect 4160 29699 4212 29708
rect 4160 29665 4169 29699
rect 4169 29665 4203 29699
rect 4203 29665 4212 29699
rect 4160 29656 4212 29665
rect 8944 29724 8996 29776
rect 6000 29699 6052 29708
rect 6000 29665 6009 29699
rect 6009 29665 6043 29699
rect 6043 29665 6052 29699
rect 6000 29656 6052 29665
rect 6276 29699 6328 29708
rect 6276 29665 6285 29699
rect 6285 29665 6319 29699
rect 6319 29665 6328 29699
rect 6276 29656 6328 29665
rect 6552 29699 6604 29708
rect 6552 29665 6561 29699
rect 6561 29665 6595 29699
rect 6595 29665 6604 29699
rect 6552 29656 6604 29665
rect 7012 29699 7064 29708
rect 7012 29665 7021 29699
rect 7021 29665 7055 29699
rect 7055 29665 7064 29699
rect 7012 29656 7064 29665
rect 8668 29656 8720 29708
rect 11244 29724 11296 29776
rect 13544 29724 13596 29776
rect 5816 29588 5868 29640
rect 6828 29631 6880 29640
rect 6828 29597 6837 29631
rect 6837 29597 6871 29631
rect 6871 29597 6880 29631
rect 6828 29588 6880 29597
rect 2504 29452 2556 29504
rect 3608 29452 3660 29504
rect 10048 29588 10100 29640
rect 10600 29699 10652 29708
rect 10600 29665 10609 29699
rect 10609 29665 10643 29699
rect 10643 29665 10652 29699
rect 10600 29656 10652 29665
rect 14556 29699 14608 29708
rect 14556 29665 14565 29699
rect 14565 29665 14599 29699
rect 14599 29665 14608 29699
rect 14556 29656 14608 29665
rect 15200 29767 15252 29776
rect 15200 29733 15209 29767
rect 15209 29733 15243 29767
rect 15243 29733 15252 29767
rect 15200 29724 15252 29733
rect 15384 29835 15436 29844
rect 15384 29801 15393 29835
rect 15393 29801 15427 29835
rect 15427 29801 15436 29835
rect 15384 29792 15436 29801
rect 16120 29835 16172 29844
rect 16120 29801 16129 29835
rect 16129 29801 16163 29835
rect 16163 29801 16172 29835
rect 16120 29792 16172 29801
rect 18512 29792 18564 29844
rect 21548 29792 21600 29844
rect 12532 29588 12584 29640
rect 12624 29588 12676 29640
rect 15200 29588 15252 29640
rect 15384 29588 15436 29640
rect 16764 29724 16816 29776
rect 17592 29699 17644 29708
rect 17592 29665 17626 29699
rect 17626 29665 17644 29699
rect 17592 29656 17644 29665
rect 21364 29724 21416 29776
rect 23664 29792 23716 29844
rect 24124 29835 24176 29844
rect 24124 29801 24133 29835
rect 24133 29801 24167 29835
rect 24167 29801 24176 29835
rect 24124 29792 24176 29801
rect 18880 29656 18932 29708
rect 20444 29656 20496 29708
rect 21456 29699 21508 29708
rect 21456 29665 21465 29699
rect 21465 29665 21499 29699
rect 21499 29665 21508 29699
rect 21456 29656 21508 29665
rect 15292 29520 15344 29572
rect 16580 29520 16632 29572
rect 16856 29520 16908 29572
rect 20076 29520 20128 29572
rect 21824 29699 21876 29708
rect 21824 29665 21833 29699
rect 21833 29665 21867 29699
rect 21867 29665 21876 29699
rect 21824 29656 21876 29665
rect 22468 29767 22520 29776
rect 22468 29733 22477 29767
rect 22477 29733 22511 29767
rect 22511 29733 22520 29767
rect 22468 29724 22520 29733
rect 22744 29724 22796 29776
rect 25044 29724 25096 29776
rect 22652 29699 22704 29708
rect 22652 29665 22661 29699
rect 22661 29665 22695 29699
rect 22695 29665 22704 29699
rect 22652 29656 22704 29665
rect 23480 29656 23532 29708
rect 24308 29588 24360 29640
rect 24492 29588 24544 29640
rect 26976 29631 27028 29640
rect 26976 29597 26985 29631
rect 26985 29597 27019 29631
rect 27019 29597 27028 29631
rect 26976 29588 27028 29597
rect 22560 29520 22612 29572
rect 8392 29452 8444 29504
rect 12256 29495 12308 29504
rect 12256 29461 12265 29495
rect 12265 29461 12299 29495
rect 12299 29461 12308 29495
rect 12256 29452 12308 29461
rect 13360 29452 13412 29504
rect 15660 29452 15712 29504
rect 16948 29495 17000 29504
rect 16948 29461 16957 29495
rect 16957 29461 16991 29495
rect 16991 29461 17000 29495
rect 16948 29452 17000 29461
rect 20260 29495 20312 29504
rect 20260 29461 20269 29495
rect 20269 29461 20303 29495
rect 20303 29461 20312 29495
rect 20260 29452 20312 29461
rect 21456 29452 21508 29504
rect 22008 29495 22060 29504
rect 22008 29461 22017 29495
rect 22017 29461 22051 29495
rect 22051 29461 22060 29495
rect 22008 29452 22060 29461
rect 22192 29495 22244 29504
rect 22192 29461 22201 29495
rect 22201 29461 22235 29495
rect 22235 29461 22244 29495
rect 22192 29452 22244 29461
rect 22928 29495 22980 29504
rect 22928 29461 22937 29495
rect 22937 29461 22971 29495
rect 22971 29461 22980 29495
rect 22928 29452 22980 29461
rect 23112 29495 23164 29504
rect 23112 29461 23121 29495
rect 23121 29461 23155 29495
rect 23155 29461 23164 29495
rect 23112 29452 23164 29461
rect 23388 29520 23440 29572
rect 25412 29520 25464 29572
rect 23572 29452 23624 29504
rect 23756 29452 23808 29504
rect 3756 29350 3808 29402
rect 3820 29350 3872 29402
rect 3884 29350 3936 29402
rect 3948 29350 4000 29402
rect 4012 29350 4064 29402
rect 10472 29350 10524 29402
rect 10536 29350 10588 29402
rect 10600 29350 10652 29402
rect 10664 29350 10716 29402
rect 10728 29350 10780 29402
rect 17188 29350 17240 29402
rect 17252 29350 17304 29402
rect 17316 29350 17368 29402
rect 17380 29350 17432 29402
rect 17444 29350 17496 29402
rect 23904 29350 23956 29402
rect 23968 29350 24020 29402
rect 24032 29350 24084 29402
rect 24096 29350 24148 29402
rect 24160 29350 24212 29402
rect 7012 29248 7064 29300
rect 8576 29291 8628 29300
rect 8576 29257 8585 29291
rect 8585 29257 8619 29291
rect 8619 29257 8628 29291
rect 8576 29248 8628 29257
rect 11428 29291 11480 29300
rect 11428 29257 11437 29291
rect 11437 29257 11471 29291
rect 11471 29257 11480 29291
rect 11428 29248 11480 29257
rect 15660 29291 15712 29300
rect 15660 29257 15669 29291
rect 15669 29257 15703 29291
rect 15703 29257 15712 29291
rect 15660 29248 15712 29257
rect 16672 29248 16724 29300
rect 18880 29248 18932 29300
rect 20352 29291 20404 29300
rect 20352 29257 20361 29291
rect 20361 29257 20395 29291
rect 20395 29257 20404 29291
rect 20352 29248 20404 29257
rect 21456 29291 21508 29300
rect 21456 29257 21465 29291
rect 21465 29257 21499 29291
rect 21499 29257 21508 29291
rect 21456 29248 21508 29257
rect 3516 29155 3568 29164
rect 3516 29121 3525 29155
rect 3525 29121 3559 29155
rect 3559 29121 3568 29155
rect 3516 29112 3568 29121
rect 3608 29044 3660 29096
rect 5724 29180 5776 29232
rect 6368 29180 6420 29232
rect 8852 29180 8904 29232
rect 10048 29180 10100 29232
rect 12532 29180 12584 29232
rect 17132 29180 17184 29232
rect 5356 29019 5408 29028
rect 5356 28985 5365 29019
rect 5365 28985 5399 29019
rect 5399 28985 5408 29019
rect 5356 28976 5408 28985
rect 5632 29044 5684 29096
rect 5724 29044 5776 29096
rect 6092 29087 6144 29096
rect 6092 29053 6101 29087
rect 6101 29053 6135 29087
rect 6135 29053 6144 29087
rect 6092 29044 6144 29053
rect 6644 28976 6696 29028
rect 8300 28976 8352 29028
rect 9312 29044 9364 29096
rect 9956 29044 10008 29096
rect 10324 29112 10376 29164
rect 10232 29087 10284 29096
rect 10232 29053 10241 29087
rect 10241 29053 10275 29087
rect 10275 29053 10284 29087
rect 10232 29044 10284 29053
rect 12348 29112 12400 29164
rect 13636 29112 13688 29164
rect 14740 29112 14792 29164
rect 18512 29112 18564 29164
rect 11704 29087 11756 29096
rect 11704 29053 11713 29087
rect 11713 29053 11747 29087
rect 11747 29053 11756 29087
rect 11704 29044 11756 29053
rect 13360 29044 13412 29096
rect 15292 29087 15344 29096
rect 15292 29053 15301 29087
rect 15301 29053 15335 29087
rect 15335 29053 15344 29087
rect 15292 29044 15344 29053
rect 15476 29087 15528 29096
rect 15476 29053 15485 29087
rect 15485 29053 15519 29087
rect 15519 29053 15528 29087
rect 15476 29044 15528 29053
rect 16028 29044 16080 29096
rect 16580 29087 16632 29096
rect 16580 29053 16589 29087
rect 16589 29053 16623 29087
rect 16623 29053 16632 29087
rect 16580 29044 16632 29053
rect 16764 29087 16816 29096
rect 16764 29053 16773 29087
rect 16773 29053 16807 29087
rect 16807 29053 16816 29087
rect 16764 29044 16816 29053
rect 18972 29112 19024 29164
rect 10968 29019 11020 29028
rect 10968 28985 10977 29019
rect 10977 28985 11011 29019
rect 11011 28985 11020 29019
rect 10968 28976 11020 28985
rect 11152 29019 11204 29028
rect 11152 28985 11161 29019
rect 11161 28985 11195 29019
rect 11195 28985 11204 29019
rect 11152 28976 11204 28985
rect 12164 28976 12216 29028
rect 13084 28976 13136 29028
rect 15844 28976 15896 29028
rect 16672 29019 16724 29028
rect 16672 28985 16681 29019
rect 16681 28985 16715 29019
rect 16715 28985 16724 29019
rect 16672 28976 16724 28985
rect 19156 29044 19208 29096
rect 20260 29112 20312 29164
rect 20904 29112 20956 29164
rect 21364 29155 21416 29164
rect 21364 29121 21373 29155
rect 21373 29121 21407 29155
rect 21407 29121 21416 29155
rect 21364 29112 21416 29121
rect 21548 29180 21600 29232
rect 23112 29291 23164 29300
rect 23112 29257 23121 29291
rect 23121 29257 23155 29291
rect 23155 29257 23164 29291
rect 23112 29248 23164 29257
rect 22744 29180 22796 29232
rect 22560 29112 22612 29164
rect 20076 29087 20128 29096
rect 20076 29053 20085 29087
rect 20085 29053 20119 29087
rect 20119 29053 20128 29087
rect 20076 29044 20128 29053
rect 21272 29087 21324 29096
rect 21272 29053 21281 29087
rect 21281 29053 21315 29087
rect 21315 29053 21324 29087
rect 21272 29044 21324 29053
rect 4988 28951 5040 28960
rect 4988 28917 4997 28951
rect 4997 28917 5031 28951
rect 5031 28917 5040 28951
rect 4988 28908 5040 28917
rect 5540 28908 5592 28960
rect 5632 28908 5684 28960
rect 8576 28951 8628 28960
rect 8576 28917 8585 28951
rect 8585 28917 8619 28951
rect 8619 28917 8628 28951
rect 8576 28908 8628 28917
rect 8760 28908 8812 28960
rect 9404 28951 9456 28960
rect 9404 28917 9413 28951
rect 9413 28917 9447 28951
rect 9447 28917 9456 28951
rect 9404 28908 9456 28917
rect 10140 28951 10192 28960
rect 10140 28917 10149 28951
rect 10149 28917 10183 28951
rect 10183 28917 10192 28951
rect 10140 28908 10192 28917
rect 11336 28951 11388 28960
rect 11336 28917 11345 28951
rect 11345 28917 11379 28951
rect 11379 28917 11388 28951
rect 11336 28908 11388 28917
rect 13268 28908 13320 28960
rect 16304 28951 16356 28960
rect 16304 28917 16329 28951
rect 16329 28917 16356 28951
rect 16304 28908 16356 28917
rect 19432 28976 19484 29028
rect 20352 28976 20404 29028
rect 22468 29044 22520 29096
rect 22928 29044 22980 29096
rect 23296 29180 23348 29232
rect 23204 29044 23256 29096
rect 23572 29248 23624 29300
rect 26976 29248 27028 29300
rect 24032 29155 24084 29164
rect 24032 29121 24041 29155
rect 24041 29121 24075 29155
rect 24075 29121 24084 29155
rect 24032 29112 24084 29121
rect 24124 29044 24176 29096
rect 25504 29087 25556 29096
rect 25504 29053 25513 29087
rect 25513 29053 25547 29087
rect 25547 29053 25556 29087
rect 25504 29044 25556 29053
rect 26148 29044 26200 29096
rect 17040 28951 17092 28960
rect 17040 28917 17049 28951
rect 17049 28917 17083 28951
rect 17083 28917 17092 28951
rect 17040 28908 17092 28917
rect 22560 28951 22612 28960
rect 24308 29019 24360 29028
rect 24308 28985 24342 29019
rect 24342 28985 24360 29019
rect 24308 28976 24360 28985
rect 24400 28976 24452 29028
rect 22560 28917 22585 28951
rect 22585 28917 22612 28951
rect 22560 28908 22612 28917
rect 22928 28951 22980 28960
rect 22928 28917 22937 28951
rect 22937 28917 22971 28951
rect 22971 28917 22980 28951
rect 22928 28908 22980 28917
rect 23388 28908 23440 28960
rect 25596 28976 25648 29028
rect 7114 28806 7166 28858
rect 7178 28806 7230 28858
rect 7242 28806 7294 28858
rect 7306 28806 7358 28858
rect 7370 28806 7422 28858
rect 13830 28806 13882 28858
rect 13894 28806 13946 28858
rect 13958 28806 14010 28858
rect 14022 28806 14074 28858
rect 14086 28806 14138 28858
rect 20546 28806 20598 28858
rect 20610 28806 20662 28858
rect 20674 28806 20726 28858
rect 20738 28806 20790 28858
rect 20802 28806 20854 28858
rect 27262 28806 27314 28858
rect 27326 28806 27378 28858
rect 27390 28806 27442 28858
rect 27454 28806 27506 28858
rect 27518 28806 27570 28858
rect 3056 28704 3108 28756
rect 3332 28704 3384 28756
rect 3516 28636 3568 28688
rect 4160 28704 4212 28756
rect 4988 28704 5040 28756
rect 5816 28747 5868 28756
rect 5816 28713 5825 28747
rect 5825 28713 5859 28747
rect 5859 28713 5868 28747
rect 5816 28704 5868 28713
rect 6828 28704 6880 28756
rect 3608 28611 3660 28620
rect 8116 28679 8168 28688
rect 8116 28645 8143 28679
rect 8143 28645 8168 28679
rect 8116 28636 8168 28645
rect 8576 28636 8628 28688
rect 3608 28577 3626 28611
rect 3626 28577 3660 28611
rect 3608 28568 3660 28577
rect 5356 28568 5408 28620
rect 6736 28611 6788 28620
rect 6736 28577 6770 28611
rect 6770 28577 6788 28611
rect 6736 28568 6788 28577
rect 7840 28568 7892 28620
rect 10324 28704 10376 28756
rect 9404 28636 9456 28688
rect 2872 28364 2924 28416
rect 5632 28364 5684 28416
rect 6460 28543 6512 28552
rect 6460 28509 6469 28543
rect 6469 28509 6503 28543
rect 6503 28509 6512 28543
rect 6460 28500 6512 28509
rect 8024 28500 8076 28552
rect 9772 28568 9824 28620
rect 11520 28636 11572 28688
rect 13728 28704 13780 28756
rect 15200 28747 15252 28756
rect 15200 28713 15225 28747
rect 15225 28713 15252 28747
rect 15200 28704 15252 28713
rect 7472 28432 7524 28484
rect 8300 28432 8352 28484
rect 8484 28432 8536 28484
rect 10232 28500 10284 28552
rect 12992 28568 13044 28620
rect 14648 28611 14700 28620
rect 14648 28577 14657 28611
rect 14657 28577 14691 28611
rect 14691 28577 14700 28611
rect 14648 28568 14700 28577
rect 15844 28636 15896 28688
rect 16304 28704 16356 28756
rect 23756 28747 23808 28756
rect 23756 28713 23765 28747
rect 23765 28713 23799 28747
rect 23799 28713 23808 28747
rect 23756 28704 23808 28713
rect 24308 28704 24360 28756
rect 25596 28747 25648 28756
rect 25596 28713 25605 28747
rect 25605 28713 25639 28747
rect 25639 28713 25648 28747
rect 25596 28704 25648 28713
rect 16580 28636 16632 28688
rect 15476 28568 15528 28620
rect 10324 28475 10376 28484
rect 10324 28441 10333 28475
rect 10333 28441 10367 28475
rect 10367 28441 10376 28475
rect 13912 28500 13964 28552
rect 15200 28500 15252 28552
rect 15384 28500 15436 28552
rect 15752 28568 15804 28620
rect 10324 28432 10376 28441
rect 10968 28432 11020 28484
rect 11244 28475 11296 28484
rect 11244 28441 11253 28475
rect 11253 28441 11287 28475
rect 11287 28441 11296 28475
rect 11244 28432 11296 28441
rect 6644 28364 6696 28416
rect 7840 28407 7892 28416
rect 7840 28373 7849 28407
rect 7849 28373 7883 28407
rect 7883 28373 7892 28407
rect 7840 28364 7892 28373
rect 10232 28364 10284 28416
rect 11060 28407 11112 28416
rect 11060 28373 11069 28407
rect 11069 28373 11103 28407
rect 11103 28373 11112 28407
rect 11060 28364 11112 28373
rect 11336 28364 11388 28416
rect 11796 28407 11848 28416
rect 11796 28373 11805 28407
rect 11805 28373 11839 28407
rect 11839 28373 11848 28407
rect 11796 28364 11848 28373
rect 13268 28407 13320 28416
rect 13268 28373 13277 28407
rect 13277 28373 13311 28407
rect 13311 28373 13320 28407
rect 13268 28364 13320 28373
rect 14280 28364 14332 28416
rect 15108 28364 15160 28416
rect 16856 28568 16908 28620
rect 17040 28611 17092 28620
rect 17040 28577 17074 28611
rect 17074 28577 17092 28611
rect 17040 28568 17092 28577
rect 17592 28568 17644 28620
rect 18420 28611 18472 28620
rect 18420 28577 18429 28611
rect 18429 28577 18463 28611
rect 18463 28577 18472 28611
rect 18420 28568 18472 28577
rect 24860 28636 24912 28688
rect 18788 28568 18840 28620
rect 19340 28568 19392 28620
rect 22284 28568 22336 28620
rect 19708 28500 19760 28552
rect 21640 28500 21692 28552
rect 22928 28568 22980 28620
rect 23388 28611 23440 28620
rect 23388 28577 23397 28611
rect 23397 28577 23431 28611
rect 23431 28577 23440 28611
rect 23388 28568 23440 28577
rect 23664 28568 23716 28620
rect 24308 28568 24360 28620
rect 25412 28611 25464 28620
rect 25412 28577 25421 28611
rect 25421 28577 25455 28611
rect 25455 28577 25464 28611
rect 25412 28568 25464 28577
rect 25044 28500 25096 28552
rect 16764 28364 16816 28416
rect 17868 28364 17920 28416
rect 18972 28364 19024 28416
rect 22376 28432 22428 28484
rect 22284 28407 22336 28416
rect 22284 28373 22293 28407
rect 22293 28373 22327 28407
rect 22327 28373 22336 28407
rect 22284 28364 22336 28373
rect 3756 28262 3808 28314
rect 3820 28262 3872 28314
rect 3884 28262 3936 28314
rect 3948 28262 4000 28314
rect 4012 28262 4064 28314
rect 10472 28262 10524 28314
rect 10536 28262 10588 28314
rect 10600 28262 10652 28314
rect 10664 28262 10716 28314
rect 10728 28262 10780 28314
rect 17188 28262 17240 28314
rect 17252 28262 17304 28314
rect 17316 28262 17368 28314
rect 17380 28262 17432 28314
rect 17444 28262 17496 28314
rect 23904 28262 23956 28314
rect 23968 28262 24020 28314
rect 24032 28262 24084 28314
rect 24096 28262 24148 28314
rect 24160 28262 24212 28314
rect 3608 28160 3660 28212
rect 6092 28203 6144 28212
rect 6092 28169 6101 28203
rect 6101 28169 6135 28203
rect 6135 28169 6144 28203
rect 6092 28160 6144 28169
rect 6736 28160 6788 28212
rect 8116 28203 8168 28212
rect 8116 28169 8125 28203
rect 8125 28169 8159 28203
rect 8159 28169 8168 28203
rect 8116 28160 8168 28169
rect 9956 28203 10008 28212
rect 9956 28169 9965 28203
rect 9965 28169 9999 28203
rect 9999 28169 10008 28203
rect 9956 28160 10008 28169
rect 10140 28203 10192 28212
rect 10140 28169 10149 28203
rect 10149 28169 10183 28203
rect 10183 28169 10192 28203
rect 10140 28160 10192 28169
rect 12992 28203 13044 28212
rect 12992 28169 13001 28203
rect 13001 28169 13035 28203
rect 13035 28169 13044 28203
rect 12992 28160 13044 28169
rect 13360 28160 13412 28212
rect 13912 28203 13964 28212
rect 13912 28169 13921 28203
rect 13921 28169 13955 28203
rect 13955 28169 13964 28203
rect 13912 28160 13964 28169
rect 10968 28092 11020 28144
rect 11152 28135 11204 28144
rect 11152 28101 11161 28135
rect 11161 28101 11195 28135
rect 11195 28101 11204 28135
rect 11152 28092 11204 28101
rect 10324 28024 10376 28076
rect 3240 27999 3292 28008
rect 3240 27965 3249 27999
rect 3249 27965 3283 27999
rect 3283 27965 3292 27999
rect 3240 27956 3292 27965
rect 4160 27956 4212 28008
rect 5356 27956 5408 28008
rect 5724 27956 5776 28008
rect 6828 27956 6880 28008
rect 7472 27956 7524 28008
rect 2688 27820 2740 27872
rect 3148 27888 3200 27940
rect 6184 27888 6236 27940
rect 6644 27888 6696 27940
rect 7840 27956 7892 28008
rect 8024 27888 8076 27940
rect 8392 27956 8444 28008
rect 10048 27956 10100 28008
rect 10876 27999 10928 28008
rect 10876 27965 10885 27999
rect 10885 27965 10919 27999
rect 10919 27965 10928 27999
rect 10876 27956 10928 27965
rect 11336 28067 11388 28076
rect 11336 28033 11345 28067
rect 11345 28033 11379 28067
rect 11379 28033 11388 28067
rect 11336 28024 11388 28033
rect 8484 27888 8536 27940
rect 8944 27931 8996 27940
rect 8944 27897 8953 27931
rect 8953 27897 8987 27931
rect 8987 27897 8996 27931
rect 8944 27888 8996 27897
rect 10324 27888 10376 27940
rect 11244 27956 11296 28008
rect 13084 27956 13136 28008
rect 11612 27931 11664 27940
rect 11612 27897 11646 27931
rect 11646 27897 11664 27931
rect 11612 27888 11664 27897
rect 2872 27820 2924 27872
rect 3332 27820 3384 27872
rect 3884 27863 3936 27872
rect 3884 27829 3893 27863
rect 3893 27829 3927 27863
rect 3927 27829 3936 27863
rect 3884 27820 3936 27829
rect 5908 27820 5960 27872
rect 6736 27863 6788 27872
rect 6736 27829 6745 27863
rect 6745 27829 6779 27863
rect 6779 27829 6788 27863
rect 6736 27820 6788 27829
rect 8576 27820 8628 27872
rect 11520 27820 11572 27872
rect 12716 27863 12768 27872
rect 12716 27829 12725 27863
rect 12725 27829 12759 27863
rect 12759 27829 12768 27863
rect 12716 27820 12768 27829
rect 13636 27888 13688 27940
rect 14648 28160 14700 28212
rect 18420 28203 18472 28212
rect 18420 28169 18429 28203
rect 18429 28169 18463 28203
rect 18463 28169 18472 28203
rect 18420 28160 18472 28169
rect 18788 28160 18840 28212
rect 20076 28160 20128 28212
rect 21272 28160 21324 28212
rect 21640 28203 21692 28212
rect 21640 28169 21649 28203
rect 21649 28169 21683 28203
rect 21683 28169 21692 28203
rect 21640 28160 21692 28169
rect 22100 28160 22152 28212
rect 22652 28160 22704 28212
rect 24216 28160 24268 28212
rect 24308 28203 24360 28212
rect 24308 28169 24317 28203
rect 24317 28169 24351 28203
rect 24351 28169 24360 28203
rect 24308 28160 24360 28169
rect 20904 28092 20956 28144
rect 15660 27999 15712 28008
rect 15660 27965 15669 27999
rect 15669 27965 15703 27999
rect 15703 27965 15712 27999
rect 15660 27956 15712 27965
rect 16856 27956 16908 28008
rect 17040 27956 17092 28008
rect 18420 27956 18472 28008
rect 18880 27999 18932 28008
rect 18880 27965 18889 27999
rect 18889 27965 18923 27999
rect 18923 27965 18932 27999
rect 18880 27956 18932 27965
rect 18972 27999 19024 28008
rect 18972 27965 18981 27999
rect 18981 27965 19015 27999
rect 19015 27965 19024 27999
rect 18972 27956 19024 27965
rect 14464 27888 14516 27940
rect 18328 27888 18380 27940
rect 19156 27956 19208 28008
rect 19708 27956 19760 28008
rect 20352 27956 20404 28008
rect 20904 27931 20956 27940
rect 20904 27897 20913 27931
rect 20913 27897 20947 27931
rect 20947 27897 20956 27931
rect 20904 27888 20956 27897
rect 21272 27931 21324 27940
rect 21272 27897 21281 27931
rect 21281 27897 21315 27931
rect 21315 27897 21324 27931
rect 21272 27888 21324 27897
rect 21456 27820 21508 27872
rect 22192 28092 22244 28144
rect 23572 28092 23624 28144
rect 22928 28024 22980 28076
rect 24584 28024 24636 28076
rect 22744 27956 22796 28008
rect 23020 27999 23072 28008
rect 23020 27965 23029 27999
rect 23029 27965 23063 27999
rect 23063 27965 23072 27999
rect 23020 27956 23072 27965
rect 23572 27956 23624 28008
rect 22652 27888 22704 27940
rect 23388 27888 23440 27940
rect 22192 27820 22244 27872
rect 23756 27888 23808 27940
rect 24216 27931 24268 27940
rect 24216 27897 24225 27931
rect 24225 27897 24259 27931
rect 24259 27897 24268 27931
rect 24216 27888 24268 27897
rect 25136 27999 25188 28008
rect 25136 27965 25145 27999
rect 25145 27965 25179 27999
rect 25179 27965 25188 27999
rect 25136 27956 25188 27965
rect 25044 27888 25096 27940
rect 23664 27820 23716 27872
rect 23848 27863 23900 27872
rect 23848 27829 23857 27863
rect 23857 27829 23891 27863
rect 23891 27829 23900 27863
rect 23848 27820 23900 27829
rect 25320 27863 25372 27872
rect 25320 27829 25329 27863
rect 25329 27829 25363 27863
rect 25363 27829 25372 27863
rect 25320 27820 25372 27829
rect 7114 27718 7166 27770
rect 7178 27718 7230 27770
rect 7242 27718 7294 27770
rect 7306 27718 7358 27770
rect 7370 27718 7422 27770
rect 13830 27718 13882 27770
rect 13894 27718 13946 27770
rect 13958 27718 14010 27770
rect 14022 27718 14074 27770
rect 14086 27718 14138 27770
rect 20546 27718 20598 27770
rect 20610 27718 20662 27770
rect 20674 27718 20726 27770
rect 20738 27718 20790 27770
rect 20802 27718 20854 27770
rect 27262 27718 27314 27770
rect 27326 27718 27378 27770
rect 27390 27718 27442 27770
rect 27454 27718 27506 27770
rect 27518 27718 27570 27770
rect 3240 27616 3292 27668
rect 6092 27616 6144 27668
rect 6920 27616 6972 27668
rect 8024 27616 8076 27668
rect 1860 27523 1912 27532
rect 1860 27489 1869 27523
rect 1869 27489 1903 27523
rect 1903 27489 1912 27523
rect 3884 27548 3936 27600
rect 5724 27548 5776 27600
rect 1860 27480 1912 27489
rect 3240 27480 3292 27532
rect 3608 27480 3660 27532
rect 5356 27523 5408 27532
rect 5356 27489 5365 27523
rect 5365 27489 5399 27523
rect 5399 27489 5408 27523
rect 5356 27480 5408 27489
rect 6828 27548 6880 27600
rect 11612 27659 11664 27668
rect 11612 27625 11621 27659
rect 11621 27625 11655 27659
rect 11655 27625 11664 27659
rect 11612 27616 11664 27625
rect 14464 27659 14516 27668
rect 14464 27625 14473 27659
rect 14473 27625 14507 27659
rect 14507 27625 14516 27659
rect 14464 27616 14516 27625
rect 15660 27616 15712 27668
rect 11152 27548 11204 27600
rect 5908 27523 5960 27532
rect 5908 27489 5917 27523
rect 5917 27489 5951 27523
rect 5951 27489 5960 27523
rect 5908 27480 5960 27489
rect 6184 27480 6236 27532
rect 7012 27480 7064 27532
rect 10876 27480 10928 27532
rect 11796 27523 11848 27532
rect 11796 27489 11805 27523
rect 11805 27489 11839 27523
rect 11839 27489 11848 27523
rect 11796 27480 11848 27489
rect 12716 27548 12768 27600
rect 16764 27548 16816 27600
rect 17592 27548 17644 27600
rect 13360 27480 13412 27532
rect 13636 27480 13688 27532
rect 14280 27523 14332 27532
rect 14280 27489 14289 27523
rect 14289 27489 14323 27523
rect 14323 27489 14332 27523
rect 14280 27480 14332 27489
rect 15108 27480 15160 27532
rect 15476 27480 15528 27532
rect 15844 27480 15896 27532
rect 16672 27480 16724 27532
rect 21364 27616 21416 27668
rect 3056 27412 3108 27464
rect 3332 27455 3384 27464
rect 3332 27421 3341 27455
rect 3341 27421 3375 27455
rect 3375 27421 3384 27455
rect 3332 27412 3384 27421
rect 5632 27412 5684 27464
rect 8392 27412 8444 27464
rect 8484 27412 8536 27464
rect 9772 27412 9824 27464
rect 17776 27523 17828 27532
rect 17776 27489 17785 27523
rect 17785 27489 17819 27523
rect 17819 27489 17828 27523
rect 17776 27480 17828 27489
rect 17960 27480 18012 27532
rect 18696 27480 18748 27532
rect 19340 27523 19392 27532
rect 19340 27489 19349 27523
rect 19349 27489 19383 27523
rect 19383 27489 19392 27523
rect 19340 27480 19392 27489
rect 19432 27480 19484 27532
rect 17040 27455 17092 27464
rect 17040 27421 17049 27455
rect 17049 27421 17083 27455
rect 17083 27421 17092 27455
rect 17040 27412 17092 27421
rect 23572 27616 23624 27668
rect 24216 27616 24268 27668
rect 22100 27548 22152 27600
rect 21548 27412 21600 27464
rect 22192 27480 22244 27532
rect 22652 27523 22704 27532
rect 22652 27489 22661 27523
rect 22661 27489 22695 27523
rect 22695 27489 22704 27523
rect 22652 27480 22704 27489
rect 22744 27523 22796 27532
rect 22744 27489 22753 27523
rect 22753 27489 22787 27523
rect 22787 27489 22796 27523
rect 22744 27480 22796 27489
rect 22836 27523 22888 27532
rect 22836 27489 22845 27523
rect 22845 27489 22879 27523
rect 22879 27489 22888 27523
rect 22836 27480 22888 27489
rect 23020 27523 23072 27532
rect 23020 27489 23029 27523
rect 23029 27489 23063 27523
rect 23063 27489 23072 27523
rect 23020 27480 23072 27489
rect 23664 27548 23716 27600
rect 24124 27548 24176 27600
rect 23480 27480 23532 27532
rect 25044 27548 25096 27600
rect 25320 27548 25372 27600
rect 26148 27480 26200 27532
rect 2044 27387 2096 27396
rect 2044 27353 2053 27387
rect 2053 27353 2087 27387
rect 2087 27353 2096 27387
rect 2044 27344 2096 27353
rect 2688 27319 2740 27328
rect 2688 27285 2697 27319
rect 2697 27285 2731 27319
rect 2731 27285 2740 27319
rect 2688 27276 2740 27285
rect 3148 27276 3200 27328
rect 4896 27319 4948 27328
rect 4896 27285 4905 27319
rect 4905 27285 4939 27319
rect 4939 27285 4948 27319
rect 4896 27276 4948 27285
rect 5172 27276 5224 27328
rect 5816 27319 5868 27328
rect 5816 27285 5825 27319
rect 5825 27285 5859 27319
rect 5859 27285 5868 27319
rect 5816 27276 5868 27285
rect 6184 27319 6236 27328
rect 6184 27285 6193 27319
rect 6193 27285 6227 27319
rect 6227 27285 6236 27319
rect 6184 27276 6236 27285
rect 9036 27319 9088 27328
rect 9036 27285 9045 27319
rect 9045 27285 9079 27319
rect 9079 27285 9088 27319
rect 9036 27276 9088 27285
rect 9128 27319 9180 27328
rect 9128 27285 9137 27319
rect 9137 27285 9171 27319
rect 9171 27285 9180 27319
rect 9128 27276 9180 27285
rect 9312 27387 9364 27396
rect 9312 27353 9321 27387
rect 9321 27353 9355 27387
rect 9355 27353 9364 27387
rect 9312 27344 9364 27353
rect 16856 27344 16908 27396
rect 17132 27344 17184 27396
rect 21180 27344 21232 27396
rect 9864 27276 9916 27328
rect 10876 27276 10928 27328
rect 11980 27319 12032 27328
rect 11980 27285 11989 27319
rect 11989 27285 12023 27319
rect 12023 27285 12032 27319
rect 11980 27276 12032 27285
rect 12992 27276 13044 27328
rect 13820 27276 13872 27328
rect 14924 27276 14976 27328
rect 15660 27276 15712 27328
rect 19248 27319 19300 27328
rect 19248 27285 19257 27319
rect 19257 27285 19291 27319
rect 19291 27285 19300 27319
rect 19248 27276 19300 27285
rect 20720 27319 20772 27328
rect 20720 27285 20729 27319
rect 20729 27285 20763 27319
rect 20763 27285 20772 27319
rect 20720 27276 20772 27285
rect 21548 27276 21600 27328
rect 23848 27344 23900 27396
rect 25136 27344 25188 27396
rect 22284 27319 22336 27328
rect 22284 27285 22293 27319
rect 22293 27285 22327 27319
rect 22327 27285 22336 27319
rect 22284 27276 22336 27285
rect 24584 27319 24636 27328
rect 24584 27285 24593 27319
rect 24593 27285 24627 27319
rect 24627 27285 24636 27319
rect 24584 27276 24636 27285
rect 3756 27174 3808 27226
rect 3820 27174 3872 27226
rect 3884 27174 3936 27226
rect 3948 27174 4000 27226
rect 4012 27174 4064 27226
rect 10472 27174 10524 27226
rect 10536 27174 10588 27226
rect 10600 27174 10652 27226
rect 10664 27174 10716 27226
rect 10728 27174 10780 27226
rect 17188 27174 17240 27226
rect 17252 27174 17304 27226
rect 17316 27174 17368 27226
rect 17380 27174 17432 27226
rect 17444 27174 17496 27226
rect 23904 27174 23956 27226
rect 23968 27174 24020 27226
rect 24032 27174 24084 27226
rect 24096 27174 24148 27226
rect 24160 27174 24212 27226
rect 2780 27072 2832 27124
rect 4160 27115 4212 27124
rect 4160 27081 4169 27115
rect 4169 27081 4203 27115
rect 4203 27081 4212 27115
rect 4160 27072 4212 27081
rect 5632 27115 5684 27124
rect 5632 27081 5641 27115
rect 5641 27081 5675 27115
rect 5675 27081 5684 27115
rect 5632 27072 5684 27081
rect 5724 27072 5776 27124
rect 3056 26936 3108 26988
rect 3240 26936 3292 26988
rect 5172 27004 5224 27056
rect 5356 26936 5408 26988
rect 848 26911 900 26920
rect 848 26877 857 26911
rect 857 26877 891 26911
rect 891 26877 900 26911
rect 848 26868 900 26877
rect 2412 26868 2464 26920
rect 1124 26843 1176 26852
rect 1124 26809 1158 26843
rect 1158 26809 1176 26843
rect 1124 26800 1176 26809
rect 1492 26800 1544 26852
rect 1860 26800 1912 26852
rect 2228 26775 2280 26784
rect 2228 26741 2237 26775
rect 2237 26741 2271 26775
rect 2271 26741 2280 26775
rect 2228 26732 2280 26741
rect 2320 26775 2372 26784
rect 2320 26741 2329 26775
rect 2329 26741 2363 26775
rect 2363 26741 2372 26775
rect 2320 26732 2372 26741
rect 4988 26911 5040 26920
rect 4988 26877 4997 26911
rect 4997 26877 5031 26911
rect 5031 26877 5040 26911
rect 4988 26868 5040 26877
rect 9312 27072 9364 27124
rect 10048 27072 10100 27124
rect 16304 27072 16356 27124
rect 17960 27072 18012 27124
rect 19432 27072 19484 27124
rect 21456 27115 21508 27124
rect 21456 27081 21465 27115
rect 21465 27081 21499 27115
rect 21499 27081 21508 27115
rect 21456 27072 21508 27081
rect 22100 27072 22152 27124
rect 22744 27072 22796 27124
rect 9128 27004 9180 27056
rect 6092 26911 6144 26920
rect 6092 26877 6101 26911
rect 6101 26877 6135 26911
rect 6135 26877 6144 26911
rect 6092 26868 6144 26877
rect 6368 26936 6420 26988
rect 6920 26979 6972 26988
rect 6920 26945 6929 26979
rect 6929 26945 6963 26979
rect 6963 26945 6972 26979
rect 6920 26936 6972 26945
rect 5724 26800 5776 26852
rect 8116 26911 8168 26920
rect 8116 26877 8125 26911
rect 8125 26877 8159 26911
rect 8159 26877 8168 26911
rect 8116 26868 8168 26877
rect 8484 26911 8536 26920
rect 8484 26877 8493 26911
rect 8493 26877 8527 26911
rect 8527 26877 8536 26911
rect 8484 26868 8536 26877
rect 9128 26911 9180 26920
rect 9128 26877 9138 26911
rect 9138 26877 9172 26911
rect 9172 26877 9180 26911
rect 9128 26868 9180 26877
rect 6920 26800 6972 26852
rect 5540 26732 5592 26784
rect 5908 26732 5960 26784
rect 6092 26732 6144 26784
rect 6276 26732 6328 26784
rect 6828 26732 6880 26784
rect 7472 26775 7524 26784
rect 7472 26741 7481 26775
rect 7481 26741 7515 26775
rect 7515 26741 7524 26775
rect 7472 26732 7524 26741
rect 9404 26843 9456 26852
rect 9404 26809 9413 26843
rect 9413 26809 9447 26843
rect 9447 26809 9456 26843
rect 9404 26800 9456 26809
rect 9772 26911 9824 26920
rect 9772 26877 9781 26911
rect 9781 26877 9815 26911
rect 9815 26877 9824 26911
rect 9772 26868 9824 26877
rect 15568 27004 15620 27056
rect 10508 26911 10560 26920
rect 10508 26877 10517 26911
rect 10517 26877 10551 26911
rect 10551 26877 10560 26911
rect 10508 26868 10560 26877
rect 10784 26868 10836 26920
rect 11060 26868 11112 26920
rect 11152 26868 11204 26920
rect 11980 26911 12032 26920
rect 10140 26800 10192 26852
rect 11980 26877 11989 26911
rect 11989 26877 12023 26911
rect 12023 26877 12032 26911
rect 11980 26868 12032 26877
rect 12808 26936 12860 26988
rect 12900 26911 12952 26920
rect 12900 26877 12909 26911
rect 12909 26877 12943 26911
rect 12943 26877 12952 26911
rect 12900 26868 12952 26877
rect 12992 26911 13044 26920
rect 12992 26877 13001 26911
rect 13001 26877 13035 26911
rect 13035 26877 13044 26911
rect 12992 26868 13044 26877
rect 10232 26775 10284 26784
rect 10232 26741 10241 26775
rect 10241 26741 10275 26775
rect 10275 26741 10284 26775
rect 10232 26732 10284 26741
rect 13360 26800 13412 26852
rect 13820 26911 13872 26920
rect 13820 26877 13829 26911
rect 13829 26877 13863 26911
rect 13863 26877 13872 26911
rect 13820 26868 13872 26877
rect 14280 26911 14332 26920
rect 14280 26877 14289 26911
rect 14289 26877 14323 26911
rect 14323 26877 14332 26911
rect 14280 26868 14332 26877
rect 14832 26911 14884 26920
rect 14832 26877 14841 26911
rect 14841 26877 14875 26911
rect 14875 26877 14884 26911
rect 14832 26868 14884 26877
rect 14924 26911 14976 26920
rect 14924 26877 14933 26911
rect 14933 26877 14967 26911
rect 14967 26877 14976 26911
rect 14924 26868 14976 26877
rect 16948 26936 17000 26988
rect 15568 26911 15620 26920
rect 15568 26877 15577 26911
rect 15577 26877 15611 26911
rect 15611 26877 15620 26911
rect 15568 26868 15620 26877
rect 15660 26911 15712 26920
rect 15660 26877 15669 26911
rect 15669 26877 15703 26911
rect 15703 26877 15712 26911
rect 15660 26868 15712 26877
rect 15844 26911 15896 26920
rect 15844 26877 15853 26911
rect 15853 26877 15887 26911
rect 15887 26877 15896 26911
rect 15844 26868 15896 26877
rect 17132 26868 17184 26920
rect 11152 26732 11204 26784
rect 11428 26732 11480 26784
rect 11612 26732 11664 26784
rect 12716 26775 12768 26784
rect 12716 26741 12725 26775
rect 12725 26741 12759 26775
rect 12759 26741 12768 26775
rect 12716 26732 12768 26741
rect 12992 26732 13044 26784
rect 15660 26732 15712 26784
rect 16764 26732 16816 26784
rect 18328 27004 18380 27056
rect 17776 26868 17828 26920
rect 18144 26911 18196 26920
rect 18144 26877 18153 26911
rect 18153 26877 18187 26911
rect 18187 26877 18196 26911
rect 18144 26868 18196 26877
rect 18420 26868 18472 26920
rect 19248 26868 19300 26920
rect 21272 26979 21324 26988
rect 21272 26945 21281 26979
rect 21281 26945 21315 26979
rect 21315 26945 21324 26979
rect 21272 26936 21324 26945
rect 17500 26843 17552 26852
rect 17500 26809 17509 26843
rect 17509 26809 17543 26843
rect 17543 26809 17552 26843
rect 17500 26800 17552 26809
rect 18236 26843 18288 26852
rect 18236 26809 18245 26843
rect 18245 26809 18279 26843
rect 18279 26809 18288 26843
rect 18236 26800 18288 26809
rect 20904 26911 20956 26920
rect 20904 26877 20913 26911
rect 20913 26877 20947 26911
rect 20947 26877 20956 26911
rect 20904 26868 20956 26877
rect 21088 26911 21140 26920
rect 21088 26877 21097 26911
rect 21097 26877 21131 26911
rect 21131 26877 21140 26911
rect 21088 26868 21140 26877
rect 21180 26911 21232 26920
rect 21180 26877 21189 26911
rect 21189 26877 21223 26911
rect 21223 26877 21232 26911
rect 21180 26868 21232 26877
rect 22468 27004 22520 27056
rect 21916 26936 21968 26988
rect 22652 26936 22704 26988
rect 21824 26800 21876 26852
rect 22100 26868 22152 26920
rect 22836 26868 22888 26920
rect 23756 26868 23808 26920
rect 24032 26843 24084 26852
rect 24032 26809 24041 26843
rect 24041 26809 24075 26843
rect 24075 26809 24084 26843
rect 25044 26868 25096 26920
rect 25320 26868 25372 26920
rect 26148 26868 26200 26920
rect 24032 26800 24084 26809
rect 20720 26732 20772 26784
rect 21916 26732 21968 26784
rect 22100 26732 22152 26784
rect 23020 26732 23072 26784
rect 25136 26775 25188 26784
rect 25136 26741 25145 26775
rect 25145 26741 25179 26775
rect 25179 26741 25188 26775
rect 25136 26732 25188 26741
rect 25596 26732 25648 26784
rect 25872 26843 25924 26852
rect 25872 26809 25906 26843
rect 25906 26809 25924 26843
rect 25872 26800 25924 26809
rect 7114 26630 7166 26682
rect 7178 26630 7230 26682
rect 7242 26630 7294 26682
rect 7306 26630 7358 26682
rect 7370 26630 7422 26682
rect 13830 26630 13882 26682
rect 13894 26630 13946 26682
rect 13958 26630 14010 26682
rect 14022 26630 14074 26682
rect 14086 26630 14138 26682
rect 20546 26630 20598 26682
rect 20610 26630 20662 26682
rect 20674 26630 20726 26682
rect 20738 26630 20790 26682
rect 20802 26630 20854 26682
rect 27262 26630 27314 26682
rect 27326 26630 27378 26682
rect 27390 26630 27442 26682
rect 27454 26630 27506 26682
rect 27518 26630 27570 26682
rect 1124 26571 1176 26580
rect 1124 26537 1133 26571
rect 1133 26537 1167 26571
rect 1167 26537 1176 26571
rect 1124 26528 1176 26537
rect 2228 26528 2280 26580
rect 2780 26571 2832 26580
rect 2780 26537 2789 26571
rect 2789 26537 2823 26571
rect 2823 26537 2832 26571
rect 2780 26528 2832 26537
rect 5632 26528 5684 26580
rect 6184 26528 6236 26580
rect 8116 26528 8168 26580
rect 11428 26571 11480 26580
rect 11428 26537 11437 26571
rect 11437 26537 11471 26571
rect 11471 26537 11480 26571
rect 11428 26528 11480 26537
rect 14280 26528 14332 26580
rect 2320 26392 2372 26444
rect 3056 26392 3108 26444
rect 3148 26435 3200 26444
rect 3148 26401 3157 26435
rect 3157 26401 3191 26435
rect 3191 26401 3200 26435
rect 3148 26392 3200 26401
rect 4344 26392 4396 26444
rect 5448 26392 5500 26444
rect 5816 26435 5868 26444
rect 5816 26401 5825 26435
rect 5825 26401 5859 26435
rect 5859 26401 5868 26435
rect 5816 26392 5868 26401
rect 3516 26324 3568 26376
rect 6092 26435 6144 26444
rect 6092 26401 6101 26435
rect 6101 26401 6135 26435
rect 6135 26401 6144 26435
rect 6092 26392 6144 26401
rect 6184 26435 6236 26444
rect 6184 26401 6193 26435
rect 6193 26401 6227 26435
rect 6227 26401 6236 26435
rect 6184 26392 6236 26401
rect 6460 26392 6512 26444
rect 8300 26392 8352 26444
rect 9956 26460 10008 26512
rect 11704 26460 11756 26512
rect 2412 26256 2464 26308
rect 3332 26256 3384 26308
rect 4160 26256 4212 26308
rect 6368 26299 6420 26308
rect 6368 26265 6377 26299
rect 6377 26265 6411 26299
rect 6411 26265 6420 26299
rect 6368 26256 6420 26265
rect 4620 26188 4672 26240
rect 4988 26188 5040 26240
rect 9220 26435 9272 26444
rect 9220 26401 9229 26435
rect 9229 26401 9263 26435
rect 9263 26401 9272 26435
rect 9220 26392 9272 26401
rect 9588 26392 9640 26444
rect 10048 26392 10100 26444
rect 10232 26392 10284 26444
rect 11612 26435 11664 26444
rect 11612 26401 11621 26435
rect 11621 26401 11655 26435
rect 11655 26401 11664 26435
rect 11612 26392 11664 26401
rect 12072 26435 12124 26444
rect 12072 26401 12081 26435
rect 12081 26401 12115 26435
rect 12115 26401 12124 26435
rect 12072 26392 12124 26401
rect 11428 26324 11480 26376
rect 12440 26392 12492 26444
rect 12716 26435 12768 26444
rect 12716 26401 12725 26435
rect 12725 26401 12759 26435
rect 12759 26401 12768 26435
rect 12716 26392 12768 26401
rect 12992 26435 13044 26444
rect 12992 26401 13001 26435
rect 13001 26401 13035 26435
rect 13035 26401 13044 26435
rect 12992 26392 13044 26401
rect 14740 26392 14792 26444
rect 15660 26435 15712 26444
rect 15660 26401 15669 26435
rect 15669 26401 15703 26435
rect 15703 26401 15712 26435
rect 15660 26392 15712 26401
rect 16580 26528 16632 26580
rect 16672 26528 16724 26580
rect 21640 26528 21692 26580
rect 22560 26528 22612 26580
rect 23756 26528 23808 26580
rect 25872 26528 25924 26580
rect 16304 26435 16356 26444
rect 16304 26401 16313 26435
rect 16313 26401 16347 26435
rect 16347 26401 16356 26435
rect 16304 26392 16356 26401
rect 16672 26435 16724 26444
rect 16672 26401 16681 26435
rect 16681 26401 16715 26435
rect 16715 26401 16724 26435
rect 16672 26392 16724 26401
rect 17868 26392 17920 26444
rect 21088 26460 21140 26512
rect 18236 26435 18288 26444
rect 18236 26401 18245 26435
rect 18245 26401 18279 26435
rect 18279 26401 18288 26435
rect 18236 26392 18288 26401
rect 10232 26256 10284 26308
rect 10508 26256 10560 26308
rect 16028 26256 16080 26308
rect 16948 26324 17000 26376
rect 17960 26324 18012 26376
rect 18420 26435 18472 26444
rect 18420 26401 18429 26435
rect 18429 26401 18463 26435
rect 18463 26401 18472 26435
rect 18420 26392 18472 26401
rect 20628 26435 20680 26444
rect 20628 26401 20637 26435
rect 20637 26401 20671 26435
rect 20671 26401 20680 26435
rect 20628 26392 20680 26401
rect 17132 26256 17184 26308
rect 18236 26256 18288 26308
rect 19340 26367 19392 26376
rect 19340 26333 19349 26367
rect 19349 26333 19383 26367
rect 19383 26333 19392 26367
rect 19340 26324 19392 26333
rect 20352 26324 20404 26376
rect 20996 26435 21048 26444
rect 20996 26401 21005 26435
rect 21005 26401 21039 26435
rect 21039 26401 21048 26435
rect 20996 26392 21048 26401
rect 21548 26435 21600 26444
rect 21548 26401 21557 26435
rect 21557 26401 21591 26435
rect 21591 26401 21600 26435
rect 21548 26392 21600 26401
rect 21824 26435 21876 26444
rect 21824 26401 21833 26435
rect 21833 26401 21867 26435
rect 21867 26401 21876 26435
rect 21824 26392 21876 26401
rect 23756 26392 23808 26444
rect 19708 26256 19760 26308
rect 6828 26188 6880 26240
rect 8576 26231 8628 26240
rect 8576 26197 8585 26231
rect 8585 26197 8619 26231
rect 8619 26197 8628 26231
rect 8576 26188 8628 26197
rect 8668 26188 8720 26240
rect 9680 26188 9732 26240
rect 10968 26188 11020 26240
rect 11888 26231 11940 26240
rect 11888 26197 11897 26231
rect 11897 26197 11931 26231
rect 11931 26197 11940 26231
rect 11888 26188 11940 26197
rect 16396 26188 16448 26240
rect 18604 26231 18656 26240
rect 18604 26197 18613 26231
rect 18613 26197 18647 26231
rect 18647 26197 18656 26231
rect 18604 26188 18656 26197
rect 20168 26188 20220 26240
rect 21456 26367 21508 26376
rect 21456 26333 21465 26367
rect 21465 26333 21499 26367
rect 21499 26333 21508 26367
rect 21456 26324 21508 26333
rect 22284 26324 22336 26376
rect 25044 26503 25096 26512
rect 25044 26469 25053 26503
rect 25053 26469 25087 26503
rect 25087 26469 25096 26503
rect 25044 26460 25096 26469
rect 25596 26435 25648 26444
rect 25596 26401 25605 26435
rect 25605 26401 25639 26435
rect 25639 26401 25648 26435
rect 25596 26392 25648 26401
rect 25044 26324 25096 26376
rect 22192 26256 22244 26308
rect 24308 26256 24360 26308
rect 20904 26231 20956 26240
rect 20904 26197 20913 26231
rect 20913 26197 20947 26231
rect 20947 26197 20956 26231
rect 20904 26188 20956 26197
rect 23388 26188 23440 26240
rect 24032 26231 24084 26240
rect 24032 26197 24041 26231
rect 24041 26197 24075 26231
rect 24075 26197 24084 26231
rect 24032 26188 24084 26197
rect 24676 26231 24728 26240
rect 24676 26197 24685 26231
rect 24685 26197 24719 26231
rect 24719 26197 24728 26231
rect 24676 26188 24728 26197
rect 3756 26086 3808 26138
rect 3820 26086 3872 26138
rect 3884 26086 3936 26138
rect 3948 26086 4000 26138
rect 4012 26086 4064 26138
rect 10472 26086 10524 26138
rect 10536 26086 10588 26138
rect 10600 26086 10652 26138
rect 10664 26086 10716 26138
rect 10728 26086 10780 26138
rect 17188 26086 17240 26138
rect 17252 26086 17304 26138
rect 17316 26086 17368 26138
rect 17380 26086 17432 26138
rect 17444 26086 17496 26138
rect 23904 26086 23956 26138
rect 23968 26086 24020 26138
rect 24032 26086 24084 26138
rect 24096 26086 24148 26138
rect 24160 26086 24212 26138
rect 7012 26027 7064 26036
rect 7012 25993 7021 26027
rect 7021 25993 7055 26027
rect 7055 25993 7064 26027
rect 7012 25984 7064 25993
rect 8576 25984 8628 26036
rect 2780 25916 2832 25968
rect 9772 25984 9824 26036
rect 10232 25984 10284 26036
rect 11704 25984 11756 26036
rect 10968 25916 11020 25968
rect 11060 25916 11112 25968
rect 14832 25984 14884 26036
rect 15844 25984 15896 26036
rect 16396 26027 16448 26036
rect 16396 25993 16405 26027
rect 16405 25993 16439 26027
rect 16439 25993 16448 26027
rect 16396 25984 16448 25993
rect 20812 25984 20864 26036
rect 20996 25984 21048 26036
rect 22008 25984 22060 26036
rect 23756 25984 23808 26036
rect 24032 26027 24084 26036
rect 24032 25993 24041 26027
rect 24041 25993 24075 26027
rect 24075 25993 24084 26027
rect 24032 25984 24084 25993
rect 24676 26027 24728 26036
rect 24676 25993 24685 26027
rect 24685 25993 24719 26027
rect 24719 25993 24728 26027
rect 24676 25984 24728 25993
rect 25044 25984 25096 26036
rect 16672 25916 16724 25968
rect 2412 25848 2464 25900
rect 2688 25848 2740 25900
rect 4988 25891 5040 25900
rect 4988 25857 4997 25891
rect 4997 25857 5031 25891
rect 5031 25857 5040 25891
rect 4988 25848 5040 25857
rect 6920 25848 6972 25900
rect 2872 25823 2924 25832
rect 2872 25789 2881 25823
rect 2881 25789 2915 25823
rect 2915 25789 2924 25823
rect 2872 25780 2924 25789
rect 4436 25780 4488 25832
rect 5080 25823 5132 25832
rect 5080 25789 5089 25823
rect 5089 25789 5123 25823
rect 5123 25789 5132 25823
rect 5080 25780 5132 25789
rect 5172 25823 5224 25832
rect 5172 25789 5181 25823
rect 5181 25789 5215 25823
rect 5215 25789 5224 25823
rect 5172 25780 5224 25789
rect 6276 25780 6328 25832
rect 7012 25780 7064 25832
rect 9404 25848 9456 25900
rect 7472 25780 7524 25832
rect 3240 25755 3292 25764
rect 3240 25721 3249 25755
rect 3249 25721 3283 25755
rect 3283 25721 3292 25755
rect 3240 25712 3292 25721
rect 3608 25712 3660 25764
rect 1860 25644 1912 25696
rect 2596 25644 2648 25696
rect 3056 25687 3108 25696
rect 3056 25653 3065 25687
rect 3065 25653 3099 25687
rect 3099 25653 3108 25687
rect 3056 25644 3108 25653
rect 4252 25644 4304 25696
rect 7840 25755 7892 25764
rect 7840 25721 7849 25755
rect 7849 25721 7883 25755
rect 7883 25721 7892 25755
rect 7840 25712 7892 25721
rect 8300 25780 8352 25832
rect 8392 25823 8444 25832
rect 8392 25789 8401 25823
rect 8401 25789 8435 25823
rect 8435 25789 8444 25823
rect 8392 25780 8444 25789
rect 8668 25823 8720 25832
rect 8668 25789 8702 25823
rect 8702 25789 8720 25823
rect 8668 25780 8720 25789
rect 10140 25823 10192 25832
rect 10140 25789 10149 25823
rect 10149 25789 10183 25823
rect 10183 25789 10192 25823
rect 10140 25780 10192 25789
rect 10876 25848 10928 25900
rect 11152 25848 11204 25900
rect 12624 25848 12676 25900
rect 14832 25848 14884 25900
rect 15752 25848 15804 25900
rect 16764 25891 16816 25900
rect 16764 25857 16773 25891
rect 16773 25857 16807 25891
rect 16807 25857 16816 25891
rect 16764 25848 16816 25857
rect 18420 25848 18472 25900
rect 18696 25891 18748 25900
rect 18696 25857 18705 25891
rect 18705 25857 18739 25891
rect 18739 25857 18748 25891
rect 18696 25848 18748 25857
rect 11244 25780 11296 25832
rect 12808 25823 12860 25832
rect 12808 25789 12817 25823
rect 12817 25789 12851 25823
rect 12851 25789 12860 25823
rect 12808 25780 12860 25789
rect 15476 25823 15528 25832
rect 15476 25789 15485 25823
rect 15485 25789 15519 25823
rect 15519 25789 15528 25823
rect 15476 25780 15528 25789
rect 16028 25780 16080 25832
rect 16580 25823 16632 25832
rect 16580 25789 16589 25823
rect 16589 25789 16623 25823
rect 16623 25789 16632 25823
rect 16580 25780 16632 25789
rect 17868 25823 17920 25832
rect 17868 25789 17877 25823
rect 17877 25789 17911 25823
rect 17911 25789 17920 25823
rect 17868 25780 17920 25789
rect 18144 25780 18196 25832
rect 18236 25823 18288 25832
rect 18236 25789 18245 25823
rect 18245 25789 18279 25823
rect 18279 25789 18288 25823
rect 18236 25780 18288 25789
rect 18604 25780 18656 25832
rect 20260 25780 20312 25832
rect 20628 25780 20680 25832
rect 7932 25644 7984 25696
rect 9220 25712 9272 25764
rect 9864 25712 9916 25764
rect 10324 25712 10376 25764
rect 13636 25712 13688 25764
rect 17960 25755 18012 25764
rect 17960 25721 17969 25755
rect 17969 25721 18003 25755
rect 18003 25721 18012 25755
rect 17960 25712 18012 25721
rect 9404 25644 9456 25696
rect 10048 25644 10100 25696
rect 12992 25644 13044 25696
rect 15016 25687 15068 25696
rect 15016 25653 15025 25687
rect 15025 25653 15059 25687
rect 15059 25653 15068 25687
rect 15016 25644 15068 25653
rect 17684 25687 17736 25696
rect 17684 25653 17693 25687
rect 17693 25653 17727 25687
rect 17727 25653 17736 25687
rect 17684 25644 17736 25653
rect 20352 25712 20404 25764
rect 21456 25916 21508 25968
rect 24308 25959 24360 25968
rect 24308 25925 24317 25959
rect 24317 25925 24351 25959
rect 24351 25925 24360 25959
rect 24308 25916 24360 25925
rect 25320 25848 25372 25900
rect 20904 25823 20956 25832
rect 20904 25789 20913 25823
rect 20913 25789 20947 25823
rect 20947 25789 20956 25823
rect 20904 25780 20956 25789
rect 20996 25823 21048 25832
rect 20996 25789 21005 25823
rect 21005 25789 21039 25823
rect 21039 25789 21048 25823
rect 20996 25780 21048 25789
rect 20168 25644 20220 25696
rect 23388 25823 23440 25832
rect 23388 25789 23406 25823
rect 23406 25789 23440 25823
rect 23388 25780 23440 25789
rect 25136 25780 25188 25832
rect 23388 25644 23440 25696
rect 24676 25687 24728 25696
rect 24676 25653 24685 25687
rect 24685 25653 24719 25687
rect 24719 25653 24728 25687
rect 24676 25644 24728 25653
rect 25044 25712 25096 25764
rect 25228 25712 25280 25764
rect 7114 25542 7166 25594
rect 7178 25542 7230 25594
rect 7242 25542 7294 25594
rect 7306 25542 7358 25594
rect 7370 25542 7422 25594
rect 13830 25542 13882 25594
rect 13894 25542 13946 25594
rect 13958 25542 14010 25594
rect 14022 25542 14074 25594
rect 14086 25542 14138 25594
rect 20546 25542 20598 25594
rect 20610 25542 20662 25594
rect 20674 25542 20726 25594
rect 20738 25542 20790 25594
rect 20802 25542 20854 25594
rect 27262 25542 27314 25594
rect 27326 25542 27378 25594
rect 27390 25542 27442 25594
rect 27454 25542 27506 25594
rect 27518 25542 27570 25594
rect 848 25347 900 25356
rect 848 25313 857 25347
rect 857 25313 891 25347
rect 891 25313 900 25347
rect 848 25304 900 25313
rect 1124 25347 1176 25356
rect 1124 25313 1158 25347
rect 1158 25313 1176 25347
rect 1124 25304 1176 25313
rect 2412 25304 2464 25356
rect 2688 25440 2740 25492
rect 4436 25483 4488 25492
rect 4436 25449 4445 25483
rect 4445 25449 4479 25483
rect 4479 25449 4488 25483
rect 4436 25440 4488 25449
rect 5540 25440 5592 25492
rect 7840 25440 7892 25492
rect 10048 25440 10100 25492
rect 3608 25372 3660 25424
rect 6920 25372 6972 25424
rect 8300 25372 8352 25424
rect 11060 25372 11112 25424
rect 11888 25372 11940 25424
rect 12072 25440 12124 25492
rect 13636 25440 13688 25492
rect 3056 25347 3108 25356
rect 3056 25313 3090 25347
rect 3090 25313 3108 25347
rect 2136 25236 2188 25288
rect 3056 25304 3108 25313
rect 4988 25347 5040 25356
rect 4988 25313 4997 25347
rect 4997 25313 5031 25347
rect 5031 25313 5040 25347
rect 4988 25304 5040 25313
rect 5080 25347 5132 25356
rect 5080 25313 5089 25347
rect 5089 25313 5123 25347
rect 5123 25313 5132 25347
rect 5080 25304 5132 25313
rect 7012 25347 7064 25356
rect 7012 25313 7021 25347
rect 7021 25313 7055 25347
rect 7055 25313 7064 25347
rect 7012 25304 7064 25313
rect 7656 25304 7708 25356
rect 4896 25236 4948 25288
rect 5356 25279 5408 25288
rect 5356 25245 5365 25279
rect 5365 25245 5399 25279
rect 5399 25245 5408 25279
rect 5356 25236 5408 25245
rect 6920 25279 6972 25288
rect 6920 25245 6929 25279
rect 6929 25245 6963 25279
rect 6963 25245 6972 25279
rect 6920 25236 6972 25245
rect 9588 25304 9640 25356
rect 9680 25347 9732 25356
rect 9680 25313 9689 25347
rect 9689 25313 9723 25347
rect 9723 25313 9732 25347
rect 9680 25304 9732 25313
rect 10140 25304 10192 25356
rect 11152 25347 11204 25356
rect 11152 25313 11161 25347
rect 11161 25313 11195 25347
rect 11195 25313 11204 25347
rect 11152 25304 11204 25313
rect 12992 25415 13044 25424
rect 12992 25381 13001 25415
rect 13001 25381 13035 25415
rect 13035 25381 13044 25415
rect 12992 25372 13044 25381
rect 14004 25304 14056 25356
rect 15016 25440 15068 25492
rect 19340 25440 19392 25492
rect 20260 25483 20312 25492
rect 20260 25449 20269 25483
rect 20269 25449 20303 25483
rect 20303 25449 20312 25483
rect 20260 25440 20312 25449
rect 21364 25483 21416 25492
rect 21364 25449 21373 25483
rect 21373 25449 21407 25483
rect 21407 25449 21416 25483
rect 21364 25440 21416 25449
rect 22100 25440 22152 25492
rect 22744 25440 22796 25492
rect 23388 25483 23440 25492
rect 23388 25449 23397 25483
rect 23397 25449 23431 25483
rect 23431 25449 23440 25483
rect 23388 25440 23440 25449
rect 17684 25372 17736 25424
rect 14924 25304 14976 25356
rect 18972 25304 19024 25356
rect 22008 25372 22060 25424
rect 24308 25440 24360 25492
rect 25136 25440 25188 25492
rect 25228 25483 25280 25492
rect 25228 25449 25237 25483
rect 25237 25449 25271 25483
rect 25271 25449 25280 25483
rect 25228 25440 25280 25449
rect 21272 25304 21324 25356
rect 22284 25347 22336 25356
rect 22284 25313 22293 25347
rect 22293 25313 22327 25347
rect 22327 25313 22336 25347
rect 22284 25304 22336 25313
rect 22468 25347 22520 25356
rect 22468 25313 22477 25347
rect 22477 25313 22511 25347
rect 22511 25313 22520 25347
rect 22468 25304 22520 25313
rect 8852 25236 8904 25288
rect 15016 25279 15068 25288
rect 15016 25245 15025 25279
rect 15025 25245 15059 25279
rect 15059 25245 15068 25279
rect 15016 25236 15068 25245
rect 17040 25236 17092 25288
rect 17776 25279 17828 25288
rect 17776 25245 17785 25279
rect 17785 25245 17819 25279
rect 17819 25245 17828 25279
rect 17776 25236 17828 25245
rect 21732 25279 21784 25288
rect 21732 25245 21741 25279
rect 21741 25245 21775 25279
rect 21775 25245 21784 25279
rect 21732 25236 21784 25245
rect 22376 25279 22428 25288
rect 22376 25245 22385 25279
rect 22385 25245 22419 25279
rect 22419 25245 22428 25279
rect 22376 25236 22428 25245
rect 24676 25415 24728 25424
rect 9680 25168 9732 25220
rect 10324 25168 10376 25220
rect 23112 25236 23164 25288
rect 23756 25236 23808 25288
rect 24676 25381 24685 25415
rect 24685 25381 24719 25415
rect 24719 25381 24728 25415
rect 24676 25372 24728 25381
rect 24860 25372 24912 25424
rect 24308 25304 24360 25356
rect 25044 25347 25096 25356
rect 25044 25313 25053 25347
rect 25053 25313 25087 25347
rect 25087 25313 25096 25347
rect 25044 25304 25096 25313
rect 25872 25304 25924 25356
rect 25412 25236 25464 25288
rect 2228 25143 2280 25152
rect 2228 25109 2237 25143
rect 2237 25109 2271 25143
rect 2271 25109 2280 25143
rect 2228 25100 2280 25109
rect 2688 25143 2740 25152
rect 2688 25109 2697 25143
rect 2697 25109 2731 25143
rect 2731 25109 2740 25143
rect 2688 25100 2740 25109
rect 4620 25143 4672 25152
rect 4620 25109 4629 25143
rect 4629 25109 4663 25143
rect 4663 25109 4672 25143
rect 4620 25100 4672 25109
rect 7564 25143 7616 25152
rect 7564 25109 7573 25143
rect 7573 25109 7607 25143
rect 7607 25109 7616 25143
rect 7564 25100 7616 25109
rect 10968 25100 11020 25152
rect 12716 25100 12768 25152
rect 17684 25100 17736 25152
rect 23664 25100 23716 25152
rect 24032 25100 24084 25152
rect 3756 24998 3808 25050
rect 3820 24998 3872 25050
rect 3884 24998 3936 25050
rect 3948 24998 4000 25050
rect 4012 24998 4064 25050
rect 10472 24998 10524 25050
rect 10536 24998 10588 25050
rect 10600 24998 10652 25050
rect 10664 24998 10716 25050
rect 10728 24998 10780 25050
rect 17188 24998 17240 25050
rect 17252 24998 17304 25050
rect 17316 24998 17368 25050
rect 17380 24998 17432 25050
rect 17444 24998 17496 25050
rect 23904 24998 23956 25050
rect 23968 24998 24020 25050
rect 24032 24998 24084 25050
rect 24096 24998 24148 25050
rect 24160 24998 24212 25050
rect 1124 24896 1176 24948
rect 1952 24896 2004 24948
rect 2596 24939 2648 24948
rect 2596 24905 2605 24939
rect 2605 24905 2639 24939
rect 2639 24905 2648 24939
rect 2596 24896 2648 24905
rect 2872 24896 2924 24948
rect 4160 24939 4212 24948
rect 4160 24905 4169 24939
rect 4169 24905 4203 24939
rect 4203 24905 4212 24939
rect 4160 24896 4212 24905
rect 5080 24896 5132 24948
rect 5356 24896 5408 24948
rect 9588 24896 9640 24948
rect 10140 24896 10192 24948
rect 11244 24896 11296 24948
rect 14556 24939 14608 24948
rect 14556 24905 14565 24939
rect 14565 24905 14599 24939
rect 14599 24905 14608 24939
rect 14556 24896 14608 24905
rect 2596 24760 2648 24812
rect 2780 24760 2832 24812
rect 3056 24760 3108 24812
rect 4988 24803 5040 24812
rect 4988 24769 4997 24803
rect 4997 24769 5031 24803
rect 5031 24769 5040 24803
rect 4988 24760 5040 24769
rect 2228 24692 2280 24744
rect 3516 24692 3568 24744
rect 1860 24667 1912 24676
rect 1860 24633 1887 24667
rect 1887 24633 1912 24667
rect 1860 24624 1912 24633
rect 2044 24667 2096 24676
rect 2044 24633 2053 24667
rect 2053 24633 2087 24667
rect 2087 24633 2096 24667
rect 2044 24624 2096 24633
rect 2688 24624 2740 24676
rect 4896 24735 4948 24744
rect 4896 24701 4905 24735
rect 4905 24701 4939 24735
rect 4939 24701 4948 24735
rect 4896 24692 4948 24701
rect 8392 24760 8444 24812
rect 10048 24760 10100 24812
rect 11152 24760 11204 24812
rect 13360 24760 13412 24812
rect 6184 24624 6236 24676
rect 7472 24692 7524 24744
rect 7840 24735 7892 24744
rect 7840 24701 7849 24735
rect 7849 24701 7883 24735
rect 7883 24701 7892 24735
rect 7840 24692 7892 24701
rect 9496 24692 9548 24744
rect 8760 24624 8812 24676
rect 9312 24624 9364 24676
rect 6276 24556 6328 24608
rect 6736 24556 6788 24608
rect 10324 24624 10376 24676
rect 14004 24692 14056 24744
rect 14464 24692 14516 24744
rect 12624 24624 12676 24676
rect 14648 24692 14700 24744
rect 15476 24896 15528 24948
rect 15752 24896 15804 24948
rect 22376 24896 22428 24948
rect 17684 24828 17736 24880
rect 17776 24828 17828 24880
rect 18144 24828 18196 24880
rect 22192 24828 22244 24880
rect 15568 24760 15620 24812
rect 15660 24735 15712 24744
rect 15660 24701 15669 24735
rect 15669 24701 15703 24735
rect 15703 24701 15712 24735
rect 15660 24692 15712 24701
rect 15936 24735 15988 24744
rect 15936 24701 15945 24735
rect 15945 24701 15979 24735
rect 15979 24701 15988 24735
rect 15936 24692 15988 24701
rect 17040 24692 17092 24744
rect 23756 24896 23808 24948
rect 11152 24556 11204 24608
rect 13360 24599 13412 24608
rect 13360 24565 13369 24599
rect 13369 24565 13403 24599
rect 13403 24565 13412 24599
rect 13360 24556 13412 24565
rect 13452 24556 13504 24608
rect 14832 24599 14884 24608
rect 14832 24565 14841 24599
rect 14841 24565 14875 24599
rect 14875 24565 14884 24599
rect 14832 24556 14884 24565
rect 15108 24599 15160 24608
rect 15108 24565 15117 24599
rect 15117 24565 15151 24599
rect 15151 24565 15160 24599
rect 15108 24556 15160 24565
rect 17960 24692 18012 24744
rect 19064 24735 19116 24744
rect 19064 24701 19073 24735
rect 19073 24701 19107 24735
rect 19107 24701 19116 24735
rect 19064 24692 19116 24701
rect 16948 24556 17000 24608
rect 18420 24624 18472 24676
rect 23112 24692 23164 24744
rect 17408 24599 17460 24608
rect 17408 24565 17417 24599
rect 17417 24565 17451 24599
rect 17451 24565 17460 24599
rect 17408 24556 17460 24565
rect 21364 24624 21416 24676
rect 21732 24624 21784 24676
rect 23756 24624 23808 24676
rect 24032 24667 24084 24676
rect 24032 24633 24057 24667
rect 24057 24633 24084 24667
rect 24492 24760 24544 24812
rect 24400 24692 24452 24744
rect 24676 24692 24728 24744
rect 24860 24735 24912 24744
rect 24860 24701 24893 24735
rect 24893 24701 24912 24735
rect 24860 24692 24912 24701
rect 24032 24624 24084 24633
rect 25320 24735 25372 24744
rect 25320 24701 25329 24735
rect 25329 24701 25363 24735
rect 25363 24701 25372 24735
rect 25320 24692 25372 24701
rect 25412 24692 25464 24744
rect 26056 24624 26108 24676
rect 20904 24556 20956 24608
rect 23388 24556 23440 24608
rect 24308 24556 24360 24608
rect 24768 24599 24820 24608
rect 24768 24565 24777 24599
rect 24777 24565 24811 24599
rect 24811 24565 24820 24599
rect 24768 24556 24820 24565
rect 25136 24556 25188 24608
rect 25780 24556 25832 24608
rect 26884 24556 26936 24608
rect 7114 24454 7166 24506
rect 7178 24454 7230 24506
rect 7242 24454 7294 24506
rect 7306 24454 7358 24506
rect 7370 24454 7422 24506
rect 13830 24454 13882 24506
rect 13894 24454 13946 24506
rect 13958 24454 14010 24506
rect 14022 24454 14074 24506
rect 14086 24454 14138 24506
rect 20546 24454 20598 24506
rect 20610 24454 20662 24506
rect 20674 24454 20726 24506
rect 20738 24454 20790 24506
rect 20802 24454 20854 24506
rect 27262 24454 27314 24506
rect 27326 24454 27378 24506
rect 27390 24454 27442 24506
rect 27454 24454 27506 24506
rect 27518 24454 27570 24506
rect 6184 24395 6236 24404
rect 6184 24361 6193 24395
rect 6193 24361 6227 24395
rect 6227 24361 6236 24395
rect 6184 24352 6236 24361
rect 6276 24352 6328 24404
rect 7840 24352 7892 24404
rect 8852 24395 8904 24404
rect 8852 24361 8861 24395
rect 8861 24361 8895 24395
rect 8895 24361 8904 24395
rect 8852 24352 8904 24361
rect 9312 24395 9364 24404
rect 9312 24361 9321 24395
rect 9321 24361 9355 24395
rect 9355 24361 9364 24395
rect 9312 24352 9364 24361
rect 9956 24352 10008 24404
rect 10324 24395 10376 24404
rect 10324 24361 10341 24395
rect 10341 24361 10376 24395
rect 10324 24352 10376 24361
rect 12624 24395 12676 24404
rect 12624 24361 12633 24395
rect 12633 24361 12667 24395
rect 12667 24361 12676 24395
rect 12624 24352 12676 24361
rect 12716 24352 12768 24404
rect 14188 24352 14240 24404
rect 15568 24395 15620 24404
rect 15568 24361 15577 24395
rect 15577 24361 15611 24395
rect 15611 24361 15620 24395
rect 15568 24352 15620 24361
rect 15660 24352 15712 24404
rect 17408 24352 17460 24404
rect 19064 24352 19116 24404
rect 22192 24352 22244 24404
rect 2596 24284 2648 24336
rect 6920 24284 6972 24336
rect 1860 24055 1912 24064
rect 1860 24021 1869 24055
rect 1869 24021 1903 24055
rect 1903 24021 1912 24055
rect 1860 24012 1912 24021
rect 2320 24216 2372 24268
rect 2872 24259 2924 24268
rect 2872 24225 2881 24259
rect 2881 24225 2915 24259
rect 2915 24225 2924 24259
rect 2872 24216 2924 24225
rect 4804 24259 4856 24268
rect 4804 24225 4813 24259
rect 4813 24225 4847 24259
rect 4847 24225 4856 24259
rect 4804 24216 4856 24225
rect 2136 24148 2188 24200
rect 3608 24080 3660 24132
rect 5448 24080 5500 24132
rect 6736 24259 6788 24268
rect 6736 24225 6745 24259
rect 6745 24225 6779 24259
rect 6779 24225 6788 24259
rect 6736 24216 6788 24225
rect 6828 24259 6880 24268
rect 6828 24225 6837 24259
rect 6837 24225 6871 24259
rect 6871 24225 6880 24259
rect 6828 24216 6880 24225
rect 7196 24259 7248 24268
rect 7196 24225 7205 24259
rect 7205 24225 7239 24259
rect 7239 24225 7248 24259
rect 7196 24216 7248 24225
rect 7564 24284 7616 24336
rect 8024 24216 8076 24268
rect 8300 24216 8352 24268
rect 9404 24216 9456 24268
rect 9680 24259 9732 24268
rect 9680 24225 9689 24259
rect 9689 24225 9723 24259
rect 9723 24225 9732 24259
rect 9680 24216 9732 24225
rect 10048 24216 10100 24268
rect 11152 24216 11204 24268
rect 13452 24284 13504 24336
rect 7380 24148 7432 24200
rect 7472 24191 7524 24200
rect 7472 24157 7481 24191
rect 7481 24157 7515 24191
rect 7515 24157 7524 24191
rect 7472 24148 7524 24157
rect 7012 24080 7064 24132
rect 7196 24080 7248 24132
rect 10232 24148 10284 24200
rect 10968 24080 11020 24132
rect 11704 24123 11756 24132
rect 11704 24089 11713 24123
rect 11713 24089 11747 24123
rect 11747 24089 11756 24123
rect 11704 24080 11756 24089
rect 13084 24259 13136 24268
rect 13084 24225 13093 24259
rect 13093 24225 13127 24259
rect 13127 24225 13136 24259
rect 13084 24216 13136 24225
rect 15936 24284 15988 24336
rect 14832 24216 14884 24268
rect 15016 24216 15068 24268
rect 16212 24216 16264 24268
rect 16396 24148 16448 24200
rect 2688 24012 2740 24064
rect 2780 24055 2832 24064
rect 2780 24021 2789 24055
rect 2789 24021 2823 24055
rect 2823 24021 2832 24055
rect 2780 24012 2832 24021
rect 4160 24012 4212 24064
rect 4896 24012 4948 24064
rect 8760 24012 8812 24064
rect 10140 24055 10192 24064
rect 10140 24021 10149 24055
rect 10149 24021 10183 24055
rect 10183 24021 10192 24055
rect 10140 24012 10192 24021
rect 10876 24012 10928 24064
rect 12992 24012 13044 24064
rect 13728 24012 13780 24064
rect 16488 24012 16540 24064
rect 18144 24148 18196 24200
rect 18972 24148 19024 24200
rect 20444 24216 20496 24268
rect 20904 24216 20956 24268
rect 20996 24216 21048 24268
rect 21824 24284 21876 24336
rect 24308 24352 24360 24404
rect 24400 24395 24452 24404
rect 24400 24361 24409 24395
rect 24409 24361 24443 24395
rect 24443 24361 24452 24395
rect 24400 24352 24452 24361
rect 25964 24352 26016 24404
rect 26056 24395 26108 24404
rect 26056 24361 26065 24395
rect 26065 24361 26099 24395
rect 26099 24361 26108 24395
rect 26056 24352 26108 24361
rect 23388 24327 23440 24336
rect 23388 24293 23397 24327
rect 23397 24293 23431 24327
rect 23431 24293 23440 24327
rect 23388 24284 23440 24293
rect 24492 24284 24544 24336
rect 24860 24327 24912 24336
rect 24860 24293 24869 24327
rect 24869 24293 24903 24327
rect 24903 24293 24912 24327
rect 24860 24284 24912 24293
rect 25228 24284 25280 24336
rect 25596 24327 25648 24336
rect 25596 24293 25605 24327
rect 25605 24293 25639 24327
rect 25639 24293 25648 24327
rect 25596 24284 25648 24293
rect 22192 24216 22244 24268
rect 23664 24259 23716 24268
rect 23664 24225 23673 24259
rect 23673 24225 23707 24259
rect 23707 24225 23716 24259
rect 23664 24216 23716 24225
rect 25136 24259 25188 24268
rect 25136 24225 25145 24259
rect 25145 24225 25179 24259
rect 25179 24225 25188 24259
rect 25136 24216 25188 24225
rect 25320 24259 25372 24268
rect 25320 24225 25329 24259
rect 25329 24225 25363 24259
rect 25363 24225 25372 24259
rect 25320 24216 25372 24225
rect 19800 24148 19852 24200
rect 20076 24191 20128 24200
rect 20076 24157 20085 24191
rect 20085 24157 20119 24191
rect 20119 24157 20128 24191
rect 20076 24148 20128 24157
rect 20812 24148 20864 24200
rect 22100 24148 22152 24200
rect 23756 24191 23808 24200
rect 23756 24157 23765 24191
rect 23765 24157 23799 24191
rect 23799 24157 23808 24191
rect 23756 24148 23808 24157
rect 17592 24055 17644 24064
rect 17592 24021 17601 24055
rect 17601 24021 17635 24055
rect 17635 24021 17644 24055
rect 17592 24012 17644 24021
rect 18880 24055 18932 24064
rect 18880 24021 18889 24055
rect 18889 24021 18923 24055
rect 18923 24021 18932 24055
rect 18880 24012 18932 24021
rect 22652 24055 22704 24064
rect 22652 24021 22661 24055
rect 22661 24021 22695 24055
rect 22695 24021 22704 24055
rect 22652 24012 22704 24021
rect 23296 24012 23348 24064
rect 26884 24259 26936 24268
rect 26884 24225 26893 24259
rect 26893 24225 26927 24259
rect 26927 24225 26936 24259
rect 26884 24216 26936 24225
rect 24492 24055 24544 24064
rect 24492 24021 24501 24055
rect 24501 24021 24535 24055
rect 24535 24021 24544 24055
rect 24492 24012 24544 24021
rect 25780 24055 25832 24064
rect 25780 24021 25789 24055
rect 25789 24021 25823 24055
rect 25823 24021 25832 24055
rect 25780 24012 25832 24021
rect 3756 23910 3808 23962
rect 3820 23910 3872 23962
rect 3884 23910 3936 23962
rect 3948 23910 4000 23962
rect 4012 23910 4064 23962
rect 10472 23910 10524 23962
rect 10536 23910 10588 23962
rect 10600 23910 10652 23962
rect 10664 23910 10716 23962
rect 10728 23910 10780 23962
rect 17188 23910 17240 23962
rect 17252 23910 17304 23962
rect 17316 23910 17368 23962
rect 17380 23910 17432 23962
rect 17444 23910 17496 23962
rect 23904 23910 23956 23962
rect 23968 23910 24020 23962
rect 24032 23910 24084 23962
rect 24096 23910 24148 23962
rect 24160 23910 24212 23962
rect 2320 23851 2372 23860
rect 2320 23817 2329 23851
rect 2329 23817 2363 23851
rect 2363 23817 2372 23851
rect 2320 23808 2372 23817
rect 2596 23808 2648 23860
rect 2044 23740 2096 23792
rect 2780 23672 2832 23724
rect 1860 23536 1912 23588
rect 2136 23579 2188 23588
rect 2136 23545 2145 23579
rect 2145 23545 2179 23579
rect 2179 23545 2188 23579
rect 2136 23536 2188 23545
rect 1124 23468 1176 23520
rect 1492 23468 1544 23520
rect 2320 23511 2372 23520
rect 2320 23477 2345 23511
rect 2345 23477 2372 23511
rect 2320 23468 2372 23477
rect 2504 23468 2556 23520
rect 4804 23808 4856 23860
rect 5172 23808 5224 23860
rect 5356 23851 5408 23860
rect 5356 23817 5365 23851
rect 5365 23817 5399 23851
rect 5399 23817 5408 23851
rect 5356 23808 5408 23817
rect 6828 23808 6880 23860
rect 10232 23808 10284 23860
rect 12900 23808 12952 23860
rect 3792 23647 3844 23656
rect 3792 23613 3801 23647
rect 3801 23613 3835 23647
rect 3835 23613 3844 23647
rect 3792 23604 3844 23613
rect 3884 23647 3936 23656
rect 3884 23613 3893 23647
rect 3893 23613 3927 23647
rect 3927 23613 3936 23647
rect 3884 23604 3936 23613
rect 7196 23740 7248 23792
rect 7564 23740 7616 23792
rect 13728 23851 13780 23860
rect 13728 23817 13737 23851
rect 13737 23817 13771 23851
rect 13771 23817 13780 23851
rect 13728 23808 13780 23817
rect 14556 23808 14608 23860
rect 14648 23851 14700 23860
rect 14648 23817 14657 23851
rect 14657 23817 14691 23851
rect 14691 23817 14700 23851
rect 14648 23808 14700 23817
rect 18144 23851 18196 23860
rect 18144 23817 18153 23851
rect 18153 23817 18187 23851
rect 18187 23817 18196 23851
rect 20812 23851 20864 23860
rect 18144 23808 18196 23817
rect 20812 23817 20821 23851
rect 20821 23817 20855 23851
rect 20855 23817 20864 23851
rect 20812 23808 20864 23817
rect 4528 23672 4580 23724
rect 2688 23536 2740 23588
rect 2872 23536 2924 23588
rect 3700 23536 3752 23588
rect 4344 23647 4396 23656
rect 4344 23613 4353 23647
rect 4353 23613 4387 23647
rect 4387 23613 4396 23647
rect 4344 23604 4396 23613
rect 4528 23579 4580 23588
rect 4528 23545 4537 23579
rect 4537 23545 4571 23579
rect 4571 23545 4580 23579
rect 4528 23536 4580 23545
rect 4620 23468 4672 23520
rect 4896 23604 4948 23656
rect 4988 23647 5040 23656
rect 4988 23613 4997 23647
rect 4997 23613 5031 23647
rect 5031 23613 5040 23647
rect 4988 23604 5040 23613
rect 5080 23647 5132 23656
rect 5080 23613 5089 23647
rect 5089 23613 5123 23647
rect 5123 23613 5132 23647
rect 5080 23604 5132 23613
rect 5448 23715 5500 23724
rect 5448 23681 5457 23715
rect 5457 23681 5491 23715
rect 5491 23681 5500 23715
rect 5448 23672 5500 23681
rect 9496 23715 9548 23724
rect 9496 23681 9505 23715
rect 9505 23681 9539 23715
rect 9539 23681 9548 23715
rect 9496 23672 9548 23681
rect 10508 23672 10560 23724
rect 10876 23672 10928 23724
rect 6460 23536 6512 23588
rect 7840 23604 7892 23656
rect 11152 23647 11204 23656
rect 11152 23613 11161 23647
rect 11161 23613 11195 23647
rect 11195 23613 11204 23647
rect 11152 23604 11204 23613
rect 11336 23647 11388 23656
rect 11336 23613 11345 23647
rect 11345 23613 11379 23647
rect 11379 23613 11388 23647
rect 11336 23604 11388 23613
rect 12808 23647 12860 23656
rect 12808 23613 12817 23647
rect 12817 23613 12851 23647
rect 12851 23613 12860 23647
rect 12808 23604 12860 23613
rect 13360 23604 13412 23656
rect 9956 23536 10008 23588
rect 11796 23536 11848 23588
rect 11888 23536 11940 23588
rect 14188 23740 14240 23792
rect 15016 23740 15068 23792
rect 15108 23715 15160 23724
rect 15108 23681 15117 23715
rect 15117 23681 15151 23715
rect 15151 23681 15160 23715
rect 15108 23672 15160 23681
rect 19800 23740 19852 23792
rect 20352 23740 20404 23792
rect 15292 23672 15344 23724
rect 17776 23672 17828 23724
rect 21272 23783 21324 23792
rect 21272 23749 21281 23783
rect 21281 23749 21315 23783
rect 21315 23749 21324 23783
rect 21272 23740 21324 23749
rect 21364 23783 21416 23792
rect 21364 23749 21373 23783
rect 21373 23749 21407 23783
rect 21407 23749 21416 23783
rect 21364 23740 21416 23749
rect 14280 23604 14332 23656
rect 16856 23604 16908 23656
rect 18328 23647 18380 23656
rect 18328 23613 18337 23647
rect 18337 23613 18371 23647
rect 18371 23613 18380 23647
rect 18328 23604 18380 23613
rect 20444 23604 20496 23656
rect 20904 23672 20956 23724
rect 7012 23468 7064 23520
rect 7380 23468 7432 23520
rect 7748 23468 7800 23520
rect 10048 23468 10100 23520
rect 12072 23468 12124 23520
rect 12440 23468 12492 23520
rect 13084 23468 13136 23520
rect 15660 23536 15712 23588
rect 16304 23536 16356 23588
rect 14464 23468 14516 23520
rect 15016 23511 15068 23520
rect 15016 23477 15025 23511
rect 15025 23477 15059 23511
rect 15059 23477 15068 23511
rect 15016 23468 15068 23477
rect 15844 23468 15896 23520
rect 20996 23647 21048 23656
rect 20996 23613 21005 23647
rect 21005 23613 21039 23647
rect 21039 23613 21048 23647
rect 20996 23604 21048 23613
rect 21088 23647 21140 23656
rect 21088 23613 21097 23647
rect 21097 23613 21131 23647
rect 21131 23613 21140 23647
rect 21088 23604 21140 23613
rect 20904 23536 20956 23588
rect 21824 23647 21876 23656
rect 21824 23613 21869 23647
rect 21869 23613 21876 23647
rect 21824 23604 21876 23613
rect 21640 23579 21692 23588
rect 21640 23545 21649 23579
rect 21649 23545 21683 23579
rect 21683 23545 21692 23579
rect 21640 23536 21692 23545
rect 20168 23511 20220 23520
rect 20168 23477 20177 23511
rect 20177 23477 20211 23511
rect 20211 23477 20220 23511
rect 20168 23468 20220 23477
rect 21088 23468 21140 23520
rect 21916 23468 21968 23520
rect 23756 23808 23808 23860
rect 23848 23808 23900 23860
rect 24400 23808 24452 23860
rect 25596 23672 25648 23724
rect 25412 23647 25464 23656
rect 25412 23613 25421 23647
rect 25421 23613 25455 23647
rect 25455 23613 25464 23647
rect 25412 23604 25464 23613
rect 25964 23647 26016 23656
rect 25964 23613 25973 23647
rect 25973 23613 26007 23647
rect 26007 23613 26016 23647
rect 25964 23604 26016 23613
rect 26700 23647 26752 23656
rect 26700 23613 26709 23647
rect 26709 23613 26743 23647
rect 26743 23613 26752 23647
rect 26700 23604 26752 23613
rect 22652 23536 22704 23588
rect 24768 23536 24820 23588
rect 22192 23468 22244 23520
rect 25780 23511 25832 23520
rect 25780 23477 25789 23511
rect 25789 23477 25823 23511
rect 25823 23477 25832 23511
rect 25780 23468 25832 23477
rect 7114 23366 7166 23418
rect 7178 23366 7230 23418
rect 7242 23366 7294 23418
rect 7306 23366 7358 23418
rect 7370 23366 7422 23418
rect 13830 23366 13882 23418
rect 13894 23366 13946 23418
rect 13958 23366 14010 23418
rect 14022 23366 14074 23418
rect 14086 23366 14138 23418
rect 20546 23366 20598 23418
rect 20610 23366 20662 23418
rect 20674 23366 20726 23418
rect 20738 23366 20790 23418
rect 20802 23366 20854 23418
rect 27262 23366 27314 23418
rect 27326 23366 27378 23418
rect 27390 23366 27442 23418
rect 27454 23366 27506 23418
rect 27518 23366 27570 23418
rect 2872 23264 2924 23316
rect 2780 23196 2832 23248
rect 1124 23171 1176 23180
rect 1124 23137 1158 23171
rect 1158 23137 1176 23171
rect 1124 23128 1176 23137
rect 2596 23128 2648 23180
rect 3056 23171 3108 23180
rect 3056 23137 3065 23171
rect 3065 23137 3099 23171
rect 3099 23137 3108 23171
rect 3056 23128 3108 23137
rect 3792 23264 3844 23316
rect 5080 23264 5132 23316
rect 6460 23307 6512 23316
rect 6460 23273 6469 23307
rect 6469 23273 6503 23307
rect 6503 23273 6512 23307
rect 6460 23264 6512 23273
rect 4160 23196 4212 23248
rect 848 23103 900 23112
rect 848 23069 857 23103
rect 857 23069 891 23103
rect 891 23069 900 23103
rect 848 23060 900 23069
rect 3332 23060 3384 23112
rect 3700 23128 3752 23180
rect 6092 23196 6144 23248
rect 7564 23264 7616 23316
rect 8576 23264 8628 23316
rect 3608 23060 3660 23112
rect 4344 23128 4396 23180
rect 3516 22992 3568 23044
rect 4436 23103 4488 23112
rect 4436 23069 4445 23103
rect 4445 23069 4479 23103
rect 4479 23069 4488 23103
rect 4436 23060 4488 23069
rect 4804 23171 4856 23180
rect 4804 23137 4813 23171
rect 4813 23137 4847 23171
rect 4847 23137 4856 23171
rect 4804 23128 4856 23137
rect 5908 23171 5960 23180
rect 5908 23137 5917 23171
rect 5917 23137 5951 23171
rect 5951 23137 5960 23171
rect 5908 23128 5960 23137
rect 6184 23171 6236 23180
rect 6184 23137 6193 23171
rect 6193 23137 6227 23171
rect 6227 23137 6236 23171
rect 6184 23128 6236 23137
rect 6736 23171 6788 23180
rect 6736 23137 6745 23171
rect 6745 23137 6779 23171
rect 6779 23137 6788 23171
rect 6736 23128 6788 23137
rect 6920 23196 6972 23248
rect 8300 23196 8352 23248
rect 8760 23196 8812 23248
rect 9956 23307 10008 23316
rect 9956 23273 9965 23307
rect 9965 23273 9999 23307
rect 9999 23273 10008 23307
rect 9956 23264 10008 23273
rect 12716 23264 12768 23316
rect 13728 23264 13780 23316
rect 15016 23264 15068 23316
rect 16672 23264 16724 23316
rect 16856 23264 16908 23316
rect 17592 23264 17644 23316
rect 18328 23264 18380 23316
rect 18880 23307 18932 23316
rect 18880 23273 18889 23307
rect 18889 23273 18923 23307
rect 18923 23273 18932 23307
rect 18880 23264 18932 23273
rect 11796 23239 11848 23248
rect 11796 23205 11805 23239
rect 11805 23205 11839 23239
rect 11839 23205 11848 23239
rect 11796 23196 11848 23205
rect 12532 23196 12584 23248
rect 14188 23196 14240 23248
rect 14556 23196 14608 23248
rect 6276 23060 6328 23112
rect 7012 23171 7064 23180
rect 7012 23137 7021 23171
rect 7021 23137 7055 23171
rect 7055 23137 7064 23171
rect 7012 23128 7064 23137
rect 7104 23171 7156 23180
rect 7104 23137 7113 23171
rect 7113 23137 7147 23171
rect 7147 23137 7156 23171
rect 7104 23128 7156 23137
rect 7564 23128 7616 23180
rect 6644 22992 6696 23044
rect 9496 23128 9548 23180
rect 10140 23171 10192 23180
rect 10140 23137 10149 23171
rect 10149 23137 10183 23171
rect 10183 23137 10192 23171
rect 10140 23128 10192 23137
rect 10324 23171 10376 23180
rect 10324 23137 10333 23171
rect 10333 23137 10367 23171
rect 10367 23137 10376 23171
rect 10324 23128 10376 23137
rect 7840 22992 7892 23044
rect 9680 23060 9732 23112
rect 10048 23060 10100 23112
rect 11888 23128 11940 23180
rect 12072 23128 12124 23180
rect 12348 23128 12400 23180
rect 12900 23171 12952 23180
rect 12900 23137 12909 23171
rect 12909 23137 12943 23171
rect 12943 23137 12952 23171
rect 12900 23128 12952 23137
rect 11428 23060 11480 23112
rect 11520 23060 11572 23112
rect 14372 23128 14424 23180
rect 16580 23196 16632 23248
rect 11336 22992 11388 23044
rect 12348 22992 12400 23044
rect 15752 23171 15804 23180
rect 15752 23137 15761 23171
rect 15761 23137 15795 23171
rect 15795 23137 15804 23171
rect 15752 23128 15804 23137
rect 16304 23128 16356 23180
rect 17684 23196 17736 23248
rect 20996 23264 21048 23316
rect 21916 23307 21968 23316
rect 21916 23273 21925 23307
rect 21925 23273 21959 23307
rect 21959 23273 21968 23307
rect 21916 23264 21968 23273
rect 18144 23128 18196 23180
rect 18788 23171 18840 23180
rect 18788 23137 18797 23171
rect 18797 23137 18831 23171
rect 18831 23137 18840 23171
rect 18788 23128 18840 23137
rect 19616 23128 19668 23180
rect 22192 23239 22244 23248
rect 22192 23205 22201 23239
rect 22201 23205 22235 23239
rect 22235 23205 22244 23239
rect 22192 23196 22244 23205
rect 16396 22992 16448 23044
rect 19340 23060 19392 23112
rect 20904 22992 20956 23044
rect 22100 23171 22152 23180
rect 22100 23137 22109 23171
rect 22109 23137 22143 23171
rect 22143 23137 22152 23171
rect 22100 23128 22152 23137
rect 22284 23171 22336 23180
rect 22284 23137 22293 23171
rect 22293 23137 22327 23171
rect 22327 23137 22336 23171
rect 22284 23128 22336 23137
rect 23296 23264 23348 23316
rect 24676 23307 24728 23316
rect 24676 23273 24685 23307
rect 24685 23273 24719 23307
rect 24719 23273 24728 23307
rect 24676 23264 24728 23273
rect 26700 23264 26752 23316
rect 23848 23171 23900 23180
rect 23848 23137 23857 23171
rect 23857 23137 23891 23171
rect 23891 23137 23900 23171
rect 23848 23128 23900 23137
rect 25136 23196 25188 23248
rect 25596 23128 25648 23180
rect 21640 23060 21692 23112
rect 24584 23060 24636 23112
rect 25044 23060 25096 23112
rect 26884 23060 26936 23112
rect 4528 22924 4580 22976
rect 9128 22924 9180 22976
rect 11704 22924 11756 22976
rect 11796 22924 11848 22976
rect 12992 22924 13044 22976
rect 13176 22924 13228 22976
rect 15476 22924 15528 22976
rect 18880 22924 18932 22976
rect 20352 22924 20404 22976
rect 22284 22924 22336 22976
rect 24492 22967 24544 22976
rect 24492 22933 24501 22967
rect 24501 22933 24535 22967
rect 24535 22933 24544 22967
rect 24492 22924 24544 22933
rect 3756 22822 3808 22874
rect 3820 22822 3872 22874
rect 3884 22822 3936 22874
rect 3948 22822 4000 22874
rect 4012 22822 4064 22874
rect 10472 22822 10524 22874
rect 10536 22822 10588 22874
rect 10600 22822 10652 22874
rect 10664 22822 10716 22874
rect 10728 22822 10780 22874
rect 17188 22822 17240 22874
rect 17252 22822 17304 22874
rect 17316 22822 17368 22874
rect 17380 22822 17432 22874
rect 17444 22822 17496 22874
rect 23904 22822 23956 22874
rect 23968 22822 24020 22874
rect 24032 22822 24084 22874
rect 24096 22822 24148 22874
rect 24160 22822 24212 22874
rect 2320 22720 2372 22772
rect 3332 22720 3384 22772
rect 3608 22720 3660 22772
rect 5264 22763 5316 22772
rect 5264 22729 5273 22763
rect 5273 22729 5307 22763
rect 5307 22729 5316 22763
rect 5264 22720 5316 22729
rect 9128 22720 9180 22772
rect 9772 22720 9824 22772
rect 4620 22652 4672 22704
rect 7104 22652 7156 22704
rect 5172 22584 5224 22636
rect 5356 22627 5408 22636
rect 5356 22593 5365 22627
rect 5365 22593 5399 22627
rect 5399 22593 5408 22627
rect 5356 22584 5408 22593
rect 7564 22584 7616 22636
rect 14280 22720 14332 22772
rect 16580 22763 16632 22772
rect 16580 22729 16589 22763
rect 16589 22729 16623 22763
rect 16623 22729 16632 22763
rect 16580 22720 16632 22729
rect 19616 22763 19668 22772
rect 19616 22729 19625 22763
rect 19625 22729 19659 22763
rect 19659 22729 19668 22763
rect 19616 22720 19668 22729
rect 26884 22763 26936 22772
rect 26884 22729 26893 22763
rect 26893 22729 26927 22763
rect 26927 22729 26936 22763
rect 26884 22720 26936 22729
rect 12992 22652 13044 22704
rect 14464 22652 14516 22704
rect 16396 22652 16448 22704
rect 2596 22559 2648 22568
rect 2596 22525 2605 22559
rect 2605 22525 2639 22559
rect 2639 22525 2648 22559
rect 2596 22516 2648 22525
rect 2872 22516 2924 22568
rect 4528 22559 4580 22568
rect 4528 22525 4537 22559
rect 4537 22525 4571 22559
rect 4571 22525 4580 22559
rect 4528 22516 4580 22525
rect 4988 22516 5040 22568
rect 5264 22516 5316 22568
rect 3148 22448 3200 22500
rect 5632 22516 5684 22568
rect 6368 22516 6420 22568
rect 7472 22516 7524 22568
rect 5908 22448 5960 22500
rect 7564 22448 7616 22500
rect 11336 22627 11388 22636
rect 11336 22593 11345 22627
rect 11345 22593 11379 22627
rect 11379 22593 11388 22627
rect 11336 22584 11388 22593
rect 11520 22627 11572 22636
rect 11520 22593 11529 22627
rect 11529 22593 11563 22627
rect 11563 22593 11572 22627
rect 11520 22584 11572 22593
rect 12256 22584 12308 22636
rect 12900 22584 12952 22636
rect 14924 22584 14976 22636
rect 17960 22627 18012 22636
rect 17960 22593 17969 22627
rect 17969 22593 18003 22627
rect 18003 22593 18012 22627
rect 17960 22584 18012 22593
rect 19340 22584 19392 22636
rect 20076 22584 20128 22636
rect 11888 22516 11940 22568
rect 12992 22559 13044 22568
rect 12992 22525 13001 22559
rect 13001 22525 13035 22559
rect 13035 22525 13044 22559
rect 12992 22516 13044 22525
rect 13176 22559 13228 22568
rect 13176 22525 13185 22559
rect 13185 22525 13219 22559
rect 13219 22525 13228 22559
rect 13176 22516 13228 22525
rect 13268 22516 13320 22568
rect 14740 22516 14792 22568
rect 15292 22516 15344 22568
rect 15476 22559 15528 22568
rect 15476 22525 15510 22559
rect 15510 22525 15528 22559
rect 15476 22516 15528 22525
rect 2688 22380 2740 22432
rect 4252 22380 4304 22432
rect 5724 22380 5776 22432
rect 6920 22423 6972 22432
rect 6920 22389 6929 22423
rect 6929 22389 6963 22423
rect 6963 22389 6972 22423
rect 6920 22380 6972 22389
rect 7012 22423 7064 22432
rect 7012 22389 7021 22423
rect 7021 22389 7055 22423
rect 7055 22389 7064 22423
rect 7012 22380 7064 22389
rect 8484 22380 8536 22432
rect 8760 22491 8812 22500
rect 8760 22457 8794 22491
rect 8794 22457 8812 22491
rect 8760 22448 8812 22457
rect 8852 22448 8904 22500
rect 11796 22448 11848 22500
rect 13360 22448 13412 22500
rect 17776 22559 17828 22568
rect 17776 22525 17785 22559
rect 17785 22525 17819 22559
rect 17819 22525 17828 22559
rect 17776 22516 17828 22525
rect 10140 22423 10192 22432
rect 10140 22389 10149 22423
rect 10149 22389 10183 22423
rect 10183 22389 10192 22423
rect 10140 22380 10192 22389
rect 10416 22380 10468 22432
rect 11244 22423 11296 22432
rect 11244 22389 11253 22423
rect 11253 22389 11287 22423
rect 11287 22389 11296 22423
rect 11244 22380 11296 22389
rect 12808 22380 12860 22432
rect 16948 22448 17000 22500
rect 17224 22448 17276 22500
rect 15476 22380 15528 22432
rect 22376 22559 22428 22568
rect 22376 22525 22385 22559
rect 22385 22525 22419 22559
rect 22419 22525 22428 22559
rect 22376 22516 22428 22525
rect 22560 22559 22612 22568
rect 22560 22525 22569 22559
rect 22569 22525 22603 22559
rect 22603 22525 22612 22559
rect 22560 22516 22612 22525
rect 25044 22584 25096 22636
rect 25412 22584 25464 22636
rect 22928 22559 22980 22568
rect 22928 22525 22937 22559
rect 22937 22525 22971 22559
rect 22971 22525 22980 22559
rect 22928 22516 22980 22525
rect 23204 22559 23256 22568
rect 23204 22525 23213 22559
rect 23213 22525 23247 22559
rect 23247 22525 23256 22559
rect 23204 22516 23256 22525
rect 23480 22516 23532 22568
rect 25780 22559 25832 22568
rect 25780 22525 25814 22559
rect 25814 22525 25832 22559
rect 25780 22516 25832 22525
rect 19524 22448 19576 22500
rect 20168 22448 20220 22500
rect 22468 22423 22520 22432
rect 22468 22389 22477 22423
rect 22477 22389 22511 22423
rect 22511 22389 22520 22423
rect 22468 22380 22520 22389
rect 22652 22380 22704 22432
rect 23020 22380 23072 22432
rect 23940 22380 23992 22432
rect 24860 22380 24912 22432
rect 7114 22278 7166 22330
rect 7178 22278 7230 22330
rect 7242 22278 7294 22330
rect 7306 22278 7358 22330
rect 7370 22278 7422 22330
rect 13830 22278 13882 22330
rect 13894 22278 13946 22330
rect 13958 22278 14010 22330
rect 14022 22278 14074 22330
rect 14086 22278 14138 22330
rect 20546 22278 20598 22330
rect 20610 22278 20662 22330
rect 20674 22278 20726 22330
rect 20738 22278 20790 22330
rect 20802 22278 20854 22330
rect 27262 22278 27314 22330
rect 27326 22278 27378 22330
rect 27390 22278 27442 22330
rect 27454 22278 27506 22330
rect 27518 22278 27570 22330
rect 3516 22176 3568 22228
rect 4988 22219 5040 22228
rect 4988 22185 4997 22219
rect 4997 22185 5031 22219
rect 5031 22185 5040 22219
rect 4988 22176 5040 22185
rect 5172 22176 5224 22228
rect 7472 22219 7524 22228
rect 7472 22185 7481 22219
rect 7481 22185 7515 22219
rect 7515 22185 7524 22219
rect 7472 22176 7524 22185
rect 8760 22176 8812 22228
rect 10232 22176 10284 22228
rect 13360 22219 13412 22228
rect 13360 22185 13369 22219
rect 13369 22185 13403 22219
rect 13403 22185 13412 22219
rect 13360 22176 13412 22185
rect 14464 22176 14516 22228
rect 2228 22040 2280 22092
rect 2596 22040 2648 22092
rect 4804 22040 4856 22092
rect 5080 22083 5132 22092
rect 5080 22049 5089 22083
rect 5089 22049 5123 22083
rect 5123 22049 5132 22083
rect 5080 22040 5132 22049
rect 6736 22040 6788 22092
rect 6920 22083 6972 22092
rect 6920 22049 6929 22083
rect 6929 22049 6963 22083
rect 6963 22049 6972 22083
rect 6920 22040 6972 22049
rect 8576 22083 8628 22092
rect 8576 22049 8594 22083
rect 8594 22049 8628 22083
rect 8576 22040 8628 22049
rect 9404 22083 9456 22092
rect 3148 21972 3200 22024
rect 3332 21972 3384 22024
rect 5356 22015 5408 22024
rect 5356 21981 5365 22015
rect 5365 21981 5399 22015
rect 5399 21981 5408 22015
rect 5356 21972 5408 21981
rect 6184 21972 6236 22024
rect 7656 21972 7708 22024
rect 8852 22015 8904 22024
rect 8852 21981 8861 22015
rect 8861 21981 8895 22015
rect 8895 21981 8904 22015
rect 8852 21972 8904 21981
rect 9404 22049 9413 22083
rect 9413 22049 9447 22083
rect 9447 22049 9456 22083
rect 9404 22040 9456 22049
rect 9496 22083 9548 22092
rect 9496 22049 9505 22083
rect 9505 22049 9539 22083
rect 9539 22049 9548 22083
rect 9496 22040 9548 22049
rect 10140 22151 10192 22160
rect 10140 22117 10149 22151
rect 10149 22117 10183 22151
rect 10183 22117 10192 22151
rect 10140 22108 10192 22117
rect 12348 22108 12400 22160
rect 5540 21904 5592 21956
rect 1400 21836 1452 21888
rect 5448 21836 5500 21888
rect 6460 21836 6512 21888
rect 10416 22083 10468 22092
rect 10416 22049 10425 22083
rect 10425 22049 10459 22083
rect 10459 22049 10468 22083
rect 10416 22040 10468 22049
rect 11336 22040 11388 22092
rect 11796 22083 11848 22092
rect 11796 22049 11805 22083
rect 11805 22049 11839 22083
rect 11839 22049 11848 22083
rect 11796 22040 11848 22049
rect 12256 22040 12308 22092
rect 10140 21972 10192 22024
rect 12348 21972 12400 22024
rect 14188 22108 14240 22160
rect 15292 22108 15344 22160
rect 16672 22176 16724 22228
rect 19524 22176 19576 22228
rect 22560 22176 22612 22228
rect 17040 22108 17092 22160
rect 17776 22108 17828 22160
rect 21732 22108 21784 22160
rect 13360 21972 13412 22024
rect 15200 21972 15252 22024
rect 16764 22040 16816 22092
rect 18880 22040 18932 22092
rect 20168 22040 20220 22092
rect 13452 21904 13504 21956
rect 15752 21904 15804 21956
rect 16120 21904 16172 21956
rect 17776 21947 17828 21956
rect 17776 21913 17785 21947
rect 17785 21913 17819 21947
rect 17819 21913 17828 21947
rect 17776 21904 17828 21913
rect 21456 21972 21508 22024
rect 22652 22108 22704 22160
rect 22744 22108 22796 22160
rect 23020 22151 23072 22160
rect 23020 22117 23045 22151
rect 23045 22117 23072 22151
rect 23204 22219 23256 22228
rect 23204 22185 23213 22219
rect 23213 22185 23247 22219
rect 23247 22185 23256 22219
rect 23204 22176 23256 22185
rect 23020 22108 23072 22117
rect 23296 22108 23348 22160
rect 22284 22040 22336 22092
rect 23940 22040 23992 22092
rect 22928 21972 22980 22024
rect 22100 21904 22152 21956
rect 22192 21947 22244 21956
rect 22192 21913 22201 21947
rect 22201 21913 22235 21947
rect 22235 21913 22244 21947
rect 22192 21904 22244 21913
rect 22560 21904 22612 21956
rect 25596 21972 25648 22024
rect 9404 21836 9456 21888
rect 9956 21879 10008 21888
rect 9956 21845 9965 21879
rect 9965 21845 9999 21879
rect 9999 21845 10008 21879
rect 9956 21836 10008 21845
rect 10324 21836 10376 21888
rect 11244 21836 11296 21888
rect 12256 21836 12308 21888
rect 13268 21836 13320 21888
rect 13728 21879 13780 21888
rect 13728 21845 13737 21879
rect 13737 21845 13771 21879
rect 13771 21845 13780 21879
rect 13728 21836 13780 21845
rect 16488 21836 16540 21888
rect 17224 21836 17276 21888
rect 20812 21836 20864 21888
rect 22744 21879 22796 21888
rect 22744 21845 22753 21879
rect 22753 21845 22787 21879
rect 22787 21845 22796 21879
rect 22744 21836 22796 21845
rect 3756 21734 3808 21786
rect 3820 21734 3872 21786
rect 3884 21734 3936 21786
rect 3948 21734 4000 21786
rect 4012 21734 4064 21786
rect 10472 21734 10524 21786
rect 10536 21734 10588 21786
rect 10600 21734 10652 21786
rect 10664 21734 10716 21786
rect 10728 21734 10780 21786
rect 17188 21734 17240 21786
rect 17252 21734 17304 21786
rect 17316 21734 17368 21786
rect 17380 21734 17432 21786
rect 17444 21734 17496 21786
rect 23904 21734 23956 21786
rect 23968 21734 24020 21786
rect 24032 21734 24084 21786
rect 24096 21734 24148 21786
rect 24160 21734 24212 21786
rect 1584 21632 1636 21684
rect 1952 21632 2004 21684
rect 4252 21632 4304 21684
rect 5908 21675 5960 21684
rect 5908 21641 5917 21675
rect 5917 21641 5951 21675
rect 5951 21641 5960 21675
rect 5908 21632 5960 21641
rect 7564 21632 7616 21684
rect 8668 21632 8720 21684
rect 9036 21632 9088 21684
rect 11336 21632 11388 21684
rect 13728 21632 13780 21684
rect 2044 21564 2096 21616
rect 848 21471 900 21480
rect 848 21437 857 21471
rect 857 21437 891 21471
rect 891 21437 900 21471
rect 848 21428 900 21437
rect 940 21360 992 21412
rect 2964 21360 3016 21412
rect 4160 21360 4212 21412
rect 5540 21564 5592 21616
rect 6736 21564 6788 21616
rect 8944 21564 8996 21616
rect 11520 21564 11572 21616
rect 7012 21496 7064 21548
rect 2596 21292 2648 21344
rect 2688 21335 2740 21344
rect 2688 21301 2697 21335
rect 2697 21301 2731 21335
rect 2731 21301 2740 21335
rect 2688 21292 2740 21301
rect 2872 21335 2924 21344
rect 2872 21301 2881 21335
rect 2881 21301 2915 21335
rect 2915 21301 2924 21335
rect 2872 21292 2924 21301
rect 3332 21292 3384 21344
rect 4712 21335 4764 21344
rect 4712 21301 4721 21335
rect 4721 21301 4755 21335
rect 4755 21301 4764 21335
rect 4712 21292 4764 21301
rect 4896 21335 4948 21344
rect 4896 21301 4923 21335
rect 4923 21301 4948 21335
rect 4896 21292 4948 21301
rect 5540 21292 5592 21344
rect 6092 21471 6144 21480
rect 6092 21437 6101 21471
rect 6101 21437 6135 21471
rect 6135 21437 6144 21471
rect 6092 21428 6144 21437
rect 6276 21471 6328 21480
rect 6276 21437 6285 21471
rect 6285 21437 6319 21471
rect 6319 21437 6328 21471
rect 6276 21428 6328 21437
rect 6460 21471 6512 21480
rect 6460 21437 6469 21471
rect 6469 21437 6503 21471
rect 6503 21437 6512 21471
rect 6460 21428 6512 21437
rect 6736 21428 6788 21480
rect 7840 21496 7892 21548
rect 11796 21496 11848 21548
rect 12072 21496 12124 21548
rect 7012 21360 7064 21412
rect 8944 21360 8996 21412
rect 11060 21360 11112 21412
rect 7472 21292 7524 21344
rect 8392 21335 8444 21344
rect 8392 21301 8401 21335
rect 8401 21301 8435 21335
rect 8435 21301 8444 21335
rect 8392 21292 8444 21301
rect 8576 21335 8628 21344
rect 8576 21301 8603 21335
rect 8603 21301 8628 21335
rect 8576 21292 8628 21301
rect 11244 21471 11296 21480
rect 11244 21437 11262 21471
rect 11262 21437 11296 21471
rect 11244 21428 11296 21437
rect 11428 21428 11480 21480
rect 12164 21471 12216 21480
rect 12164 21437 12173 21471
rect 12173 21437 12207 21471
rect 12207 21437 12216 21471
rect 12164 21428 12216 21437
rect 13728 21496 13780 21548
rect 11888 21360 11940 21412
rect 12348 21360 12400 21412
rect 12532 21292 12584 21344
rect 13084 21292 13136 21344
rect 14556 21564 14608 21616
rect 14372 21496 14424 21548
rect 20168 21632 20220 21684
rect 14740 21607 14792 21616
rect 14740 21573 14749 21607
rect 14749 21573 14783 21607
rect 14783 21573 14792 21607
rect 14740 21564 14792 21573
rect 16856 21564 16908 21616
rect 15200 21496 15252 21548
rect 21916 21564 21968 21616
rect 22376 21632 22428 21684
rect 22468 21632 22520 21684
rect 23480 21632 23532 21684
rect 22192 21564 22244 21616
rect 20352 21496 20404 21548
rect 22744 21607 22796 21616
rect 22744 21573 22753 21607
rect 22753 21573 22787 21607
rect 22787 21573 22796 21607
rect 22744 21564 22796 21573
rect 25596 21632 25648 21684
rect 15292 21428 15344 21480
rect 16120 21471 16172 21480
rect 16120 21437 16129 21471
rect 16129 21437 16163 21471
rect 16163 21437 16172 21471
rect 16120 21428 16172 21437
rect 16212 21428 16264 21480
rect 15108 21360 15160 21412
rect 15660 21292 15712 21344
rect 15936 21292 15988 21344
rect 16396 21292 16448 21344
rect 20168 21471 20220 21480
rect 20168 21437 20177 21471
rect 20177 21437 20211 21471
rect 20211 21437 20220 21471
rect 20168 21428 20220 21437
rect 20444 21471 20496 21480
rect 20444 21437 20453 21471
rect 20453 21437 20487 21471
rect 20487 21437 20496 21471
rect 20444 21428 20496 21437
rect 20812 21471 20864 21480
rect 20812 21437 20821 21471
rect 20821 21437 20855 21471
rect 20855 21437 20864 21471
rect 20812 21428 20864 21437
rect 21088 21471 21140 21480
rect 21088 21437 21097 21471
rect 21097 21437 21131 21471
rect 21131 21437 21140 21471
rect 21088 21428 21140 21437
rect 21272 21471 21324 21480
rect 21272 21437 21279 21471
rect 21279 21437 21324 21471
rect 21272 21428 21324 21437
rect 22008 21428 22060 21480
rect 17408 21403 17460 21412
rect 17408 21369 17442 21403
rect 17442 21369 17460 21403
rect 17408 21360 17460 21369
rect 17960 21360 18012 21412
rect 18420 21292 18472 21344
rect 18880 21292 18932 21344
rect 19800 21292 19852 21344
rect 20996 21360 21048 21412
rect 21916 21360 21968 21412
rect 22652 21360 22704 21412
rect 22376 21292 22428 21344
rect 23296 21292 23348 21344
rect 24860 21360 24912 21412
rect 25596 21403 25648 21412
rect 25596 21369 25630 21403
rect 25630 21369 25648 21403
rect 25596 21360 25648 21369
rect 26976 21292 27028 21344
rect 7114 21190 7166 21242
rect 7178 21190 7230 21242
rect 7242 21190 7294 21242
rect 7306 21190 7358 21242
rect 7370 21190 7422 21242
rect 13830 21190 13882 21242
rect 13894 21190 13946 21242
rect 13958 21190 14010 21242
rect 14022 21190 14074 21242
rect 14086 21190 14138 21242
rect 20546 21190 20598 21242
rect 20610 21190 20662 21242
rect 20674 21190 20726 21242
rect 20738 21190 20790 21242
rect 20802 21190 20854 21242
rect 27262 21190 27314 21242
rect 27326 21190 27378 21242
rect 27390 21190 27442 21242
rect 27454 21190 27506 21242
rect 27518 21190 27570 21242
rect 940 21131 992 21140
rect 940 21097 949 21131
rect 949 21097 983 21131
rect 983 21097 992 21131
rect 940 21088 992 21097
rect 1400 21131 1452 21140
rect 1400 21097 1427 21131
rect 1427 21097 1452 21131
rect 1400 21088 1452 21097
rect 1584 21063 1636 21072
rect 1584 21029 1593 21063
rect 1593 21029 1627 21063
rect 1627 21029 1636 21063
rect 1584 21020 1636 21029
rect 3240 21088 3292 21140
rect 4804 21063 4856 21072
rect 4804 21029 4813 21063
rect 4813 21029 4847 21063
rect 4847 21029 4856 21063
rect 4804 21020 4856 21029
rect 2872 20952 2924 21004
rect 3332 20952 3384 21004
rect 5264 21063 5316 21072
rect 5264 21029 5273 21063
rect 5273 21029 5307 21063
rect 5307 21029 5316 21063
rect 5264 21020 5316 21029
rect 6736 21020 6788 21072
rect 9772 21088 9824 21140
rect 15292 21088 15344 21140
rect 15752 21088 15804 21140
rect 8484 21063 8536 21072
rect 8484 21029 8493 21063
rect 8493 21029 8527 21063
rect 8527 21029 8536 21063
rect 8484 21020 8536 21029
rect 848 20884 900 20936
rect 2780 20884 2832 20936
rect 4160 20927 4212 20936
rect 4160 20893 4169 20927
rect 4169 20893 4203 20927
rect 4203 20893 4212 20927
rect 4160 20884 4212 20893
rect 4344 20927 4396 20936
rect 4344 20893 4353 20927
rect 4353 20893 4387 20927
rect 4387 20893 4396 20927
rect 4344 20884 4396 20893
rect 4436 20927 4488 20936
rect 4436 20893 4445 20927
rect 4445 20893 4479 20927
rect 4479 20893 4488 20927
rect 4436 20884 4488 20893
rect 4528 20927 4580 20936
rect 4528 20893 4537 20927
rect 4537 20893 4571 20927
rect 4571 20893 4580 20927
rect 4528 20884 4580 20893
rect 2964 20816 3016 20868
rect 4896 20859 4948 20868
rect 4896 20825 4905 20859
rect 4905 20825 4939 20859
rect 4939 20825 4948 20859
rect 4896 20816 4948 20825
rect 5448 20995 5500 21004
rect 5448 20961 5457 20995
rect 5457 20961 5491 20995
rect 5491 20961 5500 20995
rect 5448 20952 5500 20961
rect 6184 20952 6236 21004
rect 6828 20952 6880 21004
rect 8116 20995 8168 21004
rect 8116 20961 8134 20995
rect 8134 20961 8168 20995
rect 8116 20952 8168 20961
rect 8576 20952 8628 21004
rect 9864 21020 9916 21072
rect 11888 21063 11940 21072
rect 8760 20952 8812 21004
rect 9680 20995 9732 21004
rect 9680 20961 9689 20995
rect 9689 20961 9723 20995
rect 9723 20961 9732 20995
rect 9680 20952 9732 20961
rect 5724 20884 5776 20936
rect 8852 20884 8904 20936
rect 9588 20884 9640 20936
rect 10140 20927 10192 20936
rect 10140 20893 10149 20927
rect 10149 20893 10183 20927
rect 10183 20893 10192 20927
rect 10140 20884 10192 20893
rect 11428 20995 11480 21004
rect 11428 20961 11437 20995
rect 11437 20961 11471 20995
rect 11471 20961 11480 20995
rect 11428 20952 11480 20961
rect 7012 20859 7064 20868
rect 2412 20748 2464 20800
rect 7012 20825 7021 20859
rect 7021 20825 7055 20859
rect 7055 20825 7064 20859
rect 7012 20816 7064 20825
rect 5356 20748 5408 20800
rect 9680 20816 9732 20868
rect 11336 20884 11388 20936
rect 11888 21029 11897 21063
rect 11897 21029 11931 21063
rect 11931 21029 11940 21063
rect 11888 21020 11940 21029
rect 12164 21020 12216 21072
rect 11704 20927 11756 20936
rect 11704 20893 11713 20927
rect 11713 20893 11747 20927
rect 11747 20893 11756 20927
rect 11704 20884 11756 20893
rect 12992 20995 13044 21004
rect 12992 20961 13001 20995
rect 13001 20961 13035 20995
rect 13035 20961 13044 20995
rect 12992 20952 13044 20961
rect 13084 20995 13136 21004
rect 13084 20961 13093 20995
rect 13093 20961 13127 20995
rect 13127 20961 13136 20995
rect 13084 20952 13136 20961
rect 13360 20995 13412 21004
rect 13360 20961 13369 20995
rect 13369 20961 13403 20995
rect 13403 20961 13412 20995
rect 13360 20952 13412 20961
rect 13636 20995 13688 21004
rect 13636 20961 13670 20995
rect 13670 20961 13688 20995
rect 13636 20952 13688 20961
rect 15292 20952 15344 21004
rect 15384 20995 15436 21004
rect 15384 20961 15393 20995
rect 15393 20961 15427 20995
rect 15427 20961 15436 20995
rect 15384 20952 15436 20961
rect 15476 20995 15528 21004
rect 15476 20961 15485 20995
rect 15485 20961 15519 20995
rect 15519 20961 15528 20995
rect 15476 20952 15528 20961
rect 16212 20995 16264 21004
rect 16212 20961 16221 20995
rect 16221 20961 16255 20995
rect 16255 20961 16264 20995
rect 16212 20952 16264 20961
rect 17408 21131 17460 21140
rect 17408 21097 17417 21131
rect 17417 21097 17451 21131
rect 17451 21097 17460 21131
rect 17408 21088 17460 21097
rect 8668 20791 8720 20800
rect 8668 20757 8677 20791
rect 8677 20757 8711 20791
rect 8711 20757 8720 20791
rect 8668 20748 8720 20757
rect 8852 20791 8904 20800
rect 8852 20757 8861 20791
rect 8861 20757 8895 20791
rect 8895 20757 8904 20791
rect 8852 20748 8904 20757
rect 10232 20748 10284 20800
rect 12072 20791 12124 20800
rect 12072 20757 12081 20791
rect 12081 20757 12115 20791
rect 12115 20757 12124 20791
rect 12072 20748 12124 20757
rect 15016 20927 15068 20936
rect 15016 20893 15025 20927
rect 15025 20893 15059 20927
rect 15059 20893 15068 20927
rect 15016 20884 15068 20893
rect 15660 20884 15712 20936
rect 17040 20952 17092 21004
rect 17684 20995 17736 21004
rect 17684 20961 17693 20995
rect 17693 20961 17727 20995
rect 17727 20961 17736 20995
rect 17684 20952 17736 20961
rect 17776 20995 17828 21004
rect 17776 20961 17785 20995
rect 17785 20961 17819 20995
rect 17819 20961 17828 20995
rect 17776 20952 17828 20961
rect 17960 20995 18012 21004
rect 17960 20961 17969 20995
rect 17969 20961 18003 20995
rect 18003 20961 18012 20995
rect 17960 20952 18012 20961
rect 18880 21020 18932 21072
rect 20168 21088 20220 21140
rect 20996 21131 21048 21140
rect 20996 21097 21005 21131
rect 21005 21097 21039 21131
rect 21039 21097 21048 21131
rect 20996 21088 21048 21097
rect 21088 21088 21140 21140
rect 21364 21088 21416 21140
rect 25596 21131 25648 21140
rect 25596 21097 25605 21131
rect 25605 21097 25639 21131
rect 25639 21097 25648 21131
rect 25596 21088 25648 21097
rect 22008 21020 22060 21072
rect 22284 21020 22336 21072
rect 23296 21063 23348 21072
rect 23296 21029 23305 21063
rect 23305 21029 23339 21063
rect 23339 21029 23348 21063
rect 23296 21020 23348 21029
rect 23480 21063 23532 21072
rect 23480 21029 23505 21063
rect 23505 21029 23532 21063
rect 23480 21020 23532 21029
rect 17868 20884 17920 20936
rect 17776 20816 17828 20868
rect 18696 20995 18748 21004
rect 18696 20961 18705 20995
rect 18705 20961 18739 20995
rect 18739 20961 18748 20995
rect 18696 20952 18748 20961
rect 20444 20952 20496 21004
rect 23204 20952 23256 21004
rect 18972 20884 19024 20936
rect 22652 20884 22704 20936
rect 25044 20884 25096 20936
rect 12440 20791 12492 20800
rect 12440 20757 12449 20791
rect 12449 20757 12483 20791
rect 12483 20757 12492 20791
rect 12440 20748 12492 20757
rect 13544 20748 13596 20800
rect 13728 20748 13780 20800
rect 15752 20748 15804 20800
rect 16304 20791 16356 20800
rect 16304 20757 16313 20791
rect 16313 20757 16347 20791
rect 16347 20757 16356 20791
rect 16304 20748 16356 20757
rect 20352 20816 20404 20868
rect 19800 20748 19852 20800
rect 21456 20816 21508 20868
rect 23296 20816 23348 20868
rect 22468 20791 22520 20800
rect 22468 20757 22477 20791
rect 22477 20757 22511 20791
rect 22511 20757 22520 20791
rect 22468 20748 22520 20757
rect 23572 20748 23624 20800
rect 23756 20748 23808 20800
rect 26976 20995 27028 21004
rect 26976 20961 26985 20995
rect 26985 20961 27019 20995
rect 27019 20961 27028 20995
rect 26976 20952 27028 20961
rect 3756 20646 3808 20698
rect 3820 20646 3872 20698
rect 3884 20646 3936 20698
rect 3948 20646 4000 20698
rect 4012 20646 4064 20698
rect 10472 20646 10524 20698
rect 10536 20646 10588 20698
rect 10600 20646 10652 20698
rect 10664 20646 10716 20698
rect 10728 20646 10780 20698
rect 17188 20646 17240 20698
rect 17252 20646 17304 20698
rect 17316 20646 17368 20698
rect 17380 20646 17432 20698
rect 17444 20646 17496 20698
rect 23904 20646 23956 20698
rect 23968 20646 24020 20698
rect 24032 20646 24084 20698
rect 24096 20646 24148 20698
rect 24160 20646 24212 20698
rect 2320 20544 2372 20596
rect 2688 20544 2740 20596
rect 2044 20408 2096 20460
rect 2228 20340 2280 20392
rect 2412 20383 2464 20392
rect 2412 20349 2421 20383
rect 2421 20349 2455 20383
rect 2455 20349 2464 20383
rect 2412 20340 2464 20349
rect 1584 20272 1636 20324
rect 2688 20383 2740 20392
rect 2688 20349 2697 20383
rect 2697 20349 2731 20383
rect 2731 20349 2740 20383
rect 2688 20340 2740 20349
rect 2780 20272 2832 20324
rect 1216 20204 1268 20256
rect 1860 20247 1912 20256
rect 1860 20213 1887 20247
rect 1887 20213 1912 20247
rect 1860 20204 1912 20213
rect 2504 20204 2556 20256
rect 3332 20340 3384 20392
rect 3792 20204 3844 20256
rect 4528 20544 4580 20596
rect 5264 20544 5316 20596
rect 6736 20544 6788 20596
rect 8116 20544 8168 20596
rect 8484 20544 8536 20596
rect 11336 20587 11388 20596
rect 11336 20553 11345 20587
rect 11345 20553 11379 20587
rect 11379 20553 11388 20587
rect 11336 20544 11388 20553
rect 13636 20544 13688 20596
rect 15384 20544 15436 20596
rect 15752 20544 15804 20596
rect 4344 20476 4396 20528
rect 15844 20476 15896 20528
rect 19892 20544 19944 20596
rect 17776 20476 17828 20528
rect 4160 20408 4212 20460
rect 4252 20340 4304 20392
rect 5448 20408 5500 20460
rect 13360 20408 13412 20460
rect 17960 20408 18012 20460
rect 18696 20408 18748 20460
rect 22100 20544 22152 20596
rect 23480 20544 23532 20596
rect 20076 20408 20128 20460
rect 4896 20383 4948 20392
rect 4896 20349 4905 20383
rect 4905 20349 4939 20383
rect 4939 20349 4948 20383
rect 4896 20340 4948 20349
rect 5724 20340 5776 20392
rect 7472 20383 7524 20392
rect 7472 20349 7481 20383
rect 7481 20349 7515 20383
rect 7515 20349 7524 20383
rect 7472 20340 7524 20349
rect 8392 20340 8444 20392
rect 9680 20340 9732 20392
rect 10232 20383 10284 20392
rect 10232 20349 10266 20383
rect 10266 20349 10284 20383
rect 10232 20340 10284 20349
rect 13544 20383 13596 20392
rect 13544 20349 13553 20383
rect 13553 20349 13587 20383
rect 13587 20349 13596 20383
rect 13544 20340 13596 20349
rect 14832 20340 14884 20392
rect 16304 20340 16356 20392
rect 5540 20272 5592 20324
rect 8484 20272 8536 20324
rect 9036 20272 9088 20324
rect 7932 20204 7984 20256
rect 12624 20204 12676 20256
rect 17868 20383 17920 20392
rect 17868 20349 17877 20383
rect 17877 20349 17911 20383
rect 17911 20349 17920 20383
rect 17868 20340 17920 20349
rect 18328 20272 18380 20324
rect 19248 20272 19300 20324
rect 19708 20383 19760 20392
rect 19708 20349 19717 20383
rect 19717 20349 19751 20383
rect 19751 20349 19760 20383
rect 19708 20340 19760 20349
rect 20168 20340 20220 20392
rect 21088 20340 21140 20392
rect 15292 20204 15344 20256
rect 18052 20204 18104 20256
rect 19432 20247 19484 20256
rect 19432 20213 19441 20247
rect 19441 20213 19475 20247
rect 19475 20213 19484 20247
rect 19432 20204 19484 20213
rect 19800 20315 19852 20324
rect 19800 20281 19809 20315
rect 19809 20281 19843 20315
rect 19843 20281 19852 20315
rect 19800 20272 19852 20281
rect 20444 20272 20496 20324
rect 21456 20340 21508 20392
rect 21732 20451 21784 20460
rect 21732 20417 21741 20451
rect 21741 20417 21775 20451
rect 21775 20417 21784 20451
rect 21732 20408 21784 20417
rect 21640 20383 21692 20392
rect 21640 20349 21649 20383
rect 21649 20349 21683 20383
rect 21683 20349 21692 20383
rect 22468 20408 22520 20460
rect 21640 20340 21692 20349
rect 21916 20383 21968 20392
rect 21916 20349 21925 20383
rect 21925 20349 21959 20383
rect 21959 20349 21968 20383
rect 21916 20340 21968 20349
rect 22008 20383 22060 20392
rect 22008 20349 22017 20383
rect 22017 20349 22051 20383
rect 22051 20349 22060 20383
rect 22008 20340 22060 20349
rect 22376 20383 22428 20392
rect 22376 20349 22385 20383
rect 22385 20349 22419 20383
rect 22419 20349 22428 20383
rect 22376 20340 22428 20349
rect 22560 20383 22612 20392
rect 22560 20349 22569 20383
rect 22569 20349 22603 20383
rect 22603 20349 22612 20383
rect 22560 20340 22612 20349
rect 22744 20340 22796 20392
rect 21272 20315 21324 20324
rect 21272 20281 21281 20315
rect 21281 20281 21315 20315
rect 21315 20281 21324 20315
rect 21272 20272 21324 20281
rect 22836 20272 22888 20324
rect 23204 20315 23256 20324
rect 23204 20281 23213 20315
rect 23213 20281 23247 20315
rect 23247 20281 23256 20315
rect 23756 20340 23808 20392
rect 23204 20272 23256 20281
rect 20996 20247 21048 20256
rect 20996 20213 21005 20247
rect 21005 20213 21039 20247
rect 21039 20213 21048 20247
rect 20996 20204 21048 20213
rect 21088 20204 21140 20256
rect 21548 20204 21600 20256
rect 22744 20247 22796 20256
rect 22744 20213 22753 20247
rect 22753 20213 22787 20247
rect 22787 20213 22796 20247
rect 22744 20204 22796 20213
rect 23572 20247 23624 20256
rect 23572 20213 23581 20247
rect 23581 20213 23615 20247
rect 23615 20213 23624 20247
rect 23572 20204 23624 20213
rect 25872 20340 25924 20392
rect 27068 20272 27120 20324
rect 7114 20102 7166 20154
rect 7178 20102 7230 20154
rect 7242 20102 7294 20154
rect 7306 20102 7358 20154
rect 7370 20102 7422 20154
rect 13830 20102 13882 20154
rect 13894 20102 13946 20154
rect 13958 20102 14010 20154
rect 14022 20102 14074 20154
rect 14086 20102 14138 20154
rect 20546 20102 20598 20154
rect 20610 20102 20662 20154
rect 20674 20102 20726 20154
rect 20738 20102 20790 20154
rect 20802 20102 20854 20154
rect 27262 20102 27314 20154
rect 27326 20102 27378 20154
rect 27390 20102 27442 20154
rect 27454 20102 27506 20154
rect 27518 20102 27570 20154
rect 2228 20043 2280 20052
rect 2228 20009 2237 20043
rect 2237 20009 2271 20043
rect 2271 20009 2280 20043
rect 2228 20000 2280 20009
rect 2320 20043 2372 20052
rect 2320 20009 2329 20043
rect 2329 20009 2363 20043
rect 2363 20009 2372 20043
rect 2320 20000 2372 20009
rect 4436 20000 4488 20052
rect 9036 20043 9088 20052
rect 9036 20009 9045 20043
rect 9045 20009 9079 20043
rect 9079 20009 9088 20043
rect 9036 20000 9088 20009
rect 3700 19932 3752 19984
rect 1124 19907 1176 19916
rect 1124 19873 1158 19907
rect 1158 19873 1176 19907
rect 1124 19864 1176 19873
rect 2044 19864 2096 19916
rect 2688 19907 2740 19916
rect 2688 19873 2697 19907
rect 2697 19873 2731 19907
rect 2731 19873 2740 19907
rect 2688 19864 2740 19873
rect 2780 19907 2832 19916
rect 2780 19873 2789 19907
rect 2789 19873 2823 19907
rect 2823 19873 2832 19907
rect 2780 19864 2832 19873
rect 3332 19907 3384 19916
rect 3332 19873 3341 19907
rect 3341 19873 3375 19907
rect 3375 19873 3384 19907
rect 3332 19864 3384 19873
rect 3792 19907 3844 19916
rect 3792 19873 3801 19907
rect 3801 19873 3835 19907
rect 3835 19873 3844 19907
rect 3792 19864 3844 19873
rect 10968 20000 11020 20052
rect 12532 20000 12584 20052
rect 14832 20043 14884 20052
rect 14832 20009 14841 20043
rect 14841 20009 14875 20043
rect 14875 20009 14884 20043
rect 14832 20000 14884 20009
rect 15384 20000 15436 20052
rect 15660 20000 15712 20052
rect 848 19839 900 19848
rect 848 19805 857 19839
rect 857 19805 891 19839
rect 891 19805 900 19839
rect 848 19796 900 19805
rect 4252 19728 4304 19780
rect 4712 19907 4764 19916
rect 4712 19873 4721 19907
rect 4721 19873 4755 19907
rect 4755 19873 4764 19907
rect 4712 19864 4764 19873
rect 5080 19864 5132 19916
rect 6736 19864 6788 19916
rect 7472 19864 7524 19916
rect 4436 19796 4488 19848
rect 4896 19839 4948 19848
rect 4896 19805 4905 19839
rect 4905 19805 4939 19839
rect 4939 19805 4948 19839
rect 4896 19796 4948 19805
rect 5724 19796 5776 19848
rect 8852 19907 8904 19916
rect 8852 19873 8861 19907
rect 8861 19873 8895 19907
rect 8895 19873 8904 19907
rect 8852 19864 8904 19873
rect 9864 19864 9916 19916
rect 11428 19864 11480 19916
rect 12440 19932 12492 19984
rect 12808 19932 12860 19984
rect 15292 19932 15344 19984
rect 18696 20043 18748 20052
rect 18696 20009 18705 20043
rect 18705 20009 18739 20043
rect 18739 20009 18748 20043
rect 18696 20000 18748 20009
rect 19800 20000 19852 20052
rect 21088 20000 21140 20052
rect 12348 19864 12400 19916
rect 10048 19796 10100 19848
rect 10876 19796 10928 19848
rect 2964 19703 3016 19712
rect 2964 19669 2973 19703
rect 2973 19669 3007 19703
rect 3007 19669 3016 19703
rect 2964 19660 3016 19669
rect 5632 19660 5684 19712
rect 12716 19796 12768 19848
rect 12900 19796 12952 19848
rect 13636 19796 13688 19848
rect 12072 19771 12124 19780
rect 12072 19737 12081 19771
rect 12081 19737 12115 19771
rect 12115 19737 12124 19771
rect 12072 19728 12124 19737
rect 15660 19864 15712 19916
rect 15752 19864 15804 19916
rect 17960 19932 18012 19984
rect 17592 19907 17644 19916
rect 17592 19873 17626 19907
rect 17626 19873 17644 19907
rect 17592 19864 17644 19873
rect 20996 19932 21048 19984
rect 21640 20000 21692 20052
rect 22560 20000 22612 20052
rect 14648 19839 14700 19848
rect 14648 19805 14657 19839
rect 14657 19805 14691 19839
rect 14691 19805 14700 19839
rect 14648 19796 14700 19805
rect 16488 19796 16540 19848
rect 18972 19796 19024 19848
rect 21732 19932 21784 19984
rect 22100 19864 22152 19916
rect 22376 19932 22428 19984
rect 22652 19932 22704 19984
rect 23204 20000 23256 20052
rect 23388 19975 23440 19984
rect 23388 19941 23397 19975
rect 23397 19941 23431 19975
rect 23431 19941 23440 19975
rect 23388 19932 23440 19941
rect 23572 19796 23624 19848
rect 8392 19703 8444 19712
rect 8392 19669 8401 19703
rect 8401 19669 8435 19703
rect 8435 19669 8444 19703
rect 8392 19660 8444 19669
rect 11704 19703 11756 19712
rect 11704 19669 11713 19703
rect 11713 19669 11747 19703
rect 11747 19669 11756 19703
rect 11704 19660 11756 19669
rect 12440 19660 12492 19712
rect 13176 19660 13228 19712
rect 13820 19703 13872 19712
rect 13820 19669 13829 19703
rect 13829 19669 13863 19703
rect 13863 19669 13872 19703
rect 13820 19660 13872 19669
rect 14096 19660 14148 19712
rect 15016 19703 15068 19712
rect 15016 19669 15025 19703
rect 15025 19669 15059 19703
rect 15059 19669 15068 19703
rect 15016 19660 15068 19669
rect 15752 19703 15804 19712
rect 15752 19669 15761 19703
rect 15761 19669 15795 19703
rect 15795 19669 15804 19703
rect 15752 19660 15804 19669
rect 15844 19660 15896 19712
rect 16856 19703 16908 19712
rect 16856 19669 16865 19703
rect 16865 19669 16899 19703
rect 16899 19669 16908 19703
rect 16856 19660 16908 19669
rect 22652 19660 22704 19712
rect 22836 19660 22888 19712
rect 23020 19771 23072 19780
rect 23020 19737 23029 19771
rect 23029 19737 23063 19771
rect 23063 19737 23072 19771
rect 23020 19728 23072 19737
rect 23204 19728 23256 19780
rect 27068 19796 27120 19848
rect 3756 19558 3808 19610
rect 3820 19558 3872 19610
rect 3884 19558 3936 19610
rect 3948 19558 4000 19610
rect 4012 19558 4064 19610
rect 10472 19558 10524 19610
rect 10536 19558 10588 19610
rect 10600 19558 10652 19610
rect 10664 19558 10716 19610
rect 10728 19558 10780 19610
rect 17188 19558 17240 19610
rect 17252 19558 17304 19610
rect 17316 19558 17368 19610
rect 17380 19558 17432 19610
rect 17444 19558 17496 19610
rect 23904 19558 23956 19610
rect 23968 19558 24020 19610
rect 24032 19558 24084 19610
rect 24096 19558 24148 19610
rect 24160 19558 24212 19610
rect 1124 19456 1176 19508
rect 1492 19456 1544 19508
rect 2780 19456 2832 19508
rect 3332 19456 3384 19508
rect 4252 19499 4304 19508
rect 4252 19465 4261 19499
rect 4261 19465 4295 19499
rect 4295 19465 4304 19499
rect 4252 19456 4304 19465
rect 4436 19499 4488 19508
rect 4436 19465 4445 19499
rect 4445 19465 4479 19499
rect 4479 19465 4488 19499
rect 4436 19456 4488 19465
rect 6736 19499 6788 19508
rect 6736 19465 6745 19499
rect 6745 19465 6779 19499
rect 6779 19465 6788 19499
rect 6736 19456 6788 19465
rect 8116 19456 8168 19508
rect 12900 19499 12952 19508
rect 12900 19465 12909 19499
rect 12909 19465 12943 19499
rect 12943 19465 12952 19499
rect 12900 19456 12952 19465
rect 13176 19499 13228 19508
rect 13176 19465 13185 19499
rect 13185 19465 13219 19499
rect 13219 19465 13228 19499
rect 13176 19456 13228 19465
rect 13820 19456 13872 19508
rect 16212 19499 16264 19508
rect 16212 19465 16221 19499
rect 16221 19465 16255 19499
rect 16255 19465 16264 19499
rect 16212 19456 16264 19465
rect 17592 19456 17644 19508
rect 20168 19456 20220 19508
rect 22652 19456 22704 19508
rect 23020 19456 23072 19508
rect 2044 19431 2096 19440
rect 2044 19397 2053 19431
rect 2053 19397 2087 19431
rect 2087 19397 2096 19431
rect 2044 19388 2096 19397
rect 1216 19295 1268 19304
rect 1216 19261 1225 19295
rect 1225 19261 1259 19295
rect 1259 19261 1268 19295
rect 1216 19252 1268 19261
rect 1860 19252 1912 19304
rect 3608 19320 3660 19372
rect 5632 19363 5684 19372
rect 5632 19329 5641 19363
rect 5641 19329 5675 19363
rect 5675 19329 5684 19363
rect 5632 19320 5684 19329
rect 2504 19184 2556 19236
rect 4620 19252 4672 19304
rect 5816 19388 5868 19440
rect 5816 19295 5868 19304
rect 5816 19261 5825 19295
rect 5825 19261 5859 19295
rect 5859 19261 5868 19295
rect 5816 19252 5868 19261
rect 14648 19388 14700 19440
rect 17316 19388 17368 19440
rect 17776 19388 17828 19440
rect 22100 19388 22152 19440
rect 5632 19184 5684 19236
rect 7196 19295 7248 19304
rect 7196 19261 7205 19295
rect 7205 19261 7239 19295
rect 7239 19261 7248 19295
rect 7196 19252 7248 19261
rect 7748 19252 7800 19304
rect 11520 19295 11572 19304
rect 11520 19261 11529 19295
rect 11529 19261 11563 19295
rect 11563 19261 11572 19295
rect 11520 19252 11572 19261
rect 13360 19252 13412 19304
rect 2688 19116 2740 19168
rect 4620 19116 4672 19168
rect 5908 19116 5960 19168
rect 6460 19116 6512 19168
rect 7472 19159 7524 19168
rect 7472 19125 7497 19159
rect 7497 19125 7524 19159
rect 7472 19116 7524 19125
rect 7656 19159 7708 19168
rect 7656 19125 7665 19159
rect 7665 19125 7699 19159
rect 7699 19125 7708 19159
rect 7656 19116 7708 19125
rect 8392 19184 8444 19236
rect 8576 19227 8628 19236
rect 8576 19193 8585 19227
rect 8585 19193 8619 19227
rect 8619 19193 8628 19227
rect 8576 19184 8628 19193
rect 9496 19227 9548 19236
rect 9496 19193 9505 19227
rect 9505 19193 9539 19227
rect 9539 19193 9548 19227
rect 9496 19184 9548 19193
rect 9772 19184 9824 19236
rect 11060 19227 11112 19236
rect 11060 19193 11069 19227
rect 11069 19193 11103 19227
rect 11103 19193 11112 19227
rect 11060 19184 11112 19193
rect 12256 19184 12308 19236
rect 14096 19252 14148 19304
rect 15200 19295 15252 19304
rect 15200 19261 15209 19295
rect 15209 19261 15243 19295
rect 15243 19261 15252 19295
rect 15200 19252 15252 19261
rect 15292 19295 15344 19304
rect 15292 19261 15301 19295
rect 15301 19261 15335 19295
rect 15335 19261 15344 19295
rect 15292 19252 15344 19261
rect 15752 19252 15804 19304
rect 15844 19295 15896 19304
rect 15844 19261 15853 19295
rect 15853 19261 15887 19295
rect 15887 19261 15896 19295
rect 15844 19252 15896 19261
rect 16120 19252 16172 19304
rect 8760 19159 8812 19168
rect 8760 19125 8785 19159
rect 8785 19125 8812 19159
rect 8760 19116 8812 19125
rect 8944 19159 8996 19168
rect 8944 19125 8953 19159
rect 8953 19125 8987 19159
rect 8987 19125 8996 19159
rect 8944 19116 8996 19125
rect 12808 19116 12860 19168
rect 13360 19159 13412 19168
rect 13360 19125 13369 19159
rect 13369 19125 13403 19159
rect 13403 19125 13412 19159
rect 13360 19116 13412 19125
rect 13544 19116 13596 19168
rect 15476 19184 15528 19236
rect 16856 19252 16908 19304
rect 17868 19320 17920 19372
rect 17316 19295 17368 19304
rect 17316 19261 17325 19295
rect 17325 19261 17359 19295
rect 17359 19261 17368 19295
rect 17316 19252 17368 19261
rect 18052 19252 18104 19304
rect 18972 19252 19024 19304
rect 21180 19295 21232 19304
rect 21180 19261 21189 19295
rect 21189 19261 21223 19295
rect 21223 19261 21232 19295
rect 21180 19252 21232 19261
rect 22284 19320 22336 19372
rect 17224 19227 17276 19236
rect 17224 19193 17233 19227
rect 17233 19193 17267 19227
rect 17267 19193 17276 19227
rect 17224 19184 17276 19193
rect 17592 19227 17644 19236
rect 17592 19193 17601 19227
rect 17601 19193 17635 19227
rect 17635 19193 17644 19227
rect 17592 19184 17644 19193
rect 18512 19184 18564 19236
rect 19064 19184 19116 19236
rect 21088 19184 21140 19236
rect 15016 19159 15068 19168
rect 15016 19125 15025 19159
rect 15025 19125 15059 19159
rect 15059 19125 15068 19159
rect 15016 19116 15068 19125
rect 15752 19116 15804 19168
rect 20444 19116 20496 19168
rect 21824 19116 21876 19168
rect 22376 19295 22428 19304
rect 22376 19261 22385 19295
rect 22385 19261 22419 19295
rect 22419 19261 22428 19295
rect 22376 19252 22428 19261
rect 22836 19320 22888 19372
rect 22744 19295 22796 19304
rect 22744 19261 22753 19295
rect 22753 19261 22787 19295
rect 22787 19261 22796 19295
rect 22744 19252 22796 19261
rect 23020 19295 23072 19304
rect 23020 19261 23029 19295
rect 23029 19261 23063 19295
rect 23063 19261 23072 19295
rect 23020 19252 23072 19261
rect 23296 19252 23348 19304
rect 25136 19252 25188 19304
rect 27068 19252 27120 19304
rect 22928 19184 22980 19236
rect 23388 19227 23440 19236
rect 23388 19193 23397 19227
rect 23397 19193 23431 19227
rect 23431 19193 23440 19227
rect 23388 19184 23440 19193
rect 25780 19184 25832 19236
rect 22468 19116 22520 19168
rect 23296 19116 23348 19168
rect 24768 19116 24820 19168
rect 7114 19014 7166 19066
rect 7178 19014 7230 19066
rect 7242 19014 7294 19066
rect 7306 19014 7358 19066
rect 7370 19014 7422 19066
rect 13830 19014 13882 19066
rect 13894 19014 13946 19066
rect 13958 19014 14010 19066
rect 14022 19014 14074 19066
rect 14086 19014 14138 19066
rect 20546 19014 20598 19066
rect 20610 19014 20662 19066
rect 20674 19014 20726 19066
rect 20738 19014 20790 19066
rect 20802 19014 20854 19066
rect 27262 19014 27314 19066
rect 27326 19014 27378 19066
rect 27390 19014 27442 19066
rect 27454 19014 27506 19066
rect 27518 19014 27570 19066
rect 2504 18955 2556 18964
rect 2504 18921 2513 18955
rect 2513 18921 2547 18955
rect 2547 18921 2556 18955
rect 2504 18912 2556 18921
rect 5816 18912 5868 18964
rect 6368 18912 6420 18964
rect 8576 18912 8628 18964
rect 11060 18912 11112 18964
rect 2964 18844 3016 18896
rect 5724 18776 5776 18828
rect 6552 18844 6604 18896
rect 6000 18819 6052 18828
rect 6000 18785 6009 18819
rect 6009 18785 6043 18819
rect 6043 18785 6052 18819
rect 6000 18776 6052 18785
rect 6092 18819 6144 18828
rect 6092 18785 6101 18819
rect 6101 18785 6135 18819
rect 6135 18785 6144 18819
rect 6092 18776 6144 18785
rect 7288 18776 7340 18828
rect 8576 18776 8628 18828
rect 11520 18844 11572 18896
rect 12256 18887 12308 18896
rect 12256 18853 12265 18887
rect 12265 18853 12299 18887
rect 12299 18853 12308 18887
rect 12256 18844 12308 18853
rect 13452 18844 13504 18896
rect 13544 18887 13596 18896
rect 13544 18853 13553 18887
rect 13553 18853 13587 18887
rect 13587 18853 13596 18887
rect 13544 18844 13596 18853
rect 15200 18844 15252 18896
rect 20444 18912 20496 18964
rect 21272 18912 21324 18964
rect 21364 18912 21416 18964
rect 23020 18912 23072 18964
rect 25780 18955 25832 18964
rect 25780 18921 25789 18955
rect 25789 18921 25823 18955
rect 25823 18921 25832 18955
rect 25780 18912 25832 18921
rect 4988 18572 5040 18624
rect 9588 18708 9640 18760
rect 6460 18683 6512 18692
rect 6460 18649 6469 18683
rect 6469 18649 6503 18683
rect 6503 18649 6512 18683
rect 6460 18640 6512 18649
rect 11060 18751 11112 18760
rect 11060 18717 11069 18751
rect 11069 18717 11103 18751
rect 11103 18717 11112 18751
rect 11060 18708 11112 18717
rect 11428 18819 11480 18828
rect 11428 18785 11437 18819
rect 11437 18785 11471 18819
rect 11471 18785 11480 18819
rect 11428 18776 11480 18785
rect 11704 18819 11756 18828
rect 11704 18785 11713 18819
rect 11713 18785 11747 18819
rect 11747 18785 11756 18819
rect 11704 18776 11756 18785
rect 12440 18819 12492 18828
rect 12440 18785 12449 18819
rect 12449 18785 12483 18819
rect 12483 18785 12492 18819
rect 12440 18776 12492 18785
rect 12624 18819 12676 18828
rect 12624 18785 12633 18819
rect 12633 18785 12667 18819
rect 12667 18785 12676 18819
rect 12624 18776 12676 18785
rect 13084 18819 13136 18828
rect 13084 18785 13093 18819
rect 13093 18785 13127 18819
rect 13127 18785 13136 18819
rect 13084 18776 13136 18785
rect 13360 18819 13412 18828
rect 13360 18785 13369 18819
rect 13369 18785 13403 18819
rect 13403 18785 13412 18819
rect 13360 18776 13412 18785
rect 13636 18819 13688 18828
rect 13636 18785 13645 18819
rect 13645 18785 13679 18819
rect 13679 18785 13688 18819
rect 13636 18776 13688 18785
rect 14372 18776 14424 18828
rect 16672 18776 16724 18828
rect 17684 18776 17736 18828
rect 11612 18640 11664 18692
rect 15936 18640 15988 18692
rect 8392 18572 8444 18624
rect 11060 18572 11112 18624
rect 16120 18683 16172 18692
rect 16120 18649 16129 18683
rect 16129 18649 16163 18683
rect 16163 18649 16172 18683
rect 16120 18640 16172 18649
rect 17500 18572 17552 18624
rect 21732 18844 21784 18896
rect 19064 18776 19116 18828
rect 21364 18776 21416 18828
rect 21456 18819 21508 18828
rect 21456 18785 21465 18819
rect 21465 18785 21499 18819
rect 21499 18785 21508 18819
rect 21456 18776 21508 18785
rect 21640 18819 21692 18828
rect 21640 18785 21649 18819
rect 21649 18785 21683 18819
rect 21683 18785 21692 18819
rect 21640 18776 21692 18785
rect 21824 18819 21876 18828
rect 21824 18785 21833 18819
rect 21833 18785 21867 18819
rect 21867 18785 21876 18819
rect 21824 18776 21876 18785
rect 22284 18887 22336 18896
rect 22284 18853 22293 18887
rect 22293 18853 22327 18887
rect 22327 18853 22336 18887
rect 22284 18844 22336 18853
rect 20904 18708 20956 18760
rect 22468 18819 22520 18828
rect 22468 18785 22477 18819
rect 22477 18785 22511 18819
rect 22511 18785 22520 18819
rect 22468 18776 22520 18785
rect 22560 18751 22612 18760
rect 22560 18717 22569 18751
rect 22569 18717 22603 18751
rect 22603 18717 22612 18751
rect 22560 18708 22612 18717
rect 22744 18819 22796 18828
rect 22744 18785 22753 18819
rect 22753 18785 22787 18819
rect 22787 18785 22796 18819
rect 22744 18776 22796 18785
rect 22928 18887 22980 18896
rect 22928 18853 22937 18887
rect 22937 18853 22971 18887
rect 22971 18853 22980 18887
rect 22928 18844 22980 18853
rect 23388 18844 23440 18896
rect 23204 18819 23256 18828
rect 23204 18785 23213 18819
rect 23213 18785 23247 18819
rect 23247 18785 23256 18819
rect 23204 18776 23256 18785
rect 25504 18776 25556 18828
rect 24952 18640 25004 18692
rect 18880 18572 18932 18624
rect 19156 18572 19208 18624
rect 20904 18572 20956 18624
rect 21088 18572 21140 18624
rect 22468 18572 22520 18624
rect 22836 18572 22888 18624
rect 3756 18470 3808 18522
rect 3820 18470 3872 18522
rect 3884 18470 3936 18522
rect 3948 18470 4000 18522
rect 4012 18470 4064 18522
rect 10472 18470 10524 18522
rect 10536 18470 10588 18522
rect 10600 18470 10652 18522
rect 10664 18470 10716 18522
rect 10728 18470 10780 18522
rect 17188 18470 17240 18522
rect 17252 18470 17304 18522
rect 17316 18470 17368 18522
rect 17380 18470 17432 18522
rect 17444 18470 17496 18522
rect 23904 18470 23956 18522
rect 23968 18470 24020 18522
rect 24032 18470 24084 18522
rect 24096 18470 24148 18522
rect 24160 18470 24212 18522
rect 5080 18368 5132 18420
rect 6092 18411 6144 18420
rect 6092 18377 6101 18411
rect 6101 18377 6135 18411
rect 6135 18377 6144 18411
rect 6092 18368 6144 18377
rect 7288 18411 7340 18420
rect 7288 18377 7297 18411
rect 7297 18377 7331 18411
rect 7331 18377 7340 18411
rect 7288 18368 7340 18377
rect 8576 18411 8628 18420
rect 8576 18377 8585 18411
rect 8585 18377 8619 18411
rect 8619 18377 8628 18411
rect 8576 18368 8628 18377
rect 13176 18368 13228 18420
rect 16672 18411 16724 18420
rect 16672 18377 16681 18411
rect 16681 18377 16715 18411
rect 16715 18377 16724 18411
rect 16672 18368 16724 18377
rect 17684 18368 17736 18420
rect 18604 18368 18656 18420
rect 21180 18411 21232 18420
rect 21180 18377 21189 18411
rect 21189 18377 21223 18411
rect 21223 18377 21232 18411
rect 21180 18368 21232 18377
rect 21548 18368 21600 18420
rect 6460 18300 6512 18352
rect 5264 18232 5316 18284
rect 5632 18232 5684 18284
rect 1308 18207 1360 18216
rect 1308 18173 1317 18207
rect 1317 18173 1351 18207
rect 1351 18173 1360 18207
rect 1308 18164 1360 18173
rect 2044 18207 2096 18216
rect 2044 18173 2053 18207
rect 2053 18173 2087 18207
rect 2087 18173 2096 18207
rect 2044 18164 2096 18173
rect 2228 18207 2280 18216
rect 2228 18173 2237 18207
rect 2237 18173 2271 18207
rect 2271 18173 2280 18207
rect 2228 18164 2280 18173
rect 4528 18207 4580 18216
rect 4528 18173 4537 18207
rect 4537 18173 4571 18207
rect 4571 18173 4580 18207
rect 4528 18164 4580 18173
rect 4988 18207 5040 18216
rect 4988 18173 4997 18207
rect 4997 18173 5031 18207
rect 5031 18173 5040 18207
rect 4988 18164 5040 18173
rect 2688 18139 2740 18148
rect 2688 18105 2697 18139
rect 2697 18105 2731 18139
rect 2731 18105 2740 18139
rect 2688 18096 2740 18105
rect 4804 18139 4856 18148
rect 4804 18105 4813 18139
rect 4813 18105 4847 18139
rect 4847 18105 4856 18139
rect 5540 18207 5592 18216
rect 5540 18173 5550 18207
rect 5550 18173 5584 18207
rect 5584 18173 5592 18207
rect 6552 18232 6604 18284
rect 7564 18232 7616 18284
rect 5540 18164 5592 18173
rect 6368 18207 6420 18216
rect 6368 18173 6377 18207
rect 6377 18173 6411 18207
rect 6411 18173 6420 18207
rect 6368 18164 6420 18173
rect 7656 18164 7708 18216
rect 8944 18164 8996 18216
rect 4804 18096 4856 18105
rect 9496 18096 9548 18148
rect 9588 18096 9640 18148
rect 11244 18164 11296 18216
rect 12072 18164 12124 18216
rect 13360 18207 13412 18216
rect 13360 18173 13369 18207
rect 13369 18173 13403 18207
rect 13403 18173 13412 18207
rect 13360 18164 13412 18173
rect 14372 18207 14424 18216
rect 14372 18173 14376 18207
rect 14376 18173 14410 18207
rect 14410 18173 14424 18207
rect 14372 18164 14424 18173
rect 15752 18232 15804 18284
rect 16304 18300 16356 18352
rect 21456 18300 21508 18352
rect 16580 18232 16632 18284
rect 10968 18096 11020 18148
rect 11152 18096 11204 18148
rect 1124 18071 1176 18080
rect 1124 18037 1133 18071
rect 1133 18037 1167 18071
rect 1167 18037 1176 18071
rect 1124 18028 1176 18037
rect 1860 18071 1912 18080
rect 1860 18037 1869 18071
rect 1869 18037 1903 18071
rect 1903 18037 1912 18071
rect 1860 18028 1912 18037
rect 1952 18028 2004 18080
rect 5448 18028 5500 18080
rect 6000 18028 6052 18080
rect 6276 18071 6328 18080
rect 6276 18037 6285 18071
rect 6285 18037 6319 18071
rect 6319 18037 6328 18071
rect 6276 18028 6328 18037
rect 7840 18028 7892 18080
rect 8300 18028 8352 18080
rect 11428 18028 11480 18080
rect 12808 18096 12860 18148
rect 15016 18164 15068 18216
rect 15108 18207 15160 18216
rect 15108 18173 15117 18207
rect 15117 18173 15151 18207
rect 15151 18173 15160 18207
rect 15108 18164 15160 18173
rect 16304 18164 16356 18216
rect 17868 18232 17920 18284
rect 17684 18207 17736 18216
rect 17684 18173 17693 18207
rect 17693 18173 17727 18207
rect 17727 18173 17736 18207
rect 17684 18164 17736 18173
rect 17776 18207 17828 18216
rect 17776 18173 17785 18207
rect 17785 18173 17819 18207
rect 17819 18173 17828 18207
rect 17776 18164 17828 18173
rect 17960 18207 18012 18216
rect 17960 18173 17969 18207
rect 17969 18173 18003 18207
rect 18003 18173 18012 18207
rect 17960 18164 18012 18173
rect 18144 18207 18196 18216
rect 18144 18173 18153 18207
rect 18153 18173 18187 18207
rect 18187 18173 18196 18207
rect 18144 18164 18196 18173
rect 18972 18207 19024 18216
rect 18972 18173 18981 18207
rect 18981 18173 19015 18207
rect 19015 18173 19024 18207
rect 18972 18164 19024 18173
rect 20904 18207 20956 18216
rect 20904 18173 20913 18207
rect 20913 18173 20947 18207
rect 20947 18173 20956 18207
rect 20904 18164 20956 18173
rect 12072 18071 12124 18080
rect 12072 18037 12081 18071
rect 12081 18037 12115 18071
rect 12115 18037 12124 18071
rect 12072 18028 12124 18037
rect 13636 18071 13688 18080
rect 13636 18037 13645 18071
rect 13645 18037 13679 18071
rect 13679 18037 13688 18071
rect 13636 18028 13688 18037
rect 14188 18071 14240 18080
rect 14188 18037 14197 18071
rect 14197 18037 14231 18071
rect 14231 18037 14240 18071
rect 14188 18028 14240 18037
rect 14280 18028 14332 18080
rect 15844 18096 15896 18148
rect 16120 18096 16172 18148
rect 19432 18096 19484 18148
rect 21180 18164 21232 18216
rect 21364 18207 21416 18216
rect 21364 18173 21373 18207
rect 21373 18173 21407 18207
rect 21407 18173 21416 18207
rect 21364 18164 21416 18173
rect 22468 18368 22520 18420
rect 23296 18368 23348 18420
rect 23388 18368 23440 18420
rect 25504 18411 25556 18420
rect 25504 18377 25513 18411
rect 25513 18377 25547 18411
rect 25547 18377 25556 18411
rect 25504 18368 25556 18377
rect 24400 18300 24452 18352
rect 24860 18300 24912 18352
rect 21824 18232 21876 18284
rect 22560 18232 22612 18284
rect 23204 18275 23256 18284
rect 23204 18241 23213 18275
rect 23213 18241 23247 18275
rect 23247 18241 23256 18275
rect 23204 18232 23256 18241
rect 21732 18096 21784 18148
rect 22376 18096 22428 18148
rect 22836 18096 22888 18148
rect 15200 18028 15252 18080
rect 15292 18071 15344 18080
rect 15292 18037 15301 18071
rect 15301 18037 15335 18071
rect 15335 18037 15344 18071
rect 15292 18028 15344 18037
rect 15384 18028 15436 18080
rect 17592 18028 17644 18080
rect 17776 18028 17828 18080
rect 22100 18071 22152 18080
rect 22100 18037 22109 18071
rect 22109 18037 22143 18071
rect 22143 18037 22152 18071
rect 22100 18028 22152 18037
rect 24400 18207 24452 18216
rect 24400 18173 24409 18207
rect 24409 18173 24443 18207
rect 24443 18173 24452 18207
rect 24400 18164 24452 18173
rect 24768 18164 24820 18216
rect 27068 18207 27120 18216
rect 27068 18173 27077 18207
rect 27077 18173 27111 18207
rect 27111 18173 27120 18207
rect 27068 18164 27120 18173
rect 25136 18139 25188 18148
rect 25136 18105 25145 18139
rect 25145 18105 25179 18139
rect 25179 18105 25188 18139
rect 25136 18096 25188 18105
rect 25504 18096 25556 18148
rect 26608 18096 26660 18148
rect 23940 18028 23992 18080
rect 25780 18028 25832 18080
rect 26148 18028 26200 18080
rect 7114 17926 7166 17978
rect 7178 17926 7230 17978
rect 7242 17926 7294 17978
rect 7306 17926 7358 17978
rect 7370 17926 7422 17978
rect 13830 17926 13882 17978
rect 13894 17926 13946 17978
rect 13958 17926 14010 17978
rect 14022 17926 14074 17978
rect 14086 17926 14138 17978
rect 20546 17926 20598 17978
rect 20610 17926 20662 17978
rect 20674 17926 20726 17978
rect 20738 17926 20790 17978
rect 20802 17926 20854 17978
rect 27262 17926 27314 17978
rect 27326 17926 27378 17978
rect 27390 17926 27442 17978
rect 27454 17926 27506 17978
rect 27518 17926 27570 17978
rect 2228 17867 2280 17876
rect 2228 17833 2237 17867
rect 2237 17833 2271 17867
rect 2271 17833 2280 17867
rect 2228 17824 2280 17833
rect 4528 17824 4580 17876
rect 4804 17824 4856 17876
rect 1124 17799 1176 17808
rect 1124 17765 1158 17799
rect 1158 17765 1176 17799
rect 1124 17756 1176 17765
rect 848 17731 900 17740
rect 848 17697 857 17731
rect 857 17697 891 17731
rect 891 17697 900 17731
rect 848 17688 900 17697
rect 3056 17688 3108 17740
rect 4528 17688 4580 17740
rect 2504 17663 2556 17672
rect 2504 17629 2513 17663
rect 2513 17629 2547 17663
rect 2547 17629 2556 17663
rect 2504 17620 2556 17629
rect 2688 17663 2740 17672
rect 2688 17629 2697 17663
rect 2697 17629 2731 17663
rect 2731 17629 2740 17663
rect 2688 17620 2740 17629
rect 4160 17620 4212 17672
rect 3240 17552 3292 17604
rect 5172 17731 5224 17740
rect 5172 17697 5181 17731
rect 5181 17697 5215 17731
rect 5215 17697 5224 17731
rect 5172 17688 5224 17697
rect 5540 17756 5592 17808
rect 6460 17688 6512 17740
rect 6920 17799 6972 17808
rect 6920 17765 6929 17799
rect 6929 17765 6963 17799
rect 6963 17765 6972 17799
rect 6920 17756 6972 17765
rect 7288 17824 7340 17876
rect 10048 17867 10100 17876
rect 10048 17833 10057 17867
rect 10057 17833 10091 17867
rect 10091 17833 10100 17867
rect 10048 17824 10100 17833
rect 10968 17867 11020 17876
rect 10968 17833 10977 17867
rect 10977 17833 11011 17867
rect 11011 17833 11020 17867
rect 10968 17824 11020 17833
rect 12072 17824 12124 17876
rect 13360 17824 13412 17876
rect 7472 17756 7524 17808
rect 7472 17620 7524 17672
rect 8668 17663 8720 17672
rect 8668 17629 8677 17663
rect 8677 17629 8711 17663
rect 8711 17629 8720 17663
rect 8668 17620 8720 17629
rect 2872 17527 2924 17536
rect 2872 17493 2881 17527
rect 2881 17493 2915 17527
rect 2915 17493 2924 17527
rect 2872 17484 2924 17493
rect 3332 17527 3384 17536
rect 3332 17493 3341 17527
rect 3341 17493 3375 17527
rect 3375 17493 3384 17527
rect 3332 17484 3384 17493
rect 4344 17484 4396 17536
rect 5540 17484 5592 17536
rect 5632 17484 5684 17536
rect 7840 17552 7892 17604
rect 10232 17688 10284 17740
rect 11152 17731 11204 17740
rect 11152 17697 11161 17731
rect 11161 17697 11195 17731
rect 11195 17697 11204 17731
rect 11152 17688 11204 17697
rect 11428 17731 11480 17740
rect 11428 17697 11437 17731
rect 11437 17697 11471 17731
rect 11471 17697 11480 17731
rect 11428 17688 11480 17697
rect 11520 17731 11572 17740
rect 11520 17697 11529 17731
rect 11529 17697 11563 17731
rect 11563 17697 11572 17731
rect 11520 17688 11572 17697
rect 12440 17731 12492 17740
rect 12440 17697 12474 17731
rect 12474 17697 12492 17731
rect 12440 17688 12492 17697
rect 14280 17824 14332 17876
rect 15660 17824 15712 17876
rect 17960 17824 18012 17876
rect 21364 17824 21416 17876
rect 23204 17824 23256 17876
rect 24400 17824 24452 17876
rect 24860 17824 24912 17876
rect 26608 17867 26660 17876
rect 26608 17833 26617 17867
rect 26617 17833 26651 17867
rect 26651 17833 26660 17867
rect 26608 17824 26660 17833
rect 15292 17756 15344 17808
rect 14188 17688 14240 17740
rect 11888 17620 11940 17672
rect 11152 17552 11204 17604
rect 15108 17688 15160 17740
rect 15384 17620 15436 17672
rect 15292 17552 15344 17604
rect 15844 17688 15896 17740
rect 17868 17799 17920 17808
rect 17868 17765 17877 17799
rect 17877 17765 17911 17799
rect 17911 17765 17920 17799
rect 17868 17756 17920 17765
rect 21180 17756 21232 17808
rect 16948 17688 17000 17740
rect 18236 17688 18288 17740
rect 19156 17731 19208 17740
rect 19156 17697 19165 17731
rect 19165 17697 19199 17731
rect 19199 17697 19208 17731
rect 19156 17688 19208 17697
rect 6460 17527 6512 17536
rect 6460 17493 6469 17527
rect 6469 17493 6503 17527
rect 6503 17493 6512 17527
rect 6460 17484 6512 17493
rect 8116 17484 8168 17536
rect 9036 17484 9088 17536
rect 14740 17484 14792 17536
rect 15752 17484 15804 17536
rect 18328 17620 18380 17672
rect 19708 17731 19760 17740
rect 19708 17697 19717 17731
rect 19717 17697 19751 17731
rect 19751 17697 19760 17731
rect 19708 17688 19760 17697
rect 19892 17688 19944 17740
rect 20352 17688 20404 17740
rect 20996 17688 21048 17740
rect 21548 17731 21600 17740
rect 21548 17697 21557 17731
rect 21557 17697 21591 17731
rect 21591 17697 21600 17731
rect 21548 17688 21600 17697
rect 21640 17731 21692 17740
rect 21640 17697 21649 17731
rect 21649 17697 21683 17731
rect 21683 17697 21692 17731
rect 21640 17688 21692 17697
rect 21916 17731 21968 17740
rect 21916 17697 21925 17731
rect 21925 17697 21959 17731
rect 21959 17697 21968 17731
rect 21916 17688 21968 17697
rect 22192 17731 22244 17740
rect 22192 17697 22205 17731
rect 22205 17697 22244 17731
rect 22192 17688 22244 17697
rect 23940 17731 23992 17740
rect 23940 17697 23958 17731
rect 23958 17697 23992 17731
rect 24768 17756 24820 17808
rect 23940 17688 23992 17697
rect 24676 17688 24728 17740
rect 25688 17688 25740 17740
rect 25780 17731 25832 17740
rect 25780 17697 25789 17731
rect 25789 17697 25823 17731
rect 25823 17697 25832 17731
rect 25780 17688 25832 17697
rect 27068 17756 27120 17808
rect 25964 17731 26016 17740
rect 25964 17697 25973 17731
rect 25973 17697 26007 17731
rect 26007 17697 26016 17731
rect 25964 17688 26016 17697
rect 26148 17688 26200 17740
rect 26424 17731 26476 17740
rect 26424 17697 26433 17731
rect 26433 17697 26467 17731
rect 26467 17697 26476 17731
rect 26424 17688 26476 17697
rect 16856 17552 16908 17604
rect 19340 17552 19392 17604
rect 22100 17552 22152 17604
rect 22468 17552 22520 17604
rect 22928 17552 22980 17604
rect 24952 17552 25004 17604
rect 25044 17552 25096 17604
rect 16764 17484 16816 17536
rect 17592 17484 17644 17536
rect 19524 17484 19576 17536
rect 24308 17527 24360 17536
rect 24308 17493 24317 17527
rect 24317 17493 24351 17527
rect 24351 17493 24360 17527
rect 24308 17484 24360 17493
rect 25504 17527 25556 17536
rect 25504 17493 25513 17527
rect 25513 17493 25547 17527
rect 25547 17493 25556 17527
rect 25504 17484 25556 17493
rect 26424 17484 26476 17536
rect 3756 17382 3808 17434
rect 3820 17382 3872 17434
rect 3884 17382 3936 17434
rect 3948 17382 4000 17434
rect 4012 17382 4064 17434
rect 10472 17382 10524 17434
rect 10536 17382 10588 17434
rect 10600 17382 10652 17434
rect 10664 17382 10716 17434
rect 10728 17382 10780 17434
rect 17188 17382 17240 17434
rect 17252 17382 17304 17434
rect 17316 17382 17368 17434
rect 17380 17382 17432 17434
rect 17444 17382 17496 17434
rect 23904 17382 23956 17434
rect 23968 17382 24020 17434
rect 24032 17382 24084 17434
rect 24096 17382 24148 17434
rect 24160 17382 24212 17434
rect 1308 17323 1360 17332
rect 1308 17289 1317 17323
rect 1317 17289 1351 17323
rect 1351 17289 1360 17323
rect 1308 17280 1360 17289
rect 1492 17323 1544 17332
rect 1492 17289 1501 17323
rect 1501 17289 1535 17323
rect 1535 17289 1544 17323
rect 1492 17280 1544 17289
rect 2228 17323 2280 17332
rect 2228 17289 2237 17323
rect 2237 17289 2271 17323
rect 2271 17289 2280 17323
rect 2228 17280 2280 17289
rect 1860 17255 1912 17264
rect 1860 17221 1869 17255
rect 1869 17221 1903 17255
rect 1903 17221 1912 17255
rect 1860 17212 1912 17221
rect 2504 17255 2556 17264
rect 2504 17221 2513 17255
rect 2513 17221 2547 17255
rect 2547 17221 2556 17255
rect 2504 17212 2556 17221
rect 3056 17323 3108 17332
rect 3056 17289 3065 17323
rect 3065 17289 3099 17323
rect 3099 17289 3108 17323
rect 3056 17280 3108 17289
rect 3240 17323 3292 17332
rect 3240 17289 3249 17323
rect 3249 17289 3283 17323
rect 3283 17289 3292 17323
rect 3240 17280 3292 17289
rect 5172 17280 5224 17332
rect 5264 17280 5316 17332
rect 2688 17144 2740 17196
rect 5448 17212 5500 17264
rect 6276 17280 6328 17332
rect 8668 17280 8720 17332
rect 12440 17280 12492 17332
rect 15384 17280 15436 17332
rect 16672 17280 16724 17332
rect 18052 17280 18104 17332
rect 22100 17280 22152 17332
rect 15200 17212 15252 17264
rect 15292 17212 15344 17264
rect 5356 17144 5408 17196
rect 6552 17144 6604 17196
rect 11428 17144 11480 17196
rect 1952 17008 2004 17060
rect 4344 17119 4396 17128
rect 4344 17085 4362 17119
rect 4362 17085 4396 17119
rect 4344 17076 4396 17085
rect 2872 17051 2924 17060
rect 2872 17017 2881 17051
rect 2881 17017 2915 17051
rect 2915 17017 2924 17051
rect 2872 17008 2924 17017
rect 4896 17119 4948 17128
rect 4896 17085 4905 17119
rect 4905 17085 4939 17119
rect 4939 17085 4948 17119
rect 4896 17076 4948 17085
rect 4988 17076 5040 17128
rect 5632 17119 5684 17128
rect 5632 17085 5641 17119
rect 5641 17085 5675 17119
rect 5675 17085 5684 17119
rect 5632 17076 5684 17085
rect 6460 17119 6512 17128
rect 6460 17085 6469 17119
rect 6469 17085 6503 17119
rect 6503 17085 6512 17119
rect 6460 17076 6512 17085
rect 6644 17119 6696 17128
rect 6644 17085 6653 17119
rect 6653 17085 6687 17119
rect 6687 17085 6696 17119
rect 6644 17076 6696 17085
rect 7564 17076 7616 17128
rect 8392 17076 8444 17128
rect 9036 17119 9088 17128
rect 9036 17085 9070 17119
rect 9070 17085 9088 17119
rect 9036 17076 9088 17085
rect 6092 17008 6144 17060
rect 7656 17008 7708 17060
rect 11060 17119 11112 17128
rect 11060 17085 11069 17119
rect 11069 17085 11103 17119
rect 11103 17085 11112 17119
rect 11060 17076 11112 17085
rect 13636 17144 13688 17196
rect 15752 17187 15804 17196
rect 15752 17153 15761 17187
rect 15761 17153 15795 17187
rect 15795 17153 15804 17187
rect 15752 17144 15804 17153
rect 17960 17212 18012 17264
rect 13084 17119 13136 17128
rect 13084 17085 13093 17119
rect 13093 17085 13127 17119
rect 13127 17085 13136 17119
rect 13084 17076 13136 17085
rect 13544 17076 13596 17128
rect 12716 17008 12768 17060
rect 16856 17076 16908 17128
rect 17592 17076 17644 17128
rect 18052 17076 18104 17128
rect 18328 17119 18380 17128
rect 18328 17085 18337 17119
rect 18337 17085 18371 17119
rect 18371 17085 18380 17119
rect 18328 17076 18380 17085
rect 21548 17144 21600 17196
rect 18972 17076 19024 17128
rect 20996 17119 21048 17128
rect 20996 17085 21005 17119
rect 21005 17085 21039 17119
rect 21039 17085 21048 17119
rect 20996 17076 21048 17085
rect 21456 17119 21508 17128
rect 21456 17085 21465 17119
rect 21465 17085 21499 17119
rect 21499 17085 21508 17119
rect 21456 17076 21508 17085
rect 22284 17076 22336 17128
rect 22928 17076 22980 17128
rect 23204 17119 23256 17128
rect 23204 17085 23213 17119
rect 23213 17085 23247 17119
rect 23247 17085 23256 17119
rect 23204 17076 23256 17085
rect 17868 17008 17920 17060
rect 18236 17051 18288 17060
rect 18236 17017 18245 17051
rect 18245 17017 18279 17051
rect 18279 17017 18288 17051
rect 18236 17008 18288 17017
rect 18420 17008 18472 17060
rect 1860 16940 1912 16992
rect 4160 16940 4212 16992
rect 5356 16940 5408 16992
rect 5448 16940 5500 16992
rect 6368 16940 6420 16992
rect 10140 16983 10192 16992
rect 10140 16949 10149 16983
rect 10149 16949 10183 16983
rect 10183 16949 10192 16983
rect 10140 16940 10192 16949
rect 10324 16983 10376 16992
rect 10324 16949 10333 16983
rect 10333 16949 10367 16983
rect 10367 16949 10376 16983
rect 10324 16940 10376 16949
rect 10692 16983 10744 16992
rect 10692 16949 10701 16983
rect 10701 16949 10735 16983
rect 10735 16949 10744 16983
rect 10692 16940 10744 16949
rect 12532 16940 12584 16992
rect 13452 16940 13504 16992
rect 13820 16940 13872 16992
rect 16856 16940 16908 16992
rect 17224 16940 17276 16992
rect 19248 17008 19300 17060
rect 22008 17008 22060 17060
rect 20996 16940 21048 16992
rect 22376 16940 22428 16992
rect 23572 17008 23624 17060
rect 24124 17076 24176 17128
rect 25044 17119 25096 17128
rect 25044 17085 25053 17119
rect 25053 17085 25087 17119
rect 25087 17085 25096 17119
rect 25044 17076 25096 17085
rect 25688 17119 25740 17128
rect 25688 17085 25697 17119
rect 25697 17085 25731 17119
rect 25731 17085 25740 17119
rect 25688 17076 25740 17085
rect 24952 17008 25004 17060
rect 24400 16940 24452 16992
rect 25320 16940 25372 16992
rect 26056 17008 26108 17060
rect 7114 16838 7166 16890
rect 7178 16838 7230 16890
rect 7242 16838 7294 16890
rect 7306 16838 7358 16890
rect 7370 16838 7422 16890
rect 13830 16838 13882 16890
rect 13894 16838 13946 16890
rect 13958 16838 14010 16890
rect 14022 16838 14074 16890
rect 14086 16838 14138 16890
rect 20546 16838 20598 16890
rect 20610 16838 20662 16890
rect 20674 16838 20726 16890
rect 20738 16838 20790 16890
rect 20802 16838 20854 16890
rect 27262 16838 27314 16890
rect 27326 16838 27378 16890
rect 27390 16838 27442 16890
rect 27454 16838 27506 16890
rect 27518 16838 27570 16890
rect 1584 16736 1636 16788
rect 2412 16736 2464 16788
rect 2688 16736 2740 16788
rect 4344 16736 4396 16788
rect 4988 16736 5040 16788
rect 5448 16779 5500 16788
rect 5448 16745 5457 16779
rect 5457 16745 5491 16779
rect 5491 16745 5500 16779
rect 5448 16736 5500 16745
rect 7472 16779 7524 16788
rect 7472 16745 7481 16779
rect 7481 16745 7515 16779
rect 7515 16745 7524 16779
rect 7472 16736 7524 16745
rect 7656 16779 7708 16788
rect 7656 16745 7665 16779
rect 7665 16745 7699 16779
rect 7699 16745 7708 16779
rect 7656 16736 7708 16745
rect 8024 16779 8076 16788
rect 8024 16745 8033 16779
rect 8033 16745 8067 16779
rect 8067 16745 8076 16779
rect 8024 16736 8076 16745
rect 10140 16736 10192 16788
rect 10232 16779 10284 16788
rect 10232 16745 10241 16779
rect 10241 16745 10275 16779
rect 10275 16745 10284 16779
rect 10232 16736 10284 16745
rect 11336 16736 11388 16788
rect 12808 16736 12860 16788
rect 13728 16736 13780 16788
rect 14464 16736 14516 16788
rect 15292 16736 15344 16788
rect 2504 16643 2556 16652
rect 2504 16609 2513 16643
rect 2513 16609 2547 16643
rect 2547 16609 2556 16643
rect 2504 16600 2556 16609
rect 3332 16600 3384 16652
rect 7564 16668 7616 16720
rect 5264 16600 5316 16652
rect 6092 16643 6144 16652
rect 6092 16609 6101 16643
rect 6101 16609 6135 16643
rect 6135 16609 6144 16643
rect 6092 16600 6144 16609
rect 6368 16643 6420 16652
rect 6368 16609 6402 16643
rect 6402 16609 6420 16643
rect 6368 16600 6420 16609
rect 6644 16600 6696 16652
rect 6828 16600 6880 16652
rect 7840 16643 7892 16652
rect 7840 16609 7849 16643
rect 7849 16609 7883 16643
rect 7883 16609 7892 16643
rect 7840 16600 7892 16609
rect 10692 16668 10744 16720
rect 2596 16464 2648 16516
rect 9128 16532 9180 16584
rect 10324 16643 10376 16652
rect 10324 16609 10333 16643
rect 10333 16609 10367 16643
rect 10367 16609 10376 16643
rect 10324 16600 10376 16609
rect 12716 16668 12768 16720
rect 14188 16711 14240 16720
rect 14188 16677 14197 16711
rect 14197 16677 14231 16711
rect 14231 16677 14240 16711
rect 14188 16668 14240 16677
rect 11428 16643 11480 16652
rect 11428 16609 11437 16643
rect 11437 16609 11471 16643
rect 11471 16609 11480 16643
rect 11428 16600 11480 16609
rect 13636 16600 13688 16652
rect 14464 16643 14516 16652
rect 14464 16609 14473 16643
rect 14473 16609 14507 16643
rect 14507 16609 14516 16643
rect 14464 16600 14516 16609
rect 14740 16643 14792 16652
rect 14740 16609 14749 16643
rect 14749 16609 14783 16643
rect 14783 16609 14792 16643
rect 14740 16600 14792 16609
rect 15844 16668 15896 16720
rect 16948 16779 17000 16788
rect 16948 16745 16957 16779
rect 16957 16745 16991 16779
rect 16991 16745 17000 16779
rect 16948 16736 17000 16745
rect 17684 16736 17736 16788
rect 18328 16736 18380 16788
rect 16672 16668 16724 16720
rect 15200 16600 15252 16652
rect 15292 16643 15344 16652
rect 15292 16609 15301 16643
rect 15301 16609 15335 16643
rect 15335 16609 15344 16643
rect 15292 16600 15344 16609
rect 15568 16643 15620 16652
rect 15568 16609 15577 16643
rect 15577 16609 15611 16643
rect 15611 16609 15620 16643
rect 15568 16600 15620 16609
rect 11152 16532 11204 16584
rect 13820 16575 13872 16584
rect 13820 16541 13829 16575
rect 13829 16541 13863 16575
rect 13863 16541 13872 16575
rect 13820 16532 13872 16541
rect 15108 16575 15160 16584
rect 15108 16541 15117 16575
rect 15117 16541 15151 16575
rect 15151 16541 15160 16575
rect 15108 16532 15160 16541
rect 15936 16600 15988 16652
rect 16488 16600 16540 16652
rect 17224 16643 17276 16652
rect 17224 16609 17233 16643
rect 17233 16609 17267 16643
rect 17267 16609 17276 16643
rect 17224 16600 17276 16609
rect 17960 16668 18012 16720
rect 17592 16643 17644 16652
rect 17592 16609 17626 16643
rect 17626 16609 17644 16643
rect 17592 16600 17644 16609
rect 20352 16779 20404 16788
rect 20352 16745 20361 16779
rect 20361 16745 20395 16779
rect 20395 16745 20404 16779
rect 20352 16736 20404 16745
rect 21916 16779 21968 16788
rect 21916 16745 21925 16779
rect 21925 16745 21959 16779
rect 21959 16745 21968 16779
rect 21916 16736 21968 16745
rect 22008 16779 22060 16788
rect 22008 16745 22017 16779
rect 22017 16745 22051 16779
rect 22051 16745 22060 16779
rect 22008 16736 22060 16745
rect 24124 16779 24176 16788
rect 24124 16745 24133 16779
rect 24133 16745 24167 16779
rect 24167 16745 24176 16779
rect 24124 16736 24176 16745
rect 24676 16736 24728 16788
rect 25320 16779 25372 16788
rect 25320 16745 25329 16779
rect 25329 16745 25363 16779
rect 25363 16745 25372 16779
rect 25320 16736 25372 16745
rect 20996 16668 21048 16720
rect 19800 16600 19852 16652
rect 21548 16600 21600 16652
rect 20260 16575 20312 16584
rect 20260 16541 20269 16575
rect 20269 16541 20303 16575
rect 20303 16541 20312 16575
rect 20260 16532 20312 16541
rect 21088 16532 21140 16584
rect 2504 16396 2556 16448
rect 4896 16464 4948 16516
rect 21456 16532 21508 16584
rect 22284 16643 22336 16652
rect 22284 16609 22293 16643
rect 22293 16609 22327 16643
rect 22327 16609 22336 16643
rect 22284 16600 22336 16609
rect 22376 16643 22428 16652
rect 22376 16609 22385 16643
rect 22385 16609 22419 16643
rect 22419 16609 22428 16643
rect 22376 16600 22428 16609
rect 22928 16668 22980 16720
rect 22836 16600 22888 16652
rect 23020 16643 23072 16652
rect 23020 16609 23054 16643
rect 23054 16609 23072 16643
rect 23020 16600 23072 16609
rect 24308 16668 24360 16720
rect 24584 16668 24636 16720
rect 22652 16532 22704 16584
rect 24400 16643 24452 16652
rect 24400 16609 24409 16643
rect 24409 16609 24443 16643
rect 24443 16609 24452 16643
rect 24400 16600 24452 16609
rect 24860 16643 24912 16652
rect 24860 16609 24869 16643
rect 24869 16609 24903 16643
rect 24903 16609 24912 16643
rect 24860 16600 24912 16609
rect 26056 16779 26108 16788
rect 26056 16745 26065 16779
rect 26065 16745 26099 16779
rect 26099 16745 26108 16779
rect 26056 16736 26108 16745
rect 4160 16396 4212 16448
rect 4528 16439 4580 16448
rect 4528 16405 4537 16439
rect 4537 16405 4571 16439
rect 4571 16405 4580 16439
rect 4528 16396 4580 16405
rect 21640 16464 21692 16516
rect 9312 16439 9364 16448
rect 9312 16405 9321 16439
rect 9321 16405 9355 16439
rect 9355 16405 9364 16439
rect 9312 16396 9364 16405
rect 11060 16439 11112 16448
rect 11060 16405 11069 16439
rect 11069 16405 11103 16439
rect 11103 16405 11112 16439
rect 11060 16396 11112 16405
rect 12624 16396 12676 16448
rect 13176 16396 13228 16448
rect 15752 16439 15804 16448
rect 15752 16405 15761 16439
rect 15761 16405 15795 16439
rect 15795 16405 15804 16439
rect 15752 16396 15804 16405
rect 16764 16439 16816 16448
rect 16764 16405 16773 16439
rect 16773 16405 16807 16439
rect 16807 16405 16816 16439
rect 16764 16396 16816 16405
rect 18788 16439 18840 16448
rect 18788 16405 18797 16439
rect 18797 16405 18831 16439
rect 18831 16405 18840 16439
rect 18788 16396 18840 16405
rect 19340 16396 19392 16448
rect 24860 16396 24912 16448
rect 25504 16396 25556 16448
rect 3756 16294 3808 16346
rect 3820 16294 3872 16346
rect 3884 16294 3936 16346
rect 3948 16294 4000 16346
rect 4012 16294 4064 16346
rect 10472 16294 10524 16346
rect 10536 16294 10588 16346
rect 10600 16294 10652 16346
rect 10664 16294 10716 16346
rect 10728 16294 10780 16346
rect 17188 16294 17240 16346
rect 17252 16294 17304 16346
rect 17316 16294 17368 16346
rect 17380 16294 17432 16346
rect 17444 16294 17496 16346
rect 23904 16294 23956 16346
rect 23968 16294 24020 16346
rect 24032 16294 24084 16346
rect 24096 16294 24148 16346
rect 24160 16294 24212 16346
rect 4344 16235 4396 16244
rect 4344 16201 4353 16235
rect 4353 16201 4387 16235
rect 4387 16201 4396 16235
rect 4344 16192 4396 16201
rect 2228 16124 2280 16176
rect 2504 16124 2556 16176
rect 1860 16056 1912 16108
rect 5816 16056 5868 16108
rect 1952 15988 2004 16040
rect 2412 15988 2464 16040
rect 2504 16031 2556 16040
rect 2504 15997 2513 16031
rect 2513 15997 2547 16031
rect 2547 15997 2556 16031
rect 2504 15988 2556 15997
rect 3332 15988 3384 16040
rect 4620 15988 4672 16040
rect 4804 15988 4856 16040
rect 6460 15988 6512 16040
rect 11060 16192 11112 16244
rect 13176 16192 13228 16244
rect 15108 16192 15160 16244
rect 15568 16192 15620 16244
rect 17592 16192 17644 16244
rect 22376 16192 22428 16244
rect 23020 16235 23072 16244
rect 23020 16201 23029 16235
rect 23029 16201 23063 16235
rect 23063 16201 23072 16235
rect 23020 16192 23072 16201
rect 21456 16056 21508 16108
rect 11888 16031 11940 16040
rect 4160 15920 4212 15972
rect 9680 15920 9732 15972
rect 11888 15997 11897 16031
rect 11897 15997 11931 16031
rect 11931 15997 11940 16031
rect 11888 15988 11940 15997
rect 1492 15852 1544 15904
rect 4620 15852 4672 15904
rect 6552 15895 6604 15904
rect 6552 15861 6561 15895
rect 6561 15861 6595 15895
rect 6595 15861 6604 15895
rect 6552 15852 6604 15861
rect 12440 15920 12492 15972
rect 11244 15852 11296 15904
rect 13820 15988 13872 16040
rect 15200 16031 15252 16040
rect 15200 15997 15209 16031
rect 15209 15997 15243 16031
rect 15243 15997 15252 16031
rect 15200 15988 15252 15997
rect 13728 15963 13780 15972
rect 13728 15929 13755 15963
rect 13755 15929 13780 15963
rect 13728 15920 13780 15929
rect 14464 15920 14516 15972
rect 15660 16031 15712 16040
rect 15660 15997 15669 16031
rect 15669 15997 15703 16031
rect 15703 15997 15712 16031
rect 15660 15988 15712 15997
rect 17684 16031 17736 16040
rect 17684 15997 17693 16031
rect 17693 15997 17727 16031
rect 17727 15997 17736 16031
rect 17684 15988 17736 15997
rect 17868 16031 17920 16040
rect 17868 15997 17877 16031
rect 17877 15997 17911 16031
rect 17911 15997 17920 16031
rect 17868 15988 17920 15997
rect 18788 15988 18840 16040
rect 19248 16031 19300 16040
rect 19248 15997 19257 16031
rect 19257 15997 19291 16031
rect 19291 15997 19300 16031
rect 19248 15988 19300 15997
rect 19524 16031 19576 16040
rect 19524 15997 19558 16031
rect 19558 15997 19576 16031
rect 19524 15988 19576 15997
rect 19800 15988 19852 16040
rect 21088 16031 21140 16040
rect 21088 15997 21097 16031
rect 21097 15997 21131 16031
rect 21131 15997 21140 16031
rect 21088 15988 21140 15997
rect 21180 15988 21232 16040
rect 21640 16099 21692 16108
rect 21640 16065 21649 16099
rect 21649 16065 21683 16099
rect 21683 16065 21692 16099
rect 21640 16056 21692 16065
rect 17776 15963 17828 15972
rect 17776 15929 17785 15963
rect 17785 15929 17819 15963
rect 17819 15929 17828 15963
rect 17776 15920 17828 15929
rect 13360 15852 13412 15904
rect 21088 15852 21140 15904
rect 21732 16031 21784 16040
rect 21732 15997 21741 16031
rect 21741 15997 21775 16031
rect 21775 15997 21784 16031
rect 21732 15988 21784 15997
rect 21824 15988 21876 16040
rect 23572 16099 23624 16108
rect 23572 16065 23581 16099
rect 23581 16065 23615 16099
rect 23615 16065 23624 16099
rect 23572 16056 23624 16065
rect 22284 15920 22336 15972
rect 22652 15963 22704 15972
rect 22652 15929 22661 15963
rect 22661 15929 22695 15963
rect 22695 15929 22704 15963
rect 22652 15920 22704 15929
rect 24216 15988 24268 16040
rect 24860 16056 24912 16108
rect 24492 16031 24544 16040
rect 24492 15997 24501 16031
rect 24501 15997 24535 16031
rect 24535 15997 24544 16031
rect 24492 15988 24544 15997
rect 24584 16031 24636 16040
rect 24584 15997 24593 16031
rect 24593 15997 24627 16031
rect 24627 15997 24636 16031
rect 24584 15988 24636 15997
rect 24676 16031 24728 16040
rect 24676 15997 24685 16031
rect 24685 15997 24719 16031
rect 24719 15997 24728 16031
rect 24676 15988 24728 15997
rect 25688 15988 25740 16040
rect 24400 15852 24452 15904
rect 26240 15852 26292 15904
rect 7114 15750 7166 15802
rect 7178 15750 7230 15802
rect 7242 15750 7294 15802
rect 7306 15750 7358 15802
rect 7370 15750 7422 15802
rect 13830 15750 13882 15802
rect 13894 15750 13946 15802
rect 13958 15750 14010 15802
rect 14022 15750 14074 15802
rect 14086 15750 14138 15802
rect 20546 15750 20598 15802
rect 20610 15750 20662 15802
rect 20674 15750 20726 15802
rect 20738 15750 20790 15802
rect 20802 15750 20854 15802
rect 27262 15750 27314 15802
rect 27326 15750 27378 15802
rect 27390 15750 27442 15802
rect 27454 15750 27506 15802
rect 27518 15750 27570 15802
rect 1492 15512 1544 15564
rect 1676 15555 1728 15564
rect 1676 15521 1685 15555
rect 1685 15521 1719 15555
rect 1719 15521 1728 15555
rect 1676 15512 1728 15521
rect 1860 15555 1912 15564
rect 1860 15521 1869 15555
rect 1869 15521 1903 15555
rect 1903 15521 1912 15555
rect 1860 15512 1912 15521
rect 3332 15691 3384 15700
rect 3332 15657 3341 15691
rect 3341 15657 3375 15691
rect 3375 15657 3384 15691
rect 3332 15648 3384 15657
rect 6460 15691 6512 15700
rect 6460 15657 6469 15691
rect 6469 15657 6503 15691
rect 6503 15657 6512 15691
rect 6460 15648 6512 15657
rect 7012 15648 7064 15700
rect 3608 15580 3660 15632
rect 6184 15580 6236 15632
rect 2596 15512 2648 15564
rect 5080 15512 5132 15564
rect 1400 15376 1452 15428
rect 1216 15351 1268 15360
rect 1216 15317 1225 15351
rect 1225 15317 1259 15351
rect 1259 15317 1268 15351
rect 1216 15308 1268 15317
rect 2596 15308 2648 15360
rect 6276 15444 6328 15496
rect 8208 15512 8260 15564
rect 10324 15648 10376 15700
rect 11428 15648 11480 15700
rect 12440 15691 12492 15700
rect 12440 15657 12449 15691
rect 12449 15657 12483 15691
rect 12483 15657 12492 15691
rect 12440 15648 12492 15657
rect 9312 15580 9364 15632
rect 14464 15648 14516 15700
rect 17684 15648 17736 15700
rect 16580 15580 16632 15632
rect 17868 15580 17920 15632
rect 20260 15648 20312 15700
rect 11244 15555 11296 15564
rect 11244 15521 11253 15555
rect 11253 15521 11287 15555
rect 11287 15521 11296 15555
rect 11244 15512 11296 15521
rect 9128 15444 9180 15496
rect 9220 15444 9272 15496
rect 11336 15444 11388 15496
rect 12440 15512 12492 15564
rect 12624 15555 12676 15564
rect 12624 15521 12633 15555
rect 12633 15521 12667 15555
rect 12667 15521 12676 15555
rect 12624 15512 12676 15521
rect 12992 15555 13044 15564
rect 12992 15521 13001 15555
rect 13001 15521 13035 15555
rect 13035 15521 13044 15555
rect 12992 15512 13044 15521
rect 13360 15512 13412 15564
rect 13544 15555 13596 15564
rect 13544 15521 13553 15555
rect 13553 15521 13587 15555
rect 13587 15521 13596 15555
rect 13544 15512 13596 15521
rect 11520 15444 11572 15496
rect 15200 15444 15252 15496
rect 15568 15555 15620 15564
rect 15568 15521 15577 15555
rect 15577 15521 15611 15555
rect 15611 15521 15620 15555
rect 15568 15512 15620 15521
rect 16856 15555 16908 15564
rect 16856 15521 16865 15555
rect 16865 15521 16899 15555
rect 16899 15521 16908 15555
rect 16856 15512 16908 15521
rect 17040 15512 17092 15564
rect 17960 15444 18012 15496
rect 18696 15512 18748 15564
rect 22008 15648 22060 15700
rect 22652 15648 22704 15700
rect 23204 15648 23256 15700
rect 24492 15648 24544 15700
rect 19248 15555 19300 15564
rect 19248 15521 19257 15555
rect 19257 15521 19291 15555
rect 19291 15521 19300 15555
rect 19248 15512 19300 15521
rect 19340 15512 19392 15564
rect 21088 15512 21140 15564
rect 21824 15623 21876 15632
rect 21824 15589 21833 15623
rect 21833 15589 21867 15623
rect 21867 15589 21876 15623
rect 21824 15580 21876 15589
rect 22100 15623 22152 15632
rect 22100 15589 22109 15623
rect 22109 15589 22143 15623
rect 22143 15589 22152 15623
rect 22100 15580 22152 15589
rect 22744 15580 22796 15632
rect 22468 15512 22520 15564
rect 24400 15555 24452 15564
rect 24400 15521 24409 15555
rect 24409 15521 24443 15555
rect 24443 15521 24452 15555
rect 24400 15512 24452 15521
rect 24584 15555 24636 15564
rect 24584 15521 24593 15555
rect 24593 15521 24627 15555
rect 24627 15521 24636 15555
rect 24584 15512 24636 15521
rect 24676 15512 24728 15564
rect 21180 15444 21232 15496
rect 4528 15308 4580 15360
rect 4804 15308 4856 15360
rect 5172 15308 5224 15360
rect 5816 15308 5868 15360
rect 6276 15308 6328 15360
rect 17592 15376 17644 15428
rect 21732 15444 21784 15496
rect 23664 15444 23716 15496
rect 22928 15376 22980 15428
rect 24952 15512 25004 15564
rect 26608 15512 26660 15564
rect 26240 15487 26292 15496
rect 26240 15453 26249 15487
rect 26249 15453 26283 15487
rect 26283 15453 26292 15487
rect 26240 15444 26292 15453
rect 26976 15487 27028 15496
rect 26976 15453 26985 15487
rect 26985 15453 27019 15487
rect 27019 15453 27028 15487
rect 26976 15444 27028 15453
rect 26792 15376 26844 15428
rect 7196 15351 7248 15360
rect 7196 15317 7205 15351
rect 7205 15317 7239 15351
rect 7239 15317 7248 15351
rect 7196 15308 7248 15317
rect 7748 15308 7800 15360
rect 8484 15351 8536 15360
rect 8484 15317 8493 15351
rect 8493 15317 8527 15351
rect 8527 15317 8536 15351
rect 8484 15308 8536 15317
rect 8760 15308 8812 15360
rect 16672 15308 16724 15360
rect 17040 15308 17092 15360
rect 18880 15308 18932 15360
rect 22008 15308 22060 15360
rect 22560 15351 22612 15360
rect 22560 15317 22569 15351
rect 22569 15317 22603 15351
rect 22603 15317 22612 15351
rect 22560 15308 22612 15317
rect 26700 15308 26752 15360
rect 3756 15206 3808 15258
rect 3820 15206 3872 15258
rect 3884 15206 3936 15258
rect 3948 15206 4000 15258
rect 4012 15206 4064 15258
rect 10472 15206 10524 15258
rect 10536 15206 10588 15258
rect 10600 15206 10652 15258
rect 10664 15206 10716 15258
rect 10728 15206 10780 15258
rect 17188 15206 17240 15258
rect 17252 15206 17304 15258
rect 17316 15206 17368 15258
rect 17380 15206 17432 15258
rect 17444 15206 17496 15258
rect 23904 15206 23956 15258
rect 23968 15206 24020 15258
rect 24032 15206 24084 15258
rect 24096 15206 24148 15258
rect 24160 15206 24212 15258
rect 2504 15104 2556 15156
rect 3608 15104 3660 15156
rect 6920 15104 6972 15156
rect 7196 15104 7248 15156
rect 8116 15104 8168 15156
rect 12992 15104 13044 15156
rect 21824 15104 21876 15156
rect 23664 15147 23716 15156
rect 23664 15113 23673 15147
rect 23673 15113 23707 15147
rect 23707 15113 23716 15147
rect 23664 15104 23716 15113
rect 26332 15104 26384 15156
rect 26976 15104 27028 15156
rect 4160 14968 4212 15020
rect 1400 14900 1452 14952
rect 4620 15011 4672 15020
rect 4620 14977 4629 15011
rect 4629 14977 4663 15011
rect 4663 14977 4672 15011
rect 4620 14968 4672 14977
rect 4712 15011 4764 15020
rect 4712 14977 4721 15011
rect 4721 14977 4755 15011
rect 4755 14977 4764 15011
rect 4712 14968 4764 14977
rect 14832 15036 14884 15088
rect 1216 14832 1268 14884
rect 4528 14900 4580 14952
rect 6092 14900 6144 14952
rect 6552 14943 6604 14952
rect 6552 14909 6586 14943
rect 6586 14909 6604 14943
rect 6552 14900 6604 14909
rect 7748 14943 7800 14952
rect 7748 14909 7757 14943
rect 7757 14909 7791 14943
rect 7791 14909 7800 14943
rect 7748 14900 7800 14909
rect 7932 14943 7984 14952
rect 7932 14909 7941 14943
rect 7941 14909 7975 14943
rect 7975 14909 7984 14943
rect 7932 14900 7984 14909
rect 8392 14943 8444 14952
rect 8392 14909 8401 14943
rect 8401 14909 8435 14943
rect 8435 14909 8444 14943
rect 8392 14900 8444 14909
rect 9588 14900 9640 14952
rect 11152 14900 11204 14952
rect 12348 14968 12400 15020
rect 5172 14832 5224 14884
rect 6184 14832 6236 14884
rect 8484 14832 8536 14884
rect 12164 14832 12216 14884
rect 12624 14943 12676 14952
rect 12624 14909 12633 14943
rect 12633 14909 12667 14943
rect 12667 14909 12676 14943
rect 12624 14900 12676 14909
rect 13636 14968 13688 15020
rect 14188 14900 14240 14952
rect 14280 14900 14332 14952
rect 7748 14764 7800 14816
rect 9588 14764 9640 14816
rect 11704 14764 11756 14816
rect 13544 14832 13596 14884
rect 14832 14832 14884 14884
rect 15200 14832 15252 14884
rect 16212 14900 16264 14952
rect 21916 14968 21968 15020
rect 25044 14968 25096 15020
rect 25688 15011 25740 15020
rect 25688 14977 25697 15011
rect 25697 14977 25731 15011
rect 25731 14977 25740 15011
rect 25688 14968 25740 14977
rect 16856 14832 16908 14884
rect 12900 14764 12952 14816
rect 17960 14900 18012 14952
rect 22100 14900 22152 14952
rect 22836 14900 22888 14952
rect 21088 14832 21140 14884
rect 22560 14875 22612 14884
rect 22560 14841 22594 14875
rect 22594 14841 22612 14875
rect 22560 14832 22612 14841
rect 23296 14832 23348 14884
rect 24952 14875 25004 14884
rect 24952 14841 24961 14875
rect 24961 14841 24995 14875
rect 24995 14841 25004 14875
rect 24952 14832 25004 14841
rect 26424 14832 26476 14884
rect 17500 14764 17552 14816
rect 17960 14764 18012 14816
rect 23388 14764 23440 14816
rect 26884 14764 26936 14816
rect 7114 14662 7166 14714
rect 7178 14662 7230 14714
rect 7242 14662 7294 14714
rect 7306 14662 7358 14714
rect 7370 14662 7422 14714
rect 13830 14662 13882 14714
rect 13894 14662 13946 14714
rect 13958 14662 14010 14714
rect 14022 14662 14074 14714
rect 14086 14662 14138 14714
rect 20546 14662 20598 14714
rect 20610 14662 20662 14714
rect 20674 14662 20726 14714
rect 20738 14662 20790 14714
rect 20802 14662 20854 14714
rect 27262 14662 27314 14714
rect 27326 14662 27378 14714
rect 27390 14662 27442 14714
rect 27454 14662 27506 14714
rect 27518 14662 27570 14714
rect 2044 14560 2096 14612
rect 1676 14535 1728 14544
rect 1676 14501 1685 14535
rect 1685 14501 1719 14535
rect 1719 14501 1728 14535
rect 1676 14492 1728 14501
rect 3332 14560 3384 14612
rect 9496 14560 9548 14612
rect 16856 14603 16908 14612
rect 16856 14569 16865 14603
rect 16865 14569 16899 14603
rect 16899 14569 16908 14603
rect 16856 14560 16908 14569
rect 5080 14535 5132 14544
rect 5080 14501 5089 14535
rect 5089 14501 5123 14535
rect 5123 14501 5132 14535
rect 5080 14492 5132 14501
rect 1584 14220 1636 14272
rect 3148 14467 3200 14476
rect 3148 14433 3157 14467
rect 3157 14433 3191 14467
rect 3191 14433 3200 14467
rect 3148 14424 3200 14433
rect 3332 14467 3384 14476
rect 3332 14433 3341 14467
rect 3341 14433 3375 14467
rect 3375 14433 3384 14467
rect 3332 14424 3384 14433
rect 4804 14467 4856 14476
rect 4804 14433 4813 14467
rect 4813 14433 4847 14467
rect 4847 14433 4856 14467
rect 4804 14424 4856 14433
rect 5448 14424 5500 14476
rect 4528 14399 4580 14408
rect 4528 14365 4537 14399
rect 4537 14365 4571 14399
rect 4571 14365 4580 14399
rect 4528 14356 4580 14365
rect 7932 14492 7984 14544
rect 11336 14535 11388 14544
rect 11336 14501 11345 14535
rect 11345 14501 11379 14535
rect 11379 14501 11388 14535
rect 11336 14492 11388 14501
rect 15568 14492 15620 14544
rect 17500 14535 17552 14544
rect 17500 14501 17509 14535
rect 17509 14501 17543 14535
rect 17543 14501 17552 14535
rect 17500 14492 17552 14501
rect 22100 14535 22152 14544
rect 7656 14424 7708 14476
rect 7748 14467 7800 14476
rect 7748 14433 7757 14467
rect 7757 14433 7791 14467
rect 7791 14433 7800 14467
rect 7748 14424 7800 14433
rect 8208 14424 8260 14476
rect 7472 14356 7524 14408
rect 8760 14399 8812 14408
rect 8760 14365 8769 14399
rect 8769 14365 8803 14399
rect 8803 14365 8812 14399
rect 8760 14356 8812 14365
rect 9588 14467 9640 14476
rect 9588 14433 9597 14467
rect 9597 14433 9631 14467
rect 9631 14433 9640 14467
rect 9588 14424 9640 14433
rect 11244 14424 11296 14476
rect 11704 14467 11756 14476
rect 11704 14433 11713 14467
rect 11713 14433 11747 14467
rect 11747 14433 11756 14467
rect 11704 14424 11756 14433
rect 11888 14424 11940 14476
rect 12072 14467 12124 14476
rect 12072 14433 12106 14467
rect 12106 14433 12124 14467
rect 12072 14424 12124 14433
rect 14556 14467 14608 14476
rect 14556 14433 14590 14467
rect 14590 14433 14608 14467
rect 14556 14424 14608 14433
rect 17040 14467 17092 14476
rect 17040 14433 17049 14467
rect 17049 14433 17083 14467
rect 17083 14433 17092 14467
rect 17040 14424 17092 14433
rect 17960 14424 18012 14476
rect 18144 14424 18196 14476
rect 22100 14501 22109 14535
rect 22109 14501 22143 14535
rect 22143 14501 22152 14535
rect 22100 14492 22152 14501
rect 23020 14492 23072 14544
rect 2228 14220 2280 14272
rect 2964 14220 3016 14272
rect 5908 14220 5960 14272
rect 6184 14263 6236 14272
rect 6184 14229 6193 14263
rect 6193 14229 6227 14263
rect 6227 14229 6236 14263
rect 6184 14220 6236 14229
rect 6276 14220 6328 14272
rect 7012 14288 7064 14340
rect 9220 14331 9272 14340
rect 9220 14297 9229 14331
rect 9229 14297 9263 14331
rect 9263 14297 9272 14331
rect 9220 14288 9272 14297
rect 14280 14399 14332 14408
rect 14280 14365 14289 14399
rect 14289 14365 14323 14399
rect 14323 14365 14332 14399
rect 14280 14356 14332 14365
rect 16304 14356 16356 14408
rect 21088 14424 21140 14476
rect 21272 14467 21324 14476
rect 21272 14433 21281 14467
rect 21281 14433 21315 14467
rect 21315 14433 21324 14467
rect 21272 14424 21324 14433
rect 21732 14356 21784 14408
rect 22652 14424 22704 14476
rect 23296 14467 23348 14476
rect 23296 14433 23305 14467
rect 23305 14433 23339 14467
rect 23339 14433 23348 14467
rect 23296 14424 23348 14433
rect 23756 14560 23808 14612
rect 25044 14603 25096 14612
rect 25044 14569 25053 14603
rect 25053 14569 25087 14603
rect 25087 14569 25096 14603
rect 25044 14560 25096 14569
rect 25688 14492 25740 14544
rect 26608 14424 26660 14476
rect 23480 14356 23532 14408
rect 22008 14288 22060 14340
rect 23572 14288 23624 14340
rect 6920 14220 6972 14272
rect 13176 14263 13228 14272
rect 13176 14229 13185 14263
rect 13185 14229 13219 14263
rect 13219 14229 13228 14263
rect 13176 14220 13228 14229
rect 13268 14263 13320 14272
rect 13268 14229 13277 14263
rect 13277 14229 13311 14263
rect 13311 14229 13320 14263
rect 13268 14220 13320 14229
rect 13452 14220 13504 14272
rect 15016 14220 15068 14272
rect 16120 14263 16172 14272
rect 16120 14229 16129 14263
rect 16129 14229 16163 14263
rect 16163 14229 16172 14263
rect 16120 14220 16172 14229
rect 18696 14220 18748 14272
rect 20720 14263 20772 14272
rect 20720 14229 20729 14263
rect 20729 14229 20763 14263
rect 20763 14229 20772 14263
rect 20720 14220 20772 14229
rect 23388 14220 23440 14272
rect 24952 14356 25004 14408
rect 26884 14467 26936 14476
rect 26884 14433 26893 14467
rect 26893 14433 26927 14467
rect 26927 14433 26936 14467
rect 26884 14424 26936 14433
rect 26976 14424 27028 14476
rect 25688 14288 25740 14340
rect 25780 14220 25832 14272
rect 3756 14118 3808 14170
rect 3820 14118 3872 14170
rect 3884 14118 3936 14170
rect 3948 14118 4000 14170
rect 4012 14118 4064 14170
rect 10472 14118 10524 14170
rect 10536 14118 10588 14170
rect 10600 14118 10652 14170
rect 10664 14118 10716 14170
rect 10728 14118 10780 14170
rect 17188 14118 17240 14170
rect 17252 14118 17304 14170
rect 17316 14118 17368 14170
rect 17380 14118 17432 14170
rect 17444 14118 17496 14170
rect 23904 14118 23956 14170
rect 23968 14118 24020 14170
rect 24032 14118 24084 14170
rect 24096 14118 24148 14170
rect 24160 14118 24212 14170
rect 2228 14059 2280 14068
rect 2228 14025 2237 14059
rect 2237 14025 2271 14059
rect 2271 14025 2280 14059
rect 2228 14016 2280 14025
rect 1400 13812 1452 13864
rect 3148 14016 3200 14068
rect 10876 14016 10928 14068
rect 8484 13948 8536 14000
rect 10048 13948 10100 14000
rect 3424 13812 3476 13864
rect 4528 13812 4580 13864
rect 5172 13812 5224 13864
rect 5448 13812 5500 13864
rect 6552 13855 6604 13864
rect 6552 13821 6561 13855
rect 6561 13821 6595 13855
rect 6595 13821 6604 13855
rect 6552 13812 6604 13821
rect 6644 13812 6696 13864
rect 6828 13812 6880 13864
rect 8116 13812 8168 13864
rect 10968 13812 11020 13864
rect 12072 14016 12124 14068
rect 13268 14016 13320 14068
rect 14464 14016 14516 14068
rect 14556 14016 14608 14068
rect 15016 14016 15068 14068
rect 15108 13948 15160 14000
rect 16120 14016 16172 14068
rect 18144 14016 18196 14068
rect 1308 13744 1360 13796
rect 4160 13744 4212 13796
rect 4712 13744 4764 13796
rect 10324 13744 10376 13796
rect 1768 13676 1820 13728
rect 3884 13676 3936 13728
rect 4620 13676 4672 13728
rect 6736 13676 6788 13728
rect 7932 13676 7984 13728
rect 8944 13719 8996 13728
rect 8944 13685 8953 13719
rect 8953 13685 8987 13719
rect 8987 13685 8996 13719
rect 8944 13676 8996 13685
rect 9956 13676 10008 13728
rect 12624 13855 12676 13864
rect 12624 13821 12633 13855
rect 12633 13821 12667 13855
rect 12667 13821 12676 13855
rect 12624 13812 12676 13821
rect 11520 13787 11572 13796
rect 11520 13753 11529 13787
rect 11529 13753 11563 13787
rect 11563 13753 11572 13787
rect 11520 13744 11572 13753
rect 12164 13744 12216 13796
rect 12992 13744 13044 13796
rect 13360 13855 13412 13864
rect 13360 13821 13369 13855
rect 13369 13821 13403 13855
rect 13403 13821 13412 13855
rect 13360 13812 13412 13821
rect 14188 13880 14240 13932
rect 14280 13880 14332 13932
rect 14648 13880 14700 13932
rect 13728 13855 13780 13864
rect 13728 13821 13737 13855
rect 13737 13821 13771 13855
rect 13771 13821 13780 13855
rect 13728 13812 13780 13821
rect 15108 13812 15160 13864
rect 16764 13855 16816 13864
rect 16764 13821 16773 13855
rect 16773 13821 16807 13855
rect 16807 13821 16816 13855
rect 16764 13812 16816 13821
rect 18604 13948 18656 14000
rect 19524 13948 19576 14000
rect 21364 14016 21416 14068
rect 21732 14059 21784 14068
rect 21732 14025 21741 14059
rect 21741 14025 21775 14059
rect 21775 14025 21784 14059
rect 21732 14016 21784 14025
rect 20996 13948 21048 14000
rect 21088 13948 21140 14000
rect 14556 13744 14608 13796
rect 17592 13812 17644 13864
rect 18052 13744 18104 13796
rect 18512 13855 18564 13864
rect 18512 13821 18521 13855
rect 18521 13821 18555 13855
rect 18555 13821 18564 13855
rect 18512 13812 18564 13821
rect 18696 13855 18748 13864
rect 18696 13821 18705 13855
rect 18705 13821 18739 13855
rect 18739 13821 18748 13855
rect 18696 13812 18748 13821
rect 18972 13812 19024 13864
rect 20352 13855 20404 13864
rect 20352 13821 20361 13855
rect 20361 13821 20395 13855
rect 20395 13821 20404 13855
rect 20352 13812 20404 13821
rect 20720 13880 20772 13932
rect 22100 14016 22152 14068
rect 23204 13991 23256 14000
rect 23204 13957 23213 13991
rect 23213 13957 23247 13991
rect 23247 13957 23256 13991
rect 23204 13948 23256 13957
rect 19064 13744 19116 13796
rect 21916 13812 21968 13864
rect 23388 13812 23440 13864
rect 23756 13812 23808 13864
rect 24860 13855 24912 13864
rect 24860 13821 24869 13855
rect 24869 13821 24903 13855
rect 24903 13821 24912 13855
rect 24860 13812 24912 13821
rect 25044 13855 25096 13864
rect 25044 13821 25053 13855
rect 25053 13821 25087 13855
rect 25087 13821 25096 13855
rect 25044 13812 25096 13821
rect 25596 13812 25648 13864
rect 25780 13855 25832 13864
rect 25780 13821 25814 13855
rect 25814 13821 25832 13855
rect 25780 13812 25832 13821
rect 21272 13744 21324 13796
rect 22192 13744 22244 13796
rect 24400 13744 24452 13796
rect 11888 13676 11940 13728
rect 12440 13676 12492 13728
rect 12900 13719 12952 13728
rect 12900 13685 12927 13719
rect 12927 13685 12952 13719
rect 12900 13676 12952 13685
rect 15016 13676 15068 13728
rect 15200 13676 15252 13728
rect 16212 13719 16264 13728
rect 16212 13685 16221 13719
rect 16221 13685 16255 13719
rect 16255 13685 16264 13719
rect 16212 13676 16264 13685
rect 16948 13719 17000 13728
rect 16948 13685 16957 13719
rect 16957 13685 16991 13719
rect 16991 13685 17000 13719
rect 16948 13676 17000 13685
rect 18880 13676 18932 13728
rect 23296 13719 23348 13728
rect 23296 13685 23305 13719
rect 23305 13685 23339 13719
rect 23339 13685 23348 13719
rect 23296 13676 23348 13685
rect 23572 13676 23624 13728
rect 24584 13719 24636 13728
rect 24584 13685 24593 13719
rect 24593 13685 24627 13719
rect 24627 13685 24636 13719
rect 24584 13676 24636 13685
rect 26884 13719 26936 13728
rect 26884 13685 26893 13719
rect 26893 13685 26927 13719
rect 26927 13685 26936 13719
rect 26884 13676 26936 13685
rect 7114 13574 7166 13626
rect 7178 13574 7230 13626
rect 7242 13574 7294 13626
rect 7306 13574 7358 13626
rect 7370 13574 7422 13626
rect 13830 13574 13882 13626
rect 13894 13574 13946 13626
rect 13958 13574 14010 13626
rect 14022 13574 14074 13626
rect 14086 13574 14138 13626
rect 20546 13574 20598 13626
rect 20610 13574 20662 13626
rect 20674 13574 20726 13626
rect 20738 13574 20790 13626
rect 20802 13574 20854 13626
rect 27262 13574 27314 13626
rect 27326 13574 27378 13626
rect 27390 13574 27442 13626
rect 27454 13574 27506 13626
rect 27518 13574 27570 13626
rect 1308 13515 1360 13524
rect 1308 13481 1317 13515
rect 1317 13481 1351 13515
rect 1351 13481 1360 13515
rect 1308 13472 1360 13481
rect 3332 13515 3384 13524
rect 3332 13481 3341 13515
rect 3341 13481 3375 13515
rect 3375 13481 3384 13515
rect 3332 13472 3384 13481
rect 4160 13472 4212 13524
rect 6552 13472 6604 13524
rect 6920 13404 6972 13456
rect 12440 13472 12492 13524
rect 13452 13472 13504 13524
rect 14372 13515 14424 13524
rect 14372 13481 14399 13515
rect 14399 13481 14424 13515
rect 14372 13472 14424 13481
rect 15108 13472 15160 13524
rect 18052 13472 18104 13524
rect 18880 13515 18932 13524
rect 18880 13481 18907 13515
rect 18907 13481 18932 13515
rect 18880 13472 18932 13481
rect 3148 13379 3200 13388
rect 3148 13345 3157 13379
rect 3157 13345 3191 13379
rect 3191 13345 3200 13379
rect 3148 13336 3200 13345
rect 3424 13379 3476 13388
rect 3424 13345 3433 13379
rect 3433 13345 3467 13379
rect 3467 13345 3476 13379
rect 3424 13336 3476 13345
rect 1860 13311 1912 13320
rect 1860 13277 1869 13311
rect 1869 13277 1903 13311
rect 1903 13277 1912 13311
rect 1860 13268 1912 13277
rect 3884 13379 3936 13388
rect 3884 13345 3893 13379
rect 3893 13345 3927 13379
rect 3927 13345 3936 13379
rect 3884 13336 3936 13345
rect 6184 13336 6236 13388
rect 6276 13379 6328 13388
rect 6276 13345 6285 13379
rect 6285 13345 6319 13379
rect 6319 13345 6328 13379
rect 6276 13336 6328 13345
rect 6368 13379 6420 13388
rect 6368 13345 6377 13379
rect 6377 13345 6411 13379
rect 6411 13345 6420 13379
rect 6368 13336 6420 13345
rect 6736 13379 6788 13388
rect 6736 13345 6770 13379
rect 6770 13345 6788 13379
rect 6736 13336 6788 13345
rect 8392 13404 8444 13456
rect 13360 13404 13412 13456
rect 14188 13404 14240 13456
rect 14556 13447 14608 13456
rect 14556 13413 14565 13447
rect 14565 13413 14599 13447
rect 14599 13413 14608 13447
rect 14556 13404 14608 13413
rect 16212 13404 16264 13456
rect 16948 13404 17000 13456
rect 19064 13447 19116 13456
rect 19064 13413 19073 13447
rect 19073 13413 19107 13447
rect 19107 13413 19116 13447
rect 19064 13404 19116 13413
rect 21272 13515 21324 13524
rect 21272 13481 21281 13515
rect 21281 13481 21315 13515
rect 21315 13481 21324 13515
rect 21272 13472 21324 13481
rect 22192 13472 22244 13524
rect 9588 13379 9640 13388
rect 9588 13345 9597 13379
rect 9597 13345 9631 13379
rect 9631 13345 9640 13379
rect 9588 13336 9640 13345
rect 9864 13379 9916 13388
rect 9864 13345 9873 13379
rect 9873 13345 9907 13379
rect 9907 13345 9916 13379
rect 9864 13336 9916 13345
rect 9956 13379 10008 13388
rect 9956 13345 9965 13379
rect 9965 13345 9999 13379
rect 9999 13345 10008 13379
rect 9956 13336 10008 13345
rect 10876 13336 10928 13388
rect 11520 13336 11572 13388
rect 15660 13379 15712 13388
rect 15660 13345 15669 13379
rect 15669 13345 15703 13379
rect 15703 13345 15712 13379
rect 15660 13336 15712 13345
rect 16028 13336 16080 13388
rect 2320 13243 2372 13252
rect 2320 13209 2329 13243
rect 2329 13209 2363 13243
rect 2363 13209 2372 13243
rect 2320 13200 2372 13209
rect 2688 13175 2740 13184
rect 2688 13141 2697 13175
rect 2697 13141 2731 13175
rect 2731 13141 2740 13175
rect 2688 13132 2740 13141
rect 5816 13268 5868 13320
rect 6092 13311 6144 13320
rect 6092 13277 6101 13311
rect 6101 13277 6135 13311
rect 6135 13277 6144 13311
rect 6092 13268 6144 13277
rect 5356 13200 5408 13252
rect 13084 13268 13136 13320
rect 15384 13311 15436 13320
rect 15384 13277 15393 13311
rect 15393 13277 15427 13311
rect 15427 13277 15436 13311
rect 15384 13268 15436 13277
rect 16396 13311 16448 13320
rect 16396 13277 16405 13311
rect 16405 13277 16439 13311
rect 16439 13277 16448 13311
rect 16396 13268 16448 13277
rect 8944 13200 8996 13252
rect 15568 13200 15620 13252
rect 17684 13200 17736 13252
rect 20996 13379 21048 13388
rect 20996 13345 21005 13379
rect 21005 13345 21039 13379
rect 21039 13345 21048 13379
rect 20996 13336 21048 13345
rect 21456 13379 21508 13388
rect 21456 13345 21465 13379
rect 21465 13345 21499 13379
rect 21499 13345 21508 13379
rect 21456 13336 21508 13345
rect 21548 13379 21600 13388
rect 21548 13345 21557 13379
rect 21557 13345 21591 13379
rect 21591 13345 21600 13379
rect 21548 13336 21600 13345
rect 22744 13404 22796 13456
rect 22468 13336 22520 13388
rect 4528 13132 4580 13184
rect 5448 13132 5500 13184
rect 9312 13175 9364 13184
rect 9312 13141 9321 13175
rect 9321 13141 9355 13175
rect 9355 13141 9364 13175
rect 9312 13132 9364 13141
rect 10876 13132 10928 13184
rect 11336 13132 11388 13184
rect 12808 13132 12860 13184
rect 14280 13132 14332 13184
rect 15476 13175 15528 13184
rect 15476 13141 15485 13175
rect 15485 13141 15519 13175
rect 15519 13141 15528 13175
rect 15476 13132 15528 13141
rect 17592 13132 17644 13184
rect 20720 13311 20772 13320
rect 20720 13277 20729 13311
rect 20729 13277 20763 13311
rect 20763 13277 20772 13311
rect 20720 13268 20772 13277
rect 22100 13268 22152 13320
rect 19340 13243 19392 13252
rect 19340 13209 19349 13243
rect 19349 13209 19383 13243
rect 19383 13209 19392 13243
rect 19340 13200 19392 13209
rect 25412 13472 25464 13524
rect 26608 13472 26660 13524
rect 23572 13404 23624 13456
rect 23020 13200 23072 13252
rect 23296 13336 23348 13388
rect 24952 13404 25004 13456
rect 25688 13404 25740 13456
rect 23296 13200 23348 13252
rect 23388 13200 23440 13252
rect 26608 13336 26660 13388
rect 26884 13336 26936 13388
rect 24860 13311 24912 13320
rect 24860 13277 24869 13311
rect 24869 13277 24903 13311
rect 24903 13277 24912 13311
rect 24860 13268 24912 13277
rect 27068 13268 27120 13320
rect 24308 13132 24360 13184
rect 24952 13175 25004 13184
rect 24952 13141 24961 13175
rect 24961 13141 24995 13175
rect 24995 13141 25004 13175
rect 24952 13132 25004 13141
rect 25044 13132 25096 13184
rect 26240 13132 26292 13184
rect 3756 13030 3808 13082
rect 3820 13030 3872 13082
rect 3884 13030 3936 13082
rect 3948 13030 4000 13082
rect 4012 13030 4064 13082
rect 10472 13030 10524 13082
rect 10536 13030 10588 13082
rect 10600 13030 10652 13082
rect 10664 13030 10716 13082
rect 10728 13030 10780 13082
rect 17188 13030 17240 13082
rect 17252 13030 17304 13082
rect 17316 13030 17368 13082
rect 17380 13030 17432 13082
rect 17444 13030 17496 13082
rect 23904 13030 23956 13082
rect 23968 13030 24020 13082
rect 24032 13030 24084 13082
rect 24096 13030 24148 13082
rect 24160 13030 24212 13082
rect 1860 12928 1912 12980
rect 4528 12928 4580 12980
rect 1676 12860 1728 12912
rect 2044 12860 2096 12912
rect 2964 12860 3016 12912
rect 1768 12835 1820 12844
rect 1768 12801 1777 12835
rect 1777 12801 1811 12835
rect 1811 12801 1820 12835
rect 1768 12792 1820 12801
rect 1860 12835 1912 12844
rect 1860 12801 1869 12835
rect 1869 12801 1903 12835
rect 1903 12801 1912 12835
rect 1860 12792 1912 12801
rect 1584 12767 1636 12776
rect 1584 12733 1593 12767
rect 1593 12733 1627 12767
rect 1627 12733 1636 12767
rect 1584 12724 1636 12733
rect 2320 12724 2372 12776
rect 2780 12767 2832 12776
rect 2780 12733 2789 12767
rect 2789 12733 2823 12767
rect 2823 12733 2832 12767
rect 2780 12724 2832 12733
rect 3700 12860 3752 12912
rect 5172 12928 5224 12980
rect 4528 12835 4580 12844
rect 4528 12801 4537 12835
rect 4537 12801 4571 12835
rect 4571 12801 4580 12835
rect 4528 12792 4580 12801
rect 5448 12860 5500 12912
rect 6828 12928 6880 12980
rect 10324 12928 10376 12980
rect 10876 12928 10928 12980
rect 12164 12928 12216 12980
rect 12624 12928 12676 12980
rect 12808 12971 12860 12980
rect 12808 12937 12817 12971
rect 12817 12937 12851 12971
rect 12851 12937 12860 12971
rect 12808 12928 12860 12937
rect 15568 12928 15620 12980
rect 9588 12860 9640 12912
rect 9680 12860 9732 12912
rect 10048 12860 10100 12912
rect 10784 12860 10836 12912
rect 13084 12860 13136 12912
rect 16764 12928 16816 12980
rect 17040 12928 17092 12980
rect 20352 12971 20404 12980
rect 20352 12937 20361 12971
rect 20361 12937 20395 12971
rect 20395 12937 20404 12971
rect 20352 12928 20404 12937
rect 2872 12656 2924 12708
rect 4344 12767 4396 12776
rect 4344 12733 4353 12767
rect 4353 12733 4387 12767
rect 4387 12733 4396 12767
rect 4344 12724 4396 12733
rect 3608 12699 3660 12708
rect 3608 12665 3617 12699
rect 3617 12665 3651 12699
rect 3651 12665 3660 12699
rect 4712 12724 4764 12776
rect 4804 12699 4856 12708
rect 3608 12656 3660 12665
rect 2228 12588 2280 12640
rect 2596 12631 2648 12640
rect 2596 12597 2605 12631
rect 2605 12597 2639 12631
rect 2639 12597 2648 12631
rect 2596 12588 2648 12597
rect 3240 12631 3292 12640
rect 3240 12597 3249 12631
rect 3249 12597 3283 12631
rect 3283 12597 3292 12631
rect 3240 12588 3292 12597
rect 4252 12588 4304 12640
rect 4804 12665 4813 12699
rect 4813 12665 4847 12699
rect 4847 12665 4856 12699
rect 4804 12656 4856 12665
rect 6368 12767 6420 12776
rect 6368 12733 6377 12767
rect 6377 12733 6411 12767
rect 6411 12733 6420 12767
rect 6368 12724 6420 12733
rect 6552 12767 6604 12776
rect 6552 12733 6561 12767
rect 6561 12733 6595 12767
rect 6595 12733 6604 12767
rect 6552 12724 6604 12733
rect 8944 12792 8996 12844
rect 9312 12792 9364 12844
rect 9496 12792 9548 12844
rect 9864 12792 9916 12844
rect 8852 12656 8904 12708
rect 9680 12656 9732 12708
rect 6000 12588 6052 12640
rect 6184 12588 6236 12640
rect 9772 12588 9824 12640
rect 10324 12588 10376 12640
rect 10784 12656 10836 12708
rect 11888 12724 11940 12776
rect 13084 12767 13136 12776
rect 13084 12733 13093 12767
rect 13093 12733 13127 12767
rect 13127 12733 13136 12767
rect 13084 12724 13136 12733
rect 13452 12724 13504 12776
rect 16396 12792 16448 12844
rect 20720 12835 20772 12844
rect 20720 12801 20729 12835
rect 20729 12801 20763 12835
rect 20763 12801 20772 12835
rect 20720 12792 20772 12801
rect 22836 12971 22888 12980
rect 22836 12937 22845 12971
rect 22845 12937 22879 12971
rect 22879 12937 22888 12971
rect 22836 12928 22888 12937
rect 23020 12928 23072 12980
rect 24860 12928 24912 12980
rect 27068 12971 27120 12980
rect 27068 12937 27077 12971
rect 27077 12937 27111 12971
rect 27111 12937 27120 12971
rect 27068 12928 27120 12937
rect 14648 12724 14700 12776
rect 17592 12767 17644 12776
rect 17592 12733 17601 12767
rect 17601 12733 17635 12767
rect 17635 12733 17644 12767
rect 17592 12724 17644 12733
rect 17684 12767 17736 12776
rect 17684 12733 17693 12767
rect 17693 12733 17727 12767
rect 17727 12733 17736 12767
rect 17684 12724 17736 12733
rect 18604 12724 18656 12776
rect 19340 12724 19392 12776
rect 21456 12724 21508 12776
rect 21824 12724 21876 12776
rect 22652 12792 22704 12844
rect 23296 12792 23348 12844
rect 23756 12860 23808 12912
rect 25596 12792 25648 12844
rect 11520 12656 11572 12708
rect 12440 12656 12492 12708
rect 12900 12656 12952 12708
rect 12992 12699 13044 12708
rect 12992 12665 13001 12699
rect 13001 12665 13035 12699
rect 13035 12665 13044 12699
rect 12992 12656 13044 12665
rect 14188 12656 14240 12708
rect 15476 12699 15528 12708
rect 15476 12665 15510 12699
rect 15510 12665 15528 12699
rect 15476 12656 15528 12665
rect 10968 12588 11020 12640
rect 11336 12588 11388 12640
rect 11704 12588 11756 12640
rect 13084 12588 13136 12640
rect 15384 12588 15436 12640
rect 16120 12656 16172 12708
rect 17960 12699 18012 12708
rect 17960 12665 17969 12699
rect 17969 12665 18003 12699
rect 18003 12665 18012 12699
rect 17960 12656 18012 12665
rect 19248 12656 19300 12708
rect 24952 12767 25004 12776
rect 24952 12733 24970 12767
rect 24970 12733 25004 12767
rect 24952 12724 25004 12733
rect 22744 12656 22796 12708
rect 26240 12724 26292 12776
rect 25228 12656 25280 12708
rect 15844 12588 15896 12640
rect 20076 12631 20128 12640
rect 20076 12597 20085 12631
rect 20085 12597 20119 12631
rect 20119 12597 20128 12631
rect 20076 12588 20128 12597
rect 22652 12631 22704 12640
rect 22652 12597 22661 12631
rect 22661 12597 22695 12631
rect 22695 12597 22704 12631
rect 22652 12588 22704 12597
rect 23296 12588 23348 12640
rect 26056 12588 26108 12640
rect 7114 12486 7166 12538
rect 7178 12486 7230 12538
rect 7242 12486 7294 12538
rect 7306 12486 7358 12538
rect 7370 12486 7422 12538
rect 13830 12486 13882 12538
rect 13894 12486 13946 12538
rect 13958 12486 14010 12538
rect 14022 12486 14074 12538
rect 14086 12486 14138 12538
rect 20546 12486 20598 12538
rect 20610 12486 20662 12538
rect 20674 12486 20726 12538
rect 20738 12486 20790 12538
rect 20802 12486 20854 12538
rect 27262 12486 27314 12538
rect 27326 12486 27378 12538
rect 27390 12486 27442 12538
rect 27454 12486 27506 12538
rect 27518 12486 27570 12538
rect 2136 12384 2188 12436
rect 1400 12316 1452 12368
rect 2596 12359 2648 12368
rect 1124 12291 1176 12300
rect 1124 12257 1158 12291
rect 1158 12257 1176 12291
rect 1124 12248 1176 12257
rect 2596 12325 2630 12359
rect 2630 12325 2648 12359
rect 2596 12316 2648 12325
rect 3700 12427 3752 12436
rect 3700 12393 3709 12427
rect 3709 12393 3743 12427
rect 3743 12393 3752 12427
rect 3700 12384 3752 12393
rect 4344 12384 4396 12436
rect 5172 12384 5224 12436
rect 7748 12316 7800 12368
rect 11520 12427 11572 12436
rect 11520 12393 11529 12427
rect 11529 12393 11563 12427
rect 11563 12393 11572 12427
rect 11520 12384 11572 12393
rect 12256 12384 12308 12436
rect 13452 12427 13504 12436
rect 13452 12393 13461 12427
rect 13461 12393 13495 12427
rect 13495 12393 13504 12427
rect 13452 12384 13504 12393
rect 14188 12384 14240 12436
rect 14280 12384 14332 12436
rect 15660 12427 15712 12436
rect 15660 12393 15669 12427
rect 15669 12393 15703 12427
rect 15703 12393 15712 12427
rect 15660 12384 15712 12393
rect 19248 12427 19300 12436
rect 19248 12393 19257 12427
rect 19257 12393 19291 12427
rect 19291 12393 19300 12427
rect 19248 12384 19300 12393
rect 9588 12359 9640 12368
rect 9588 12325 9597 12359
rect 9597 12325 9631 12359
rect 9631 12325 9640 12359
rect 9588 12316 9640 12325
rect 9772 12359 9824 12368
rect 9772 12325 9797 12359
rect 9797 12325 9824 12359
rect 9772 12316 9824 12325
rect 9956 12316 10008 12368
rect 3424 12248 3476 12300
rect 3608 12248 3660 12300
rect 4252 12291 4304 12300
rect 4252 12257 4261 12291
rect 4261 12257 4295 12291
rect 4295 12257 4304 12291
rect 4252 12248 4304 12257
rect 4620 12248 4672 12300
rect 5356 12248 5408 12300
rect 5908 12248 5960 12300
rect 4804 12180 4856 12232
rect 7012 12112 7064 12164
rect 2228 12087 2280 12096
rect 2228 12053 2237 12087
rect 2237 12053 2271 12087
rect 2271 12053 2280 12087
rect 2228 12044 2280 12053
rect 4160 12044 4212 12096
rect 7564 12044 7616 12096
rect 9588 12180 9640 12232
rect 11336 12291 11388 12300
rect 11336 12257 11345 12291
rect 11345 12257 11379 12291
rect 11379 12257 11388 12291
rect 11336 12248 11388 12257
rect 11428 12291 11480 12300
rect 11428 12257 11437 12291
rect 11437 12257 11471 12291
rect 11471 12257 11480 12291
rect 11428 12248 11480 12257
rect 11704 12291 11756 12300
rect 11704 12257 11713 12291
rect 11713 12257 11747 12291
rect 11747 12257 11756 12291
rect 11704 12248 11756 12257
rect 12164 12248 12216 12300
rect 12716 12248 12768 12300
rect 14832 12359 14884 12368
rect 14832 12325 14841 12359
rect 14841 12325 14875 12359
rect 14875 12325 14884 12359
rect 14832 12316 14884 12325
rect 11888 12180 11940 12232
rect 14280 12291 14332 12300
rect 14280 12257 14289 12291
rect 14289 12257 14323 12291
rect 14323 12257 14332 12291
rect 14280 12248 14332 12257
rect 14464 12248 14516 12300
rect 19708 12316 19760 12368
rect 16212 12248 16264 12300
rect 18512 12248 18564 12300
rect 18972 12248 19024 12300
rect 21640 12248 21692 12300
rect 22652 12384 22704 12436
rect 9128 12044 9180 12096
rect 10232 12044 10284 12096
rect 10324 12044 10376 12096
rect 12256 12044 12308 12096
rect 15568 12180 15620 12232
rect 16028 12180 16080 12232
rect 17868 12180 17920 12232
rect 19708 12180 19760 12232
rect 20076 12180 20128 12232
rect 23204 12359 23256 12368
rect 23204 12325 23213 12359
rect 23213 12325 23247 12359
rect 23247 12325 23256 12359
rect 23204 12316 23256 12325
rect 23388 12427 23440 12436
rect 23388 12393 23397 12427
rect 23397 12393 23431 12427
rect 23431 12393 23440 12427
rect 23388 12384 23440 12393
rect 23480 12384 23532 12436
rect 25044 12384 25096 12436
rect 25228 12427 25280 12436
rect 25228 12393 25237 12427
rect 25237 12393 25271 12427
rect 25271 12393 25280 12427
rect 25228 12384 25280 12393
rect 26424 12427 26476 12436
rect 26424 12393 26433 12427
rect 26433 12393 26467 12427
rect 26467 12393 26476 12427
rect 26424 12384 26476 12393
rect 24308 12316 24360 12368
rect 25412 12316 25464 12368
rect 22468 12248 22520 12300
rect 24400 12248 24452 12300
rect 22100 12180 22152 12232
rect 25688 12291 25740 12300
rect 25688 12257 25697 12291
rect 25697 12257 25731 12291
rect 25731 12257 25740 12291
rect 25688 12248 25740 12257
rect 26976 12316 27028 12368
rect 26056 12248 26108 12300
rect 26700 12291 26752 12300
rect 26700 12257 26709 12291
rect 26709 12257 26743 12291
rect 26743 12257 26752 12291
rect 26700 12248 26752 12257
rect 26148 12180 26200 12232
rect 13636 12112 13688 12164
rect 18144 12044 18196 12096
rect 19156 12044 19208 12096
rect 24584 12112 24636 12164
rect 25688 12112 25740 12164
rect 26884 12291 26936 12300
rect 26884 12257 26893 12291
rect 26893 12257 26927 12291
rect 26927 12257 26936 12291
rect 26884 12248 26936 12257
rect 22560 12087 22612 12096
rect 22560 12053 22569 12087
rect 22569 12053 22603 12087
rect 22603 12053 22612 12087
rect 22560 12044 22612 12053
rect 23204 12044 23256 12096
rect 3756 11942 3808 11994
rect 3820 11942 3872 11994
rect 3884 11942 3936 11994
rect 3948 11942 4000 11994
rect 4012 11942 4064 11994
rect 10472 11942 10524 11994
rect 10536 11942 10588 11994
rect 10600 11942 10652 11994
rect 10664 11942 10716 11994
rect 10728 11942 10780 11994
rect 17188 11942 17240 11994
rect 17252 11942 17304 11994
rect 17316 11942 17368 11994
rect 17380 11942 17432 11994
rect 17444 11942 17496 11994
rect 23904 11942 23956 11994
rect 23968 11942 24020 11994
rect 24032 11942 24084 11994
rect 24096 11942 24148 11994
rect 24160 11942 24212 11994
rect 1124 11840 1176 11892
rect 3608 11840 3660 11892
rect 4344 11840 4396 11892
rect 4804 11840 4856 11892
rect 5908 11840 5960 11892
rect 6920 11840 6972 11892
rect 2228 11704 2280 11756
rect 1400 11636 1452 11688
rect 6644 11704 6696 11756
rect 7472 11883 7524 11892
rect 7472 11849 7481 11883
rect 7481 11849 7515 11883
rect 7515 11849 7524 11883
rect 7472 11840 7524 11849
rect 9588 11883 9640 11892
rect 9588 11849 9597 11883
rect 9597 11849 9631 11883
rect 9631 11849 9640 11883
rect 9588 11840 9640 11849
rect 12716 11840 12768 11892
rect 13268 11840 13320 11892
rect 13452 11840 13504 11892
rect 15660 11840 15712 11892
rect 16212 11840 16264 11892
rect 17868 11883 17920 11892
rect 17868 11849 17877 11883
rect 17877 11849 17911 11883
rect 17911 11849 17920 11883
rect 17868 11840 17920 11849
rect 18144 11883 18196 11892
rect 18144 11849 18153 11883
rect 18153 11849 18187 11883
rect 18187 11849 18196 11883
rect 18144 11840 18196 11849
rect 18972 11883 19024 11892
rect 18972 11849 18981 11883
rect 18981 11849 19015 11883
rect 19015 11849 19024 11883
rect 18972 11840 19024 11849
rect 19156 11883 19208 11892
rect 19156 11849 19165 11883
rect 19165 11849 19199 11883
rect 19199 11849 19208 11883
rect 19156 11840 19208 11849
rect 21824 11883 21876 11892
rect 21824 11849 21833 11883
rect 21833 11849 21867 11883
rect 21867 11849 21876 11883
rect 21824 11840 21876 11849
rect 24768 11840 24820 11892
rect 20996 11772 21048 11824
rect 23112 11772 23164 11824
rect 3424 11636 3476 11688
rect 5356 11636 5408 11688
rect 4068 11568 4120 11620
rect 1860 11500 1912 11552
rect 3424 11543 3476 11552
rect 3424 11509 3451 11543
rect 3451 11509 3476 11543
rect 3424 11500 3476 11509
rect 6736 11636 6788 11688
rect 7564 11679 7616 11688
rect 7564 11645 7573 11679
rect 7573 11645 7607 11679
rect 7607 11645 7616 11679
rect 7564 11636 7616 11645
rect 8208 11636 8260 11688
rect 11888 11704 11940 11756
rect 6552 11568 6604 11620
rect 10416 11568 10468 11620
rect 12532 11636 12584 11688
rect 14556 11636 14608 11688
rect 16396 11704 16448 11756
rect 21088 11704 21140 11756
rect 22100 11704 22152 11756
rect 19064 11636 19116 11688
rect 19708 11679 19760 11688
rect 19708 11645 19717 11679
rect 19717 11645 19751 11679
rect 19751 11645 19760 11679
rect 19708 11636 19760 11645
rect 19984 11679 20036 11688
rect 19984 11645 19993 11679
rect 19993 11645 20027 11679
rect 20027 11645 20036 11679
rect 19984 11636 20036 11645
rect 12900 11611 12952 11620
rect 6920 11500 6972 11552
rect 9404 11500 9456 11552
rect 11336 11500 11388 11552
rect 12532 11543 12584 11552
rect 12532 11509 12541 11543
rect 12541 11509 12575 11543
rect 12575 11509 12584 11543
rect 12532 11500 12584 11509
rect 12900 11577 12927 11611
rect 12927 11577 12952 11611
rect 12900 11568 12952 11577
rect 12992 11568 13044 11620
rect 13636 11568 13688 11620
rect 14740 11568 14792 11620
rect 15384 11568 15436 11620
rect 16948 11568 17000 11620
rect 18328 11611 18380 11620
rect 18328 11577 18337 11611
rect 18337 11577 18371 11611
rect 18371 11577 18380 11611
rect 18328 11568 18380 11577
rect 14372 11500 14424 11552
rect 15568 11500 15620 11552
rect 17132 11500 17184 11552
rect 18880 11500 18932 11552
rect 19616 11543 19668 11552
rect 19616 11509 19625 11543
rect 19625 11509 19659 11543
rect 19659 11509 19668 11543
rect 19616 11500 19668 11509
rect 20352 11500 20404 11552
rect 21732 11679 21784 11688
rect 21732 11645 21741 11679
rect 21741 11645 21775 11679
rect 21775 11645 21784 11679
rect 21732 11636 21784 11645
rect 22284 11636 22336 11688
rect 22376 11679 22428 11688
rect 22376 11645 22385 11679
rect 22385 11645 22419 11679
rect 22419 11645 22428 11679
rect 22376 11636 22428 11645
rect 20904 11500 20956 11552
rect 22008 11568 22060 11620
rect 22560 11679 22612 11688
rect 22560 11645 22569 11679
rect 22569 11645 22603 11679
rect 22603 11645 22612 11679
rect 22560 11636 22612 11645
rect 22836 11500 22888 11552
rect 23020 11543 23072 11552
rect 23020 11509 23029 11543
rect 23029 11509 23063 11543
rect 23063 11509 23072 11543
rect 23020 11500 23072 11509
rect 23204 11611 23256 11620
rect 23204 11577 23213 11611
rect 23213 11577 23247 11611
rect 23247 11577 23256 11611
rect 23204 11568 23256 11577
rect 23664 11568 23716 11620
rect 25688 11840 25740 11892
rect 26608 11840 26660 11892
rect 26976 11840 27028 11892
rect 24952 11679 25004 11688
rect 24952 11645 24961 11679
rect 24961 11645 24995 11679
rect 24995 11645 25004 11679
rect 24952 11636 25004 11645
rect 25136 11679 25188 11688
rect 25136 11645 25145 11679
rect 25145 11645 25179 11679
rect 25179 11645 25188 11679
rect 25136 11636 25188 11645
rect 25596 11704 25648 11756
rect 23480 11500 23532 11552
rect 24492 11500 24544 11552
rect 24584 11500 24636 11552
rect 26424 11636 26476 11688
rect 7114 11398 7166 11450
rect 7178 11398 7230 11450
rect 7242 11398 7294 11450
rect 7306 11398 7358 11450
rect 7370 11398 7422 11450
rect 13830 11398 13882 11450
rect 13894 11398 13946 11450
rect 13958 11398 14010 11450
rect 14022 11398 14074 11450
rect 14086 11398 14138 11450
rect 20546 11398 20598 11450
rect 20610 11398 20662 11450
rect 20674 11398 20726 11450
rect 20738 11398 20790 11450
rect 20802 11398 20854 11450
rect 27262 11398 27314 11450
rect 27326 11398 27378 11450
rect 27390 11398 27442 11450
rect 27454 11398 27506 11450
rect 27518 11398 27570 11450
rect 1400 11339 1452 11348
rect 1400 11305 1409 11339
rect 1409 11305 1443 11339
rect 1443 11305 1452 11339
rect 1400 11296 1452 11305
rect 3240 11296 3292 11348
rect 6736 11339 6788 11348
rect 6736 11305 6745 11339
rect 6745 11305 6779 11339
rect 6779 11305 6788 11339
rect 6736 11296 6788 11305
rect 6920 11296 6972 11348
rect 9128 11296 9180 11348
rect 8852 11228 8904 11280
rect 1676 11160 1728 11212
rect 1860 11203 1912 11212
rect 1860 11169 1869 11203
rect 1869 11169 1903 11203
rect 1903 11169 1912 11203
rect 1860 11160 1912 11169
rect 4344 11160 4396 11212
rect 6644 11160 6696 11212
rect 6828 11160 6880 11212
rect 7012 11203 7064 11212
rect 7012 11169 7021 11203
rect 7021 11169 7055 11203
rect 7055 11169 7064 11203
rect 7012 11160 7064 11169
rect 7564 11160 7616 11212
rect 2320 11092 2372 11144
rect 3424 11092 3476 11144
rect 6092 11092 6144 11144
rect 2780 11024 2832 11076
rect 7012 11024 7064 11076
rect 8208 11092 8260 11144
rect 8944 11024 8996 11076
rect 9956 11296 10008 11348
rect 10416 11339 10468 11348
rect 10416 11305 10425 11339
rect 10425 11305 10459 11339
rect 10459 11305 10468 11339
rect 10416 11296 10468 11305
rect 9588 11228 9640 11280
rect 11888 11296 11940 11348
rect 12532 11296 12584 11348
rect 9864 11160 9916 11212
rect 10232 11203 10284 11212
rect 10232 11169 10241 11203
rect 10241 11169 10275 11203
rect 10275 11169 10284 11203
rect 10232 11160 10284 11169
rect 11612 11160 11664 11212
rect 13636 11228 13688 11280
rect 13452 11203 13504 11212
rect 13452 11169 13486 11203
rect 13486 11169 13504 11203
rect 13452 11160 13504 11169
rect 15292 11296 15344 11348
rect 15384 11339 15436 11348
rect 15384 11305 15393 11339
rect 15393 11305 15427 11339
rect 15427 11305 15436 11339
rect 15384 11296 15436 11305
rect 14280 11228 14332 11280
rect 9220 11092 9272 11144
rect 15292 11135 15344 11144
rect 15292 11101 15301 11135
rect 15301 11101 15335 11135
rect 15335 11101 15344 11135
rect 15292 11092 15344 11101
rect 15568 11203 15620 11212
rect 15568 11169 15577 11203
rect 15577 11169 15611 11203
rect 15611 11169 15620 11203
rect 15568 11160 15620 11169
rect 16948 11339 17000 11348
rect 16948 11305 16957 11339
rect 16957 11305 16991 11339
rect 16991 11305 17000 11339
rect 16948 11296 17000 11305
rect 16580 11228 16632 11280
rect 16120 11203 16172 11212
rect 16120 11169 16129 11203
rect 16129 11169 16163 11203
rect 16163 11169 16172 11203
rect 16120 11160 16172 11169
rect 16212 11160 16264 11212
rect 17132 11203 17184 11212
rect 17132 11169 17141 11203
rect 17141 11169 17175 11203
rect 17175 11169 17184 11203
rect 17132 11160 17184 11169
rect 17868 11160 17920 11212
rect 19984 11296 20036 11348
rect 20444 11296 20496 11348
rect 21732 11296 21784 11348
rect 22008 11296 22060 11348
rect 22468 11339 22520 11348
rect 22468 11305 22477 11339
rect 22477 11305 22511 11339
rect 22511 11305 22520 11339
rect 22468 11296 22520 11305
rect 19616 11271 19668 11280
rect 19616 11237 19625 11271
rect 19625 11237 19659 11271
rect 19659 11237 19668 11271
rect 19616 11228 19668 11237
rect 20812 11271 20864 11280
rect 20812 11237 20830 11271
rect 20830 11237 20864 11271
rect 20812 11228 20864 11237
rect 21548 11228 21600 11280
rect 23204 11296 23256 11348
rect 23480 11296 23532 11348
rect 23572 11296 23624 11348
rect 24584 11296 24636 11348
rect 26148 11296 26200 11348
rect 23020 11228 23072 11280
rect 20076 11160 20128 11212
rect 22008 11160 22060 11212
rect 27068 11203 27120 11212
rect 27068 11169 27077 11203
rect 27077 11169 27111 11203
rect 27111 11169 27120 11203
rect 27068 11160 27120 11169
rect 18420 11092 18472 11144
rect 9772 11024 9824 11076
rect 10324 11024 10376 11076
rect 10968 11024 11020 11076
rect 2504 10956 2556 11008
rect 2688 10956 2740 11008
rect 6184 10999 6236 11008
rect 6184 10965 6193 10999
rect 6193 10965 6227 10999
rect 6227 10965 6236 10999
rect 6184 10956 6236 10965
rect 9128 10956 9180 11008
rect 9312 10956 9364 11008
rect 12900 10956 12952 11008
rect 14648 10999 14700 11008
rect 14648 10965 14657 10999
rect 14657 10965 14691 10999
rect 14691 10965 14700 10999
rect 14648 10956 14700 10965
rect 16120 10999 16172 11008
rect 16120 10965 16129 10999
rect 16129 10965 16163 10999
rect 16163 10965 16172 10999
rect 16120 10956 16172 10965
rect 17868 10956 17920 11008
rect 17960 10956 18012 11008
rect 22376 11092 22428 11144
rect 25596 11092 25648 11144
rect 26056 11135 26108 11144
rect 26056 11101 26065 11135
rect 26065 11101 26099 11135
rect 26099 11101 26108 11135
rect 26056 11092 26108 11101
rect 23572 11024 23624 11076
rect 20444 10956 20496 11008
rect 21640 10956 21692 11008
rect 22192 10956 22244 11008
rect 23664 10956 23716 11008
rect 25412 10956 25464 11008
rect 27068 10956 27120 11008
rect 3756 10854 3808 10906
rect 3820 10854 3872 10906
rect 3884 10854 3936 10906
rect 3948 10854 4000 10906
rect 4012 10854 4064 10906
rect 10472 10854 10524 10906
rect 10536 10854 10588 10906
rect 10600 10854 10652 10906
rect 10664 10854 10716 10906
rect 10728 10854 10780 10906
rect 17188 10854 17240 10906
rect 17252 10854 17304 10906
rect 17316 10854 17368 10906
rect 17380 10854 17432 10906
rect 17444 10854 17496 10906
rect 23904 10854 23956 10906
rect 23968 10854 24020 10906
rect 24032 10854 24084 10906
rect 24096 10854 24148 10906
rect 24160 10854 24212 10906
rect 3516 10795 3568 10804
rect 3516 10761 3525 10795
rect 3525 10761 3559 10795
rect 3559 10761 3568 10795
rect 3516 10752 3568 10761
rect 6184 10752 6236 10804
rect 11336 10752 11388 10804
rect 12992 10752 13044 10804
rect 13452 10752 13504 10804
rect 14648 10752 14700 10804
rect 2964 10616 3016 10668
rect 2596 10548 2648 10600
rect 2780 10591 2832 10600
rect 2780 10557 2789 10591
rect 2789 10557 2823 10591
rect 2823 10557 2832 10591
rect 2780 10548 2832 10557
rect 3424 10548 3476 10600
rect 4804 10591 4856 10600
rect 4804 10557 4813 10591
rect 4813 10557 4847 10591
rect 4847 10557 4856 10591
rect 4804 10548 4856 10557
rect 3516 10523 3568 10532
rect 3516 10489 3525 10523
rect 3525 10489 3559 10523
rect 3559 10489 3568 10523
rect 3516 10480 3568 10489
rect 9772 10684 9824 10736
rect 11244 10684 11296 10736
rect 7012 10659 7064 10668
rect 7012 10625 7021 10659
rect 7021 10625 7055 10659
rect 7055 10625 7064 10659
rect 7012 10616 7064 10625
rect 6000 10548 6052 10600
rect 6644 10591 6696 10600
rect 6644 10557 6653 10591
rect 6653 10557 6687 10591
rect 6687 10557 6696 10591
rect 6644 10548 6696 10557
rect 6828 10548 6880 10600
rect 8944 10591 8996 10600
rect 8944 10557 8953 10591
rect 8953 10557 8987 10591
rect 8987 10557 8996 10591
rect 8944 10548 8996 10557
rect 9128 10548 9180 10600
rect 9220 10591 9272 10600
rect 9220 10557 9229 10591
rect 9229 10557 9263 10591
rect 9263 10557 9272 10591
rect 9220 10548 9272 10557
rect 9312 10591 9364 10600
rect 9312 10557 9321 10591
rect 9321 10557 9355 10591
rect 9355 10557 9364 10591
rect 9312 10548 9364 10557
rect 9864 10616 9916 10668
rect 9496 10548 9548 10600
rect 10324 10591 10376 10600
rect 10324 10557 10333 10591
rect 10333 10557 10367 10591
rect 10367 10557 10376 10591
rect 10324 10548 10376 10557
rect 10876 10591 10928 10600
rect 10876 10557 10885 10591
rect 10885 10557 10919 10591
rect 10919 10557 10928 10591
rect 10876 10548 10928 10557
rect 11244 10548 11296 10600
rect 12256 10684 12308 10736
rect 18880 10752 18932 10804
rect 20076 10795 20128 10804
rect 20076 10761 20085 10795
rect 20085 10761 20119 10795
rect 20119 10761 20128 10795
rect 20076 10752 20128 10761
rect 21088 10752 21140 10804
rect 25412 10795 25464 10804
rect 25412 10761 25421 10795
rect 25421 10761 25455 10795
rect 25455 10761 25464 10795
rect 25412 10752 25464 10761
rect 26884 10795 26936 10804
rect 12808 10616 12860 10668
rect 12900 10659 12952 10668
rect 12900 10625 12909 10659
rect 12909 10625 12943 10659
rect 12943 10625 12952 10659
rect 12900 10616 12952 10625
rect 12992 10616 13044 10668
rect 7656 10480 7708 10532
rect 12164 10591 12216 10600
rect 12164 10557 12173 10591
rect 12173 10557 12207 10591
rect 12207 10557 12216 10591
rect 12164 10548 12216 10557
rect 12072 10480 12124 10532
rect 13268 10591 13320 10600
rect 13268 10557 13277 10591
rect 13277 10557 13311 10591
rect 13311 10557 13320 10591
rect 13268 10548 13320 10557
rect 14004 10591 14056 10600
rect 14004 10557 14013 10591
rect 14013 10557 14047 10591
rect 14047 10557 14056 10591
rect 14004 10548 14056 10557
rect 14280 10548 14332 10600
rect 14740 10548 14792 10600
rect 15384 10548 15436 10600
rect 2320 10412 2372 10464
rect 2964 10455 3016 10464
rect 2964 10421 2973 10455
rect 2973 10421 3007 10455
rect 3007 10421 3016 10455
rect 2964 10412 3016 10421
rect 3608 10412 3660 10464
rect 5080 10412 5132 10464
rect 6276 10412 6328 10464
rect 7472 10455 7524 10464
rect 7472 10421 7481 10455
rect 7481 10421 7515 10455
rect 7515 10421 7524 10455
rect 7472 10412 7524 10421
rect 8852 10412 8904 10464
rect 8944 10412 8996 10464
rect 10140 10455 10192 10464
rect 10140 10421 10149 10455
rect 10149 10421 10183 10455
rect 10183 10421 10192 10455
rect 10140 10412 10192 10421
rect 11060 10412 11112 10464
rect 11152 10412 11204 10464
rect 12256 10412 12308 10464
rect 14556 10523 14608 10532
rect 14556 10489 14565 10523
rect 14565 10489 14599 10523
rect 14599 10489 14608 10523
rect 14556 10480 14608 10489
rect 15660 10591 15712 10600
rect 15660 10557 15669 10591
rect 15669 10557 15703 10591
rect 15703 10557 15712 10591
rect 15660 10548 15712 10557
rect 15844 10591 15896 10600
rect 15844 10557 15853 10591
rect 15853 10557 15887 10591
rect 15887 10557 15896 10591
rect 15844 10548 15896 10557
rect 16212 10548 16264 10600
rect 16028 10523 16080 10532
rect 16028 10489 16037 10523
rect 16037 10489 16071 10523
rect 16071 10489 16080 10523
rect 16028 10480 16080 10489
rect 17040 10684 17092 10736
rect 17040 10591 17092 10600
rect 17040 10557 17049 10591
rect 17049 10557 17083 10591
rect 17083 10557 17092 10591
rect 17040 10548 17092 10557
rect 17960 10684 18012 10736
rect 20444 10684 20496 10736
rect 26884 10761 26893 10795
rect 26893 10761 26927 10795
rect 26927 10761 26936 10795
rect 26884 10752 26936 10761
rect 17776 10616 17828 10668
rect 22100 10659 22152 10668
rect 22100 10625 22109 10659
rect 22109 10625 22143 10659
rect 22143 10625 22152 10659
rect 22100 10616 22152 10625
rect 22468 10616 22520 10668
rect 22836 10616 22888 10668
rect 17868 10591 17920 10600
rect 17868 10557 17877 10591
rect 17877 10557 17911 10591
rect 17911 10557 17920 10591
rect 17868 10548 17920 10557
rect 14372 10455 14424 10464
rect 14372 10421 14399 10455
rect 14399 10421 14424 10455
rect 14372 10412 14424 10421
rect 15384 10455 15436 10464
rect 15384 10421 15393 10455
rect 15393 10421 15427 10455
rect 15427 10421 15436 10455
rect 15384 10412 15436 10421
rect 17224 10455 17276 10464
rect 17224 10421 17233 10455
rect 17233 10421 17267 10455
rect 17267 10421 17276 10455
rect 17224 10412 17276 10421
rect 18236 10548 18288 10600
rect 18420 10591 18472 10600
rect 18420 10557 18429 10591
rect 18429 10557 18463 10591
rect 18463 10557 18472 10591
rect 18420 10548 18472 10557
rect 20352 10591 20404 10600
rect 20352 10557 20361 10591
rect 20361 10557 20395 10591
rect 20395 10557 20404 10591
rect 20352 10548 20404 10557
rect 20996 10548 21048 10600
rect 22008 10591 22060 10600
rect 22008 10557 22017 10591
rect 22017 10557 22051 10591
rect 22051 10557 22060 10591
rect 22008 10548 22060 10557
rect 18512 10480 18564 10532
rect 19892 10480 19944 10532
rect 23296 10591 23348 10600
rect 23296 10557 23305 10591
rect 23305 10557 23339 10591
rect 23339 10557 23348 10591
rect 23296 10548 23348 10557
rect 24308 10616 24360 10668
rect 24768 10616 24820 10668
rect 23572 10548 23624 10600
rect 25320 10548 25372 10600
rect 25596 10548 25648 10600
rect 23848 10480 23900 10532
rect 24768 10480 24820 10532
rect 17960 10455 18012 10464
rect 17960 10421 17969 10455
rect 17969 10421 18003 10455
rect 18003 10421 18012 10455
rect 17960 10412 18012 10421
rect 24860 10455 24912 10464
rect 24860 10421 24869 10455
rect 24869 10421 24903 10455
rect 24903 10421 24912 10455
rect 24860 10412 24912 10421
rect 24952 10455 25004 10464
rect 24952 10421 24961 10455
rect 24961 10421 24995 10455
rect 24995 10421 25004 10455
rect 24952 10412 25004 10421
rect 25504 10412 25556 10464
rect 7114 10310 7166 10362
rect 7178 10310 7230 10362
rect 7242 10310 7294 10362
rect 7306 10310 7358 10362
rect 7370 10310 7422 10362
rect 13830 10310 13882 10362
rect 13894 10310 13946 10362
rect 13958 10310 14010 10362
rect 14022 10310 14074 10362
rect 14086 10310 14138 10362
rect 20546 10310 20598 10362
rect 20610 10310 20662 10362
rect 20674 10310 20726 10362
rect 20738 10310 20790 10362
rect 20802 10310 20854 10362
rect 27262 10310 27314 10362
rect 27326 10310 27378 10362
rect 27390 10310 27442 10362
rect 27454 10310 27506 10362
rect 27518 10310 27570 10362
rect 2596 10072 2648 10124
rect 2872 10140 2924 10192
rect 3332 10208 3384 10260
rect 4804 10208 4856 10260
rect 6644 10208 6696 10260
rect 7472 10208 7524 10260
rect 2320 10047 2372 10056
rect 2320 10013 2329 10047
rect 2329 10013 2363 10047
rect 2363 10013 2372 10047
rect 2320 10004 2372 10013
rect 2688 10004 2740 10056
rect 4896 10072 4948 10124
rect 6276 10115 6328 10124
rect 6276 10081 6285 10115
rect 6285 10081 6319 10115
rect 6319 10081 6328 10115
rect 6276 10072 6328 10081
rect 6920 10115 6972 10124
rect 6920 10081 6929 10115
rect 6929 10081 6963 10115
rect 6963 10081 6972 10115
rect 6920 10072 6972 10081
rect 4252 10047 4304 10056
rect 4252 10013 4261 10047
rect 4261 10013 4295 10047
rect 4295 10013 4304 10047
rect 4252 10004 4304 10013
rect 6828 10004 6880 10056
rect 7656 10140 7708 10192
rect 10140 10140 10192 10192
rect 8024 10047 8076 10056
rect 8024 10013 8033 10047
rect 8033 10013 8067 10047
rect 8067 10013 8076 10047
rect 8024 10004 8076 10013
rect 8668 10115 8720 10124
rect 8668 10081 8677 10115
rect 8677 10081 8711 10115
rect 8711 10081 8720 10115
rect 8668 10072 8720 10081
rect 2688 9911 2740 9920
rect 2688 9877 2697 9911
rect 2697 9877 2731 9911
rect 2731 9877 2740 9911
rect 2688 9868 2740 9877
rect 3516 9868 3568 9920
rect 8484 9936 8536 9988
rect 8760 10004 8812 10056
rect 8944 10115 8996 10124
rect 8944 10081 8953 10115
rect 8953 10081 8987 10115
rect 8987 10081 8996 10115
rect 8944 10072 8996 10081
rect 9128 10115 9180 10124
rect 9128 10081 9137 10115
rect 9137 10081 9171 10115
rect 9171 10081 9180 10115
rect 9128 10072 9180 10081
rect 10048 10072 10100 10124
rect 10324 10208 10376 10260
rect 11612 10208 11664 10260
rect 11888 10251 11940 10260
rect 11888 10217 11897 10251
rect 11897 10217 11931 10251
rect 11931 10217 11940 10251
rect 11888 10208 11940 10217
rect 14188 10208 14240 10260
rect 10416 10140 10468 10192
rect 11336 10183 11388 10192
rect 11336 10149 11345 10183
rect 11345 10149 11379 10183
rect 11379 10149 11388 10183
rect 11336 10140 11388 10149
rect 12348 10140 12400 10192
rect 9220 10004 9272 10056
rect 9404 10047 9456 10056
rect 9404 10013 9413 10047
rect 9413 10013 9447 10047
rect 9447 10013 9456 10047
rect 9404 10004 9456 10013
rect 6920 9868 6972 9920
rect 8392 9911 8444 9920
rect 8392 9877 8401 9911
rect 8401 9877 8435 9911
rect 8435 9877 8444 9911
rect 8392 9868 8444 9877
rect 9036 9868 9088 9920
rect 9772 9868 9824 9920
rect 10324 9868 10376 9920
rect 10876 9868 10928 9920
rect 11152 9911 11204 9920
rect 11152 9877 11161 9911
rect 11161 9877 11195 9911
rect 11195 9877 11204 9911
rect 11152 9868 11204 9877
rect 11888 10072 11940 10124
rect 11980 10115 12032 10124
rect 11980 10081 11989 10115
rect 11989 10081 12023 10115
rect 12023 10081 12032 10115
rect 11980 10072 12032 10081
rect 12808 10140 12860 10192
rect 13268 10140 13320 10192
rect 12992 10115 13044 10124
rect 12992 10081 13001 10115
rect 13001 10081 13035 10115
rect 13035 10081 13044 10115
rect 12992 10072 13044 10081
rect 13176 10115 13228 10124
rect 13176 10081 13185 10115
rect 13185 10081 13219 10115
rect 13219 10081 13228 10115
rect 13176 10072 13228 10081
rect 14648 10115 14700 10124
rect 14648 10081 14657 10115
rect 14657 10081 14691 10115
rect 14691 10081 14700 10115
rect 14648 10072 14700 10081
rect 15844 10208 15896 10260
rect 16028 10208 16080 10260
rect 15292 10140 15344 10192
rect 17040 10208 17092 10260
rect 18328 10208 18380 10260
rect 12532 10004 12584 10056
rect 14556 10004 14608 10056
rect 16028 10072 16080 10124
rect 17960 10140 18012 10192
rect 16212 10115 16264 10124
rect 16212 10081 16221 10115
rect 16221 10081 16255 10115
rect 16255 10081 16264 10115
rect 16212 10072 16264 10081
rect 18420 10140 18472 10192
rect 18880 10208 18932 10260
rect 23296 10208 23348 10260
rect 23480 10208 23532 10260
rect 21548 10140 21600 10192
rect 15568 10004 15620 10056
rect 15660 10047 15712 10056
rect 15660 10013 15669 10047
rect 15669 10013 15703 10047
rect 15703 10013 15712 10047
rect 15660 10004 15712 10013
rect 18144 10115 18196 10124
rect 18144 10081 18153 10115
rect 18153 10081 18187 10115
rect 18187 10081 18196 10115
rect 18144 10072 18196 10081
rect 17776 10047 17828 10056
rect 17776 10013 17785 10047
rect 17785 10013 17819 10047
rect 17819 10013 17828 10047
rect 17776 10004 17828 10013
rect 18512 10047 18564 10056
rect 18512 10013 18521 10047
rect 18521 10013 18555 10047
rect 18555 10013 18564 10047
rect 18512 10004 18564 10013
rect 12256 9911 12308 9920
rect 12256 9877 12265 9911
rect 12265 9877 12299 9911
rect 12299 9877 12308 9911
rect 12256 9868 12308 9877
rect 16396 9936 16448 9988
rect 12900 9868 12952 9920
rect 13268 9868 13320 9920
rect 14924 9868 14976 9920
rect 15200 9868 15252 9920
rect 17040 9868 17092 9920
rect 20076 10115 20128 10124
rect 20076 10081 20085 10115
rect 20085 10081 20119 10115
rect 20119 10081 20128 10115
rect 20076 10072 20128 10081
rect 22284 10072 22336 10124
rect 22560 10115 22612 10124
rect 22560 10081 22569 10115
rect 22569 10081 22603 10115
rect 22603 10081 22612 10115
rect 22560 10072 22612 10081
rect 22836 10115 22888 10124
rect 22836 10081 22845 10115
rect 22845 10081 22879 10115
rect 22879 10081 22888 10115
rect 22836 10072 22888 10081
rect 23020 10115 23072 10124
rect 23020 10081 23029 10115
rect 23029 10081 23063 10115
rect 23063 10081 23072 10115
rect 23020 10072 23072 10081
rect 23388 10072 23440 10124
rect 24308 10115 24360 10124
rect 24308 10081 24317 10115
rect 24317 10081 24351 10115
rect 24351 10081 24360 10115
rect 24308 10072 24360 10081
rect 24492 10115 24544 10124
rect 24492 10081 24501 10115
rect 24501 10081 24535 10115
rect 24535 10081 24544 10115
rect 24492 10072 24544 10081
rect 24584 10115 24636 10124
rect 24584 10081 24593 10115
rect 24593 10081 24627 10115
rect 24627 10081 24636 10115
rect 24584 10072 24636 10081
rect 24860 10140 24912 10192
rect 25136 10140 25188 10192
rect 26148 10208 26200 10260
rect 26424 10251 26476 10260
rect 26424 10217 26433 10251
rect 26433 10217 26467 10251
rect 26467 10217 26476 10251
rect 26424 10208 26476 10217
rect 26976 10115 27028 10124
rect 26976 10081 26985 10115
rect 26985 10081 27019 10115
rect 27019 10081 27028 10115
rect 26976 10072 27028 10081
rect 25136 10004 25188 10056
rect 23848 9936 23900 9988
rect 24584 9936 24636 9988
rect 26056 9936 26108 9988
rect 22100 9911 22152 9920
rect 22100 9877 22109 9911
rect 22109 9877 22143 9911
rect 22143 9877 22152 9911
rect 22100 9868 22152 9877
rect 23756 9868 23808 9920
rect 3756 9766 3808 9818
rect 3820 9766 3872 9818
rect 3884 9766 3936 9818
rect 3948 9766 4000 9818
rect 4012 9766 4064 9818
rect 10472 9766 10524 9818
rect 10536 9766 10588 9818
rect 10600 9766 10652 9818
rect 10664 9766 10716 9818
rect 10728 9766 10780 9818
rect 17188 9766 17240 9818
rect 17252 9766 17304 9818
rect 17316 9766 17368 9818
rect 17380 9766 17432 9818
rect 17444 9766 17496 9818
rect 23904 9766 23956 9818
rect 23968 9766 24020 9818
rect 24032 9766 24084 9818
rect 24096 9766 24148 9818
rect 24160 9766 24212 9818
rect 3332 9664 3384 9716
rect 4896 9707 4948 9716
rect 4896 9673 4905 9707
rect 4905 9673 4939 9707
rect 4939 9673 4948 9707
rect 4896 9664 4948 9673
rect 7564 9664 7616 9716
rect 12440 9664 12492 9716
rect 13176 9664 13228 9716
rect 2964 9639 3016 9648
rect 2964 9605 2973 9639
rect 2973 9605 3007 9639
rect 3007 9605 3016 9639
rect 2964 9596 3016 9605
rect 7748 9596 7800 9648
rect 12072 9596 12124 9648
rect 12164 9596 12216 9648
rect 14648 9664 14700 9716
rect 15200 9707 15252 9716
rect 15200 9673 15209 9707
rect 15209 9673 15243 9707
rect 15243 9673 15252 9707
rect 15200 9664 15252 9673
rect 15384 9664 15436 9716
rect 18236 9664 18288 9716
rect 22284 9664 22336 9716
rect 23664 9707 23716 9716
rect 23664 9673 23673 9707
rect 23673 9673 23707 9707
rect 23707 9673 23716 9707
rect 23664 9664 23716 9673
rect 15660 9596 15712 9648
rect 2688 9528 2740 9580
rect 2320 9460 2372 9512
rect 2504 9460 2556 9512
rect 2872 9460 2924 9512
rect 9404 9528 9456 9580
rect 3608 9460 3660 9512
rect 4804 9460 4856 9512
rect 5080 9503 5132 9512
rect 5080 9469 5089 9503
rect 5089 9469 5123 9503
rect 5123 9469 5132 9503
rect 5080 9460 5132 9469
rect 7840 9503 7892 9512
rect 7840 9469 7849 9503
rect 7849 9469 7883 9503
rect 7883 9469 7892 9503
rect 7840 9460 7892 9469
rect 1952 9435 2004 9444
rect 1952 9401 1961 9435
rect 1961 9401 1995 9435
rect 1995 9401 2004 9435
rect 1952 9392 2004 9401
rect 2780 9392 2832 9444
rect 2964 9324 3016 9376
rect 3424 9324 3476 9376
rect 6920 9392 6972 9444
rect 7472 9324 7524 9376
rect 8760 9503 8812 9512
rect 8760 9469 8769 9503
rect 8769 9469 8803 9503
rect 8803 9469 8812 9503
rect 8760 9460 8812 9469
rect 9128 9460 9180 9512
rect 9588 9503 9640 9512
rect 9588 9469 9597 9503
rect 9597 9469 9631 9503
rect 9631 9469 9640 9503
rect 9588 9460 9640 9469
rect 11060 9528 11112 9580
rect 10324 9460 10376 9512
rect 8668 9324 8720 9376
rect 8944 9324 8996 9376
rect 11336 9367 11388 9376
rect 11336 9333 11345 9367
rect 11345 9333 11379 9367
rect 11379 9333 11388 9367
rect 11336 9324 11388 9333
rect 12348 9528 12400 9580
rect 11704 9460 11756 9512
rect 11980 9460 12032 9512
rect 12164 9503 12216 9512
rect 12164 9469 12173 9503
rect 12173 9469 12207 9503
rect 12207 9469 12216 9503
rect 12164 9460 12216 9469
rect 12440 9503 12492 9512
rect 12440 9469 12449 9503
rect 12449 9469 12483 9503
rect 12483 9469 12492 9503
rect 12440 9460 12492 9469
rect 13084 9528 13136 9580
rect 15568 9528 15620 9580
rect 12900 9503 12952 9512
rect 12900 9469 12909 9503
rect 12909 9469 12943 9503
rect 12943 9469 12952 9503
rect 12900 9460 12952 9469
rect 12992 9503 13044 9512
rect 12992 9469 13001 9503
rect 13001 9469 13035 9503
rect 13035 9469 13044 9503
rect 12992 9460 13044 9469
rect 13176 9503 13228 9512
rect 13176 9469 13185 9503
rect 13185 9469 13219 9503
rect 13219 9469 13228 9503
rect 13176 9460 13228 9469
rect 13268 9503 13320 9512
rect 13268 9469 13277 9503
rect 13277 9469 13311 9503
rect 13311 9469 13320 9503
rect 13268 9460 13320 9469
rect 13636 9460 13688 9512
rect 16304 9528 16356 9580
rect 15936 9460 15988 9512
rect 11980 9367 12032 9376
rect 11980 9333 11989 9367
rect 11989 9333 12023 9367
rect 12023 9333 12032 9367
rect 11980 9324 12032 9333
rect 12716 9367 12768 9376
rect 12716 9333 12725 9367
rect 12725 9333 12759 9367
rect 12759 9333 12768 9367
rect 12716 9324 12768 9333
rect 12808 9324 12860 9376
rect 12992 9324 13044 9376
rect 13544 9324 13596 9376
rect 14372 9392 14424 9444
rect 15384 9435 15436 9444
rect 15384 9401 15393 9435
rect 15393 9401 15427 9435
rect 15427 9401 15436 9435
rect 15384 9392 15436 9401
rect 16396 9503 16448 9512
rect 16396 9469 16405 9503
rect 16405 9469 16439 9503
rect 16439 9469 16448 9503
rect 16396 9460 16448 9469
rect 22376 9639 22428 9648
rect 22376 9605 22385 9639
rect 22385 9605 22419 9639
rect 22419 9605 22428 9639
rect 25136 9664 25188 9716
rect 25504 9707 25556 9716
rect 25504 9673 25513 9707
rect 25513 9673 25547 9707
rect 25547 9673 25556 9707
rect 25504 9664 25556 9673
rect 22376 9596 22428 9605
rect 18696 9503 18748 9512
rect 18696 9469 18705 9503
rect 18705 9469 18739 9503
rect 18739 9469 18748 9503
rect 18696 9460 18748 9469
rect 19524 9460 19576 9512
rect 20996 9503 21048 9512
rect 20996 9469 21005 9503
rect 21005 9469 21039 9503
rect 21039 9469 21048 9503
rect 20996 9460 21048 9469
rect 22100 9460 22152 9512
rect 22652 9460 22704 9512
rect 27068 9639 27120 9648
rect 27068 9605 27077 9639
rect 27077 9605 27111 9639
rect 27111 9605 27120 9639
rect 27068 9596 27120 9605
rect 23572 9571 23624 9580
rect 23572 9537 23581 9571
rect 23581 9537 23615 9571
rect 23615 9537 23624 9571
rect 23572 9528 23624 9537
rect 24124 9528 24176 9580
rect 24308 9528 24360 9580
rect 16948 9392 17000 9444
rect 15016 9367 15068 9376
rect 15016 9333 15025 9367
rect 15025 9333 15059 9367
rect 15059 9333 15068 9367
rect 15016 9324 15068 9333
rect 15752 9324 15804 9376
rect 15936 9324 15988 9376
rect 18788 9367 18840 9376
rect 18788 9333 18797 9367
rect 18797 9333 18831 9367
rect 18831 9333 18840 9367
rect 18788 9324 18840 9333
rect 19616 9324 19668 9376
rect 19984 9392 20036 9444
rect 21916 9392 21968 9444
rect 24676 9460 24728 9512
rect 25044 9503 25096 9512
rect 25044 9469 25053 9503
rect 25053 9469 25087 9503
rect 25087 9469 25096 9503
rect 25044 9460 25096 9469
rect 25136 9503 25188 9512
rect 25136 9469 25145 9503
rect 25145 9469 25179 9503
rect 25179 9469 25188 9503
rect 25136 9460 25188 9469
rect 25228 9503 25280 9512
rect 25228 9469 25237 9503
rect 25237 9469 25271 9503
rect 25271 9469 25280 9503
rect 25228 9460 25280 9469
rect 25596 9460 25648 9512
rect 26240 9460 26292 9512
rect 24952 9392 25004 9444
rect 21364 9324 21416 9376
rect 22192 9324 22244 9376
rect 24676 9324 24728 9376
rect 25780 9392 25832 9444
rect 25136 9324 25188 9376
rect 26056 9324 26108 9376
rect 7114 9222 7166 9274
rect 7178 9222 7230 9274
rect 7242 9222 7294 9274
rect 7306 9222 7358 9274
rect 7370 9222 7422 9274
rect 13830 9222 13882 9274
rect 13894 9222 13946 9274
rect 13958 9222 14010 9274
rect 14022 9222 14074 9274
rect 14086 9222 14138 9274
rect 20546 9222 20598 9274
rect 20610 9222 20662 9274
rect 20674 9222 20726 9274
rect 20738 9222 20790 9274
rect 20802 9222 20854 9274
rect 27262 9222 27314 9274
rect 27326 9222 27378 9274
rect 27390 9222 27442 9274
rect 27454 9222 27506 9274
rect 27518 9222 27570 9274
rect 1400 9120 1452 9172
rect 4160 9120 4212 9172
rect 2688 9095 2740 9104
rect 2688 9061 2715 9095
rect 2715 9061 2740 9095
rect 2688 9052 2740 9061
rect 2872 9095 2924 9104
rect 2872 9061 2881 9095
rect 2881 9061 2915 9095
rect 2915 9061 2924 9095
rect 2872 9052 2924 9061
rect 1124 9027 1176 9036
rect 1124 8993 1158 9027
rect 1158 8993 1176 9027
rect 1124 8984 1176 8993
rect 2320 8984 2372 9036
rect 1952 8916 2004 8968
rect 2136 8848 2188 8900
rect 2780 8848 2832 8900
rect 2964 8959 3016 8968
rect 2964 8925 2973 8959
rect 2973 8925 3007 8959
rect 3007 8925 3016 8959
rect 2964 8916 3016 8925
rect 3148 9027 3200 9036
rect 3148 8993 3160 9027
rect 3160 8993 3194 9027
rect 3194 8993 3200 9027
rect 12164 9120 12216 9172
rect 13544 9120 13596 9172
rect 14188 9120 14240 9172
rect 19984 9163 20036 9172
rect 19984 9129 19993 9163
rect 19993 9129 20027 9163
rect 20027 9129 20036 9163
rect 19984 9120 20036 9129
rect 22652 9163 22704 9172
rect 22652 9129 22661 9163
rect 22661 9129 22695 9163
rect 22695 9129 22704 9163
rect 22652 9120 22704 9129
rect 3148 8984 3200 8993
rect 7472 8984 7524 9036
rect 8024 8984 8076 9036
rect 7012 8916 7064 8968
rect 8668 8916 8720 8968
rect 9036 9027 9088 9036
rect 9036 8993 9045 9027
rect 9045 8993 9079 9027
rect 9079 8993 9088 9027
rect 9036 8984 9088 8993
rect 9220 8984 9272 9036
rect 10876 9052 10928 9104
rect 11336 9052 11388 9104
rect 10324 8984 10376 9036
rect 9312 8916 9364 8968
rect 7840 8848 7892 8900
rect 9588 8848 9640 8900
rect 12808 9027 12860 9036
rect 12808 8993 12817 9027
rect 12817 8993 12851 9027
rect 12851 8993 12860 9027
rect 12808 8984 12860 8993
rect 13084 9027 13136 9036
rect 13084 8993 13093 9027
rect 13093 8993 13127 9027
rect 13127 8993 13136 9027
rect 13084 8984 13136 8993
rect 15016 9052 15068 9104
rect 15384 9052 15436 9104
rect 16304 9052 16356 9104
rect 18696 9052 18748 9104
rect 14188 8984 14240 9036
rect 14372 9027 14424 9036
rect 14372 8993 14381 9027
rect 14381 8993 14415 9027
rect 14415 8993 14424 9027
rect 14372 8984 14424 8993
rect 13176 8916 13228 8968
rect 15660 9027 15712 9036
rect 15660 8993 15669 9027
rect 15669 8993 15703 9027
rect 15703 8993 15712 9027
rect 15660 8984 15712 8993
rect 15844 9027 15896 9036
rect 15844 8993 15853 9027
rect 15853 8993 15887 9027
rect 15887 8993 15896 9027
rect 15844 8984 15896 8993
rect 15936 9027 15988 9036
rect 15936 8993 15945 9027
rect 15945 8993 15979 9027
rect 15979 8993 15988 9027
rect 15936 8984 15988 8993
rect 17592 8984 17644 9036
rect 19616 9052 19668 9104
rect 20168 9027 20220 9036
rect 20168 8993 20177 9027
rect 20177 8993 20211 9027
rect 20211 8993 20220 9027
rect 20168 8984 20220 8993
rect 20444 9027 20496 9036
rect 20444 8993 20453 9027
rect 20453 8993 20487 9027
rect 20487 8993 20496 9027
rect 20444 8984 20496 8993
rect 20996 9052 21048 9104
rect 21272 9052 21324 9104
rect 22008 9052 22060 9104
rect 21364 8984 21416 9036
rect 21824 8984 21876 9036
rect 23756 9027 23808 9036
rect 23756 8993 23774 9027
rect 23774 8993 23808 9027
rect 23756 8984 23808 8993
rect 2504 8823 2556 8832
rect 2504 8789 2513 8823
rect 2513 8789 2547 8823
rect 2547 8789 2556 8823
rect 2504 8780 2556 8789
rect 2596 8780 2648 8832
rect 3056 8780 3108 8832
rect 8300 8780 8352 8832
rect 10232 8780 10284 8832
rect 12348 8823 12400 8832
rect 12348 8789 12357 8823
rect 12357 8789 12391 8823
rect 12391 8789 12400 8823
rect 12348 8780 12400 8789
rect 12440 8780 12492 8832
rect 15752 8916 15804 8968
rect 16764 8916 16816 8968
rect 17040 8959 17092 8968
rect 17040 8925 17049 8959
rect 17049 8925 17083 8959
rect 17083 8925 17092 8959
rect 17040 8916 17092 8925
rect 19064 8916 19116 8968
rect 19248 8916 19300 8968
rect 19432 8916 19484 8968
rect 19892 8959 19944 8968
rect 19892 8925 19901 8959
rect 19901 8925 19935 8959
rect 19935 8925 19944 8959
rect 19892 8916 19944 8925
rect 20076 8916 20128 8968
rect 24124 9027 24176 9036
rect 24124 8993 24133 9027
rect 24133 8993 24167 9027
rect 24167 8993 24176 9027
rect 24124 8984 24176 8993
rect 24308 9027 24360 9036
rect 24308 8993 24317 9027
rect 24317 8993 24351 9027
rect 24351 8993 24360 9027
rect 24308 8984 24360 8993
rect 24584 9120 24636 9172
rect 25136 9120 25188 9172
rect 25780 9120 25832 9172
rect 25964 9120 26016 9172
rect 24860 9052 24912 9104
rect 25228 9052 25280 9104
rect 20812 8848 20864 8900
rect 16856 8780 16908 8832
rect 18880 8780 18932 8832
rect 19892 8780 19944 8832
rect 24676 8916 24728 8968
rect 26148 8984 26200 9036
rect 26240 9027 26292 9036
rect 26240 8993 26249 9027
rect 26249 8993 26283 9027
rect 26283 8993 26292 9027
rect 26240 8984 26292 8993
rect 26884 8984 26936 9036
rect 24124 8780 24176 8832
rect 24952 8780 25004 8832
rect 26056 8848 26108 8900
rect 26424 8780 26476 8832
rect 3756 8678 3808 8730
rect 3820 8678 3872 8730
rect 3884 8678 3936 8730
rect 3948 8678 4000 8730
rect 4012 8678 4064 8730
rect 10472 8678 10524 8730
rect 10536 8678 10588 8730
rect 10600 8678 10652 8730
rect 10664 8678 10716 8730
rect 10728 8678 10780 8730
rect 17188 8678 17240 8730
rect 17252 8678 17304 8730
rect 17316 8678 17368 8730
rect 17380 8678 17432 8730
rect 17444 8678 17496 8730
rect 23904 8678 23956 8730
rect 23968 8678 24020 8730
rect 24032 8678 24084 8730
rect 24096 8678 24148 8730
rect 24160 8678 24212 8730
rect 1124 8619 1176 8628
rect 1124 8585 1133 8619
rect 1133 8585 1167 8619
rect 1167 8585 1176 8619
rect 1124 8576 1176 8585
rect 2596 8576 2648 8628
rect 2780 8619 2832 8628
rect 2780 8585 2789 8619
rect 2789 8585 2823 8619
rect 2823 8585 2832 8619
rect 2780 8576 2832 8585
rect 3240 8576 3292 8628
rect 3056 8508 3108 8560
rect 2504 8440 2556 8492
rect 5080 8576 5132 8628
rect 6552 8508 6604 8560
rect 8484 8508 8536 8560
rect 11152 8576 11204 8628
rect 11704 8619 11756 8628
rect 11704 8585 11713 8619
rect 11713 8585 11747 8619
rect 11747 8585 11756 8619
rect 11704 8576 11756 8585
rect 13084 8576 13136 8628
rect 14188 8619 14240 8628
rect 14188 8585 14197 8619
rect 14197 8585 14231 8619
rect 14231 8585 14240 8619
rect 14188 8576 14240 8585
rect 10508 8508 10560 8560
rect 13728 8508 13780 8560
rect 2136 8415 2188 8424
rect 2136 8381 2145 8415
rect 2145 8381 2179 8415
rect 2179 8381 2188 8415
rect 2136 8372 2188 8381
rect 2596 8372 2648 8424
rect 3056 8415 3108 8424
rect 3056 8381 3065 8415
rect 3065 8381 3099 8415
rect 3099 8381 3108 8415
rect 3056 8372 3108 8381
rect 4160 8372 4212 8424
rect 4896 8415 4948 8424
rect 4896 8381 4905 8415
rect 4905 8381 4939 8415
rect 4939 8381 4948 8415
rect 4896 8372 4948 8381
rect 9312 8440 9364 8492
rect 13636 8440 13688 8492
rect 2688 8304 2740 8356
rect 4252 8304 4304 8356
rect 5816 8304 5868 8356
rect 6920 8372 6972 8424
rect 9588 8372 9640 8424
rect 10600 8372 10652 8424
rect 10232 8304 10284 8356
rect 10324 8304 10376 8356
rect 10508 8347 10560 8356
rect 10508 8313 10517 8347
rect 10517 8313 10551 8347
rect 10551 8313 10560 8347
rect 10508 8304 10560 8313
rect 7012 8236 7064 8288
rect 8024 8236 8076 8288
rect 11152 8304 11204 8356
rect 11888 8347 11940 8356
rect 11888 8313 11915 8347
rect 11915 8313 11940 8347
rect 11888 8304 11940 8313
rect 12256 8372 12308 8424
rect 12348 8372 12400 8424
rect 12992 8372 13044 8424
rect 15108 8508 15160 8560
rect 14648 8440 14700 8492
rect 16948 8440 17000 8492
rect 14832 8372 14884 8424
rect 14280 8304 14332 8356
rect 15292 8415 15344 8424
rect 15292 8381 15301 8415
rect 15301 8381 15335 8415
rect 15335 8381 15344 8415
rect 15292 8372 15344 8381
rect 15384 8417 15436 8424
rect 15384 8383 15393 8417
rect 15393 8383 15427 8417
rect 15427 8383 15436 8417
rect 15384 8372 15436 8383
rect 15568 8415 15620 8424
rect 15568 8381 15577 8415
rect 15577 8381 15611 8415
rect 15611 8381 15620 8415
rect 15568 8372 15620 8381
rect 16488 8415 16540 8424
rect 16488 8381 16497 8415
rect 16497 8381 16531 8415
rect 16531 8381 16540 8415
rect 16488 8372 16540 8381
rect 17592 8576 17644 8628
rect 18696 8576 18748 8628
rect 19524 8619 19576 8628
rect 19524 8585 19533 8619
rect 19533 8585 19567 8619
rect 19567 8585 19576 8619
rect 19524 8576 19576 8585
rect 20444 8576 20496 8628
rect 22560 8576 22612 8628
rect 17960 8508 18012 8560
rect 19248 8508 19300 8560
rect 19432 8440 19484 8492
rect 20168 8440 20220 8492
rect 18696 8415 18748 8424
rect 18696 8381 18705 8415
rect 18705 8381 18739 8415
rect 18739 8381 18748 8415
rect 18696 8372 18748 8381
rect 18880 8415 18932 8424
rect 18880 8381 18889 8415
rect 18889 8381 18923 8415
rect 18923 8381 18932 8415
rect 18880 8372 18932 8381
rect 19064 8372 19116 8424
rect 14372 8279 14424 8288
rect 14372 8245 14381 8279
rect 14381 8245 14415 8279
rect 14415 8245 14424 8279
rect 14372 8236 14424 8245
rect 14740 8236 14792 8288
rect 18328 8347 18380 8356
rect 18328 8313 18337 8347
rect 18337 8313 18371 8347
rect 18371 8313 18380 8347
rect 18328 8304 18380 8313
rect 19616 8415 19668 8424
rect 19616 8381 19625 8415
rect 19625 8381 19659 8415
rect 19659 8381 19668 8415
rect 19616 8372 19668 8381
rect 19892 8372 19944 8424
rect 20076 8415 20128 8424
rect 20076 8381 20085 8415
rect 20085 8381 20119 8415
rect 20119 8381 20128 8415
rect 20076 8372 20128 8381
rect 20812 8415 20864 8424
rect 20812 8381 20821 8415
rect 20821 8381 20855 8415
rect 20855 8381 20864 8415
rect 20812 8372 20864 8381
rect 24032 8440 24084 8492
rect 21640 8372 21692 8424
rect 21732 8415 21784 8424
rect 21732 8381 21741 8415
rect 21741 8381 21775 8415
rect 21775 8381 21784 8415
rect 21732 8372 21784 8381
rect 23388 8415 23440 8424
rect 23388 8381 23397 8415
rect 23397 8381 23431 8415
rect 23431 8381 23440 8415
rect 23388 8372 23440 8381
rect 21824 8304 21876 8356
rect 24400 8372 24452 8424
rect 24952 8415 25004 8424
rect 24952 8381 24970 8415
rect 24970 8381 25004 8415
rect 24952 8372 25004 8381
rect 25596 8415 25648 8424
rect 23572 8347 23624 8356
rect 23572 8313 23581 8347
rect 23581 8313 23615 8347
rect 23615 8313 23624 8347
rect 23572 8304 23624 8313
rect 24124 8304 24176 8356
rect 25044 8304 25096 8356
rect 25596 8381 25605 8415
rect 25605 8381 25639 8415
rect 25639 8381 25648 8415
rect 25596 8372 25648 8381
rect 25688 8304 25740 8356
rect 16396 8236 16448 8288
rect 21364 8279 21416 8288
rect 21364 8245 21373 8279
rect 21373 8245 21407 8279
rect 21407 8245 21416 8279
rect 21364 8236 21416 8245
rect 21548 8236 21600 8288
rect 23480 8236 23532 8288
rect 24768 8236 24820 8288
rect 25320 8236 25372 8288
rect 26884 8236 26936 8288
rect 7114 8134 7166 8186
rect 7178 8134 7230 8186
rect 7242 8134 7294 8186
rect 7306 8134 7358 8186
rect 7370 8134 7422 8186
rect 13830 8134 13882 8186
rect 13894 8134 13946 8186
rect 13958 8134 14010 8186
rect 14022 8134 14074 8186
rect 14086 8134 14138 8186
rect 20546 8134 20598 8186
rect 20610 8134 20662 8186
rect 20674 8134 20726 8186
rect 20738 8134 20790 8186
rect 20802 8134 20854 8186
rect 27262 8134 27314 8186
rect 27326 8134 27378 8186
rect 27390 8134 27442 8186
rect 27454 8134 27506 8186
rect 27518 8134 27570 8186
rect 10508 8032 10560 8084
rect 10600 8075 10652 8084
rect 10600 8041 10609 8075
rect 10609 8041 10643 8075
rect 10643 8041 10652 8075
rect 10600 8032 10652 8041
rect 3148 7896 3200 7948
rect 4896 7964 4948 8016
rect 4436 7939 4488 7948
rect 4436 7905 4445 7939
rect 4445 7905 4479 7939
rect 4479 7905 4488 7939
rect 4436 7896 4488 7905
rect 6000 7939 6052 7948
rect 6000 7905 6009 7939
rect 6009 7905 6043 7939
rect 6043 7905 6052 7939
rect 6000 7896 6052 7905
rect 6644 8007 6696 8016
rect 6644 7973 6653 8007
rect 6653 7973 6687 8007
rect 6687 7973 6696 8007
rect 6644 7964 6696 7973
rect 7012 7964 7064 8016
rect 3240 7828 3292 7880
rect 4252 7803 4304 7812
rect 4252 7769 4261 7803
rect 4261 7769 4295 7803
rect 4295 7769 4304 7803
rect 4252 7760 4304 7769
rect 5816 7803 5868 7812
rect 5816 7769 5825 7803
rect 5825 7769 5859 7803
rect 5859 7769 5868 7803
rect 5816 7760 5868 7769
rect 6276 7803 6328 7812
rect 6276 7769 6285 7803
rect 6285 7769 6319 7803
rect 6319 7769 6328 7803
rect 6276 7760 6328 7769
rect 6920 7760 6972 7812
rect 8852 7803 8904 7812
rect 8852 7769 8861 7803
rect 8861 7769 8895 7803
rect 8895 7769 8904 7803
rect 8852 7760 8904 7769
rect 1124 7692 1176 7744
rect 2872 7692 2924 7744
rect 8116 7692 8168 7744
rect 8208 7692 8260 7744
rect 9312 7896 9364 7948
rect 9772 7896 9824 7948
rect 9128 7871 9180 7880
rect 9128 7837 9137 7871
rect 9137 7837 9171 7871
rect 9171 7837 9180 7871
rect 9128 7828 9180 7837
rect 10876 7896 10928 7948
rect 12348 7871 12400 7880
rect 12348 7837 12357 7871
rect 12357 7837 12391 7871
rect 12391 7837 12400 7871
rect 12348 7828 12400 7837
rect 12256 7760 12308 7812
rect 13176 7964 13228 8016
rect 14280 7964 14332 8016
rect 13636 7939 13688 7948
rect 13636 7905 13645 7939
rect 13645 7905 13679 7939
rect 13679 7905 13688 7939
rect 13636 7896 13688 7905
rect 13912 7939 13964 7948
rect 13912 7905 13946 7939
rect 13946 7905 13964 7939
rect 13912 7896 13964 7905
rect 15108 7939 15160 7948
rect 15108 7905 15117 7939
rect 15117 7905 15151 7939
rect 15151 7905 15160 7939
rect 15108 7896 15160 7905
rect 15292 7939 15344 7948
rect 15292 7905 15301 7939
rect 15301 7905 15335 7939
rect 15335 7905 15344 7939
rect 15292 7896 15344 7905
rect 15568 7939 15620 7948
rect 15568 7905 15577 7939
rect 15577 7905 15611 7939
rect 15611 7905 15620 7939
rect 15568 7896 15620 7905
rect 15660 7896 15712 7948
rect 17040 7964 17092 8016
rect 16396 7939 16448 7948
rect 16396 7905 16430 7939
rect 16430 7905 16448 7939
rect 16396 7896 16448 7905
rect 18328 8032 18380 8084
rect 20904 8032 20956 8084
rect 21916 7964 21968 8016
rect 13176 7871 13228 7880
rect 13176 7837 13185 7871
rect 13185 7837 13219 7871
rect 13219 7837 13228 7871
rect 13176 7828 13228 7837
rect 13360 7871 13412 7880
rect 13360 7837 13369 7871
rect 13369 7837 13403 7871
rect 13403 7837 13412 7871
rect 13360 7828 13412 7837
rect 17684 7871 17736 7880
rect 17684 7837 17693 7871
rect 17693 7837 17727 7871
rect 17727 7837 17736 7871
rect 17684 7828 17736 7837
rect 18788 7871 18840 7880
rect 18788 7837 18797 7871
rect 18797 7837 18831 7871
rect 18831 7837 18840 7871
rect 18788 7828 18840 7837
rect 19616 7939 19668 7948
rect 19616 7905 19625 7939
rect 19625 7905 19659 7939
rect 19659 7905 19668 7939
rect 19616 7896 19668 7905
rect 14740 7760 14792 7812
rect 15476 7760 15528 7812
rect 11336 7735 11388 7744
rect 11336 7701 11345 7735
rect 11345 7701 11379 7735
rect 11379 7701 11388 7735
rect 11336 7692 11388 7701
rect 12072 7692 12124 7744
rect 14004 7692 14056 7744
rect 14556 7692 14608 7744
rect 17776 7692 17828 7744
rect 18144 7760 18196 7812
rect 19708 7828 19760 7880
rect 20076 7896 20128 7948
rect 20260 7896 20312 7948
rect 19984 7828 20036 7880
rect 19524 7760 19576 7812
rect 20904 7939 20956 7948
rect 20904 7905 20913 7939
rect 20913 7905 20947 7939
rect 20947 7905 20956 7939
rect 20904 7896 20956 7905
rect 21364 7896 21416 7948
rect 21548 7939 21600 7948
rect 21548 7905 21582 7939
rect 21582 7905 21600 7939
rect 21548 7896 21600 7905
rect 23020 8032 23072 8084
rect 24032 8075 24084 8084
rect 24032 8041 24041 8075
rect 24041 8041 24075 8075
rect 24075 8041 24084 8075
rect 24032 8032 24084 8041
rect 24308 8032 24360 8084
rect 24860 8075 24912 8084
rect 24860 8041 24869 8075
rect 24869 8041 24903 8075
rect 24903 8041 24912 8075
rect 24860 8032 24912 8041
rect 25688 8032 25740 8084
rect 21272 7871 21324 7880
rect 21272 7837 21281 7871
rect 21281 7837 21315 7871
rect 21315 7837 21324 7871
rect 21272 7828 21324 7837
rect 23388 7896 23440 7948
rect 23480 7939 23532 7948
rect 23480 7905 23489 7939
rect 23489 7905 23523 7939
rect 23523 7905 23532 7939
rect 23480 7896 23532 7905
rect 23572 7896 23624 7948
rect 24124 7964 24176 8016
rect 24492 7964 24544 8016
rect 25320 7964 25372 8016
rect 24032 7939 24084 7948
rect 24032 7905 24041 7939
rect 24041 7905 24075 7939
rect 24075 7905 24084 7939
rect 24032 7896 24084 7905
rect 24768 7896 24820 7948
rect 25872 7939 25924 7948
rect 25872 7905 25881 7939
rect 25881 7905 25915 7939
rect 25915 7905 25924 7939
rect 25872 7896 25924 7905
rect 26056 8032 26108 8084
rect 26424 8075 26476 8084
rect 26424 8041 26433 8075
rect 26433 8041 26467 8075
rect 26467 8041 26476 8075
rect 26424 8032 26476 8041
rect 26240 7939 26292 7948
rect 26240 7905 26249 7939
rect 26249 7905 26283 7939
rect 26283 7905 26292 7939
rect 26240 7896 26292 7905
rect 27068 7939 27120 7948
rect 27068 7905 27077 7939
rect 27077 7905 27111 7939
rect 27111 7905 27120 7939
rect 27068 7896 27120 7905
rect 26792 7828 26844 7880
rect 20904 7760 20956 7812
rect 18420 7692 18472 7744
rect 18880 7692 18932 7744
rect 21916 7692 21968 7744
rect 3756 7590 3808 7642
rect 3820 7590 3872 7642
rect 3884 7590 3936 7642
rect 3948 7590 4000 7642
rect 4012 7590 4064 7642
rect 10472 7590 10524 7642
rect 10536 7590 10588 7642
rect 10600 7590 10652 7642
rect 10664 7590 10716 7642
rect 10728 7590 10780 7642
rect 17188 7590 17240 7642
rect 17252 7590 17304 7642
rect 17316 7590 17368 7642
rect 17380 7590 17432 7642
rect 17444 7590 17496 7642
rect 23904 7590 23956 7642
rect 23968 7590 24020 7642
rect 24032 7590 24084 7642
rect 24096 7590 24148 7642
rect 24160 7590 24212 7642
rect 2136 7488 2188 7540
rect 2596 7531 2648 7540
rect 2596 7497 2605 7531
rect 2605 7497 2639 7531
rect 2639 7497 2648 7531
rect 2596 7488 2648 7497
rect 3240 7531 3292 7540
rect 3240 7497 3249 7531
rect 3249 7497 3283 7531
rect 3283 7497 3292 7531
rect 3240 7488 3292 7497
rect 4436 7531 4488 7540
rect 4436 7497 4445 7531
rect 4445 7497 4479 7531
rect 4479 7497 4488 7531
rect 4436 7488 4488 7497
rect 6000 7488 6052 7540
rect 6644 7488 6696 7540
rect 9128 7488 9180 7540
rect 9588 7488 9640 7540
rect 10232 7488 10284 7540
rect 8024 7420 8076 7472
rect 8852 7420 8904 7472
rect 3332 7352 3384 7404
rect 4896 7352 4948 7404
rect 1400 7284 1452 7336
rect 1676 7284 1728 7336
rect 2596 7284 2648 7336
rect 3516 7327 3568 7336
rect 3516 7293 3525 7327
rect 3525 7293 3559 7327
rect 3559 7293 3568 7327
rect 3516 7284 3568 7293
rect 1124 7259 1176 7268
rect 1124 7225 1158 7259
rect 1158 7225 1176 7259
rect 1124 7216 1176 7225
rect 3240 7216 3292 7268
rect 4068 7259 4120 7268
rect 4068 7225 4077 7259
rect 4077 7225 4111 7259
rect 4111 7225 4120 7259
rect 4068 7216 4120 7225
rect 2228 7191 2280 7200
rect 2228 7157 2237 7191
rect 2237 7157 2271 7191
rect 2271 7157 2280 7191
rect 2228 7148 2280 7157
rect 4252 7191 4304 7200
rect 4252 7157 4277 7191
rect 4277 7157 4304 7191
rect 4620 7284 4672 7336
rect 4804 7327 4856 7336
rect 4804 7293 4813 7327
rect 4813 7293 4847 7327
rect 4847 7293 4856 7327
rect 4804 7284 4856 7293
rect 4988 7327 5040 7336
rect 4988 7293 4997 7327
rect 4997 7293 5031 7327
rect 5031 7293 5040 7327
rect 4988 7284 5040 7293
rect 6276 7352 6328 7404
rect 6000 7284 6052 7336
rect 6460 7327 6512 7336
rect 6460 7293 6469 7327
rect 6469 7293 6503 7327
rect 6503 7293 6512 7327
rect 6460 7284 6512 7293
rect 6920 7352 6972 7404
rect 6736 7284 6788 7336
rect 6828 7327 6880 7336
rect 6828 7293 6837 7327
rect 6837 7293 6871 7327
rect 6871 7293 6880 7327
rect 6828 7284 6880 7293
rect 7656 7352 7708 7404
rect 9404 7352 9456 7404
rect 4252 7148 4304 7157
rect 4712 7148 4764 7200
rect 5908 7191 5960 7200
rect 5908 7157 5917 7191
rect 5917 7157 5951 7191
rect 5951 7157 5960 7191
rect 5908 7148 5960 7157
rect 7748 7216 7800 7268
rect 8208 7327 8260 7336
rect 8208 7293 8217 7327
rect 8217 7293 8251 7327
rect 8251 7293 8260 7327
rect 8208 7284 8260 7293
rect 8576 7259 8628 7268
rect 7012 7148 7064 7200
rect 7840 7148 7892 7200
rect 8576 7225 8585 7259
rect 8585 7225 8619 7259
rect 8619 7225 8628 7259
rect 8576 7216 8628 7225
rect 9680 7327 9732 7336
rect 9680 7293 9689 7327
rect 9689 7293 9723 7327
rect 9723 7293 9732 7327
rect 9680 7284 9732 7293
rect 9772 7327 9824 7336
rect 9772 7293 9781 7327
rect 9781 7293 9815 7327
rect 9815 7293 9824 7327
rect 9772 7284 9824 7293
rect 13176 7488 13228 7540
rect 12256 7420 12308 7472
rect 13912 7488 13964 7540
rect 14188 7488 14240 7540
rect 15660 7531 15712 7540
rect 15660 7497 15669 7531
rect 15669 7497 15703 7531
rect 15703 7497 15712 7531
rect 15660 7488 15712 7497
rect 16304 7488 16356 7540
rect 16488 7488 16540 7540
rect 11336 7284 11388 7336
rect 14004 7395 14056 7404
rect 14004 7361 14013 7395
rect 14013 7361 14047 7395
rect 14047 7361 14056 7395
rect 14004 7352 14056 7361
rect 12072 7327 12124 7336
rect 12072 7293 12081 7327
rect 12081 7293 12115 7327
rect 12115 7293 12124 7327
rect 12072 7284 12124 7293
rect 12532 7327 12584 7336
rect 12532 7293 12541 7327
rect 12541 7293 12575 7327
rect 12575 7293 12584 7327
rect 12532 7284 12584 7293
rect 14556 7352 14608 7404
rect 12348 7216 12400 7268
rect 9680 7148 9732 7200
rect 10324 7191 10376 7200
rect 10324 7157 10333 7191
rect 10333 7157 10367 7191
rect 10367 7157 10376 7191
rect 10324 7148 10376 7157
rect 11336 7148 11388 7200
rect 11704 7148 11756 7200
rect 14372 7284 14424 7336
rect 15016 7327 15068 7336
rect 15016 7293 15025 7327
rect 15025 7293 15059 7327
rect 15059 7293 15068 7327
rect 15016 7284 15068 7293
rect 15200 7284 15252 7336
rect 15568 7284 15620 7336
rect 16948 7327 17000 7336
rect 16948 7293 16957 7327
rect 16957 7293 16991 7327
rect 16991 7293 17000 7327
rect 16948 7284 17000 7293
rect 17040 7327 17092 7336
rect 17040 7293 17049 7327
rect 17049 7293 17083 7327
rect 17083 7293 17092 7327
rect 17040 7284 17092 7293
rect 17132 7327 17184 7336
rect 17132 7293 17141 7327
rect 17141 7293 17175 7327
rect 17175 7293 17184 7327
rect 17132 7284 17184 7293
rect 18420 7488 18472 7540
rect 17868 7420 17920 7472
rect 17960 7420 18012 7472
rect 18880 7531 18932 7540
rect 18880 7497 18889 7531
rect 18889 7497 18923 7531
rect 18923 7497 18932 7531
rect 18880 7488 18932 7497
rect 19524 7531 19576 7540
rect 19524 7497 19533 7531
rect 19533 7497 19567 7531
rect 19567 7497 19576 7531
rect 19524 7488 19576 7497
rect 20904 7488 20956 7540
rect 21640 7531 21692 7540
rect 21640 7497 21649 7531
rect 21649 7497 21683 7531
rect 21683 7497 21692 7531
rect 21640 7488 21692 7497
rect 21732 7531 21784 7540
rect 21732 7497 21741 7531
rect 21741 7497 21775 7531
rect 21775 7497 21784 7531
rect 21732 7488 21784 7497
rect 25872 7488 25924 7540
rect 18788 7352 18840 7404
rect 19616 7420 19668 7472
rect 16672 7216 16724 7268
rect 18144 7327 18196 7336
rect 18144 7293 18153 7327
rect 18153 7293 18187 7327
rect 18187 7293 18196 7327
rect 18144 7284 18196 7293
rect 18236 7327 18288 7336
rect 18236 7293 18245 7327
rect 18245 7293 18279 7327
rect 18279 7293 18288 7327
rect 18236 7284 18288 7293
rect 19708 7327 19760 7336
rect 17776 7216 17828 7268
rect 19708 7293 19717 7327
rect 19717 7293 19751 7327
rect 19751 7293 19760 7327
rect 19708 7284 19760 7293
rect 19984 7327 20036 7336
rect 19984 7293 19993 7327
rect 19993 7293 20027 7327
rect 20027 7293 20036 7327
rect 19984 7284 20036 7293
rect 20076 7284 20128 7336
rect 21916 7395 21968 7404
rect 21916 7361 21925 7395
rect 21925 7361 21959 7395
rect 21959 7361 21968 7395
rect 21916 7352 21968 7361
rect 26884 7395 26936 7404
rect 26884 7361 26893 7395
rect 26893 7361 26927 7395
rect 26927 7361 26936 7395
rect 26884 7352 26936 7361
rect 22008 7327 22060 7336
rect 13084 7148 13136 7200
rect 16212 7191 16264 7200
rect 16212 7157 16221 7191
rect 16221 7157 16255 7191
rect 16255 7157 16264 7191
rect 16212 7148 16264 7157
rect 19064 7259 19116 7268
rect 19064 7225 19073 7259
rect 19073 7225 19107 7259
rect 19107 7225 19116 7259
rect 19064 7216 19116 7225
rect 21180 7216 21232 7268
rect 22008 7293 22017 7327
rect 22017 7293 22051 7327
rect 22051 7293 22060 7327
rect 22008 7284 22060 7293
rect 23020 7284 23072 7336
rect 23296 7327 23348 7336
rect 23296 7293 23305 7327
rect 23305 7293 23339 7327
rect 23339 7293 23348 7327
rect 23296 7284 23348 7293
rect 23572 7327 23624 7336
rect 23572 7293 23581 7327
rect 23581 7293 23615 7327
rect 23615 7293 23624 7327
rect 23572 7284 23624 7293
rect 24584 7284 24636 7336
rect 19524 7148 19576 7200
rect 23756 7216 23808 7268
rect 21916 7148 21968 7200
rect 22560 7148 22612 7200
rect 25044 7216 25096 7268
rect 26056 7191 26108 7200
rect 26056 7157 26065 7191
rect 26065 7157 26099 7191
rect 26099 7157 26108 7191
rect 26056 7148 26108 7157
rect 7114 7046 7166 7098
rect 7178 7046 7230 7098
rect 7242 7046 7294 7098
rect 7306 7046 7358 7098
rect 7370 7046 7422 7098
rect 13830 7046 13882 7098
rect 13894 7046 13946 7098
rect 13958 7046 14010 7098
rect 14022 7046 14074 7098
rect 14086 7046 14138 7098
rect 20546 7046 20598 7098
rect 20610 7046 20662 7098
rect 20674 7046 20726 7098
rect 20738 7046 20790 7098
rect 20802 7046 20854 7098
rect 27262 7046 27314 7098
rect 27326 7046 27378 7098
rect 27390 7046 27442 7098
rect 27454 7046 27506 7098
rect 27518 7046 27570 7098
rect 2136 6987 2188 6996
rect 2136 6953 2145 6987
rect 2145 6953 2179 6987
rect 2179 6953 2188 6987
rect 2136 6944 2188 6953
rect 5908 6944 5960 6996
rect 2596 6876 2648 6928
rect 2136 6808 2188 6860
rect 2228 6851 2280 6860
rect 2228 6817 2237 6851
rect 2237 6817 2271 6851
rect 2271 6817 2280 6851
rect 2228 6808 2280 6817
rect 2688 6740 2740 6792
rect 2964 6851 3016 6860
rect 2964 6817 2973 6851
rect 2973 6817 3007 6851
rect 3007 6817 3016 6851
rect 2964 6808 3016 6817
rect 3332 6919 3384 6928
rect 3332 6885 3341 6919
rect 3341 6885 3375 6919
rect 3375 6885 3384 6919
rect 3332 6876 3384 6885
rect 3240 6851 3292 6860
rect 3240 6817 3249 6851
rect 3249 6817 3283 6851
rect 3283 6817 3292 6851
rect 3240 6808 3292 6817
rect 3608 6851 3660 6860
rect 3608 6817 3617 6851
rect 3617 6817 3651 6851
rect 3651 6817 3660 6851
rect 3608 6808 3660 6817
rect 4252 6851 4304 6860
rect 4252 6817 4261 6851
rect 4261 6817 4295 6851
rect 4295 6817 4304 6851
rect 4252 6808 4304 6817
rect 4896 6851 4948 6860
rect 4896 6817 4905 6851
rect 4905 6817 4939 6851
rect 4939 6817 4948 6851
rect 4896 6808 4948 6817
rect 4988 6851 5040 6860
rect 4988 6817 4997 6851
rect 4997 6817 5031 6851
rect 5031 6817 5040 6851
rect 4988 6808 5040 6817
rect 5080 6851 5132 6860
rect 5080 6817 5089 6851
rect 5089 6817 5123 6851
rect 5123 6817 5132 6851
rect 5080 6808 5132 6817
rect 5264 6851 5316 6860
rect 5264 6817 5273 6851
rect 5273 6817 5307 6851
rect 5307 6817 5316 6851
rect 5264 6808 5316 6817
rect 6000 6808 6052 6860
rect 6828 6944 6880 6996
rect 6920 6944 6972 6996
rect 7656 6987 7708 6996
rect 7656 6953 7665 6987
rect 7665 6953 7699 6987
rect 7699 6953 7708 6987
rect 7656 6944 7708 6953
rect 3148 6672 3200 6724
rect 4620 6783 4672 6792
rect 4620 6749 4629 6783
rect 4629 6749 4663 6783
rect 4663 6749 4672 6783
rect 4620 6740 4672 6749
rect 4804 6740 4856 6792
rect 6460 6851 6512 6860
rect 6460 6817 6469 6851
rect 6469 6817 6503 6851
rect 6503 6817 6512 6851
rect 6460 6808 6512 6817
rect 7012 6876 7064 6928
rect 11704 6944 11756 6996
rect 12532 6944 12584 6996
rect 13360 6944 13412 6996
rect 16212 6944 16264 6996
rect 8668 6876 8720 6928
rect 6644 6851 6696 6860
rect 6644 6817 6653 6851
rect 6653 6817 6687 6851
rect 6687 6817 6696 6851
rect 6644 6808 6696 6817
rect 6828 6851 6880 6860
rect 6828 6817 6837 6851
rect 6837 6817 6871 6851
rect 6871 6817 6880 6851
rect 6828 6808 6880 6817
rect 9312 6808 9364 6860
rect 11336 6876 11388 6928
rect 19064 6944 19116 6996
rect 19616 6987 19668 6996
rect 19616 6953 19625 6987
rect 19625 6953 19659 6987
rect 19659 6953 19668 6987
rect 19616 6944 19668 6953
rect 19708 6944 19760 6996
rect 24492 6944 24544 6996
rect 17684 6876 17736 6928
rect 11520 6808 11572 6860
rect 12532 6808 12584 6860
rect 13084 6851 13136 6860
rect 13084 6817 13093 6851
rect 13093 6817 13127 6851
rect 13127 6817 13136 6851
rect 13084 6808 13136 6817
rect 6736 6740 6788 6792
rect 12164 6740 12216 6792
rect 12348 6740 12400 6792
rect 14188 6808 14240 6860
rect 16672 6851 16724 6860
rect 16672 6817 16681 6851
rect 16681 6817 16715 6851
rect 16715 6817 16724 6851
rect 16672 6808 16724 6817
rect 16948 6851 17000 6860
rect 16948 6817 16957 6851
rect 16957 6817 16991 6851
rect 16991 6817 17000 6851
rect 16948 6808 17000 6817
rect 17040 6851 17092 6860
rect 17040 6817 17049 6851
rect 17049 6817 17083 6851
rect 17083 6817 17092 6851
rect 17040 6808 17092 6817
rect 17132 6740 17184 6792
rect 17776 6851 17828 6860
rect 17776 6817 17785 6851
rect 17785 6817 17819 6851
rect 17819 6817 17828 6851
rect 17776 6808 17828 6817
rect 17960 6808 18012 6860
rect 18420 6851 18472 6860
rect 18420 6817 18443 6851
rect 18443 6817 18472 6851
rect 18420 6808 18472 6817
rect 21180 6876 21232 6928
rect 21456 6876 21508 6928
rect 22008 6876 22060 6928
rect 20260 6851 20312 6860
rect 17684 6740 17736 6792
rect 18052 6740 18104 6792
rect 18144 6783 18196 6792
rect 18144 6749 18153 6783
rect 18153 6749 18187 6783
rect 18187 6749 18196 6783
rect 18144 6740 18196 6749
rect 20260 6817 20269 6851
rect 20269 6817 20303 6851
rect 20303 6817 20312 6851
rect 20260 6808 20312 6817
rect 23296 6851 23348 6860
rect 23296 6817 23305 6851
rect 23305 6817 23339 6851
rect 23339 6817 23348 6851
rect 23296 6808 23348 6817
rect 23572 6851 23624 6860
rect 23572 6817 23581 6851
rect 23581 6817 23615 6851
rect 23615 6817 23624 6851
rect 23572 6808 23624 6817
rect 23756 6851 23808 6860
rect 23756 6817 23765 6851
rect 23765 6817 23799 6851
rect 23799 6817 23808 6851
rect 23756 6808 23808 6817
rect 7840 6672 7892 6724
rect 3516 6604 3568 6656
rect 7748 6604 7800 6656
rect 9036 6604 9088 6656
rect 14648 6672 14700 6724
rect 17592 6672 17644 6724
rect 24768 6851 24820 6860
rect 24768 6817 24777 6851
rect 24777 6817 24811 6851
rect 24811 6817 24820 6851
rect 24768 6808 24820 6817
rect 25320 6876 25372 6928
rect 25136 6851 25188 6860
rect 25136 6817 25145 6851
rect 25145 6817 25179 6851
rect 25179 6817 25188 6851
rect 25136 6808 25188 6817
rect 25228 6851 25280 6860
rect 25228 6817 25237 6851
rect 25237 6817 25271 6851
rect 25271 6817 25280 6851
rect 25228 6808 25280 6817
rect 25412 6851 25464 6860
rect 25412 6817 25421 6851
rect 25421 6817 25455 6851
rect 25455 6817 25464 6851
rect 25412 6808 25464 6817
rect 26424 6944 26476 6996
rect 25964 6851 26016 6860
rect 25964 6817 25973 6851
rect 25973 6817 26007 6851
rect 26007 6817 26016 6851
rect 25964 6808 26016 6817
rect 26148 6851 26200 6860
rect 26148 6817 26157 6851
rect 26157 6817 26191 6851
rect 26191 6817 26200 6851
rect 26148 6808 26200 6817
rect 26792 6851 26844 6860
rect 26792 6817 26801 6851
rect 26801 6817 26835 6851
rect 26835 6817 26844 6851
rect 26792 6808 26844 6817
rect 12348 6647 12400 6656
rect 12348 6613 12357 6647
rect 12357 6613 12391 6647
rect 12391 6613 12400 6647
rect 12348 6604 12400 6613
rect 13268 6647 13320 6656
rect 13268 6613 13277 6647
rect 13277 6613 13311 6647
rect 13311 6613 13320 6647
rect 13268 6604 13320 6613
rect 18420 6604 18472 6656
rect 22560 6672 22612 6724
rect 23020 6715 23072 6724
rect 23020 6681 23029 6715
rect 23029 6681 23063 6715
rect 23063 6681 23072 6715
rect 23020 6672 23072 6681
rect 25228 6672 25280 6724
rect 21640 6604 21692 6656
rect 24768 6604 24820 6656
rect 25136 6604 25188 6656
rect 25688 6647 25740 6656
rect 25688 6613 25697 6647
rect 25697 6613 25731 6647
rect 25731 6613 25740 6647
rect 25688 6604 25740 6613
rect 3756 6502 3808 6554
rect 3820 6502 3872 6554
rect 3884 6502 3936 6554
rect 3948 6502 4000 6554
rect 4012 6502 4064 6554
rect 10472 6502 10524 6554
rect 10536 6502 10588 6554
rect 10600 6502 10652 6554
rect 10664 6502 10716 6554
rect 10728 6502 10780 6554
rect 17188 6502 17240 6554
rect 17252 6502 17304 6554
rect 17316 6502 17368 6554
rect 17380 6502 17432 6554
rect 17444 6502 17496 6554
rect 23904 6502 23956 6554
rect 23968 6502 24020 6554
rect 24032 6502 24084 6554
rect 24096 6502 24148 6554
rect 24160 6502 24212 6554
rect 4620 6400 4672 6452
rect 6000 6443 6052 6452
rect 6000 6409 6009 6443
rect 6009 6409 6043 6443
rect 6043 6409 6052 6443
rect 6000 6400 6052 6409
rect 9956 6400 10008 6452
rect 11520 6443 11572 6452
rect 11520 6409 11529 6443
rect 11529 6409 11563 6443
rect 11563 6409 11572 6443
rect 11520 6400 11572 6409
rect 3608 6375 3660 6384
rect 3608 6341 3617 6375
rect 3617 6341 3651 6375
rect 3651 6341 3660 6375
rect 3608 6332 3660 6341
rect 5264 6332 5316 6384
rect 9220 6332 9272 6384
rect 3516 6196 3568 6248
rect 4528 6196 4580 6248
rect 4712 6196 4764 6248
rect 5080 6264 5132 6316
rect 4896 6239 4948 6248
rect 4896 6205 4905 6239
rect 4905 6205 4939 6239
rect 4939 6205 4948 6239
rect 4896 6196 4948 6205
rect 5632 6196 5684 6248
rect 6828 6264 6880 6316
rect 2964 6128 3016 6180
rect 3608 6128 3660 6180
rect 4068 6171 4120 6180
rect 4068 6137 4077 6171
rect 4077 6137 4111 6171
rect 4111 6137 4120 6171
rect 4068 6128 4120 6137
rect 6184 6196 6236 6248
rect 7472 6196 7524 6248
rect 8116 6196 8168 6248
rect 6552 6128 6604 6180
rect 7012 6128 7064 6180
rect 3700 6103 3752 6112
rect 3700 6069 3709 6103
rect 3709 6069 3743 6103
rect 3743 6069 3752 6103
rect 3700 6060 3752 6069
rect 8668 6128 8720 6180
rect 9036 6196 9088 6248
rect 10324 6332 10376 6384
rect 9864 6239 9916 6248
rect 9864 6205 9873 6239
rect 9873 6205 9907 6239
rect 9907 6205 9916 6239
rect 9864 6196 9916 6205
rect 9956 6239 10008 6248
rect 9956 6205 9965 6239
rect 9965 6205 9999 6239
rect 9999 6205 10008 6239
rect 9956 6196 10008 6205
rect 10048 6239 10100 6248
rect 10048 6205 10057 6239
rect 10057 6205 10091 6239
rect 10091 6205 10100 6239
rect 10048 6196 10100 6205
rect 10508 6196 10560 6248
rect 12532 6443 12584 6452
rect 12532 6409 12541 6443
rect 12541 6409 12575 6443
rect 12575 6409 12584 6443
rect 12532 6400 12584 6409
rect 16304 6400 16356 6452
rect 23296 6400 23348 6452
rect 24400 6443 24452 6452
rect 24400 6409 24409 6443
rect 24409 6409 24443 6443
rect 24443 6409 24452 6443
rect 24400 6400 24452 6409
rect 24584 6443 24636 6452
rect 24584 6409 24593 6443
rect 24593 6409 24627 6443
rect 24627 6409 24636 6443
rect 24584 6400 24636 6409
rect 25320 6443 25372 6452
rect 25320 6409 25329 6443
rect 25329 6409 25363 6443
rect 25363 6409 25372 6443
rect 25320 6400 25372 6409
rect 25412 6400 25464 6452
rect 12348 6332 12400 6384
rect 9404 6128 9456 6180
rect 7748 6103 7800 6112
rect 7748 6069 7773 6103
rect 7773 6069 7800 6103
rect 7748 6060 7800 6069
rect 7932 6103 7984 6112
rect 7932 6069 7941 6103
rect 7941 6069 7975 6103
rect 7975 6069 7984 6103
rect 7932 6060 7984 6069
rect 9864 6060 9916 6112
rect 11520 6196 11572 6248
rect 11796 6239 11848 6248
rect 11796 6205 11805 6239
rect 11805 6205 11839 6239
rect 11839 6205 11848 6239
rect 11796 6196 11848 6205
rect 12256 6239 12308 6248
rect 12256 6205 12265 6239
rect 12265 6205 12299 6239
rect 12299 6205 12308 6239
rect 12256 6196 12308 6205
rect 12348 6239 12400 6248
rect 12348 6205 12357 6239
rect 12357 6205 12391 6239
rect 12391 6205 12400 6239
rect 12348 6196 12400 6205
rect 15752 6332 15804 6384
rect 13268 6264 13320 6316
rect 13176 6239 13228 6248
rect 13176 6205 13185 6239
rect 13185 6205 13219 6239
rect 13219 6205 13228 6239
rect 13176 6196 13228 6205
rect 21272 6264 21324 6316
rect 23572 6264 23624 6316
rect 15292 6171 15344 6180
rect 15292 6137 15301 6171
rect 15301 6137 15335 6171
rect 15335 6137 15344 6171
rect 15292 6128 15344 6137
rect 15476 6171 15528 6180
rect 15476 6137 15485 6171
rect 15485 6137 15519 6171
rect 15519 6137 15528 6171
rect 16580 6239 16632 6248
rect 16580 6205 16589 6239
rect 16589 6205 16623 6239
rect 16623 6205 16632 6239
rect 16580 6196 16632 6205
rect 17040 6196 17092 6248
rect 17132 6196 17184 6248
rect 17868 6196 17920 6248
rect 21640 6196 21692 6248
rect 22928 6196 22980 6248
rect 25136 6196 25188 6248
rect 25964 6264 26016 6316
rect 26056 6196 26108 6248
rect 15476 6128 15528 6137
rect 17776 6128 17828 6180
rect 12164 6103 12216 6112
rect 12164 6069 12173 6103
rect 12173 6069 12207 6103
rect 12207 6069 12216 6103
rect 12164 6060 12216 6069
rect 13544 6103 13596 6112
rect 13544 6069 13553 6103
rect 13553 6069 13587 6103
rect 13587 6069 13596 6103
rect 13544 6060 13596 6069
rect 15200 6060 15252 6112
rect 15568 6103 15620 6112
rect 15568 6069 15577 6103
rect 15577 6069 15611 6103
rect 15611 6069 15620 6103
rect 15568 6060 15620 6069
rect 16028 6103 16080 6112
rect 16028 6069 16037 6103
rect 16037 6069 16071 6103
rect 16071 6069 16080 6103
rect 16028 6060 16080 6069
rect 16488 6060 16540 6112
rect 17224 6103 17276 6112
rect 17224 6069 17233 6103
rect 17233 6069 17267 6103
rect 17267 6069 17276 6103
rect 17224 6060 17276 6069
rect 17592 6060 17644 6112
rect 23112 6103 23164 6112
rect 23112 6069 23121 6103
rect 23121 6069 23155 6103
rect 23155 6069 23164 6103
rect 25688 6128 25740 6180
rect 25964 6171 26016 6180
rect 25964 6137 25973 6171
rect 25973 6137 26007 6171
rect 26007 6137 26016 6171
rect 25964 6128 26016 6137
rect 23112 6060 23164 6069
rect 7114 5958 7166 6010
rect 7178 5958 7230 6010
rect 7242 5958 7294 6010
rect 7306 5958 7358 6010
rect 7370 5958 7422 6010
rect 13830 5958 13882 6010
rect 13894 5958 13946 6010
rect 13958 5958 14010 6010
rect 14022 5958 14074 6010
rect 14086 5958 14138 6010
rect 20546 5958 20598 6010
rect 20610 5958 20662 6010
rect 20674 5958 20726 6010
rect 20738 5958 20790 6010
rect 20802 5958 20854 6010
rect 27262 5958 27314 6010
rect 27326 5958 27378 6010
rect 27390 5958 27442 6010
rect 27454 5958 27506 6010
rect 27518 5958 27570 6010
rect 3424 5856 3476 5908
rect 4896 5856 4948 5908
rect 5632 5899 5684 5908
rect 5632 5865 5641 5899
rect 5641 5865 5675 5899
rect 5675 5865 5684 5899
rect 5632 5856 5684 5865
rect 3700 5788 3752 5840
rect 3056 5763 3108 5772
rect 3056 5729 3065 5763
rect 3065 5729 3099 5763
rect 3099 5729 3108 5763
rect 3056 5720 3108 5729
rect 4160 5720 4212 5772
rect 4252 5763 4304 5772
rect 4252 5729 4261 5763
rect 4261 5729 4295 5763
rect 4295 5729 4304 5763
rect 4252 5720 4304 5729
rect 4528 5763 4580 5772
rect 4528 5729 4537 5763
rect 4537 5729 4571 5763
rect 4571 5729 4580 5763
rect 4528 5720 4580 5729
rect 4896 5763 4948 5772
rect 4896 5729 4905 5763
rect 4905 5729 4939 5763
rect 4939 5729 4948 5763
rect 4896 5720 4948 5729
rect 6184 5720 6236 5772
rect 6276 5763 6328 5772
rect 6276 5729 6285 5763
rect 6285 5729 6319 5763
rect 6319 5729 6328 5763
rect 6276 5720 6328 5729
rect 8208 5763 8260 5772
rect 9312 5788 9364 5840
rect 10048 5899 10100 5908
rect 10048 5865 10057 5899
rect 10057 5865 10091 5899
rect 10091 5865 10100 5899
rect 10048 5856 10100 5865
rect 10508 5899 10560 5908
rect 10508 5865 10517 5899
rect 10517 5865 10551 5899
rect 10551 5865 10560 5899
rect 10508 5856 10560 5865
rect 11796 5856 11848 5908
rect 12348 5856 12400 5908
rect 13176 5856 13228 5908
rect 8208 5729 8226 5763
rect 8226 5729 8260 5763
rect 8208 5720 8260 5729
rect 8852 5763 8904 5772
rect 8852 5729 8886 5763
rect 8886 5729 8904 5763
rect 8852 5720 8904 5729
rect 10140 5720 10192 5772
rect 13544 5788 13596 5840
rect 14188 5899 14240 5908
rect 14188 5865 14197 5899
rect 14197 5865 14231 5899
rect 14231 5865 14240 5899
rect 14188 5856 14240 5865
rect 15476 5856 15528 5908
rect 16488 5899 16540 5908
rect 16488 5865 16497 5899
rect 16497 5865 16531 5899
rect 16531 5865 16540 5899
rect 16488 5856 16540 5865
rect 14556 5788 14608 5840
rect 15568 5788 15620 5840
rect 15476 5763 15528 5772
rect 15476 5729 15494 5763
rect 15494 5729 15528 5763
rect 15476 5720 15528 5729
rect 16028 5720 16080 5772
rect 17224 5788 17276 5840
rect 15752 5695 15804 5704
rect 15752 5661 15761 5695
rect 15761 5661 15795 5695
rect 15795 5661 15804 5695
rect 15752 5652 15804 5661
rect 17776 5788 17828 5840
rect 17868 5831 17920 5840
rect 17868 5797 17877 5831
rect 17877 5797 17911 5831
rect 17911 5797 17920 5831
rect 17868 5788 17920 5797
rect 19984 5763 20036 5772
rect 19984 5729 19993 5763
rect 19993 5729 20027 5763
rect 20027 5729 20036 5763
rect 19984 5720 20036 5729
rect 21824 5856 21876 5908
rect 23020 5899 23072 5908
rect 23020 5865 23029 5899
rect 23029 5865 23063 5899
rect 23063 5865 23072 5899
rect 23020 5856 23072 5865
rect 25228 5856 25280 5908
rect 21548 5788 21600 5840
rect 21916 5831 21968 5840
rect 21732 5763 21784 5772
rect 21732 5729 21741 5763
rect 21741 5729 21775 5763
rect 21775 5729 21784 5763
rect 21732 5720 21784 5729
rect 7012 5627 7064 5636
rect 7012 5593 7021 5627
rect 7021 5593 7055 5627
rect 7055 5593 7064 5627
rect 7012 5584 7064 5593
rect 7196 5584 7248 5636
rect 19708 5695 19760 5704
rect 19708 5661 19717 5695
rect 19717 5661 19751 5695
rect 19751 5661 19760 5695
rect 19708 5652 19760 5661
rect 21916 5797 21925 5831
rect 21925 5797 21959 5831
rect 21959 5797 21968 5831
rect 21916 5788 21968 5797
rect 24676 5831 24728 5840
rect 24676 5797 24685 5831
rect 24685 5797 24719 5831
rect 24719 5797 24728 5831
rect 24676 5788 24728 5797
rect 22928 5763 22980 5772
rect 22928 5729 22937 5763
rect 22937 5729 22971 5763
rect 22971 5729 22980 5763
rect 22928 5720 22980 5729
rect 23112 5763 23164 5772
rect 23112 5729 23121 5763
rect 23121 5729 23155 5763
rect 23155 5729 23164 5763
rect 23112 5720 23164 5729
rect 25228 5763 25280 5772
rect 25228 5729 25237 5763
rect 25237 5729 25271 5763
rect 25271 5729 25280 5763
rect 25228 5720 25280 5729
rect 25412 5720 25464 5772
rect 25688 5763 25740 5772
rect 25688 5729 25697 5763
rect 25697 5729 25731 5763
rect 25731 5729 25740 5763
rect 25688 5720 25740 5729
rect 1124 5516 1176 5568
rect 2412 5559 2464 5568
rect 2412 5525 2421 5559
rect 2421 5525 2455 5559
rect 2455 5525 2464 5559
rect 2412 5516 2464 5525
rect 3148 5559 3200 5568
rect 3148 5525 3157 5559
rect 3157 5525 3191 5559
rect 3191 5525 3200 5559
rect 3148 5516 3200 5525
rect 7472 5516 7524 5568
rect 12532 5516 12584 5568
rect 16304 5516 16356 5568
rect 16580 5516 16632 5568
rect 17960 5584 18012 5636
rect 24308 5627 24360 5636
rect 24308 5593 24317 5627
rect 24317 5593 24351 5627
rect 24351 5593 24360 5627
rect 24308 5584 24360 5593
rect 18880 5516 18932 5568
rect 19340 5559 19392 5568
rect 19340 5525 19349 5559
rect 19349 5525 19383 5559
rect 19383 5525 19392 5559
rect 19340 5516 19392 5525
rect 20904 5559 20956 5568
rect 20904 5525 20913 5559
rect 20913 5525 20947 5559
rect 20947 5525 20956 5559
rect 20904 5516 20956 5525
rect 22560 5559 22612 5568
rect 22560 5525 22569 5559
rect 22569 5525 22603 5559
rect 22603 5525 22612 5559
rect 22560 5516 22612 5525
rect 24584 5516 24636 5568
rect 24768 5516 24820 5568
rect 25320 5516 25372 5568
rect 3756 5414 3808 5466
rect 3820 5414 3872 5466
rect 3884 5414 3936 5466
rect 3948 5414 4000 5466
rect 4012 5414 4064 5466
rect 10472 5414 10524 5466
rect 10536 5414 10588 5466
rect 10600 5414 10652 5466
rect 10664 5414 10716 5466
rect 10728 5414 10780 5466
rect 17188 5414 17240 5466
rect 17252 5414 17304 5466
rect 17316 5414 17368 5466
rect 17380 5414 17432 5466
rect 17444 5414 17496 5466
rect 23904 5414 23956 5466
rect 23968 5414 24020 5466
rect 24032 5414 24084 5466
rect 24096 5414 24148 5466
rect 24160 5414 24212 5466
rect 3056 5355 3108 5364
rect 3056 5321 3065 5355
rect 3065 5321 3099 5355
rect 3099 5321 3108 5355
rect 3056 5312 3108 5321
rect 4252 5312 4304 5364
rect 6276 5355 6328 5364
rect 6276 5321 6285 5355
rect 6285 5321 6319 5355
rect 6319 5321 6328 5355
rect 6276 5312 6328 5321
rect 6460 5312 6512 5364
rect 4804 5244 4856 5296
rect 1676 5219 1728 5228
rect 1676 5185 1685 5219
rect 1685 5185 1719 5219
rect 1719 5185 1728 5219
rect 1676 5176 1728 5185
rect 6092 5219 6144 5228
rect 6092 5185 6101 5219
rect 6101 5185 6135 5219
rect 6135 5185 6144 5219
rect 6920 5244 6972 5296
rect 7748 5312 7800 5364
rect 8208 5312 8260 5364
rect 8852 5312 8904 5364
rect 11796 5312 11848 5364
rect 14556 5355 14608 5364
rect 14556 5321 14565 5355
rect 14565 5321 14599 5355
rect 14599 5321 14608 5355
rect 14556 5312 14608 5321
rect 15200 5312 15252 5364
rect 15476 5312 15528 5364
rect 15752 5312 15804 5364
rect 6092 5176 6144 5185
rect 2412 5108 2464 5160
rect 3056 5108 3108 5160
rect 4988 5108 5040 5160
rect 5264 5151 5316 5160
rect 5264 5117 5273 5151
rect 5273 5117 5307 5151
rect 5307 5117 5316 5151
rect 5264 5108 5316 5117
rect 3332 5040 3384 5092
rect 4252 5040 4304 5092
rect 1400 5015 1452 5024
rect 1400 4981 1409 5015
rect 1409 4981 1443 5015
rect 1443 4981 1452 5015
rect 1400 4972 1452 4981
rect 3608 5015 3660 5024
rect 3608 4981 3617 5015
rect 3617 4981 3651 5015
rect 3651 4981 3660 5015
rect 3608 4972 3660 4981
rect 5908 5108 5960 5160
rect 6184 5151 6236 5160
rect 6184 5117 6193 5151
rect 6193 5117 6227 5151
rect 6227 5117 6236 5151
rect 6184 5108 6236 5117
rect 7840 5244 7892 5296
rect 8300 5244 8352 5296
rect 11888 5244 11940 5296
rect 12348 5244 12400 5296
rect 7196 5176 7248 5228
rect 7472 5151 7524 5160
rect 7472 5117 7481 5151
rect 7481 5117 7515 5151
rect 7515 5117 7524 5151
rect 7472 5108 7524 5117
rect 7932 5108 7984 5160
rect 9220 5151 9272 5160
rect 9220 5117 9229 5151
rect 9229 5117 9263 5151
rect 9263 5117 9272 5151
rect 9220 5108 9272 5117
rect 10784 5108 10836 5160
rect 11980 5108 12032 5160
rect 12532 5108 12584 5160
rect 12624 5151 12676 5160
rect 12624 5117 12633 5151
rect 12633 5117 12667 5151
rect 12667 5117 12676 5151
rect 12624 5108 12676 5117
rect 12716 5108 12768 5160
rect 13452 5108 13504 5160
rect 13728 5108 13780 5160
rect 7012 5040 7064 5092
rect 7564 5040 7616 5092
rect 11336 5040 11388 5092
rect 14648 5040 14700 5092
rect 15568 5176 15620 5228
rect 18144 5312 18196 5364
rect 17868 5244 17920 5296
rect 19708 5244 19760 5296
rect 6184 4972 6236 5024
rect 12716 4972 12768 5024
rect 15200 4972 15252 5024
rect 16304 5108 16356 5160
rect 18328 5176 18380 5228
rect 18880 5219 18932 5228
rect 18880 5185 18889 5219
rect 18889 5185 18923 5219
rect 18923 5185 18932 5219
rect 18880 5176 18932 5185
rect 21732 5312 21784 5364
rect 21824 5355 21876 5364
rect 21824 5321 21833 5355
rect 21833 5321 21867 5355
rect 21867 5321 21876 5355
rect 21824 5312 21876 5321
rect 23664 5244 23716 5296
rect 22560 5219 22612 5228
rect 22560 5185 22569 5219
rect 22569 5185 22603 5219
rect 22603 5185 22612 5219
rect 22560 5176 22612 5185
rect 24308 5312 24360 5364
rect 24676 5219 24728 5228
rect 24676 5185 24685 5219
rect 24685 5185 24719 5219
rect 24719 5185 24728 5219
rect 24676 5176 24728 5185
rect 25044 5219 25096 5228
rect 25044 5185 25053 5219
rect 25053 5185 25087 5219
rect 25087 5185 25096 5219
rect 25044 5176 25096 5185
rect 18144 5151 18196 5160
rect 18144 5117 18153 5151
rect 18153 5117 18187 5151
rect 18187 5117 18196 5151
rect 18144 5108 18196 5117
rect 19156 5151 19208 5160
rect 19156 5117 19165 5151
rect 19165 5117 19199 5151
rect 19199 5117 19208 5151
rect 19156 5108 19208 5117
rect 20904 5108 20956 5160
rect 21732 5151 21784 5160
rect 21732 5117 21741 5151
rect 21741 5117 21775 5151
rect 21775 5117 21784 5151
rect 21732 5108 21784 5117
rect 21916 5151 21968 5160
rect 21916 5117 21925 5151
rect 21925 5117 21959 5151
rect 21959 5117 21968 5151
rect 21916 5108 21968 5117
rect 22100 5108 22152 5160
rect 23204 5108 23256 5160
rect 24584 5151 24636 5160
rect 24584 5117 24593 5151
rect 24593 5117 24627 5151
rect 24627 5117 24636 5151
rect 24584 5108 24636 5117
rect 25320 5151 25372 5160
rect 25320 5117 25354 5151
rect 25354 5117 25372 5151
rect 25320 5108 25372 5117
rect 18052 5015 18104 5024
rect 18052 4981 18061 5015
rect 18061 4981 18095 5015
rect 18095 4981 18104 5015
rect 18052 4972 18104 4981
rect 19892 5015 19944 5024
rect 19892 4981 19901 5015
rect 19901 4981 19935 5015
rect 19935 4981 19944 5015
rect 19892 4972 19944 4981
rect 24400 4972 24452 5024
rect 25688 4972 25740 5024
rect 7114 4870 7166 4922
rect 7178 4870 7230 4922
rect 7242 4870 7294 4922
rect 7306 4870 7358 4922
rect 7370 4870 7422 4922
rect 13830 4870 13882 4922
rect 13894 4870 13946 4922
rect 13958 4870 14010 4922
rect 14022 4870 14074 4922
rect 14086 4870 14138 4922
rect 20546 4870 20598 4922
rect 20610 4870 20662 4922
rect 20674 4870 20726 4922
rect 20738 4870 20790 4922
rect 20802 4870 20854 4922
rect 27262 4870 27314 4922
rect 27326 4870 27378 4922
rect 27390 4870 27442 4922
rect 27454 4870 27506 4922
rect 27518 4870 27570 4922
rect 2136 4811 2188 4820
rect 2136 4777 2145 4811
rect 2145 4777 2179 4811
rect 2179 4777 2188 4811
rect 2136 4768 2188 4777
rect 2964 4811 3016 4820
rect 2964 4777 2973 4811
rect 2973 4777 3007 4811
rect 3007 4777 3016 4811
rect 2964 4768 3016 4777
rect 3332 4768 3384 4820
rect 1124 4675 1176 4684
rect 1124 4641 1133 4675
rect 1133 4641 1167 4675
rect 1167 4641 1176 4675
rect 1124 4632 1176 4641
rect 1400 4675 1452 4684
rect 1400 4641 1409 4675
rect 1409 4641 1443 4675
rect 1443 4641 1452 4675
rect 1400 4632 1452 4641
rect 3608 4700 3660 4752
rect 4896 4811 4948 4820
rect 4896 4777 4905 4811
rect 4905 4777 4939 4811
rect 4939 4777 4948 4811
rect 4896 4768 4948 4777
rect 4988 4811 5040 4820
rect 4988 4777 4997 4811
rect 4997 4777 5031 4811
rect 5031 4777 5040 4811
rect 4988 4768 5040 4777
rect 5908 4768 5960 4820
rect 6000 4743 6052 4752
rect 6000 4709 6009 4743
rect 6009 4709 6043 4743
rect 6043 4709 6052 4743
rect 6000 4700 6052 4709
rect 6460 4743 6512 4752
rect 3148 4675 3200 4684
rect 3148 4641 3157 4675
rect 3157 4641 3191 4675
rect 3191 4641 3200 4675
rect 3148 4632 3200 4641
rect 4712 4675 4764 4684
rect 4712 4641 4721 4675
rect 4721 4641 4755 4675
rect 4755 4641 4764 4675
rect 4712 4632 4764 4641
rect 5172 4675 5224 4684
rect 5172 4641 5181 4675
rect 5181 4641 5215 4675
rect 5215 4641 5224 4675
rect 5172 4632 5224 4641
rect 6460 4709 6469 4743
rect 6469 4709 6503 4743
rect 6503 4709 6512 4743
rect 6460 4700 6512 4709
rect 7748 4768 7800 4820
rect 8300 4768 8352 4820
rect 8576 4768 8628 4820
rect 10784 4811 10836 4820
rect 10784 4777 10793 4811
rect 10793 4777 10827 4811
rect 10827 4777 10836 4811
rect 10784 4768 10836 4777
rect 12624 4768 12676 4820
rect 13728 4768 13780 4820
rect 14832 4768 14884 4820
rect 18696 4768 18748 4820
rect 19156 4811 19208 4820
rect 19156 4777 19165 4811
rect 19165 4777 19199 4811
rect 19199 4777 19208 4811
rect 19156 4768 19208 4777
rect 20260 4811 20312 4820
rect 20260 4777 20269 4811
rect 20269 4777 20303 4811
rect 20303 4777 20312 4811
rect 20260 4768 20312 4777
rect 7564 4632 7616 4684
rect 6920 4539 6972 4548
rect 6920 4505 6929 4539
rect 6929 4505 6963 4539
rect 6963 4505 6972 4539
rect 6920 4496 6972 4505
rect 7104 4496 7156 4548
rect 11152 4632 11204 4684
rect 11244 4675 11296 4684
rect 11244 4641 11253 4675
rect 11253 4641 11287 4675
rect 11287 4641 11296 4675
rect 11244 4632 11296 4641
rect 11888 4700 11940 4752
rect 11980 4700 12032 4752
rect 12716 4743 12768 4752
rect 12716 4709 12725 4743
rect 12725 4709 12759 4743
rect 12759 4709 12768 4743
rect 12716 4700 12768 4709
rect 19340 4700 19392 4752
rect 22928 4768 22980 4820
rect 23204 4811 23256 4820
rect 23204 4777 23213 4811
rect 23213 4777 23247 4811
rect 23247 4777 23256 4811
rect 23204 4768 23256 4777
rect 24400 4811 24452 4820
rect 24400 4777 24409 4811
rect 24409 4777 24443 4811
rect 24443 4777 24452 4811
rect 24400 4768 24452 4777
rect 24584 4768 24636 4820
rect 11520 4675 11572 4684
rect 11520 4641 11529 4675
rect 11529 4641 11563 4675
rect 11563 4641 11572 4675
rect 11520 4632 11572 4641
rect 13176 4675 13228 4684
rect 13176 4641 13185 4675
rect 13185 4641 13219 4675
rect 13219 4641 13228 4675
rect 13176 4632 13228 4641
rect 13452 4675 13504 4684
rect 13452 4641 13461 4675
rect 13461 4641 13495 4675
rect 13495 4641 13504 4675
rect 13452 4632 13504 4641
rect 14464 4675 14516 4684
rect 14464 4641 14473 4675
rect 14473 4641 14507 4675
rect 14507 4641 14516 4675
rect 14464 4632 14516 4641
rect 17960 4632 18012 4684
rect 18052 4675 18104 4684
rect 18052 4641 18061 4675
rect 18061 4641 18095 4675
rect 18095 4641 18104 4675
rect 18052 4632 18104 4641
rect 18972 4675 19024 4684
rect 18972 4641 18981 4675
rect 18981 4641 19015 4675
rect 19015 4641 19024 4675
rect 18972 4632 19024 4641
rect 20720 4632 20772 4684
rect 21824 4675 21876 4684
rect 21824 4641 21833 4675
rect 21833 4641 21867 4675
rect 21867 4641 21876 4675
rect 21824 4632 21876 4641
rect 25412 4700 25464 4752
rect 25688 4700 25740 4752
rect 23388 4675 23440 4684
rect 23388 4641 23397 4675
rect 23397 4641 23431 4675
rect 23431 4641 23440 4675
rect 23388 4632 23440 4641
rect 24768 4632 24820 4684
rect 11796 4607 11848 4616
rect 11796 4573 11805 4607
rect 11805 4573 11839 4607
rect 11839 4573 11848 4607
rect 11796 4564 11848 4573
rect 11888 4607 11940 4616
rect 11888 4573 11897 4607
rect 11897 4573 11931 4607
rect 11931 4573 11940 4607
rect 11888 4564 11940 4573
rect 11060 4496 11112 4548
rect 11244 4496 11296 4548
rect 22100 4607 22152 4616
rect 22100 4573 22109 4607
rect 22109 4573 22143 4607
rect 22143 4573 22152 4607
rect 22100 4564 22152 4573
rect 12348 4496 12400 4548
rect 25228 4496 25280 4548
rect 2964 4428 3016 4480
rect 6092 4428 6144 4480
rect 9404 4471 9456 4480
rect 9404 4437 9413 4471
rect 9413 4437 9447 4471
rect 9447 4437 9456 4471
rect 9404 4428 9456 4437
rect 9680 4471 9732 4480
rect 9680 4437 9689 4471
rect 9689 4437 9723 4471
rect 9723 4437 9732 4471
rect 9680 4428 9732 4437
rect 16304 4428 16356 4480
rect 24492 4428 24544 4480
rect 3756 4326 3808 4378
rect 3820 4326 3872 4378
rect 3884 4326 3936 4378
rect 3948 4326 4000 4378
rect 4012 4326 4064 4378
rect 10472 4326 10524 4378
rect 10536 4326 10588 4378
rect 10600 4326 10652 4378
rect 10664 4326 10716 4378
rect 10728 4326 10780 4378
rect 17188 4326 17240 4378
rect 17252 4326 17304 4378
rect 17316 4326 17368 4378
rect 17380 4326 17432 4378
rect 17444 4326 17496 4378
rect 23904 4326 23956 4378
rect 23968 4326 24020 4378
rect 24032 4326 24084 4378
rect 24096 4326 24148 4378
rect 24160 4326 24212 4378
rect 4252 4267 4304 4276
rect 4252 4233 4261 4267
rect 4261 4233 4295 4267
rect 4295 4233 4304 4267
rect 4252 4224 4304 4233
rect 7564 4267 7616 4276
rect 7564 4233 7573 4267
rect 7573 4233 7607 4267
rect 7607 4233 7616 4267
rect 7564 4224 7616 4233
rect 11060 4267 11112 4276
rect 11060 4233 11069 4267
rect 11069 4233 11103 4267
rect 11103 4233 11112 4267
rect 11060 4224 11112 4233
rect 11244 4267 11296 4276
rect 11244 4233 11253 4267
rect 11253 4233 11287 4267
rect 11287 4233 11296 4267
rect 11244 4224 11296 4233
rect 13176 4224 13228 4276
rect 2964 4088 3016 4140
rect 2872 4063 2924 4072
rect 2872 4029 2881 4063
rect 2881 4029 2915 4063
rect 2915 4029 2924 4063
rect 2872 4020 2924 4029
rect 3424 4020 3476 4072
rect 4896 4156 4948 4208
rect 5264 4156 5316 4208
rect 11520 4156 11572 4208
rect 12072 4156 12124 4208
rect 14464 4224 14516 4276
rect 18972 4224 19024 4276
rect 22376 4267 22428 4276
rect 22376 4233 22385 4267
rect 22385 4233 22419 4267
rect 22419 4233 22428 4267
rect 22376 4224 22428 4233
rect 23388 4224 23440 4276
rect 25412 4224 25464 4276
rect 4160 3952 4212 4004
rect 6184 4020 6236 4072
rect 7012 4020 7064 4072
rect 7656 4020 7708 4072
rect 9404 4131 9456 4140
rect 9404 4097 9413 4131
rect 9413 4097 9447 4131
rect 9447 4097 9456 4131
rect 9404 4088 9456 4097
rect 7840 4063 7892 4072
rect 7840 4029 7849 4063
rect 7849 4029 7883 4063
rect 7883 4029 7892 4063
rect 7840 4020 7892 4029
rect 8024 4063 8076 4072
rect 8024 4029 8033 4063
rect 8033 4029 8067 4063
rect 8067 4029 8076 4063
rect 8024 4020 8076 4029
rect 8116 4063 8168 4072
rect 8116 4029 8125 4063
rect 8125 4029 8159 4063
rect 8159 4029 8168 4063
rect 8116 4020 8168 4029
rect 8760 4063 8812 4072
rect 2320 3884 2372 3936
rect 3240 3884 3292 3936
rect 6000 3884 6052 3936
rect 6920 3952 6972 4004
rect 8760 4029 8769 4063
rect 8769 4029 8803 4063
rect 8803 4029 8812 4063
rect 8760 4020 8812 4029
rect 9036 4063 9088 4072
rect 9036 4029 9045 4063
rect 9045 4029 9079 4063
rect 9079 4029 9088 4063
rect 9036 4020 9088 4029
rect 11152 4088 11204 4140
rect 8576 3995 8628 4004
rect 8576 3961 8585 3995
rect 8585 3961 8619 3995
rect 8619 3961 8628 3995
rect 11244 4020 11296 4072
rect 11796 4020 11848 4072
rect 12348 4020 12400 4072
rect 12808 4063 12860 4072
rect 12808 4029 12817 4063
rect 12817 4029 12851 4063
rect 12851 4029 12860 4063
rect 12808 4020 12860 4029
rect 8576 3952 8628 3961
rect 13728 3952 13780 4004
rect 14188 4020 14240 4072
rect 14740 4020 14792 4072
rect 16304 4131 16356 4140
rect 16304 4097 16313 4131
rect 16313 4097 16347 4131
rect 16347 4097 16356 4131
rect 16304 4088 16356 4097
rect 18328 4088 18380 4140
rect 19248 4156 19300 4208
rect 7564 3884 7616 3936
rect 10876 3884 10928 3936
rect 11152 3884 11204 3936
rect 12716 3927 12768 3936
rect 12716 3893 12725 3927
rect 12725 3893 12759 3927
rect 12759 3893 12768 3927
rect 12716 3884 12768 3893
rect 12808 3884 12860 3936
rect 15476 4063 15528 4072
rect 15476 4029 15485 4063
rect 15485 4029 15519 4063
rect 15519 4029 15528 4063
rect 15476 4020 15528 4029
rect 15936 4063 15988 4072
rect 15936 4029 15945 4063
rect 15945 4029 15979 4063
rect 15979 4029 15988 4063
rect 15936 4020 15988 4029
rect 16488 4020 16540 4072
rect 16764 4020 16816 4072
rect 17408 3995 17460 4004
rect 15200 3884 15252 3936
rect 17408 3961 17417 3995
rect 17417 3961 17451 3995
rect 17451 3961 17460 3995
rect 17408 3952 17460 3961
rect 18236 4020 18288 4072
rect 18696 4063 18748 4072
rect 18696 4029 18705 4063
rect 18705 4029 18739 4063
rect 18739 4029 18748 4063
rect 18696 4020 18748 4029
rect 18788 4020 18840 4072
rect 18972 4020 19024 4072
rect 20720 4131 20772 4140
rect 20720 4097 20729 4131
rect 20729 4097 20763 4131
rect 20763 4097 20772 4131
rect 20720 4088 20772 4097
rect 21364 4088 21416 4140
rect 18512 3952 18564 4004
rect 20168 3952 20220 4004
rect 20444 3952 20496 4004
rect 22192 4063 22244 4072
rect 22192 4029 22201 4063
rect 22201 4029 22235 4063
rect 22235 4029 22244 4063
rect 22192 4020 22244 4029
rect 22928 4020 22980 4072
rect 23204 4063 23256 4072
rect 23204 4029 23213 4063
rect 23213 4029 23247 4063
rect 23247 4029 23256 4063
rect 23204 4020 23256 4029
rect 23756 4020 23808 4072
rect 16304 3884 16356 3936
rect 17040 3884 17092 3936
rect 17868 3884 17920 3936
rect 18328 3927 18380 3936
rect 18328 3893 18337 3927
rect 18337 3893 18371 3927
rect 18371 3893 18380 3927
rect 18328 3884 18380 3893
rect 19984 3884 20036 3936
rect 22376 3884 22428 3936
rect 23388 3884 23440 3936
rect 7114 3782 7166 3834
rect 7178 3782 7230 3834
rect 7242 3782 7294 3834
rect 7306 3782 7358 3834
rect 7370 3782 7422 3834
rect 13830 3782 13882 3834
rect 13894 3782 13946 3834
rect 13958 3782 14010 3834
rect 14022 3782 14074 3834
rect 14086 3782 14138 3834
rect 20546 3782 20598 3834
rect 20610 3782 20662 3834
rect 20674 3782 20726 3834
rect 20738 3782 20790 3834
rect 20802 3782 20854 3834
rect 27262 3782 27314 3834
rect 27326 3782 27378 3834
rect 27390 3782 27442 3834
rect 27454 3782 27506 3834
rect 27518 3782 27570 3834
rect 2872 3680 2924 3732
rect 4252 3612 4304 3664
rect 5172 3680 5224 3732
rect 7012 3612 7064 3664
rect 3608 3587 3660 3596
rect 3608 3553 3617 3587
rect 3617 3553 3651 3587
rect 3651 3553 3660 3587
rect 3608 3544 3660 3553
rect 4068 3544 4120 3596
rect 4160 3587 4212 3596
rect 4160 3553 4169 3587
rect 4169 3553 4203 3587
rect 4203 3553 4212 3587
rect 4160 3544 4212 3553
rect 6092 3587 6144 3596
rect 6092 3553 6101 3587
rect 6101 3553 6135 3587
rect 6135 3553 6144 3587
rect 6092 3544 6144 3553
rect 6276 3587 6328 3596
rect 6276 3553 6285 3587
rect 6285 3553 6319 3587
rect 6319 3553 6328 3587
rect 6276 3544 6328 3553
rect 6828 3587 6880 3596
rect 6828 3553 6837 3587
rect 6837 3553 6871 3587
rect 6871 3553 6880 3587
rect 6828 3544 6880 3553
rect 6552 3476 6604 3528
rect 3516 3408 3568 3460
rect 5356 3408 5408 3460
rect 7288 3408 7340 3460
rect 4804 3383 4856 3392
rect 4804 3349 4813 3383
rect 4813 3349 4847 3383
rect 4847 3349 4856 3383
rect 4804 3340 4856 3349
rect 8024 3680 8076 3732
rect 7840 3612 7892 3664
rect 7656 3587 7708 3596
rect 7656 3553 7665 3587
rect 7665 3553 7699 3587
rect 7699 3553 7708 3587
rect 7656 3544 7708 3553
rect 8760 3612 8812 3664
rect 8576 3544 8628 3596
rect 9680 3680 9732 3732
rect 10140 3723 10192 3732
rect 10140 3689 10149 3723
rect 10149 3689 10183 3723
rect 10183 3689 10192 3723
rect 10140 3680 10192 3689
rect 12808 3680 12860 3732
rect 14188 3680 14240 3732
rect 15476 3723 15528 3732
rect 15476 3689 15501 3723
rect 15501 3689 15528 3723
rect 15476 3680 15528 3689
rect 15936 3723 15988 3732
rect 15936 3689 15945 3723
rect 15945 3689 15979 3723
rect 15979 3689 15988 3723
rect 15936 3680 15988 3689
rect 16488 3723 16540 3732
rect 16488 3689 16497 3723
rect 16497 3689 16531 3723
rect 16531 3689 16540 3723
rect 16488 3680 16540 3689
rect 17408 3680 17460 3732
rect 12716 3612 12768 3664
rect 10968 3587 11020 3596
rect 10968 3553 10977 3587
rect 10977 3553 11011 3587
rect 11011 3553 11020 3587
rect 10968 3544 11020 3553
rect 11152 3587 11204 3596
rect 11152 3553 11161 3587
rect 11161 3553 11195 3587
rect 11195 3553 11204 3587
rect 11152 3544 11204 3553
rect 11980 3544 12032 3596
rect 8024 3340 8076 3392
rect 11060 3383 11112 3392
rect 11060 3349 11069 3383
rect 11069 3349 11103 3383
rect 11103 3349 11112 3383
rect 11060 3340 11112 3349
rect 15108 3612 15160 3664
rect 17040 3612 17092 3664
rect 17868 3655 17920 3664
rect 17868 3621 17877 3655
rect 17877 3621 17911 3655
rect 17911 3621 17920 3655
rect 17868 3612 17920 3621
rect 18328 3680 18380 3732
rect 18880 3723 18932 3732
rect 18880 3689 18889 3723
rect 18889 3689 18923 3723
rect 18923 3689 18932 3723
rect 18880 3680 18932 3689
rect 20444 3680 20496 3732
rect 21824 3723 21876 3732
rect 21824 3689 21833 3723
rect 21833 3689 21867 3723
rect 21867 3689 21876 3723
rect 21824 3680 21876 3689
rect 25136 3680 25188 3732
rect 18696 3612 18748 3664
rect 13452 3587 13504 3596
rect 13452 3553 13461 3587
rect 13461 3553 13495 3587
rect 13495 3553 13504 3587
rect 13452 3544 13504 3553
rect 14188 3544 14240 3596
rect 15384 3544 15436 3596
rect 16304 3587 16356 3596
rect 16304 3553 16313 3587
rect 16313 3553 16347 3587
rect 16347 3553 16356 3587
rect 16304 3544 16356 3553
rect 18788 3587 18840 3596
rect 18788 3553 18797 3587
rect 18797 3553 18831 3587
rect 18831 3553 18840 3587
rect 18788 3544 18840 3553
rect 18972 3587 19024 3596
rect 18972 3553 18981 3587
rect 18981 3553 19015 3587
rect 19015 3553 19024 3587
rect 18972 3544 19024 3553
rect 19156 3544 19208 3596
rect 20168 3587 20220 3596
rect 20168 3553 20177 3587
rect 20177 3553 20211 3587
rect 20211 3553 20220 3587
rect 20168 3544 20220 3553
rect 23112 3612 23164 3664
rect 12808 3383 12860 3392
rect 12808 3349 12817 3383
rect 12817 3349 12851 3383
rect 12851 3349 12860 3383
rect 12808 3340 12860 3349
rect 14280 3476 14332 3528
rect 17960 3476 18012 3528
rect 18144 3476 18196 3528
rect 18604 3476 18656 3528
rect 19248 3476 19300 3528
rect 16304 3408 16356 3460
rect 18236 3408 18288 3460
rect 18972 3408 19024 3460
rect 20720 3587 20772 3596
rect 20720 3553 20729 3587
rect 20729 3553 20763 3587
rect 20763 3553 20772 3587
rect 20720 3544 20772 3553
rect 20628 3476 20680 3528
rect 22560 3544 22612 3596
rect 23204 3544 23256 3596
rect 24768 3587 24820 3596
rect 24768 3553 24777 3587
rect 24777 3553 24811 3587
rect 24811 3553 24820 3587
rect 24768 3544 24820 3553
rect 22836 3476 22888 3528
rect 21640 3408 21692 3460
rect 15476 3383 15528 3392
rect 15476 3349 15485 3383
rect 15485 3349 15519 3383
rect 15519 3349 15528 3383
rect 15476 3340 15528 3349
rect 16396 3340 16448 3392
rect 20444 3340 20496 3392
rect 20628 3340 20680 3392
rect 21364 3383 21416 3392
rect 21364 3349 21373 3383
rect 21373 3349 21407 3383
rect 21407 3349 21416 3383
rect 21364 3340 21416 3349
rect 22100 3340 22152 3392
rect 22928 3340 22980 3392
rect 23664 3383 23716 3392
rect 23664 3349 23673 3383
rect 23673 3349 23707 3383
rect 23707 3349 23716 3383
rect 23664 3340 23716 3349
rect 25044 3340 25096 3392
rect 3756 3238 3808 3290
rect 3820 3238 3872 3290
rect 3884 3238 3936 3290
rect 3948 3238 4000 3290
rect 4012 3238 4064 3290
rect 10472 3238 10524 3290
rect 10536 3238 10588 3290
rect 10600 3238 10652 3290
rect 10664 3238 10716 3290
rect 10728 3238 10780 3290
rect 17188 3238 17240 3290
rect 17252 3238 17304 3290
rect 17316 3238 17368 3290
rect 17380 3238 17432 3290
rect 17444 3238 17496 3290
rect 23904 3238 23956 3290
rect 23968 3238 24020 3290
rect 24032 3238 24084 3290
rect 24096 3238 24148 3290
rect 24160 3238 24212 3290
rect 4252 3179 4304 3188
rect 4252 3145 4261 3179
rect 4261 3145 4295 3179
rect 4295 3145 4304 3179
rect 4252 3136 4304 3145
rect 4712 3136 4764 3188
rect 4804 3136 4856 3188
rect 5172 3179 5224 3188
rect 5172 3145 5181 3179
rect 5181 3145 5215 3179
rect 5215 3145 5224 3179
rect 5172 3136 5224 3145
rect 6828 3136 6880 3188
rect 9956 3136 10008 3188
rect 10968 3136 11020 3188
rect 13452 3136 13504 3188
rect 13728 3179 13780 3188
rect 13728 3145 13737 3179
rect 13737 3145 13771 3179
rect 13771 3145 13780 3179
rect 13728 3136 13780 3145
rect 14280 3179 14332 3188
rect 14280 3145 14289 3179
rect 14289 3145 14323 3179
rect 14323 3145 14332 3179
rect 14280 3136 14332 3145
rect 14832 3136 14884 3188
rect 3608 3068 3660 3120
rect 4620 3068 4672 3120
rect 6092 3068 6144 3120
rect 8024 3068 8076 3120
rect 10232 3068 10284 3120
rect 12072 3068 12124 3120
rect 3148 2932 3200 2984
rect 3516 2975 3568 2984
rect 3516 2941 3525 2975
rect 3525 2941 3559 2975
rect 3559 2941 3568 2975
rect 3516 2932 3568 2941
rect 6276 3043 6328 3052
rect 1216 2796 1268 2848
rect 4804 2975 4856 2984
rect 4804 2941 4813 2975
rect 4813 2941 4847 2975
rect 4847 2941 4856 2975
rect 4804 2932 4856 2941
rect 4988 2975 5040 2984
rect 4988 2941 4997 2975
rect 4997 2941 5031 2975
rect 5031 2941 5040 2975
rect 4988 2932 5040 2941
rect 6276 3009 6285 3043
rect 6285 3009 6319 3043
rect 6319 3009 6328 3043
rect 6276 3000 6328 3009
rect 5264 2932 5316 2984
rect 5356 2975 5408 2984
rect 5356 2941 5365 2975
rect 5365 2941 5399 2975
rect 5399 2941 5408 2975
rect 5356 2932 5408 2941
rect 5540 2864 5592 2916
rect 6460 2975 6512 2984
rect 6460 2941 6499 2975
rect 6499 2941 6512 2975
rect 6460 2932 6512 2941
rect 6920 2975 6972 2984
rect 6920 2941 6929 2975
rect 6929 2941 6963 2975
rect 6963 2941 6972 2975
rect 6920 2932 6972 2941
rect 7748 2932 7800 2984
rect 7932 2932 7984 2984
rect 8300 2932 8352 2984
rect 11152 3000 11204 3052
rect 10968 2932 11020 2984
rect 11336 2932 11388 2984
rect 12072 2932 12124 2984
rect 12808 2975 12860 2984
rect 12808 2941 12817 2975
rect 12817 2941 12851 2975
rect 12851 2941 12860 2975
rect 12808 2932 12860 2941
rect 9956 2907 10008 2916
rect 9956 2873 9965 2907
rect 9965 2873 9999 2907
rect 9999 2873 10008 2907
rect 9956 2864 10008 2873
rect 7932 2839 7984 2848
rect 7932 2805 7941 2839
rect 7941 2805 7975 2839
rect 7975 2805 7984 2839
rect 7932 2796 7984 2805
rect 9680 2796 9732 2848
rect 11796 2907 11848 2916
rect 11796 2873 11805 2907
rect 11805 2873 11839 2907
rect 11839 2873 11848 2907
rect 11796 2864 11848 2873
rect 13544 2975 13596 2984
rect 13544 2941 13553 2975
rect 13553 2941 13587 2975
rect 13587 2941 13596 2975
rect 13544 2932 13596 2941
rect 14740 3068 14792 3120
rect 15384 3136 15436 3188
rect 15476 3068 15528 3120
rect 18420 3136 18472 3188
rect 18788 3136 18840 3188
rect 20076 3136 20128 3188
rect 21824 3136 21876 3188
rect 21916 3136 21968 3188
rect 22100 3136 22152 3188
rect 22560 3136 22612 3188
rect 22928 3136 22980 3188
rect 17684 3068 17736 3120
rect 20628 3111 20680 3120
rect 20628 3077 20637 3111
rect 20637 3077 20671 3111
rect 20671 3077 20680 3111
rect 20628 3068 20680 3077
rect 23388 3136 23440 3188
rect 23940 3136 23992 3188
rect 24308 3179 24360 3188
rect 24308 3145 24317 3179
rect 24317 3145 24351 3179
rect 24351 3145 24360 3179
rect 24308 3136 24360 3145
rect 24768 3179 24820 3188
rect 24768 3145 24777 3179
rect 24777 3145 24811 3179
rect 24811 3145 24820 3179
rect 24768 3136 24820 3145
rect 15384 3043 15436 3052
rect 15384 3009 15393 3043
rect 15393 3009 15427 3043
rect 15427 3009 15436 3043
rect 15384 3000 15436 3009
rect 16396 3043 16448 3052
rect 16396 3009 16405 3043
rect 16405 3009 16439 3043
rect 16439 3009 16448 3043
rect 16396 3000 16448 3009
rect 18144 3000 18196 3052
rect 10140 2796 10192 2848
rect 10968 2839 11020 2848
rect 10968 2805 10977 2839
rect 10977 2805 11011 2839
rect 11011 2805 11020 2839
rect 10968 2796 11020 2805
rect 11612 2796 11664 2848
rect 13636 2864 13688 2916
rect 13912 2864 13964 2916
rect 14280 2975 14332 2984
rect 14280 2941 14289 2975
rect 14289 2941 14323 2975
rect 14323 2941 14332 2975
rect 14280 2932 14332 2941
rect 14464 2975 14516 2984
rect 14464 2941 14473 2975
rect 14473 2941 14507 2975
rect 14507 2941 14516 2975
rect 14464 2932 14516 2941
rect 15936 2932 15988 2984
rect 15108 2907 15160 2916
rect 15108 2873 15117 2907
rect 15117 2873 15151 2907
rect 15151 2873 15160 2907
rect 15108 2864 15160 2873
rect 16856 2932 16908 2984
rect 18972 3000 19024 3052
rect 20444 3000 20496 3052
rect 18788 2975 18840 2984
rect 18788 2941 18798 2975
rect 18798 2941 18832 2975
rect 18832 2941 18840 2975
rect 18788 2932 18840 2941
rect 19156 2932 19208 2984
rect 20168 2932 20220 2984
rect 21640 2975 21692 2984
rect 21640 2941 21649 2975
rect 21649 2941 21683 2975
rect 21683 2941 21692 2975
rect 21640 2932 21692 2941
rect 22008 3043 22060 3052
rect 22008 3009 22017 3043
rect 22017 3009 22051 3043
rect 22051 3009 22060 3043
rect 22008 3000 22060 3009
rect 12716 2839 12768 2848
rect 12716 2805 12725 2839
rect 12725 2805 12759 2839
rect 12759 2805 12768 2839
rect 12716 2796 12768 2805
rect 14188 2796 14240 2848
rect 16120 2796 16172 2848
rect 18420 2907 18472 2916
rect 18420 2873 18429 2907
rect 18429 2873 18463 2907
rect 18463 2873 18472 2907
rect 18420 2864 18472 2873
rect 21824 2932 21876 2984
rect 22836 3000 22888 3052
rect 18052 2839 18104 2848
rect 18052 2805 18061 2839
rect 18061 2805 18095 2839
rect 18095 2805 18104 2839
rect 18052 2796 18104 2805
rect 18788 2796 18840 2848
rect 21916 2864 21968 2916
rect 20352 2796 20404 2848
rect 23664 2932 23716 2984
rect 23112 2864 23164 2916
rect 24216 2932 24268 2984
rect 25320 3000 25372 3052
rect 25044 2975 25096 2984
rect 25044 2941 25053 2975
rect 25053 2941 25087 2975
rect 25087 2941 25096 2975
rect 25044 2932 25096 2941
rect 25136 2796 25188 2848
rect 7114 2694 7166 2746
rect 7178 2694 7230 2746
rect 7242 2694 7294 2746
rect 7306 2694 7358 2746
rect 7370 2694 7422 2746
rect 13830 2694 13882 2746
rect 13894 2694 13946 2746
rect 13958 2694 14010 2746
rect 14022 2694 14074 2746
rect 14086 2694 14138 2746
rect 20546 2694 20598 2746
rect 20610 2694 20662 2746
rect 20674 2694 20726 2746
rect 20738 2694 20790 2746
rect 20802 2694 20854 2746
rect 27262 2694 27314 2746
rect 27326 2694 27378 2746
rect 27390 2694 27442 2746
rect 27454 2694 27506 2746
rect 27518 2694 27570 2746
rect 4804 2592 4856 2644
rect 3424 2499 3476 2508
rect 3424 2465 3433 2499
rect 3433 2465 3467 2499
rect 3467 2465 3476 2499
rect 3424 2456 3476 2465
rect 3148 2388 3200 2440
rect 4068 2456 4120 2508
rect 4528 2499 4580 2508
rect 4528 2465 4537 2499
rect 4537 2465 4571 2499
rect 4571 2465 4580 2499
rect 4528 2456 4580 2465
rect 4712 2499 4764 2508
rect 4712 2465 4721 2499
rect 4721 2465 4755 2499
rect 4755 2465 4764 2499
rect 4712 2456 4764 2465
rect 4896 2456 4948 2508
rect 8116 2592 8168 2644
rect 6092 2524 6144 2576
rect 6828 2524 6880 2576
rect 6920 2524 6972 2576
rect 5264 2456 5316 2508
rect 6184 2456 6236 2508
rect 7564 2499 7616 2508
rect 7564 2465 7573 2499
rect 7573 2465 7607 2499
rect 7607 2465 7616 2499
rect 7564 2456 7616 2465
rect 7932 2456 7984 2508
rect 8024 2499 8076 2508
rect 8024 2465 8033 2499
rect 8033 2465 8067 2499
rect 8067 2465 8076 2499
rect 8024 2456 8076 2465
rect 8300 2456 8352 2508
rect 9496 2456 9548 2508
rect 9680 2499 9732 2508
rect 9680 2465 9689 2499
rect 9689 2465 9723 2499
rect 9723 2465 9732 2499
rect 9680 2456 9732 2465
rect 10140 2499 10192 2508
rect 10140 2465 10149 2499
rect 10149 2465 10183 2499
rect 10183 2465 10192 2499
rect 10140 2456 10192 2465
rect 10232 2499 10284 2508
rect 10232 2465 10241 2499
rect 10241 2465 10275 2499
rect 10275 2465 10284 2499
rect 10232 2456 10284 2465
rect 4068 2320 4120 2372
rect 6000 2388 6052 2440
rect 6920 2431 6972 2440
rect 6920 2397 6929 2431
rect 6929 2397 6963 2431
rect 6963 2397 6972 2431
rect 6920 2388 6972 2397
rect 7012 2388 7064 2440
rect 11060 2456 11112 2508
rect 12900 2592 12952 2644
rect 11244 2388 11296 2440
rect 11612 2499 11664 2508
rect 11612 2465 11621 2499
rect 11621 2465 11655 2499
rect 11655 2465 11664 2499
rect 11612 2456 11664 2465
rect 11796 2499 11848 2508
rect 11796 2465 11805 2499
rect 11805 2465 11839 2499
rect 11839 2465 11848 2499
rect 11796 2456 11848 2465
rect 15936 2635 15988 2644
rect 15936 2601 15945 2635
rect 15945 2601 15979 2635
rect 15979 2601 15988 2635
rect 15936 2592 15988 2601
rect 18144 2592 18196 2644
rect 20076 2592 20128 2644
rect 23112 2592 23164 2644
rect 13544 2388 13596 2440
rect 13636 2388 13688 2440
rect 14280 2456 14332 2508
rect 15476 2456 15528 2508
rect 16120 2499 16172 2508
rect 16120 2465 16129 2499
rect 16129 2465 16163 2499
rect 16163 2465 16172 2499
rect 16120 2456 16172 2465
rect 16304 2456 16356 2508
rect 18052 2524 18104 2576
rect 17960 2499 18012 2508
rect 17960 2465 17969 2499
rect 17969 2465 18003 2499
rect 18003 2465 18012 2499
rect 17960 2456 18012 2465
rect 18144 2499 18196 2508
rect 18144 2465 18153 2499
rect 18153 2465 18187 2499
rect 18187 2465 18196 2499
rect 18144 2456 18196 2465
rect 18604 2499 18656 2508
rect 18604 2465 18613 2499
rect 18613 2465 18647 2499
rect 18647 2465 18656 2499
rect 18604 2456 18656 2465
rect 18788 2499 18840 2508
rect 18788 2465 18797 2499
rect 18797 2465 18831 2499
rect 18831 2465 18840 2499
rect 18788 2456 18840 2465
rect 18972 2456 19024 2508
rect 12716 2320 12768 2372
rect 18052 2320 18104 2372
rect 20076 2499 20128 2508
rect 20076 2465 20085 2499
rect 20085 2465 20119 2499
rect 20119 2465 20128 2499
rect 20076 2456 20128 2465
rect 20444 2524 20496 2576
rect 20352 2456 20404 2508
rect 20720 2456 20772 2508
rect 22008 2456 22060 2508
rect 22284 2456 22336 2508
rect 24308 2592 24360 2644
rect 22192 2320 22244 2372
rect 23664 2320 23716 2372
rect 24216 2320 24268 2372
rect 4160 2252 4212 2304
rect 4988 2252 5040 2304
rect 5540 2252 5592 2304
rect 5908 2252 5960 2304
rect 6276 2252 6328 2304
rect 8208 2252 8260 2304
rect 9680 2295 9732 2304
rect 9680 2261 9689 2295
rect 9689 2261 9723 2295
rect 9723 2261 9732 2295
rect 9680 2252 9732 2261
rect 9956 2252 10008 2304
rect 10232 2295 10284 2304
rect 10232 2261 10241 2295
rect 10241 2261 10275 2295
rect 10275 2261 10284 2295
rect 10232 2252 10284 2261
rect 11244 2252 11296 2304
rect 11336 2252 11388 2304
rect 11888 2252 11940 2304
rect 12256 2252 12308 2304
rect 15200 2252 15252 2304
rect 16304 2295 16356 2304
rect 16304 2261 16313 2295
rect 16313 2261 16347 2295
rect 16347 2261 16356 2295
rect 16304 2252 16356 2261
rect 16580 2295 16632 2304
rect 16580 2261 16589 2295
rect 16589 2261 16623 2295
rect 16623 2261 16632 2295
rect 16580 2252 16632 2261
rect 17684 2295 17736 2304
rect 17684 2261 17693 2295
rect 17693 2261 17727 2295
rect 17727 2261 17736 2295
rect 17684 2252 17736 2261
rect 18512 2252 18564 2304
rect 18972 2252 19024 2304
rect 19064 2295 19116 2304
rect 19064 2261 19073 2295
rect 19073 2261 19107 2295
rect 19107 2261 19116 2295
rect 19064 2252 19116 2261
rect 19800 2252 19852 2304
rect 20260 2295 20312 2304
rect 20260 2261 20269 2295
rect 20269 2261 20303 2295
rect 20303 2261 20312 2295
rect 20260 2252 20312 2261
rect 21548 2252 21600 2304
rect 23020 2295 23072 2304
rect 23020 2261 23029 2295
rect 23029 2261 23063 2295
rect 23063 2261 23072 2295
rect 23020 2252 23072 2261
rect 3756 2150 3808 2202
rect 3820 2150 3872 2202
rect 3884 2150 3936 2202
rect 3948 2150 4000 2202
rect 4012 2150 4064 2202
rect 10472 2150 10524 2202
rect 10536 2150 10588 2202
rect 10600 2150 10652 2202
rect 10664 2150 10716 2202
rect 10728 2150 10780 2202
rect 17188 2150 17240 2202
rect 17252 2150 17304 2202
rect 17316 2150 17368 2202
rect 17380 2150 17432 2202
rect 17444 2150 17496 2202
rect 23904 2150 23956 2202
rect 23968 2150 24020 2202
rect 24032 2150 24084 2202
rect 24096 2150 24148 2202
rect 24160 2150 24212 2202
rect 940 1887 992 1896
rect 940 1853 949 1887
rect 949 1853 983 1887
rect 983 1853 992 1887
rect 940 1844 992 1853
rect 1768 1844 1820 1896
rect 2136 1887 2188 1896
rect 2136 1853 2145 1887
rect 2145 1853 2179 1887
rect 2179 1853 2188 1887
rect 2136 1844 2188 1853
rect 3148 1844 3200 1896
rect 4712 1912 4764 1964
rect 3516 1887 3568 1896
rect 3516 1853 3525 1887
rect 3525 1853 3559 1887
rect 3559 1853 3568 1887
rect 3516 1844 3568 1853
rect 4252 1887 4304 1896
rect 4252 1853 4261 1887
rect 4261 1853 4295 1887
rect 4295 1853 4304 1887
rect 4252 1844 4304 1853
rect 4528 1887 4580 1896
rect 4528 1853 4537 1887
rect 4537 1853 4571 1887
rect 4571 1853 4580 1887
rect 4528 1844 4580 1853
rect 4620 1887 4672 1896
rect 4620 1853 4629 1887
rect 4629 1853 4663 1887
rect 4663 1853 4672 1887
rect 4620 1844 4672 1853
rect 6000 2048 6052 2100
rect 10968 2048 11020 2100
rect 6920 1980 6972 2032
rect 6276 1955 6328 1964
rect 6276 1921 6285 1955
rect 6285 1921 6319 1955
rect 6319 1921 6328 1955
rect 6276 1912 6328 1921
rect 5264 1844 5316 1896
rect 5448 1776 5500 1828
rect 6552 1887 6604 1896
rect 6552 1853 6561 1887
rect 6561 1853 6595 1887
rect 6595 1853 6604 1887
rect 6552 1844 6604 1853
rect 7472 1844 7524 1896
rect 9036 1887 9088 1896
rect 9036 1853 9045 1887
rect 9045 1853 9079 1887
rect 9079 1853 9088 1887
rect 9036 1844 9088 1853
rect 10232 1912 10284 1964
rect 18880 2048 18932 2100
rect 20628 1980 20680 2032
rect 10048 1844 10100 1896
rect 10876 1887 10928 1896
rect 10876 1853 10885 1887
rect 10885 1853 10919 1887
rect 10919 1853 10928 1887
rect 10876 1844 10928 1853
rect 11060 1887 11112 1896
rect 11060 1853 11069 1887
rect 11069 1853 11103 1887
rect 11103 1853 11112 1887
rect 11060 1844 11112 1853
rect 11888 1887 11940 1896
rect 11888 1853 11897 1887
rect 11897 1853 11931 1887
rect 11931 1853 11940 1887
rect 11888 1844 11940 1853
rect 12716 1887 12768 1896
rect 12716 1853 12725 1887
rect 12725 1853 12759 1887
rect 12759 1853 12768 1887
rect 12716 1844 12768 1853
rect 12900 1844 12952 1896
rect 14464 1912 14516 1964
rect 15200 1955 15252 1964
rect 15200 1921 15209 1955
rect 15209 1921 15243 1955
rect 15243 1921 15252 1955
rect 15200 1912 15252 1921
rect 6644 1776 6696 1828
rect 11796 1776 11848 1828
rect 13544 1887 13596 1896
rect 13544 1853 13553 1887
rect 13553 1853 13587 1887
rect 13587 1853 13596 1887
rect 13544 1844 13596 1853
rect 14188 1844 14240 1896
rect 14556 1887 14608 1896
rect 14556 1853 14565 1887
rect 14565 1853 14599 1887
rect 14599 1853 14608 1887
rect 14556 1844 14608 1853
rect 15476 1887 15528 1896
rect 15476 1853 15485 1887
rect 15485 1853 15519 1887
rect 15519 1853 15528 1887
rect 15476 1844 15528 1853
rect 16120 1844 16172 1896
rect 16396 1887 16448 1896
rect 16396 1853 16405 1887
rect 16405 1853 16439 1887
rect 16439 1853 16448 1887
rect 16396 1844 16448 1853
rect 17316 1844 17368 1896
rect 17592 1844 17644 1896
rect 17868 1887 17920 1896
rect 17868 1853 17877 1887
rect 17877 1853 17911 1887
rect 17911 1853 17920 1887
rect 17868 1844 17920 1853
rect 18696 1887 18748 1896
rect 18696 1853 18705 1887
rect 18705 1853 18739 1887
rect 18739 1853 18748 1887
rect 18696 1844 18748 1853
rect 19248 1844 19300 1896
rect 19800 1887 19852 1896
rect 19800 1853 19809 1887
rect 19809 1853 19843 1887
rect 19843 1853 19852 1887
rect 19800 1844 19852 1853
rect 20444 1844 20496 1896
rect 22284 2048 22336 2100
rect 22376 1980 22428 2032
rect 23572 1912 23624 1964
rect 24860 1912 24912 1964
rect 21364 1844 21416 1896
rect 22192 1844 22244 1896
rect 22468 1844 22520 1896
rect 23388 1844 23440 1896
rect 23756 1844 23808 1896
rect 24308 1844 24360 1896
rect 24952 1844 25004 1896
rect 25228 1844 25280 1896
rect 2964 1708 3016 1760
rect 3608 1751 3660 1760
rect 3608 1717 3617 1751
rect 3617 1717 3651 1751
rect 3651 1717 3660 1751
rect 3608 1708 3660 1717
rect 4528 1708 4580 1760
rect 4804 1708 4856 1760
rect 12992 1708 13044 1760
rect 13176 1751 13228 1760
rect 13176 1717 13185 1751
rect 13185 1717 13219 1751
rect 13219 1717 13228 1751
rect 13176 1708 13228 1717
rect 7114 1606 7166 1658
rect 7178 1606 7230 1658
rect 7242 1606 7294 1658
rect 7306 1606 7358 1658
rect 7370 1606 7422 1658
rect 13830 1606 13882 1658
rect 13894 1606 13946 1658
rect 13958 1606 14010 1658
rect 14022 1606 14074 1658
rect 14086 1606 14138 1658
rect 20546 1606 20598 1658
rect 20610 1606 20662 1658
rect 20674 1606 20726 1658
rect 20738 1606 20790 1658
rect 20802 1606 20854 1658
rect 27262 1606 27314 1658
rect 27326 1606 27378 1658
rect 27390 1606 27442 1658
rect 27454 1606 27506 1658
rect 27518 1606 27570 1658
rect 1216 1411 1268 1420
rect 1216 1377 1225 1411
rect 1225 1377 1259 1411
rect 1259 1377 1268 1411
rect 1216 1368 1268 1377
rect 2320 1436 2372 1488
rect 3516 1436 3568 1488
rect 2964 1411 3016 1420
rect 2964 1377 2973 1411
rect 2973 1377 3007 1411
rect 3007 1377 3016 1411
rect 2964 1368 3016 1377
rect 3608 1411 3660 1420
rect 3608 1377 3617 1411
rect 3617 1377 3651 1411
rect 3651 1377 3660 1411
rect 3608 1368 3660 1377
rect 4436 1411 4488 1420
rect 4436 1377 4445 1411
rect 4445 1377 4479 1411
rect 4479 1377 4488 1411
rect 4436 1368 4488 1377
rect 4804 1411 4856 1420
rect 4804 1377 4813 1411
rect 4813 1377 4847 1411
rect 4847 1377 4856 1411
rect 4804 1368 4856 1377
rect 5632 1411 5684 1420
rect 5632 1377 5641 1411
rect 5641 1377 5675 1411
rect 5675 1377 5684 1411
rect 5632 1368 5684 1377
rect 3240 1343 3292 1352
rect 3240 1309 3249 1343
rect 3249 1309 3283 1343
rect 3283 1309 3292 1343
rect 3240 1300 3292 1309
rect 3332 1343 3384 1352
rect 3332 1309 3341 1343
rect 3341 1309 3375 1343
rect 3375 1309 3384 1343
rect 3332 1300 3384 1309
rect 1308 1164 1360 1216
rect 5448 1300 5500 1352
rect 6920 1368 6972 1420
rect 7012 1411 7064 1420
rect 7012 1377 7021 1411
rect 7021 1377 7055 1411
rect 7055 1377 7064 1411
rect 7012 1368 7064 1377
rect 8392 1504 8444 1556
rect 8208 1411 8260 1420
rect 8208 1377 8217 1411
rect 8217 1377 8251 1411
rect 8251 1377 8260 1411
rect 8208 1368 8260 1377
rect 8944 1368 8996 1420
rect 9956 1411 10008 1420
rect 9956 1377 9965 1411
rect 9965 1377 9999 1411
rect 9999 1377 10008 1411
rect 9956 1368 10008 1377
rect 11152 1504 11204 1556
rect 17776 1504 17828 1556
rect 11060 1436 11112 1488
rect 17040 1436 17092 1488
rect 7932 1343 7984 1352
rect 7932 1309 7941 1343
rect 7941 1309 7975 1343
rect 7975 1309 7984 1343
rect 7932 1300 7984 1309
rect 11336 1368 11388 1420
rect 12072 1411 12124 1420
rect 12072 1377 12081 1411
rect 12081 1377 12115 1411
rect 12115 1377 12124 1411
rect 12072 1368 12124 1377
rect 12992 1411 13044 1420
rect 12992 1377 13001 1411
rect 13001 1377 13035 1411
rect 13035 1377 13044 1411
rect 12992 1368 13044 1377
rect 13544 1368 13596 1420
rect 13728 1368 13780 1420
rect 14464 1411 14516 1420
rect 14464 1377 14473 1411
rect 14473 1377 14507 1411
rect 14507 1377 14516 1411
rect 14464 1368 14516 1377
rect 14556 1411 14608 1420
rect 14556 1377 14565 1411
rect 14565 1377 14599 1411
rect 14599 1377 14608 1411
rect 14556 1368 14608 1377
rect 14832 1411 14884 1420
rect 14832 1377 14841 1411
rect 14841 1377 14875 1411
rect 14875 1377 14884 1411
rect 14832 1368 14884 1377
rect 15568 1368 15620 1420
rect 16304 1368 16356 1420
rect 16764 1368 16816 1420
rect 17316 1411 17368 1420
rect 17316 1377 17325 1411
rect 17325 1377 17359 1411
rect 17359 1377 17368 1411
rect 17316 1368 17368 1377
rect 17868 1436 17920 1488
rect 18512 1436 18564 1488
rect 19064 1436 19116 1488
rect 13360 1343 13412 1352
rect 13360 1309 13369 1343
rect 13369 1309 13403 1343
rect 13403 1309 13412 1343
rect 13360 1300 13412 1309
rect 18880 1368 18932 1420
rect 22284 1436 22336 1488
rect 20076 1368 20128 1420
rect 21548 1411 21600 1420
rect 21548 1377 21557 1411
rect 21557 1377 21591 1411
rect 21591 1377 21600 1411
rect 21548 1368 21600 1377
rect 21640 1368 21692 1420
rect 22468 1411 22520 1420
rect 22468 1377 22477 1411
rect 22477 1377 22511 1411
rect 22511 1377 22520 1411
rect 22468 1368 22520 1377
rect 22928 1436 22980 1488
rect 22836 1368 22888 1420
rect 24308 1368 24360 1420
rect 24860 1411 24912 1420
rect 24860 1377 24869 1411
rect 24869 1377 24903 1411
rect 24903 1377 24912 1411
rect 24860 1368 24912 1377
rect 25136 1411 25188 1420
rect 25136 1377 25145 1411
rect 25145 1377 25179 1411
rect 25179 1377 25188 1411
rect 25136 1368 25188 1377
rect 25504 1368 25556 1420
rect 19248 1300 19300 1352
rect 21272 1343 21324 1352
rect 21272 1309 21281 1343
rect 21281 1309 21315 1343
rect 21315 1309 21324 1343
rect 21272 1300 21324 1309
rect 23388 1300 23440 1352
rect 5448 1164 5500 1216
rect 6736 1164 6788 1216
rect 6828 1164 6880 1216
rect 9404 1164 9456 1216
rect 13728 1164 13780 1216
rect 19984 1164 20036 1216
rect 3756 1062 3808 1114
rect 3820 1062 3872 1114
rect 3884 1062 3936 1114
rect 3948 1062 4000 1114
rect 4012 1062 4064 1114
rect 10472 1062 10524 1114
rect 10536 1062 10588 1114
rect 10600 1062 10652 1114
rect 10664 1062 10716 1114
rect 10728 1062 10780 1114
rect 17188 1062 17240 1114
rect 17252 1062 17304 1114
rect 17316 1062 17368 1114
rect 17380 1062 17432 1114
rect 17444 1062 17496 1114
rect 23904 1062 23956 1114
rect 23968 1062 24020 1114
rect 24032 1062 24084 1114
rect 24096 1062 24148 1114
rect 24160 1062 24212 1114
rect 940 960 992 1012
rect 1308 960 1360 1012
rect 3332 960 3384 1012
rect 5448 1003 5500 1012
rect 5448 969 5457 1003
rect 5457 969 5491 1003
rect 5491 969 5500 1003
rect 5448 960 5500 969
rect 7932 1003 7984 1012
rect 7932 969 7941 1003
rect 7941 969 7975 1003
rect 7975 969 7984 1003
rect 7932 960 7984 969
rect 9036 1003 9088 1012
rect 9036 969 9045 1003
rect 9045 969 9079 1003
rect 9079 969 9088 1003
rect 9036 960 9088 969
rect 13360 960 13412 1012
rect 21272 1003 21324 1012
rect 21272 969 21281 1003
rect 21281 969 21315 1003
rect 21315 969 21324 1003
rect 21272 960 21324 969
rect 21364 960 21416 1012
rect 23572 960 23624 1012
rect 3240 892 3292 944
rect 2136 756 2188 808
rect 4160 824 4212 876
rect 4252 867 4304 876
rect 4252 833 4261 867
rect 4261 833 4295 867
rect 4295 833 4304 867
rect 4252 824 4304 833
rect 6736 867 6788 876
rect 6736 833 6745 867
rect 6745 833 6779 867
rect 6779 833 6788 867
rect 6736 824 6788 833
rect 9404 867 9456 876
rect 9404 833 9413 867
rect 9413 833 9447 867
rect 9447 833 9456 867
rect 9404 824 9456 833
rect 10876 824 10928 876
rect 12256 867 12308 876
rect 12256 833 12265 867
rect 12265 833 12299 867
rect 12299 833 12308 867
rect 12256 824 12308 833
rect 18696 867 18748 876
rect 18696 833 18705 867
rect 18705 833 18739 867
rect 18739 833 18748 867
rect 18696 824 18748 833
rect 19984 867 20036 876
rect 19984 833 19993 867
rect 19993 833 20027 867
rect 20027 833 20036 867
rect 19984 824 20036 833
rect 23756 824 23808 876
rect 2872 756 2924 808
rect 4528 799 4580 808
rect 4528 765 4537 799
rect 4537 765 4571 799
rect 4571 765 4580 799
rect 4528 756 4580 765
rect 5080 756 5132 808
rect 5908 756 5960 808
rect 7840 799 7892 808
rect 7840 765 7849 799
rect 7849 765 7883 799
rect 7883 765 7892 799
rect 7840 756 7892 765
rect 9680 799 9732 808
rect 9680 765 9689 799
rect 9689 765 9723 799
rect 9723 765 9732 799
rect 9680 756 9732 765
rect 10600 756 10652 808
rect 11244 799 11296 808
rect 11244 765 11253 799
rect 11253 765 11287 799
rect 11287 765 11296 799
rect 11244 756 11296 765
rect 11704 756 11756 808
rect 13176 756 13228 808
rect 13360 799 13412 808
rect 13360 765 13369 799
rect 13369 765 13403 799
rect 13403 765 13412 799
rect 13360 756 13412 765
rect 14188 756 14240 808
rect 14280 799 14332 808
rect 14280 765 14289 799
rect 14289 765 14323 799
rect 14323 765 14332 799
rect 14280 756 14332 765
rect 15016 756 15068 808
rect 16396 756 16448 808
rect 16580 756 16632 808
rect 17224 756 17276 808
rect 17592 756 17644 808
rect 17684 799 17736 808
rect 17684 765 17693 799
rect 17693 765 17727 799
rect 17727 765 17736 799
rect 17684 756 17736 765
rect 18328 756 18380 808
rect 18972 799 19024 808
rect 18972 765 18981 799
rect 18981 765 19015 799
rect 19015 765 19024 799
rect 18972 756 19024 765
rect 19432 756 19484 808
rect 20260 799 20312 808
rect 20260 765 20269 799
rect 20269 765 20303 799
rect 20303 765 20312 799
rect 20260 756 20312 765
rect 21088 799 21140 808
rect 21088 765 21097 799
rect 21097 765 21131 799
rect 21131 765 21140 799
rect 21088 756 21140 765
rect 22376 756 22428 808
rect 22560 756 22612 808
rect 23296 799 23348 808
rect 23296 765 23305 799
rect 23305 765 23339 799
rect 23339 765 23348 799
rect 23296 756 23348 765
rect 23664 756 23716 808
rect 24492 756 24544 808
rect 25228 756 25280 808
rect 25320 799 25372 808
rect 25320 765 25329 799
rect 25329 765 25363 799
rect 25363 765 25372 799
rect 25320 756 25372 765
rect 26056 756 26108 808
rect 7114 518 7166 570
rect 7178 518 7230 570
rect 7242 518 7294 570
rect 7306 518 7358 570
rect 7370 518 7422 570
rect 13830 518 13882 570
rect 13894 518 13946 570
rect 13958 518 14010 570
rect 14022 518 14074 570
rect 14086 518 14138 570
rect 20546 518 20598 570
rect 20610 518 20662 570
rect 20674 518 20726 570
rect 20738 518 20790 570
rect 20802 518 20854 570
rect 27262 518 27314 570
rect 27326 518 27378 570
rect 27390 518 27442 570
rect 27454 518 27506 570
rect 27518 518 27570 570
rect 20444 416 20496 468
rect 20628 416 20680 468
<< metal2 >>
rect 1398 31600 1454 32000
rect 2870 31600 2926 32000
rect 4342 31600 4398 32000
rect 5814 31600 5870 32000
rect 7286 31600 7342 32000
rect 7392 31606 7604 31634
rect 1412 29850 1440 31600
rect 2884 30138 2912 31600
rect 3756 30492 4064 30501
rect 3756 30490 3762 30492
rect 3818 30490 3842 30492
rect 3898 30490 3922 30492
rect 3978 30490 4002 30492
rect 4058 30490 4064 30492
rect 3818 30438 3820 30490
rect 4000 30438 4002 30490
rect 3756 30436 3762 30438
rect 3818 30436 3842 30438
rect 3898 30436 3922 30438
rect 3978 30436 4002 30438
rect 4058 30436 4064 30438
rect 3756 30427 4064 30436
rect 4356 30326 4384 31600
rect 5632 30796 5684 30802
rect 5632 30738 5684 30744
rect 4344 30320 4396 30326
rect 4344 30262 4396 30268
rect 3240 30184 3292 30190
rect 2780 30116 2832 30122
rect 2884 30110 3004 30138
rect 3240 30126 3292 30132
rect 5540 30184 5592 30190
rect 5540 30126 5592 30132
rect 2780 30058 2832 30064
rect 1400 29844 1452 29850
rect 1400 29786 1452 29792
rect 2504 29504 2556 29510
rect 2504 29446 2556 29452
rect 1860 27532 1912 27538
rect 1860 27474 1912 27480
rect 848 26920 900 26926
rect 848 26862 900 26868
rect 860 25362 888 26862
rect 1872 26858 1900 27474
rect 2044 27396 2096 27402
rect 2044 27338 2096 27344
rect 1124 26852 1176 26858
rect 1124 26794 1176 26800
rect 1492 26852 1544 26858
rect 1492 26794 1544 26800
rect 1860 26852 1912 26858
rect 1860 26794 1912 26800
rect 1136 26586 1164 26794
rect 1124 26580 1176 26586
rect 1124 26522 1176 26528
rect 848 25356 900 25362
rect 848 25298 900 25304
rect 1124 25356 1176 25362
rect 1124 25298 1176 25304
rect 1136 24954 1164 25298
rect 1124 24948 1176 24954
rect 1124 24890 1176 24896
rect 1504 23526 1532 26794
rect 1860 25696 1912 25702
rect 1860 25638 1912 25644
rect 1872 24682 1900 25638
rect 1952 24948 2004 24954
rect 1952 24890 2004 24896
rect 1860 24676 1912 24682
rect 1860 24618 1912 24624
rect 1860 24064 1912 24070
rect 1964 24052 1992 24890
rect 2056 24682 2084 27338
rect 2412 26920 2464 26926
rect 2412 26862 2464 26868
rect 2228 26784 2280 26790
rect 2228 26726 2280 26732
rect 2320 26784 2372 26790
rect 2320 26726 2372 26732
rect 2240 26586 2268 26726
rect 2228 26580 2280 26586
rect 2228 26522 2280 26528
rect 2332 26450 2360 26726
rect 2320 26444 2372 26450
rect 2320 26386 2372 26392
rect 2424 26314 2452 26862
rect 2412 26308 2464 26314
rect 2412 26250 2464 26256
rect 2424 25906 2452 26250
rect 2412 25900 2464 25906
rect 2412 25842 2464 25848
rect 2424 25362 2452 25842
rect 2412 25356 2464 25362
rect 2412 25298 2464 25304
rect 2136 25288 2188 25294
rect 2136 25230 2188 25236
rect 2044 24676 2096 24682
rect 2044 24618 2096 24624
rect 1912 24024 1992 24052
rect 1860 24006 1912 24012
rect 1872 23594 1900 24006
rect 2056 23882 2084 24618
rect 2148 24206 2176 25230
rect 2228 25152 2280 25158
rect 2228 25094 2280 25100
rect 2240 24750 2268 25094
rect 2228 24744 2280 24750
rect 2228 24686 2280 24692
rect 2320 24268 2372 24274
rect 2424 24256 2452 25298
rect 2372 24228 2452 24256
rect 2320 24210 2372 24216
rect 2136 24200 2188 24206
rect 2136 24142 2188 24148
rect 1964 23854 2084 23882
rect 1860 23588 1912 23594
rect 1860 23530 1912 23536
rect 1124 23520 1176 23526
rect 1124 23462 1176 23468
rect 1492 23520 1544 23526
rect 1492 23462 1544 23468
rect 1136 23186 1164 23462
rect 1124 23180 1176 23186
rect 1124 23122 1176 23128
rect 848 23112 900 23118
rect 848 23054 900 23060
rect 860 21486 888 23054
rect 1400 21888 1452 21894
rect 1400 21830 1452 21836
rect 848 21480 900 21486
rect 848 21422 900 21428
rect 860 20942 888 21422
rect 940 21412 992 21418
rect 940 21354 992 21360
rect 952 21146 980 21354
rect 1412 21146 1440 21830
rect 940 21140 992 21146
rect 940 21082 992 21088
rect 1400 21140 1452 21146
rect 1400 21082 1452 21088
rect 848 20936 900 20942
rect 848 20878 900 20884
rect 860 19854 888 20878
rect 1216 20256 1268 20262
rect 1216 20198 1268 20204
rect 1124 19916 1176 19922
rect 1124 19858 1176 19864
rect 848 19848 900 19854
rect 848 19790 900 19796
rect 860 17746 888 19790
rect 1136 19514 1164 19858
rect 1124 19508 1176 19514
rect 1124 19450 1176 19456
rect 1228 19310 1256 20198
rect 1504 19514 1532 23462
rect 1964 21690 1992 23854
rect 2044 23792 2096 23798
rect 2044 23734 2096 23740
rect 1584 21684 1636 21690
rect 1584 21626 1636 21632
rect 1952 21684 2004 21690
rect 1952 21626 2004 21632
rect 1596 21078 1624 21626
rect 2056 21622 2084 23734
rect 2148 23594 2176 24142
rect 2332 23866 2360 24210
rect 2516 24154 2544 29446
rect 2688 27872 2740 27878
rect 2688 27814 2740 27820
rect 2700 27334 2728 27814
rect 2688 27328 2740 27334
rect 2688 27270 2740 27276
rect 2792 27282 2820 30058
rect 2976 30054 3004 30110
rect 2964 30048 3016 30054
rect 2964 29990 3016 29996
rect 3252 29782 3280 30126
rect 4344 30116 4396 30122
rect 4344 30058 4396 30064
rect 3424 30048 3476 30054
rect 3424 29990 3476 29996
rect 3240 29776 3292 29782
rect 3240 29718 3292 29724
rect 3332 29708 3384 29714
rect 3332 29650 3384 29656
rect 3344 28762 3372 29650
rect 3056 28756 3108 28762
rect 3056 28698 3108 28704
rect 3332 28756 3384 28762
rect 3332 28698 3384 28704
rect 2872 28416 2924 28422
rect 2872 28358 2924 28364
rect 2884 27878 2912 28358
rect 2872 27872 2924 27878
rect 2872 27814 2924 27820
rect 3068 27470 3096 28698
rect 3240 28008 3292 28014
rect 3240 27950 3292 27956
rect 3148 27940 3200 27946
rect 3148 27882 3200 27888
rect 3160 27554 3188 27882
rect 3252 27674 3280 27950
rect 3332 27872 3384 27878
rect 3332 27814 3384 27820
rect 3240 27668 3292 27674
rect 3240 27610 3292 27616
rect 3160 27538 3280 27554
rect 3160 27532 3292 27538
rect 3160 27526 3240 27532
rect 3240 27474 3292 27480
rect 3056 27464 3108 27470
rect 3056 27406 3108 27412
rect 3148 27328 3200 27334
rect 2792 27254 3004 27282
rect 3148 27270 3200 27276
rect 2780 27124 2832 27130
rect 2780 27066 2832 27072
rect 2792 26586 2820 27066
rect 2780 26580 2832 26586
rect 2780 26522 2832 26528
rect 2780 25968 2832 25974
rect 2780 25910 2832 25916
rect 2688 25900 2740 25906
rect 2688 25842 2740 25848
rect 2596 25696 2648 25702
rect 2596 25638 2648 25644
rect 2608 24954 2636 25638
rect 2700 25498 2728 25842
rect 2688 25492 2740 25498
rect 2688 25434 2740 25440
rect 2688 25152 2740 25158
rect 2688 25094 2740 25100
rect 2596 24948 2648 24954
rect 2596 24890 2648 24896
rect 2596 24812 2648 24818
rect 2596 24754 2648 24760
rect 2608 24342 2636 24754
rect 2700 24682 2728 25094
rect 2792 24818 2820 25910
rect 2872 25832 2924 25838
rect 2872 25774 2924 25780
rect 2884 24954 2912 25774
rect 2872 24948 2924 24954
rect 2872 24890 2924 24896
rect 2780 24812 2832 24818
rect 2780 24754 2832 24760
rect 2688 24676 2740 24682
rect 2688 24618 2740 24624
rect 2596 24336 2648 24342
rect 2596 24278 2648 24284
rect 2424 24126 2544 24154
rect 2320 23860 2372 23866
rect 2320 23802 2372 23808
rect 2136 23588 2188 23594
rect 2136 23530 2188 23536
rect 2320 23520 2372 23526
rect 2320 23462 2372 23468
rect 2332 22778 2360 23462
rect 2320 22772 2372 22778
rect 2320 22714 2372 22720
rect 2424 22658 2452 24126
rect 2608 23866 2636 24278
rect 2872 24268 2924 24274
rect 2872 24210 2924 24216
rect 2688 24064 2740 24070
rect 2688 24006 2740 24012
rect 2780 24064 2832 24070
rect 2780 24006 2832 24012
rect 2596 23860 2648 23866
rect 2596 23802 2648 23808
rect 2504 23520 2556 23526
rect 2504 23462 2556 23468
rect 2148 22630 2452 22658
rect 2044 21616 2096 21622
rect 2044 21558 2096 21564
rect 1584 21072 1636 21078
rect 1584 21014 1636 21020
rect 1596 20330 1624 21014
rect 2056 20466 2084 21558
rect 2044 20460 2096 20466
rect 2044 20402 2096 20408
rect 1584 20324 1636 20330
rect 1584 20266 1636 20272
rect 1492 19508 1544 19514
rect 1492 19450 1544 19456
rect 1216 19304 1268 19310
rect 1216 19246 1268 19252
rect 1308 18216 1360 18222
rect 1308 18158 1360 18164
rect 1124 18080 1176 18086
rect 1124 18022 1176 18028
rect 1136 17814 1164 18022
rect 1124 17808 1176 17814
rect 1124 17750 1176 17756
rect 848 17740 900 17746
rect 848 17682 900 17688
rect 1320 17338 1348 18158
rect 1504 17338 1532 19450
rect 1308 17332 1360 17338
rect 1308 17274 1360 17280
rect 1492 17332 1544 17338
rect 1492 17274 1544 17280
rect 1596 16794 1624 20266
rect 1860 20256 1912 20262
rect 1860 20198 1912 20204
rect 1872 19310 1900 20198
rect 2056 19922 2084 20402
rect 2044 19916 2096 19922
rect 2044 19858 2096 19864
rect 2044 19440 2096 19446
rect 2044 19382 2096 19388
rect 1860 19304 1912 19310
rect 1860 19246 1912 19252
rect 2056 18222 2084 19382
rect 2044 18216 2096 18222
rect 2044 18158 2096 18164
rect 1860 18080 1912 18086
rect 1860 18022 1912 18028
rect 1952 18080 2004 18086
rect 1952 18022 2004 18028
rect 1872 17270 1900 18022
rect 1860 17264 1912 17270
rect 1860 17206 1912 17212
rect 1872 16998 1900 17206
rect 1964 17066 1992 18022
rect 1952 17060 2004 17066
rect 1952 17002 2004 17008
rect 1860 16992 1912 16998
rect 1860 16934 1912 16940
rect 1584 16788 1636 16794
rect 1584 16730 1636 16736
rect 1872 16266 1900 16934
rect 1872 16238 1992 16266
rect 1860 16108 1912 16114
rect 1860 16050 1912 16056
rect 1492 15904 1544 15910
rect 1492 15846 1544 15852
rect 1504 15570 1532 15846
rect 1674 15600 1730 15609
rect 1492 15564 1544 15570
rect 1872 15570 1900 16050
rect 1964 16046 1992 16238
rect 1952 16040 2004 16046
rect 1952 15982 2004 15988
rect 1674 15535 1676 15544
rect 1492 15506 1544 15512
rect 1728 15535 1730 15544
rect 1860 15564 1912 15570
rect 1676 15506 1728 15512
rect 1860 15506 1912 15512
rect 1400 15428 1452 15434
rect 1400 15370 1452 15376
rect 1216 15360 1268 15366
rect 1216 15302 1268 15308
rect 1228 14890 1256 15302
rect 1412 14958 1440 15370
rect 1400 14952 1452 14958
rect 1400 14894 1452 14900
rect 1216 14884 1268 14890
rect 1216 14826 1268 14832
rect 1412 13870 1440 14894
rect 1688 14550 1716 15506
rect 1872 14770 1900 15506
rect 1872 14742 1992 14770
rect 1676 14544 1728 14550
rect 1676 14486 1728 14492
rect 1584 14272 1636 14278
rect 1584 14214 1636 14220
rect 1400 13864 1452 13870
rect 1400 13806 1452 13812
rect 1308 13796 1360 13802
rect 1308 13738 1360 13744
rect 1320 13530 1348 13738
rect 1308 13524 1360 13530
rect 1308 13466 1360 13472
rect 1412 12374 1440 13806
rect 1596 12782 1624 14214
rect 1768 13728 1820 13734
rect 1768 13670 1820 13676
rect 1676 12912 1728 12918
rect 1676 12854 1728 12860
rect 1584 12776 1636 12782
rect 1584 12718 1636 12724
rect 1400 12368 1452 12374
rect 1400 12310 1452 12316
rect 1124 12300 1176 12306
rect 1124 12242 1176 12248
rect 1136 11898 1164 12242
rect 1124 11892 1176 11898
rect 1124 11834 1176 11840
rect 1400 11688 1452 11694
rect 1400 11630 1452 11636
rect 1412 11354 1440 11630
rect 1400 11348 1452 11354
rect 1400 11290 1452 11296
rect 1688 11218 1716 12854
rect 1780 12850 1808 13670
rect 1860 13320 1912 13326
rect 1860 13262 1912 13268
rect 1872 12986 1900 13262
rect 1860 12980 1912 12986
rect 1860 12922 1912 12928
rect 1964 12866 1992 14742
rect 2044 14612 2096 14618
rect 2044 14554 2096 14560
rect 2056 12918 2084 14554
rect 1872 12850 1992 12866
rect 2044 12912 2096 12918
rect 2044 12854 2096 12860
rect 1768 12844 1820 12850
rect 1768 12786 1820 12792
rect 1860 12844 1992 12850
rect 1912 12838 1992 12844
rect 1860 12786 1912 12792
rect 2148 12442 2176 22630
rect 2228 22094 2280 22098
rect 2516 22094 2544 23462
rect 2608 23186 2636 23802
rect 2700 23594 2728 24006
rect 2792 23730 2820 24006
rect 2780 23724 2832 23730
rect 2780 23666 2832 23672
rect 2688 23588 2740 23594
rect 2688 23530 2740 23536
rect 2792 23254 2820 23666
rect 2884 23594 2912 24210
rect 2872 23588 2924 23594
rect 2872 23530 2924 23536
rect 2884 23322 2912 23530
rect 2872 23316 2924 23322
rect 2872 23258 2924 23264
rect 2780 23248 2832 23254
rect 2780 23190 2832 23196
rect 2596 23180 2648 23186
rect 2596 23122 2648 23128
rect 2608 22574 2636 23122
rect 2884 22574 2912 23258
rect 2596 22568 2648 22574
rect 2596 22510 2648 22516
rect 2872 22568 2924 22574
rect 2872 22510 2924 22516
rect 2688 22432 2740 22438
rect 2688 22374 2740 22380
rect 2228 22092 2544 22094
rect 2280 22066 2544 22092
rect 2228 22034 2280 22040
rect 2412 20800 2464 20806
rect 2412 20742 2464 20748
rect 2320 20596 2372 20602
rect 2320 20538 2372 20544
rect 2228 20392 2280 20398
rect 2228 20334 2280 20340
rect 2240 20058 2268 20334
rect 2332 20058 2360 20538
rect 2424 20398 2452 20742
rect 2412 20392 2464 20398
rect 2412 20334 2464 20340
rect 2516 20262 2544 22066
rect 2596 22094 2648 22098
rect 2700 22094 2728 22374
rect 2596 22092 2728 22094
rect 2648 22066 2728 22092
rect 2596 22034 2648 22040
rect 2608 21350 2636 22034
rect 2976 21570 3004 27254
rect 3056 26988 3108 26994
rect 3056 26930 3108 26936
rect 3068 26450 3096 26930
rect 3160 26450 3188 27270
rect 3252 26994 3280 27474
rect 3344 27470 3372 27814
rect 3332 27464 3384 27470
rect 3332 27406 3384 27412
rect 3240 26988 3292 26994
rect 3240 26930 3292 26936
rect 3056 26444 3108 26450
rect 3056 26386 3108 26392
rect 3148 26444 3200 26450
rect 3148 26386 3200 26392
rect 3344 26314 3372 27406
rect 3332 26308 3384 26314
rect 3332 26250 3384 26256
rect 3240 25764 3292 25770
rect 3240 25706 3292 25712
rect 3056 25696 3108 25702
rect 3056 25638 3108 25644
rect 3068 25362 3096 25638
rect 3056 25356 3108 25362
rect 3056 25298 3108 25304
rect 3056 24812 3108 24818
rect 3056 24754 3108 24760
rect 3068 23186 3096 24754
rect 3056 23180 3108 23186
rect 3056 23122 3108 23128
rect 3148 22500 3200 22506
rect 3148 22442 3200 22448
rect 3160 22030 3188 22442
rect 3148 22024 3200 22030
rect 3148 21966 3200 21972
rect 2976 21542 3188 21570
rect 2964 21412 3016 21418
rect 2964 21354 3016 21360
rect 2596 21344 2648 21350
rect 2596 21286 2648 21292
rect 2688 21344 2740 21350
rect 2688 21286 2740 21292
rect 2872 21344 2924 21350
rect 2872 21286 2924 21292
rect 2608 20482 2636 21286
rect 2700 20602 2728 21286
rect 2884 21010 2912 21286
rect 2872 21004 2924 21010
rect 2872 20946 2924 20952
rect 2780 20936 2832 20942
rect 2780 20878 2832 20884
rect 2688 20596 2740 20602
rect 2688 20538 2740 20544
rect 2608 20454 2728 20482
rect 2700 20398 2728 20454
rect 2688 20392 2740 20398
rect 2688 20334 2740 20340
rect 2792 20330 2820 20878
rect 2976 20874 3004 21354
rect 2964 20868 3016 20874
rect 2964 20810 3016 20816
rect 2780 20324 2832 20330
rect 2780 20266 2832 20272
rect 2504 20256 2556 20262
rect 2504 20198 2556 20204
rect 2228 20052 2280 20058
rect 2228 19994 2280 20000
rect 2320 20052 2372 20058
rect 2320 19994 2372 20000
rect 2688 19916 2740 19922
rect 2688 19858 2740 19864
rect 2780 19916 2832 19922
rect 2780 19858 2832 19864
rect 2504 19236 2556 19242
rect 2504 19178 2556 19184
rect 2516 18970 2544 19178
rect 2700 19174 2728 19858
rect 2792 19514 2820 19858
rect 2964 19712 3016 19718
rect 2964 19654 3016 19660
rect 2780 19508 2832 19514
rect 2780 19450 2832 19456
rect 2688 19168 2740 19174
rect 2688 19110 2740 19116
rect 2504 18964 2556 18970
rect 2504 18906 2556 18912
rect 2976 18902 3004 19654
rect 2964 18896 3016 18902
rect 2964 18838 3016 18844
rect 2228 18216 2280 18222
rect 2228 18158 2280 18164
rect 2240 17882 2268 18158
rect 2688 18148 2740 18154
rect 2688 18090 2740 18096
rect 2228 17876 2280 17882
rect 2228 17818 2280 17824
rect 2700 17678 2728 18090
rect 3056 17740 3108 17746
rect 3056 17682 3108 17688
rect 2504 17672 2556 17678
rect 2504 17614 2556 17620
rect 2688 17672 2740 17678
rect 2688 17614 2740 17620
rect 2516 17354 2544 17614
rect 2872 17536 2924 17542
rect 2872 17478 2924 17484
rect 2228 17332 2280 17338
rect 2424 17326 2544 17354
rect 2424 17320 2452 17326
rect 2280 17292 2452 17320
rect 2228 17274 2280 17280
rect 2240 16182 2268 17274
rect 2504 17264 2556 17270
rect 2504 17206 2556 17212
rect 2412 16788 2464 16794
rect 2412 16730 2464 16736
rect 2228 16176 2280 16182
rect 2228 16118 2280 16124
rect 2424 16046 2452 16730
rect 2516 16658 2544 17206
rect 2688 17196 2740 17202
rect 2688 17138 2740 17144
rect 2700 16794 2728 17138
rect 2884 17066 2912 17478
rect 3068 17338 3096 17682
rect 3056 17332 3108 17338
rect 3056 17274 3108 17280
rect 3160 17218 3188 21542
rect 3252 21146 3280 25706
rect 3332 23112 3384 23118
rect 3332 23054 3384 23060
rect 3344 22778 3372 23054
rect 3332 22772 3384 22778
rect 3332 22714 3384 22720
rect 3436 22094 3464 29990
rect 4356 29850 4384 30058
rect 4344 29844 4396 29850
rect 4344 29786 4396 29792
rect 5552 29782 5580 30126
rect 3516 29776 3568 29782
rect 3516 29718 3568 29724
rect 5540 29776 5592 29782
rect 5540 29718 5592 29724
rect 3528 29170 3556 29718
rect 4160 29708 4212 29714
rect 4160 29650 4212 29656
rect 3608 29504 3660 29510
rect 3608 29446 3660 29452
rect 3516 29164 3568 29170
rect 3516 29106 3568 29112
rect 3528 28694 3556 29106
rect 3620 29102 3648 29446
rect 3756 29404 4064 29413
rect 3756 29402 3762 29404
rect 3818 29402 3842 29404
rect 3898 29402 3922 29404
rect 3978 29402 4002 29404
rect 4058 29402 4064 29404
rect 3818 29350 3820 29402
rect 4000 29350 4002 29402
rect 3756 29348 3762 29350
rect 3818 29348 3842 29350
rect 3898 29348 3922 29350
rect 3978 29348 4002 29350
rect 4058 29348 4064 29350
rect 3756 29339 4064 29348
rect 3608 29096 3660 29102
rect 3608 29038 3660 29044
rect 4172 28762 4200 29650
rect 5644 29102 5672 30738
rect 5828 30122 5856 31600
rect 7300 31498 7328 31600
rect 7392 31498 7420 31606
rect 7300 31470 7420 31498
rect 7114 31036 7422 31045
rect 7114 31034 7120 31036
rect 7176 31034 7200 31036
rect 7256 31034 7280 31036
rect 7336 31034 7360 31036
rect 7416 31034 7422 31036
rect 7176 30982 7178 31034
rect 7358 30982 7360 31034
rect 7114 30980 7120 30982
rect 7176 30980 7200 30982
rect 7256 30980 7280 30982
rect 7336 30980 7360 30982
rect 7416 30980 7422 30982
rect 7114 30971 7422 30980
rect 7576 30802 7604 31606
rect 8758 31600 8814 32000
rect 10230 31600 10286 32000
rect 11702 31600 11758 32000
rect 13174 31600 13230 32000
rect 14646 31600 14702 32000
rect 16118 31600 16174 32000
rect 17590 31600 17646 32000
rect 17696 31606 18000 31634
rect 8772 30802 8800 31600
rect 10140 30864 10192 30870
rect 10140 30806 10192 30812
rect 7564 30796 7616 30802
rect 7564 30738 7616 30744
rect 8760 30796 8812 30802
rect 8760 30738 8812 30744
rect 6920 30728 6972 30734
rect 6840 30676 6920 30682
rect 6840 30670 6972 30676
rect 8024 30728 8076 30734
rect 8024 30670 8076 30676
rect 6368 30660 6420 30666
rect 6368 30602 6420 30608
rect 6840 30654 6960 30670
rect 6276 30592 6328 30598
rect 6276 30534 6328 30540
rect 5816 30116 5868 30122
rect 5816 30058 5868 30064
rect 6092 30048 6144 30054
rect 6092 29990 6144 29996
rect 6000 29708 6052 29714
rect 6000 29650 6052 29656
rect 5816 29640 5868 29646
rect 5816 29582 5868 29588
rect 5724 29232 5776 29238
rect 5724 29174 5776 29180
rect 5736 29102 5764 29174
rect 5632 29096 5684 29102
rect 5632 29038 5684 29044
rect 5724 29096 5776 29102
rect 5724 29038 5776 29044
rect 5356 29028 5408 29034
rect 5356 28970 5408 28976
rect 4988 28960 5040 28966
rect 4988 28902 5040 28908
rect 5000 28762 5028 28902
rect 4160 28756 4212 28762
rect 4160 28698 4212 28704
rect 4988 28756 5040 28762
rect 4988 28698 5040 28704
rect 3516 28688 3568 28694
rect 3516 28630 3568 28636
rect 5368 28626 5396 28970
rect 5540 28960 5592 28966
rect 5540 28902 5592 28908
rect 5632 28960 5684 28966
rect 5632 28902 5684 28908
rect 3608 28620 3660 28626
rect 3608 28562 3660 28568
rect 5356 28620 5408 28626
rect 5356 28562 5408 28568
rect 3620 28218 3648 28562
rect 3756 28316 4064 28325
rect 3756 28314 3762 28316
rect 3818 28314 3842 28316
rect 3898 28314 3922 28316
rect 3978 28314 4002 28316
rect 4058 28314 4064 28316
rect 3818 28262 3820 28314
rect 4000 28262 4002 28314
rect 3756 28260 3762 28262
rect 3818 28260 3842 28262
rect 3898 28260 3922 28262
rect 3978 28260 4002 28262
rect 4058 28260 4064 28262
rect 3756 28251 4064 28260
rect 3608 28212 3660 28218
rect 3608 28154 3660 28160
rect 5368 28014 5396 28562
rect 4160 28008 4212 28014
rect 4160 27950 4212 27956
rect 5356 28008 5408 28014
rect 5356 27950 5408 27956
rect 3884 27872 3936 27878
rect 3884 27814 3936 27820
rect 3896 27606 3924 27814
rect 3884 27600 3936 27606
rect 3884 27542 3936 27548
rect 3608 27532 3660 27538
rect 3608 27474 3660 27480
rect 3516 26376 3568 26382
rect 3516 26318 3568 26324
rect 3528 24750 3556 26318
rect 3620 25770 3648 27474
rect 3756 27228 4064 27237
rect 3756 27226 3762 27228
rect 3818 27226 3842 27228
rect 3898 27226 3922 27228
rect 3978 27226 4002 27228
rect 4058 27226 4064 27228
rect 3818 27174 3820 27226
rect 4000 27174 4002 27226
rect 3756 27172 3762 27174
rect 3818 27172 3842 27174
rect 3898 27172 3922 27174
rect 3978 27172 4002 27174
rect 4058 27172 4064 27174
rect 3756 27163 4064 27172
rect 4172 27130 4200 27950
rect 5368 27538 5396 27950
rect 5356 27532 5408 27538
rect 5356 27474 5408 27480
rect 4896 27328 4948 27334
rect 4896 27270 4948 27276
rect 5172 27328 5224 27334
rect 5172 27270 5224 27276
rect 4160 27124 4212 27130
rect 4160 27066 4212 27072
rect 4908 26908 4936 27270
rect 5184 27062 5212 27270
rect 5172 27056 5224 27062
rect 5172 26998 5224 27004
rect 5368 26994 5396 27474
rect 5356 26988 5408 26994
rect 5356 26930 5408 26936
rect 4988 26920 5040 26926
rect 4908 26880 4988 26908
rect 4344 26444 4396 26450
rect 4344 26386 4396 26392
rect 4160 26308 4212 26314
rect 4160 26250 4212 26256
rect 3756 26140 4064 26149
rect 3756 26138 3762 26140
rect 3818 26138 3842 26140
rect 3898 26138 3922 26140
rect 3978 26138 4002 26140
rect 4058 26138 4064 26140
rect 3818 26086 3820 26138
rect 4000 26086 4002 26138
rect 3756 26084 3762 26086
rect 3818 26084 3842 26086
rect 3898 26084 3922 26086
rect 3978 26084 4002 26086
rect 4058 26084 4064 26086
rect 3756 26075 4064 26084
rect 4172 25922 4200 26250
rect 4080 25894 4200 25922
rect 3608 25764 3660 25770
rect 3608 25706 3660 25712
rect 3620 25430 3648 25706
rect 3608 25424 3660 25430
rect 3608 25366 3660 25372
rect 3516 24744 3568 24750
rect 3516 24686 3568 24692
rect 3620 24138 3648 25366
rect 4080 25140 4108 25894
rect 4252 25696 4304 25702
rect 4252 25638 4304 25644
rect 4080 25112 4200 25140
rect 3756 25052 4064 25061
rect 3756 25050 3762 25052
rect 3818 25050 3842 25052
rect 3898 25050 3922 25052
rect 3978 25050 4002 25052
rect 4058 25050 4064 25052
rect 3818 24998 3820 25050
rect 4000 24998 4002 25050
rect 3756 24996 3762 24998
rect 3818 24996 3842 24998
rect 3898 24996 3922 24998
rect 3978 24996 4002 24998
rect 4058 24996 4064 24998
rect 3756 24987 4064 24996
rect 4172 24954 4200 25112
rect 4160 24948 4212 24954
rect 4160 24890 4212 24896
rect 3608 24132 3660 24138
rect 3608 24074 3660 24080
rect 4160 24064 4212 24070
rect 4160 24006 4212 24012
rect 3756 23964 4064 23973
rect 3756 23962 3762 23964
rect 3818 23962 3842 23964
rect 3898 23962 3922 23964
rect 3978 23962 4002 23964
rect 4058 23962 4064 23964
rect 3818 23910 3820 23962
rect 4000 23910 4002 23962
rect 3756 23908 3762 23910
rect 3818 23908 3842 23910
rect 3898 23908 3922 23910
rect 3978 23908 4002 23910
rect 4058 23908 4064 23910
rect 3756 23899 4064 23908
rect 3792 23656 3844 23662
rect 3790 23624 3792 23633
rect 3884 23656 3936 23662
rect 3844 23624 3846 23633
rect 3700 23588 3752 23594
rect 4172 23644 4200 24006
rect 3936 23616 4200 23644
rect 3884 23598 3936 23604
rect 3790 23559 3846 23568
rect 3700 23530 3752 23536
rect 3712 23186 3740 23530
rect 3804 23322 3832 23559
rect 3792 23316 3844 23322
rect 3792 23258 3844 23264
rect 4172 23254 4200 23616
rect 4160 23248 4212 23254
rect 4160 23190 4212 23196
rect 3700 23180 3752 23186
rect 3700 23122 3752 23128
rect 3608 23112 3660 23118
rect 3608 23054 3660 23060
rect 3516 23044 3568 23050
rect 3516 22986 3568 22992
rect 3528 22234 3556 22986
rect 3620 22778 3648 23054
rect 3756 22876 4064 22885
rect 3756 22874 3762 22876
rect 3818 22874 3842 22876
rect 3898 22874 3922 22876
rect 3978 22874 4002 22876
rect 4058 22874 4064 22876
rect 3818 22822 3820 22874
rect 4000 22822 4002 22874
rect 3756 22820 3762 22822
rect 3818 22820 3842 22822
rect 3898 22820 3922 22822
rect 3978 22820 4002 22822
rect 4058 22820 4064 22822
rect 3756 22811 4064 22820
rect 3608 22772 3660 22778
rect 3608 22714 3660 22720
rect 4264 22438 4292 25638
rect 4356 23662 4384 26386
rect 4620 26240 4672 26246
rect 4620 26182 4672 26188
rect 4436 25832 4488 25838
rect 4436 25774 4488 25780
rect 4448 25498 4476 25774
rect 4436 25492 4488 25498
rect 4436 25434 4488 25440
rect 4632 25158 4660 26182
rect 4908 25294 4936 26880
rect 4988 26862 5040 26868
rect 5552 26790 5580 28902
rect 5644 28422 5672 28902
rect 5632 28416 5684 28422
rect 5632 28358 5684 28364
rect 5736 28014 5764 29038
rect 5828 28762 5856 29582
rect 5816 28756 5868 28762
rect 5816 28698 5868 28704
rect 5724 28008 5776 28014
rect 5724 27950 5776 27956
rect 5736 27606 5764 27950
rect 5908 27872 5960 27878
rect 5908 27814 5960 27820
rect 5724 27600 5776 27606
rect 5724 27542 5776 27548
rect 5632 27464 5684 27470
rect 5632 27406 5684 27412
rect 5644 27130 5672 27406
rect 5736 27130 5764 27542
rect 5920 27538 5948 27814
rect 5908 27532 5960 27538
rect 5908 27474 5960 27480
rect 5816 27328 5868 27334
rect 5816 27270 5868 27276
rect 5632 27124 5684 27130
rect 5632 27066 5684 27072
rect 5724 27124 5776 27130
rect 5724 27066 5776 27072
rect 5540 26784 5592 26790
rect 5540 26726 5592 26732
rect 5644 26586 5672 27066
rect 5724 26852 5776 26858
rect 5724 26794 5776 26800
rect 5632 26580 5684 26586
rect 5632 26522 5684 26528
rect 5448 26444 5500 26450
rect 5500 26404 5580 26432
rect 5448 26386 5500 26392
rect 4988 26240 5040 26246
rect 4988 26182 5040 26188
rect 5000 25906 5028 26182
rect 4988 25900 5040 25906
rect 4988 25842 5040 25848
rect 5080 25832 5132 25838
rect 5080 25774 5132 25780
rect 5172 25832 5224 25838
rect 5172 25774 5224 25780
rect 5092 25362 5120 25774
rect 4988 25356 5040 25362
rect 4988 25298 5040 25304
rect 5080 25356 5132 25362
rect 5080 25298 5132 25304
rect 4896 25288 4948 25294
rect 4896 25230 4948 25236
rect 4620 25152 4672 25158
rect 4620 25094 4672 25100
rect 4908 24750 4936 25230
rect 5000 24818 5028 25298
rect 5092 24954 5120 25298
rect 5080 24948 5132 24954
rect 5080 24890 5132 24896
rect 4988 24812 5040 24818
rect 4988 24754 5040 24760
rect 4896 24744 4948 24750
rect 4896 24686 4948 24692
rect 4804 24268 4856 24274
rect 4804 24210 4856 24216
rect 4816 23866 4844 24210
rect 4896 24064 4948 24070
rect 4896 24006 4948 24012
rect 4804 23860 4856 23866
rect 4804 23802 4856 23808
rect 4528 23724 4580 23730
rect 4528 23666 4580 23672
rect 4344 23656 4396 23662
rect 4344 23598 4396 23604
rect 4356 23186 4384 23598
rect 4540 23594 4568 23666
rect 4908 23662 4936 24006
rect 5184 23866 5212 25774
rect 5552 25498 5580 26404
rect 5540 25492 5592 25498
rect 5540 25434 5592 25440
rect 5356 25288 5408 25294
rect 5356 25230 5408 25236
rect 5368 24954 5396 25230
rect 5356 24948 5408 24954
rect 5356 24890 5408 24896
rect 5736 24426 5764 26794
rect 5828 26450 5856 27270
rect 5908 26784 5960 26790
rect 5908 26726 5960 26732
rect 5816 26444 5868 26450
rect 5816 26386 5868 26392
rect 5920 26353 5948 26726
rect 5906 26344 5962 26353
rect 5906 26279 5962 26288
rect 5552 24398 5764 24426
rect 5448 24132 5500 24138
rect 5448 24074 5500 24080
rect 5172 23860 5224 23866
rect 5172 23802 5224 23808
rect 5356 23860 5408 23866
rect 5356 23802 5408 23808
rect 4896 23656 4948 23662
rect 4988 23656 5040 23662
rect 4896 23598 4948 23604
rect 4986 23624 4988 23633
rect 5080 23656 5132 23662
rect 5040 23624 5042 23633
rect 4528 23588 4580 23594
rect 4448 23548 4528 23576
rect 4344 23180 4396 23186
rect 4344 23122 4396 23128
rect 4448 23118 4476 23548
rect 5080 23598 5132 23604
rect 4986 23559 5042 23568
rect 4528 23530 4580 23536
rect 4620 23520 4672 23526
rect 4672 23480 4844 23508
rect 4620 23462 4672 23468
rect 4816 23186 4844 23480
rect 5092 23322 5120 23598
rect 5080 23316 5132 23322
rect 5080 23258 5132 23264
rect 4804 23180 4856 23186
rect 4804 23122 4856 23128
rect 4436 23112 4488 23118
rect 4436 23054 4488 23060
rect 4528 22976 4580 22982
rect 4528 22918 4580 22924
rect 4540 22574 4568 22918
rect 5264 22772 5316 22778
rect 5264 22714 5316 22720
rect 4620 22704 4672 22710
rect 4620 22646 4672 22652
rect 4528 22568 4580 22574
rect 4528 22510 4580 22516
rect 4252 22432 4304 22438
rect 4252 22374 4304 22380
rect 3516 22228 3568 22234
rect 3516 22170 3568 22176
rect 3436 22066 3556 22094
rect 3332 22024 3384 22030
rect 3332 21966 3384 21972
rect 3344 21350 3372 21966
rect 3332 21344 3384 21350
rect 3332 21286 3384 21292
rect 3240 21140 3292 21146
rect 3240 21082 3292 21088
rect 3344 21010 3372 21286
rect 3332 21004 3384 21010
rect 3332 20946 3384 20952
rect 3332 20392 3384 20398
rect 3332 20334 3384 20340
rect 3344 19922 3372 20334
rect 3332 19916 3384 19922
rect 3332 19858 3384 19864
rect 3344 19514 3372 19858
rect 3332 19508 3384 19514
rect 3332 19450 3384 19456
rect 3240 17604 3292 17610
rect 3240 17546 3292 17552
rect 3252 17338 3280 17546
rect 3332 17536 3384 17542
rect 3332 17478 3384 17484
rect 3240 17332 3292 17338
rect 3240 17274 3292 17280
rect 3068 17190 3188 17218
rect 2872 17060 2924 17066
rect 2872 17002 2924 17008
rect 2688 16788 2740 16794
rect 2688 16730 2740 16736
rect 2504 16652 2556 16658
rect 2504 16594 2556 16600
rect 2596 16516 2648 16522
rect 2596 16458 2648 16464
rect 2504 16448 2556 16454
rect 2504 16390 2556 16396
rect 2516 16182 2544 16390
rect 2504 16176 2556 16182
rect 2504 16118 2556 16124
rect 2516 16046 2544 16118
rect 2412 16040 2464 16046
rect 2412 15982 2464 15988
rect 2504 16040 2556 16046
rect 2504 15982 2556 15988
rect 2516 15162 2544 15982
rect 2608 15570 2636 16458
rect 2596 15564 2648 15570
rect 2596 15506 2648 15512
rect 2608 15366 2636 15506
rect 2596 15360 2648 15366
rect 2596 15302 2648 15308
rect 2504 15156 2556 15162
rect 2504 15098 2556 15104
rect 2228 14272 2280 14278
rect 2964 14272 3016 14278
rect 2228 14214 2280 14220
rect 2884 14232 2964 14260
rect 2240 14074 2268 14214
rect 2228 14068 2280 14074
rect 2228 14010 2280 14016
rect 2320 13252 2372 13258
rect 2320 13194 2372 13200
rect 2332 12782 2360 13194
rect 2688 13184 2740 13190
rect 2688 13126 2740 13132
rect 2320 12776 2372 12782
rect 2320 12718 2372 12724
rect 2228 12640 2280 12646
rect 2228 12582 2280 12588
rect 2136 12436 2188 12442
rect 2136 12378 2188 12384
rect 2240 12102 2268 12582
rect 2228 12096 2280 12102
rect 2228 12038 2280 12044
rect 2240 11762 2268 12038
rect 2228 11756 2280 11762
rect 2228 11698 2280 11704
rect 1860 11552 1912 11558
rect 1860 11494 1912 11500
rect 1872 11218 1900 11494
rect 1676 11212 1728 11218
rect 1676 11154 1728 11160
rect 1860 11212 1912 11218
rect 1860 11154 1912 11160
rect 2332 11150 2360 12718
rect 2596 12640 2648 12646
rect 2596 12582 2648 12588
rect 2608 12374 2636 12582
rect 2596 12368 2648 12374
rect 2596 12310 2648 12316
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 2700 11014 2728 13126
rect 2780 12776 2832 12782
rect 2780 12718 2832 12724
rect 2792 11082 2820 12718
rect 2884 12714 2912 14232
rect 2964 14214 3016 14220
rect 2964 12912 3016 12918
rect 2964 12854 3016 12860
rect 2872 12708 2924 12714
rect 2872 12650 2924 12656
rect 2780 11076 2832 11082
rect 2780 11018 2832 11024
rect 2504 11008 2556 11014
rect 2504 10950 2556 10956
rect 2688 11008 2740 11014
rect 2688 10950 2740 10956
rect 2320 10464 2372 10470
rect 2320 10406 2372 10412
rect 2332 10062 2360 10406
rect 2320 10056 2372 10062
rect 2318 10024 2320 10033
rect 2372 10024 2374 10033
rect 2318 9959 2374 9968
rect 2516 9518 2544 10950
rect 2976 10674 3004 12854
rect 2964 10668 3016 10674
rect 2964 10610 3016 10616
rect 2596 10600 2648 10606
rect 2596 10542 2648 10548
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 2608 10130 2636 10542
rect 2792 10282 2820 10542
rect 2964 10464 3016 10470
rect 2964 10406 3016 10412
rect 3068 10418 3096 17190
rect 3344 16658 3372 17478
rect 3332 16652 3384 16658
rect 3332 16594 3384 16600
rect 3332 16040 3384 16046
rect 3332 15982 3384 15988
rect 3344 15706 3372 15982
rect 3332 15700 3384 15706
rect 3332 15642 3384 15648
rect 3344 14618 3372 15642
rect 3332 14612 3384 14618
rect 3332 14554 3384 14560
rect 3344 14482 3372 14554
rect 3148 14476 3200 14482
rect 3148 14418 3200 14424
rect 3332 14476 3384 14482
rect 3332 14418 3384 14424
rect 3160 14074 3188 14418
rect 3148 14068 3200 14074
rect 3148 14010 3200 14016
rect 3160 13394 3188 14010
rect 3344 13530 3372 14418
rect 3424 13864 3476 13870
rect 3424 13806 3476 13812
rect 3332 13524 3384 13530
rect 3332 13466 3384 13472
rect 3436 13394 3464 13806
rect 3148 13388 3200 13394
rect 3148 13330 3200 13336
rect 3424 13388 3476 13394
rect 3424 13330 3476 13336
rect 3240 12640 3292 12646
rect 3240 12582 3292 12588
rect 3252 11354 3280 12582
rect 3424 12300 3476 12306
rect 3424 12242 3476 12248
rect 3436 11694 3464 12242
rect 3424 11688 3476 11694
rect 3424 11630 3476 11636
rect 3424 11552 3476 11558
rect 3424 11494 3476 11500
rect 3240 11348 3292 11354
rect 3240 11290 3292 11296
rect 3436 11150 3464 11494
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 3528 10810 3556 22066
rect 3756 21788 4064 21797
rect 3756 21786 3762 21788
rect 3818 21786 3842 21788
rect 3898 21786 3922 21788
rect 3978 21786 4002 21788
rect 4058 21786 4064 21788
rect 3818 21734 3820 21786
rect 4000 21734 4002 21786
rect 3756 21732 3762 21734
rect 3818 21732 3842 21734
rect 3898 21732 3922 21734
rect 3978 21732 4002 21734
rect 4058 21732 4064 21734
rect 3756 21723 4064 21732
rect 4252 21684 4304 21690
rect 4252 21626 4304 21632
rect 4160 21412 4212 21418
rect 4160 21354 4212 21360
rect 4172 20942 4200 21354
rect 4160 20936 4212 20942
rect 4160 20878 4212 20884
rect 3756 20700 4064 20709
rect 3756 20698 3762 20700
rect 3818 20698 3842 20700
rect 3898 20698 3922 20700
rect 3978 20698 4002 20700
rect 4058 20698 4064 20700
rect 3818 20646 3820 20698
rect 4000 20646 4002 20698
rect 3756 20644 3762 20646
rect 3818 20644 3842 20646
rect 3898 20644 3922 20646
rect 3978 20644 4002 20646
rect 4058 20644 4064 20646
rect 3756 20635 4064 20644
rect 4172 20466 4200 20878
rect 4160 20460 4212 20466
rect 4160 20402 4212 20408
rect 4264 20398 4292 21626
rect 4344 20936 4396 20942
rect 4344 20878 4396 20884
rect 4436 20936 4488 20942
rect 4436 20878 4488 20884
rect 4528 20936 4580 20942
rect 4528 20878 4580 20884
rect 4356 20534 4384 20878
rect 4344 20528 4396 20534
rect 4344 20470 4396 20476
rect 4252 20392 4304 20398
rect 4252 20334 4304 20340
rect 3792 20256 3844 20262
rect 3792 20198 3844 20204
rect 3700 19984 3752 19990
rect 3620 19944 3700 19972
rect 3620 19378 3648 19944
rect 3700 19926 3752 19932
rect 3804 19922 3832 20198
rect 4448 20058 4476 20878
rect 4540 20602 4568 20878
rect 4528 20596 4580 20602
rect 4528 20538 4580 20544
rect 4436 20052 4488 20058
rect 4436 19994 4488 20000
rect 3792 19916 3844 19922
rect 3792 19858 3844 19864
rect 4436 19848 4488 19854
rect 4436 19790 4488 19796
rect 4252 19780 4304 19786
rect 4252 19722 4304 19728
rect 3756 19612 4064 19621
rect 3756 19610 3762 19612
rect 3818 19610 3842 19612
rect 3898 19610 3922 19612
rect 3978 19610 4002 19612
rect 4058 19610 4064 19612
rect 3818 19558 3820 19610
rect 4000 19558 4002 19610
rect 3756 19556 3762 19558
rect 3818 19556 3842 19558
rect 3898 19556 3922 19558
rect 3978 19556 4002 19558
rect 4058 19556 4064 19558
rect 3756 19547 4064 19556
rect 4264 19514 4292 19722
rect 4448 19514 4476 19790
rect 4252 19508 4304 19514
rect 4252 19450 4304 19456
rect 4436 19508 4488 19514
rect 4436 19450 4488 19456
rect 3608 19372 3660 19378
rect 3608 19314 3660 19320
rect 4632 19310 4660 22646
rect 5172 22636 5224 22642
rect 5172 22578 5224 22584
rect 4988 22568 5040 22574
rect 4988 22510 5040 22516
rect 5000 22234 5028 22510
rect 5184 22234 5212 22578
rect 5276 22574 5304 22714
rect 5368 22642 5396 23802
rect 5460 23730 5488 24074
rect 5448 23724 5500 23730
rect 5448 23666 5500 23672
rect 5356 22636 5408 22642
rect 5356 22578 5408 22584
rect 5264 22568 5316 22574
rect 5264 22510 5316 22516
rect 4988 22228 5040 22234
rect 4988 22170 5040 22176
rect 5172 22228 5224 22234
rect 5172 22170 5224 22176
rect 4804 22092 4856 22098
rect 4804 22034 4856 22040
rect 5080 22092 5132 22098
rect 5080 22034 5132 22040
rect 4712 21344 4764 21350
rect 4712 21286 4764 21292
rect 4724 19922 4752 21286
rect 4816 21078 4844 22034
rect 4896 21344 4948 21350
rect 4896 21286 4948 21292
rect 4804 21072 4856 21078
rect 4804 21014 4856 21020
rect 4908 20874 4936 21286
rect 4896 20868 4948 20874
rect 4896 20810 4948 20816
rect 4896 20392 4948 20398
rect 4896 20334 4948 20340
rect 4712 19916 4764 19922
rect 4712 19858 4764 19864
rect 4908 19854 4936 20334
rect 5092 19922 5120 22034
rect 5356 22024 5408 22030
rect 5354 21992 5356 22001
rect 5408 21992 5410 22001
rect 5552 21962 5580 24398
rect 5920 23186 5948 26279
rect 5908 23180 5960 23186
rect 5828 23140 5908 23168
rect 5632 22568 5684 22574
rect 5632 22510 5684 22516
rect 5354 21927 5410 21936
rect 5540 21956 5592 21962
rect 5264 21072 5316 21078
rect 5264 21014 5316 21020
rect 5276 20602 5304 21014
rect 5368 20806 5396 21927
rect 5540 21898 5592 21904
rect 5448 21888 5500 21894
rect 5448 21830 5500 21836
rect 5460 21010 5488 21830
rect 5552 21622 5580 21898
rect 5540 21616 5592 21622
rect 5540 21558 5592 21564
rect 5540 21344 5592 21350
rect 5540 21286 5592 21292
rect 5448 21004 5500 21010
rect 5448 20946 5500 20952
rect 5356 20800 5408 20806
rect 5356 20742 5408 20748
rect 5264 20596 5316 20602
rect 5264 20538 5316 20544
rect 5460 20466 5488 20946
rect 5448 20460 5500 20466
rect 5448 20402 5500 20408
rect 5552 20330 5580 21286
rect 5644 21026 5672 22510
rect 5724 22432 5776 22438
rect 5724 22374 5776 22380
rect 5736 21128 5764 22374
rect 5828 21298 5856 23140
rect 5908 23122 5960 23128
rect 5908 22500 5960 22506
rect 5908 22442 5960 22448
rect 5920 21690 5948 22442
rect 5908 21684 5960 21690
rect 5908 21626 5960 21632
rect 5828 21270 5948 21298
rect 5736 21100 5856 21128
rect 5644 20998 5764 21026
rect 5736 20942 5764 20998
rect 5724 20936 5776 20942
rect 5724 20878 5776 20884
rect 5736 20398 5764 20878
rect 5724 20392 5776 20398
rect 5724 20334 5776 20340
rect 5540 20324 5592 20330
rect 5540 20266 5592 20272
rect 5080 19916 5132 19922
rect 5080 19858 5132 19864
rect 4896 19848 4948 19854
rect 4896 19790 4948 19796
rect 4620 19304 4672 19310
rect 4620 19246 4672 19252
rect 4620 19168 4672 19174
rect 4620 19110 4672 19116
rect 3756 18524 4064 18533
rect 3756 18522 3762 18524
rect 3818 18522 3842 18524
rect 3898 18522 3922 18524
rect 3978 18522 4002 18524
rect 4058 18522 4064 18524
rect 3818 18470 3820 18522
rect 4000 18470 4002 18522
rect 3756 18468 3762 18470
rect 3818 18468 3842 18470
rect 3898 18468 3922 18470
rect 3978 18468 4002 18470
rect 4058 18468 4064 18470
rect 3756 18459 4064 18468
rect 4528 18216 4580 18222
rect 4528 18158 4580 18164
rect 4540 17882 4568 18158
rect 4528 17876 4580 17882
rect 4528 17818 4580 17824
rect 4528 17740 4580 17746
rect 4528 17682 4580 17688
rect 4160 17672 4212 17678
rect 4160 17614 4212 17620
rect 3756 17436 4064 17445
rect 3756 17434 3762 17436
rect 3818 17434 3842 17436
rect 3898 17434 3922 17436
rect 3978 17434 4002 17436
rect 4058 17434 4064 17436
rect 3818 17382 3820 17434
rect 4000 17382 4002 17434
rect 3756 17380 3762 17382
rect 3818 17380 3842 17382
rect 3898 17380 3922 17382
rect 3978 17380 4002 17382
rect 4058 17380 4064 17382
rect 3756 17371 4064 17380
rect 4172 16998 4200 17614
rect 4344 17536 4396 17542
rect 4344 17478 4396 17484
rect 4356 17134 4384 17478
rect 4344 17128 4396 17134
rect 4344 17070 4396 17076
rect 4160 16992 4212 16998
rect 4160 16934 4212 16940
rect 4172 16454 4200 16934
rect 4344 16788 4396 16794
rect 4344 16730 4396 16736
rect 4160 16448 4212 16454
rect 4160 16390 4212 16396
rect 3756 16348 4064 16357
rect 3756 16346 3762 16348
rect 3818 16346 3842 16348
rect 3898 16346 3922 16348
rect 3978 16346 4002 16348
rect 4058 16346 4064 16348
rect 3818 16294 3820 16346
rect 4000 16294 4002 16346
rect 3756 16292 3762 16294
rect 3818 16292 3842 16294
rect 3898 16292 3922 16294
rect 3978 16292 4002 16294
rect 4058 16292 4064 16294
rect 3756 16283 4064 16292
rect 4356 16250 4384 16730
rect 4540 16454 4568 17682
rect 4528 16448 4580 16454
rect 4528 16390 4580 16396
rect 4344 16244 4396 16250
rect 4344 16186 4396 16192
rect 4632 16046 4660 19110
rect 4988 18624 5040 18630
rect 4988 18566 5040 18572
rect 5000 18222 5028 18566
rect 5092 18426 5120 19858
rect 5736 19854 5764 20334
rect 5724 19848 5776 19854
rect 5724 19790 5776 19796
rect 5632 19712 5684 19718
rect 5632 19654 5684 19660
rect 5644 19378 5672 19654
rect 5632 19372 5684 19378
rect 5632 19314 5684 19320
rect 5632 19236 5684 19242
rect 5460 19196 5632 19224
rect 5080 18420 5132 18426
rect 5080 18362 5132 18368
rect 5264 18284 5316 18290
rect 5264 18226 5316 18232
rect 4988 18216 5040 18222
rect 4988 18158 5040 18164
rect 4804 18148 4856 18154
rect 4804 18090 4856 18096
rect 4816 17882 4844 18090
rect 4804 17876 4856 17882
rect 4804 17818 4856 17824
rect 5172 17740 5224 17746
rect 5172 17682 5224 17688
rect 5184 17338 5212 17682
rect 5276 17338 5304 18226
rect 5460 18086 5488 19196
rect 5632 19178 5684 19184
rect 5736 18834 5764 19790
rect 5828 19446 5856 21100
rect 5816 19440 5868 19446
rect 5816 19382 5868 19388
rect 5816 19304 5868 19310
rect 5816 19246 5868 19252
rect 5828 18970 5856 19246
rect 5920 19174 5948 21270
rect 5908 19168 5960 19174
rect 5908 19110 5960 19116
rect 5816 18964 5868 18970
rect 6012 18952 6040 29650
rect 6104 29102 6132 29990
rect 6288 29714 6316 30534
rect 6380 30054 6408 30602
rect 6840 30274 6868 30654
rect 6920 30592 6972 30598
rect 6920 30534 6972 30540
rect 6460 30252 6512 30258
rect 6460 30194 6512 30200
rect 6656 30246 6868 30274
rect 6368 30048 6420 30054
rect 6368 29990 6420 29996
rect 6276 29708 6328 29714
rect 6276 29650 6328 29656
rect 6380 29238 6408 29990
rect 6368 29232 6420 29238
rect 6368 29174 6420 29180
rect 6092 29096 6144 29102
rect 6092 29038 6144 29044
rect 6472 28558 6500 30194
rect 6552 29708 6604 29714
rect 6552 29650 6604 29656
rect 6460 28552 6512 28558
rect 6460 28494 6512 28500
rect 6092 28212 6144 28218
rect 6092 28154 6144 28160
rect 6104 27674 6132 28154
rect 6184 27940 6236 27946
rect 6184 27882 6236 27888
rect 6092 27668 6144 27674
rect 6092 27610 6144 27616
rect 6104 26926 6132 27610
rect 6196 27538 6224 27882
rect 6184 27532 6236 27538
rect 6236 27492 6316 27520
rect 6184 27474 6236 27480
rect 6184 27328 6236 27334
rect 6184 27270 6236 27276
rect 6092 26920 6144 26926
rect 6092 26862 6144 26868
rect 6092 26784 6144 26790
rect 6092 26726 6144 26732
rect 6104 26450 6132 26726
rect 6196 26586 6224 27270
rect 6288 26790 6316 27492
rect 6368 26988 6420 26994
rect 6368 26930 6420 26936
rect 6276 26784 6328 26790
rect 6276 26726 6328 26732
rect 6184 26580 6236 26586
rect 6184 26522 6236 26528
rect 6196 26450 6224 26522
rect 6092 26444 6144 26450
rect 6092 26386 6144 26392
rect 6184 26444 6236 26450
rect 6380 26432 6408 26930
rect 6472 26450 6500 28494
rect 6184 26386 6236 26392
rect 6288 26404 6408 26432
rect 6460 26444 6512 26450
rect 6288 25838 6316 26404
rect 6460 26386 6512 26392
rect 6368 26308 6420 26314
rect 6368 26250 6420 26256
rect 6276 25832 6328 25838
rect 6276 25774 6328 25780
rect 6184 24676 6236 24682
rect 6184 24618 6236 24624
rect 6196 24410 6224 24618
rect 6276 24608 6328 24614
rect 6276 24550 6328 24556
rect 6288 24410 6316 24550
rect 6184 24404 6236 24410
rect 6184 24346 6236 24352
rect 6276 24404 6328 24410
rect 6276 24346 6328 24352
rect 6092 23248 6144 23254
rect 6092 23190 6144 23196
rect 6182 23216 6238 23225
rect 6104 21486 6132 23190
rect 6182 23151 6184 23160
rect 6236 23151 6238 23160
rect 6184 23122 6236 23128
rect 6276 23112 6328 23118
rect 6276 23054 6328 23060
rect 6184 22024 6236 22030
rect 6184 21966 6236 21972
rect 6092 21480 6144 21486
rect 6092 21422 6144 21428
rect 6196 21010 6224 21966
rect 6288 21486 6316 23054
rect 6380 22574 6408 26250
rect 6460 23588 6512 23594
rect 6460 23530 6512 23536
rect 6472 23322 6500 23530
rect 6460 23316 6512 23322
rect 6460 23258 6512 23264
rect 6368 22568 6420 22574
rect 6368 22510 6420 22516
rect 6564 22094 6592 29650
rect 6656 29034 6684 30246
rect 6932 30190 6960 30534
rect 8036 30394 8064 30670
rect 8760 30660 8812 30666
rect 8760 30602 8812 30608
rect 8024 30388 8076 30394
rect 8024 30330 8076 30336
rect 6920 30184 6972 30190
rect 6920 30126 6972 30132
rect 7114 29948 7422 29957
rect 7114 29946 7120 29948
rect 7176 29946 7200 29948
rect 7256 29946 7280 29948
rect 7336 29946 7360 29948
rect 7416 29946 7422 29948
rect 7176 29894 7178 29946
rect 7358 29894 7360 29946
rect 7114 29892 7120 29894
rect 7176 29892 7200 29894
rect 7256 29892 7280 29894
rect 7336 29892 7360 29894
rect 7416 29892 7422 29894
rect 7114 29883 7422 29892
rect 7012 29708 7064 29714
rect 7012 29650 7064 29656
rect 6828 29640 6880 29646
rect 6828 29582 6880 29588
rect 6644 29028 6696 29034
rect 6644 28970 6696 28976
rect 6656 28422 6684 28970
rect 6840 28762 6868 29582
rect 7024 29306 7052 29650
rect 7012 29300 7064 29306
rect 7012 29242 7064 29248
rect 7114 28860 7422 28869
rect 7114 28858 7120 28860
rect 7176 28858 7200 28860
rect 7256 28858 7280 28860
rect 7336 28858 7360 28860
rect 7416 28858 7422 28860
rect 7176 28806 7178 28858
rect 7358 28806 7360 28858
rect 7114 28804 7120 28806
rect 7176 28804 7200 28806
rect 7256 28804 7280 28806
rect 7336 28804 7360 28806
rect 7416 28804 7422 28806
rect 7114 28795 7422 28804
rect 6828 28756 6880 28762
rect 6828 28698 6880 28704
rect 6736 28620 6788 28626
rect 6736 28562 6788 28568
rect 6644 28416 6696 28422
rect 6644 28358 6696 28364
rect 6656 27946 6684 28358
rect 6748 28218 6776 28562
rect 6736 28212 6788 28218
rect 6736 28154 6788 28160
rect 6840 28014 6868 28698
rect 7840 28620 7892 28626
rect 7840 28562 7892 28568
rect 7472 28484 7524 28490
rect 7472 28426 7524 28432
rect 7484 28014 7512 28426
rect 7852 28422 7880 28562
rect 8036 28558 8064 30330
rect 8484 30252 8536 30258
rect 8484 30194 8536 30200
rect 8300 30184 8352 30190
rect 8300 30126 8352 30132
rect 8312 29034 8340 30126
rect 8392 29504 8444 29510
rect 8496 29492 8524 30194
rect 8576 30048 8628 30054
rect 8576 29990 8628 29996
rect 8668 30048 8720 30054
rect 8668 29990 8720 29996
rect 8444 29464 8524 29492
rect 8392 29446 8444 29452
rect 8300 29028 8352 29034
rect 8300 28970 8352 28976
rect 8116 28688 8168 28694
rect 8116 28630 8168 28636
rect 8024 28552 8076 28558
rect 8024 28494 8076 28500
rect 7840 28416 7892 28422
rect 7840 28358 7892 28364
rect 7852 28014 7880 28358
rect 6828 28008 6880 28014
rect 6828 27950 6880 27956
rect 7472 28008 7524 28014
rect 7472 27950 7524 27956
rect 7840 28008 7892 28014
rect 7840 27950 7892 27956
rect 6644 27940 6696 27946
rect 6644 27882 6696 27888
rect 6656 23361 6684 27882
rect 6736 27872 6788 27878
rect 6736 27814 6788 27820
rect 6748 26353 6776 27814
rect 6840 27606 6868 27950
rect 8036 27946 8064 28494
rect 8128 28218 8156 28630
rect 8312 28490 8340 28970
rect 8300 28484 8352 28490
rect 8300 28426 8352 28432
rect 8404 28370 8432 29446
rect 8588 29306 8616 29990
rect 8680 29714 8708 29990
rect 8668 29708 8720 29714
rect 8668 29650 8720 29656
rect 8576 29300 8628 29306
rect 8576 29242 8628 29248
rect 8772 28966 8800 30602
rect 9680 30592 9732 30598
rect 9680 30534 9732 30540
rect 9692 30274 9720 30534
rect 9416 30246 9720 30274
rect 9416 30190 9444 30246
rect 8852 30184 8904 30190
rect 8852 30126 8904 30132
rect 9128 30184 9180 30190
rect 9128 30126 9180 30132
rect 9404 30184 9456 30190
rect 9404 30126 9456 30132
rect 8864 29238 8892 30126
rect 9140 29850 9168 30126
rect 9312 30048 9364 30054
rect 9312 29990 9364 29996
rect 9128 29844 9180 29850
rect 9128 29786 9180 29792
rect 8944 29776 8996 29782
rect 8944 29718 8996 29724
rect 8852 29232 8904 29238
rect 8852 29174 8904 29180
rect 8576 28960 8628 28966
rect 8576 28902 8628 28908
rect 8760 28960 8812 28966
rect 8760 28902 8812 28908
rect 8588 28694 8616 28902
rect 8576 28688 8628 28694
rect 8576 28630 8628 28636
rect 8484 28484 8536 28490
rect 8484 28426 8536 28432
rect 8496 28370 8524 28426
rect 8404 28342 8524 28370
rect 8116 28212 8168 28218
rect 8116 28154 8168 28160
rect 8404 28014 8432 28342
rect 8392 28008 8444 28014
rect 8392 27950 8444 27956
rect 8024 27940 8076 27946
rect 8024 27882 8076 27888
rect 7114 27772 7422 27781
rect 7114 27770 7120 27772
rect 7176 27770 7200 27772
rect 7256 27770 7280 27772
rect 7336 27770 7360 27772
rect 7416 27770 7422 27772
rect 7176 27718 7178 27770
rect 7358 27718 7360 27770
rect 7114 27716 7120 27718
rect 7176 27716 7200 27718
rect 7256 27716 7280 27718
rect 7336 27716 7360 27718
rect 7416 27716 7422 27718
rect 7114 27707 7422 27716
rect 8036 27674 8064 27882
rect 6920 27668 6972 27674
rect 6920 27610 6972 27616
rect 8024 27668 8076 27674
rect 8024 27610 8076 27616
rect 6828 27600 6880 27606
rect 6828 27542 6880 27548
rect 6932 26994 6960 27610
rect 7012 27532 7064 27538
rect 7012 27474 7064 27480
rect 6920 26988 6972 26994
rect 6920 26930 6972 26936
rect 6920 26852 6972 26858
rect 6920 26794 6972 26800
rect 6828 26784 6880 26790
rect 6828 26726 6880 26732
rect 6734 26344 6790 26353
rect 6734 26279 6790 26288
rect 6840 26246 6868 26726
rect 6828 26240 6880 26246
rect 6828 26182 6880 26188
rect 6932 25906 6960 26794
rect 7024 26042 7052 27474
rect 8404 27470 8432 27950
rect 8484 27940 8536 27946
rect 8484 27882 8536 27888
rect 8496 27470 8524 27882
rect 8588 27878 8616 28630
rect 8956 27946 8984 29718
rect 9324 29102 9352 29990
rect 10152 29850 10180 30806
rect 10244 30802 10272 31600
rect 11716 30802 11744 31600
rect 10232 30796 10284 30802
rect 10232 30738 10284 30744
rect 11704 30796 11756 30802
rect 11704 30738 11756 30744
rect 12072 30796 12124 30802
rect 12072 30738 12124 30744
rect 11244 30660 11296 30666
rect 11244 30602 11296 30608
rect 10324 30592 10376 30598
rect 10324 30534 10376 30540
rect 11060 30592 11112 30598
rect 11060 30534 11112 30540
rect 10336 29850 10364 30534
rect 10472 30492 10780 30501
rect 10472 30490 10478 30492
rect 10534 30490 10558 30492
rect 10614 30490 10638 30492
rect 10694 30490 10718 30492
rect 10774 30490 10780 30492
rect 10534 30438 10536 30490
rect 10716 30438 10718 30490
rect 10472 30436 10478 30438
rect 10534 30436 10558 30438
rect 10614 30436 10638 30438
rect 10694 30436 10718 30438
rect 10774 30436 10780 30438
rect 10472 30427 10780 30436
rect 11072 30190 11100 30534
rect 11256 30190 11284 30602
rect 11704 30592 11756 30598
rect 11704 30534 11756 30540
rect 11336 30252 11388 30258
rect 11336 30194 11388 30200
rect 11060 30184 11112 30190
rect 11060 30126 11112 30132
rect 11244 30184 11296 30190
rect 11244 30126 11296 30132
rect 10600 30048 10652 30054
rect 10600 29990 10652 29996
rect 10876 30048 10928 30054
rect 10876 29990 10928 29996
rect 10140 29844 10192 29850
rect 10140 29786 10192 29792
rect 10324 29844 10376 29850
rect 10324 29786 10376 29792
rect 10048 29640 10100 29646
rect 10048 29582 10100 29588
rect 10060 29238 10088 29582
rect 10048 29232 10100 29238
rect 10048 29174 10100 29180
rect 9312 29096 9364 29102
rect 9312 29038 9364 29044
rect 9956 29096 10008 29102
rect 9956 29038 10008 29044
rect 9324 28506 9352 29038
rect 9404 28960 9456 28966
rect 9404 28902 9456 28908
rect 9416 28694 9444 28902
rect 9404 28688 9456 28694
rect 9404 28630 9456 28636
rect 9772 28620 9824 28626
rect 9772 28562 9824 28568
rect 9324 28478 9444 28506
rect 8944 27940 8996 27946
rect 8944 27882 8996 27888
rect 8576 27872 8628 27878
rect 8576 27814 8628 27820
rect 8392 27464 8444 27470
rect 8392 27406 8444 27412
rect 8484 27464 8536 27470
rect 8484 27406 8536 27412
rect 8116 26920 8168 26926
rect 8116 26862 8168 26868
rect 7472 26784 7524 26790
rect 7472 26726 7524 26732
rect 7114 26684 7422 26693
rect 7114 26682 7120 26684
rect 7176 26682 7200 26684
rect 7256 26682 7280 26684
rect 7336 26682 7360 26684
rect 7416 26682 7422 26684
rect 7176 26630 7178 26682
rect 7358 26630 7360 26682
rect 7114 26628 7120 26630
rect 7176 26628 7200 26630
rect 7256 26628 7280 26630
rect 7336 26628 7360 26630
rect 7416 26628 7422 26630
rect 7114 26619 7422 26628
rect 7012 26036 7064 26042
rect 7012 25978 7064 25984
rect 6920 25900 6972 25906
rect 6920 25842 6972 25848
rect 6932 25430 6960 25842
rect 7484 25838 7512 26726
rect 8128 26586 8156 26862
rect 8116 26580 8168 26586
rect 8116 26522 8168 26528
rect 8300 26444 8352 26450
rect 8300 26386 8352 26392
rect 8312 25838 8340 26386
rect 8404 25838 8432 27406
rect 8496 26926 8524 27406
rect 9312 27396 9364 27402
rect 9312 27338 9364 27344
rect 9036 27328 9088 27334
rect 9036 27270 9088 27276
rect 9128 27328 9180 27334
rect 9128 27270 9180 27276
rect 8484 26920 8536 26926
rect 9048 26908 9076 27270
rect 9140 27062 9168 27270
rect 9324 27130 9352 27338
rect 9312 27124 9364 27130
rect 9312 27066 9364 27072
rect 9128 27056 9180 27062
rect 9128 26998 9180 27004
rect 9128 26920 9180 26926
rect 9048 26880 9128 26908
rect 8484 26862 8536 26868
rect 9128 26862 9180 26868
rect 9416 26858 9444 28478
rect 9784 27470 9812 28562
rect 9968 28218 9996 29038
rect 9956 28212 10008 28218
rect 9956 28154 10008 28160
rect 10060 28014 10088 29174
rect 10336 29170 10364 29786
rect 10612 29714 10640 29990
rect 10600 29708 10652 29714
rect 10600 29650 10652 29656
rect 10472 29404 10780 29413
rect 10472 29402 10478 29404
rect 10534 29402 10558 29404
rect 10614 29402 10638 29404
rect 10694 29402 10718 29404
rect 10774 29402 10780 29404
rect 10534 29350 10536 29402
rect 10716 29350 10718 29402
rect 10472 29348 10478 29350
rect 10534 29348 10558 29350
rect 10614 29348 10638 29350
rect 10694 29348 10718 29350
rect 10774 29348 10780 29350
rect 10472 29339 10780 29348
rect 10324 29164 10376 29170
rect 10324 29106 10376 29112
rect 10232 29096 10284 29102
rect 10232 29038 10284 29044
rect 10140 28960 10192 28966
rect 10140 28902 10192 28908
rect 10152 28218 10180 28902
rect 10244 28558 10272 29038
rect 10336 28762 10364 29106
rect 10324 28756 10376 28762
rect 10324 28698 10376 28704
rect 10232 28552 10284 28558
rect 10232 28494 10284 28500
rect 10244 28422 10272 28494
rect 10324 28484 10376 28490
rect 10324 28426 10376 28432
rect 10232 28416 10284 28422
rect 10232 28358 10284 28364
rect 10140 28212 10192 28218
rect 10140 28154 10192 28160
rect 10336 28082 10364 28426
rect 10472 28316 10780 28325
rect 10472 28314 10478 28316
rect 10534 28314 10558 28316
rect 10614 28314 10638 28316
rect 10694 28314 10718 28316
rect 10774 28314 10780 28316
rect 10534 28262 10536 28314
rect 10716 28262 10718 28314
rect 10472 28260 10478 28262
rect 10534 28260 10558 28262
rect 10614 28260 10638 28262
rect 10694 28260 10718 28262
rect 10774 28260 10780 28262
rect 10472 28251 10780 28260
rect 10324 28076 10376 28082
rect 10324 28018 10376 28024
rect 10888 28014 10916 29990
rect 11072 29850 11100 30126
rect 11060 29844 11112 29850
rect 11060 29786 11112 29792
rect 11256 29782 11284 30126
rect 11244 29776 11296 29782
rect 11244 29718 11296 29724
rect 11348 29050 11376 30194
rect 11428 30116 11480 30122
rect 11428 30058 11480 30064
rect 11440 29306 11468 30058
rect 11428 29300 11480 29306
rect 11428 29242 11480 29248
rect 11716 29102 11744 30534
rect 12084 30394 12112 30738
rect 12716 30728 12768 30734
rect 12716 30670 12768 30676
rect 12728 30394 12756 30670
rect 12072 30388 12124 30394
rect 12072 30330 12124 30336
rect 12716 30388 12768 30394
rect 12716 30330 12768 30336
rect 12728 29850 12756 30330
rect 13188 30190 13216 31600
rect 13830 31036 14138 31045
rect 13830 31034 13836 31036
rect 13892 31034 13916 31036
rect 13972 31034 13996 31036
rect 14052 31034 14076 31036
rect 14132 31034 14138 31036
rect 13892 30982 13894 31034
rect 14074 30982 14076 31034
rect 13830 30980 13836 30982
rect 13892 30980 13916 30982
rect 13972 30980 13996 30982
rect 14052 30980 14076 30982
rect 14132 30980 14138 30982
rect 13830 30971 14138 30980
rect 14660 30802 14688 31600
rect 16132 30870 16160 31600
rect 17604 31498 17632 31600
rect 17696 31498 17724 31606
rect 17604 31470 17724 31498
rect 16672 31136 16724 31142
rect 16672 31078 16724 31084
rect 16120 30864 16172 30870
rect 16120 30806 16172 30812
rect 16684 30802 16712 31078
rect 17972 30870 18000 31606
rect 19062 31600 19118 32000
rect 19168 31606 19380 31634
rect 19076 31498 19104 31600
rect 19168 31498 19196 31606
rect 19076 31470 19196 31498
rect 19352 30870 19380 31606
rect 20534 31600 20590 32000
rect 20640 31606 20944 31634
rect 20548 31498 20576 31600
rect 20640 31498 20668 31606
rect 20548 31470 20668 31498
rect 19432 31136 19484 31142
rect 19432 31078 19484 31084
rect 19444 30938 19472 31078
rect 20546 31036 20854 31045
rect 20546 31034 20552 31036
rect 20608 31034 20632 31036
rect 20688 31034 20712 31036
rect 20768 31034 20792 31036
rect 20848 31034 20854 31036
rect 20608 30982 20610 31034
rect 20790 30982 20792 31034
rect 20546 30980 20552 30982
rect 20608 30980 20632 30982
rect 20688 30980 20712 30982
rect 20768 30980 20792 30982
rect 20848 30980 20854 30982
rect 20546 30971 20854 30980
rect 19432 30932 19484 30938
rect 19432 30874 19484 30880
rect 20916 30870 20944 31606
rect 22006 31600 22062 32000
rect 23478 31600 23534 32000
rect 24950 31600 25006 32000
rect 26422 31600 26478 32000
rect 22020 30954 22048 31600
rect 22020 30926 22140 30954
rect 22112 30870 22140 30926
rect 17960 30864 18012 30870
rect 17682 30832 17738 30841
rect 14188 30796 14240 30802
rect 14188 30738 14240 30744
rect 14648 30796 14700 30802
rect 14648 30738 14700 30744
rect 16672 30796 16724 30802
rect 19156 30864 19208 30870
rect 17960 30806 18012 30812
rect 19062 30832 19118 30841
rect 17682 30767 17684 30776
rect 16672 30738 16724 30744
rect 17736 30767 17738 30776
rect 17776 30796 17828 30802
rect 17684 30738 17736 30744
rect 17776 30738 17828 30744
rect 18052 30796 18104 30802
rect 18052 30738 18104 30744
rect 18788 30796 18840 30802
rect 19156 30806 19208 30812
rect 19340 30864 19392 30870
rect 19340 30806 19392 30812
rect 20904 30864 20956 30870
rect 20904 30806 20956 30812
rect 22100 30864 22152 30870
rect 22100 30806 22152 30812
rect 18788 30738 18840 30744
rect 18984 30776 19062 30784
rect 18984 30756 19064 30776
rect 13636 30592 13688 30598
rect 13636 30534 13688 30540
rect 14004 30592 14056 30598
rect 14004 30534 14056 30540
rect 13176 30184 13228 30190
rect 13176 30126 13228 30132
rect 13176 30048 13228 30054
rect 13176 29990 13228 29996
rect 13544 30048 13596 30054
rect 13544 29990 13596 29996
rect 12716 29844 12768 29850
rect 12716 29786 12768 29792
rect 12532 29640 12584 29646
rect 12532 29582 12584 29588
rect 12624 29640 12676 29646
rect 12624 29582 12676 29588
rect 12256 29504 12308 29510
rect 12256 29446 12308 29452
rect 11704 29096 11756 29102
rect 10968 29028 11020 29034
rect 10968 28970 11020 28976
rect 11152 29028 11204 29034
rect 11348 29022 11468 29050
rect 11704 29038 11756 29044
rect 11152 28970 11204 28976
rect 10980 28490 11008 28970
rect 10968 28484 11020 28490
rect 10968 28426 11020 28432
rect 10980 28150 11008 28426
rect 11060 28416 11112 28422
rect 11060 28358 11112 28364
rect 10968 28144 11020 28150
rect 10968 28086 11020 28092
rect 10048 28008 10100 28014
rect 10048 27950 10100 27956
rect 10876 28008 10928 28014
rect 10876 27950 10928 27956
rect 10324 27940 10376 27946
rect 10324 27882 10376 27888
rect 9772 27464 9824 27470
rect 9772 27406 9824 27412
rect 9864 27328 9916 27334
rect 9864 27270 9916 27276
rect 9772 26920 9824 26926
rect 9772 26862 9824 26868
rect 9404 26852 9456 26858
rect 9404 26794 9456 26800
rect 9220 26444 9272 26450
rect 9220 26386 9272 26392
rect 8576 26240 8628 26246
rect 8576 26182 8628 26188
rect 8668 26240 8720 26246
rect 8668 26182 8720 26188
rect 8588 26042 8616 26182
rect 8576 26036 8628 26042
rect 8576 25978 8628 25984
rect 8680 25838 8708 26182
rect 7012 25832 7064 25838
rect 7012 25774 7064 25780
rect 7472 25832 7524 25838
rect 7472 25774 7524 25780
rect 8300 25832 8352 25838
rect 8300 25774 8352 25780
rect 8392 25832 8444 25838
rect 8392 25774 8444 25780
rect 8668 25832 8720 25838
rect 8668 25774 8720 25780
rect 6920 25424 6972 25430
rect 6920 25366 6972 25372
rect 6932 25294 6960 25366
rect 7024 25362 7052 25774
rect 7840 25764 7892 25770
rect 7840 25706 7892 25712
rect 7114 25596 7422 25605
rect 7114 25594 7120 25596
rect 7176 25594 7200 25596
rect 7256 25594 7280 25596
rect 7336 25594 7360 25596
rect 7416 25594 7422 25596
rect 7176 25542 7178 25594
rect 7358 25542 7360 25594
rect 7114 25540 7120 25542
rect 7176 25540 7200 25542
rect 7256 25540 7280 25542
rect 7336 25540 7360 25542
rect 7416 25540 7422 25542
rect 7114 25531 7422 25540
rect 7852 25498 7880 25706
rect 7932 25696 7984 25702
rect 7932 25638 7984 25644
rect 7840 25492 7892 25498
rect 7840 25434 7892 25440
rect 7012 25356 7064 25362
rect 7012 25298 7064 25304
rect 7656 25356 7708 25362
rect 7656 25298 7708 25304
rect 6920 25288 6972 25294
rect 6920 25230 6972 25236
rect 6736 24608 6788 24614
rect 6736 24550 6788 24556
rect 6748 24274 6776 24550
rect 6932 24342 6960 25230
rect 6920 24336 6972 24342
rect 6920 24278 6972 24284
rect 6736 24268 6788 24274
rect 6736 24210 6788 24216
rect 6828 24268 6880 24274
rect 6828 24210 6880 24216
rect 6840 23866 6868 24210
rect 6828 23860 6880 23866
rect 6828 23802 6880 23808
rect 6642 23352 6698 23361
rect 6642 23287 6698 23296
rect 6932 23254 6960 24278
rect 7024 24138 7052 25298
rect 7564 25152 7616 25158
rect 7564 25094 7616 25100
rect 7472 24744 7524 24750
rect 7472 24686 7524 24692
rect 7114 24508 7422 24517
rect 7114 24506 7120 24508
rect 7176 24506 7200 24508
rect 7256 24506 7280 24508
rect 7336 24506 7360 24508
rect 7416 24506 7422 24508
rect 7176 24454 7178 24506
rect 7358 24454 7360 24506
rect 7114 24452 7120 24454
rect 7176 24452 7200 24454
rect 7256 24452 7280 24454
rect 7336 24452 7360 24454
rect 7416 24452 7422 24454
rect 7114 24443 7422 24452
rect 7196 24268 7248 24274
rect 7196 24210 7248 24216
rect 7208 24138 7236 24210
rect 7484 24206 7512 24686
rect 7576 24342 7604 25094
rect 7564 24336 7616 24342
rect 7564 24278 7616 24284
rect 7380 24200 7432 24206
rect 7380 24142 7432 24148
rect 7472 24200 7524 24206
rect 7472 24142 7524 24148
rect 7012 24132 7064 24138
rect 7012 24074 7064 24080
rect 7196 24132 7248 24138
rect 7196 24074 7248 24080
rect 7208 23798 7236 24074
rect 7196 23792 7248 23798
rect 7196 23734 7248 23740
rect 7392 23526 7420 24142
rect 7564 23792 7616 23798
rect 7564 23734 7616 23740
rect 7012 23520 7064 23526
rect 7012 23462 7064 23468
rect 7380 23520 7432 23526
rect 7380 23462 7432 23468
rect 6920 23248 6972 23254
rect 6920 23190 6972 23196
rect 7024 23186 7052 23462
rect 7114 23420 7422 23429
rect 7114 23418 7120 23420
rect 7176 23418 7200 23420
rect 7256 23418 7280 23420
rect 7336 23418 7360 23420
rect 7416 23418 7422 23420
rect 7176 23366 7178 23418
rect 7358 23366 7360 23418
rect 7114 23364 7120 23366
rect 7176 23364 7200 23366
rect 7256 23364 7280 23366
rect 7336 23364 7360 23366
rect 7416 23364 7422 23366
rect 7114 23355 7422 23364
rect 7576 23322 7604 23734
rect 7564 23316 7616 23322
rect 7564 23258 7616 23264
rect 7576 23186 7604 23258
rect 6736 23180 6788 23186
rect 6656 23140 6736 23168
rect 6656 23050 6684 23140
rect 6736 23122 6788 23128
rect 7012 23180 7064 23186
rect 7012 23122 7064 23128
rect 7104 23180 7156 23186
rect 7104 23122 7156 23128
rect 7564 23180 7616 23186
rect 7564 23122 7616 23128
rect 6644 23044 6696 23050
rect 6644 22986 6696 22992
rect 6380 22066 6592 22094
rect 6276 21480 6328 21486
rect 6276 21422 6328 21428
rect 6184 21004 6236 21010
rect 6184 20946 6236 20952
rect 6380 19122 6408 22066
rect 6460 21888 6512 21894
rect 6460 21830 6512 21836
rect 6472 21486 6500 21830
rect 6460 21480 6512 21486
rect 6460 21422 6512 21428
rect 5816 18906 5868 18912
rect 5920 18924 6040 18952
rect 6196 19094 6408 19122
rect 6460 19168 6512 19174
rect 6460 19110 6512 19116
rect 5724 18828 5776 18834
rect 5724 18770 5776 18776
rect 5632 18284 5684 18290
rect 5632 18226 5684 18232
rect 5540 18216 5592 18222
rect 5540 18158 5592 18164
rect 5448 18080 5500 18086
rect 5448 18022 5500 18028
rect 5172 17332 5224 17338
rect 5172 17274 5224 17280
rect 5264 17332 5316 17338
rect 5264 17274 5316 17280
rect 4896 17128 4948 17134
rect 4896 17070 4948 17076
rect 4988 17128 5040 17134
rect 4988 17070 5040 17076
rect 4908 16522 4936 17070
rect 5000 16794 5028 17070
rect 4988 16788 5040 16794
rect 4988 16730 5040 16736
rect 5276 16658 5304 17274
rect 5460 17270 5488 18022
rect 5552 17814 5580 18158
rect 5540 17808 5592 17814
rect 5540 17750 5592 17756
rect 5644 17626 5672 18226
rect 5552 17598 5672 17626
rect 5552 17542 5580 17598
rect 5540 17536 5592 17542
rect 5540 17478 5592 17484
rect 5632 17536 5684 17542
rect 5632 17478 5684 17484
rect 5448 17264 5500 17270
rect 5448 17206 5500 17212
rect 5356 17196 5408 17202
rect 5356 17138 5408 17144
rect 5368 16998 5396 17138
rect 5644 17134 5672 17478
rect 5632 17128 5684 17134
rect 5632 17070 5684 17076
rect 5356 16992 5408 16998
rect 5356 16934 5408 16940
rect 5448 16992 5500 16998
rect 5448 16934 5500 16940
rect 5460 16794 5488 16934
rect 5448 16788 5500 16794
rect 5448 16730 5500 16736
rect 5264 16652 5316 16658
rect 5264 16594 5316 16600
rect 4896 16516 4948 16522
rect 4896 16458 4948 16464
rect 5816 16108 5868 16114
rect 5816 16050 5868 16056
rect 4620 16040 4672 16046
rect 4804 16040 4856 16046
rect 4672 16000 4752 16028
rect 4620 15982 4672 15988
rect 4160 15972 4212 15978
rect 4160 15914 4212 15920
rect 3608 15632 3660 15638
rect 3608 15574 3660 15580
rect 3620 15162 3648 15574
rect 3756 15260 4064 15269
rect 3756 15258 3762 15260
rect 3818 15258 3842 15260
rect 3898 15258 3922 15260
rect 3978 15258 4002 15260
rect 4058 15258 4064 15260
rect 3818 15206 3820 15258
rect 4000 15206 4002 15258
rect 3756 15204 3762 15206
rect 3818 15204 3842 15206
rect 3898 15204 3922 15206
rect 3978 15204 4002 15206
rect 4058 15204 4064 15206
rect 3756 15195 4064 15204
rect 3608 15156 3660 15162
rect 3608 15098 3660 15104
rect 4172 15026 4200 15914
rect 4620 15904 4672 15910
rect 4620 15846 4672 15852
rect 4528 15360 4580 15366
rect 4528 15302 4580 15308
rect 4160 15020 4212 15026
rect 4160 14962 4212 14968
rect 4540 14958 4568 15302
rect 4632 15026 4660 15846
rect 4724 15026 4752 16000
rect 4804 15982 4856 15988
rect 4816 15366 4844 15982
rect 5080 15564 5132 15570
rect 5080 15506 5132 15512
rect 4804 15360 4856 15366
rect 4804 15302 4856 15308
rect 4620 15020 4672 15026
rect 4620 14962 4672 14968
rect 4712 15020 4764 15026
rect 4712 14962 4764 14968
rect 4528 14952 4580 14958
rect 4528 14894 4580 14900
rect 4540 14414 4568 14894
rect 4816 14482 4844 15302
rect 5092 14550 5120 15506
rect 5828 15366 5856 16050
rect 5172 15360 5224 15366
rect 5172 15302 5224 15308
rect 5816 15360 5868 15366
rect 5816 15302 5868 15308
rect 5184 14890 5212 15302
rect 5172 14884 5224 14890
rect 5172 14826 5224 14832
rect 5080 14544 5132 14550
rect 5828 14498 5856 15302
rect 5080 14486 5132 14492
rect 5460 14482 5856 14498
rect 4804 14476 4856 14482
rect 4804 14418 4856 14424
rect 5448 14476 5856 14482
rect 5500 14470 5856 14476
rect 5448 14418 5500 14424
rect 4528 14408 4580 14414
rect 4528 14350 4580 14356
rect 3756 14172 4064 14181
rect 3756 14170 3762 14172
rect 3818 14170 3842 14172
rect 3898 14170 3922 14172
rect 3978 14170 4002 14172
rect 4058 14170 4064 14172
rect 3818 14118 3820 14170
rect 4000 14118 4002 14170
rect 3756 14116 3762 14118
rect 3818 14116 3842 14118
rect 3898 14116 3922 14118
rect 3978 14116 4002 14118
rect 4058 14116 4064 14118
rect 3756 14107 4064 14116
rect 4540 13870 4568 14350
rect 4528 13864 4580 13870
rect 4528 13806 4580 13812
rect 5172 13864 5224 13870
rect 5172 13806 5224 13812
rect 5448 13864 5500 13870
rect 5448 13806 5500 13812
rect 4160 13796 4212 13802
rect 4160 13738 4212 13744
rect 3884 13728 3936 13734
rect 3884 13670 3936 13676
rect 3896 13394 3924 13670
rect 4172 13530 4200 13738
rect 4160 13524 4212 13530
rect 4160 13466 4212 13472
rect 3884 13388 3936 13394
rect 3884 13330 3936 13336
rect 4540 13190 4568 13806
rect 4712 13796 4764 13802
rect 4712 13738 4764 13744
rect 4620 13728 4672 13734
rect 4620 13670 4672 13676
rect 4528 13184 4580 13190
rect 4528 13126 4580 13132
rect 3756 13084 4064 13093
rect 3756 13082 3762 13084
rect 3818 13082 3842 13084
rect 3898 13082 3922 13084
rect 3978 13082 4002 13084
rect 4058 13082 4064 13084
rect 3818 13030 3820 13082
rect 4000 13030 4002 13082
rect 3756 13028 3762 13030
rect 3818 13028 3842 13030
rect 3898 13028 3922 13030
rect 3978 13028 4002 13030
rect 4058 13028 4064 13030
rect 3756 13019 4064 13028
rect 4528 12980 4580 12986
rect 4528 12922 4580 12928
rect 3700 12912 3752 12918
rect 3700 12854 3752 12860
rect 3608 12708 3660 12714
rect 3608 12650 3660 12656
rect 3620 12306 3648 12650
rect 3712 12442 3740 12854
rect 4540 12850 4568 12922
rect 4528 12844 4580 12850
rect 4528 12786 4580 12792
rect 4344 12776 4396 12782
rect 4344 12718 4396 12724
rect 4252 12640 4304 12646
rect 4252 12582 4304 12588
rect 3700 12436 3752 12442
rect 3700 12378 3752 12384
rect 3608 12300 3660 12306
rect 3608 12242 3660 12248
rect 3712 12186 3740 12378
rect 4264 12306 4292 12582
rect 4356 12442 4384 12718
rect 4344 12436 4396 12442
rect 4344 12378 4396 12384
rect 4252 12300 4304 12306
rect 4252 12242 4304 12248
rect 3620 12158 3740 12186
rect 3620 11898 3648 12158
rect 4160 12096 4212 12102
rect 4160 12038 4212 12044
rect 3756 11996 4064 12005
rect 3756 11994 3762 11996
rect 3818 11994 3842 11996
rect 3898 11994 3922 11996
rect 3978 11994 4002 11996
rect 4058 11994 4064 11996
rect 3818 11942 3820 11994
rect 4000 11942 4002 11994
rect 3756 11940 3762 11942
rect 3818 11940 3842 11942
rect 3898 11940 3922 11942
rect 3978 11940 4002 11942
rect 4058 11940 4064 11942
rect 3756 11931 4064 11940
rect 3608 11892 3660 11898
rect 3608 11834 3660 11840
rect 4172 11642 4200 12038
rect 4356 11898 4384 12378
rect 4632 12306 4660 13670
rect 4724 12782 4752 13738
rect 5184 12986 5212 13806
rect 5356 13252 5408 13258
rect 5356 13194 5408 13200
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 4712 12776 4764 12782
rect 4712 12718 4764 12724
rect 4620 12300 4672 12306
rect 4620 12242 4672 12248
rect 4344 11892 4396 11898
rect 4344 11834 4396 11840
rect 4080 11626 4200 11642
rect 4068 11620 4200 11626
rect 4120 11614 4200 11620
rect 4068 11562 4120 11568
rect 4356 11218 4384 11834
rect 4344 11212 4396 11218
rect 4344 11154 4396 11160
rect 3756 10908 4064 10917
rect 3756 10906 3762 10908
rect 3818 10906 3842 10908
rect 3898 10906 3922 10908
rect 3978 10906 4002 10908
rect 4058 10906 4064 10908
rect 3818 10854 3820 10906
rect 4000 10854 4002 10906
rect 3756 10852 3762 10854
rect 3818 10852 3842 10854
rect 3898 10852 3922 10854
rect 3978 10852 4002 10854
rect 4058 10852 4064 10854
rect 3756 10843 4064 10852
rect 3516 10804 3568 10810
rect 3516 10746 3568 10752
rect 3424 10600 3476 10606
rect 3424 10542 3476 10548
rect 2700 10254 2820 10282
rect 2596 10124 2648 10130
rect 2596 10066 2648 10072
rect 2320 9512 2372 9518
rect 2320 9454 2372 9460
rect 2504 9512 2556 9518
rect 2504 9454 2556 9460
rect 2608 9466 2636 10066
rect 2700 10062 2728 10254
rect 2872 10192 2924 10198
rect 2870 10160 2872 10169
rect 2924 10160 2926 10169
rect 2870 10095 2926 10104
rect 2688 10056 2740 10062
rect 2740 10016 2820 10044
rect 2688 9998 2740 10004
rect 2688 9920 2740 9926
rect 2688 9862 2740 9868
rect 2700 9586 2728 9862
rect 2688 9580 2740 9586
rect 2688 9522 2740 9528
rect 1952 9444 2004 9450
rect 1952 9386 2004 9392
rect 1400 9172 1452 9178
rect 1400 9114 1452 9120
rect 1124 9036 1176 9042
rect 1124 8978 1176 8984
rect 1136 8634 1164 8978
rect 1124 8628 1176 8634
rect 1124 8570 1176 8576
rect 1124 7744 1176 7750
rect 1124 7686 1176 7692
rect 1136 7274 1164 7686
rect 1412 7342 1440 9114
rect 1964 8974 1992 9386
rect 2332 9042 2360 9454
rect 2608 9438 2728 9466
rect 2792 9450 2820 10016
rect 2976 9654 3004 10406
rect 3068 10390 3280 10418
rect 3146 10024 3202 10033
rect 3146 9959 3202 9968
rect 2964 9648 3016 9654
rect 2964 9590 3016 9596
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 2700 9110 2728 9438
rect 2780 9444 2832 9450
rect 2780 9386 2832 9392
rect 2884 9110 2912 9454
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 2688 9104 2740 9110
rect 2688 9046 2740 9052
rect 2872 9104 2924 9110
rect 2872 9046 2924 9052
rect 2320 9036 2372 9042
rect 2320 8978 2372 8984
rect 1952 8968 2004 8974
rect 1952 8910 2004 8916
rect 2136 8900 2188 8906
rect 2136 8842 2188 8848
rect 2148 8430 2176 8842
rect 2136 8424 2188 8430
rect 2136 8366 2188 8372
rect 2136 7540 2188 7546
rect 2136 7482 2188 7488
rect 1400 7336 1452 7342
rect 1400 7278 1452 7284
rect 1676 7336 1728 7342
rect 1676 7278 1728 7284
rect 1124 7268 1176 7274
rect 1124 7210 1176 7216
rect 1124 5568 1176 5574
rect 1124 5510 1176 5516
rect 1136 4690 1164 5510
rect 1688 5234 1716 7278
rect 2148 7002 2176 7482
rect 2228 7200 2280 7206
rect 2228 7142 2280 7148
rect 2136 6996 2188 7002
rect 2136 6938 2188 6944
rect 2240 6866 2268 7142
rect 2136 6860 2188 6866
rect 2136 6802 2188 6808
rect 2228 6860 2280 6866
rect 2228 6802 2280 6808
rect 1676 5228 1728 5234
rect 1676 5170 1728 5176
rect 1400 5024 1452 5030
rect 1400 4966 1452 4972
rect 1412 4690 1440 4966
rect 2148 4826 2176 6802
rect 2136 4820 2188 4826
rect 2136 4762 2188 4768
rect 1124 4684 1176 4690
rect 1124 4626 1176 4632
rect 1400 4684 1452 4690
rect 1400 4626 1452 4632
rect 2332 3942 2360 8978
rect 2504 8832 2556 8838
rect 2504 8774 2556 8780
rect 2596 8832 2648 8838
rect 2596 8774 2648 8780
rect 2516 8498 2544 8774
rect 2608 8634 2636 8774
rect 2596 8628 2648 8634
rect 2596 8570 2648 8576
rect 2504 8492 2556 8498
rect 2504 8434 2556 8440
rect 2596 8424 2648 8430
rect 2596 8366 2648 8372
rect 2608 7546 2636 8366
rect 2700 8362 2728 9046
rect 2780 8900 2832 8906
rect 2780 8842 2832 8848
rect 2792 8634 2820 8842
rect 2780 8628 2832 8634
rect 2780 8570 2832 8576
rect 2688 8356 2740 8362
rect 2688 8298 2740 8304
rect 2792 8242 2820 8570
rect 2700 8214 2820 8242
rect 2596 7540 2648 7546
rect 2596 7482 2648 7488
rect 2596 7336 2648 7342
rect 2596 7278 2648 7284
rect 2608 6934 2636 7278
rect 2596 6928 2648 6934
rect 2596 6870 2648 6876
rect 2700 6798 2728 8214
rect 2884 7750 2912 9046
rect 2976 8974 3004 9318
rect 3160 9042 3188 9959
rect 3148 9036 3200 9042
rect 3148 8978 3200 8984
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 3056 8832 3108 8838
rect 3056 8774 3108 8780
rect 3068 8566 3096 8774
rect 3252 8634 3280 10390
rect 3332 10260 3384 10266
rect 3332 10202 3384 10208
rect 3344 9722 3372 10202
rect 3332 9716 3384 9722
rect 3332 9658 3384 9664
rect 3436 9382 3464 10542
rect 3516 10532 3568 10538
rect 3516 10474 3568 10480
rect 3528 9926 3556 10474
rect 3608 10464 3660 10470
rect 3608 10406 3660 10412
rect 3516 9920 3568 9926
rect 3516 9862 3568 9868
rect 3620 9518 3648 10406
rect 4250 10160 4306 10169
rect 4250 10095 4306 10104
rect 4264 10062 4292 10095
rect 4252 10056 4304 10062
rect 4252 9998 4304 10004
rect 3756 9820 4064 9829
rect 3756 9818 3762 9820
rect 3818 9818 3842 9820
rect 3898 9818 3922 9820
rect 3978 9818 4002 9820
rect 4058 9818 4064 9820
rect 3818 9766 3820 9818
rect 4000 9766 4002 9818
rect 3756 9764 3762 9766
rect 3818 9764 3842 9766
rect 3898 9764 3922 9766
rect 3978 9764 4002 9766
rect 4058 9764 4064 9766
rect 3756 9755 4064 9764
rect 4264 9674 4292 9998
rect 4172 9646 4292 9674
rect 3608 9512 3660 9518
rect 3608 9454 3660 9460
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3240 8628 3292 8634
rect 3240 8570 3292 8576
rect 3056 8560 3108 8566
rect 3056 8502 3108 8508
rect 3068 8430 3096 8502
rect 3056 8424 3108 8430
rect 3056 8366 3108 8372
rect 3148 7948 3200 7954
rect 3148 7890 3200 7896
rect 2872 7744 2924 7750
rect 2872 7686 2924 7692
rect 2964 6860 3016 6866
rect 2964 6802 3016 6808
rect 2688 6792 2740 6798
rect 2688 6734 2740 6740
rect 2976 6186 3004 6802
rect 3160 6730 3188 7890
rect 3240 7880 3292 7886
rect 3240 7822 3292 7828
rect 3252 7546 3280 7822
rect 3240 7540 3292 7546
rect 3240 7482 3292 7488
rect 3332 7404 3384 7410
rect 3332 7346 3384 7352
rect 3240 7268 3292 7274
rect 3240 7210 3292 7216
rect 3252 6866 3280 7210
rect 3344 6934 3372 7346
rect 3332 6928 3384 6934
rect 3332 6870 3384 6876
rect 3240 6860 3292 6866
rect 3240 6802 3292 6808
rect 3148 6724 3200 6730
rect 3148 6666 3200 6672
rect 2964 6180 3016 6186
rect 2964 6122 3016 6128
rect 2412 5568 2464 5574
rect 2412 5510 2464 5516
rect 2424 5166 2452 5510
rect 2412 5160 2464 5166
rect 2412 5102 2464 5108
rect 2976 4826 3004 6122
rect 3056 5772 3108 5778
rect 3056 5714 3108 5720
rect 3068 5370 3096 5714
rect 3148 5568 3200 5574
rect 3252 5556 3280 6802
rect 3436 5914 3464 9318
rect 4172 9178 4200 9646
rect 4160 9172 4212 9178
rect 4160 9114 4212 9120
rect 3756 8732 4064 8741
rect 3756 8730 3762 8732
rect 3818 8730 3842 8732
rect 3898 8730 3922 8732
rect 3978 8730 4002 8732
rect 4058 8730 4064 8732
rect 3818 8678 3820 8730
rect 4000 8678 4002 8730
rect 3756 8676 3762 8678
rect 3818 8676 3842 8678
rect 3898 8676 3922 8678
rect 3978 8676 4002 8678
rect 4058 8676 4064 8678
rect 3756 8667 4064 8676
rect 4172 8430 4200 9114
rect 4160 8424 4212 8430
rect 4160 8366 4212 8372
rect 4252 8356 4304 8362
rect 4252 8298 4304 8304
rect 4264 7818 4292 8298
rect 4436 7948 4488 7954
rect 4436 7890 4488 7896
rect 4252 7812 4304 7818
rect 4252 7754 4304 7760
rect 3756 7644 4064 7653
rect 3756 7642 3762 7644
rect 3818 7642 3842 7644
rect 3898 7642 3922 7644
rect 3978 7642 4002 7644
rect 4058 7642 4064 7644
rect 3818 7590 3820 7642
rect 4000 7590 4002 7642
rect 3756 7588 3762 7590
rect 3818 7588 3842 7590
rect 3898 7588 3922 7590
rect 3978 7588 4002 7590
rect 4058 7588 4064 7590
rect 3756 7579 4064 7588
rect 4448 7546 4476 7890
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 3516 7336 3568 7342
rect 4620 7336 4672 7342
rect 3568 7296 3648 7324
rect 3516 7278 3568 7284
rect 3620 6866 3648 7296
rect 4620 7278 4672 7284
rect 4068 7268 4120 7274
rect 4068 7210 4120 7216
rect 3608 6860 3660 6866
rect 3608 6802 3660 6808
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3528 6254 3556 6598
rect 3620 6390 3648 6802
rect 4080 6746 4108 7210
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 4264 6866 4292 7142
rect 4252 6860 4304 6866
rect 4252 6802 4304 6808
rect 4632 6798 4660 7278
rect 4724 7206 4752 12718
rect 4804 12708 4856 12714
rect 4804 12650 4856 12656
rect 4816 12238 4844 12650
rect 5184 12442 5212 12922
rect 5172 12436 5224 12442
rect 5172 12378 5224 12384
rect 5368 12306 5396 13194
rect 5460 13190 5488 13806
rect 5828 13326 5856 14470
rect 5920 14278 5948 18924
rect 6000 18828 6052 18834
rect 6000 18770 6052 18776
rect 6092 18828 6144 18834
rect 6092 18770 6144 18776
rect 6012 18086 6040 18770
rect 6104 18426 6132 18770
rect 6092 18420 6144 18426
rect 6092 18362 6144 18368
rect 6000 18080 6052 18086
rect 6000 18022 6052 18028
rect 6196 17184 6224 19094
rect 6368 18964 6420 18970
rect 6368 18906 6420 18912
rect 6380 18222 6408 18906
rect 6472 18698 6500 19110
rect 6552 18896 6604 18902
rect 6552 18838 6604 18844
rect 6460 18692 6512 18698
rect 6460 18634 6512 18640
rect 6472 18358 6500 18634
rect 6460 18352 6512 18358
rect 6460 18294 6512 18300
rect 6368 18216 6420 18222
rect 6368 18158 6420 18164
rect 6276 18080 6328 18086
rect 6276 18022 6328 18028
rect 6288 17338 6316 18022
rect 6472 17746 6500 18294
rect 6564 18290 6592 18838
rect 6552 18284 6604 18290
rect 6552 18226 6604 18232
rect 6460 17740 6512 17746
rect 6460 17682 6512 17688
rect 6460 17536 6512 17542
rect 6460 17478 6512 17484
rect 6276 17332 6328 17338
rect 6276 17274 6328 17280
rect 6012 17156 6224 17184
rect 5908 14272 5960 14278
rect 5908 14214 5960 14220
rect 5816 13320 5868 13326
rect 5816 13262 5868 13268
rect 5448 13184 5500 13190
rect 5448 13126 5500 13132
rect 5460 12918 5488 13126
rect 5448 12912 5500 12918
rect 5448 12854 5500 12860
rect 6012 12646 6040 17156
rect 6472 17134 6500 17478
rect 6564 17202 6592 18226
rect 6552 17196 6604 17202
rect 6552 17138 6604 17144
rect 6656 17134 6684 22986
rect 7116 22710 7144 23122
rect 7104 22704 7156 22710
rect 7104 22646 7156 22652
rect 7576 22642 7604 23122
rect 7564 22636 7616 22642
rect 7564 22578 7616 22584
rect 7472 22568 7524 22574
rect 7472 22510 7524 22516
rect 6920 22432 6972 22438
rect 6920 22374 6972 22380
rect 7012 22432 7064 22438
rect 7012 22374 7064 22380
rect 6932 22098 6960 22374
rect 6736 22092 6788 22098
rect 6736 22034 6788 22040
rect 6920 22092 6972 22098
rect 6920 22034 6972 22040
rect 6748 21622 6776 22034
rect 6736 21616 6788 21622
rect 6736 21558 6788 21564
rect 7024 21554 7052 22374
rect 7114 22332 7422 22341
rect 7114 22330 7120 22332
rect 7176 22330 7200 22332
rect 7256 22330 7280 22332
rect 7336 22330 7360 22332
rect 7416 22330 7422 22332
rect 7176 22278 7178 22330
rect 7358 22278 7360 22330
rect 7114 22276 7120 22278
rect 7176 22276 7200 22278
rect 7256 22276 7280 22278
rect 7336 22276 7360 22278
rect 7416 22276 7422 22278
rect 7114 22267 7422 22276
rect 7484 22234 7512 22510
rect 7564 22500 7616 22506
rect 7564 22442 7616 22448
rect 7472 22228 7524 22234
rect 7472 22170 7524 22176
rect 7576 21690 7604 22442
rect 7668 22030 7696 25298
rect 7840 24744 7892 24750
rect 7840 24686 7892 24692
rect 7852 24410 7880 24686
rect 7840 24404 7892 24410
rect 7840 24346 7892 24352
rect 7840 23656 7892 23662
rect 7840 23598 7892 23604
rect 7748 23520 7800 23526
rect 7748 23462 7800 23468
rect 7760 23225 7788 23462
rect 7746 23216 7802 23225
rect 7746 23151 7802 23160
rect 7656 22024 7708 22030
rect 7656 21966 7708 21972
rect 7564 21684 7616 21690
rect 7564 21626 7616 21632
rect 7012 21548 7064 21554
rect 7012 21490 7064 21496
rect 6736 21480 6788 21486
rect 6736 21422 6788 21428
rect 6748 21078 6776 21422
rect 7012 21412 7064 21418
rect 7012 21354 7064 21360
rect 6736 21072 6788 21078
rect 6736 21014 6788 21020
rect 6748 20602 6776 21014
rect 6828 21004 6880 21010
rect 6828 20946 6880 20952
rect 6736 20596 6788 20602
rect 6736 20538 6788 20544
rect 6736 19916 6788 19922
rect 6736 19858 6788 19864
rect 6748 19514 6776 19858
rect 6736 19508 6788 19514
rect 6736 19450 6788 19456
rect 6460 17128 6512 17134
rect 6460 17070 6512 17076
rect 6644 17128 6696 17134
rect 6644 17070 6696 17076
rect 6092 17060 6144 17066
rect 6092 17002 6144 17008
rect 6104 16658 6132 17002
rect 6368 16992 6420 16998
rect 6368 16934 6420 16940
rect 6380 16658 6408 16934
rect 6840 16658 6868 20946
rect 7024 20874 7052 21354
rect 7472 21344 7524 21350
rect 7472 21286 7524 21292
rect 7114 21244 7422 21253
rect 7114 21242 7120 21244
rect 7176 21242 7200 21244
rect 7256 21242 7280 21244
rect 7336 21242 7360 21244
rect 7416 21242 7422 21244
rect 7176 21190 7178 21242
rect 7358 21190 7360 21242
rect 7114 21188 7120 21190
rect 7176 21188 7200 21190
rect 7256 21188 7280 21190
rect 7336 21188 7360 21190
rect 7416 21188 7422 21190
rect 7114 21179 7422 21188
rect 7012 20868 7064 20874
rect 7012 20810 7064 20816
rect 7484 20398 7512 21286
rect 7472 20392 7524 20398
rect 7472 20334 7524 20340
rect 7114 20156 7422 20165
rect 7114 20154 7120 20156
rect 7176 20154 7200 20156
rect 7256 20154 7280 20156
rect 7336 20154 7360 20156
rect 7416 20154 7422 20156
rect 7176 20102 7178 20154
rect 7358 20102 7360 20154
rect 7114 20100 7120 20102
rect 7176 20100 7200 20102
rect 7256 20100 7280 20102
rect 7336 20100 7360 20102
rect 7416 20100 7422 20102
rect 7114 20091 7422 20100
rect 7484 19922 7512 20334
rect 7472 19916 7524 19922
rect 7472 19858 7524 19864
rect 7484 19394 7512 19858
rect 7208 19366 7604 19394
rect 7208 19310 7236 19366
rect 7196 19304 7248 19310
rect 7196 19246 7248 19252
rect 7472 19168 7524 19174
rect 7472 19110 7524 19116
rect 7114 19068 7422 19077
rect 7114 19066 7120 19068
rect 7176 19066 7200 19068
rect 7256 19066 7280 19068
rect 7336 19066 7360 19068
rect 7416 19066 7422 19068
rect 7176 19014 7178 19066
rect 7358 19014 7360 19066
rect 7114 19012 7120 19014
rect 7176 19012 7200 19014
rect 7256 19012 7280 19014
rect 7336 19012 7360 19014
rect 7416 19012 7422 19014
rect 7114 19003 7422 19012
rect 7288 18828 7340 18834
rect 7288 18770 7340 18776
rect 7300 18426 7328 18770
rect 7288 18420 7340 18426
rect 7288 18362 7340 18368
rect 7114 17980 7422 17989
rect 7114 17978 7120 17980
rect 7176 17978 7200 17980
rect 7256 17978 7280 17980
rect 7336 17978 7360 17980
rect 7416 17978 7422 17980
rect 7176 17926 7178 17978
rect 7358 17926 7360 17978
rect 7114 17924 7120 17926
rect 7176 17924 7200 17926
rect 7256 17924 7280 17926
rect 7336 17924 7360 17926
rect 7416 17924 7422 17926
rect 7114 17915 7422 17924
rect 7288 17876 7340 17882
rect 7024 17836 7288 17864
rect 6920 17808 6972 17814
rect 7024 17796 7052 17836
rect 7288 17818 7340 17824
rect 7484 17814 7512 19110
rect 7576 18290 7604 19366
rect 7760 19310 7788 23151
rect 7852 23050 7880 23598
rect 7840 23044 7892 23050
rect 7840 22986 7892 22992
rect 7840 21548 7892 21554
rect 7840 21490 7892 21496
rect 7748 19304 7800 19310
rect 7748 19246 7800 19252
rect 7656 19168 7708 19174
rect 7656 19110 7708 19116
rect 7564 18284 7616 18290
rect 7564 18226 7616 18232
rect 6972 17768 7052 17796
rect 7472 17808 7524 17814
rect 6920 17750 6972 17756
rect 7472 17750 7524 17756
rect 7472 17672 7524 17678
rect 7472 17614 7524 17620
rect 7114 16892 7422 16901
rect 7114 16890 7120 16892
rect 7176 16890 7200 16892
rect 7256 16890 7280 16892
rect 7336 16890 7360 16892
rect 7416 16890 7422 16892
rect 7176 16838 7178 16890
rect 7358 16838 7360 16890
rect 7114 16836 7120 16838
rect 7176 16836 7200 16838
rect 7256 16836 7280 16838
rect 7336 16836 7360 16838
rect 7416 16836 7422 16838
rect 7114 16827 7422 16836
rect 7484 16794 7512 17614
rect 7576 17134 7604 18226
rect 7668 18222 7696 19110
rect 7656 18216 7708 18222
rect 7656 18158 7708 18164
rect 7852 18086 7880 21490
rect 7944 20262 7972 25638
rect 8300 25424 8352 25430
rect 8300 25366 8352 25372
rect 8312 24274 8340 25366
rect 8404 24818 8432 25774
rect 9232 25770 9260 26386
rect 9416 25906 9444 26794
rect 9588 26444 9640 26450
rect 9588 26386 9640 26392
rect 9404 25900 9456 25906
rect 9404 25842 9456 25848
rect 9220 25764 9272 25770
rect 9220 25706 9272 25712
rect 9404 25696 9456 25702
rect 9404 25638 9456 25644
rect 8852 25288 8904 25294
rect 8852 25230 8904 25236
rect 8392 24812 8444 24818
rect 8392 24754 8444 24760
rect 8760 24676 8812 24682
rect 8864 24664 8892 25230
rect 8812 24636 8892 24664
rect 8760 24618 8812 24624
rect 8864 24410 8892 24636
rect 9312 24676 9364 24682
rect 9312 24618 9364 24624
rect 9324 24410 9352 24618
rect 8852 24404 8904 24410
rect 8852 24346 8904 24352
rect 9312 24404 9364 24410
rect 9312 24346 9364 24352
rect 9416 24274 9444 25638
rect 9600 25362 9628 26386
rect 9680 26240 9732 26246
rect 9680 26182 9732 26188
rect 9692 25362 9720 26182
rect 9784 26042 9812 26862
rect 9772 26036 9824 26042
rect 9772 25978 9824 25984
rect 9876 25888 9904 27270
rect 10048 27124 10100 27130
rect 10048 27066 10100 27072
rect 9956 26512 10008 26518
rect 9956 26454 10008 26460
rect 9784 25860 9904 25888
rect 9588 25356 9640 25362
rect 9588 25298 9640 25304
rect 9680 25356 9732 25362
rect 9680 25298 9732 25304
rect 9600 24954 9628 25298
rect 9680 25220 9732 25226
rect 9680 25162 9732 25168
rect 9588 24948 9640 24954
rect 9588 24890 9640 24896
rect 9496 24744 9548 24750
rect 9496 24686 9548 24692
rect 8024 24268 8076 24274
rect 8024 24210 8076 24216
rect 8300 24268 8352 24274
rect 8300 24210 8352 24216
rect 9404 24268 9456 24274
rect 9404 24210 9456 24216
rect 7932 20256 7984 20262
rect 7932 20198 7984 20204
rect 7840 18080 7892 18086
rect 7840 18022 7892 18028
rect 7840 17604 7892 17610
rect 7840 17546 7892 17552
rect 7564 17128 7616 17134
rect 7564 17070 7616 17076
rect 7472 16788 7524 16794
rect 7472 16730 7524 16736
rect 7576 16726 7604 17070
rect 7656 17060 7708 17066
rect 7656 17002 7708 17008
rect 7668 16794 7696 17002
rect 7656 16788 7708 16794
rect 7656 16730 7708 16736
rect 7564 16720 7616 16726
rect 7564 16662 7616 16668
rect 7852 16658 7880 17546
rect 8036 16794 8064 24210
rect 8760 24064 8812 24070
rect 8760 24006 8812 24012
rect 8576 23316 8628 23322
rect 8576 23258 8628 23264
rect 8300 23248 8352 23254
rect 8300 23190 8352 23196
rect 8116 21004 8168 21010
rect 8116 20946 8168 20952
rect 8128 20602 8156 20946
rect 8116 20596 8168 20602
rect 8116 20538 8168 20544
rect 8116 19508 8168 19514
rect 8116 19450 8168 19456
rect 8128 17542 8156 19450
rect 8312 18086 8340 23190
rect 8484 22432 8536 22438
rect 8484 22374 8536 22380
rect 8392 21344 8444 21350
rect 8496 21332 8524 22374
rect 8588 22098 8616 23258
rect 8772 23254 8800 24006
rect 9508 23730 9536 24686
rect 9692 24274 9720 25162
rect 9680 24268 9732 24274
rect 9680 24210 9732 24216
rect 9496 23724 9548 23730
rect 9496 23666 9548 23672
rect 8760 23248 8812 23254
rect 8760 23190 8812 23196
rect 9508 23186 9536 23666
rect 9496 23180 9548 23186
rect 9496 23122 9548 23128
rect 9680 23112 9732 23118
rect 9680 23054 9732 23060
rect 9128 22976 9180 22982
rect 9128 22918 9180 22924
rect 9140 22778 9168 22918
rect 9128 22772 9180 22778
rect 9128 22714 9180 22720
rect 8760 22500 8812 22506
rect 8760 22442 8812 22448
rect 8852 22500 8904 22506
rect 8852 22442 8904 22448
rect 8772 22234 8800 22442
rect 8760 22228 8812 22234
rect 8760 22170 8812 22176
rect 8576 22092 8628 22098
rect 8576 22034 8628 22040
rect 8864 22030 8892 22442
rect 9140 22094 9168 22714
rect 9048 22066 9168 22094
rect 9404 22092 9456 22098
rect 8852 22024 8904 22030
rect 8852 21966 8904 21972
rect 8668 21684 8720 21690
rect 8668 21626 8720 21632
rect 8576 21344 8628 21350
rect 8496 21304 8576 21332
rect 8392 21286 8444 21292
rect 8576 21286 8628 21292
rect 8404 20398 8432 21286
rect 8484 21072 8536 21078
rect 8484 21014 8536 21020
rect 8496 20602 8524 21014
rect 8588 21010 8616 21286
rect 8576 21004 8628 21010
rect 8576 20946 8628 20952
rect 8680 20806 8708 21626
rect 8760 21004 8812 21010
rect 8760 20946 8812 20952
rect 8668 20800 8720 20806
rect 8668 20742 8720 20748
rect 8484 20596 8536 20602
rect 8484 20538 8536 20544
rect 8392 20392 8444 20398
rect 8392 20334 8444 20340
rect 8496 20330 8524 20538
rect 8484 20324 8536 20330
rect 8484 20266 8536 20272
rect 8392 19712 8444 19718
rect 8392 19654 8444 19660
rect 8404 19242 8432 19654
rect 8392 19236 8444 19242
rect 8392 19178 8444 19184
rect 8576 19236 8628 19242
rect 8576 19178 8628 19184
rect 8588 18970 8616 19178
rect 8772 19174 8800 20946
rect 8864 20942 8892 21966
rect 9048 21690 9076 22066
rect 9404 22034 9456 22040
rect 9496 22094 9548 22098
rect 9692 22094 9720 23054
rect 9784 22778 9812 25860
rect 9864 25764 9916 25770
rect 9864 25706 9916 25712
rect 9772 22772 9824 22778
rect 9772 22714 9824 22720
rect 9876 22094 9904 25706
rect 9968 25480 9996 26454
rect 10060 26450 10088 27066
rect 10140 26852 10192 26858
rect 10140 26794 10192 26800
rect 10048 26444 10100 26450
rect 10048 26386 10100 26392
rect 10060 25702 10088 26386
rect 10152 25838 10180 26794
rect 10232 26784 10284 26790
rect 10232 26726 10284 26732
rect 10244 26450 10272 26726
rect 10232 26444 10284 26450
rect 10232 26386 10284 26392
rect 10232 26308 10284 26314
rect 10232 26250 10284 26256
rect 10244 26042 10272 26250
rect 10232 26036 10284 26042
rect 10232 25978 10284 25984
rect 10140 25832 10192 25838
rect 10140 25774 10192 25780
rect 10048 25696 10100 25702
rect 10048 25638 10100 25644
rect 10048 25492 10100 25498
rect 9968 25452 10048 25480
rect 9968 24410 9996 25452
rect 10048 25434 10100 25440
rect 10152 25362 10180 25774
rect 10140 25356 10192 25362
rect 10140 25298 10192 25304
rect 10152 24954 10180 25298
rect 10140 24948 10192 24954
rect 10140 24890 10192 24896
rect 10048 24812 10100 24818
rect 10048 24754 10100 24760
rect 9956 24404 10008 24410
rect 9956 24346 10008 24352
rect 10060 24274 10088 24754
rect 10048 24268 10100 24274
rect 10048 24210 10100 24216
rect 9956 23588 10008 23594
rect 9956 23530 10008 23536
rect 9968 23322 9996 23530
rect 10060 23526 10088 24210
rect 10244 24206 10272 25978
rect 10336 25770 10364 27882
rect 10888 27538 10916 27950
rect 10876 27532 10928 27538
rect 10876 27474 10928 27480
rect 10876 27328 10928 27334
rect 10876 27270 10928 27276
rect 10472 27228 10780 27237
rect 10472 27226 10478 27228
rect 10534 27226 10558 27228
rect 10614 27226 10638 27228
rect 10694 27226 10718 27228
rect 10774 27226 10780 27228
rect 10534 27174 10536 27226
rect 10716 27174 10718 27226
rect 10472 27172 10478 27174
rect 10534 27172 10558 27174
rect 10614 27172 10638 27174
rect 10694 27172 10718 27174
rect 10774 27172 10780 27174
rect 10472 27163 10780 27172
rect 10508 26920 10560 26926
rect 10508 26862 10560 26868
rect 10784 26920 10836 26926
rect 10888 26908 10916 27270
rect 11072 26926 11100 28358
rect 11164 28150 11192 28970
rect 11336 28960 11388 28966
rect 11336 28902 11388 28908
rect 11244 28484 11296 28490
rect 11244 28426 11296 28432
rect 11152 28144 11204 28150
rect 11152 28086 11204 28092
rect 11164 27606 11192 28086
rect 11256 28014 11284 28426
rect 11348 28422 11376 28902
rect 11336 28416 11388 28422
rect 11336 28358 11388 28364
rect 11440 28098 11468 29022
rect 12164 29028 12216 29034
rect 12164 28970 12216 28976
rect 11520 28688 11572 28694
rect 11520 28630 11572 28636
rect 11348 28082 11468 28098
rect 11336 28076 11468 28082
rect 11388 28070 11468 28076
rect 11336 28018 11388 28024
rect 11244 28008 11296 28014
rect 11244 27950 11296 27956
rect 11532 27878 11560 28630
rect 11796 28416 11848 28422
rect 11796 28358 11848 28364
rect 11612 27940 11664 27946
rect 11612 27882 11664 27888
rect 11520 27872 11572 27878
rect 11520 27814 11572 27820
rect 11624 27674 11652 27882
rect 11612 27668 11664 27674
rect 11612 27610 11664 27616
rect 11152 27600 11204 27606
rect 11152 27542 11204 27548
rect 11808 27538 11836 28358
rect 11796 27532 11848 27538
rect 11796 27474 11848 27480
rect 11980 27328 12032 27334
rect 11980 27270 12032 27276
rect 11992 26926 12020 27270
rect 10836 26880 10916 26908
rect 10784 26862 10836 26868
rect 10520 26314 10548 26862
rect 10508 26308 10560 26314
rect 10508 26250 10560 26256
rect 10472 26140 10780 26149
rect 10472 26138 10478 26140
rect 10534 26138 10558 26140
rect 10614 26138 10638 26140
rect 10694 26138 10718 26140
rect 10774 26138 10780 26140
rect 10534 26086 10536 26138
rect 10716 26086 10718 26138
rect 10472 26084 10478 26086
rect 10534 26084 10558 26086
rect 10614 26084 10638 26086
rect 10694 26084 10718 26086
rect 10774 26084 10780 26086
rect 10472 26075 10780 26084
rect 10888 25906 10916 26880
rect 11060 26920 11112 26926
rect 11060 26862 11112 26868
rect 11152 26920 11204 26926
rect 11152 26862 11204 26868
rect 11980 26920 12032 26926
rect 11980 26862 12032 26868
rect 11164 26790 11192 26862
rect 11152 26784 11204 26790
rect 11428 26784 11480 26790
rect 11204 26744 11284 26772
rect 11152 26726 11204 26732
rect 10968 26240 11020 26246
rect 10968 26182 11020 26188
rect 10980 25974 11008 26182
rect 10968 25968 11020 25974
rect 10968 25910 11020 25916
rect 11060 25968 11112 25974
rect 11060 25910 11112 25916
rect 10876 25900 10928 25906
rect 10876 25842 10928 25848
rect 10324 25764 10376 25770
rect 10324 25706 10376 25712
rect 10324 25220 10376 25226
rect 10324 25162 10376 25168
rect 10336 24682 10364 25162
rect 10980 25158 11008 25910
rect 11072 25430 11100 25910
rect 11152 25900 11204 25906
rect 11152 25842 11204 25848
rect 11060 25424 11112 25430
rect 11060 25366 11112 25372
rect 11164 25362 11192 25842
rect 11256 25838 11284 26744
rect 11428 26726 11480 26732
rect 11612 26784 11664 26790
rect 11612 26726 11664 26732
rect 11440 26586 11468 26726
rect 11428 26580 11480 26586
rect 11428 26522 11480 26528
rect 11624 26450 11652 26726
rect 11704 26512 11756 26518
rect 11704 26454 11756 26460
rect 11612 26444 11664 26450
rect 11612 26386 11664 26392
rect 11428 26376 11480 26382
rect 11428 26318 11480 26324
rect 11244 25832 11296 25838
rect 11244 25774 11296 25780
rect 11152 25356 11204 25362
rect 11152 25298 11204 25304
rect 10968 25152 11020 25158
rect 10968 25094 11020 25100
rect 10472 25052 10780 25061
rect 10472 25050 10478 25052
rect 10534 25050 10558 25052
rect 10614 25050 10638 25052
rect 10694 25050 10718 25052
rect 10774 25050 10780 25052
rect 10534 24998 10536 25050
rect 10716 24998 10718 25050
rect 10472 24996 10478 24998
rect 10534 24996 10558 24998
rect 10614 24996 10638 24998
rect 10694 24996 10718 24998
rect 10774 24996 10780 24998
rect 10472 24987 10780 24996
rect 10324 24676 10376 24682
rect 10324 24618 10376 24624
rect 10324 24404 10376 24410
rect 10324 24346 10376 24352
rect 10232 24200 10284 24206
rect 10232 24142 10284 24148
rect 10140 24064 10192 24070
rect 10140 24006 10192 24012
rect 10048 23520 10100 23526
rect 10048 23462 10100 23468
rect 9956 23316 10008 23322
rect 9956 23258 10008 23264
rect 10060 23118 10088 23462
rect 10152 23186 10180 24006
rect 10244 23866 10272 24142
rect 10232 23860 10284 23866
rect 10232 23802 10284 23808
rect 10336 23338 10364 24346
rect 10980 24256 11008 25094
rect 11164 24818 11192 25298
rect 11256 24954 11284 25774
rect 11244 24948 11296 24954
rect 11244 24890 11296 24896
rect 11152 24812 11204 24818
rect 11152 24754 11204 24760
rect 11164 24614 11192 24754
rect 11152 24608 11204 24614
rect 11152 24550 11204 24556
rect 10888 24228 11008 24256
rect 11152 24268 11204 24274
rect 10888 24070 10916 24228
rect 11152 24210 11204 24216
rect 10968 24132 11020 24138
rect 10968 24074 11020 24080
rect 10876 24064 10928 24070
rect 10876 24006 10928 24012
rect 10472 23964 10780 23973
rect 10472 23962 10478 23964
rect 10534 23962 10558 23964
rect 10614 23962 10638 23964
rect 10694 23962 10718 23964
rect 10774 23962 10780 23964
rect 10534 23910 10536 23962
rect 10716 23910 10718 23962
rect 10472 23908 10478 23910
rect 10534 23908 10558 23910
rect 10614 23908 10638 23910
rect 10694 23908 10718 23910
rect 10774 23908 10780 23910
rect 10472 23899 10780 23908
rect 10888 23730 10916 24006
rect 10508 23724 10560 23730
rect 10508 23666 10560 23672
rect 10876 23724 10928 23730
rect 10876 23666 10928 23672
rect 10244 23310 10364 23338
rect 10140 23180 10192 23186
rect 10140 23122 10192 23128
rect 10048 23112 10100 23118
rect 10048 23054 10100 23060
rect 10140 22432 10192 22438
rect 10140 22374 10192 22380
rect 10152 22166 10180 22374
rect 10244 22234 10272 23310
rect 10322 23216 10378 23225
rect 10322 23151 10324 23160
rect 10376 23151 10378 23160
rect 10324 23122 10376 23128
rect 10520 23066 10548 23666
rect 10336 23038 10548 23066
rect 10232 22228 10284 22234
rect 10232 22170 10284 22176
rect 10140 22160 10192 22166
rect 10140 22102 10192 22108
rect 9496 22092 9720 22094
rect 9548 22066 9720 22092
rect 9784 22066 9904 22094
rect 9496 22034 9548 22040
rect 9416 21894 9444 22034
rect 9404 21888 9456 21894
rect 9404 21830 9456 21836
rect 9036 21684 9088 21690
rect 9036 21626 9088 21632
rect 8944 21616 8996 21622
rect 8944 21558 8996 21564
rect 8956 21418 8984 21558
rect 8944 21412 8996 21418
rect 8944 21354 8996 21360
rect 9784 21146 9812 22066
rect 10140 22024 10192 22030
rect 10140 21966 10192 21972
rect 9956 21888 10008 21894
rect 9956 21830 10008 21836
rect 9772 21140 9824 21146
rect 9772 21082 9824 21088
rect 9678 21040 9734 21049
rect 9678 20975 9680 20984
rect 9732 20975 9734 20984
rect 9680 20946 9732 20952
rect 8852 20936 8904 20942
rect 8852 20878 8904 20884
rect 9588 20936 9640 20942
rect 9588 20878 9640 20884
rect 8852 20800 8904 20806
rect 8852 20742 8904 20748
rect 8864 19922 8892 20742
rect 9600 20380 9628 20878
rect 9680 20868 9732 20874
rect 9680 20810 9732 20816
rect 9692 20505 9720 20810
rect 9678 20496 9734 20505
rect 9678 20431 9734 20440
rect 9680 20392 9732 20398
rect 9600 20352 9680 20380
rect 9036 20324 9088 20330
rect 9036 20266 9088 20272
rect 9048 20058 9076 20266
rect 9036 20052 9088 20058
rect 9036 19994 9088 20000
rect 8852 19916 8904 19922
rect 8852 19858 8904 19864
rect 9496 19236 9548 19242
rect 9496 19178 9548 19184
rect 8760 19168 8812 19174
rect 8760 19110 8812 19116
rect 8944 19168 8996 19174
rect 8944 19110 8996 19116
rect 8576 18964 8628 18970
rect 8576 18906 8628 18912
rect 8576 18828 8628 18834
rect 8576 18770 8628 18776
rect 8392 18624 8444 18630
rect 8392 18566 8444 18572
rect 8300 18080 8352 18086
rect 8300 18022 8352 18028
rect 8404 17898 8432 18566
rect 8588 18426 8616 18770
rect 8576 18420 8628 18426
rect 8576 18362 8628 18368
rect 8956 18222 8984 19110
rect 8944 18216 8996 18222
rect 8944 18158 8996 18164
rect 9508 18154 9536 19178
rect 9600 18766 9628 20352
rect 9680 20334 9732 20340
rect 9784 19242 9812 21082
rect 9864 21072 9916 21078
rect 9864 21014 9916 21020
rect 9876 19922 9904 21014
rect 9864 19916 9916 19922
rect 9864 19858 9916 19864
rect 9772 19236 9824 19242
rect 9772 19178 9824 19184
rect 9588 18760 9640 18766
rect 9588 18702 9640 18708
rect 9600 18154 9628 18702
rect 9496 18148 9548 18154
rect 9496 18090 9548 18096
rect 9588 18148 9640 18154
rect 9588 18090 9640 18096
rect 8312 17870 8432 17898
rect 8116 17536 8168 17542
rect 8116 17478 8168 17484
rect 8024 16788 8076 16794
rect 8024 16730 8076 16736
rect 6092 16652 6144 16658
rect 6092 16594 6144 16600
rect 6368 16652 6420 16658
rect 6368 16594 6420 16600
rect 6644 16652 6696 16658
rect 6644 16594 6696 16600
rect 6828 16652 6880 16658
rect 6828 16594 6880 16600
rect 7840 16652 7892 16658
rect 7840 16594 7892 16600
rect 6104 14958 6132 16594
rect 6460 16040 6512 16046
rect 6460 15982 6512 15988
rect 6472 15706 6500 15982
rect 6552 15904 6604 15910
rect 6552 15846 6604 15852
rect 6460 15700 6512 15706
rect 6460 15642 6512 15648
rect 6184 15632 6236 15638
rect 6184 15574 6236 15580
rect 6092 14952 6144 14958
rect 6092 14894 6144 14900
rect 6196 14890 6224 15574
rect 6276 15496 6328 15502
rect 6276 15438 6328 15444
rect 6288 15366 6316 15438
rect 6276 15360 6328 15366
rect 6276 15302 6328 15308
rect 6564 14958 6592 15846
rect 6552 14952 6604 14958
rect 6552 14894 6604 14900
rect 6184 14884 6236 14890
rect 6184 14826 6236 14832
rect 6196 14278 6224 14826
rect 6184 14272 6236 14278
rect 6184 14214 6236 14220
rect 6276 14272 6328 14278
rect 6276 14214 6328 14220
rect 6288 13394 6316 14214
rect 6656 13870 6684 16594
rect 7114 15804 7422 15813
rect 7114 15802 7120 15804
rect 7176 15802 7200 15804
rect 7256 15802 7280 15804
rect 7336 15802 7360 15804
rect 7416 15802 7422 15804
rect 7176 15750 7178 15802
rect 7358 15750 7360 15802
rect 7114 15748 7120 15750
rect 7176 15748 7200 15750
rect 7256 15748 7280 15750
rect 7336 15748 7360 15750
rect 7416 15748 7422 15750
rect 7114 15739 7422 15748
rect 7012 15700 7064 15706
rect 7012 15642 7064 15648
rect 6920 15156 6972 15162
rect 6920 15098 6972 15104
rect 6932 14278 6960 15098
rect 7024 14346 7052 15642
rect 7196 15360 7248 15366
rect 7196 15302 7248 15308
rect 7748 15360 7800 15366
rect 7748 15302 7800 15308
rect 7208 15162 7236 15302
rect 7196 15156 7248 15162
rect 7196 15098 7248 15104
rect 7760 14958 7788 15302
rect 8128 15162 8156 17478
rect 8208 15564 8260 15570
rect 8312 15552 8340 17870
rect 8668 17672 8720 17678
rect 8668 17614 8720 17620
rect 8680 17338 8708 17614
rect 9036 17536 9088 17542
rect 9036 17478 9088 17484
rect 8668 17332 8720 17338
rect 8668 17274 8720 17280
rect 9048 17134 9076 17478
rect 8392 17128 8444 17134
rect 8392 17070 8444 17076
rect 9036 17128 9088 17134
rect 9036 17070 9088 17076
rect 8260 15524 8340 15552
rect 8208 15506 8260 15512
rect 8116 15156 8168 15162
rect 8116 15098 8168 15104
rect 7748 14952 7800 14958
rect 7748 14894 7800 14900
rect 7932 14952 7984 14958
rect 7932 14894 7984 14900
rect 7748 14816 7800 14822
rect 7748 14758 7800 14764
rect 7114 14716 7422 14725
rect 7114 14714 7120 14716
rect 7176 14714 7200 14716
rect 7256 14714 7280 14716
rect 7336 14714 7360 14716
rect 7416 14714 7422 14716
rect 7176 14662 7178 14714
rect 7358 14662 7360 14714
rect 7114 14660 7120 14662
rect 7176 14660 7200 14662
rect 7256 14660 7280 14662
rect 7336 14660 7360 14662
rect 7416 14660 7422 14662
rect 7114 14651 7422 14660
rect 7760 14482 7788 14758
rect 7944 14550 7972 14894
rect 7932 14544 7984 14550
rect 7932 14486 7984 14492
rect 7656 14476 7708 14482
rect 7656 14418 7708 14424
rect 7748 14476 7800 14482
rect 7748 14418 7800 14424
rect 7472 14408 7524 14414
rect 7472 14350 7524 14356
rect 7012 14340 7064 14346
rect 7012 14282 7064 14288
rect 6920 14272 6972 14278
rect 6920 14214 6972 14220
rect 6552 13864 6604 13870
rect 6552 13806 6604 13812
rect 6644 13864 6696 13870
rect 6644 13806 6696 13812
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6564 13530 6592 13806
rect 6736 13728 6788 13734
rect 6736 13670 6788 13676
rect 6552 13524 6604 13530
rect 6552 13466 6604 13472
rect 6748 13394 6776 13670
rect 6184 13388 6236 13394
rect 6184 13330 6236 13336
rect 6276 13388 6328 13394
rect 6276 13330 6328 13336
rect 6368 13388 6420 13394
rect 6368 13330 6420 13336
rect 6736 13388 6788 13394
rect 6736 13330 6788 13336
rect 6092 13320 6144 13326
rect 6092 13262 6144 13268
rect 6000 12640 6052 12646
rect 6000 12582 6052 12588
rect 5356 12300 5408 12306
rect 5356 12242 5408 12248
rect 5908 12300 5960 12306
rect 5908 12242 5960 12248
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 4816 11898 4844 12174
rect 4804 11892 4856 11898
rect 4804 11834 4856 11840
rect 5368 11694 5396 12242
rect 5920 11898 5948 12242
rect 5908 11892 5960 11898
rect 5908 11834 5960 11840
rect 5356 11688 5408 11694
rect 5356 11630 5408 11636
rect 6104 11150 6132 13262
rect 6196 12646 6224 13330
rect 6184 12640 6236 12646
rect 6184 12582 6236 12588
rect 6288 12458 6316 13330
rect 6380 12782 6408 13330
rect 6840 12986 6868 13806
rect 7114 13628 7422 13637
rect 7114 13626 7120 13628
rect 7176 13626 7200 13628
rect 7256 13626 7280 13628
rect 7336 13626 7360 13628
rect 7416 13626 7422 13628
rect 7176 13574 7178 13626
rect 7358 13574 7360 13626
rect 7114 13572 7120 13574
rect 7176 13572 7200 13574
rect 7256 13572 7280 13574
rect 7336 13572 7360 13574
rect 7416 13572 7422 13574
rect 7114 13563 7422 13572
rect 6920 13456 6972 13462
rect 6920 13398 6972 13404
rect 6828 12980 6880 12986
rect 6828 12922 6880 12928
rect 6368 12776 6420 12782
rect 6368 12718 6420 12724
rect 6552 12776 6604 12782
rect 6552 12718 6604 12724
rect 6564 12458 6592 12718
rect 6288 12430 6592 12458
rect 6564 11626 6592 12430
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 6552 11620 6604 11626
rect 6552 11562 6604 11568
rect 6656 11218 6684 11698
rect 6736 11688 6788 11694
rect 6736 11630 6788 11636
rect 6748 11354 6776 11630
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 6840 11218 6868 12922
rect 6932 11898 6960 13398
rect 7114 12540 7422 12549
rect 7114 12538 7120 12540
rect 7176 12538 7200 12540
rect 7256 12538 7280 12540
rect 7336 12538 7360 12540
rect 7416 12538 7422 12540
rect 7176 12486 7178 12538
rect 7358 12486 7360 12538
rect 7114 12484 7120 12486
rect 7176 12484 7200 12486
rect 7256 12484 7280 12486
rect 7336 12484 7360 12486
rect 7416 12484 7422 12486
rect 7114 12475 7422 12484
rect 7012 12164 7064 12170
rect 7012 12106 7064 12112
rect 6920 11892 6972 11898
rect 6920 11834 6972 11840
rect 6920 11552 6972 11558
rect 6920 11494 6972 11500
rect 6932 11354 6960 11494
rect 6920 11348 6972 11354
rect 6920 11290 6972 11296
rect 6644 11212 6696 11218
rect 6644 11154 6696 11160
rect 6828 11212 6880 11218
rect 6828 11154 6880 11160
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 6656 11098 6684 11154
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 6000 10600 6052 10606
rect 6104 10588 6132 11086
rect 6656 11070 6776 11098
rect 6184 11008 6236 11014
rect 6184 10950 6236 10956
rect 6196 10810 6224 10950
rect 6184 10804 6236 10810
rect 6184 10746 6236 10752
rect 6052 10560 6132 10588
rect 6644 10600 6696 10606
rect 6000 10542 6052 10548
rect 6748 10588 6776 11070
rect 6828 10600 6880 10606
rect 6748 10560 6828 10588
rect 6644 10542 6696 10548
rect 6828 10542 6880 10548
rect 4816 10266 4844 10542
rect 5080 10464 5132 10470
rect 5080 10406 5132 10412
rect 6276 10464 6328 10470
rect 6276 10406 6328 10412
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 4816 9518 4844 10202
rect 4896 10124 4948 10130
rect 4896 10066 4948 10072
rect 4908 9722 4936 10066
rect 4896 9716 4948 9722
rect 4896 9658 4948 9664
rect 5092 9518 5120 10406
rect 6288 10130 6316 10406
rect 6656 10266 6684 10542
rect 6644 10260 6696 10266
rect 6644 10202 6696 10208
rect 6276 10124 6328 10130
rect 6276 10066 6328 10072
rect 6840 10062 6868 10542
rect 6932 10130 6960 11290
rect 7024 11218 7052 12106
rect 7484 11898 7512 14350
rect 7564 12096 7616 12102
rect 7564 12038 7616 12044
rect 7472 11892 7524 11898
rect 7472 11834 7524 11840
rect 7576 11694 7604 12038
rect 7564 11688 7616 11694
rect 7564 11630 7616 11636
rect 7114 11452 7422 11461
rect 7114 11450 7120 11452
rect 7176 11450 7200 11452
rect 7256 11450 7280 11452
rect 7336 11450 7360 11452
rect 7416 11450 7422 11452
rect 7176 11398 7178 11450
rect 7358 11398 7360 11450
rect 7114 11396 7120 11398
rect 7176 11396 7200 11398
rect 7256 11396 7280 11398
rect 7336 11396 7360 11398
rect 7416 11396 7422 11398
rect 7114 11387 7422 11396
rect 7576 11218 7604 11630
rect 7012 11212 7064 11218
rect 7012 11154 7064 11160
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 7012 11076 7064 11082
rect 7012 11018 7064 11024
rect 7024 10674 7052 11018
rect 7012 10668 7064 10674
rect 7012 10610 7064 10616
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 4804 9512 4856 9518
rect 4804 9454 4856 9460
rect 5080 9512 5132 9518
rect 5080 9454 5132 9460
rect 6932 9450 6960 9862
rect 6920 9444 6972 9450
rect 6920 9386 6972 9392
rect 7024 8974 7052 10610
rect 7668 10538 7696 14418
rect 8128 13870 8156 15098
rect 8404 14958 8432 17070
rect 9508 16697 9536 18090
rect 9494 16688 9550 16697
rect 9494 16623 9550 16632
rect 9128 16584 9180 16590
rect 9128 16526 9180 16532
rect 9140 15502 9168 16526
rect 9312 16448 9364 16454
rect 9312 16390 9364 16396
rect 9324 15638 9352 16390
rect 9312 15632 9364 15638
rect 9312 15574 9364 15580
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 9220 15496 9272 15502
rect 9220 15438 9272 15444
rect 8484 15360 8536 15366
rect 8484 15302 8536 15308
rect 8760 15360 8812 15366
rect 8760 15302 8812 15308
rect 8392 14952 8444 14958
rect 8392 14894 8444 14900
rect 8208 14476 8260 14482
rect 8208 14418 8260 14424
rect 8116 13864 8168 13870
rect 8116 13806 8168 13812
rect 7932 13728 7984 13734
rect 7932 13670 7984 13676
rect 7748 12368 7800 12374
rect 7748 12310 7800 12316
rect 7656 10532 7708 10538
rect 7656 10474 7708 10480
rect 7472 10464 7524 10470
rect 7472 10406 7524 10412
rect 7114 10364 7422 10373
rect 7114 10362 7120 10364
rect 7176 10362 7200 10364
rect 7256 10362 7280 10364
rect 7336 10362 7360 10364
rect 7416 10362 7422 10364
rect 7176 10310 7178 10362
rect 7358 10310 7360 10362
rect 7114 10308 7120 10310
rect 7176 10308 7200 10310
rect 7256 10308 7280 10310
rect 7336 10308 7360 10310
rect 7416 10308 7422 10310
rect 7114 10299 7422 10308
rect 7484 10266 7512 10406
rect 7472 10260 7524 10266
rect 7472 10202 7524 10208
rect 7668 10198 7696 10474
rect 7656 10192 7708 10198
rect 7656 10134 7708 10140
rect 7564 9716 7616 9722
rect 7564 9658 7616 9664
rect 7472 9376 7524 9382
rect 7472 9318 7524 9324
rect 7114 9276 7422 9285
rect 7114 9274 7120 9276
rect 7176 9274 7200 9276
rect 7256 9274 7280 9276
rect 7336 9274 7360 9276
rect 7416 9274 7422 9276
rect 7176 9222 7178 9274
rect 7358 9222 7360 9274
rect 7114 9220 7120 9222
rect 7176 9220 7200 9222
rect 7256 9220 7280 9222
rect 7336 9220 7360 9222
rect 7416 9220 7422 9222
rect 7114 9211 7422 9220
rect 7484 9042 7512 9318
rect 7472 9036 7524 9042
rect 7472 8978 7524 8984
rect 7012 8968 7064 8974
rect 7012 8910 7064 8916
rect 5080 8628 5132 8634
rect 5080 8570 5132 8576
rect 4896 8424 4948 8430
rect 4896 8366 4948 8372
rect 4908 8022 4936 8366
rect 4896 8016 4948 8022
rect 4896 7958 4948 7964
rect 4896 7404 4948 7410
rect 4896 7346 4948 7352
rect 4804 7336 4856 7342
rect 4804 7278 4856 7284
rect 4712 7200 4764 7206
rect 4712 7142 4764 7148
rect 4816 6798 4844 7278
rect 4908 6866 4936 7346
rect 4988 7336 5040 7342
rect 4988 7278 5040 7284
rect 5000 6866 5028 7278
rect 5092 6866 5120 8570
rect 6552 8560 6604 8566
rect 6552 8502 6604 8508
rect 5816 8356 5868 8362
rect 5816 8298 5868 8304
rect 5828 7818 5856 8298
rect 6000 7948 6052 7954
rect 6000 7890 6052 7896
rect 5816 7812 5868 7818
rect 5816 7754 5868 7760
rect 6012 7546 6040 7890
rect 6276 7812 6328 7818
rect 6276 7754 6328 7760
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 6288 7410 6316 7754
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 6000 7336 6052 7342
rect 6000 7278 6052 7284
rect 6460 7336 6512 7342
rect 6460 7278 6512 7284
rect 5908 7200 5960 7206
rect 5908 7142 5960 7148
rect 5920 7002 5948 7142
rect 5908 6996 5960 7002
rect 5908 6938 5960 6944
rect 6012 6866 6040 7278
rect 6472 6866 6500 7278
rect 4896 6860 4948 6866
rect 4896 6802 4948 6808
rect 4988 6860 5040 6866
rect 4988 6802 5040 6808
rect 5080 6860 5132 6866
rect 5080 6802 5132 6808
rect 5264 6860 5316 6866
rect 5264 6802 5316 6808
rect 6000 6860 6052 6866
rect 6000 6802 6052 6808
rect 6460 6860 6512 6866
rect 6460 6802 6512 6808
rect 6564 6848 6592 8502
rect 6920 8424 6972 8430
rect 6920 8366 6972 8372
rect 6644 8016 6696 8022
rect 6644 7958 6696 7964
rect 6656 7546 6684 7958
rect 6932 7818 6960 8366
rect 7012 8288 7064 8294
rect 7012 8230 7064 8236
rect 7024 8022 7052 8230
rect 7114 8188 7422 8197
rect 7114 8186 7120 8188
rect 7176 8186 7200 8188
rect 7256 8186 7280 8188
rect 7336 8186 7360 8188
rect 7416 8186 7422 8188
rect 7176 8134 7178 8186
rect 7358 8134 7360 8186
rect 7114 8132 7120 8134
rect 7176 8132 7200 8134
rect 7256 8132 7280 8134
rect 7336 8132 7360 8134
rect 7416 8132 7422 8134
rect 7114 8123 7422 8132
rect 7012 8016 7064 8022
rect 7012 7958 7064 7964
rect 6920 7812 6972 7818
rect 6920 7754 6972 7760
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6644 6860 6696 6866
rect 6564 6820 6644 6848
rect 4620 6792 4672 6798
rect 4080 6718 4200 6746
rect 4620 6734 4672 6740
rect 4804 6792 4856 6798
rect 4804 6734 4856 6740
rect 3756 6556 4064 6565
rect 3756 6554 3762 6556
rect 3818 6554 3842 6556
rect 3898 6554 3922 6556
rect 3978 6554 4002 6556
rect 4058 6554 4064 6556
rect 3818 6502 3820 6554
rect 4000 6502 4002 6554
rect 3756 6500 3762 6502
rect 3818 6500 3842 6502
rect 3898 6500 3922 6502
rect 3978 6500 4002 6502
rect 4058 6500 4064 6502
rect 3756 6491 4064 6500
rect 4172 6440 4200 6718
rect 4632 6458 4660 6734
rect 4080 6412 4200 6440
rect 4620 6452 4672 6458
rect 3608 6384 3660 6390
rect 3608 6326 3660 6332
rect 3516 6248 3568 6254
rect 3516 6190 3568 6196
rect 3620 6186 3648 6326
rect 4080 6186 4108 6412
rect 4620 6394 4672 6400
rect 5092 6322 5120 6802
rect 5276 6390 5304 6802
rect 6012 6458 6040 6802
rect 6000 6452 6052 6458
rect 6000 6394 6052 6400
rect 5264 6384 5316 6390
rect 5264 6326 5316 6332
rect 5080 6316 5132 6322
rect 5080 6258 5132 6264
rect 4528 6248 4580 6254
rect 4528 6190 4580 6196
rect 4712 6248 4764 6254
rect 4896 6248 4948 6254
rect 4764 6196 4844 6202
rect 4712 6190 4844 6196
rect 4896 6190 4948 6196
rect 5632 6248 5684 6254
rect 5632 6190 5684 6196
rect 6184 6248 6236 6254
rect 6184 6190 6236 6196
rect 3608 6180 3660 6186
rect 3608 6122 3660 6128
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 3700 6112 3752 6118
rect 3700 6054 3752 6060
rect 3424 5908 3476 5914
rect 3424 5850 3476 5856
rect 3712 5846 3740 6054
rect 3700 5840 3752 5846
rect 3700 5782 3752 5788
rect 4540 5778 4568 6190
rect 4724 6174 4844 6190
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 4252 5772 4304 5778
rect 4252 5714 4304 5720
rect 4528 5772 4580 5778
rect 4528 5714 4580 5720
rect 3200 5528 3280 5556
rect 3148 5510 3200 5516
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 3068 5166 3096 5306
rect 3056 5160 3108 5166
rect 3056 5102 3108 5108
rect 2964 4820 3016 4826
rect 2964 4762 3016 4768
rect 3160 4690 3188 5510
rect 3756 5468 4064 5477
rect 3756 5466 3762 5468
rect 3818 5466 3842 5468
rect 3898 5466 3922 5468
rect 3978 5466 4002 5468
rect 4058 5466 4064 5468
rect 3818 5414 3820 5466
rect 4000 5414 4002 5466
rect 3756 5412 3762 5414
rect 3818 5412 3842 5414
rect 3898 5412 3922 5414
rect 3978 5412 4002 5414
rect 4058 5412 4064 5414
rect 3756 5403 4064 5412
rect 4172 5250 4200 5714
rect 4264 5370 4292 5714
rect 4252 5364 4304 5370
rect 4252 5306 4304 5312
rect 4816 5302 4844 6174
rect 4908 5914 4936 6190
rect 5644 5914 5672 6190
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 5632 5908 5684 5914
rect 5632 5850 5684 5856
rect 6196 5778 6224 6190
rect 6564 6186 6592 6820
rect 6644 6802 6696 6808
rect 6748 6798 6776 7278
rect 6840 7002 6868 7278
rect 6932 7002 6960 7346
rect 7012 7200 7064 7206
rect 7012 7142 7064 7148
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 7024 6934 7052 7142
rect 7114 7100 7422 7109
rect 7114 7098 7120 7100
rect 7176 7098 7200 7100
rect 7256 7098 7280 7100
rect 7336 7098 7360 7100
rect 7416 7098 7422 7100
rect 7176 7046 7178 7098
rect 7358 7046 7360 7098
rect 7114 7044 7120 7046
rect 7176 7044 7200 7046
rect 7256 7044 7280 7046
rect 7336 7044 7360 7046
rect 7416 7044 7422 7046
rect 7114 7035 7422 7044
rect 7012 6928 7064 6934
rect 7012 6870 7064 6876
rect 6828 6860 6880 6866
rect 6828 6802 6880 6808
rect 6736 6792 6788 6798
rect 6736 6734 6788 6740
rect 6840 6322 6868 6802
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 6552 6180 6604 6186
rect 6552 6122 6604 6128
rect 7012 6180 7064 6186
rect 7012 6122 7064 6128
rect 4896 5772 4948 5778
rect 4896 5714 4948 5720
rect 6184 5772 6236 5778
rect 6184 5714 6236 5720
rect 6276 5772 6328 5778
rect 6276 5714 6328 5720
rect 4804 5296 4856 5302
rect 4172 5222 4292 5250
rect 4804 5238 4856 5244
rect 4264 5098 4292 5222
rect 3332 5092 3384 5098
rect 3332 5034 3384 5040
rect 4252 5092 4304 5098
rect 4252 5034 4304 5040
rect 3344 4826 3372 5034
rect 3608 5024 3660 5030
rect 3608 4966 3660 4972
rect 3332 4820 3384 4826
rect 3332 4762 3384 4768
rect 3620 4758 3648 4966
rect 3608 4752 3660 4758
rect 3608 4694 3660 4700
rect 3148 4684 3200 4690
rect 3148 4626 3200 4632
rect 2964 4480 3016 4486
rect 2964 4422 3016 4428
rect 2976 4146 3004 4422
rect 3756 4380 4064 4389
rect 3756 4378 3762 4380
rect 3818 4378 3842 4380
rect 3898 4378 3922 4380
rect 3978 4378 4002 4380
rect 4058 4378 4064 4380
rect 3818 4326 3820 4378
rect 4000 4326 4002 4378
rect 3756 4324 3762 4326
rect 3818 4324 3842 4326
rect 3898 4324 3922 4326
rect 3978 4324 4002 4326
rect 4058 4324 4064 4326
rect 3756 4315 4064 4324
rect 4264 4282 4292 5034
rect 4908 4826 4936 5714
rect 6288 5370 6316 5714
rect 7024 5642 7052 6122
rect 7114 6012 7422 6021
rect 7114 6010 7120 6012
rect 7176 6010 7200 6012
rect 7256 6010 7280 6012
rect 7336 6010 7360 6012
rect 7416 6010 7422 6012
rect 7176 5958 7178 6010
rect 7358 5958 7360 6010
rect 7114 5956 7120 5958
rect 7176 5956 7200 5958
rect 7256 5956 7280 5958
rect 7336 5956 7360 5958
rect 7416 5956 7422 5958
rect 7114 5947 7422 5956
rect 7012 5636 7064 5642
rect 7012 5578 7064 5584
rect 7196 5636 7248 5642
rect 7196 5578 7248 5584
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 6460 5364 6512 5370
rect 6460 5306 6512 5312
rect 6092 5228 6144 5234
rect 6092 5170 6144 5176
rect 4988 5160 5040 5166
rect 4988 5102 5040 5108
rect 5264 5160 5316 5166
rect 5264 5102 5316 5108
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 5000 4826 5028 5102
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 4988 4820 5040 4826
rect 4988 4762 5040 4768
rect 4712 4684 4764 4690
rect 4712 4626 4764 4632
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 4252 4276 4304 4282
rect 4252 4218 4304 4224
rect 2964 4140 3016 4146
rect 2964 4082 3016 4088
rect 2872 4072 2924 4078
rect 2872 4014 2924 4020
rect 3424 4072 3476 4078
rect 3424 4014 3476 4020
rect 2320 3936 2372 3942
rect 2320 3878 2372 3884
rect 2884 3738 2912 4014
rect 3240 3936 3292 3942
rect 3436 3924 3464 4014
rect 4160 4004 4212 4010
rect 4160 3946 4212 3952
rect 3292 3896 3464 3924
rect 3240 3878 3292 3884
rect 2872 3732 2924 3738
rect 2872 3674 2924 3680
rect 4172 3602 4200 3946
rect 4252 3664 4304 3670
rect 4252 3606 4304 3612
rect 3608 3596 3660 3602
rect 3608 3538 3660 3544
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 4160 3596 4212 3602
rect 4160 3538 4212 3544
rect 3516 3460 3568 3466
rect 3516 3402 3568 3408
rect 3528 2990 3556 3402
rect 3620 3126 3648 3538
rect 4080 3380 4108 3538
rect 4080 3352 4200 3380
rect 3756 3292 4064 3301
rect 3756 3290 3762 3292
rect 3818 3290 3842 3292
rect 3898 3290 3922 3292
rect 3978 3290 4002 3292
rect 4058 3290 4064 3292
rect 3818 3238 3820 3290
rect 4000 3238 4002 3290
rect 3756 3236 3762 3238
rect 3818 3236 3842 3238
rect 3898 3236 3922 3238
rect 3978 3236 4002 3238
rect 4058 3236 4064 3238
rect 3756 3227 4064 3236
rect 3608 3120 3660 3126
rect 4172 3074 4200 3352
rect 4264 3194 4292 3606
rect 4724 3194 4752 4626
rect 4896 4208 4948 4214
rect 4896 4150 4948 4156
rect 4804 3392 4856 3398
rect 4804 3334 4856 3340
rect 4816 3194 4844 3334
rect 4252 3188 4304 3194
rect 4252 3130 4304 3136
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 3608 3062 3660 3068
rect 4080 3046 4200 3074
rect 4620 3120 4672 3126
rect 4908 3074 4936 4150
rect 5184 3738 5212 4626
rect 5276 4214 5304 5102
rect 5920 4826 5948 5102
rect 5908 4820 5960 4826
rect 5908 4762 5960 4768
rect 6000 4752 6052 4758
rect 6000 4694 6052 4700
rect 5264 4208 5316 4214
rect 5264 4150 5316 4156
rect 6012 3942 6040 4694
rect 6104 4486 6132 5170
rect 6184 5160 6236 5166
rect 6184 5102 6236 5108
rect 6196 5030 6224 5102
rect 6184 5024 6236 5030
rect 6184 4966 6236 4972
rect 6092 4480 6144 4486
rect 6092 4422 6144 4428
rect 6196 4078 6224 4966
rect 6472 4758 6500 5306
rect 6920 5296 6972 5302
rect 6920 5238 6972 5244
rect 6460 4752 6512 4758
rect 6460 4694 6512 4700
rect 6184 4072 6236 4078
rect 6184 4014 6236 4020
rect 6000 3936 6052 3942
rect 6000 3878 6052 3884
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 5356 3460 5408 3466
rect 5356 3402 5408 3408
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 4620 3062 4672 3068
rect 3148 2984 3200 2990
rect 3148 2926 3200 2932
rect 3516 2984 3568 2990
rect 3516 2926 3568 2932
rect 1216 2848 1268 2854
rect 1216 2790 1268 2796
rect 940 1896 992 1902
rect 940 1838 992 1844
rect 952 1018 980 1838
rect 1228 1426 1256 2790
rect 3160 2446 3188 2926
rect 3424 2508 3476 2514
rect 3424 2450 3476 2456
rect 3148 2440 3200 2446
rect 3148 2382 3200 2388
rect 3160 1902 3188 2382
rect 1768 1896 1820 1902
rect 1768 1838 1820 1844
rect 2136 1896 2188 1902
rect 2136 1838 2188 1844
rect 3148 1896 3200 1902
rect 3148 1838 3200 1844
rect 1216 1420 1268 1426
rect 1216 1362 1268 1368
rect 1308 1216 1360 1222
rect 1308 1158 1360 1164
rect 1320 1018 1348 1158
rect 940 1012 992 1018
rect 940 954 992 960
rect 1308 1012 1360 1018
rect 1308 954 1360 960
rect 1780 400 1808 1838
rect 2148 814 2176 1838
rect 2964 1760 3016 1766
rect 2964 1702 3016 1708
rect 2320 1488 2372 1494
rect 2320 1430 2372 1436
rect 2136 808 2188 814
rect 2136 750 2188 756
rect 2332 400 2360 1430
rect 2976 1426 3004 1702
rect 2964 1420 3016 1426
rect 2964 1362 3016 1368
rect 3240 1352 3292 1358
rect 3240 1294 3292 1300
rect 3332 1352 3384 1358
rect 3332 1294 3384 1300
rect 3252 950 3280 1294
rect 3344 1018 3372 1294
rect 3332 1012 3384 1018
rect 3332 954 3384 960
rect 3240 944 3292 950
rect 3240 886 3292 892
rect 2872 808 2924 814
rect 2872 750 2924 756
rect 2884 400 2912 750
rect 3436 400 3464 2450
rect 3528 1902 3556 2926
rect 4080 2514 4108 3046
rect 4068 2508 4120 2514
rect 4068 2450 4120 2456
rect 4528 2508 4580 2514
rect 4528 2450 4580 2456
rect 4080 2378 4108 2450
rect 4068 2372 4120 2378
rect 4068 2314 4120 2320
rect 4160 2304 4212 2310
rect 4160 2246 4212 2252
rect 3756 2204 4064 2213
rect 3756 2202 3762 2204
rect 3818 2202 3842 2204
rect 3898 2202 3922 2204
rect 3978 2202 4002 2204
rect 4058 2202 4064 2204
rect 3818 2150 3820 2202
rect 4000 2150 4002 2202
rect 3756 2148 3762 2150
rect 3818 2148 3842 2150
rect 3898 2148 3922 2150
rect 3978 2148 4002 2150
rect 4058 2148 4064 2150
rect 3756 2139 4064 2148
rect 3516 1896 3568 1902
rect 3516 1838 3568 1844
rect 3608 1760 3660 1766
rect 3608 1702 3660 1708
rect 3516 1488 3568 1494
rect 3516 1430 3568 1436
rect 1766 0 1822 400
rect 2318 0 2374 400
rect 2870 0 2926 400
rect 3422 0 3478 400
rect 3528 354 3556 1430
rect 3620 1426 3648 1702
rect 3608 1420 3660 1426
rect 3608 1362 3660 1368
rect 3756 1116 4064 1125
rect 3756 1114 3762 1116
rect 3818 1114 3842 1116
rect 3898 1114 3922 1116
rect 3978 1114 4002 1116
rect 4058 1114 4064 1116
rect 3818 1062 3820 1114
rect 4000 1062 4002 1114
rect 3756 1060 3762 1062
rect 3818 1060 3842 1062
rect 3898 1060 3922 1062
rect 3978 1060 4002 1062
rect 4058 1060 4064 1062
rect 3756 1051 4064 1060
rect 4172 882 4200 2246
rect 4540 1902 4568 2450
rect 4632 1902 4660 3062
rect 4724 3046 4936 3074
rect 4724 2514 4752 3046
rect 4804 2984 4856 2990
rect 4804 2926 4856 2932
rect 4988 2984 5040 2990
rect 4988 2926 5040 2932
rect 4816 2650 4844 2926
rect 4804 2644 4856 2650
rect 4804 2586 4856 2592
rect 4712 2508 4764 2514
rect 4712 2450 4764 2456
rect 4896 2508 4948 2514
rect 4896 2450 4948 2456
rect 4908 1986 4936 2450
rect 5000 2310 5028 2926
rect 4988 2304 5040 2310
rect 4988 2246 5040 2252
rect 4724 1970 4936 1986
rect 4712 1964 4936 1970
rect 4764 1958 4936 1964
rect 4712 1906 4764 1912
rect 4252 1896 4304 1902
rect 4252 1838 4304 1844
rect 4528 1896 4580 1902
rect 4528 1838 4580 1844
rect 4620 1896 4672 1902
rect 5184 1884 5212 3130
rect 5368 2990 5396 3402
rect 5264 2984 5316 2990
rect 5264 2926 5316 2932
rect 5356 2984 5408 2990
rect 5356 2926 5408 2932
rect 5276 2514 5304 2926
rect 5540 2916 5592 2922
rect 5540 2858 5592 2864
rect 5264 2508 5316 2514
rect 5264 2450 5316 2456
rect 5552 2310 5580 2858
rect 6012 2446 6040 3878
rect 6092 3596 6144 3602
rect 6092 3538 6144 3544
rect 6276 3596 6328 3602
rect 6276 3538 6328 3544
rect 6104 3126 6132 3538
rect 6092 3120 6144 3126
rect 6092 3062 6144 3068
rect 6104 2582 6132 3062
rect 6288 3058 6316 3538
rect 6276 3052 6328 3058
rect 6276 2994 6328 3000
rect 6472 2990 6500 4694
rect 6932 4554 6960 5238
rect 7208 5234 7236 5578
rect 7484 5574 7512 6190
rect 7472 5568 7524 5574
rect 7472 5510 7524 5516
rect 7196 5228 7248 5234
rect 7196 5170 7248 5176
rect 7484 5166 7512 5510
rect 7472 5160 7524 5166
rect 7472 5102 7524 5108
rect 7576 5098 7604 9658
rect 7760 9654 7788 12310
rect 7748 9648 7800 9654
rect 7748 9590 7800 9596
rect 7840 9512 7892 9518
rect 7840 9454 7892 9460
rect 7852 8906 7880 9454
rect 7944 8922 7972 13670
rect 8220 11694 8248 14418
rect 8404 13462 8432 14894
rect 8496 14890 8524 15302
rect 8484 14884 8536 14890
rect 8484 14826 8536 14832
rect 8772 14414 8800 15302
rect 8760 14408 8812 14414
rect 8760 14350 8812 14356
rect 9232 14346 9260 15438
rect 9508 14618 9536 16623
rect 9600 15960 9628 18090
rect 9680 15972 9732 15978
rect 9600 15932 9680 15960
rect 9600 14958 9628 15932
rect 9680 15914 9732 15920
rect 9588 14952 9640 14958
rect 9588 14894 9640 14900
rect 9588 14816 9640 14822
rect 9588 14758 9640 14764
rect 9496 14612 9548 14618
rect 9496 14554 9548 14560
rect 9600 14482 9628 14758
rect 9588 14476 9640 14482
rect 9588 14418 9640 14424
rect 9220 14340 9272 14346
rect 9220 14282 9272 14288
rect 8484 14000 8536 14006
rect 8484 13942 8536 13948
rect 8392 13456 8444 13462
rect 8392 13398 8444 13404
rect 8496 12434 8524 13942
rect 9968 13818 9996 21830
rect 10046 21040 10102 21049
rect 10046 20975 10102 20984
rect 10060 19854 10088 20975
rect 10152 20942 10180 21966
rect 10336 21894 10364 23038
rect 10472 22876 10780 22885
rect 10472 22874 10478 22876
rect 10534 22874 10558 22876
rect 10614 22874 10638 22876
rect 10694 22874 10718 22876
rect 10774 22874 10780 22876
rect 10534 22822 10536 22874
rect 10716 22822 10718 22874
rect 10472 22820 10478 22822
rect 10534 22820 10558 22822
rect 10614 22820 10638 22822
rect 10694 22820 10718 22822
rect 10774 22820 10780 22822
rect 10472 22811 10780 22820
rect 10416 22432 10468 22438
rect 10416 22374 10468 22380
rect 10428 22098 10456 22374
rect 10416 22092 10468 22098
rect 10416 22034 10468 22040
rect 10324 21888 10376 21894
rect 10324 21830 10376 21836
rect 10472 21788 10780 21797
rect 10472 21786 10478 21788
rect 10534 21786 10558 21788
rect 10614 21786 10638 21788
rect 10694 21786 10718 21788
rect 10774 21786 10780 21788
rect 10534 21734 10536 21786
rect 10716 21734 10718 21786
rect 10472 21732 10478 21734
rect 10534 21732 10558 21734
rect 10614 21732 10638 21734
rect 10694 21732 10718 21734
rect 10774 21732 10780 21734
rect 10472 21723 10780 21732
rect 10140 20936 10192 20942
rect 10140 20878 10192 20884
rect 10048 19848 10100 19854
rect 10048 19790 10100 19796
rect 10046 17912 10102 17921
rect 10046 17847 10048 17856
rect 10100 17847 10102 17856
rect 10048 17818 10100 17824
rect 10152 17762 10180 20878
rect 10232 20800 10284 20806
rect 10232 20742 10284 20748
rect 10244 20398 10272 20742
rect 10472 20700 10780 20709
rect 10472 20698 10478 20700
rect 10534 20698 10558 20700
rect 10614 20698 10638 20700
rect 10694 20698 10718 20700
rect 10774 20698 10780 20700
rect 10534 20646 10536 20698
rect 10716 20646 10718 20698
rect 10472 20644 10478 20646
rect 10534 20644 10558 20646
rect 10614 20644 10638 20646
rect 10694 20644 10718 20646
rect 10774 20644 10780 20646
rect 10472 20635 10780 20644
rect 10232 20392 10284 20398
rect 10232 20334 10284 20340
rect 10980 20058 11008 24074
rect 11164 23662 11192 24210
rect 11152 23656 11204 23662
rect 11152 23598 11204 23604
rect 11336 23656 11388 23662
rect 11336 23598 11388 23604
rect 11348 23050 11376 23598
rect 11440 23118 11468 26318
rect 11716 26042 11744 26454
rect 12072 26444 12124 26450
rect 12072 26386 12124 26392
rect 11888 26240 11940 26246
rect 11888 26182 11940 26188
rect 11704 26036 11756 26042
rect 11704 25978 11756 25984
rect 11900 25430 11928 26182
rect 12084 25498 12112 26386
rect 12072 25492 12124 25498
rect 12072 25434 12124 25440
rect 11888 25424 11940 25430
rect 11888 25366 11940 25372
rect 11704 24132 11756 24138
rect 11704 24074 11756 24080
rect 11428 23112 11480 23118
rect 11428 23054 11480 23060
rect 11520 23112 11572 23118
rect 11520 23054 11572 23060
rect 11336 23044 11388 23050
rect 11336 22986 11388 22992
rect 11348 22760 11376 22986
rect 11348 22732 11468 22760
rect 11336 22636 11388 22642
rect 11336 22578 11388 22584
rect 11244 22432 11296 22438
rect 11244 22374 11296 22380
rect 11256 22137 11284 22374
rect 11242 22128 11298 22137
rect 11348 22098 11376 22578
rect 11242 22063 11298 22072
rect 11336 22092 11388 22098
rect 11336 22034 11388 22040
rect 11058 21992 11114 22001
rect 11058 21927 11114 21936
rect 11072 21418 11100 21927
rect 11244 21888 11296 21894
rect 11244 21830 11296 21836
rect 11256 21486 11284 21830
rect 11348 21690 11376 22034
rect 11336 21684 11388 21690
rect 11336 21626 11388 21632
rect 11440 21486 11468 22732
rect 11532 22642 11560 23054
rect 11716 22982 11744 24074
rect 11796 23588 11848 23594
rect 11796 23530 11848 23536
rect 11888 23588 11940 23594
rect 11888 23530 11940 23536
rect 11808 23254 11836 23530
rect 11796 23248 11848 23254
rect 11796 23190 11848 23196
rect 11900 23186 11928 23530
rect 12072 23520 12124 23526
rect 12072 23462 12124 23468
rect 12084 23186 12112 23462
rect 11888 23180 11940 23186
rect 11888 23122 11940 23128
rect 12072 23180 12124 23186
rect 12072 23122 12124 23128
rect 12176 23066 12204 28970
rect 11992 23038 12204 23066
rect 11704 22976 11756 22982
rect 11704 22918 11756 22924
rect 11796 22976 11848 22982
rect 11796 22918 11848 22924
rect 11520 22636 11572 22642
rect 11520 22578 11572 22584
rect 11532 22094 11560 22578
rect 11808 22506 11836 22918
rect 11888 22568 11940 22574
rect 11888 22510 11940 22516
rect 11796 22500 11848 22506
rect 11796 22442 11848 22448
rect 11532 22066 11744 22094
rect 11520 21616 11572 21622
rect 11520 21558 11572 21564
rect 11244 21480 11296 21486
rect 11244 21422 11296 21428
rect 11428 21480 11480 21486
rect 11428 21422 11480 21428
rect 11060 21412 11112 21418
rect 11060 21354 11112 21360
rect 11532 21332 11560 21558
rect 11440 21304 11560 21332
rect 11440 21010 11468 21304
rect 11428 21004 11480 21010
rect 11428 20946 11480 20952
rect 11336 20936 11388 20942
rect 11336 20878 11388 20884
rect 11348 20602 11376 20878
rect 11336 20596 11388 20602
rect 11336 20538 11388 20544
rect 10968 20052 11020 20058
rect 11440 20040 11468 20946
rect 11716 20942 11744 22066
rect 11796 22092 11848 22098
rect 11796 22034 11848 22040
rect 11808 21554 11836 22034
rect 11796 21548 11848 21554
rect 11796 21490 11848 21496
rect 11900 21418 11928 22510
rect 11888 21412 11940 21418
rect 11888 21354 11940 21360
rect 11900 21078 11928 21354
rect 11888 21072 11940 21078
rect 11888 21014 11940 21020
rect 11704 20936 11756 20942
rect 11704 20878 11756 20884
rect 11992 20505 12020 23038
rect 12268 22642 12296 29446
rect 12544 29238 12572 29582
rect 12532 29232 12584 29238
rect 12532 29174 12584 29180
rect 12348 29164 12400 29170
rect 12348 29106 12400 29112
rect 12360 23186 12388 29106
rect 12440 26444 12492 26450
rect 12440 26386 12492 26392
rect 12452 23526 12480 26386
rect 12636 25906 12664 29582
rect 13084 29028 13136 29034
rect 13084 28970 13136 28976
rect 12992 28620 13044 28626
rect 12992 28562 13044 28568
rect 13004 28218 13032 28562
rect 12992 28212 13044 28218
rect 12992 28154 13044 28160
rect 13096 28014 13124 28970
rect 13084 28008 13136 28014
rect 13084 27950 13136 27956
rect 12716 27872 12768 27878
rect 12716 27814 12768 27820
rect 12728 27606 12756 27814
rect 12716 27600 12768 27606
rect 12716 27542 12768 27548
rect 12992 27328 13044 27334
rect 12992 27270 13044 27276
rect 12808 26988 12860 26994
rect 12808 26930 12860 26936
rect 12716 26784 12768 26790
rect 12716 26726 12768 26732
rect 12728 26450 12756 26726
rect 12716 26444 12768 26450
rect 12716 26386 12768 26392
rect 12624 25900 12676 25906
rect 12624 25842 12676 25848
rect 12820 25838 12848 26930
rect 13004 26926 13032 27270
rect 12900 26920 12952 26926
rect 12900 26862 12952 26868
rect 12992 26920 13044 26926
rect 12992 26862 13044 26868
rect 12808 25832 12860 25838
rect 12808 25774 12860 25780
rect 12820 25242 12848 25774
rect 12728 25214 12848 25242
rect 12728 25158 12756 25214
rect 12716 25152 12768 25158
rect 12716 25094 12768 25100
rect 12624 24676 12676 24682
rect 12624 24618 12676 24624
rect 12636 24410 12664 24618
rect 12624 24404 12676 24410
rect 12624 24346 12676 24352
rect 12716 24404 12768 24410
rect 12716 24346 12768 24352
rect 12530 23624 12586 23633
rect 12530 23559 12586 23568
rect 12440 23520 12492 23526
rect 12440 23462 12492 23468
rect 12544 23254 12572 23559
rect 12728 23322 12756 24346
rect 12912 23866 12940 26862
rect 12992 26784 13044 26790
rect 12992 26726 13044 26732
rect 13004 26450 13032 26726
rect 12992 26444 13044 26450
rect 12992 26386 13044 26392
rect 12992 25696 13044 25702
rect 12992 25638 13044 25644
rect 13004 25430 13032 25638
rect 12992 25424 13044 25430
rect 12992 25366 13044 25372
rect 13188 24392 13216 29990
rect 13556 29782 13584 29990
rect 13544 29776 13596 29782
rect 13544 29718 13596 29724
rect 13360 29504 13412 29510
rect 13360 29446 13412 29452
rect 13372 29102 13400 29446
rect 13648 29170 13676 30534
rect 13728 30184 13780 30190
rect 13728 30126 13780 30132
rect 13636 29164 13688 29170
rect 13636 29106 13688 29112
rect 13360 29096 13412 29102
rect 13360 29038 13412 29044
rect 13268 28960 13320 28966
rect 13268 28902 13320 28908
rect 13280 28422 13308 28902
rect 13268 28416 13320 28422
rect 13268 28358 13320 28364
rect 13372 28218 13400 29038
rect 13740 28762 13768 30126
rect 14016 30122 14044 30534
rect 14004 30116 14056 30122
rect 14004 30058 14056 30064
rect 13830 29948 14138 29957
rect 13830 29946 13836 29948
rect 13892 29946 13916 29948
rect 13972 29946 13996 29948
rect 14052 29946 14076 29948
rect 14132 29946 14138 29948
rect 13892 29894 13894 29946
rect 14074 29894 14076 29946
rect 13830 29892 13836 29894
rect 13892 29892 13916 29894
rect 13972 29892 13996 29894
rect 14052 29892 14076 29894
rect 14132 29892 14138 29894
rect 13830 29883 14138 29892
rect 13830 28860 14138 28869
rect 13830 28858 13836 28860
rect 13892 28858 13916 28860
rect 13972 28858 13996 28860
rect 14052 28858 14076 28860
rect 14132 28858 14138 28860
rect 13892 28806 13894 28858
rect 14074 28806 14076 28858
rect 13830 28804 13836 28806
rect 13892 28804 13916 28806
rect 13972 28804 13996 28806
rect 14052 28804 14076 28806
rect 14132 28804 14138 28806
rect 13830 28795 14138 28804
rect 13728 28756 13780 28762
rect 13728 28698 13780 28704
rect 13912 28552 13964 28558
rect 13912 28494 13964 28500
rect 13924 28218 13952 28494
rect 13360 28212 13412 28218
rect 13360 28154 13412 28160
rect 13912 28212 13964 28218
rect 13912 28154 13964 28160
rect 13372 27538 13400 28154
rect 13636 27940 13688 27946
rect 13636 27882 13688 27888
rect 13648 27538 13676 27882
rect 13830 27772 14138 27781
rect 13830 27770 13836 27772
rect 13892 27770 13916 27772
rect 13972 27770 13996 27772
rect 14052 27770 14076 27772
rect 14132 27770 14138 27772
rect 13892 27718 13894 27770
rect 14074 27718 14076 27770
rect 13830 27716 13836 27718
rect 13892 27716 13916 27718
rect 13972 27716 13996 27718
rect 14052 27716 14076 27718
rect 14132 27716 14138 27718
rect 13830 27707 14138 27716
rect 13360 27532 13412 27538
rect 13360 27474 13412 27480
rect 13636 27532 13688 27538
rect 13636 27474 13688 27480
rect 13820 27328 13872 27334
rect 13820 27270 13872 27276
rect 13832 26926 13860 27270
rect 13820 26920 13872 26926
rect 13820 26862 13872 26868
rect 13360 26852 13412 26858
rect 13360 26794 13412 26800
rect 13372 24818 13400 26794
rect 13830 26684 14138 26693
rect 13830 26682 13836 26684
rect 13892 26682 13916 26684
rect 13972 26682 13996 26684
rect 14052 26682 14076 26684
rect 14132 26682 14138 26684
rect 13892 26630 13894 26682
rect 14074 26630 14076 26682
rect 13830 26628 13836 26630
rect 13892 26628 13916 26630
rect 13972 26628 13996 26630
rect 14052 26628 14076 26630
rect 14132 26628 14138 26630
rect 13830 26619 14138 26628
rect 14200 26489 14228 30738
rect 17788 30598 17816 30738
rect 14740 30592 14792 30598
rect 14740 30534 14792 30540
rect 16764 30592 16816 30598
rect 16764 30534 16816 30540
rect 17592 30592 17644 30598
rect 17776 30592 17828 30598
rect 17592 30534 17644 30540
rect 17696 30552 17776 30580
rect 14556 30048 14608 30054
rect 14556 29990 14608 29996
rect 14568 29850 14596 29990
rect 14556 29844 14608 29850
rect 14556 29786 14608 29792
rect 14568 29714 14596 29786
rect 14556 29708 14608 29714
rect 14556 29650 14608 29656
rect 14752 29170 14780 30534
rect 16028 30320 16080 30326
rect 16028 30262 16080 30268
rect 15384 30184 15436 30190
rect 15384 30126 15436 30132
rect 15396 29850 15424 30126
rect 15108 29844 15160 29850
rect 15108 29786 15160 29792
rect 15384 29844 15436 29850
rect 15384 29786 15436 29792
rect 14740 29164 14792 29170
rect 14740 29106 14792 29112
rect 14648 28620 14700 28626
rect 14648 28562 14700 28568
rect 14280 28416 14332 28422
rect 14280 28358 14332 28364
rect 14292 27538 14320 28358
rect 14660 28218 14688 28562
rect 14648 28212 14700 28218
rect 14648 28154 14700 28160
rect 14464 27940 14516 27946
rect 14464 27882 14516 27888
rect 14476 27674 14504 27882
rect 14464 27668 14516 27674
rect 14464 27610 14516 27616
rect 14280 27532 14332 27538
rect 14280 27474 14332 27480
rect 14280 26920 14332 26926
rect 14280 26862 14332 26868
rect 14292 26586 14320 26862
rect 14280 26580 14332 26586
rect 14280 26522 14332 26528
rect 14186 26480 14242 26489
rect 14752 26450 14780 29106
rect 15120 28422 15148 29786
rect 15200 29776 15252 29782
rect 15252 29724 15424 29730
rect 15200 29718 15424 29724
rect 15212 29702 15424 29718
rect 15396 29646 15424 29702
rect 15200 29640 15252 29646
rect 15200 29582 15252 29588
rect 15384 29640 15436 29646
rect 15384 29582 15436 29588
rect 15212 28762 15240 29582
rect 15292 29572 15344 29578
rect 15292 29514 15344 29520
rect 15304 29102 15332 29514
rect 15292 29096 15344 29102
rect 15292 29038 15344 29044
rect 15200 28756 15252 28762
rect 15200 28698 15252 28704
rect 15212 28558 15240 28698
rect 15396 28558 15424 29582
rect 15660 29504 15712 29510
rect 15660 29446 15712 29452
rect 15672 29306 15700 29446
rect 15660 29300 15712 29306
rect 15660 29242 15712 29248
rect 16040 29102 16068 30262
rect 16120 30184 16172 30190
rect 16120 30126 16172 30132
rect 16132 29850 16160 30126
rect 16120 29844 16172 29850
rect 16120 29786 16172 29792
rect 16776 29782 16804 30534
rect 17188 30492 17496 30501
rect 17188 30490 17194 30492
rect 17250 30490 17274 30492
rect 17330 30490 17354 30492
rect 17410 30490 17434 30492
rect 17490 30490 17496 30492
rect 17250 30438 17252 30490
rect 17432 30438 17434 30490
rect 17188 30436 17194 30438
rect 17250 30436 17274 30438
rect 17330 30436 17354 30438
rect 17410 30436 17434 30438
rect 17490 30436 17496 30438
rect 17188 30427 17496 30436
rect 16856 30116 16908 30122
rect 16856 30058 16908 30064
rect 16764 29776 16816 29782
rect 16764 29718 16816 29724
rect 16868 29578 16896 30058
rect 17604 29714 17632 30534
rect 17592 29708 17644 29714
rect 17592 29650 17644 29656
rect 16580 29572 16632 29578
rect 16580 29514 16632 29520
rect 16856 29572 16908 29578
rect 16856 29514 16908 29520
rect 16592 29102 16620 29514
rect 16672 29300 16724 29306
rect 16672 29242 16724 29248
rect 15476 29096 15528 29102
rect 15476 29038 15528 29044
rect 16028 29096 16080 29102
rect 16028 29038 16080 29044
rect 16580 29096 16632 29102
rect 16580 29038 16632 29044
rect 15488 28626 15516 29038
rect 15844 29028 15896 29034
rect 15844 28970 15896 28976
rect 15856 28694 15884 28970
rect 16304 28960 16356 28966
rect 16304 28902 16356 28908
rect 16316 28762 16344 28902
rect 16304 28756 16356 28762
rect 16304 28698 16356 28704
rect 16592 28694 16620 29038
rect 16684 29034 16712 29242
rect 16764 29096 16816 29102
rect 16764 29038 16816 29044
rect 16672 29028 16724 29034
rect 16672 28970 16724 28976
rect 15844 28688 15896 28694
rect 15844 28630 15896 28636
rect 16580 28688 16632 28694
rect 16580 28630 16632 28636
rect 15476 28620 15528 28626
rect 15476 28562 15528 28568
rect 15752 28620 15804 28626
rect 15752 28562 15804 28568
rect 15200 28552 15252 28558
rect 15200 28494 15252 28500
rect 15384 28552 15436 28558
rect 15384 28494 15436 28500
rect 15108 28416 15160 28422
rect 15108 28358 15160 28364
rect 15120 27538 15148 28358
rect 15488 27538 15516 28562
rect 15660 28008 15712 28014
rect 15660 27950 15712 27956
rect 15672 27674 15700 27950
rect 15660 27668 15712 27674
rect 15660 27610 15712 27616
rect 15108 27532 15160 27538
rect 15108 27474 15160 27480
rect 15476 27532 15528 27538
rect 15476 27474 15528 27480
rect 14924 27328 14976 27334
rect 14924 27270 14976 27276
rect 15660 27328 15712 27334
rect 15660 27270 15712 27276
rect 14936 26926 14964 27270
rect 15568 27056 15620 27062
rect 15568 26998 15620 27004
rect 15580 26926 15608 26998
rect 15672 26926 15700 27270
rect 14832 26920 14884 26926
rect 14832 26862 14884 26868
rect 14924 26920 14976 26926
rect 14924 26862 14976 26868
rect 15568 26920 15620 26926
rect 15568 26862 15620 26868
rect 15660 26920 15712 26926
rect 15660 26862 15712 26868
rect 14186 26415 14242 26424
rect 14740 26444 14792 26450
rect 13636 25764 13688 25770
rect 13636 25706 13688 25712
rect 13648 25498 13676 25706
rect 13830 25596 14138 25605
rect 13830 25594 13836 25596
rect 13892 25594 13916 25596
rect 13972 25594 13996 25596
rect 14052 25594 14076 25596
rect 14132 25594 14138 25596
rect 13892 25542 13894 25594
rect 14074 25542 14076 25594
rect 13830 25540 13836 25542
rect 13892 25540 13916 25542
rect 13972 25540 13996 25542
rect 14052 25540 14076 25542
rect 14132 25540 14138 25542
rect 13830 25531 14138 25540
rect 13636 25492 13688 25498
rect 13636 25434 13688 25440
rect 14004 25356 14056 25362
rect 14004 25298 14056 25304
rect 13360 24812 13412 24818
rect 13360 24754 13412 24760
rect 13372 24614 13400 24754
rect 14016 24750 14044 25298
rect 14004 24744 14056 24750
rect 14004 24686 14056 24692
rect 13360 24608 13412 24614
rect 13360 24550 13412 24556
rect 13452 24608 13504 24614
rect 13452 24550 13504 24556
rect 13188 24364 13308 24392
rect 13084 24268 13136 24274
rect 13084 24210 13136 24216
rect 12992 24064 13044 24070
rect 12992 24006 13044 24012
rect 12900 23860 12952 23866
rect 12900 23802 12952 23808
rect 12808 23656 12860 23662
rect 12808 23598 12860 23604
rect 12716 23316 12768 23322
rect 12716 23258 12768 23264
rect 12532 23248 12584 23254
rect 12532 23190 12584 23196
rect 12348 23180 12400 23186
rect 12348 23122 12400 23128
rect 12348 23044 12400 23050
rect 12348 22986 12400 22992
rect 12256 22636 12308 22642
rect 12256 22578 12308 22584
rect 12268 22098 12296 22578
rect 12360 22166 12388 22986
rect 12348 22160 12400 22166
rect 12348 22102 12400 22108
rect 12256 22092 12308 22098
rect 12176 22052 12256 22080
rect 12072 21548 12124 21554
rect 12072 21490 12124 21496
rect 12084 20806 12112 21490
rect 12176 21486 12204 22052
rect 12256 22034 12308 22040
rect 12348 22024 12400 22030
rect 12348 21966 12400 21972
rect 12256 21888 12308 21894
rect 12256 21830 12308 21836
rect 12164 21480 12216 21486
rect 12164 21422 12216 21428
rect 12176 21078 12204 21422
rect 12164 21072 12216 21078
rect 12164 21014 12216 21020
rect 12072 20800 12124 20806
rect 12072 20742 12124 20748
rect 11978 20496 12034 20505
rect 11978 20431 12034 20440
rect 10968 19994 11020 20000
rect 11348 20012 11468 20040
rect 10876 19848 10928 19854
rect 10876 19790 10928 19796
rect 10472 19612 10780 19621
rect 10472 19610 10478 19612
rect 10534 19610 10558 19612
rect 10614 19610 10638 19612
rect 10694 19610 10718 19612
rect 10774 19610 10780 19612
rect 10534 19558 10536 19610
rect 10716 19558 10718 19610
rect 10472 19556 10478 19558
rect 10534 19556 10558 19558
rect 10614 19556 10638 19558
rect 10694 19556 10718 19558
rect 10774 19556 10780 19558
rect 10472 19547 10780 19556
rect 10472 18524 10780 18533
rect 10472 18522 10478 18524
rect 10534 18522 10558 18524
rect 10614 18522 10638 18524
rect 10694 18522 10718 18524
rect 10774 18522 10780 18524
rect 10534 18470 10536 18522
rect 10716 18470 10718 18522
rect 10472 18468 10478 18470
rect 10534 18468 10558 18470
rect 10614 18468 10638 18470
rect 10694 18468 10718 18470
rect 10774 18468 10780 18470
rect 10472 18459 10780 18468
rect 10060 17734 10180 17762
rect 10232 17740 10284 17746
rect 10060 14006 10088 17734
rect 10232 17682 10284 17688
rect 10140 16992 10192 16998
rect 10140 16934 10192 16940
rect 10152 16794 10180 16934
rect 10244 16794 10272 17682
rect 10472 17436 10780 17445
rect 10472 17434 10478 17436
rect 10534 17434 10558 17436
rect 10614 17434 10638 17436
rect 10694 17434 10718 17436
rect 10774 17434 10780 17436
rect 10534 17382 10536 17434
rect 10716 17382 10718 17434
rect 10472 17380 10478 17382
rect 10534 17380 10558 17382
rect 10614 17380 10638 17382
rect 10694 17380 10718 17382
rect 10774 17380 10780 17382
rect 10472 17371 10780 17380
rect 10324 16992 10376 16998
rect 10324 16934 10376 16940
rect 10692 16992 10744 16998
rect 10692 16934 10744 16940
rect 10140 16788 10192 16794
rect 10140 16730 10192 16736
rect 10232 16788 10284 16794
rect 10232 16730 10284 16736
rect 10336 16658 10364 16934
rect 10704 16726 10732 16934
rect 10692 16720 10744 16726
rect 10692 16662 10744 16668
rect 10324 16652 10376 16658
rect 10324 16594 10376 16600
rect 10336 15706 10364 16594
rect 10472 16348 10780 16357
rect 10472 16346 10478 16348
rect 10534 16346 10558 16348
rect 10614 16346 10638 16348
rect 10694 16346 10718 16348
rect 10774 16346 10780 16348
rect 10534 16294 10536 16346
rect 10716 16294 10718 16346
rect 10472 16292 10478 16294
rect 10534 16292 10558 16294
rect 10614 16292 10638 16294
rect 10694 16292 10718 16294
rect 10774 16292 10780 16294
rect 10472 16283 10780 16292
rect 10324 15700 10376 15706
rect 10324 15642 10376 15648
rect 10472 15260 10780 15269
rect 10472 15258 10478 15260
rect 10534 15258 10558 15260
rect 10614 15258 10638 15260
rect 10694 15258 10718 15260
rect 10774 15258 10780 15260
rect 10534 15206 10536 15258
rect 10716 15206 10718 15258
rect 10472 15204 10478 15206
rect 10534 15204 10558 15206
rect 10614 15204 10638 15206
rect 10694 15204 10718 15206
rect 10774 15204 10780 15206
rect 10472 15195 10780 15204
rect 10472 14172 10780 14181
rect 10472 14170 10478 14172
rect 10534 14170 10558 14172
rect 10614 14170 10638 14172
rect 10694 14170 10718 14172
rect 10774 14170 10780 14172
rect 10534 14118 10536 14170
rect 10716 14118 10718 14170
rect 10472 14116 10478 14118
rect 10534 14116 10558 14118
rect 10614 14116 10638 14118
rect 10694 14116 10718 14118
rect 10774 14116 10780 14118
rect 10472 14107 10780 14116
rect 10888 14074 10916 19790
rect 11060 19236 11112 19242
rect 11060 19178 11112 19184
rect 11072 18970 11100 19178
rect 11060 18964 11112 18970
rect 11060 18906 11112 18912
rect 11060 18760 11112 18766
rect 11060 18702 11112 18708
rect 11072 18630 11100 18702
rect 11060 18624 11112 18630
rect 11060 18566 11112 18572
rect 10968 18148 11020 18154
rect 10968 18090 11020 18096
rect 10980 17882 11008 18090
rect 10968 17876 11020 17882
rect 10968 17818 11020 17824
rect 11072 17134 11100 18566
rect 11244 18216 11296 18222
rect 11244 18158 11296 18164
rect 11152 18148 11204 18154
rect 11152 18090 11204 18096
rect 11164 17746 11192 18090
rect 11152 17740 11204 17746
rect 11152 17682 11204 17688
rect 11256 17626 11284 18158
rect 11164 17610 11284 17626
rect 11152 17604 11284 17610
rect 11204 17598 11284 17604
rect 11152 17546 11204 17552
rect 11060 17128 11112 17134
rect 11060 17070 11112 17076
rect 11164 16590 11192 17546
rect 11348 16794 11376 20012
rect 11428 19916 11480 19922
rect 11428 19858 11480 19864
rect 11440 18834 11468 19858
rect 12072 19780 12124 19786
rect 12072 19722 12124 19728
rect 11704 19712 11756 19718
rect 11704 19654 11756 19660
rect 11520 19304 11572 19310
rect 11520 19246 11572 19252
rect 11532 18902 11560 19246
rect 11520 18896 11572 18902
rect 11520 18838 11572 18844
rect 11716 18834 11744 19654
rect 11428 18828 11480 18834
rect 11428 18770 11480 18776
rect 11704 18828 11756 18834
rect 11704 18770 11756 18776
rect 11612 18692 11664 18698
rect 11612 18634 11664 18640
rect 11428 18080 11480 18086
rect 11428 18022 11480 18028
rect 11440 17746 11468 18022
rect 11428 17740 11480 17746
rect 11428 17682 11480 17688
rect 11520 17740 11572 17746
rect 11624 17728 11652 18634
rect 12084 18222 12112 19722
rect 12268 19394 12296 21830
rect 12360 21418 12388 21966
rect 12348 21412 12400 21418
rect 12348 21354 12400 21360
rect 12544 21350 12572 23190
rect 12820 22438 12848 23598
rect 12900 23180 12952 23186
rect 12900 23122 12952 23128
rect 12912 22642 12940 23122
rect 13004 23066 13032 24006
rect 13096 23526 13124 24210
rect 13280 23633 13308 24364
rect 13464 24342 13492 24550
rect 13830 24508 14138 24517
rect 13830 24506 13836 24508
rect 13892 24506 13916 24508
rect 13972 24506 13996 24508
rect 14052 24506 14076 24508
rect 14132 24506 14138 24508
rect 13892 24454 13894 24506
rect 14074 24454 14076 24506
rect 13830 24452 13836 24454
rect 13892 24452 13916 24454
rect 13972 24452 13996 24454
rect 14052 24452 14076 24454
rect 14132 24452 14138 24454
rect 13830 24443 14138 24452
rect 14200 24410 14228 26415
rect 14740 26386 14792 26392
rect 14844 26042 14872 26862
rect 15382 26344 15438 26353
rect 15382 26279 15438 26288
rect 14832 26036 14884 26042
rect 14832 25978 14884 25984
rect 14844 25906 14872 25978
rect 14832 25900 14884 25906
rect 14832 25842 14884 25848
rect 15016 25696 15068 25702
rect 15016 25638 15068 25644
rect 15028 25498 15056 25638
rect 15016 25492 15068 25498
rect 15016 25434 15068 25440
rect 14924 25356 14976 25362
rect 14924 25298 14976 25304
rect 14556 24948 14608 24954
rect 14556 24890 14608 24896
rect 14464 24744 14516 24750
rect 14464 24686 14516 24692
rect 14188 24404 14240 24410
rect 14188 24346 14240 24352
rect 13452 24336 13504 24342
rect 13452 24278 13504 24284
rect 13728 24064 13780 24070
rect 13728 24006 13780 24012
rect 13740 23866 13768 24006
rect 13728 23860 13780 23866
rect 13728 23802 13780 23808
rect 14188 23792 14240 23798
rect 14188 23734 14240 23740
rect 13360 23656 13412 23662
rect 13266 23624 13322 23633
rect 13360 23598 13412 23604
rect 13266 23559 13322 23568
rect 13084 23520 13136 23526
rect 13084 23462 13136 23468
rect 13004 23038 13124 23066
rect 12992 22976 13044 22982
rect 12992 22918 13044 22924
rect 13004 22710 13032 22918
rect 12992 22704 13044 22710
rect 12992 22646 13044 22652
rect 12900 22636 12952 22642
rect 12900 22578 12952 22584
rect 12808 22432 12860 22438
rect 12808 22374 12860 22380
rect 12912 22094 12940 22578
rect 12992 22568 13044 22574
rect 12992 22510 13044 22516
rect 12728 22066 12940 22094
rect 12532 21344 12584 21350
rect 12532 21286 12584 21292
rect 12440 20800 12492 20806
rect 12440 20742 12492 20748
rect 12452 19990 12480 20742
rect 12624 20256 12676 20262
rect 12624 20198 12676 20204
rect 12532 20052 12584 20058
rect 12532 19994 12584 20000
rect 12440 19984 12492 19990
rect 12440 19926 12492 19932
rect 12348 19916 12400 19922
rect 12348 19858 12400 19864
rect 12176 19366 12296 19394
rect 12072 18216 12124 18222
rect 12072 18158 12124 18164
rect 12072 18080 12124 18086
rect 12072 18022 12124 18028
rect 12084 17882 12112 18022
rect 12072 17876 12124 17882
rect 12072 17818 12124 17824
rect 11572 17700 11652 17728
rect 11520 17682 11572 17688
rect 11440 17202 11468 17682
rect 11428 17196 11480 17202
rect 11428 17138 11480 17144
rect 11336 16788 11388 16794
rect 11336 16730 11388 16736
rect 11428 16652 11480 16658
rect 11428 16594 11480 16600
rect 11152 16584 11204 16590
rect 11152 16526 11204 16532
rect 11060 16448 11112 16454
rect 11060 16390 11112 16396
rect 11072 16250 11100 16390
rect 11060 16244 11112 16250
rect 11060 16186 11112 16192
rect 11164 14958 11192 16526
rect 11244 15904 11296 15910
rect 11244 15846 11296 15852
rect 11256 15570 11284 15846
rect 11440 15706 11468 16594
rect 11428 15700 11480 15706
rect 11428 15642 11480 15648
rect 11244 15564 11296 15570
rect 11244 15506 11296 15512
rect 11532 15502 11560 17682
rect 11888 17672 11940 17678
rect 11888 17614 11940 17620
rect 11900 16046 11928 17614
rect 11888 16040 11940 16046
rect 11888 15982 11940 15988
rect 11336 15496 11388 15502
rect 11336 15438 11388 15444
rect 11520 15496 11572 15502
rect 11520 15438 11572 15444
rect 11242 15192 11298 15201
rect 11242 15127 11298 15136
rect 11152 14952 11204 14958
rect 11152 14894 11204 14900
rect 11256 14482 11284 15127
rect 11348 14550 11376 15438
rect 12176 14890 12204 19366
rect 12256 19236 12308 19242
rect 12256 19178 12308 19184
rect 12268 18902 12296 19178
rect 12256 18896 12308 18902
rect 12256 18838 12308 18844
rect 12360 15026 12388 19858
rect 12440 19712 12492 19718
rect 12440 19654 12492 19660
rect 12452 18834 12480 19654
rect 12440 18828 12492 18834
rect 12440 18770 12492 18776
rect 12440 17740 12492 17746
rect 12440 17682 12492 17688
rect 12452 17338 12480 17682
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 12544 16998 12572 19994
rect 12636 18834 12664 20198
rect 12728 19854 12756 22066
rect 13004 21010 13032 22510
rect 13096 22094 13124 23038
rect 13176 22976 13228 22982
rect 13176 22918 13228 22924
rect 13188 22574 13216 22918
rect 13176 22568 13228 22574
rect 13176 22510 13228 22516
rect 13268 22568 13320 22574
rect 13268 22510 13320 22516
rect 13096 22066 13216 22094
rect 13084 21344 13136 21350
rect 13084 21286 13136 21292
rect 13096 21010 13124 21286
rect 12992 21004 13044 21010
rect 12992 20946 13044 20952
rect 13084 21004 13136 21010
rect 13084 20946 13136 20952
rect 12808 19984 12860 19990
rect 12808 19926 12860 19932
rect 12716 19848 12768 19854
rect 12716 19790 12768 19796
rect 12820 19174 12848 19926
rect 12900 19848 12952 19854
rect 12900 19790 12952 19796
rect 12912 19514 12940 19790
rect 13188 19718 13216 22066
rect 13280 21894 13308 22510
rect 13372 22506 13400 23598
rect 13830 23420 14138 23429
rect 13830 23418 13836 23420
rect 13892 23418 13916 23420
rect 13972 23418 13996 23420
rect 14052 23418 14076 23420
rect 14132 23418 14138 23420
rect 13892 23366 13894 23418
rect 14074 23366 14076 23418
rect 13830 23364 13836 23366
rect 13892 23364 13916 23366
rect 13972 23364 13996 23366
rect 14052 23364 14076 23366
rect 14132 23364 14138 23366
rect 13830 23355 14138 23364
rect 13728 23316 13780 23322
rect 13728 23258 13780 23264
rect 13360 22500 13412 22506
rect 13360 22442 13412 22448
rect 13372 22234 13400 22442
rect 13360 22228 13412 22234
rect 13360 22170 13412 22176
rect 13360 22024 13412 22030
rect 13360 21966 13412 21972
rect 13268 21888 13320 21894
rect 13268 21830 13320 21836
rect 13372 21010 13400 21966
rect 13452 21956 13504 21962
rect 13452 21898 13504 21904
rect 13464 21457 13492 21898
rect 13740 21894 13768 23258
rect 14200 23254 14228 23734
rect 14280 23656 14332 23662
rect 14280 23598 14332 23604
rect 14188 23248 14240 23254
rect 14188 23190 14240 23196
rect 14292 22778 14320 23598
rect 14476 23526 14504 24686
rect 14568 23866 14596 24890
rect 14648 24744 14700 24750
rect 14648 24686 14700 24692
rect 14660 23866 14688 24686
rect 14832 24608 14884 24614
rect 14832 24550 14884 24556
rect 14844 24274 14872 24550
rect 14832 24268 14884 24274
rect 14832 24210 14884 24216
rect 14556 23860 14608 23866
rect 14556 23802 14608 23808
rect 14648 23860 14700 23866
rect 14648 23802 14700 23808
rect 14464 23520 14516 23526
rect 14464 23462 14516 23468
rect 14372 23180 14424 23186
rect 14372 23122 14424 23128
rect 14280 22772 14332 22778
rect 14280 22714 14332 22720
rect 13830 22332 14138 22341
rect 13830 22330 13836 22332
rect 13892 22330 13916 22332
rect 13972 22330 13996 22332
rect 14052 22330 14076 22332
rect 14132 22330 14138 22332
rect 13892 22278 13894 22330
rect 14074 22278 14076 22330
rect 13830 22276 13836 22278
rect 13892 22276 13916 22278
rect 13972 22276 13996 22278
rect 14052 22276 14076 22278
rect 14132 22276 14138 22278
rect 13830 22267 14138 22276
rect 14188 22160 14240 22166
rect 14188 22102 14240 22108
rect 13728 21888 13780 21894
rect 13728 21830 13780 21836
rect 13740 21690 13768 21830
rect 13728 21684 13780 21690
rect 13728 21626 13780 21632
rect 13728 21548 13780 21554
rect 13728 21490 13780 21496
rect 13450 21448 13506 21457
rect 13450 21383 13506 21392
rect 13360 21004 13412 21010
rect 13360 20946 13412 20952
rect 13372 20466 13400 20946
rect 13360 20460 13412 20466
rect 13360 20402 13412 20408
rect 13176 19712 13228 19718
rect 13176 19654 13228 19660
rect 13188 19514 13216 19654
rect 12900 19508 12952 19514
rect 12900 19450 12952 19456
rect 13176 19508 13228 19514
rect 13176 19450 13228 19456
rect 12808 19168 12860 19174
rect 12808 19110 12860 19116
rect 12624 18828 12676 18834
rect 12624 18770 12676 18776
rect 12820 18154 12848 19110
rect 13084 18828 13136 18834
rect 13084 18770 13136 18776
rect 12808 18148 12860 18154
rect 12808 18090 12860 18096
rect 12716 17060 12768 17066
rect 12716 17002 12768 17008
rect 12532 16992 12584 16998
rect 12532 16934 12584 16940
rect 12728 16726 12756 17002
rect 12820 16794 12848 18090
rect 13096 17134 13124 18770
rect 13188 18426 13216 19450
rect 13372 19310 13400 20402
rect 13360 19304 13412 19310
rect 13360 19246 13412 19252
rect 13360 19168 13412 19174
rect 13360 19110 13412 19116
rect 13372 18834 13400 19110
rect 13464 18902 13492 21383
rect 13636 21004 13688 21010
rect 13636 20946 13688 20952
rect 13544 20800 13596 20806
rect 13544 20742 13596 20748
rect 13556 20398 13584 20742
rect 13648 20602 13676 20946
rect 13740 20806 13768 21490
rect 13830 21244 14138 21253
rect 13830 21242 13836 21244
rect 13892 21242 13916 21244
rect 13972 21242 13996 21244
rect 14052 21242 14076 21244
rect 14132 21242 14138 21244
rect 13892 21190 13894 21242
rect 14074 21190 14076 21242
rect 13830 21188 13836 21190
rect 13892 21188 13916 21190
rect 13972 21188 13996 21190
rect 14052 21188 14076 21190
rect 14132 21188 14138 21190
rect 13830 21179 14138 21188
rect 13728 20800 13780 20806
rect 13728 20742 13780 20748
rect 13636 20596 13688 20602
rect 13636 20538 13688 20544
rect 13544 20392 13596 20398
rect 13544 20334 13596 20340
rect 13636 19848 13688 19854
rect 13636 19790 13688 19796
rect 13544 19168 13596 19174
rect 13544 19110 13596 19116
rect 13556 18902 13584 19110
rect 13452 18896 13504 18902
rect 13452 18838 13504 18844
rect 13544 18896 13596 18902
rect 13544 18838 13596 18844
rect 13648 18834 13676 19790
rect 13360 18828 13412 18834
rect 13360 18770 13412 18776
rect 13636 18828 13688 18834
rect 13636 18770 13688 18776
rect 13176 18420 13228 18426
rect 13176 18362 13228 18368
rect 13084 17128 13136 17134
rect 13084 17070 13136 17076
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 12716 16720 12768 16726
rect 12716 16662 12768 16668
rect 12624 16448 12676 16454
rect 12624 16390 12676 16396
rect 12440 15972 12492 15978
rect 12440 15914 12492 15920
rect 12452 15706 12480 15914
rect 12440 15700 12492 15706
rect 12440 15642 12492 15648
rect 12636 15570 12664 16390
rect 12440 15564 12492 15570
rect 12440 15506 12492 15512
rect 12624 15564 12676 15570
rect 12624 15506 12676 15512
rect 12992 15564 13044 15570
rect 13096 15552 13124 17070
rect 13188 16454 13216 18362
rect 13360 18216 13412 18222
rect 13360 18158 13412 18164
rect 13372 17882 13400 18158
rect 13636 18080 13688 18086
rect 13636 18022 13688 18028
rect 13360 17876 13412 17882
rect 13360 17818 13412 17824
rect 13648 17202 13676 18022
rect 13636 17196 13688 17202
rect 13636 17138 13688 17144
rect 13544 17128 13596 17134
rect 13544 17070 13596 17076
rect 13452 16992 13504 16998
rect 13452 16934 13504 16940
rect 13176 16448 13228 16454
rect 13176 16390 13228 16396
rect 13188 16250 13216 16390
rect 13176 16244 13228 16250
rect 13176 16186 13228 16192
rect 13360 15904 13412 15910
rect 13360 15846 13412 15852
rect 13372 15570 13400 15846
rect 13044 15524 13124 15552
rect 13360 15564 13412 15570
rect 12992 15506 13044 15512
rect 13360 15506 13412 15512
rect 12348 15020 12400 15026
rect 12348 14962 12400 14968
rect 12164 14884 12216 14890
rect 12164 14826 12216 14832
rect 11704 14816 11756 14822
rect 11704 14758 11756 14764
rect 11336 14544 11388 14550
rect 11336 14486 11388 14492
rect 11716 14482 11744 14758
rect 11244 14476 11296 14482
rect 11244 14418 11296 14424
rect 11704 14476 11756 14482
rect 11704 14418 11756 14424
rect 11888 14476 11940 14482
rect 11888 14418 11940 14424
rect 12072 14476 12124 14482
rect 12072 14418 12124 14424
rect 10876 14068 10928 14074
rect 10876 14010 10928 14016
rect 10048 14000 10100 14006
rect 10048 13942 10100 13948
rect 9968 13790 10088 13818
rect 8944 13728 8996 13734
rect 8944 13670 8996 13676
rect 9956 13728 10008 13734
rect 9956 13670 10008 13676
rect 8956 13258 8984 13670
rect 9968 13394 9996 13670
rect 9588 13388 9640 13394
rect 9588 13330 9640 13336
rect 9864 13388 9916 13394
rect 9864 13330 9916 13336
rect 9956 13388 10008 13394
rect 9956 13330 10008 13336
rect 8944 13252 8996 13258
rect 8944 13194 8996 13200
rect 8956 12850 8984 13194
rect 9312 13184 9364 13190
rect 9312 13126 9364 13132
rect 9324 12850 9352 13126
rect 9600 12918 9628 13330
rect 9588 12912 9640 12918
rect 9588 12854 9640 12860
rect 9680 12912 9732 12918
rect 9680 12854 9732 12860
rect 8944 12844 8996 12850
rect 8944 12786 8996 12792
rect 9312 12844 9364 12850
rect 9312 12786 9364 12792
rect 9496 12844 9548 12850
rect 9496 12786 9548 12792
rect 8852 12708 8904 12714
rect 8852 12650 8904 12656
rect 8496 12406 8616 12434
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 8220 11150 8248 11630
rect 8208 11144 8260 11150
rect 8208 11086 8260 11092
rect 8024 10056 8076 10062
rect 8024 9998 8076 10004
rect 8036 9042 8064 9998
rect 8484 9988 8536 9994
rect 8484 9930 8536 9936
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 7840 8900 7892 8906
rect 7944 8894 8064 8922
rect 7840 8842 7892 8848
rect 8036 8294 8064 8894
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 8024 8288 8076 8294
rect 8024 8230 8076 8236
rect 8036 7478 8064 8230
rect 8116 7744 8168 7750
rect 8116 7686 8168 7692
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 8024 7472 8076 7478
rect 8024 7414 8076 7420
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7668 7002 7696 7346
rect 7748 7268 7800 7274
rect 7748 7210 7800 7216
rect 7656 6996 7708 7002
rect 7656 6938 7708 6944
rect 7760 6662 7788 7210
rect 7840 7200 7892 7206
rect 7840 7142 7892 7148
rect 7852 6730 7880 7142
rect 7840 6724 7892 6730
rect 7840 6666 7892 6672
rect 7748 6656 7800 6662
rect 7748 6598 7800 6604
rect 7852 6474 7880 6666
rect 7760 6446 7880 6474
rect 7760 6118 7788 6446
rect 8128 6254 8156 7686
rect 8220 7342 8248 7686
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 8116 6248 8168 6254
rect 8116 6190 8168 6196
rect 7748 6112 7800 6118
rect 7748 6054 7800 6060
rect 7932 6112 7984 6118
rect 7932 6054 7984 6060
rect 7760 5370 7788 6054
rect 7748 5364 7800 5370
rect 7748 5306 7800 5312
rect 7840 5296 7892 5302
rect 7840 5238 7892 5244
rect 7012 5092 7064 5098
rect 7012 5034 7064 5040
rect 7564 5092 7616 5098
rect 7564 5034 7616 5040
rect 6920 4548 6972 4554
rect 6920 4490 6972 4496
rect 7024 4078 7052 5034
rect 7114 4924 7422 4933
rect 7114 4922 7120 4924
rect 7176 4922 7200 4924
rect 7256 4922 7280 4924
rect 7336 4922 7360 4924
rect 7416 4922 7422 4924
rect 7176 4870 7178 4922
rect 7358 4870 7360 4922
rect 7114 4868 7120 4870
rect 7176 4868 7200 4870
rect 7256 4868 7280 4870
rect 7336 4868 7360 4870
rect 7416 4868 7422 4870
rect 7114 4859 7422 4868
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 7564 4684 7616 4690
rect 7564 4626 7616 4632
rect 7104 4548 7156 4554
rect 7104 4490 7156 4496
rect 7012 4072 7064 4078
rect 7012 4014 7064 4020
rect 6920 4004 6972 4010
rect 6920 3946 6972 3952
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6460 2984 6512 2990
rect 6460 2926 6512 2932
rect 6092 2576 6144 2582
rect 6092 2518 6144 2524
rect 6184 2508 6236 2514
rect 6184 2450 6236 2456
rect 6000 2440 6052 2446
rect 6000 2382 6052 2388
rect 5540 2304 5592 2310
rect 5540 2246 5592 2252
rect 5908 2304 5960 2310
rect 5908 2246 5960 2252
rect 5264 1896 5316 1902
rect 5184 1856 5264 1884
rect 4620 1838 4672 1844
rect 5264 1838 5316 1844
rect 4264 882 4292 1838
rect 5448 1828 5500 1834
rect 5448 1770 5500 1776
rect 4528 1760 4580 1766
rect 4528 1702 4580 1708
rect 4804 1760 4856 1766
rect 4804 1702 4856 1708
rect 4436 1420 4488 1426
rect 4436 1362 4488 1368
rect 4160 876 4212 882
rect 4160 818 4212 824
rect 4252 876 4304 882
rect 4252 818 4304 824
rect 4448 626 4476 1362
rect 4540 814 4568 1702
rect 4816 1426 4844 1702
rect 4804 1420 4856 1426
rect 4804 1362 4856 1368
rect 5460 1358 5488 1770
rect 5632 1420 5684 1426
rect 5632 1362 5684 1368
rect 5448 1352 5500 1358
rect 5448 1294 5500 1300
rect 5448 1216 5500 1222
rect 5448 1158 5500 1164
rect 5460 1018 5488 1158
rect 5448 1012 5500 1018
rect 5448 954 5500 960
rect 4528 808 4580 814
rect 4528 750 4580 756
rect 5080 808 5132 814
rect 5080 750 5132 756
rect 4448 598 4568 626
rect 3896 462 4016 490
rect 3896 354 3924 462
rect 3988 400 4016 462
rect 4540 400 4568 598
rect 5092 400 5120 750
rect 5644 400 5672 1362
rect 5920 814 5948 2246
rect 6012 2106 6040 2382
rect 6000 2100 6052 2106
rect 6000 2042 6052 2048
rect 5908 808 5960 814
rect 5908 750 5960 756
rect 6196 400 6224 2450
rect 6276 2304 6328 2310
rect 6276 2246 6328 2252
rect 6288 1970 6316 2246
rect 6276 1964 6328 1970
rect 6276 1906 6328 1912
rect 6564 1902 6592 3470
rect 6840 3194 6868 3538
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 6840 2582 6868 3130
rect 6932 2990 6960 3946
rect 7116 3924 7144 4490
rect 7576 4282 7604 4626
rect 7564 4276 7616 4282
rect 7564 4218 7616 4224
rect 7656 4072 7708 4078
rect 7656 4014 7708 4020
rect 7024 3896 7144 3924
rect 7564 3936 7616 3942
rect 7024 3670 7052 3896
rect 7564 3878 7616 3884
rect 7114 3836 7422 3845
rect 7114 3834 7120 3836
rect 7176 3834 7200 3836
rect 7256 3834 7280 3836
rect 7336 3834 7360 3836
rect 7416 3834 7422 3836
rect 7176 3782 7178 3834
rect 7358 3782 7360 3834
rect 7114 3780 7120 3782
rect 7176 3780 7200 3782
rect 7256 3780 7280 3782
rect 7336 3780 7360 3782
rect 7416 3780 7422 3782
rect 7114 3771 7422 3780
rect 7012 3664 7064 3670
rect 7012 3606 7064 3612
rect 7576 3482 7604 3878
rect 7668 3602 7696 4014
rect 7656 3596 7708 3602
rect 7656 3538 7708 3544
rect 7300 3466 7604 3482
rect 7288 3460 7604 3466
rect 7340 3454 7604 3460
rect 7288 3402 7340 3408
rect 6920 2984 6972 2990
rect 6920 2926 6972 2932
rect 6932 2582 6960 2926
rect 7114 2748 7422 2757
rect 7114 2746 7120 2748
rect 7176 2746 7200 2748
rect 7256 2746 7280 2748
rect 7336 2746 7360 2748
rect 7416 2746 7422 2748
rect 7176 2694 7178 2746
rect 7358 2694 7360 2746
rect 7114 2692 7120 2694
rect 7176 2692 7200 2694
rect 7256 2692 7280 2694
rect 7336 2692 7360 2694
rect 7416 2692 7422 2694
rect 7114 2683 7422 2692
rect 6828 2576 6880 2582
rect 6828 2518 6880 2524
rect 6920 2576 6972 2582
rect 6920 2518 6972 2524
rect 7576 2514 7604 3454
rect 7760 2990 7788 4762
rect 7852 4078 7880 5238
rect 7944 5166 7972 6054
rect 8208 5772 8260 5778
rect 8208 5714 8260 5720
rect 8220 5370 8248 5714
rect 8208 5364 8260 5370
rect 8208 5306 8260 5312
rect 8312 5302 8340 8774
rect 8300 5296 8352 5302
rect 8300 5238 8352 5244
rect 7932 5160 7984 5166
rect 7932 5102 7984 5108
rect 8300 4820 8352 4826
rect 8404 4808 8432 9862
rect 8496 8566 8524 9930
rect 8484 8560 8536 8566
rect 8484 8502 8536 8508
rect 8588 7426 8616 12406
rect 8864 11286 8892 12650
rect 9128 12096 9180 12102
rect 9128 12038 9180 12044
rect 9140 11354 9168 12038
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 9128 11348 9180 11354
rect 9128 11290 9180 11296
rect 8852 11280 8904 11286
rect 8852 11222 8904 11228
rect 8944 11076 8996 11082
rect 8944 11018 8996 11024
rect 8956 10606 8984 11018
rect 9140 11014 9168 11290
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 9128 11008 9180 11014
rect 9128 10950 9180 10956
rect 9140 10606 9168 10950
rect 9232 10606 9260 11086
rect 9312 11008 9364 11014
rect 9312 10950 9364 10956
rect 9324 10606 9352 10950
rect 8944 10600 8996 10606
rect 8944 10542 8996 10548
rect 9128 10600 9180 10606
rect 9128 10542 9180 10548
rect 9220 10600 9272 10606
rect 9220 10542 9272 10548
rect 9312 10600 9364 10606
rect 9312 10542 9364 10548
rect 8852 10464 8904 10470
rect 8852 10406 8904 10412
rect 8944 10464 8996 10470
rect 8944 10406 8996 10412
rect 8668 10124 8720 10130
rect 8668 10066 8720 10072
rect 8680 9382 8708 10066
rect 8760 10056 8812 10062
rect 8760 9998 8812 10004
rect 8772 9518 8800 9998
rect 8760 9512 8812 9518
rect 8760 9454 8812 9460
rect 8668 9376 8720 9382
rect 8668 9318 8720 9324
rect 8680 8974 8708 9318
rect 8668 8968 8720 8974
rect 8668 8910 8720 8916
rect 8864 7936 8892 10406
rect 8956 10130 8984 10406
rect 9140 10130 9168 10542
rect 8944 10124 8996 10130
rect 8944 10066 8996 10072
rect 9128 10124 9180 10130
rect 9128 10066 9180 10072
rect 9036 9920 9088 9926
rect 9036 9862 9088 9868
rect 8944 9376 8996 9382
rect 8944 9318 8996 9324
rect 8772 7908 8892 7936
rect 8588 7398 8708 7426
rect 8576 7268 8628 7274
rect 8576 7210 8628 7216
rect 8588 4826 8616 7210
rect 8680 6934 8708 7398
rect 8668 6928 8720 6934
rect 8668 6870 8720 6876
rect 8680 6186 8708 6870
rect 8668 6180 8720 6186
rect 8668 6122 8720 6128
rect 8352 4780 8432 4808
rect 8576 4820 8628 4826
rect 8300 4762 8352 4768
rect 8576 4762 8628 4768
rect 8772 4078 8800 7908
rect 8852 7812 8904 7818
rect 8852 7754 8904 7760
rect 8864 7478 8892 7754
rect 8852 7472 8904 7478
rect 8852 7414 8904 7420
rect 8852 5772 8904 5778
rect 8852 5714 8904 5720
rect 8864 5370 8892 5714
rect 8852 5364 8904 5370
rect 8852 5306 8904 5312
rect 7840 4072 7892 4078
rect 7840 4014 7892 4020
rect 8024 4072 8076 4078
rect 8024 4014 8076 4020
rect 8116 4072 8168 4078
rect 8116 4014 8168 4020
rect 8760 4072 8812 4078
rect 8956 4060 8984 9318
rect 9048 9042 9076 9862
rect 9140 9518 9168 10066
rect 9220 10056 9272 10062
rect 9324 10044 9352 10542
rect 9416 10146 9444 11494
rect 9508 10606 9536 12786
rect 9692 12714 9720 12854
rect 9876 12850 9904 13330
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 9680 12708 9732 12714
rect 9680 12650 9732 12656
rect 9692 12434 9720 12650
rect 9772 12640 9824 12646
rect 9772 12582 9824 12588
rect 9600 12406 9720 12434
rect 9600 12374 9628 12406
rect 9784 12374 9812 12582
rect 9588 12368 9640 12374
rect 9588 12310 9640 12316
rect 9772 12368 9824 12374
rect 9772 12310 9824 12316
rect 9588 12232 9640 12238
rect 9588 12174 9640 12180
rect 9600 11898 9628 12174
rect 9588 11892 9640 11898
rect 9588 11834 9640 11840
rect 9600 11286 9628 11834
rect 9588 11280 9640 11286
rect 9588 11222 9640 11228
rect 9784 11082 9812 12310
rect 9876 11218 9904 12786
rect 9968 12434 9996 13330
rect 10060 12918 10088 13790
rect 10324 13796 10376 13802
rect 10324 13738 10376 13744
rect 10336 12986 10364 13738
rect 10888 13394 10916 14010
rect 10968 13864 11020 13870
rect 10968 13806 11020 13812
rect 10876 13388 10928 13394
rect 10876 13330 10928 13336
rect 10876 13184 10928 13190
rect 10876 13126 10928 13132
rect 10472 13084 10780 13093
rect 10472 13082 10478 13084
rect 10534 13082 10558 13084
rect 10614 13082 10638 13084
rect 10694 13082 10718 13084
rect 10774 13082 10780 13084
rect 10534 13030 10536 13082
rect 10716 13030 10718 13082
rect 10472 13028 10478 13030
rect 10534 13028 10558 13030
rect 10614 13028 10638 13030
rect 10694 13028 10718 13030
rect 10774 13028 10780 13030
rect 10472 13019 10780 13028
rect 10888 12986 10916 13126
rect 10324 12980 10376 12986
rect 10324 12922 10376 12928
rect 10876 12980 10928 12986
rect 10876 12922 10928 12928
rect 10048 12912 10100 12918
rect 10048 12854 10100 12860
rect 10784 12912 10836 12918
rect 10784 12854 10836 12860
rect 10796 12714 10824 12854
rect 10784 12708 10836 12714
rect 10784 12650 10836 12656
rect 10980 12646 11008 13806
rect 10324 12640 10376 12646
rect 10324 12582 10376 12588
rect 10968 12640 11020 12646
rect 10968 12582 11020 12588
rect 9968 12406 10088 12434
rect 9956 12368 10008 12374
rect 9956 12310 10008 12316
rect 9968 11354 9996 12310
rect 9956 11348 10008 11354
rect 9956 11290 10008 11296
rect 9864 11212 9916 11218
rect 9864 11154 9916 11160
rect 9772 11076 9824 11082
rect 9772 11018 9824 11024
rect 9772 10736 9824 10742
rect 9772 10678 9824 10684
rect 9496 10600 9548 10606
rect 9496 10542 9548 10548
rect 9416 10118 9536 10146
rect 9272 10016 9352 10044
rect 9404 10056 9456 10062
rect 9220 9998 9272 10004
rect 9404 9998 9456 10004
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 9232 9042 9260 9998
rect 9416 9586 9444 9998
rect 9404 9580 9456 9586
rect 9324 9540 9404 9568
rect 9036 9036 9088 9042
rect 9036 8978 9088 8984
rect 9220 9036 9272 9042
rect 9220 8978 9272 8984
rect 9324 8974 9352 9540
rect 9404 9522 9456 9528
rect 9508 9500 9536 10118
rect 9784 9926 9812 10678
rect 9876 10674 9904 11154
rect 9864 10668 9916 10674
rect 9864 10610 9916 10616
rect 10060 10130 10088 12406
rect 10336 12102 10364 12582
rect 10232 12096 10284 12102
rect 10232 12038 10284 12044
rect 10324 12096 10376 12102
rect 10324 12038 10376 12044
rect 10244 11218 10272 12038
rect 10472 11996 10780 12005
rect 10472 11994 10478 11996
rect 10534 11994 10558 11996
rect 10614 11994 10638 11996
rect 10694 11994 10718 11996
rect 10774 11994 10780 11996
rect 10534 11942 10536 11994
rect 10716 11942 10718 11994
rect 10472 11940 10478 11942
rect 10534 11940 10558 11942
rect 10614 11940 10638 11942
rect 10694 11940 10718 11942
rect 10774 11940 10780 11942
rect 10472 11931 10780 11940
rect 10416 11620 10468 11626
rect 10416 11562 10468 11568
rect 10428 11354 10456 11562
rect 10416 11348 10468 11354
rect 10416 11290 10468 11296
rect 10232 11212 10284 11218
rect 10232 11154 10284 11160
rect 10980 11082 11008 12582
rect 10324 11076 10376 11082
rect 10324 11018 10376 11024
rect 10968 11076 11020 11082
rect 10968 11018 11020 11024
rect 10336 10690 10364 11018
rect 10472 10908 10780 10917
rect 10472 10906 10478 10908
rect 10534 10906 10558 10908
rect 10614 10906 10638 10908
rect 10694 10906 10718 10908
rect 10774 10906 10780 10908
rect 10534 10854 10536 10906
rect 10716 10854 10718 10906
rect 10472 10852 10478 10854
rect 10534 10852 10558 10854
rect 10614 10852 10638 10854
rect 10694 10852 10718 10854
rect 10774 10852 10780 10854
rect 10472 10843 10780 10852
rect 11256 10742 11284 14418
rect 11520 13796 11572 13802
rect 11520 13738 11572 13744
rect 11532 13394 11560 13738
rect 11900 13734 11928 14418
rect 12084 14074 12112 14418
rect 12072 14068 12124 14074
rect 12072 14010 12124 14016
rect 12176 13802 12204 14826
rect 12452 14770 12480 15506
rect 13004 15162 13032 15506
rect 12992 15156 13044 15162
rect 12992 15098 13044 15104
rect 12624 14952 12676 14958
rect 12624 14894 12676 14900
rect 12360 14742 12480 14770
rect 12164 13796 12216 13802
rect 12164 13738 12216 13744
rect 11888 13728 11940 13734
rect 11888 13670 11940 13676
rect 11520 13388 11572 13394
rect 11520 13330 11572 13336
rect 11336 13184 11388 13190
rect 11336 13126 11388 13132
rect 11348 12646 11376 13126
rect 11900 12782 11928 13670
rect 12164 12980 12216 12986
rect 12164 12922 12216 12928
rect 11888 12776 11940 12782
rect 11888 12718 11940 12724
rect 11520 12708 11572 12714
rect 11520 12650 11572 12656
rect 11336 12640 11388 12646
rect 11388 12600 11468 12628
rect 11336 12582 11388 12588
rect 11440 12306 11468 12600
rect 11532 12442 11560 12650
rect 11704 12640 11756 12646
rect 11704 12582 11756 12588
rect 11520 12436 11572 12442
rect 11520 12378 11572 12384
rect 11716 12306 11744 12582
rect 11336 12300 11388 12306
rect 11336 12242 11388 12248
rect 11428 12300 11480 12306
rect 11428 12242 11480 12248
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 11348 11558 11376 12242
rect 11900 12238 11928 12718
rect 12176 12306 12204 12922
rect 12256 12436 12308 12442
rect 12360 12434 12388 14742
rect 12636 13870 12664 14894
rect 12900 14816 12952 14822
rect 12900 14758 12952 14764
rect 12624 13864 12676 13870
rect 12624 13806 12676 13812
rect 12440 13728 12492 13734
rect 12440 13670 12492 13676
rect 12452 13530 12480 13670
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12636 12986 12664 13806
rect 12912 13734 12940 14758
rect 13464 14278 13492 16934
rect 13556 15570 13584 17070
rect 13740 16980 13768 20742
rect 13830 20156 14138 20165
rect 13830 20154 13836 20156
rect 13892 20154 13916 20156
rect 13972 20154 13996 20156
rect 14052 20154 14076 20156
rect 14132 20154 14138 20156
rect 13892 20102 13894 20154
rect 14074 20102 14076 20154
rect 13830 20100 13836 20102
rect 13892 20100 13916 20102
rect 13972 20100 13996 20102
rect 14052 20100 14076 20102
rect 14132 20100 14138 20102
rect 13830 20091 14138 20100
rect 13820 19712 13872 19718
rect 13820 19654 13872 19660
rect 14096 19712 14148 19718
rect 14096 19654 14148 19660
rect 13832 19514 13860 19654
rect 13820 19508 13872 19514
rect 13820 19450 13872 19456
rect 14108 19310 14136 19654
rect 14200 19417 14228 22102
rect 14384 21554 14412 23122
rect 14476 22710 14504 23462
rect 14556 23248 14608 23254
rect 14556 23190 14608 23196
rect 14464 22704 14516 22710
rect 14464 22646 14516 22652
rect 14464 22228 14516 22234
rect 14464 22170 14516 22176
rect 14372 21548 14424 21554
rect 14372 21490 14424 21496
rect 14186 19408 14242 19417
rect 14186 19343 14242 19352
rect 14096 19304 14148 19310
rect 14096 19246 14148 19252
rect 13830 19068 14138 19077
rect 13830 19066 13836 19068
rect 13892 19066 13916 19068
rect 13972 19066 13996 19068
rect 14052 19066 14076 19068
rect 14132 19066 14138 19068
rect 13892 19014 13894 19066
rect 14074 19014 14076 19066
rect 13830 19012 13836 19014
rect 13892 19012 13916 19014
rect 13972 19012 13996 19014
rect 14052 19012 14076 19014
rect 14132 19012 14138 19014
rect 13830 19003 14138 19012
rect 14372 18828 14424 18834
rect 14372 18770 14424 18776
rect 14384 18222 14412 18770
rect 14372 18216 14424 18222
rect 14372 18158 14424 18164
rect 14188 18080 14240 18086
rect 14188 18022 14240 18028
rect 14280 18080 14332 18086
rect 14280 18022 14332 18028
rect 13830 17980 14138 17989
rect 13830 17978 13836 17980
rect 13892 17978 13916 17980
rect 13972 17978 13996 17980
rect 14052 17978 14076 17980
rect 14132 17978 14138 17980
rect 13892 17926 13894 17978
rect 14074 17926 14076 17978
rect 13830 17924 13836 17926
rect 13892 17924 13916 17926
rect 13972 17924 13996 17926
rect 14052 17924 14076 17926
rect 14132 17924 14138 17926
rect 13830 17915 14138 17924
rect 14200 17746 14228 18022
rect 14292 17882 14320 18022
rect 14280 17876 14332 17882
rect 14280 17818 14332 17824
rect 14188 17740 14240 17746
rect 14188 17682 14240 17688
rect 13820 16992 13872 16998
rect 13740 16952 13820 16980
rect 13740 16946 13768 16952
rect 13648 16918 13768 16946
rect 13820 16934 13872 16940
rect 13648 16658 13676 16918
rect 13830 16892 14138 16901
rect 13830 16890 13836 16892
rect 13892 16890 13916 16892
rect 13972 16890 13996 16892
rect 14052 16890 14076 16892
rect 14132 16890 14138 16892
rect 13892 16838 13894 16890
rect 14074 16838 14076 16890
rect 13830 16836 13836 16838
rect 13892 16836 13916 16838
rect 13972 16836 13996 16838
rect 14052 16836 14076 16838
rect 14132 16836 14138 16838
rect 13830 16827 14138 16836
rect 14476 16794 14504 22170
rect 14568 21622 14596 23190
rect 14936 22642 14964 25298
rect 15016 25288 15068 25294
rect 15016 25230 15068 25236
rect 15028 24274 15056 25230
rect 15108 24608 15160 24614
rect 15108 24550 15160 24556
rect 15016 24268 15068 24274
rect 15016 24210 15068 24216
rect 15028 23798 15056 24210
rect 15016 23792 15068 23798
rect 15016 23734 15068 23740
rect 15120 23730 15148 24550
rect 15108 23724 15160 23730
rect 15108 23666 15160 23672
rect 15292 23724 15344 23730
rect 15292 23666 15344 23672
rect 15016 23520 15068 23526
rect 15016 23462 15068 23468
rect 15028 23322 15056 23462
rect 15016 23316 15068 23322
rect 15016 23258 15068 23264
rect 14924 22636 14976 22642
rect 14924 22578 14976 22584
rect 14740 22568 14792 22574
rect 14740 22510 14792 22516
rect 14752 21622 14780 22510
rect 14936 22094 14964 22578
rect 15304 22574 15332 23666
rect 15396 23474 15424 26279
rect 15476 25832 15528 25838
rect 15476 25774 15528 25780
rect 15488 24954 15516 25774
rect 15476 24948 15528 24954
rect 15476 24890 15528 24896
rect 15580 24818 15608 26862
rect 15660 26784 15712 26790
rect 15660 26726 15712 26732
rect 15672 26450 15700 26726
rect 15660 26444 15712 26450
rect 15660 26386 15712 26392
rect 15764 25906 15792 28562
rect 15856 27538 15884 28630
rect 16684 27538 16712 28970
rect 16776 28422 16804 29038
rect 16868 28626 16896 29514
rect 16948 29504 17000 29510
rect 16948 29446 17000 29452
rect 16856 28620 16908 28626
rect 16856 28562 16908 28568
rect 16764 28416 16816 28422
rect 16764 28358 16816 28364
rect 16868 28014 16896 28562
rect 16856 28008 16908 28014
rect 16856 27950 16908 27956
rect 16764 27600 16816 27606
rect 16764 27542 16816 27548
rect 15844 27532 15896 27538
rect 15844 27474 15896 27480
rect 16672 27532 16724 27538
rect 16672 27474 16724 27480
rect 16304 27124 16356 27130
rect 16304 27066 16356 27072
rect 15844 26920 15896 26926
rect 15844 26862 15896 26868
rect 15856 26042 15884 26862
rect 16316 26450 16344 27066
rect 16776 26790 16804 27542
rect 16856 27396 16908 27402
rect 16856 27338 16908 27344
rect 16764 26784 16816 26790
rect 16764 26726 16816 26732
rect 16580 26580 16632 26586
rect 16580 26522 16632 26528
rect 16672 26580 16724 26586
rect 16672 26522 16724 26528
rect 16304 26444 16356 26450
rect 16304 26386 16356 26392
rect 16028 26308 16080 26314
rect 16028 26250 16080 26256
rect 15844 26036 15896 26042
rect 15844 25978 15896 25984
rect 15752 25900 15804 25906
rect 15752 25842 15804 25848
rect 16040 25838 16068 26250
rect 16396 26240 16448 26246
rect 16396 26182 16448 26188
rect 16408 26042 16436 26182
rect 16396 26036 16448 26042
rect 16396 25978 16448 25984
rect 16592 25838 16620 26522
rect 16684 26450 16712 26522
rect 16672 26444 16724 26450
rect 16672 26386 16724 26392
rect 16684 26353 16712 26386
rect 16670 26344 16726 26353
rect 16670 26279 16726 26288
rect 16672 25968 16724 25974
rect 16670 25936 16672 25945
rect 16724 25936 16726 25945
rect 16776 25906 16804 26726
rect 16670 25871 16726 25880
rect 16764 25900 16816 25906
rect 16764 25842 16816 25848
rect 16028 25832 16080 25838
rect 16028 25774 16080 25780
rect 16580 25832 16632 25838
rect 16868 25786 16896 27338
rect 16960 26994 16988 29446
rect 17188 29404 17496 29413
rect 17188 29402 17194 29404
rect 17250 29402 17274 29404
rect 17330 29402 17354 29404
rect 17410 29402 17434 29404
rect 17490 29402 17496 29404
rect 17250 29350 17252 29402
rect 17432 29350 17434 29402
rect 17188 29348 17194 29350
rect 17250 29348 17274 29350
rect 17330 29348 17354 29350
rect 17410 29348 17434 29350
rect 17490 29348 17496 29350
rect 17188 29339 17496 29348
rect 17132 29232 17184 29238
rect 17132 29174 17184 29180
rect 17040 28960 17092 28966
rect 17040 28902 17092 28908
rect 17052 28626 17080 28902
rect 17040 28620 17092 28626
rect 17040 28562 17092 28568
rect 17144 28404 17172 29174
rect 17592 28620 17644 28626
rect 17592 28562 17644 28568
rect 17052 28376 17172 28404
rect 17052 28098 17080 28376
rect 17188 28316 17496 28325
rect 17188 28314 17194 28316
rect 17250 28314 17274 28316
rect 17330 28314 17354 28316
rect 17410 28314 17434 28316
rect 17490 28314 17496 28316
rect 17250 28262 17252 28314
rect 17432 28262 17434 28314
rect 17188 28260 17194 28262
rect 17250 28260 17274 28262
rect 17330 28260 17354 28262
rect 17410 28260 17434 28262
rect 17490 28260 17496 28262
rect 17188 28251 17496 28260
rect 17052 28070 17172 28098
rect 17040 28008 17092 28014
rect 17040 27950 17092 27956
rect 17052 27470 17080 27950
rect 17040 27464 17092 27470
rect 17040 27406 17092 27412
rect 16948 26988 17000 26994
rect 16948 26930 17000 26936
rect 16948 26376 17000 26382
rect 16948 26318 17000 26324
rect 16580 25774 16632 25780
rect 15752 24948 15804 24954
rect 15752 24890 15804 24896
rect 15568 24812 15620 24818
rect 15568 24754 15620 24760
rect 15580 24410 15608 24754
rect 15660 24744 15712 24750
rect 15660 24686 15712 24692
rect 15672 24410 15700 24686
rect 15568 24404 15620 24410
rect 15568 24346 15620 24352
rect 15660 24404 15712 24410
rect 15660 24346 15712 24352
rect 15660 23588 15712 23594
rect 15660 23530 15712 23536
rect 15396 23446 15608 23474
rect 15382 23216 15438 23225
rect 15382 23151 15438 23160
rect 15292 22568 15344 22574
rect 15212 22528 15292 22556
rect 14936 22066 15148 22094
rect 14556 21616 14608 21622
rect 14556 21558 14608 21564
rect 14740 21616 14792 21622
rect 14740 21558 14792 21564
rect 15120 21418 15148 22066
rect 15212 22030 15240 22528
rect 15292 22510 15344 22516
rect 15396 22420 15424 23151
rect 15476 22976 15528 22982
rect 15476 22918 15528 22924
rect 15488 22574 15516 22918
rect 15476 22568 15528 22574
rect 15476 22510 15528 22516
rect 15476 22432 15528 22438
rect 15396 22392 15476 22420
rect 15476 22374 15528 22380
rect 15292 22160 15344 22166
rect 15292 22102 15344 22108
rect 15200 22024 15252 22030
rect 15200 21966 15252 21972
rect 15212 21554 15240 21966
rect 15200 21548 15252 21554
rect 15200 21490 15252 21496
rect 15304 21486 15332 22102
rect 15292 21480 15344 21486
rect 15292 21422 15344 21428
rect 15108 21412 15160 21418
rect 15108 21354 15160 21360
rect 15304 21146 15332 21422
rect 15292 21140 15344 21146
rect 15292 21082 15344 21088
rect 15488 21010 15516 22374
rect 15292 21004 15344 21010
rect 15292 20946 15344 20952
rect 15384 21004 15436 21010
rect 15384 20946 15436 20952
rect 15476 21004 15528 21010
rect 15476 20946 15528 20952
rect 15016 20936 15068 20942
rect 15016 20878 15068 20884
rect 14832 20392 14884 20398
rect 14832 20334 14884 20340
rect 14844 20058 14872 20334
rect 14832 20052 14884 20058
rect 14832 19994 14884 20000
rect 14648 19848 14700 19854
rect 14648 19790 14700 19796
rect 14660 19446 14688 19790
rect 15028 19718 15056 20878
rect 15304 20262 15332 20946
rect 15396 20602 15424 20946
rect 15384 20596 15436 20602
rect 15384 20538 15436 20544
rect 15292 20256 15344 20262
rect 15292 20198 15344 20204
rect 15304 19990 15332 20198
rect 15384 20052 15436 20058
rect 15384 19994 15436 20000
rect 15292 19984 15344 19990
rect 15292 19926 15344 19932
rect 15016 19712 15068 19718
rect 15016 19654 15068 19660
rect 14648 19440 14700 19446
rect 14648 19382 14700 19388
rect 15304 19310 15332 19926
rect 15200 19304 15252 19310
rect 15200 19246 15252 19252
rect 15292 19304 15344 19310
rect 15292 19246 15344 19252
rect 15016 19168 15068 19174
rect 15016 19110 15068 19116
rect 15028 18222 15056 19110
rect 15212 18902 15240 19246
rect 15200 18896 15252 18902
rect 15200 18838 15252 18844
rect 15304 18748 15332 19246
rect 15212 18720 15332 18748
rect 15016 18216 15068 18222
rect 15108 18216 15160 18222
rect 15016 18158 15068 18164
rect 15106 18184 15108 18193
rect 15160 18184 15162 18193
rect 15106 18119 15162 18128
rect 15212 18086 15240 18720
rect 15396 18086 15424 19994
rect 15488 19242 15516 20946
rect 15580 19904 15608 23446
rect 15672 21350 15700 23530
rect 15764 23186 15792 24890
rect 15936 24744 15988 24750
rect 15936 24686 15988 24692
rect 15948 24342 15976 24686
rect 15936 24336 15988 24342
rect 15936 24278 15988 24284
rect 15844 23520 15896 23526
rect 15844 23462 15896 23468
rect 15752 23180 15804 23186
rect 15752 23122 15804 23128
rect 15764 21962 15792 23122
rect 15856 23089 15884 23462
rect 15842 23080 15898 23089
rect 15842 23015 15898 23024
rect 15752 21956 15804 21962
rect 15752 21898 15804 21904
rect 15660 21344 15712 21350
rect 15660 21286 15712 21292
rect 15752 21140 15804 21146
rect 15752 21082 15804 21088
rect 15660 20936 15712 20942
rect 15660 20878 15712 20884
rect 15672 20058 15700 20878
rect 15764 20806 15792 21082
rect 15752 20800 15804 20806
rect 15752 20742 15804 20748
rect 15752 20596 15804 20602
rect 15752 20538 15804 20544
rect 15660 20052 15712 20058
rect 15660 19994 15712 20000
rect 15764 19922 15792 20538
rect 15856 20534 15884 23015
rect 15936 21344 15988 21350
rect 15936 21286 15988 21292
rect 15844 20528 15896 20534
rect 15844 20470 15896 20476
rect 15660 19916 15712 19922
rect 15580 19876 15660 19904
rect 15660 19858 15712 19864
rect 15752 19916 15804 19922
rect 15752 19858 15804 19864
rect 15672 19825 15700 19858
rect 15658 19816 15714 19825
rect 15658 19751 15714 19760
rect 15764 19718 15792 19858
rect 15752 19712 15804 19718
rect 15752 19654 15804 19660
rect 15844 19712 15896 19718
rect 15844 19654 15896 19660
rect 15764 19310 15792 19654
rect 15856 19310 15884 19654
rect 15752 19304 15804 19310
rect 15752 19246 15804 19252
rect 15844 19304 15896 19310
rect 15844 19246 15896 19252
rect 15476 19236 15528 19242
rect 15476 19178 15528 19184
rect 15752 19168 15804 19174
rect 15752 19110 15804 19116
rect 15764 18290 15792 19110
rect 15752 18284 15804 18290
rect 15752 18226 15804 18232
rect 15200 18080 15252 18086
rect 15200 18022 15252 18028
rect 15292 18080 15344 18086
rect 15292 18022 15344 18028
rect 15384 18080 15436 18086
rect 15384 18022 15436 18028
rect 15304 17814 15332 18022
rect 15292 17808 15344 17814
rect 15292 17750 15344 17756
rect 15108 17740 15160 17746
rect 15108 17682 15160 17688
rect 14740 17536 14792 17542
rect 14740 17478 14792 17484
rect 13728 16788 13780 16794
rect 13728 16730 13780 16736
rect 14464 16788 14516 16794
rect 14464 16730 14516 16736
rect 13636 16652 13688 16658
rect 13636 16594 13688 16600
rect 13544 15564 13596 15570
rect 13544 15506 13596 15512
rect 13556 14890 13584 15506
rect 13648 15026 13676 16594
rect 13740 15978 13768 16730
rect 14188 16720 14240 16726
rect 14188 16662 14240 16668
rect 13820 16584 13872 16590
rect 13820 16526 13872 16532
rect 13832 16046 13860 16526
rect 13820 16040 13872 16046
rect 13820 15982 13872 15988
rect 13728 15972 13780 15978
rect 13728 15914 13780 15920
rect 13830 15804 14138 15813
rect 13830 15802 13836 15804
rect 13892 15802 13916 15804
rect 13972 15802 13996 15804
rect 14052 15802 14076 15804
rect 14132 15802 14138 15804
rect 13892 15750 13894 15802
rect 14074 15750 14076 15802
rect 13830 15748 13836 15750
rect 13892 15748 13916 15750
rect 13972 15748 13996 15750
rect 14052 15748 14076 15750
rect 14132 15748 14138 15750
rect 13830 15739 14138 15748
rect 13636 15020 13688 15026
rect 13636 14962 13688 14968
rect 14200 14958 14228 16662
rect 14752 16658 14780 17478
rect 14464 16652 14516 16658
rect 14464 16594 14516 16600
rect 14740 16652 14792 16658
rect 14740 16594 14792 16600
rect 14476 15978 14504 16594
rect 15120 16590 15148 17682
rect 15396 17678 15424 18022
rect 15660 17876 15712 17882
rect 15660 17818 15712 17824
rect 15384 17672 15436 17678
rect 15384 17614 15436 17620
rect 15292 17604 15344 17610
rect 15292 17546 15344 17552
rect 15304 17270 15332 17546
rect 15396 17338 15424 17614
rect 15384 17332 15436 17338
rect 15384 17274 15436 17280
rect 15200 17264 15252 17270
rect 15200 17206 15252 17212
rect 15292 17264 15344 17270
rect 15292 17206 15344 17212
rect 15212 16658 15240 17206
rect 15304 16794 15332 17206
rect 15292 16788 15344 16794
rect 15292 16730 15344 16736
rect 15304 16658 15332 16730
rect 15200 16652 15252 16658
rect 15200 16594 15252 16600
rect 15292 16652 15344 16658
rect 15292 16594 15344 16600
rect 15568 16652 15620 16658
rect 15568 16594 15620 16600
rect 15108 16584 15160 16590
rect 15108 16526 15160 16532
rect 15120 16250 15148 16526
rect 15108 16244 15160 16250
rect 15108 16186 15160 16192
rect 15212 16046 15240 16594
rect 15580 16250 15608 16594
rect 15568 16244 15620 16250
rect 15568 16186 15620 16192
rect 15672 16046 15700 17818
rect 15764 17728 15792 18226
rect 15856 18154 15884 19246
rect 15948 18698 15976 21286
rect 15936 18692 15988 18698
rect 15936 18634 15988 18640
rect 15844 18148 15896 18154
rect 15844 18090 15896 18096
rect 15844 17740 15896 17746
rect 15764 17700 15844 17728
rect 15844 17682 15896 17688
rect 15752 17536 15804 17542
rect 15752 17478 15804 17484
rect 15764 17202 15792 17478
rect 15752 17196 15804 17202
rect 15752 17138 15804 17144
rect 15856 16726 15884 17682
rect 15844 16720 15896 16726
rect 15844 16662 15896 16668
rect 15934 16688 15990 16697
rect 15934 16623 15936 16632
rect 15988 16623 15990 16632
rect 15936 16594 15988 16600
rect 15752 16448 15804 16454
rect 15752 16390 15804 16396
rect 15200 16040 15252 16046
rect 15200 15982 15252 15988
rect 15660 16040 15712 16046
rect 15660 15982 15712 15988
rect 14464 15972 14516 15978
rect 14464 15914 14516 15920
rect 14476 15706 14504 15914
rect 14464 15700 14516 15706
rect 14464 15642 14516 15648
rect 15568 15564 15620 15570
rect 15764 15552 15792 16390
rect 15620 15524 15792 15552
rect 15568 15506 15620 15512
rect 15200 15496 15252 15502
rect 15200 15438 15252 15444
rect 14832 15088 14884 15094
rect 14832 15030 14884 15036
rect 14188 14952 14240 14958
rect 14188 14894 14240 14900
rect 14280 14952 14332 14958
rect 14280 14894 14332 14900
rect 13544 14884 13596 14890
rect 13544 14826 13596 14832
rect 13830 14716 14138 14725
rect 13830 14714 13836 14716
rect 13892 14714 13916 14716
rect 13972 14714 13996 14716
rect 14052 14714 14076 14716
rect 14132 14714 14138 14716
rect 13892 14662 13894 14714
rect 14074 14662 14076 14714
rect 13830 14660 13836 14662
rect 13892 14660 13916 14662
rect 13972 14660 13996 14662
rect 14052 14660 14076 14662
rect 14132 14660 14138 14662
rect 13830 14651 14138 14660
rect 13176 14272 13228 14278
rect 13176 14214 13228 14220
rect 13268 14272 13320 14278
rect 13268 14214 13320 14220
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 12992 13796 13044 13802
rect 12992 13738 13044 13744
rect 12900 13728 12952 13734
rect 12900 13670 12952 13676
rect 12808 13184 12860 13190
rect 12808 13126 12860 13132
rect 12820 12986 12848 13126
rect 12624 12980 12676 12986
rect 12544 12940 12624 12968
rect 12440 12708 12492 12714
rect 12440 12650 12492 12656
rect 12308 12406 12388 12434
rect 12256 12378 12308 12384
rect 12164 12300 12216 12306
rect 11992 12260 12164 12288
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11900 11762 11928 12174
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 11888 11348 11940 11354
rect 11888 11290 11940 11296
rect 11612 11212 11664 11218
rect 11612 11154 11664 11160
rect 11336 10804 11388 10810
rect 11336 10746 11388 10752
rect 11244 10736 11296 10742
rect 10336 10662 10456 10690
rect 11244 10678 11296 10684
rect 10324 10600 10376 10606
rect 10324 10542 10376 10548
rect 10140 10464 10192 10470
rect 10140 10406 10192 10412
rect 10152 10198 10180 10406
rect 10336 10266 10364 10542
rect 10324 10260 10376 10266
rect 10324 10202 10376 10208
rect 10428 10198 10456 10662
rect 10876 10600 10928 10606
rect 10876 10542 10928 10548
rect 11244 10600 11296 10606
rect 11244 10542 11296 10548
rect 10140 10192 10192 10198
rect 10140 10134 10192 10140
rect 10416 10192 10468 10198
rect 10416 10134 10468 10140
rect 10048 10124 10100 10130
rect 10048 10066 10100 10072
rect 10888 9926 10916 10542
rect 11060 10464 11112 10470
rect 11060 10406 11112 10412
rect 11152 10464 11204 10470
rect 11152 10406 11204 10412
rect 9772 9920 9824 9926
rect 9772 9862 9824 9868
rect 10324 9920 10376 9926
rect 10324 9862 10376 9868
rect 10876 9920 10928 9926
rect 10876 9862 10928 9868
rect 9588 9512 9640 9518
rect 9508 9472 9588 9500
rect 9588 9454 9640 9460
rect 9312 8968 9364 8974
rect 9312 8910 9364 8916
rect 9324 8498 9352 8910
rect 9600 8906 9628 9454
rect 9588 8900 9640 8906
rect 9588 8842 9640 8848
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 9324 7954 9352 8434
rect 9588 8424 9640 8430
rect 9588 8366 9640 8372
rect 9312 7948 9364 7954
rect 9312 7890 9364 7896
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9140 7546 9168 7822
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 9324 6866 9352 7890
rect 9600 7546 9628 8366
rect 9784 7954 9812 9862
rect 10336 9518 10364 9862
rect 10472 9820 10780 9829
rect 10472 9818 10478 9820
rect 10534 9818 10558 9820
rect 10614 9818 10638 9820
rect 10694 9818 10718 9820
rect 10774 9818 10780 9820
rect 10534 9766 10536 9818
rect 10716 9766 10718 9818
rect 10472 9764 10478 9766
rect 10534 9764 10558 9766
rect 10614 9764 10638 9766
rect 10694 9764 10718 9766
rect 10774 9764 10780 9766
rect 10472 9755 10780 9764
rect 11072 9586 11100 10406
rect 11164 9926 11192 10406
rect 11152 9920 11204 9926
rect 11152 9862 11204 9868
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 10324 9512 10376 9518
rect 10324 9454 10376 9460
rect 10876 9104 10928 9110
rect 10876 9046 10928 9052
rect 10324 9036 10376 9042
rect 10324 8978 10376 8984
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 10244 8362 10272 8774
rect 10336 8362 10364 8978
rect 10472 8732 10780 8741
rect 10472 8730 10478 8732
rect 10534 8730 10558 8732
rect 10614 8730 10638 8732
rect 10694 8730 10718 8732
rect 10774 8730 10780 8732
rect 10534 8678 10536 8730
rect 10716 8678 10718 8730
rect 10472 8676 10478 8678
rect 10534 8676 10558 8678
rect 10614 8676 10638 8678
rect 10694 8676 10718 8678
rect 10774 8676 10780 8678
rect 10472 8667 10780 8676
rect 10508 8560 10560 8566
rect 10508 8502 10560 8508
rect 10520 8362 10548 8502
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 10232 8356 10284 8362
rect 10232 8298 10284 8304
rect 10324 8356 10376 8362
rect 10324 8298 10376 8304
rect 10508 8356 10560 8362
rect 10508 8298 10560 8304
rect 9772 7948 9824 7954
rect 9772 7890 9824 7896
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9404 7404 9456 7410
rect 9404 7346 9456 7352
rect 9312 6860 9364 6866
rect 9312 6802 9364 6808
rect 9036 6656 9088 6662
rect 9036 6598 9088 6604
rect 9048 6254 9076 6598
rect 9220 6384 9272 6390
rect 9220 6326 9272 6332
rect 9036 6248 9088 6254
rect 9036 6190 9088 6196
rect 9232 5166 9260 6326
rect 9324 5846 9352 6802
rect 9416 6186 9444 7346
rect 9784 7342 9812 7890
rect 10244 7546 10272 8298
rect 10520 8090 10548 8298
rect 10612 8090 10640 8366
rect 10508 8084 10560 8090
rect 10508 8026 10560 8032
rect 10600 8084 10652 8090
rect 10600 8026 10652 8032
rect 10888 7954 10916 9046
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11164 8362 11192 8570
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 10876 7948 10928 7954
rect 10876 7890 10928 7896
rect 10472 7644 10780 7653
rect 10472 7642 10478 7644
rect 10534 7642 10558 7644
rect 10614 7642 10638 7644
rect 10694 7642 10718 7644
rect 10774 7642 10780 7644
rect 10534 7590 10536 7642
rect 10716 7590 10718 7642
rect 10472 7588 10478 7590
rect 10534 7588 10558 7590
rect 10614 7588 10638 7590
rect 10694 7588 10718 7590
rect 10774 7588 10780 7590
rect 10472 7579 10780 7588
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 9680 7336 9732 7342
rect 9680 7278 9732 7284
rect 9772 7336 9824 7342
rect 9772 7278 9824 7284
rect 9692 7206 9720 7278
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 10324 7200 10376 7206
rect 10324 7142 10376 7148
rect 9956 6452 10008 6458
rect 9956 6394 10008 6400
rect 9968 6254 9996 6394
rect 10336 6390 10364 7142
rect 10472 6556 10780 6565
rect 10472 6554 10478 6556
rect 10534 6554 10558 6556
rect 10614 6554 10638 6556
rect 10694 6554 10718 6556
rect 10774 6554 10780 6556
rect 10534 6502 10536 6554
rect 10716 6502 10718 6554
rect 10472 6500 10478 6502
rect 10534 6500 10558 6502
rect 10614 6500 10638 6502
rect 10694 6500 10718 6502
rect 10774 6500 10780 6502
rect 10472 6491 10780 6500
rect 10324 6384 10376 6390
rect 10324 6326 10376 6332
rect 9864 6248 9916 6254
rect 9864 6190 9916 6196
rect 9956 6248 10008 6254
rect 9956 6190 10008 6196
rect 10048 6248 10100 6254
rect 10048 6190 10100 6196
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 9404 6180 9456 6186
rect 9404 6122 9456 6128
rect 9876 6118 9904 6190
rect 9864 6112 9916 6118
rect 9864 6054 9916 6060
rect 10060 5914 10088 6190
rect 10520 5914 10548 6190
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 10508 5908 10560 5914
rect 10508 5850 10560 5856
rect 9312 5840 9364 5846
rect 9312 5782 9364 5788
rect 10140 5772 10192 5778
rect 10140 5714 10192 5720
rect 9220 5160 9272 5166
rect 9220 5102 9272 5108
rect 9404 4480 9456 4486
rect 9404 4422 9456 4428
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9416 4146 9444 4422
rect 9404 4140 9456 4146
rect 9404 4082 9456 4088
rect 9036 4072 9088 4078
rect 8956 4032 9036 4060
rect 8760 4014 8812 4020
rect 9036 4014 9088 4020
rect 7852 3670 7880 4014
rect 8036 3738 8064 4014
rect 8024 3732 8076 3738
rect 8024 3674 8076 3680
rect 7840 3664 7892 3670
rect 7840 3606 7892 3612
rect 7748 2984 7800 2990
rect 7852 2972 7880 3606
rect 8024 3392 8076 3398
rect 8024 3334 8076 3340
rect 8036 3126 8064 3334
rect 8024 3120 8076 3126
rect 8024 3062 8076 3068
rect 7932 2984 7984 2990
rect 7852 2944 7932 2972
rect 7748 2926 7800 2932
rect 7932 2926 7984 2932
rect 7932 2848 7984 2854
rect 7932 2790 7984 2796
rect 7944 2514 7972 2790
rect 8036 2514 8064 3062
rect 8128 2650 8156 4014
rect 8576 4004 8628 4010
rect 8576 3946 8628 3952
rect 8588 3602 8616 3946
rect 8772 3670 8800 4014
rect 9692 3738 9720 4422
rect 10152 3738 10180 5714
rect 10472 5468 10780 5477
rect 10472 5466 10478 5468
rect 10534 5466 10558 5468
rect 10614 5466 10638 5468
rect 10694 5466 10718 5468
rect 10774 5466 10780 5468
rect 10534 5414 10536 5466
rect 10716 5414 10718 5466
rect 10472 5412 10478 5414
rect 10534 5412 10558 5414
rect 10614 5412 10638 5414
rect 10694 5412 10718 5414
rect 10774 5412 10780 5414
rect 10472 5403 10780 5412
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 10796 4826 10824 5102
rect 10784 4820 10836 4826
rect 10784 4762 10836 4768
rect 10472 4380 10780 4389
rect 10472 4378 10478 4380
rect 10534 4378 10558 4380
rect 10614 4378 10638 4380
rect 10694 4378 10718 4380
rect 10774 4378 10780 4380
rect 10534 4326 10536 4378
rect 10716 4326 10718 4378
rect 10472 4324 10478 4326
rect 10534 4324 10558 4326
rect 10614 4324 10638 4326
rect 10694 4324 10718 4326
rect 10774 4324 10780 4326
rect 10472 4315 10780 4324
rect 10888 3942 10916 7890
rect 11256 4808 11284 10542
rect 11348 10198 11376 10746
rect 11624 10266 11652 11154
rect 11900 10266 11928 11290
rect 11612 10260 11664 10266
rect 11612 10202 11664 10208
rect 11888 10260 11940 10266
rect 11888 10202 11940 10208
rect 11336 10192 11388 10198
rect 11336 10134 11388 10140
rect 11992 10130 12020 12260
rect 12164 12242 12216 12248
rect 12268 12102 12296 12378
rect 12452 12322 12480 12650
rect 12360 12294 12480 12322
rect 12256 12096 12308 12102
rect 12256 12038 12308 12044
rect 12256 10736 12308 10742
rect 12084 10684 12256 10690
rect 12084 10678 12308 10684
rect 12084 10662 12296 10678
rect 12084 10538 12112 10662
rect 12164 10600 12216 10606
rect 12162 10568 12164 10577
rect 12216 10568 12218 10577
rect 12072 10532 12124 10538
rect 12162 10503 12218 10512
rect 12072 10474 12124 10480
rect 12256 10464 12308 10470
rect 12256 10406 12308 10412
rect 11888 10124 11940 10130
rect 11888 10066 11940 10072
rect 11980 10124 12032 10130
rect 11980 10066 12032 10072
rect 11704 9512 11756 9518
rect 11704 9454 11756 9460
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 11348 9110 11376 9318
rect 11336 9104 11388 9110
rect 11336 9046 11388 9052
rect 11716 8634 11744 9454
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 11900 8362 11928 10066
rect 11992 9518 12020 10066
rect 12268 9926 12296 10406
rect 12360 10198 12388 12294
rect 12544 11694 12572 12940
rect 12624 12922 12676 12928
rect 12808 12980 12860 12986
rect 12808 12922 12860 12928
rect 12912 12714 12940 13670
rect 13004 12714 13032 13738
rect 13084 13320 13136 13326
rect 13084 13262 13136 13268
rect 13096 12918 13124 13262
rect 13084 12912 13136 12918
rect 13084 12854 13136 12860
rect 13096 12782 13124 12854
rect 13084 12776 13136 12782
rect 13084 12718 13136 12724
rect 12900 12708 12952 12714
rect 12900 12650 12952 12656
rect 12992 12708 13044 12714
rect 12992 12650 13044 12656
rect 12716 12300 12768 12306
rect 12716 12242 12768 12248
rect 12728 11898 12756 12242
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 12532 11688 12584 11694
rect 12532 11630 12584 11636
rect 12912 11626 12940 12650
rect 13004 11626 13032 12650
rect 13084 12640 13136 12646
rect 13084 12582 13136 12588
rect 12900 11620 12952 11626
rect 12900 11562 12952 11568
rect 12992 11620 13044 11626
rect 12992 11562 13044 11568
rect 12532 11552 12584 11558
rect 12532 11494 12584 11500
rect 12544 11354 12572 11494
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 12900 11008 12952 11014
rect 12900 10950 12952 10956
rect 12912 10674 12940 10950
rect 13004 10810 13032 11562
rect 12992 10804 13044 10810
rect 12992 10746 13044 10752
rect 13004 10674 13032 10746
rect 12808 10668 12860 10674
rect 12808 10610 12860 10616
rect 12900 10668 12952 10674
rect 12900 10610 12952 10616
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 12438 10568 12494 10577
rect 12438 10503 12494 10512
rect 12348 10192 12400 10198
rect 12348 10134 12400 10140
rect 12346 10024 12402 10033
rect 12346 9959 12402 9968
rect 12256 9920 12308 9926
rect 12256 9862 12308 9868
rect 12072 9648 12124 9654
rect 12070 9616 12072 9625
rect 12164 9648 12216 9654
rect 12124 9616 12126 9625
rect 12164 9590 12216 9596
rect 12070 9551 12126 9560
rect 12176 9518 12204 9590
rect 12360 9586 12388 9959
rect 12452 9722 12480 10503
rect 12820 10198 12848 10610
rect 12808 10192 12860 10198
rect 12808 10134 12860 10140
rect 12992 10124 13044 10130
rect 12992 10066 13044 10072
rect 12532 10056 12584 10062
rect 12532 9998 12584 10004
rect 12622 10024 12678 10033
rect 12440 9716 12492 9722
rect 12440 9658 12492 9664
rect 12348 9580 12400 9586
rect 12348 9522 12400 9528
rect 12452 9518 12480 9658
rect 11980 9512 12032 9518
rect 11980 9454 12032 9460
rect 12164 9512 12216 9518
rect 12164 9454 12216 9460
rect 12440 9512 12492 9518
rect 12440 9454 12492 9460
rect 11980 9376 12032 9382
rect 11980 9318 12032 9324
rect 11888 8356 11940 8362
rect 11888 8298 11940 8304
rect 11336 7744 11388 7750
rect 11336 7686 11388 7692
rect 11348 7342 11376 7686
rect 11336 7336 11388 7342
rect 11336 7278 11388 7284
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 11704 7200 11756 7206
rect 11704 7142 11756 7148
rect 11348 6934 11376 7142
rect 11716 7002 11744 7142
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 11336 6928 11388 6934
rect 11336 6870 11388 6876
rect 11520 6860 11572 6866
rect 11520 6802 11572 6808
rect 11532 6458 11560 6802
rect 11520 6452 11572 6458
rect 11520 6394 11572 6400
rect 11532 6254 11560 6394
rect 11520 6248 11572 6254
rect 11520 6190 11572 6196
rect 11796 6248 11848 6254
rect 11796 6190 11848 6196
rect 11808 5914 11836 6190
rect 11796 5908 11848 5914
rect 11796 5850 11848 5856
rect 11808 5370 11836 5850
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 11888 5296 11940 5302
rect 11888 5238 11940 5244
rect 11336 5092 11388 5098
rect 11336 5034 11388 5040
rect 11164 4780 11284 4808
rect 11164 4690 11192 4780
rect 11152 4684 11204 4690
rect 11152 4626 11204 4632
rect 11244 4684 11296 4690
rect 11348 4672 11376 5034
rect 11900 4758 11928 5238
rect 11992 5166 12020 9318
rect 12176 9178 12204 9454
rect 12164 9172 12216 9178
rect 12164 9114 12216 9120
rect 12544 8922 12572 9998
rect 12622 9959 12678 9968
rect 12636 9081 12664 9959
rect 12900 9920 12952 9926
rect 12900 9862 12952 9868
rect 12912 9518 12940 9862
rect 13004 9518 13032 10066
rect 13096 9586 13124 12582
rect 13188 10130 13216 14214
rect 13280 14074 13308 14214
rect 13268 14068 13320 14074
rect 13268 14010 13320 14016
rect 13360 13864 13412 13870
rect 13360 13806 13412 13812
rect 13372 13462 13400 13806
rect 13464 13530 13492 14214
rect 13726 13968 13782 13977
rect 14200 13938 14228 14894
rect 14292 14414 14320 14894
rect 14844 14890 14872 15030
rect 15212 14890 15240 15438
rect 14832 14884 14884 14890
rect 14832 14826 14884 14832
rect 15200 14884 15252 14890
rect 15200 14826 15252 14832
rect 14556 14476 14608 14482
rect 14556 14418 14608 14424
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 14292 13938 14320 14350
rect 14568 14074 14596 14418
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 14556 14068 14608 14074
rect 14556 14010 14608 14016
rect 13726 13903 13782 13912
rect 14188 13932 14240 13938
rect 13740 13870 13768 13903
rect 14188 13874 14240 13880
rect 14280 13932 14332 13938
rect 14280 13874 14332 13880
rect 13728 13864 13780 13870
rect 13728 13806 13780 13812
rect 13452 13524 13504 13530
rect 13452 13466 13504 13472
rect 13360 13456 13412 13462
rect 13360 13398 13412 13404
rect 13452 12776 13504 12782
rect 13452 12718 13504 12724
rect 13464 12442 13492 12718
rect 13452 12436 13504 12442
rect 13452 12378 13504 12384
rect 13464 11898 13492 12378
rect 13636 12164 13688 12170
rect 13636 12106 13688 12112
rect 13268 11892 13320 11898
rect 13268 11834 13320 11840
rect 13452 11892 13504 11898
rect 13452 11834 13504 11840
rect 13280 10606 13308 11834
rect 13648 11626 13676 12106
rect 13636 11620 13688 11626
rect 13636 11562 13688 11568
rect 13636 11280 13688 11286
rect 13636 11222 13688 11228
rect 13452 11212 13504 11218
rect 13452 11154 13504 11160
rect 13464 10810 13492 11154
rect 13452 10804 13504 10810
rect 13452 10746 13504 10752
rect 13268 10600 13320 10606
rect 13268 10542 13320 10548
rect 13280 10198 13308 10542
rect 13268 10192 13320 10198
rect 13268 10134 13320 10140
rect 13176 10124 13228 10130
rect 13176 10066 13228 10072
rect 13268 9920 13320 9926
rect 13268 9862 13320 9868
rect 13176 9716 13228 9722
rect 13176 9658 13228 9664
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 13188 9518 13216 9658
rect 13280 9518 13308 9862
rect 13648 9518 13676 11222
rect 12900 9512 12952 9518
rect 12900 9454 12952 9460
rect 12992 9512 13044 9518
rect 12992 9454 13044 9460
rect 13176 9512 13228 9518
rect 13176 9454 13228 9460
rect 13268 9512 13320 9518
rect 13268 9454 13320 9460
rect 13636 9512 13688 9518
rect 13636 9454 13688 9460
rect 13004 9382 13032 9454
rect 12716 9376 12768 9382
rect 12716 9318 12768 9324
rect 12808 9376 12860 9382
rect 12808 9318 12860 9324
rect 12992 9376 13044 9382
rect 12992 9318 13044 9324
rect 12622 9072 12678 9081
rect 12622 9007 12678 9016
rect 12268 8894 12572 8922
rect 12268 8430 12296 8894
rect 12348 8832 12400 8838
rect 12348 8774 12400 8780
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12360 8430 12388 8774
rect 12256 8424 12308 8430
rect 12256 8366 12308 8372
rect 12348 8424 12400 8430
rect 12348 8366 12400 8372
rect 12348 7880 12400 7886
rect 12348 7822 12400 7828
rect 12256 7812 12308 7818
rect 12256 7754 12308 7760
rect 12072 7744 12124 7750
rect 12072 7686 12124 7692
rect 12084 7342 12112 7686
rect 12268 7478 12296 7754
rect 12256 7472 12308 7478
rect 12256 7414 12308 7420
rect 12072 7336 12124 7342
rect 12072 7278 12124 7284
rect 12164 6792 12216 6798
rect 12164 6734 12216 6740
rect 12176 6118 12204 6734
rect 12268 6254 12296 7414
rect 12360 7274 12388 7822
rect 12348 7268 12400 7274
rect 12348 7210 12400 7216
rect 12360 6798 12388 7210
rect 12348 6792 12400 6798
rect 12348 6734 12400 6740
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 12360 6390 12388 6598
rect 12348 6384 12400 6390
rect 12348 6326 12400 6332
rect 12256 6248 12308 6254
rect 12256 6190 12308 6196
rect 12348 6248 12400 6254
rect 12348 6190 12400 6196
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 12360 5914 12388 6190
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 12452 5386 12480 8774
rect 12532 7336 12584 7342
rect 12532 7278 12584 7284
rect 12544 7002 12572 7278
rect 12532 6996 12584 7002
rect 12532 6938 12584 6944
rect 12532 6860 12584 6866
rect 12532 6802 12584 6808
rect 12544 6458 12572 6802
rect 12532 6452 12584 6458
rect 12532 6394 12584 6400
rect 12532 5568 12584 5574
rect 12532 5510 12584 5516
rect 12360 5358 12480 5386
rect 12360 5302 12388 5358
rect 12348 5296 12400 5302
rect 12348 5238 12400 5244
rect 12544 5166 12572 5510
rect 12728 5166 12756 9318
rect 12820 9042 12848 9318
rect 12808 9036 12860 9042
rect 12808 8978 12860 8984
rect 13004 8430 13032 9318
rect 13084 9036 13136 9042
rect 13084 8978 13136 8984
rect 13096 8634 13124 8978
rect 13188 8974 13216 9454
rect 13544 9376 13596 9382
rect 13544 9318 13596 9324
rect 13556 9178 13584 9318
rect 13544 9172 13596 9178
rect 13544 9114 13596 9120
rect 13176 8968 13228 8974
rect 13176 8910 13228 8916
rect 13084 8628 13136 8634
rect 13084 8570 13136 8576
rect 13648 8498 13676 9454
rect 13740 8566 13768 13806
rect 13830 13628 14138 13637
rect 13830 13626 13836 13628
rect 13892 13626 13916 13628
rect 13972 13626 13996 13628
rect 14052 13626 14076 13628
rect 14132 13626 14138 13628
rect 13892 13574 13894 13626
rect 14074 13574 14076 13626
rect 13830 13572 13836 13574
rect 13892 13572 13916 13574
rect 13972 13572 13996 13574
rect 14052 13572 14076 13574
rect 14132 13572 14138 13574
rect 13830 13563 14138 13572
rect 14200 13462 14228 13874
rect 14372 13524 14424 13530
rect 14372 13466 14424 13472
rect 14188 13456 14240 13462
rect 14188 13398 14240 13404
rect 14280 13184 14332 13190
rect 14280 13126 14332 13132
rect 14188 12708 14240 12714
rect 14188 12650 14240 12656
rect 13830 12540 14138 12549
rect 13830 12538 13836 12540
rect 13892 12538 13916 12540
rect 13972 12538 13996 12540
rect 14052 12538 14076 12540
rect 14132 12538 14138 12540
rect 13892 12486 13894 12538
rect 14074 12486 14076 12538
rect 13830 12484 13836 12486
rect 13892 12484 13916 12486
rect 13972 12484 13996 12486
rect 14052 12484 14076 12486
rect 14132 12484 14138 12486
rect 13830 12475 14138 12484
rect 14200 12442 14228 12650
rect 14292 12442 14320 13126
rect 14188 12436 14240 12442
rect 14188 12378 14240 12384
rect 14280 12436 14332 12442
rect 14280 12378 14332 12384
rect 14280 12300 14332 12306
rect 14280 12242 14332 12248
rect 13830 11452 14138 11461
rect 13830 11450 13836 11452
rect 13892 11450 13916 11452
rect 13972 11450 13996 11452
rect 14052 11450 14076 11452
rect 14132 11450 14138 11452
rect 13892 11398 13894 11450
rect 14074 11398 14076 11450
rect 13830 11396 13836 11398
rect 13892 11396 13916 11398
rect 13972 11396 13996 11398
rect 14052 11396 14076 11398
rect 14132 11396 14138 11398
rect 13830 11387 14138 11396
rect 14292 11286 14320 12242
rect 14384 11558 14412 13466
rect 14476 12306 14504 14010
rect 14648 13932 14700 13938
rect 14648 13874 14700 13880
rect 14556 13796 14608 13802
rect 14556 13738 14608 13744
rect 14568 13462 14596 13738
rect 14556 13456 14608 13462
rect 14556 13398 14608 13404
rect 14464 12300 14516 12306
rect 14464 12242 14516 12248
rect 14568 11694 14596 13398
rect 14660 12782 14688 13874
rect 14648 12776 14700 12782
rect 14648 12718 14700 12724
rect 14844 12374 14872 14826
rect 15580 14550 15608 15506
rect 15568 14544 15620 14550
rect 15568 14486 15620 14492
rect 15016 14272 15068 14278
rect 15016 14214 15068 14220
rect 15028 14074 15056 14214
rect 15016 14068 15068 14074
rect 15016 14010 15068 14016
rect 15028 13734 15056 14010
rect 15108 14000 15160 14006
rect 15108 13942 15160 13948
rect 15120 13870 15148 13942
rect 15108 13864 15160 13870
rect 15108 13806 15160 13812
rect 15016 13728 15068 13734
rect 15200 13728 15252 13734
rect 15016 13670 15068 13676
rect 15120 13688 15200 13716
rect 15120 13530 15148 13688
rect 15200 13670 15252 13676
rect 15108 13524 15160 13530
rect 15108 13466 15160 13472
rect 16040 13394 16068 25774
rect 16212 24268 16264 24274
rect 16212 24210 16264 24216
rect 16224 22137 16252 24210
rect 16396 24200 16448 24206
rect 16396 24142 16448 24148
rect 16304 23588 16356 23594
rect 16304 23530 16356 23536
rect 16316 23186 16344 23530
rect 16304 23180 16356 23186
rect 16304 23122 16356 23128
rect 16408 23050 16436 24142
rect 16488 24064 16540 24070
rect 16488 24006 16540 24012
rect 16396 23044 16448 23050
rect 16396 22986 16448 22992
rect 16408 22710 16436 22986
rect 16396 22704 16448 22710
rect 16396 22646 16448 22652
rect 16210 22128 16266 22137
rect 16500 22094 16528 24006
rect 16592 23254 16620 25774
rect 16776 25758 16896 25786
rect 16672 23316 16724 23322
rect 16672 23258 16724 23264
rect 16580 23248 16632 23254
rect 16580 23190 16632 23196
rect 16592 22778 16620 23190
rect 16580 22772 16632 22778
rect 16580 22714 16632 22720
rect 16684 22234 16712 23258
rect 16672 22228 16724 22234
rect 16672 22170 16724 22176
rect 16210 22063 16266 22072
rect 16408 22066 16528 22094
rect 16120 21956 16172 21962
rect 16120 21898 16172 21904
rect 16132 21486 16160 21898
rect 16120 21480 16172 21486
rect 16212 21480 16264 21486
rect 16120 21422 16172 21428
rect 16210 21448 16212 21457
rect 16264 21448 16266 21457
rect 16132 19394 16160 21422
rect 16210 21383 16266 21392
rect 16408 21350 16436 22066
rect 16488 21888 16540 21894
rect 16488 21830 16540 21836
rect 16396 21344 16448 21350
rect 16396 21286 16448 21292
rect 16212 21004 16264 21010
rect 16212 20946 16264 20952
rect 16224 19514 16252 20946
rect 16304 20800 16356 20806
rect 16304 20742 16356 20748
rect 16316 20398 16344 20742
rect 16304 20392 16356 20398
rect 16304 20334 16356 20340
rect 16500 19854 16528 21830
rect 16488 19848 16540 19854
rect 16488 19790 16540 19796
rect 16212 19508 16264 19514
rect 16212 19450 16264 19456
rect 16132 19366 16252 19394
rect 16120 19304 16172 19310
rect 16120 19246 16172 19252
rect 16132 18698 16160 19246
rect 16120 18692 16172 18698
rect 16120 18634 16172 18640
rect 16132 18193 16160 18634
rect 16118 18184 16174 18193
rect 16118 18119 16120 18128
rect 16172 18119 16174 18128
rect 16120 18090 16172 18096
rect 16224 14958 16252 19366
rect 16304 18352 16356 18358
rect 16304 18294 16356 18300
rect 16316 18222 16344 18294
rect 16304 18216 16356 18222
rect 16304 18158 16356 18164
rect 16500 16658 16528 19790
rect 16684 19530 16712 22170
rect 16776 22098 16804 25758
rect 16960 24614 16988 26318
rect 17052 25294 17080 27406
rect 17144 27402 17172 28070
rect 17604 27606 17632 28562
rect 17592 27600 17644 27606
rect 17592 27542 17644 27548
rect 17132 27396 17184 27402
rect 17132 27338 17184 27344
rect 17188 27228 17496 27237
rect 17188 27226 17194 27228
rect 17250 27226 17274 27228
rect 17330 27226 17354 27228
rect 17410 27226 17434 27228
rect 17490 27226 17496 27228
rect 17250 27174 17252 27226
rect 17432 27174 17434 27226
rect 17188 27172 17194 27174
rect 17250 27172 17274 27174
rect 17330 27172 17354 27174
rect 17410 27172 17434 27174
rect 17490 27172 17496 27174
rect 17188 27163 17496 27172
rect 17132 26920 17184 26926
rect 17132 26862 17184 26868
rect 17144 26314 17172 26862
rect 17500 26852 17552 26858
rect 17500 26794 17552 26800
rect 17132 26308 17184 26314
rect 17132 26250 17184 26256
rect 17512 26234 17540 26794
rect 17512 26206 17632 26234
rect 17188 26140 17496 26149
rect 17188 26138 17194 26140
rect 17250 26138 17274 26140
rect 17330 26138 17354 26140
rect 17410 26138 17434 26140
rect 17490 26138 17496 26140
rect 17250 26086 17252 26138
rect 17432 26086 17434 26138
rect 17188 26084 17194 26086
rect 17250 26084 17274 26086
rect 17330 26084 17354 26086
rect 17410 26084 17434 26086
rect 17490 26084 17496 26086
rect 17188 26075 17496 26084
rect 17604 25945 17632 26206
rect 17590 25936 17646 25945
rect 17590 25871 17646 25880
rect 17696 25786 17724 30552
rect 17776 30534 17828 30540
rect 18064 30326 18092 30738
rect 18800 30682 18828 30738
rect 18708 30654 18828 30682
rect 18708 30598 18736 30654
rect 18696 30592 18748 30598
rect 18696 30534 18748 30540
rect 18052 30320 18104 30326
rect 18052 30262 18104 30268
rect 18512 30184 18564 30190
rect 18512 30126 18564 30132
rect 18524 29850 18552 30126
rect 18512 29844 18564 29850
rect 18512 29786 18564 29792
rect 18512 29164 18564 29170
rect 18512 29106 18564 29112
rect 18420 28620 18472 28626
rect 18420 28562 18472 28568
rect 17868 28416 17920 28422
rect 17868 28358 17920 28364
rect 17776 27532 17828 27538
rect 17776 27474 17828 27480
rect 17788 27441 17816 27474
rect 17774 27432 17830 27441
rect 17774 27367 17830 27376
rect 17776 26920 17828 26926
rect 17776 26862 17828 26868
rect 17788 25820 17816 26862
rect 17880 26450 17908 28358
rect 18432 28218 18460 28562
rect 18420 28212 18472 28218
rect 18420 28154 18472 28160
rect 18420 28008 18472 28014
rect 18420 27950 18472 27956
rect 18328 27940 18380 27946
rect 18328 27882 18380 27888
rect 17960 27532 18012 27538
rect 17960 27474 18012 27480
rect 17972 27130 18000 27474
rect 17960 27124 18012 27130
rect 17960 27066 18012 27072
rect 18340 27062 18368 27882
rect 18328 27056 18380 27062
rect 18328 26998 18380 27004
rect 18144 26920 18196 26926
rect 18144 26862 18196 26868
rect 17958 26480 18014 26489
rect 17868 26444 17920 26450
rect 17958 26415 18014 26424
rect 18156 26432 18184 26862
rect 18236 26852 18288 26858
rect 18236 26794 18288 26800
rect 18248 26761 18276 26794
rect 18234 26752 18290 26761
rect 18234 26687 18290 26696
rect 18236 26444 18288 26450
rect 17868 26386 17920 26392
rect 17972 26382 18000 26415
rect 18156 26404 18236 26432
rect 17960 26376 18012 26382
rect 17960 26318 18012 26324
rect 18156 25838 18184 26404
rect 18340 26432 18368 26998
rect 18432 26926 18460 27950
rect 18420 26920 18472 26926
rect 18420 26862 18472 26868
rect 18432 26450 18460 26862
rect 18524 26761 18552 29106
rect 18708 28098 18736 30534
rect 18880 29708 18932 29714
rect 18880 29650 18932 29656
rect 18892 29306 18920 29650
rect 18880 29300 18932 29306
rect 18880 29242 18932 29248
rect 18984 29170 19012 30756
rect 19116 30767 19118 30776
rect 19064 30738 19116 30744
rect 18972 29164 19024 29170
rect 18892 29124 18972 29152
rect 18788 28620 18840 28626
rect 18788 28562 18840 28568
rect 18800 28218 18828 28562
rect 18788 28212 18840 28218
rect 18788 28154 18840 28160
rect 18708 28070 18828 28098
rect 18696 27532 18748 27538
rect 18696 27474 18748 27480
rect 18510 26752 18566 26761
rect 18510 26687 18566 26696
rect 18288 26404 18368 26432
rect 18420 26444 18472 26450
rect 18236 26386 18288 26392
rect 18420 26386 18472 26392
rect 18236 26308 18288 26314
rect 18236 26250 18288 26256
rect 18248 25838 18276 26250
rect 18432 25906 18460 26386
rect 18420 25900 18472 25906
rect 18420 25842 18472 25848
rect 17868 25832 17920 25838
rect 17788 25792 17868 25820
rect 17604 25758 17724 25786
rect 17868 25774 17920 25780
rect 18144 25832 18196 25838
rect 18144 25774 18196 25780
rect 18236 25832 18288 25838
rect 18236 25774 18288 25780
rect 17040 25288 17092 25294
rect 17040 25230 17092 25236
rect 17052 24750 17080 25230
rect 17188 25052 17496 25061
rect 17188 25050 17194 25052
rect 17250 25050 17274 25052
rect 17330 25050 17354 25052
rect 17410 25050 17434 25052
rect 17490 25050 17496 25052
rect 17250 24998 17252 25050
rect 17432 24998 17434 25050
rect 17188 24996 17194 24998
rect 17250 24996 17274 24998
rect 17330 24996 17354 24998
rect 17410 24996 17434 24998
rect 17490 24996 17496 24998
rect 17188 24987 17496 24996
rect 17040 24744 17092 24750
rect 17040 24686 17092 24692
rect 16948 24608 17000 24614
rect 16948 24550 17000 24556
rect 17408 24608 17460 24614
rect 17408 24550 17460 24556
rect 17420 24410 17448 24550
rect 17408 24404 17460 24410
rect 17408 24346 17460 24352
rect 17604 24154 17632 25758
rect 17684 25696 17736 25702
rect 17684 25638 17736 25644
rect 17696 25430 17724 25638
rect 17684 25424 17736 25430
rect 17684 25366 17736 25372
rect 17776 25288 17828 25294
rect 17776 25230 17828 25236
rect 17684 25152 17736 25158
rect 17684 25094 17736 25100
rect 17696 24886 17724 25094
rect 17788 24886 17816 25230
rect 17684 24880 17736 24886
rect 17684 24822 17736 24828
rect 17776 24880 17828 24886
rect 17776 24822 17828 24828
rect 17604 24126 17724 24154
rect 17592 24064 17644 24070
rect 17592 24006 17644 24012
rect 17188 23964 17496 23973
rect 17188 23962 17194 23964
rect 17250 23962 17274 23964
rect 17330 23962 17354 23964
rect 17410 23962 17434 23964
rect 17490 23962 17496 23964
rect 17250 23910 17252 23962
rect 17432 23910 17434 23962
rect 17188 23908 17194 23910
rect 17250 23908 17274 23910
rect 17330 23908 17354 23910
rect 17410 23908 17434 23910
rect 17490 23908 17496 23910
rect 17188 23899 17496 23908
rect 16856 23656 16908 23662
rect 16856 23598 16908 23604
rect 16868 23322 16896 23598
rect 17604 23322 17632 24006
rect 16856 23316 16908 23322
rect 16856 23258 16908 23264
rect 17592 23316 17644 23322
rect 17592 23258 17644 23264
rect 17696 23254 17724 24126
rect 17788 23730 17816 24822
rect 17880 24732 17908 25774
rect 17960 25764 18012 25770
rect 17960 25706 18012 25712
rect 17972 25673 18000 25706
rect 17958 25664 18014 25673
rect 17958 25599 18014 25608
rect 18156 24886 18184 25774
rect 18144 24880 18196 24886
rect 18144 24822 18196 24828
rect 17960 24744 18012 24750
rect 17880 24704 17960 24732
rect 17960 24686 18012 24692
rect 17776 23724 17828 23730
rect 17776 23666 17828 23672
rect 17684 23248 17736 23254
rect 17684 23190 17736 23196
rect 17188 22876 17496 22885
rect 17188 22874 17194 22876
rect 17250 22874 17274 22876
rect 17330 22874 17354 22876
rect 17410 22874 17434 22876
rect 17490 22874 17496 22876
rect 17250 22822 17252 22874
rect 17432 22822 17434 22874
rect 17188 22820 17194 22822
rect 17250 22820 17274 22822
rect 17330 22820 17354 22822
rect 17410 22820 17434 22822
rect 17490 22820 17496 22822
rect 17188 22811 17496 22820
rect 17972 22642 18000 24686
rect 18420 24676 18472 24682
rect 18420 24618 18472 24624
rect 18144 24200 18196 24206
rect 18144 24142 18196 24148
rect 18156 23866 18184 24142
rect 18144 23860 18196 23866
rect 18144 23802 18196 23808
rect 18328 23656 18380 23662
rect 18328 23598 18380 23604
rect 18340 23322 18368 23598
rect 18328 23316 18380 23322
rect 18328 23258 18380 23264
rect 18144 23180 18196 23186
rect 18144 23122 18196 23128
rect 17960 22636 18012 22642
rect 17960 22578 18012 22584
rect 17776 22568 17828 22574
rect 17776 22510 17828 22516
rect 16948 22500 17000 22506
rect 16948 22442 17000 22448
rect 17224 22500 17276 22506
rect 17224 22442 17276 22448
rect 16764 22092 16816 22098
rect 16960 22094 16988 22442
rect 17040 22160 17092 22166
rect 17040 22102 17092 22108
rect 16764 22034 16816 22040
rect 16868 22066 16988 22094
rect 16868 21622 16896 22066
rect 16856 21616 16908 21622
rect 16856 21558 16908 21564
rect 16868 19802 16896 21558
rect 17052 21049 17080 22102
rect 17236 21894 17264 22442
rect 17788 22166 17816 22510
rect 17776 22160 17828 22166
rect 18156 22137 18184 23122
rect 17776 22102 17828 22108
rect 18142 22128 18198 22137
rect 18432 22094 18460 24618
rect 18142 22063 18198 22072
rect 18340 22066 18460 22094
rect 17774 21992 17830 22001
rect 17774 21927 17776 21936
rect 17828 21927 17830 21936
rect 17776 21898 17828 21904
rect 17224 21888 17276 21894
rect 17224 21830 17276 21836
rect 17188 21788 17496 21797
rect 17188 21786 17194 21788
rect 17250 21786 17274 21788
rect 17330 21786 17354 21788
rect 17410 21786 17434 21788
rect 17490 21786 17496 21788
rect 17250 21734 17252 21786
rect 17432 21734 17434 21786
rect 17188 21732 17194 21734
rect 17250 21732 17274 21734
rect 17330 21732 17354 21734
rect 17410 21732 17434 21734
rect 17490 21732 17496 21734
rect 17188 21723 17496 21732
rect 17408 21412 17460 21418
rect 17408 21354 17460 21360
rect 17960 21412 18012 21418
rect 17960 21354 18012 21360
rect 17420 21146 17448 21354
rect 17408 21140 17460 21146
rect 17408 21082 17460 21088
rect 17038 21040 17094 21049
rect 17972 21010 18000 21354
rect 17038 20975 17040 20984
rect 17092 20975 17094 20984
rect 17684 21004 17736 21010
rect 17040 20946 17092 20952
rect 17684 20946 17736 20952
rect 17776 21004 17828 21010
rect 17776 20946 17828 20952
rect 17960 21004 18012 21010
rect 17960 20946 18012 20952
rect 17188 20700 17496 20709
rect 17188 20698 17194 20700
rect 17250 20698 17274 20700
rect 17330 20698 17354 20700
rect 17410 20698 17434 20700
rect 17490 20698 17496 20700
rect 17250 20646 17252 20698
rect 17432 20646 17434 20698
rect 17188 20644 17194 20646
rect 17250 20644 17274 20646
rect 17330 20644 17354 20646
rect 17410 20644 17434 20646
rect 17490 20644 17496 20646
rect 17188 20635 17496 20644
rect 17592 19916 17644 19922
rect 17592 19858 17644 19864
rect 16868 19774 17080 19802
rect 16856 19712 16908 19718
rect 16856 19654 16908 19660
rect 16592 19502 16712 19530
rect 16592 18290 16620 19502
rect 16868 19310 16896 19654
rect 16856 19304 16908 19310
rect 16762 19272 16818 19281
rect 16856 19246 16908 19252
rect 16762 19207 16818 19216
rect 16672 18828 16724 18834
rect 16672 18770 16724 18776
rect 16684 18426 16712 18770
rect 16672 18420 16724 18426
rect 16672 18362 16724 18368
rect 16580 18284 16632 18290
rect 16580 18226 16632 18232
rect 16776 17626 16804 19207
rect 16948 17740 17000 17746
rect 16948 17682 17000 17688
rect 16592 17598 16804 17626
rect 16856 17604 16908 17610
rect 16488 16652 16540 16658
rect 16488 16594 16540 16600
rect 16592 15638 16620 17598
rect 16856 17546 16908 17552
rect 16764 17536 16816 17542
rect 16764 17478 16816 17484
rect 16672 17332 16724 17338
rect 16672 17274 16724 17280
rect 16684 16726 16712 17274
rect 16672 16720 16724 16726
rect 16672 16662 16724 16668
rect 16580 15632 16632 15638
rect 16580 15574 16632 15580
rect 16212 14952 16264 14958
rect 16212 14894 16264 14900
rect 16304 14408 16356 14414
rect 16304 14350 16356 14356
rect 16120 14272 16172 14278
rect 16120 14214 16172 14220
rect 16132 14074 16160 14214
rect 16120 14068 16172 14074
rect 16120 14010 16172 14016
rect 16212 13728 16264 13734
rect 16212 13670 16264 13676
rect 16224 13462 16252 13670
rect 16212 13456 16264 13462
rect 16212 13398 16264 13404
rect 15660 13388 15712 13394
rect 15660 13330 15712 13336
rect 16028 13388 16080 13394
rect 16028 13330 16080 13336
rect 15384 13320 15436 13326
rect 15384 13262 15436 13268
rect 15396 12646 15424 13262
rect 15568 13252 15620 13258
rect 15568 13194 15620 13200
rect 15476 13184 15528 13190
rect 15476 13126 15528 13132
rect 15488 12714 15516 13126
rect 15580 12986 15608 13194
rect 15568 12980 15620 12986
rect 15568 12922 15620 12928
rect 15476 12708 15528 12714
rect 15476 12650 15528 12656
rect 15384 12640 15436 12646
rect 15384 12582 15436 12588
rect 14832 12368 14884 12374
rect 14832 12310 14884 12316
rect 15580 12238 15608 12922
rect 15672 12442 15700 13330
rect 15844 12640 15896 12646
rect 15844 12582 15896 12588
rect 15660 12436 15712 12442
rect 15660 12378 15712 12384
rect 15568 12232 15620 12238
rect 15568 12174 15620 12180
rect 15660 11892 15712 11898
rect 15660 11834 15712 11840
rect 14556 11688 14608 11694
rect 14556 11630 14608 11636
rect 14740 11620 14792 11626
rect 14740 11562 14792 11568
rect 15384 11620 15436 11626
rect 15384 11562 15436 11568
rect 14372 11552 14424 11558
rect 14372 11494 14424 11500
rect 14280 11280 14332 11286
rect 14280 11222 14332 11228
rect 14002 10704 14058 10713
rect 14002 10639 14058 10648
rect 14016 10606 14044 10639
rect 14292 10606 14320 11222
rect 14004 10600 14056 10606
rect 14004 10542 14056 10548
rect 14280 10600 14332 10606
rect 14280 10542 14332 10548
rect 14016 10452 14044 10542
rect 14016 10424 14228 10452
rect 13830 10364 14138 10373
rect 13830 10362 13836 10364
rect 13892 10362 13916 10364
rect 13972 10362 13996 10364
rect 14052 10362 14076 10364
rect 14132 10362 14138 10364
rect 13892 10310 13894 10362
rect 14074 10310 14076 10362
rect 13830 10308 13836 10310
rect 13892 10308 13916 10310
rect 13972 10308 13996 10310
rect 14052 10308 14076 10310
rect 14132 10308 14138 10310
rect 13830 10299 14138 10308
rect 14200 10266 14228 10424
rect 14188 10260 14240 10266
rect 14188 10202 14240 10208
rect 14186 9616 14242 9625
rect 14186 9551 14242 9560
rect 13830 9276 14138 9285
rect 13830 9274 13836 9276
rect 13892 9274 13916 9276
rect 13972 9274 13996 9276
rect 14052 9274 14076 9276
rect 14132 9274 14138 9276
rect 13892 9222 13894 9274
rect 14074 9222 14076 9274
rect 13830 9220 13836 9222
rect 13892 9220 13916 9222
rect 13972 9220 13996 9222
rect 14052 9220 14076 9222
rect 14132 9220 14138 9222
rect 13830 9211 14138 9220
rect 14200 9178 14228 9551
rect 14188 9172 14240 9178
rect 14188 9114 14240 9120
rect 14186 9072 14242 9081
rect 14186 9007 14188 9016
rect 14240 9007 14242 9016
rect 14292 9024 14320 10542
rect 14384 10470 14412 11494
rect 14648 11008 14700 11014
rect 14648 10950 14700 10956
rect 14660 10810 14688 10950
rect 14648 10804 14700 10810
rect 14648 10746 14700 10752
rect 14752 10606 14780 11562
rect 15396 11354 15424 11562
rect 15568 11552 15620 11558
rect 15568 11494 15620 11500
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15384 11348 15436 11354
rect 15384 11290 15436 11296
rect 15304 11150 15332 11290
rect 15580 11218 15608 11494
rect 15568 11212 15620 11218
rect 15568 11154 15620 11160
rect 15292 11144 15344 11150
rect 15292 11086 15344 11092
rect 14740 10600 14792 10606
rect 14740 10542 14792 10548
rect 14556 10532 14608 10538
rect 14556 10474 14608 10480
rect 14372 10464 14424 10470
rect 14372 10406 14424 10412
rect 14384 9450 14412 10406
rect 14568 10062 14596 10474
rect 15304 10198 15332 11086
rect 15672 10606 15700 11834
rect 15856 10606 15884 12582
rect 16040 12238 16068 13330
rect 16120 12708 16172 12714
rect 16120 12650 16172 12656
rect 16028 12232 16080 12238
rect 16028 12174 16080 12180
rect 16132 11218 16160 12650
rect 16224 12306 16252 13398
rect 16212 12300 16264 12306
rect 16212 12242 16264 12248
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 16224 11218 16252 11834
rect 16120 11212 16172 11218
rect 16120 11154 16172 11160
rect 16212 11212 16264 11218
rect 16212 11154 16264 11160
rect 16120 11008 16172 11014
rect 16120 10950 16172 10956
rect 15384 10600 15436 10606
rect 15660 10600 15712 10606
rect 15436 10548 15516 10554
rect 15384 10542 15516 10548
rect 15660 10542 15712 10548
rect 15844 10600 15896 10606
rect 15844 10542 15896 10548
rect 15396 10526 15516 10542
rect 15384 10464 15436 10470
rect 15384 10406 15436 10412
rect 15292 10192 15344 10198
rect 15292 10134 15344 10140
rect 14648 10124 14700 10130
rect 14648 10066 14700 10072
rect 14556 10056 14608 10062
rect 14556 9998 14608 10004
rect 14660 9722 14688 10066
rect 14924 9920 14976 9926
rect 14924 9862 14976 9868
rect 15200 9920 15252 9926
rect 15200 9862 15252 9868
rect 14648 9716 14700 9722
rect 14648 9658 14700 9664
rect 14372 9444 14424 9450
rect 14372 9386 14424 9392
rect 14372 9036 14424 9042
rect 14292 8996 14372 9024
rect 14188 8978 14240 8984
rect 14372 8978 14424 8984
rect 14188 8628 14240 8634
rect 14188 8570 14240 8576
rect 13728 8560 13780 8566
rect 13728 8502 13780 8508
rect 13636 8492 13688 8498
rect 13636 8434 13688 8440
rect 12992 8424 13044 8430
rect 12992 8366 13044 8372
rect 13176 8016 13228 8022
rect 13176 7958 13228 7964
rect 13188 7886 13216 7958
rect 13648 7954 13676 8434
rect 13830 8188 14138 8197
rect 13830 8186 13836 8188
rect 13892 8186 13916 8188
rect 13972 8186 13996 8188
rect 14052 8186 14076 8188
rect 14132 8186 14138 8188
rect 13892 8134 13894 8186
rect 14074 8134 14076 8186
rect 13830 8132 13836 8134
rect 13892 8132 13916 8134
rect 13972 8132 13996 8134
rect 14052 8132 14076 8134
rect 14132 8132 14138 8134
rect 13830 8123 14138 8132
rect 13636 7948 13688 7954
rect 13636 7890 13688 7896
rect 13912 7948 13964 7954
rect 13912 7890 13964 7896
rect 13176 7880 13228 7886
rect 13176 7822 13228 7828
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 13188 7546 13216 7822
rect 13176 7540 13228 7546
rect 13176 7482 13228 7488
rect 13084 7200 13136 7206
rect 13084 7142 13136 7148
rect 13096 6866 13124 7142
rect 13372 7002 13400 7822
rect 13924 7546 13952 7890
rect 14004 7744 14056 7750
rect 14004 7686 14056 7692
rect 13912 7540 13964 7546
rect 13912 7482 13964 7488
rect 14016 7410 14044 7686
rect 14200 7546 14228 8570
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14280 8356 14332 8362
rect 14280 8298 14332 8304
rect 14292 8022 14320 8298
rect 14372 8288 14424 8294
rect 14372 8230 14424 8236
rect 14280 8016 14332 8022
rect 14280 7958 14332 7964
rect 14188 7540 14240 7546
rect 14188 7482 14240 7488
rect 14004 7404 14056 7410
rect 14004 7346 14056 7352
rect 14384 7342 14412 8230
rect 14556 7744 14608 7750
rect 14556 7686 14608 7692
rect 14568 7410 14596 7686
rect 14556 7404 14608 7410
rect 14556 7346 14608 7352
rect 14372 7336 14424 7342
rect 14372 7278 14424 7284
rect 13830 7100 14138 7109
rect 13830 7098 13836 7100
rect 13892 7098 13916 7100
rect 13972 7098 13996 7100
rect 14052 7098 14076 7100
rect 14132 7098 14138 7100
rect 13892 7046 13894 7098
rect 14074 7046 14076 7098
rect 13830 7044 13836 7046
rect 13892 7044 13916 7046
rect 13972 7044 13996 7046
rect 14052 7044 14076 7046
rect 14132 7044 14138 7046
rect 13830 7035 14138 7044
rect 13360 6996 13412 7002
rect 13360 6938 13412 6944
rect 13084 6860 13136 6866
rect 13084 6802 13136 6808
rect 14188 6860 14240 6866
rect 14188 6802 14240 6808
rect 13268 6656 13320 6662
rect 13268 6598 13320 6604
rect 13280 6322 13308 6598
rect 13268 6316 13320 6322
rect 13268 6258 13320 6264
rect 13176 6248 13228 6254
rect 13176 6190 13228 6196
rect 13188 5914 13216 6190
rect 13544 6112 13596 6118
rect 13544 6054 13596 6060
rect 13176 5908 13228 5914
rect 13176 5850 13228 5856
rect 13556 5846 13584 6054
rect 13830 6012 14138 6021
rect 13830 6010 13836 6012
rect 13892 6010 13916 6012
rect 13972 6010 13996 6012
rect 14052 6010 14076 6012
rect 14132 6010 14138 6012
rect 13892 5958 13894 6010
rect 14074 5958 14076 6010
rect 13830 5956 13836 5958
rect 13892 5956 13916 5958
rect 13972 5956 13996 5958
rect 14052 5956 14076 5958
rect 14132 5956 14138 5958
rect 13830 5947 14138 5956
rect 14200 5914 14228 6802
rect 14660 6730 14688 8434
rect 14832 8424 14884 8430
rect 14830 8392 14832 8401
rect 14884 8392 14886 8401
rect 14830 8327 14886 8336
rect 14740 8288 14792 8294
rect 14740 8230 14792 8236
rect 14752 7818 14780 8230
rect 14740 7812 14792 7818
rect 14740 7754 14792 7760
rect 14648 6724 14700 6730
rect 14648 6666 14700 6672
rect 14188 5908 14240 5914
rect 14188 5850 14240 5856
rect 13544 5840 13596 5846
rect 13544 5782 13596 5788
rect 14556 5840 14608 5846
rect 14556 5782 14608 5788
rect 14568 5370 14596 5782
rect 14556 5364 14608 5370
rect 14556 5306 14608 5312
rect 11980 5160 12032 5166
rect 11980 5102 12032 5108
rect 12532 5160 12584 5166
rect 12532 5102 12584 5108
rect 12624 5160 12676 5166
rect 12624 5102 12676 5108
rect 12716 5160 12768 5166
rect 12716 5102 12768 5108
rect 13452 5160 13504 5166
rect 13452 5102 13504 5108
rect 13728 5160 13780 5166
rect 13728 5102 13780 5108
rect 11992 4758 12020 5102
rect 12636 4826 12664 5102
rect 12716 5024 12768 5030
rect 12716 4966 12768 4972
rect 12624 4820 12676 4826
rect 12624 4762 12676 4768
rect 12728 4758 12756 4966
rect 11888 4752 11940 4758
rect 11888 4694 11940 4700
rect 11980 4752 12032 4758
rect 11980 4694 12032 4700
rect 12716 4752 12768 4758
rect 12716 4694 12768 4700
rect 11296 4644 11376 4672
rect 11244 4626 11296 4632
rect 11060 4548 11112 4554
rect 11060 4490 11112 4496
rect 11072 4282 11100 4490
rect 11060 4276 11112 4282
rect 11060 4218 11112 4224
rect 11164 4146 11192 4626
rect 11244 4548 11296 4554
rect 11244 4490 11296 4496
rect 11256 4282 11284 4490
rect 11244 4276 11296 4282
rect 11244 4218 11296 4224
rect 11152 4140 11204 4146
rect 11152 4082 11204 4088
rect 11164 4026 11192 4082
rect 10980 3998 11192 4026
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 10876 3936 10928 3942
rect 10876 3878 10928 3884
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 8760 3664 8812 3670
rect 8760 3606 8812 3612
rect 10980 3602 11008 3998
rect 11152 3936 11204 3942
rect 11072 3896 11152 3924
rect 8576 3596 8628 3602
rect 8576 3538 8628 3544
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 10472 3292 10780 3301
rect 10472 3290 10478 3292
rect 10534 3290 10558 3292
rect 10614 3290 10638 3292
rect 10694 3290 10718 3292
rect 10774 3290 10780 3292
rect 10534 3238 10536 3290
rect 10716 3238 10718 3290
rect 10472 3236 10478 3238
rect 10534 3236 10558 3238
rect 10614 3236 10638 3238
rect 10694 3236 10718 3238
rect 10774 3236 10780 3238
rect 10472 3227 10780 3236
rect 10980 3194 11008 3538
rect 11072 3398 11100 3896
rect 11152 3878 11204 3884
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 11060 3392 11112 3398
rect 11060 3334 11112 3340
rect 9956 3188 10008 3194
rect 9956 3130 10008 3136
rect 10968 3188 11020 3194
rect 10968 3130 11020 3136
rect 8300 2984 8352 2990
rect 8300 2926 8352 2932
rect 8116 2644 8168 2650
rect 8116 2586 8168 2592
rect 8312 2514 8340 2926
rect 9968 2922 9996 3130
rect 10232 3120 10284 3126
rect 10232 3062 10284 3068
rect 9956 2916 10008 2922
rect 9956 2858 10008 2864
rect 9680 2848 9732 2854
rect 9680 2790 9732 2796
rect 10140 2848 10192 2854
rect 10140 2790 10192 2796
rect 9692 2514 9720 2790
rect 10152 2514 10180 2790
rect 10244 2514 10272 3062
rect 10980 2990 11008 3130
rect 10968 2984 11020 2990
rect 10968 2926 11020 2932
rect 10968 2848 11020 2854
rect 10968 2790 11020 2796
rect 7564 2508 7616 2514
rect 7564 2450 7616 2456
rect 7932 2508 7984 2514
rect 7932 2450 7984 2456
rect 8024 2508 8076 2514
rect 8024 2450 8076 2456
rect 8300 2508 8352 2514
rect 8300 2450 8352 2456
rect 9496 2508 9548 2514
rect 9496 2450 9548 2456
rect 9680 2508 9732 2514
rect 9680 2450 9732 2456
rect 10140 2508 10192 2514
rect 10140 2450 10192 2456
rect 10232 2508 10284 2514
rect 10232 2450 10284 2456
rect 6920 2440 6972 2446
rect 6920 2382 6972 2388
rect 7012 2440 7064 2446
rect 7012 2382 7064 2388
rect 6932 2122 6960 2382
rect 6840 2094 6960 2122
rect 6552 1896 6604 1902
rect 6552 1838 6604 1844
rect 6644 1828 6696 1834
rect 6644 1770 6696 1776
rect 6656 762 6684 1770
rect 6840 1222 6868 2094
rect 6920 2032 6972 2038
rect 6920 1974 6972 1980
rect 6932 1426 6960 1974
rect 7024 1426 7052 2382
rect 8208 2304 8260 2310
rect 8208 2246 8260 2252
rect 7472 1896 7524 1902
rect 7472 1838 7524 1844
rect 7114 1660 7422 1669
rect 7114 1658 7120 1660
rect 7176 1658 7200 1660
rect 7256 1658 7280 1660
rect 7336 1658 7360 1660
rect 7416 1658 7422 1660
rect 7176 1606 7178 1658
rect 7358 1606 7360 1658
rect 7114 1604 7120 1606
rect 7176 1604 7200 1606
rect 7256 1604 7280 1606
rect 7336 1604 7360 1606
rect 7416 1604 7422 1606
rect 7114 1595 7422 1604
rect 6920 1420 6972 1426
rect 6920 1362 6972 1368
rect 7012 1420 7064 1426
rect 7012 1362 7064 1368
rect 6736 1216 6788 1222
rect 6736 1158 6788 1164
rect 6828 1216 6880 1222
rect 6828 1158 6880 1164
rect 6748 882 6776 1158
rect 6736 876 6788 882
rect 6736 818 6788 824
rect 6656 734 6776 762
rect 6748 400 6776 734
rect 7114 572 7422 581
rect 7114 570 7120 572
rect 7176 570 7200 572
rect 7256 570 7280 572
rect 7336 570 7360 572
rect 7416 570 7422 572
rect 7176 518 7178 570
rect 7358 518 7360 570
rect 7114 516 7120 518
rect 7176 516 7200 518
rect 7256 516 7280 518
rect 7336 516 7360 518
rect 7416 516 7422 518
rect 7114 507 7422 516
rect 7484 456 7512 1838
rect 8220 1426 8248 2246
rect 9036 1896 9088 1902
rect 9036 1838 9088 1844
rect 8392 1556 8444 1562
rect 8392 1498 8444 1504
rect 8208 1420 8260 1426
rect 8208 1362 8260 1368
rect 7932 1352 7984 1358
rect 7932 1294 7984 1300
rect 7944 1018 7972 1294
rect 7932 1012 7984 1018
rect 7932 954 7984 960
rect 7840 808 7892 814
rect 7840 750 7892 756
rect 7300 428 7512 456
rect 7300 400 7328 428
rect 7852 400 7880 750
rect 8404 400 8432 1498
rect 8944 1420 8996 1426
rect 8944 1362 8996 1368
rect 8956 400 8984 1362
rect 9048 1018 9076 1838
rect 9404 1216 9456 1222
rect 9404 1158 9456 1164
rect 9036 1012 9088 1018
rect 9036 954 9088 960
rect 9416 882 9444 1158
rect 9404 876 9456 882
rect 9404 818 9456 824
rect 9508 400 9536 2450
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 9956 2304 10008 2310
rect 9956 2246 10008 2252
rect 10232 2304 10284 2310
rect 10232 2246 10284 2252
rect 9692 814 9720 2246
rect 9968 1426 9996 2246
rect 10244 1970 10272 2246
rect 10472 2204 10780 2213
rect 10472 2202 10478 2204
rect 10534 2202 10558 2204
rect 10614 2202 10638 2204
rect 10694 2202 10718 2204
rect 10774 2202 10780 2204
rect 10534 2150 10536 2202
rect 10716 2150 10718 2202
rect 10472 2148 10478 2150
rect 10534 2148 10558 2150
rect 10614 2148 10638 2150
rect 10694 2148 10718 2150
rect 10774 2148 10780 2150
rect 10472 2139 10780 2148
rect 10980 2106 11008 2790
rect 11072 2514 11100 3334
rect 11164 3058 11192 3538
rect 11152 3052 11204 3058
rect 11152 2994 11204 3000
rect 11060 2508 11112 2514
rect 11060 2450 11112 2456
rect 11256 2446 11284 4014
rect 11348 2990 11376 4644
rect 11520 4684 11572 4690
rect 11520 4626 11572 4632
rect 11532 4214 11560 4626
rect 11900 4622 11928 4694
rect 13464 4690 13492 5102
rect 13740 4826 13768 5102
rect 14660 5098 14688 6666
rect 14648 5092 14700 5098
rect 14648 5034 14700 5040
rect 13830 4924 14138 4933
rect 13830 4922 13836 4924
rect 13892 4922 13916 4924
rect 13972 4922 13996 4924
rect 14052 4922 14076 4924
rect 14132 4922 14138 4924
rect 13892 4870 13894 4922
rect 14074 4870 14076 4922
rect 13830 4868 13836 4870
rect 13892 4868 13916 4870
rect 13972 4868 13996 4870
rect 14052 4868 14076 4870
rect 14132 4868 14138 4870
rect 13830 4859 14138 4868
rect 14844 4826 14872 8327
rect 13728 4820 13780 4826
rect 13728 4762 13780 4768
rect 14832 4820 14884 4826
rect 14832 4762 14884 4768
rect 13176 4684 13228 4690
rect 13176 4626 13228 4632
rect 13452 4684 13504 4690
rect 13452 4626 13504 4632
rect 14464 4684 14516 4690
rect 14464 4626 14516 4632
rect 11796 4616 11848 4622
rect 11796 4558 11848 4564
rect 11888 4616 11940 4622
rect 11888 4558 11940 4564
rect 11520 4208 11572 4214
rect 11520 4150 11572 4156
rect 11808 4078 11836 4558
rect 11796 4072 11848 4078
rect 11796 4014 11848 4020
rect 11900 3618 11928 4558
rect 12348 4548 12400 4554
rect 12348 4490 12400 4496
rect 12072 4208 12124 4214
rect 12072 4150 12124 4156
rect 11900 3602 12020 3618
rect 11900 3596 12032 3602
rect 11900 3590 11980 3596
rect 11980 3538 12032 3544
rect 12084 3126 12112 4150
rect 12360 4078 12388 4490
rect 13188 4282 13216 4626
rect 14476 4282 14504 4626
rect 13176 4276 13228 4282
rect 13176 4218 13228 4224
rect 14464 4276 14516 4282
rect 14464 4218 14516 4224
rect 12348 4072 12400 4078
rect 12348 4014 12400 4020
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 14188 4072 14240 4078
rect 14188 4014 14240 4020
rect 14740 4072 14792 4078
rect 14740 4014 14792 4020
rect 12820 3942 12848 4014
rect 13728 4004 13780 4010
rect 13728 3946 13780 3952
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 12808 3936 12860 3942
rect 12808 3878 12860 3884
rect 12728 3670 12756 3878
rect 12820 3738 12848 3878
rect 12808 3732 12860 3738
rect 12808 3674 12860 3680
rect 12716 3664 12768 3670
rect 12716 3606 12768 3612
rect 13452 3596 13504 3602
rect 13452 3538 13504 3544
rect 12808 3392 12860 3398
rect 12808 3334 12860 3340
rect 12072 3120 12124 3126
rect 12072 3062 12124 3068
rect 12084 2990 12112 3062
rect 12820 2990 12848 3334
rect 13464 3194 13492 3538
rect 13740 3194 13768 3946
rect 13830 3836 14138 3845
rect 13830 3834 13836 3836
rect 13892 3834 13916 3836
rect 13972 3834 13996 3836
rect 14052 3834 14076 3836
rect 14132 3834 14138 3836
rect 13892 3782 13894 3834
rect 14074 3782 14076 3834
rect 13830 3780 13836 3782
rect 13892 3780 13916 3782
rect 13972 3780 13996 3782
rect 14052 3780 14076 3782
rect 14132 3780 14138 3782
rect 13830 3771 14138 3780
rect 14200 3738 14228 4014
rect 14188 3732 14240 3738
rect 14188 3674 14240 3680
rect 14188 3596 14240 3602
rect 14188 3538 14240 3544
rect 13452 3188 13504 3194
rect 13452 3130 13504 3136
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 13542 3088 13598 3097
rect 13542 3023 13598 3032
rect 13556 2990 13584 3023
rect 11336 2984 11388 2990
rect 11334 2952 11336 2961
rect 12072 2984 12124 2990
rect 11388 2952 11390 2961
rect 12072 2926 12124 2932
rect 12808 2984 12860 2990
rect 12808 2926 12860 2932
rect 13544 2984 13596 2990
rect 13544 2926 13596 2932
rect 11334 2887 11390 2896
rect 11796 2916 11848 2922
rect 11796 2858 11848 2864
rect 11612 2848 11664 2854
rect 11612 2790 11664 2796
rect 11624 2514 11652 2790
rect 11808 2514 11836 2858
rect 12716 2848 12768 2854
rect 12716 2790 12768 2796
rect 11612 2508 11664 2514
rect 11612 2450 11664 2456
rect 11796 2508 11848 2514
rect 11796 2450 11848 2456
rect 11244 2440 11296 2446
rect 11244 2382 11296 2388
rect 11244 2304 11296 2310
rect 11244 2246 11296 2252
rect 11336 2304 11388 2310
rect 11336 2246 11388 2252
rect 10968 2100 11020 2106
rect 10968 2042 11020 2048
rect 10232 1964 10284 1970
rect 10232 1906 10284 1912
rect 10048 1896 10100 1902
rect 10048 1838 10100 1844
rect 10876 1896 10928 1902
rect 10876 1838 10928 1844
rect 11060 1896 11112 1902
rect 11060 1838 11112 1844
rect 9956 1420 10008 1426
rect 9956 1362 10008 1368
rect 9680 808 9732 814
rect 9680 750 9732 756
rect 10060 400 10088 1838
rect 10472 1116 10780 1125
rect 10472 1114 10478 1116
rect 10534 1114 10558 1116
rect 10614 1114 10638 1116
rect 10694 1114 10718 1116
rect 10774 1114 10780 1116
rect 10534 1062 10536 1114
rect 10716 1062 10718 1114
rect 10472 1060 10478 1062
rect 10534 1060 10558 1062
rect 10614 1060 10638 1062
rect 10694 1060 10718 1062
rect 10774 1060 10780 1062
rect 10472 1051 10780 1060
rect 10888 882 10916 1838
rect 11072 1494 11100 1838
rect 11152 1556 11204 1562
rect 11152 1498 11204 1504
rect 11060 1488 11112 1494
rect 11060 1430 11112 1436
rect 10876 876 10928 882
rect 10876 818 10928 824
rect 10600 808 10652 814
rect 10600 750 10652 756
rect 10612 400 10640 750
rect 11164 400 11192 1498
rect 11256 814 11284 2246
rect 11348 1426 11376 2246
rect 11808 1834 11836 2450
rect 12728 2378 12756 2790
rect 12900 2644 12952 2650
rect 12900 2586 12952 2592
rect 12716 2372 12768 2378
rect 12716 2314 12768 2320
rect 11888 2304 11940 2310
rect 11888 2246 11940 2252
rect 12256 2304 12308 2310
rect 12256 2246 12308 2252
rect 11900 1902 11928 2246
rect 11888 1896 11940 1902
rect 11888 1838 11940 1844
rect 11796 1828 11848 1834
rect 11796 1770 11848 1776
rect 11336 1420 11388 1426
rect 11336 1362 11388 1368
rect 12072 1420 12124 1426
rect 12072 1362 12124 1368
rect 11244 808 11296 814
rect 11244 750 11296 756
rect 11704 808 11756 814
rect 11704 750 11756 756
rect 12084 762 12112 1362
rect 12268 882 12296 2246
rect 12912 1902 12940 2586
rect 13556 2446 13584 2926
rect 13636 2916 13688 2922
rect 13636 2858 13688 2864
rect 13648 2446 13676 2858
rect 13544 2440 13596 2446
rect 13544 2382 13596 2388
rect 13636 2440 13688 2446
rect 13636 2382 13688 2388
rect 12716 1896 12768 1902
rect 12900 1896 12952 1902
rect 12768 1856 12848 1884
rect 12716 1838 12768 1844
rect 12256 876 12308 882
rect 12256 818 12308 824
rect 11716 400 11744 750
rect 12084 734 12296 762
rect 12268 400 12296 734
rect 12820 400 12848 1856
rect 12900 1838 12952 1844
rect 13544 1896 13596 1902
rect 13544 1838 13596 1844
rect 12992 1760 13044 1766
rect 12992 1702 13044 1708
rect 13176 1760 13228 1766
rect 13176 1702 13228 1708
rect 13004 1426 13032 1702
rect 12992 1420 13044 1426
rect 12992 1362 13044 1368
rect 13188 814 13216 1702
rect 13556 1426 13584 1838
rect 13740 1426 13768 3130
rect 13910 2952 13966 2961
rect 13910 2887 13912 2896
rect 13964 2887 13966 2896
rect 13912 2858 13964 2864
rect 14200 2854 14228 3538
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 14292 3194 14320 3470
rect 14280 3188 14332 3194
rect 14280 3130 14332 3136
rect 14752 3126 14780 4014
rect 14936 3890 14964 9862
rect 15212 9722 15240 9862
rect 15396 9722 15424 10406
rect 15200 9716 15252 9722
rect 15200 9658 15252 9664
rect 15384 9716 15436 9722
rect 15384 9658 15436 9664
rect 15384 9444 15436 9450
rect 15488 9432 15516 10526
rect 15672 10146 15700 10542
rect 15856 10266 15884 10542
rect 16028 10532 16080 10538
rect 16028 10474 16080 10480
rect 16040 10266 16068 10474
rect 15844 10260 15896 10266
rect 15844 10202 15896 10208
rect 16028 10260 16080 10266
rect 16028 10202 16080 10208
rect 15580 10118 15700 10146
rect 15580 10062 15608 10118
rect 15568 10056 15620 10062
rect 15568 9998 15620 10004
rect 15660 10056 15712 10062
rect 15660 9998 15712 10004
rect 15580 9586 15608 9998
rect 15672 9654 15700 9998
rect 15660 9648 15712 9654
rect 15660 9590 15712 9596
rect 15568 9580 15620 9586
rect 15568 9522 15620 9528
rect 15436 9404 15516 9432
rect 15384 9386 15436 9392
rect 15016 9376 15068 9382
rect 15016 9318 15068 9324
rect 15028 9110 15056 9318
rect 15396 9110 15424 9386
rect 15016 9104 15068 9110
rect 15016 9046 15068 9052
rect 15384 9104 15436 9110
rect 15384 9046 15436 9052
rect 15580 9024 15608 9522
rect 15856 9500 15884 10202
rect 16028 10124 16080 10130
rect 16132 10112 16160 10950
rect 16212 10600 16264 10606
rect 16212 10542 16264 10548
rect 16224 10130 16252 10542
rect 16080 10084 16160 10112
rect 16212 10124 16264 10130
rect 16028 10066 16080 10072
rect 16212 10066 16264 10072
rect 16316 9586 16344 14350
rect 16396 13320 16448 13326
rect 16396 13262 16448 13268
rect 16408 12850 16436 13262
rect 16396 12844 16448 12850
rect 16396 12786 16448 12792
rect 16408 11762 16436 12786
rect 16396 11756 16448 11762
rect 16396 11698 16448 11704
rect 16592 11286 16620 15574
rect 16684 15366 16712 16662
rect 16776 16454 16804 17478
rect 16868 17134 16896 17546
rect 16856 17128 16908 17134
rect 16856 17070 16908 17076
rect 16856 16992 16908 16998
rect 16856 16934 16908 16940
rect 16764 16448 16816 16454
rect 16764 16390 16816 16396
rect 16868 15570 16896 16934
rect 16960 16794 16988 17682
rect 16948 16788 17000 16794
rect 16948 16730 17000 16736
rect 17052 15570 17080 19774
rect 17188 19612 17496 19621
rect 17188 19610 17194 19612
rect 17250 19610 17274 19612
rect 17330 19610 17354 19612
rect 17410 19610 17434 19612
rect 17490 19610 17496 19612
rect 17250 19558 17252 19610
rect 17432 19558 17434 19610
rect 17188 19556 17194 19558
rect 17250 19556 17274 19558
rect 17330 19556 17354 19558
rect 17410 19556 17434 19558
rect 17490 19556 17496 19558
rect 17188 19547 17496 19556
rect 17604 19514 17632 19858
rect 17592 19508 17644 19514
rect 17592 19450 17644 19456
rect 17316 19440 17368 19446
rect 17316 19382 17368 19388
rect 17328 19310 17356 19382
rect 17316 19304 17368 19310
rect 17222 19272 17278 19281
rect 17316 19246 17368 19252
rect 17590 19272 17646 19281
rect 17222 19207 17224 19216
rect 17276 19207 17278 19216
rect 17590 19207 17592 19216
rect 17224 19178 17276 19184
rect 17644 19207 17646 19216
rect 17592 19178 17644 19184
rect 17696 18986 17724 20946
rect 17788 20874 17816 20946
rect 17868 20936 17920 20942
rect 17868 20878 17920 20884
rect 17776 20868 17828 20874
rect 17776 20810 17828 20816
rect 17788 20534 17816 20810
rect 17776 20528 17828 20534
rect 17776 20470 17828 20476
rect 17788 19446 17816 20470
rect 17880 20398 17908 20878
rect 17960 20460 18012 20466
rect 17960 20402 18012 20408
rect 17868 20392 17920 20398
rect 17868 20334 17920 20340
rect 17776 19440 17828 19446
rect 17776 19382 17828 19388
rect 17604 18958 17724 18986
rect 17604 18714 17632 18958
rect 17684 18828 17736 18834
rect 17684 18770 17736 18776
rect 17512 18686 17632 18714
rect 17512 18630 17540 18686
rect 17500 18624 17552 18630
rect 17500 18566 17552 18572
rect 17188 18524 17496 18533
rect 17188 18522 17194 18524
rect 17250 18522 17274 18524
rect 17330 18522 17354 18524
rect 17410 18522 17434 18524
rect 17490 18522 17496 18524
rect 17250 18470 17252 18522
rect 17432 18470 17434 18522
rect 17188 18468 17194 18470
rect 17250 18468 17274 18470
rect 17330 18468 17354 18470
rect 17410 18468 17434 18470
rect 17490 18468 17496 18470
rect 17188 18459 17496 18468
rect 17604 18086 17632 18686
rect 17696 18426 17724 18770
rect 17684 18420 17736 18426
rect 17684 18362 17736 18368
rect 17682 18320 17738 18329
rect 17682 18255 17738 18264
rect 17696 18222 17724 18255
rect 17788 18222 17816 19382
rect 17880 19378 17908 20334
rect 17972 19990 18000 20402
rect 18052 20256 18104 20262
rect 18052 20198 18104 20204
rect 17960 19984 18012 19990
rect 17960 19926 18012 19932
rect 17868 19372 17920 19378
rect 17868 19314 17920 19320
rect 17880 18290 17908 19314
rect 18064 19310 18092 20198
rect 18052 19304 18104 19310
rect 18052 19246 18104 19252
rect 17868 18284 17920 18290
rect 17868 18226 17920 18232
rect 18156 18222 18184 22063
rect 18234 20496 18290 20505
rect 18234 20431 18290 20440
rect 17684 18216 17736 18222
rect 17684 18158 17736 18164
rect 17776 18216 17828 18222
rect 17776 18158 17828 18164
rect 17960 18216 18012 18222
rect 17960 18158 18012 18164
rect 18144 18216 18196 18222
rect 18144 18158 18196 18164
rect 17592 18080 17644 18086
rect 17592 18022 17644 18028
rect 17776 18080 17828 18086
rect 17776 18022 17828 18028
rect 17592 17536 17644 17542
rect 17592 17478 17644 17484
rect 17188 17436 17496 17445
rect 17188 17434 17194 17436
rect 17250 17434 17274 17436
rect 17330 17434 17354 17436
rect 17410 17434 17434 17436
rect 17490 17434 17496 17436
rect 17250 17382 17252 17434
rect 17432 17382 17434 17434
rect 17188 17380 17194 17382
rect 17250 17380 17274 17382
rect 17330 17380 17354 17382
rect 17410 17380 17434 17382
rect 17490 17380 17496 17382
rect 17188 17371 17496 17380
rect 17604 17134 17632 17478
rect 17592 17128 17644 17134
rect 17592 17070 17644 17076
rect 17224 16992 17276 16998
rect 17224 16934 17276 16940
rect 17236 16658 17264 16934
rect 17684 16788 17736 16794
rect 17684 16730 17736 16736
rect 17224 16652 17276 16658
rect 17224 16594 17276 16600
rect 17592 16652 17644 16658
rect 17592 16594 17644 16600
rect 17188 16348 17496 16357
rect 17188 16346 17194 16348
rect 17250 16346 17274 16348
rect 17330 16346 17354 16348
rect 17410 16346 17434 16348
rect 17490 16346 17496 16348
rect 17250 16294 17252 16346
rect 17432 16294 17434 16346
rect 17188 16292 17194 16294
rect 17250 16292 17274 16294
rect 17330 16292 17354 16294
rect 17410 16292 17434 16294
rect 17490 16292 17496 16294
rect 17188 16283 17496 16292
rect 17604 16250 17632 16594
rect 17592 16244 17644 16250
rect 17592 16186 17644 16192
rect 17696 16046 17724 16730
rect 17684 16040 17736 16046
rect 17684 15982 17736 15988
rect 17696 15706 17724 15982
rect 17788 15978 17816 18022
rect 17972 17882 18000 18158
rect 17960 17876 18012 17882
rect 17960 17818 18012 17824
rect 17868 17808 17920 17814
rect 17868 17750 17920 17756
rect 17880 17066 17908 17750
rect 18248 17746 18276 20431
rect 18340 20330 18368 22066
rect 18420 21344 18472 21350
rect 18420 21286 18472 21292
rect 18328 20324 18380 20330
rect 18328 20266 18380 20272
rect 18236 17740 18288 17746
rect 18236 17682 18288 17688
rect 18328 17672 18380 17678
rect 18328 17614 18380 17620
rect 18052 17332 18104 17338
rect 18052 17274 18104 17280
rect 17960 17264 18012 17270
rect 17960 17206 18012 17212
rect 17868 17060 17920 17066
rect 17868 17002 17920 17008
rect 17880 16046 17908 17002
rect 17972 16726 18000 17206
rect 18064 17134 18092 17274
rect 18340 17134 18368 17614
rect 18052 17128 18104 17134
rect 18052 17070 18104 17076
rect 18328 17128 18380 17134
rect 18328 17070 18380 17076
rect 18236 17060 18288 17066
rect 18236 17002 18288 17008
rect 17960 16720 18012 16726
rect 17960 16662 18012 16668
rect 17868 16040 17920 16046
rect 17868 15982 17920 15988
rect 17776 15972 17828 15978
rect 17776 15914 17828 15920
rect 17684 15700 17736 15706
rect 17684 15642 17736 15648
rect 16856 15564 16908 15570
rect 16856 15506 16908 15512
rect 17040 15564 17092 15570
rect 17040 15506 17092 15512
rect 17592 15428 17644 15434
rect 17592 15370 17644 15376
rect 16672 15360 16724 15366
rect 16672 15302 16724 15308
rect 17040 15360 17092 15366
rect 17040 15302 17092 15308
rect 16856 14884 16908 14890
rect 16856 14826 16908 14832
rect 16868 14618 16896 14826
rect 16856 14612 16908 14618
rect 16856 14554 16908 14560
rect 17052 14482 17080 15302
rect 17188 15260 17496 15269
rect 17188 15258 17194 15260
rect 17250 15258 17274 15260
rect 17330 15258 17354 15260
rect 17410 15258 17434 15260
rect 17490 15258 17496 15260
rect 17250 15206 17252 15258
rect 17432 15206 17434 15258
rect 17188 15204 17194 15206
rect 17250 15204 17274 15206
rect 17330 15204 17354 15206
rect 17410 15204 17434 15206
rect 17490 15204 17496 15206
rect 17188 15195 17496 15204
rect 17500 14816 17552 14822
rect 17500 14758 17552 14764
rect 17512 14550 17540 14758
rect 17500 14544 17552 14550
rect 17500 14486 17552 14492
rect 17040 14476 17092 14482
rect 17040 14418 17092 14424
rect 17188 14172 17496 14181
rect 17188 14170 17194 14172
rect 17250 14170 17274 14172
rect 17330 14170 17354 14172
rect 17410 14170 17434 14172
rect 17490 14170 17496 14172
rect 17250 14118 17252 14170
rect 17432 14118 17434 14170
rect 17188 14116 17194 14118
rect 17250 14116 17274 14118
rect 17330 14116 17354 14118
rect 17410 14116 17434 14118
rect 17490 14116 17496 14118
rect 17188 14107 17496 14116
rect 17604 13870 17632 15370
rect 16764 13864 16816 13870
rect 16764 13806 16816 13812
rect 17592 13864 17644 13870
rect 17592 13806 17644 13812
rect 16776 12986 16804 13806
rect 16948 13728 17000 13734
rect 16948 13670 17000 13676
rect 16960 13462 16988 13670
rect 16948 13456 17000 13462
rect 16948 13398 17000 13404
rect 17684 13252 17736 13258
rect 17684 13194 17736 13200
rect 17592 13184 17644 13190
rect 17592 13126 17644 13132
rect 17188 13084 17496 13093
rect 17188 13082 17194 13084
rect 17250 13082 17274 13084
rect 17330 13082 17354 13084
rect 17410 13082 17434 13084
rect 17490 13082 17496 13084
rect 17250 13030 17252 13082
rect 17432 13030 17434 13082
rect 17188 13028 17194 13030
rect 17250 13028 17274 13030
rect 17330 13028 17354 13030
rect 17410 13028 17434 13030
rect 17490 13028 17496 13030
rect 17188 13019 17496 13028
rect 16764 12980 16816 12986
rect 16764 12922 16816 12928
rect 17040 12980 17092 12986
rect 17040 12922 17092 12928
rect 16948 11620 17000 11626
rect 16948 11562 17000 11568
rect 16960 11354 16988 11562
rect 16948 11348 17000 11354
rect 16948 11290 17000 11296
rect 16580 11280 16632 11286
rect 16580 11222 16632 11228
rect 17052 10742 17080 12922
rect 17604 12782 17632 13126
rect 17696 12782 17724 13194
rect 17592 12776 17644 12782
rect 17592 12718 17644 12724
rect 17684 12776 17736 12782
rect 17684 12718 17736 12724
rect 17188 11996 17496 12005
rect 17188 11994 17194 11996
rect 17250 11994 17274 11996
rect 17330 11994 17354 11996
rect 17410 11994 17434 11996
rect 17490 11994 17496 11996
rect 17250 11942 17252 11994
rect 17432 11942 17434 11994
rect 17188 11940 17194 11942
rect 17250 11940 17274 11942
rect 17330 11940 17354 11942
rect 17410 11940 17434 11942
rect 17490 11940 17496 11942
rect 17188 11931 17496 11940
rect 17132 11552 17184 11558
rect 17132 11494 17184 11500
rect 17144 11218 17172 11494
rect 17132 11212 17184 11218
rect 17132 11154 17184 11160
rect 17188 10908 17496 10917
rect 17188 10906 17194 10908
rect 17250 10906 17274 10908
rect 17330 10906 17354 10908
rect 17410 10906 17434 10908
rect 17490 10906 17496 10908
rect 17250 10854 17252 10906
rect 17432 10854 17434 10906
rect 17188 10852 17194 10854
rect 17250 10852 17274 10854
rect 17330 10852 17354 10854
rect 17410 10852 17434 10854
rect 17490 10852 17496 10854
rect 17188 10843 17496 10852
rect 17788 10849 17816 15914
rect 17880 15638 17908 15982
rect 17868 15632 17920 15638
rect 17868 15574 17920 15580
rect 17960 15496 18012 15502
rect 17960 15438 18012 15444
rect 17972 14958 18000 15438
rect 17960 14952 18012 14958
rect 17960 14894 18012 14900
rect 17960 14816 18012 14822
rect 17960 14758 18012 14764
rect 17972 14482 18000 14758
rect 17960 14476 18012 14482
rect 17960 14418 18012 14424
rect 18144 14476 18196 14482
rect 18144 14418 18196 14424
rect 18156 14074 18184 14418
rect 18144 14068 18196 14074
rect 18144 14010 18196 14016
rect 18052 13796 18104 13802
rect 18052 13738 18104 13744
rect 18064 13530 18092 13738
rect 18052 13524 18104 13530
rect 18052 13466 18104 13472
rect 17960 12708 18012 12714
rect 17960 12650 18012 12656
rect 17868 12232 17920 12238
rect 17868 12174 17920 12180
rect 17880 11898 17908 12174
rect 17868 11892 17920 11898
rect 17868 11834 17920 11840
rect 17880 11218 17908 11834
rect 17868 11212 17920 11218
rect 17868 11154 17920 11160
rect 17972 11014 18000 12650
rect 18144 12096 18196 12102
rect 18144 12038 18196 12044
rect 18156 11898 18184 12038
rect 18144 11892 18196 11898
rect 18144 11834 18196 11840
rect 17868 11008 17920 11014
rect 17868 10950 17920 10956
rect 17960 11008 18012 11014
rect 18248 10962 18276 17002
rect 18340 16794 18368 17070
rect 18432 17066 18460 21286
rect 18524 19242 18552 26687
rect 18604 26240 18656 26246
rect 18604 26182 18656 26188
rect 18616 25838 18644 26182
rect 18708 25906 18736 27474
rect 18696 25900 18748 25906
rect 18696 25842 18748 25848
rect 18604 25832 18656 25838
rect 18604 25774 18656 25780
rect 18800 23186 18828 28070
rect 18892 28014 18920 29124
rect 18972 29106 19024 29112
rect 19168 29102 19196 30806
rect 23492 30802 23520 31600
rect 22928 30796 22980 30802
rect 22928 30738 22980 30744
rect 23480 30796 23532 30802
rect 23480 30738 23532 30744
rect 20444 30728 20496 30734
rect 20444 30670 20496 30676
rect 19432 30660 19484 30666
rect 19432 30602 19484 30608
rect 19248 30592 19300 30598
rect 19248 30534 19300 30540
rect 19260 30122 19288 30534
rect 19248 30116 19300 30122
rect 19248 30058 19300 30064
rect 19340 30116 19392 30122
rect 19340 30058 19392 30064
rect 19156 29096 19208 29102
rect 19156 29038 19208 29044
rect 18972 28416 19024 28422
rect 18972 28358 19024 28364
rect 18984 28014 19012 28358
rect 19168 28014 19196 29038
rect 19352 28626 19380 30058
rect 19444 29034 19472 30602
rect 20456 30258 20484 30670
rect 22376 30592 22428 30598
rect 22376 30534 22428 30540
rect 22560 30592 22612 30598
rect 22560 30534 22612 30540
rect 21548 30320 21600 30326
rect 21548 30262 21600 30268
rect 20444 30252 20496 30258
rect 20444 30194 20496 30200
rect 20456 29714 20484 30194
rect 21560 30122 21588 30262
rect 21824 30252 21876 30258
rect 21824 30194 21876 30200
rect 21548 30116 21600 30122
rect 21548 30058 21600 30064
rect 21364 30048 21416 30054
rect 21364 29990 21416 29996
rect 21456 30048 21508 30054
rect 21456 29990 21508 29996
rect 20546 29948 20854 29957
rect 20546 29946 20552 29948
rect 20608 29946 20632 29948
rect 20688 29946 20712 29948
rect 20768 29946 20792 29948
rect 20848 29946 20854 29948
rect 20608 29894 20610 29946
rect 20790 29894 20792 29946
rect 20546 29892 20552 29894
rect 20608 29892 20632 29894
rect 20688 29892 20712 29894
rect 20768 29892 20792 29894
rect 20848 29892 20854 29894
rect 20546 29883 20854 29892
rect 21376 29782 21404 29990
rect 21364 29776 21416 29782
rect 21364 29718 21416 29724
rect 20444 29708 20496 29714
rect 20444 29650 20496 29656
rect 20076 29572 20128 29578
rect 20076 29514 20128 29520
rect 20088 29102 20116 29514
rect 20260 29504 20312 29510
rect 20260 29446 20312 29452
rect 20272 29170 20300 29446
rect 20352 29300 20404 29306
rect 20352 29242 20404 29248
rect 20260 29164 20312 29170
rect 20260 29106 20312 29112
rect 20076 29096 20128 29102
rect 20076 29038 20128 29044
rect 19432 29028 19484 29034
rect 19484 28988 19564 29016
rect 19432 28970 19484 28976
rect 19340 28620 19392 28626
rect 19340 28562 19392 28568
rect 18880 28008 18932 28014
rect 18880 27950 18932 27956
rect 18972 28008 19024 28014
rect 18972 27950 19024 27956
rect 19156 28008 19208 28014
rect 19156 27950 19208 27956
rect 18984 25362 19012 27950
rect 19352 27538 19380 28562
rect 19340 27532 19392 27538
rect 19340 27474 19392 27480
rect 19432 27532 19484 27538
rect 19432 27474 19484 27480
rect 19248 27328 19300 27334
rect 19248 27270 19300 27276
rect 19260 26926 19288 27270
rect 19444 27130 19472 27474
rect 19432 27124 19484 27130
rect 19432 27066 19484 27072
rect 19248 26920 19300 26926
rect 19248 26862 19300 26868
rect 19340 26376 19392 26382
rect 19340 26318 19392 26324
rect 19352 25498 19380 26318
rect 19340 25492 19392 25498
rect 19340 25434 19392 25440
rect 18972 25356 19024 25362
rect 18972 25298 19024 25304
rect 18984 24206 19012 25298
rect 19064 24744 19116 24750
rect 19064 24686 19116 24692
rect 19076 24410 19104 24686
rect 19064 24404 19116 24410
rect 19064 24346 19116 24352
rect 18972 24200 19024 24206
rect 18972 24142 19024 24148
rect 18880 24064 18932 24070
rect 18880 24006 18932 24012
rect 18892 23322 18920 24006
rect 18880 23316 18932 23322
rect 18880 23258 18932 23264
rect 18788 23180 18840 23186
rect 18788 23122 18840 23128
rect 19340 23112 19392 23118
rect 19340 23054 19392 23060
rect 18880 22976 18932 22982
rect 18880 22918 18932 22924
rect 18892 22098 18920 22918
rect 19352 22642 19380 23054
rect 19340 22636 19392 22642
rect 19340 22578 19392 22584
rect 19536 22506 19564 28988
rect 19708 28552 19760 28558
rect 19708 28494 19760 28500
rect 19720 28014 19748 28494
rect 20088 28218 20116 29038
rect 20364 29034 20392 29242
rect 21376 29170 21404 29718
rect 21468 29714 21496 29990
rect 21560 29850 21588 30058
rect 21548 29844 21600 29850
rect 21548 29786 21600 29792
rect 21836 29714 21864 30194
rect 22284 30184 22336 30190
rect 22284 30126 22336 30132
rect 22008 30048 22060 30054
rect 22008 29990 22060 29996
rect 21456 29708 21508 29714
rect 21456 29650 21508 29656
rect 21824 29708 21876 29714
rect 21824 29650 21876 29656
rect 22020 29510 22048 29990
rect 21456 29504 21508 29510
rect 21456 29446 21508 29452
rect 22008 29504 22060 29510
rect 22008 29446 22060 29452
rect 22192 29504 22244 29510
rect 22192 29446 22244 29452
rect 21468 29306 21496 29446
rect 21456 29300 21508 29306
rect 21456 29242 21508 29248
rect 21548 29232 21600 29238
rect 21548 29174 21600 29180
rect 20904 29164 20956 29170
rect 20904 29106 20956 29112
rect 21364 29164 21416 29170
rect 21364 29106 21416 29112
rect 20352 29028 20404 29034
rect 20352 28970 20404 28976
rect 20076 28212 20128 28218
rect 20076 28154 20128 28160
rect 20364 28014 20392 28970
rect 20546 28860 20854 28869
rect 20546 28858 20552 28860
rect 20608 28858 20632 28860
rect 20688 28858 20712 28860
rect 20768 28858 20792 28860
rect 20848 28858 20854 28860
rect 20608 28806 20610 28858
rect 20790 28806 20792 28858
rect 20546 28804 20552 28806
rect 20608 28804 20632 28806
rect 20688 28804 20712 28806
rect 20768 28804 20792 28806
rect 20848 28804 20854 28806
rect 20546 28795 20854 28804
rect 20916 28150 20944 29106
rect 21272 29096 21324 29102
rect 21272 29038 21324 29044
rect 21284 28218 21312 29038
rect 21272 28212 21324 28218
rect 21272 28154 21324 28160
rect 20904 28144 20956 28150
rect 20904 28086 20956 28092
rect 19708 28008 19760 28014
rect 19708 27950 19760 27956
rect 20352 28008 20404 28014
rect 20352 27950 20404 27956
rect 20916 27946 20944 28086
rect 20904 27940 20956 27946
rect 20904 27882 20956 27888
rect 21272 27940 21324 27946
rect 21272 27882 21324 27888
rect 20546 27772 20854 27781
rect 20546 27770 20552 27772
rect 20608 27770 20632 27772
rect 20688 27770 20712 27772
rect 20768 27770 20792 27772
rect 20848 27770 20854 27772
rect 20608 27718 20610 27770
rect 20790 27718 20792 27770
rect 20546 27716 20552 27718
rect 20608 27716 20632 27718
rect 20688 27716 20712 27718
rect 20768 27716 20792 27718
rect 20848 27716 20854 27718
rect 20546 27707 20854 27716
rect 21180 27396 21232 27402
rect 21180 27338 21232 27344
rect 20720 27328 20772 27334
rect 20720 27270 20772 27276
rect 20732 26790 20760 27270
rect 21192 26926 21220 27338
rect 21284 26994 21312 27882
rect 21456 27872 21508 27878
rect 21456 27814 21508 27820
rect 21364 27668 21416 27674
rect 21364 27610 21416 27616
rect 21272 26988 21324 26994
rect 21272 26930 21324 26936
rect 20904 26920 20956 26926
rect 20904 26862 20956 26868
rect 21088 26920 21140 26926
rect 21088 26862 21140 26868
rect 21180 26920 21232 26926
rect 21180 26862 21232 26868
rect 20720 26784 20772 26790
rect 20720 26726 20772 26732
rect 20546 26684 20854 26693
rect 20546 26682 20552 26684
rect 20608 26682 20632 26684
rect 20688 26682 20712 26684
rect 20768 26682 20792 26684
rect 20848 26682 20854 26684
rect 20608 26630 20610 26682
rect 20790 26630 20792 26682
rect 20546 26628 20552 26630
rect 20608 26628 20632 26630
rect 20688 26628 20712 26630
rect 20768 26628 20792 26630
rect 20848 26628 20854 26630
rect 20546 26619 20854 26628
rect 20628 26444 20680 26450
rect 20916 26432 20944 26862
rect 21100 26518 21128 26862
rect 21088 26512 21140 26518
rect 21088 26454 21140 26460
rect 20628 26386 20680 26392
rect 20824 26404 20944 26432
rect 20996 26444 21048 26450
rect 20352 26376 20404 26382
rect 20352 26318 20404 26324
rect 19708 26308 19760 26314
rect 19708 26250 19760 26256
rect 19616 23180 19668 23186
rect 19616 23122 19668 23128
rect 19628 22778 19656 23122
rect 19616 22772 19668 22778
rect 19616 22714 19668 22720
rect 19524 22500 19576 22506
rect 19524 22442 19576 22448
rect 19536 22234 19564 22442
rect 19524 22228 19576 22234
rect 19524 22170 19576 22176
rect 18880 22092 18932 22098
rect 18932 22052 19012 22080
rect 18880 22034 18932 22040
rect 18880 21344 18932 21350
rect 18880 21286 18932 21292
rect 18892 21078 18920 21286
rect 18880 21072 18932 21078
rect 18880 21014 18932 21020
rect 18696 21004 18748 21010
rect 18616 20964 18696 20992
rect 18512 19236 18564 19242
rect 18512 19178 18564 19184
rect 18616 18426 18644 20964
rect 18696 20946 18748 20952
rect 18984 20942 19012 22052
rect 18972 20936 19024 20942
rect 18972 20878 19024 20884
rect 18696 20460 18748 20466
rect 18696 20402 18748 20408
rect 18708 20058 18736 20402
rect 18696 20052 18748 20058
rect 18696 19994 18748 20000
rect 18984 19854 19012 20878
rect 19720 20398 19748 26250
rect 20168 26240 20220 26246
rect 20168 26182 20220 26188
rect 20180 25702 20208 26182
rect 20260 25832 20312 25838
rect 20260 25774 20312 25780
rect 20168 25696 20220 25702
rect 20168 25638 20220 25644
rect 20272 25498 20300 25774
rect 20364 25770 20392 26318
rect 20640 25838 20668 26386
rect 20824 26042 20852 26404
rect 20996 26386 21048 26392
rect 20904 26240 20956 26246
rect 20904 26182 20956 26188
rect 20812 26036 20864 26042
rect 20812 25978 20864 25984
rect 20916 25838 20944 26182
rect 21008 26042 21036 26386
rect 20996 26036 21048 26042
rect 20996 25978 21048 25984
rect 21008 25838 21036 25978
rect 20628 25832 20680 25838
rect 20628 25774 20680 25780
rect 20904 25832 20956 25838
rect 20904 25774 20956 25780
rect 20996 25832 21048 25838
rect 20996 25774 21048 25780
rect 20352 25764 20404 25770
rect 20352 25706 20404 25712
rect 20546 25596 20854 25605
rect 20546 25594 20552 25596
rect 20608 25594 20632 25596
rect 20688 25594 20712 25596
rect 20768 25594 20792 25596
rect 20848 25594 20854 25596
rect 20608 25542 20610 25594
rect 20790 25542 20792 25594
rect 20546 25540 20552 25542
rect 20608 25540 20632 25542
rect 20688 25540 20712 25542
rect 20768 25540 20792 25542
rect 20848 25540 20854 25542
rect 20546 25531 20854 25540
rect 21376 25498 21404 27610
rect 21468 27130 21496 27814
rect 21560 27470 21588 29174
rect 21640 28552 21692 28558
rect 21640 28494 21692 28500
rect 21652 28218 21680 28494
rect 21640 28212 21692 28218
rect 21640 28154 21692 28160
rect 22100 28212 22152 28218
rect 22100 28154 22152 28160
rect 22112 27690 22140 28154
rect 22204 28150 22232 29446
rect 22296 29073 22324 30126
rect 22282 29064 22338 29073
rect 22282 28999 22338 29008
rect 22296 28626 22324 28999
rect 22284 28620 22336 28626
rect 22284 28562 22336 28568
rect 22388 28490 22416 30534
rect 22572 30190 22600 30534
rect 22560 30184 22612 30190
rect 22560 30126 22612 30132
rect 22468 29776 22520 29782
rect 22468 29718 22520 29724
rect 22744 29776 22796 29782
rect 22744 29718 22796 29724
rect 22480 29102 22508 29718
rect 22652 29708 22704 29714
rect 22652 29650 22704 29656
rect 22560 29572 22612 29578
rect 22560 29514 22612 29520
rect 22572 29170 22600 29514
rect 22560 29164 22612 29170
rect 22560 29106 22612 29112
rect 22468 29096 22520 29102
rect 22468 29038 22520 29044
rect 22560 28960 22612 28966
rect 22560 28902 22612 28908
rect 22376 28484 22428 28490
rect 22376 28426 22428 28432
rect 22284 28416 22336 28422
rect 22284 28358 22336 28364
rect 22192 28144 22244 28150
rect 22192 28086 22244 28092
rect 22192 27872 22244 27878
rect 22192 27814 22244 27820
rect 22020 27662 22140 27690
rect 21548 27464 21600 27470
rect 21548 27406 21600 27412
rect 21548 27328 21600 27334
rect 21548 27270 21600 27276
rect 21456 27124 21508 27130
rect 21456 27066 21508 27072
rect 21560 26450 21588 27270
rect 21916 26988 21968 26994
rect 21916 26930 21968 26936
rect 21824 26852 21876 26858
rect 21824 26794 21876 26800
rect 21640 26580 21692 26586
rect 21640 26522 21692 26528
rect 21548 26444 21600 26450
rect 21548 26386 21600 26392
rect 21456 26376 21508 26382
rect 21456 26318 21508 26324
rect 21468 25974 21496 26318
rect 21456 25968 21508 25974
rect 21456 25910 21508 25916
rect 20260 25492 20312 25498
rect 20260 25434 20312 25440
rect 21364 25492 21416 25498
rect 21364 25434 21416 25440
rect 21272 25356 21324 25362
rect 21272 25298 21324 25304
rect 20904 24608 20956 24614
rect 20904 24550 20956 24556
rect 20546 24508 20854 24517
rect 20546 24506 20552 24508
rect 20608 24506 20632 24508
rect 20688 24506 20712 24508
rect 20768 24506 20792 24508
rect 20848 24506 20854 24508
rect 20608 24454 20610 24506
rect 20790 24454 20792 24506
rect 20546 24452 20552 24454
rect 20608 24452 20632 24454
rect 20688 24452 20712 24454
rect 20768 24452 20792 24454
rect 20848 24452 20854 24454
rect 20546 24443 20854 24452
rect 20916 24274 20944 24550
rect 20444 24268 20496 24274
rect 20444 24210 20496 24216
rect 20904 24268 20956 24274
rect 20904 24210 20956 24216
rect 20996 24268 21048 24274
rect 20996 24210 21048 24216
rect 19800 24200 19852 24206
rect 19800 24142 19852 24148
rect 20076 24200 20128 24206
rect 20076 24142 20128 24148
rect 19812 23798 19840 24142
rect 19800 23792 19852 23798
rect 19800 23734 19852 23740
rect 20088 22642 20116 24142
rect 20352 23792 20404 23798
rect 20352 23734 20404 23740
rect 20168 23520 20220 23526
rect 20168 23462 20220 23468
rect 20076 22636 20128 22642
rect 20076 22578 20128 22584
rect 20180 22506 20208 23462
rect 20364 22982 20392 23734
rect 20456 23662 20484 24210
rect 20812 24200 20864 24206
rect 20812 24142 20864 24148
rect 20824 23866 20852 24142
rect 20812 23860 20864 23866
rect 20812 23802 20864 23808
rect 20916 23730 20944 24210
rect 20904 23724 20956 23730
rect 20904 23666 20956 23672
rect 21008 23662 21036 24210
rect 21284 23798 21312 25298
rect 21364 24676 21416 24682
rect 21364 24618 21416 24624
rect 21376 23798 21404 24618
rect 21272 23792 21324 23798
rect 21272 23734 21324 23740
rect 21364 23792 21416 23798
rect 21364 23734 21416 23740
rect 21652 23746 21680 26522
rect 21836 26450 21864 26794
rect 21928 26790 21956 26930
rect 21916 26784 21968 26790
rect 21916 26726 21968 26732
rect 21824 26444 21876 26450
rect 21824 26386 21876 26392
rect 22020 26234 22048 27662
rect 22100 27600 22152 27606
rect 22100 27542 22152 27548
rect 22112 27130 22140 27542
rect 22204 27538 22232 27814
rect 22192 27532 22244 27538
rect 22192 27474 22244 27480
rect 22100 27124 22152 27130
rect 22100 27066 22152 27072
rect 22100 26920 22152 26926
rect 22100 26862 22152 26868
rect 22112 26790 22140 26862
rect 22100 26784 22152 26790
rect 22100 26726 22152 26732
rect 22204 26314 22232 27474
rect 22296 27334 22324 28358
rect 22284 27328 22336 27334
rect 22284 27270 22336 27276
rect 22468 27056 22520 27062
rect 22468 26998 22520 27004
rect 22284 26376 22336 26382
rect 22284 26318 22336 26324
rect 22192 26308 22244 26314
rect 22192 26250 22244 26256
rect 22020 26206 22140 26234
rect 22008 26036 22060 26042
rect 22008 25978 22060 25984
rect 22020 25430 22048 25978
rect 22112 25498 22140 26206
rect 22100 25492 22152 25498
rect 22100 25434 22152 25440
rect 22008 25424 22060 25430
rect 22008 25366 22060 25372
rect 22296 25362 22324 26318
rect 22480 25362 22508 26998
rect 22572 26586 22600 28902
rect 22664 28218 22692 29650
rect 22756 29238 22784 29718
rect 22940 29510 22968 30738
rect 23572 30728 23624 30734
rect 23572 30670 23624 30676
rect 23204 30048 23256 30054
rect 23204 29990 23256 29996
rect 22928 29504 22980 29510
rect 22928 29446 22980 29452
rect 23112 29504 23164 29510
rect 23112 29446 23164 29452
rect 23124 29306 23152 29446
rect 23112 29300 23164 29306
rect 23112 29242 23164 29248
rect 22744 29232 22796 29238
rect 22744 29174 22796 29180
rect 23216 29102 23244 29990
rect 23480 29708 23532 29714
rect 23480 29650 23532 29656
rect 23388 29572 23440 29578
rect 23388 29514 23440 29520
rect 23296 29232 23348 29238
rect 23294 29200 23296 29209
rect 23348 29200 23350 29209
rect 23294 29135 23350 29144
rect 22928 29096 22980 29102
rect 23204 29096 23256 29102
rect 22980 29056 23204 29084
rect 22928 29038 22980 29044
rect 23204 29038 23256 29044
rect 23400 28966 23428 29514
rect 22928 28960 22980 28966
rect 22928 28902 22980 28908
rect 23388 28960 23440 28966
rect 23388 28902 23440 28908
rect 22940 28626 22968 28902
rect 23400 28626 23428 28902
rect 22928 28620 22980 28626
rect 22928 28562 22980 28568
rect 23388 28620 23440 28626
rect 23388 28562 23440 28568
rect 22652 28212 22704 28218
rect 22652 28154 22704 28160
rect 22940 28082 22968 28562
rect 23492 28234 23520 29650
rect 23584 29510 23612 30670
rect 23904 30492 24212 30501
rect 23904 30490 23910 30492
rect 23966 30490 23990 30492
rect 24046 30490 24070 30492
rect 24126 30490 24150 30492
rect 24206 30490 24212 30492
rect 23966 30438 23968 30490
rect 24148 30438 24150 30490
rect 23904 30436 23910 30438
rect 23966 30436 23990 30438
rect 24046 30436 24070 30438
rect 24126 30436 24150 30438
rect 24206 30436 24212 30438
rect 23904 30427 24212 30436
rect 23664 30320 23716 30326
rect 23664 30262 23716 30268
rect 23676 29850 23704 30262
rect 24400 30252 24452 30258
rect 24400 30194 24452 30200
rect 24124 30184 24176 30190
rect 24124 30126 24176 30132
rect 24136 29850 24164 30126
rect 23664 29844 23716 29850
rect 23664 29786 23716 29792
rect 24124 29844 24176 29850
rect 24124 29786 24176 29792
rect 23572 29504 23624 29510
rect 23572 29446 23624 29452
rect 23572 29300 23624 29306
rect 23572 29242 23624 29248
rect 23584 29209 23612 29242
rect 23570 29200 23626 29209
rect 23570 29135 23626 29144
rect 23676 28626 23704 29786
rect 24308 29640 24360 29646
rect 24308 29582 24360 29588
rect 23756 29504 23808 29510
rect 23756 29446 23808 29452
rect 23768 28762 23796 29446
rect 23904 29404 24212 29413
rect 23904 29402 23910 29404
rect 23966 29402 23990 29404
rect 24046 29402 24070 29404
rect 24126 29402 24150 29404
rect 24206 29402 24212 29404
rect 23966 29350 23968 29402
rect 24148 29350 24150 29402
rect 23904 29348 23910 29350
rect 23966 29348 23990 29350
rect 24046 29348 24070 29350
rect 24126 29348 24150 29350
rect 24206 29348 24212 29350
rect 23904 29339 24212 29348
rect 24320 29186 24348 29582
rect 24032 29164 24084 29170
rect 24032 29106 24084 29112
rect 24136 29158 24348 29186
rect 24044 29073 24072 29106
rect 24136 29102 24164 29158
rect 24124 29096 24176 29102
rect 24030 29064 24086 29073
rect 24124 29038 24176 29044
rect 24412 29034 24440 30194
rect 24492 29640 24544 29646
rect 24492 29582 24544 29588
rect 24030 28999 24086 29008
rect 24308 29028 24360 29034
rect 24308 28970 24360 28976
rect 24400 29028 24452 29034
rect 24400 28970 24452 28976
rect 24320 28762 24348 28970
rect 23756 28756 23808 28762
rect 23756 28698 23808 28704
rect 24308 28756 24360 28762
rect 24308 28698 24360 28704
rect 23664 28620 23716 28626
rect 23664 28562 23716 28568
rect 24308 28620 24360 28626
rect 24308 28562 24360 28568
rect 23904 28316 24212 28325
rect 23904 28314 23910 28316
rect 23966 28314 23990 28316
rect 24046 28314 24070 28316
rect 24126 28314 24150 28316
rect 24206 28314 24212 28316
rect 23966 28262 23968 28314
rect 24148 28262 24150 28314
rect 23904 28260 23910 28262
rect 23966 28260 23990 28262
rect 24046 28260 24070 28262
rect 24126 28260 24150 28262
rect 24206 28260 24212 28262
rect 23904 28251 24212 28260
rect 23492 28206 23796 28234
rect 24320 28218 24348 28562
rect 22928 28076 22980 28082
rect 22928 28018 22980 28024
rect 22744 28008 22796 28014
rect 22744 27950 22796 27956
rect 23020 28008 23072 28014
rect 23492 27962 23520 28206
rect 23572 28144 23624 28150
rect 23572 28086 23624 28092
rect 23584 28014 23612 28086
rect 23020 27950 23072 27956
rect 22652 27940 22704 27946
rect 22652 27882 22704 27888
rect 22664 27538 22692 27882
rect 22756 27538 22784 27950
rect 23032 27538 23060 27950
rect 23400 27946 23520 27962
rect 23572 28008 23624 28014
rect 23572 27950 23624 27956
rect 23388 27940 23520 27946
rect 23440 27934 23520 27940
rect 23388 27882 23440 27888
rect 23492 27538 23520 27934
rect 23584 27674 23612 27950
rect 23768 27946 23796 28206
rect 24216 28212 24268 28218
rect 24216 28154 24268 28160
rect 24308 28212 24360 28218
rect 24308 28154 24360 28160
rect 24228 28098 24256 28154
rect 24412 28098 24440 28970
rect 24136 28070 24440 28098
rect 23756 27940 23808 27946
rect 23756 27882 23808 27888
rect 23664 27872 23716 27878
rect 23664 27814 23716 27820
rect 23848 27872 23900 27878
rect 23848 27814 23900 27820
rect 23572 27668 23624 27674
rect 23572 27610 23624 27616
rect 23676 27606 23704 27814
rect 23664 27600 23716 27606
rect 23664 27542 23716 27548
rect 22652 27532 22704 27538
rect 22652 27474 22704 27480
rect 22744 27532 22796 27538
rect 22744 27474 22796 27480
rect 22836 27532 22888 27538
rect 22836 27474 22888 27480
rect 23020 27532 23072 27538
rect 23020 27474 23072 27480
rect 23480 27532 23532 27538
rect 23480 27474 23532 27480
rect 22664 26994 22692 27474
rect 22756 27130 22784 27474
rect 22744 27124 22796 27130
rect 22744 27066 22796 27072
rect 22652 26988 22704 26994
rect 22652 26930 22704 26936
rect 22848 26926 22876 27474
rect 22836 26920 22888 26926
rect 22836 26862 22888 26868
rect 23032 26790 23060 27474
rect 23860 27418 23888 27814
rect 24136 27606 24164 28070
rect 24216 27940 24268 27946
rect 24216 27882 24268 27888
rect 24228 27674 24256 27882
rect 24216 27668 24268 27674
rect 24216 27610 24268 27616
rect 24124 27600 24176 27606
rect 24124 27542 24176 27548
rect 23768 27402 23888 27418
rect 23768 27396 23900 27402
rect 23768 27390 23848 27396
rect 23768 26926 23796 27390
rect 23848 27338 23900 27344
rect 23904 27228 24212 27237
rect 23904 27226 23910 27228
rect 23966 27226 23990 27228
rect 24046 27226 24070 27228
rect 24126 27226 24150 27228
rect 24206 27226 24212 27228
rect 23966 27174 23968 27226
rect 24148 27174 24150 27226
rect 23904 27172 23910 27174
rect 23966 27172 23990 27174
rect 24046 27172 24070 27174
rect 24126 27172 24150 27174
rect 24206 27172 24212 27174
rect 23904 27163 24212 27172
rect 23756 26920 23808 26926
rect 23756 26862 23808 26868
rect 23020 26784 23072 26790
rect 23020 26726 23072 26732
rect 23768 26586 23796 26862
rect 24032 26852 24084 26858
rect 24032 26794 24084 26800
rect 22560 26580 22612 26586
rect 22560 26522 22612 26528
rect 23756 26580 23808 26586
rect 23756 26522 23808 26528
rect 23756 26444 23808 26450
rect 23756 26386 23808 26392
rect 23388 26240 23440 26246
rect 23388 26182 23440 26188
rect 23400 25838 23428 26182
rect 23768 26042 23796 26386
rect 24044 26246 24072 26794
rect 24308 26308 24360 26314
rect 24308 26250 24360 26256
rect 24032 26240 24084 26246
rect 24032 26182 24084 26188
rect 23904 26140 24212 26149
rect 23904 26138 23910 26140
rect 23966 26138 23990 26140
rect 24046 26138 24070 26140
rect 24126 26138 24150 26140
rect 24206 26138 24212 26140
rect 23966 26086 23968 26138
rect 24148 26086 24150 26138
rect 23904 26084 23910 26086
rect 23966 26084 23990 26086
rect 24046 26084 24070 26086
rect 24126 26084 24150 26086
rect 24206 26084 24212 26086
rect 23904 26075 24212 26084
rect 23756 26036 23808 26042
rect 23756 25978 23808 25984
rect 24032 26036 24084 26042
rect 24032 25978 24084 25984
rect 23388 25832 23440 25838
rect 23388 25774 23440 25780
rect 23388 25696 23440 25702
rect 23388 25638 23440 25644
rect 23400 25498 23428 25638
rect 22744 25492 22796 25498
rect 22744 25434 22796 25440
rect 23388 25492 23440 25498
rect 23388 25434 23440 25440
rect 22284 25356 22336 25362
rect 22284 25298 22336 25304
rect 22468 25356 22520 25362
rect 22468 25298 22520 25304
rect 21732 25288 21784 25294
rect 21732 25230 21784 25236
rect 22376 25288 22428 25294
rect 22376 25230 22428 25236
rect 21744 24682 21772 25230
rect 22388 24954 22416 25230
rect 22376 24948 22428 24954
rect 22376 24890 22428 24896
rect 22192 24880 22244 24886
rect 22192 24822 22244 24828
rect 21732 24676 21784 24682
rect 21732 24618 21784 24624
rect 22204 24410 22232 24822
rect 22192 24404 22244 24410
rect 22192 24346 22244 24352
rect 21824 24336 21876 24342
rect 21824 24278 21876 24284
rect 21652 23718 21772 23746
rect 20444 23656 20496 23662
rect 20444 23598 20496 23604
rect 20996 23656 21048 23662
rect 20996 23598 21048 23604
rect 21088 23656 21140 23662
rect 21088 23598 21140 23604
rect 20904 23588 20956 23594
rect 20904 23530 20956 23536
rect 20546 23420 20854 23429
rect 20546 23418 20552 23420
rect 20608 23418 20632 23420
rect 20688 23418 20712 23420
rect 20768 23418 20792 23420
rect 20848 23418 20854 23420
rect 20608 23366 20610 23418
rect 20790 23366 20792 23418
rect 20546 23364 20552 23366
rect 20608 23364 20632 23366
rect 20688 23364 20712 23366
rect 20768 23364 20792 23366
rect 20848 23364 20854 23366
rect 20546 23355 20854 23364
rect 20916 23050 20944 23530
rect 21008 23322 21036 23598
rect 21100 23526 21128 23598
rect 21640 23588 21692 23594
rect 21640 23530 21692 23536
rect 21088 23520 21140 23526
rect 21088 23462 21140 23468
rect 20996 23316 21048 23322
rect 20996 23258 21048 23264
rect 21652 23118 21680 23530
rect 21640 23112 21692 23118
rect 21640 23054 21692 23060
rect 20904 23044 20956 23050
rect 20904 22986 20956 22992
rect 20352 22976 20404 22982
rect 20352 22918 20404 22924
rect 20168 22500 20220 22506
rect 20168 22442 20220 22448
rect 20546 22332 20854 22341
rect 20546 22330 20552 22332
rect 20608 22330 20632 22332
rect 20688 22330 20712 22332
rect 20768 22330 20792 22332
rect 20848 22330 20854 22332
rect 20608 22278 20610 22330
rect 20790 22278 20792 22330
rect 20546 22276 20552 22278
rect 20608 22276 20632 22278
rect 20688 22276 20712 22278
rect 20768 22276 20792 22278
rect 20848 22276 20854 22278
rect 20546 22267 20854 22276
rect 21744 22166 21772 23718
rect 21836 23662 21864 24278
rect 22192 24268 22244 24274
rect 22192 24210 22244 24216
rect 22100 24200 22152 24206
rect 22100 24142 22152 24148
rect 21824 23656 21876 23662
rect 21824 23598 21876 23604
rect 21916 23520 21968 23526
rect 21916 23462 21968 23468
rect 21928 23322 21956 23462
rect 21916 23316 21968 23322
rect 21916 23258 21968 23264
rect 22112 23186 22140 24142
rect 22204 23526 22232 24210
rect 22652 24064 22704 24070
rect 22652 24006 22704 24012
rect 22664 23594 22692 24006
rect 22652 23588 22704 23594
rect 22652 23530 22704 23536
rect 22192 23520 22244 23526
rect 22192 23462 22244 23468
rect 22204 23254 22232 23462
rect 22192 23248 22244 23254
rect 22192 23190 22244 23196
rect 22100 23180 22152 23186
rect 22100 23122 22152 23128
rect 22284 23180 22336 23186
rect 22284 23122 22336 23128
rect 22296 22982 22324 23122
rect 22284 22976 22336 22982
rect 22284 22918 22336 22924
rect 22376 22568 22428 22574
rect 22376 22510 22428 22516
rect 22560 22568 22612 22574
rect 22560 22510 22612 22516
rect 21732 22160 21784 22166
rect 21732 22102 21784 22108
rect 20168 22092 20220 22098
rect 20168 22034 20220 22040
rect 22284 22092 22336 22098
rect 22284 22034 22336 22040
rect 20180 21690 20208 22034
rect 21456 22024 21508 22030
rect 21456 21966 21508 21972
rect 20812 21888 20864 21894
rect 20812 21830 20864 21836
rect 20168 21684 20220 21690
rect 20168 21626 20220 21632
rect 20352 21548 20404 21554
rect 20352 21490 20404 21496
rect 20168 21480 20220 21486
rect 20168 21422 20220 21428
rect 19800 21344 19852 21350
rect 19800 21286 19852 21292
rect 19812 20806 19840 21286
rect 20180 21146 20208 21422
rect 20168 21140 20220 21146
rect 20168 21082 20220 21088
rect 20364 20874 20392 21490
rect 20824 21486 20852 21830
rect 20444 21480 20496 21486
rect 20444 21422 20496 21428
rect 20812 21480 20864 21486
rect 20812 21422 20864 21428
rect 21088 21480 21140 21486
rect 21088 21422 21140 21428
rect 21272 21480 21324 21486
rect 21272 21422 21324 21428
rect 20456 21010 20484 21422
rect 20996 21412 21048 21418
rect 20996 21354 21048 21360
rect 20546 21244 20854 21253
rect 20546 21242 20552 21244
rect 20608 21242 20632 21244
rect 20688 21242 20712 21244
rect 20768 21242 20792 21244
rect 20848 21242 20854 21244
rect 20608 21190 20610 21242
rect 20790 21190 20792 21242
rect 20546 21188 20552 21190
rect 20608 21188 20632 21190
rect 20688 21188 20712 21190
rect 20768 21188 20792 21190
rect 20848 21188 20854 21190
rect 20546 21179 20854 21188
rect 21008 21146 21036 21354
rect 21100 21146 21128 21422
rect 20996 21140 21048 21146
rect 20996 21082 21048 21088
rect 21088 21140 21140 21146
rect 21284 21128 21312 21422
rect 21364 21140 21416 21146
rect 21284 21100 21364 21128
rect 21088 21082 21140 21088
rect 21364 21082 21416 21088
rect 20444 21004 20496 21010
rect 20444 20946 20496 20952
rect 20352 20868 20404 20874
rect 20352 20810 20404 20816
rect 19800 20800 19852 20806
rect 19800 20742 19852 20748
rect 19708 20392 19760 20398
rect 19708 20334 19760 20340
rect 19812 20330 19840 20742
rect 19892 20596 19944 20602
rect 19944 20556 20116 20584
rect 19892 20538 19944 20544
rect 19248 20324 19300 20330
rect 19248 20266 19300 20272
rect 19800 20324 19852 20330
rect 19800 20266 19852 20272
rect 18972 19848 19024 19854
rect 18972 19790 19024 19796
rect 18984 19310 19012 19790
rect 19260 19360 19288 20266
rect 19432 20256 19484 20262
rect 19432 20198 19484 20204
rect 19260 19332 19380 19360
rect 18972 19304 19024 19310
rect 18972 19246 19024 19252
rect 18880 18624 18932 18630
rect 18984 18578 19012 19246
rect 19064 19236 19116 19242
rect 19064 19178 19116 19184
rect 19076 18834 19104 19178
rect 19064 18828 19116 18834
rect 19064 18770 19116 18776
rect 18932 18572 19012 18578
rect 18880 18566 19012 18572
rect 18892 18550 19012 18566
rect 18604 18420 18656 18426
rect 18604 18362 18656 18368
rect 18420 17060 18472 17066
rect 18420 17002 18472 17008
rect 18328 16788 18380 16794
rect 18328 16730 18380 16736
rect 18616 15552 18644 18362
rect 18984 18222 19012 18550
rect 18972 18216 19024 18222
rect 18972 18158 19024 18164
rect 18984 17134 19012 18158
rect 18972 17128 19024 17134
rect 18972 17070 19024 17076
rect 19076 16980 19104 18770
rect 19156 18624 19208 18630
rect 19156 18566 19208 18572
rect 19168 17746 19196 18566
rect 19352 17898 19380 19332
rect 19444 18154 19472 20198
rect 19812 20058 19840 20266
rect 19800 20052 19852 20058
rect 19800 19994 19852 20000
rect 19432 18148 19484 18154
rect 19432 18090 19484 18096
rect 19352 17870 19472 17898
rect 19156 17740 19208 17746
rect 19156 17682 19208 17688
rect 19340 17604 19392 17610
rect 19444 17592 19472 17870
rect 19904 17746 19932 20538
rect 20088 20466 20116 20556
rect 20076 20460 20128 20466
rect 20076 20402 20128 20408
rect 20168 20392 20220 20398
rect 20168 20334 20220 20340
rect 20180 19514 20208 20334
rect 20456 20330 20484 20946
rect 21468 20874 21496 21966
rect 22100 21956 22152 21962
rect 22100 21898 22152 21904
rect 22192 21956 22244 21962
rect 22192 21898 22244 21904
rect 21916 21616 21968 21622
rect 21916 21558 21968 21564
rect 21928 21418 21956 21558
rect 22008 21480 22060 21486
rect 22008 21422 22060 21428
rect 22112 21434 22140 21898
rect 22204 21622 22232 21898
rect 22192 21616 22244 21622
rect 22192 21558 22244 21564
rect 21916 21412 21968 21418
rect 21916 21354 21968 21360
rect 21456 20868 21508 20874
rect 21456 20810 21508 20816
rect 21732 20460 21784 20466
rect 21732 20402 21784 20408
rect 21088 20392 21140 20398
rect 21456 20392 21508 20398
rect 21140 20340 21312 20346
rect 21088 20334 21312 20340
rect 21456 20334 21508 20340
rect 21640 20392 21692 20398
rect 21640 20334 21692 20340
rect 21100 20330 21312 20334
rect 20444 20324 20496 20330
rect 21100 20324 21324 20330
rect 21100 20318 21272 20324
rect 20444 20266 20496 20272
rect 21272 20266 21324 20272
rect 20996 20256 21048 20262
rect 20996 20198 21048 20204
rect 21088 20256 21140 20262
rect 21088 20198 21140 20204
rect 20546 20156 20854 20165
rect 20546 20154 20552 20156
rect 20608 20154 20632 20156
rect 20688 20154 20712 20156
rect 20768 20154 20792 20156
rect 20848 20154 20854 20156
rect 20608 20102 20610 20154
rect 20790 20102 20792 20154
rect 20546 20100 20552 20102
rect 20608 20100 20632 20102
rect 20688 20100 20712 20102
rect 20768 20100 20792 20102
rect 20848 20100 20854 20102
rect 20546 20091 20854 20100
rect 21008 19990 21036 20198
rect 21100 20058 21128 20198
rect 21088 20052 21140 20058
rect 21088 19994 21140 20000
rect 20996 19984 21048 19990
rect 20996 19926 21048 19932
rect 20168 19508 20220 19514
rect 20168 19450 20220 19456
rect 21180 19304 21232 19310
rect 21180 19246 21232 19252
rect 21088 19236 21140 19242
rect 21088 19178 21140 19184
rect 20444 19168 20496 19174
rect 20444 19110 20496 19116
rect 20456 18970 20484 19110
rect 20546 19068 20854 19077
rect 20546 19066 20552 19068
rect 20608 19066 20632 19068
rect 20688 19066 20712 19068
rect 20768 19066 20792 19068
rect 20848 19066 20854 19068
rect 20608 19014 20610 19066
rect 20790 19014 20792 19066
rect 20546 19012 20552 19014
rect 20608 19012 20632 19014
rect 20688 19012 20712 19014
rect 20768 19012 20792 19014
rect 20848 19012 20854 19014
rect 20546 19003 20854 19012
rect 20444 18964 20496 18970
rect 20444 18906 20496 18912
rect 20904 18760 20956 18766
rect 20904 18702 20956 18708
rect 20916 18630 20944 18702
rect 21100 18630 21128 19178
rect 20904 18624 20956 18630
rect 20904 18566 20956 18572
rect 21088 18624 21140 18630
rect 21088 18566 21140 18572
rect 20916 18222 20944 18566
rect 21192 18426 21220 19246
rect 21272 18964 21324 18970
rect 21272 18906 21324 18912
rect 21364 18964 21416 18970
rect 21364 18906 21416 18912
rect 21180 18420 21232 18426
rect 21180 18362 21232 18368
rect 20904 18216 20956 18222
rect 20904 18158 20956 18164
rect 21180 18216 21232 18222
rect 21180 18158 21232 18164
rect 20546 17980 20854 17989
rect 20546 17978 20552 17980
rect 20608 17978 20632 17980
rect 20688 17978 20712 17980
rect 20768 17978 20792 17980
rect 20848 17978 20854 17980
rect 20608 17926 20610 17978
rect 20790 17926 20792 17978
rect 20546 17924 20552 17926
rect 20608 17924 20632 17926
rect 20688 17924 20712 17926
rect 20768 17924 20792 17926
rect 20848 17924 20854 17926
rect 20546 17915 20854 17924
rect 21192 17814 21220 18158
rect 21180 17808 21232 17814
rect 21180 17750 21232 17756
rect 19708 17740 19760 17746
rect 19708 17682 19760 17688
rect 19892 17740 19944 17746
rect 19892 17682 19944 17688
rect 20352 17740 20404 17746
rect 20352 17682 20404 17688
rect 20996 17740 21048 17746
rect 20996 17682 21048 17688
rect 19392 17564 19472 17592
rect 19340 17546 19392 17552
rect 19248 17060 19300 17066
rect 19248 17002 19300 17008
rect 18984 16952 19104 16980
rect 18788 16448 18840 16454
rect 18788 16390 18840 16396
rect 18800 16046 18828 16390
rect 18788 16040 18840 16046
rect 18788 15982 18840 15988
rect 18696 15564 18748 15570
rect 18616 15524 18696 15552
rect 18616 14006 18644 15524
rect 18696 15506 18748 15512
rect 18880 15360 18932 15366
rect 18880 15302 18932 15308
rect 18696 14272 18748 14278
rect 18696 14214 18748 14220
rect 18604 14000 18656 14006
rect 18604 13942 18656 13948
rect 18708 13870 18736 14214
rect 18512 13864 18564 13870
rect 18696 13864 18748 13870
rect 18512 13806 18564 13812
rect 18616 13824 18696 13852
rect 18524 12306 18552 13806
rect 18616 12782 18644 13824
rect 18696 13806 18748 13812
rect 18892 13734 18920 15302
rect 18984 13870 19012 16952
rect 19260 16046 19288 17002
rect 19340 16448 19392 16454
rect 19340 16390 19392 16396
rect 19248 16040 19300 16046
rect 19248 15982 19300 15988
rect 19260 15570 19288 15982
rect 19352 15570 19380 16390
rect 19444 15892 19472 17564
rect 19524 17536 19576 17542
rect 19524 17478 19576 17484
rect 19536 16046 19564 17478
rect 19524 16040 19576 16046
rect 19524 15982 19576 15988
rect 19444 15864 19564 15892
rect 19248 15564 19300 15570
rect 19248 15506 19300 15512
rect 19340 15564 19392 15570
rect 19340 15506 19392 15512
rect 19536 14006 19564 15864
rect 19524 14000 19576 14006
rect 19524 13942 19576 13948
rect 18972 13864 19024 13870
rect 18972 13806 19024 13812
rect 19064 13796 19116 13802
rect 19064 13738 19116 13744
rect 18880 13728 18932 13734
rect 18880 13670 18932 13676
rect 18892 13530 18920 13670
rect 18880 13524 18932 13530
rect 18880 13466 18932 13472
rect 18604 12776 18656 12782
rect 18604 12718 18656 12724
rect 18512 12300 18564 12306
rect 18432 12260 18512 12288
rect 18328 11620 18380 11626
rect 18328 11562 18380 11568
rect 17960 10950 18012 10956
rect 17774 10840 17830 10849
rect 17774 10775 17830 10784
rect 17040 10736 17092 10742
rect 17040 10678 17092 10684
rect 17776 10668 17828 10674
rect 17776 10610 17828 10616
rect 17040 10600 17092 10606
rect 17040 10542 17092 10548
rect 17222 10568 17278 10577
rect 17052 10266 17080 10542
rect 17222 10503 17278 10512
rect 17236 10470 17264 10503
rect 17224 10464 17276 10470
rect 17224 10406 17276 10412
rect 17040 10260 17092 10266
rect 17040 10202 17092 10208
rect 17788 10062 17816 10610
rect 17880 10606 17908 10950
rect 17972 10742 18000 10950
rect 18156 10934 18276 10962
rect 17960 10736 18012 10742
rect 17960 10678 18012 10684
rect 17868 10600 17920 10606
rect 17868 10542 17920 10548
rect 17960 10464 18012 10470
rect 17960 10406 18012 10412
rect 17972 10198 18000 10406
rect 17960 10192 18012 10198
rect 17960 10134 18012 10140
rect 18156 10130 18184 10934
rect 18234 10840 18290 10849
rect 18234 10775 18290 10784
rect 18248 10606 18276 10775
rect 18236 10600 18288 10606
rect 18236 10542 18288 10548
rect 18340 10266 18368 11562
rect 18432 11150 18460 12260
rect 18512 12242 18564 12248
rect 18892 11558 18920 13466
rect 19076 13462 19104 13738
rect 19064 13456 19116 13462
rect 19064 13398 19116 13404
rect 18972 12300 19024 12306
rect 18972 12242 19024 12248
rect 18984 11898 19012 12242
rect 18972 11892 19024 11898
rect 18972 11834 19024 11840
rect 19076 11694 19104 13398
rect 19340 13252 19392 13258
rect 19340 13194 19392 13200
rect 19352 12782 19380 13194
rect 19340 12776 19392 12782
rect 19340 12718 19392 12724
rect 19248 12708 19300 12714
rect 19248 12650 19300 12656
rect 19260 12442 19288 12650
rect 19248 12436 19300 12442
rect 19248 12378 19300 12384
rect 19720 12374 19748 17682
rect 20364 16794 20392 17682
rect 21008 17134 21036 17682
rect 20996 17128 21048 17134
rect 20996 17070 21048 17076
rect 21008 16998 21036 17070
rect 20996 16992 21048 16998
rect 20996 16934 21048 16940
rect 20546 16892 20854 16901
rect 20546 16890 20552 16892
rect 20608 16890 20632 16892
rect 20688 16890 20712 16892
rect 20768 16890 20792 16892
rect 20848 16890 20854 16892
rect 20608 16838 20610 16890
rect 20790 16838 20792 16890
rect 20546 16836 20552 16838
rect 20608 16836 20632 16838
rect 20688 16836 20712 16838
rect 20768 16836 20792 16838
rect 20848 16836 20854 16838
rect 20546 16827 20854 16836
rect 20352 16788 20404 16794
rect 20352 16730 20404 16736
rect 21008 16726 21036 16934
rect 20996 16720 21048 16726
rect 20996 16662 21048 16668
rect 19800 16652 19852 16658
rect 19800 16594 19852 16600
rect 19812 16046 19840 16594
rect 20260 16584 20312 16590
rect 20260 16526 20312 16532
rect 21088 16584 21140 16590
rect 21088 16526 21140 16532
rect 19800 16040 19852 16046
rect 19800 15982 19852 15988
rect 20272 15706 20300 16526
rect 21100 16046 21128 16526
rect 21088 16040 21140 16046
rect 21088 15982 21140 15988
rect 21180 16040 21232 16046
rect 21180 15982 21232 15988
rect 21100 15910 21128 15982
rect 21088 15904 21140 15910
rect 21088 15846 21140 15852
rect 20546 15804 20854 15813
rect 20546 15802 20552 15804
rect 20608 15802 20632 15804
rect 20688 15802 20712 15804
rect 20768 15802 20792 15804
rect 20848 15802 20854 15804
rect 20608 15750 20610 15802
rect 20790 15750 20792 15802
rect 20546 15748 20552 15750
rect 20608 15748 20632 15750
rect 20688 15748 20712 15750
rect 20768 15748 20792 15750
rect 20848 15748 20854 15750
rect 20546 15739 20854 15748
rect 20260 15700 20312 15706
rect 20260 15642 20312 15648
rect 21100 15570 21128 15846
rect 21088 15564 21140 15570
rect 21088 15506 21140 15512
rect 21192 15502 21220 15982
rect 21180 15496 21232 15502
rect 21180 15438 21232 15444
rect 21088 14884 21140 14890
rect 21088 14826 21140 14832
rect 20546 14716 20854 14725
rect 20546 14714 20552 14716
rect 20608 14714 20632 14716
rect 20688 14714 20712 14716
rect 20768 14714 20792 14716
rect 20848 14714 20854 14716
rect 20608 14662 20610 14714
rect 20790 14662 20792 14714
rect 20546 14660 20552 14662
rect 20608 14660 20632 14662
rect 20688 14660 20712 14662
rect 20768 14660 20792 14662
rect 20848 14660 20854 14662
rect 20546 14651 20854 14660
rect 21100 14482 21128 14826
rect 21284 14482 21312 18906
rect 21376 18834 21404 18906
rect 21468 18834 21496 20334
rect 21548 20256 21600 20262
rect 21548 20198 21600 20204
rect 21364 18828 21416 18834
rect 21364 18770 21416 18776
rect 21456 18828 21508 18834
rect 21560 18816 21588 20198
rect 21652 20058 21680 20334
rect 21640 20052 21692 20058
rect 21640 19994 21692 20000
rect 21744 19990 21772 20402
rect 21928 20398 21956 21354
rect 22020 21078 22048 21422
rect 22112 21406 22232 21434
rect 22008 21072 22060 21078
rect 22008 21014 22060 21020
rect 22020 20398 22048 21014
rect 22100 20596 22152 20602
rect 22100 20538 22152 20544
rect 21916 20392 21968 20398
rect 21916 20334 21968 20340
rect 22008 20392 22060 20398
rect 22008 20334 22060 20340
rect 21732 19984 21784 19990
rect 21732 19926 21784 19932
rect 22112 19922 22140 20538
rect 22100 19916 22152 19922
rect 22100 19858 22152 19864
rect 22112 19446 22140 19858
rect 22100 19440 22152 19446
rect 22100 19382 22152 19388
rect 21824 19168 21876 19174
rect 21824 19110 21876 19116
rect 21732 18896 21784 18902
rect 21732 18838 21784 18844
rect 21640 18828 21692 18834
rect 21560 18788 21640 18816
rect 21456 18770 21508 18776
rect 21640 18770 21692 18776
rect 21548 18420 21600 18426
rect 21600 18380 21680 18408
rect 21548 18362 21600 18368
rect 21456 18352 21508 18358
rect 21456 18294 21508 18300
rect 21364 18216 21416 18222
rect 21364 18158 21416 18164
rect 21376 17882 21404 18158
rect 21364 17876 21416 17882
rect 21364 17818 21416 17824
rect 21468 17134 21496 18294
rect 21652 17746 21680 18380
rect 21744 18154 21772 18838
rect 21836 18834 21864 19110
rect 21824 18828 21876 18834
rect 21824 18770 21876 18776
rect 21824 18284 21876 18290
rect 21824 18226 21876 18232
rect 21732 18148 21784 18154
rect 21732 18090 21784 18096
rect 21548 17740 21600 17746
rect 21548 17682 21600 17688
rect 21640 17740 21692 17746
rect 21640 17682 21692 17688
rect 21560 17202 21588 17682
rect 21548 17196 21600 17202
rect 21548 17138 21600 17144
rect 21456 17128 21508 17134
rect 21456 17070 21508 17076
rect 21560 16658 21588 17138
rect 21836 16674 21864 18226
rect 22100 18080 22152 18086
rect 22100 18022 22152 18028
rect 21916 17740 21968 17746
rect 21916 17682 21968 17688
rect 21928 16794 21956 17682
rect 22112 17610 22140 18022
rect 22204 17746 22232 21406
rect 22296 21078 22324 22034
rect 22388 21690 22416 22510
rect 22468 22432 22520 22438
rect 22468 22374 22520 22380
rect 22480 21690 22508 22374
rect 22572 22234 22600 22510
rect 22652 22432 22704 22438
rect 22652 22374 22704 22380
rect 22560 22228 22612 22234
rect 22560 22170 22612 22176
rect 22572 21962 22600 22170
rect 22664 22166 22692 22374
rect 22756 22166 22784 25434
rect 23112 25288 23164 25294
rect 23112 25230 23164 25236
rect 23756 25288 23808 25294
rect 23756 25230 23808 25236
rect 23124 24750 23152 25230
rect 23664 25152 23716 25158
rect 23664 25094 23716 25100
rect 23112 24744 23164 24750
rect 23112 24686 23164 24692
rect 22928 22568 22980 22574
rect 22928 22510 22980 22516
rect 22652 22160 22704 22166
rect 22652 22102 22704 22108
rect 22744 22160 22796 22166
rect 22744 22102 22796 22108
rect 22560 21956 22612 21962
rect 22560 21898 22612 21904
rect 22376 21684 22428 21690
rect 22376 21626 22428 21632
rect 22468 21684 22520 21690
rect 22468 21626 22520 21632
rect 22664 21418 22692 22102
rect 22940 22030 22968 22510
rect 23020 22432 23072 22438
rect 23020 22374 23072 22380
rect 23032 22166 23060 22374
rect 23020 22160 23072 22166
rect 23020 22102 23072 22108
rect 22928 22024 22980 22030
rect 22928 21966 22980 21972
rect 22744 21888 22796 21894
rect 22744 21830 22796 21836
rect 22756 21622 22784 21830
rect 22744 21616 22796 21622
rect 22744 21558 22796 21564
rect 22652 21412 22704 21418
rect 22652 21354 22704 21360
rect 22376 21344 22428 21350
rect 22376 21286 22428 21292
rect 22284 21072 22336 21078
rect 22284 21014 22336 21020
rect 22388 20398 22416 21286
rect 22664 20942 22692 21354
rect 22652 20936 22704 20942
rect 22652 20878 22704 20884
rect 22468 20800 22520 20806
rect 22468 20742 22520 20748
rect 22480 20466 22508 20742
rect 22468 20460 22520 20466
rect 22468 20402 22520 20408
rect 22756 20398 22784 21558
rect 22376 20392 22428 20398
rect 22376 20334 22428 20340
rect 22560 20392 22612 20398
rect 22744 20392 22796 20398
rect 22560 20334 22612 20340
rect 22664 20352 22744 20380
rect 22572 20058 22600 20334
rect 22560 20052 22612 20058
rect 22560 19994 22612 20000
rect 22664 19990 22692 20352
rect 22744 20334 22796 20340
rect 22836 20324 22888 20330
rect 22836 20266 22888 20272
rect 22744 20256 22796 20262
rect 22744 20198 22796 20204
rect 22376 19984 22428 19990
rect 22376 19926 22428 19932
rect 22652 19984 22704 19990
rect 22652 19926 22704 19932
rect 22284 19372 22336 19378
rect 22284 19314 22336 19320
rect 22296 18902 22324 19314
rect 22388 19310 22416 19926
rect 22652 19712 22704 19718
rect 22652 19654 22704 19660
rect 22664 19514 22692 19654
rect 22652 19508 22704 19514
rect 22652 19450 22704 19456
rect 22376 19304 22428 19310
rect 22376 19246 22428 19252
rect 22468 19168 22520 19174
rect 22468 19110 22520 19116
rect 22284 18896 22336 18902
rect 22284 18838 22336 18844
rect 22480 18834 22508 19110
rect 22468 18828 22520 18834
rect 22468 18770 22520 18776
rect 22560 18760 22612 18766
rect 22560 18702 22612 18708
rect 22468 18624 22520 18630
rect 22468 18566 22520 18572
rect 22480 18426 22508 18566
rect 22468 18420 22520 18426
rect 22468 18362 22520 18368
rect 22480 18272 22508 18362
rect 22572 18290 22600 18702
rect 22296 18244 22508 18272
rect 22560 18284 22612 18290
rect 22192 17740 22244 17746
rect 22192 17682 22244 17688
rect 22100 17604 22152 17610
rect 22100 17546 22152 17552
rect 22112 17338 22140 17546
rect 22100 17332 22152 17338
rect 22100 17274 22152 17280
rect 22296 17134 22324 18244
rect 22560 18226 22612 18232
rect 22664 18170 22692 19450
rect 22756 19310 22784 20198
rect 22848 19718 22876 20266
rect 23020 19780 23072 19786
rect 23020 19722 23072 19728
rect 22836 19712 22888 19718
rect 22836 19654 22888 19660
rect 23032 19514 23060 19722
rect 23020 19508 23072 19514
rect 23020 19450 23072 19456
rect 22836 19372 22888 19378
rect 22836 19314 22888 19320
rect 22744 19304 22796 19310
rect 22744 19246 22796 19252
rect 22744 18828 22796 18834
rect 22744 18770 22796 18776
rect 22756 18272 22784 18770
rect 22848 18630 22876 19314
rect 23020 19304 23072 19310
rect 23020 19246 23072 19252
rect 22928 19236 22980 19242
rect 22928 19178 22980 19184
rect 22940 18902 22968 19178
rect 23032 18970 23060 19246
rect 23020 18964 23072 18970
rect 23020 18906 23072 18912
rect 22928 18896 22980 18902
rect 22928 18838 22980 18844
rect 22836 18624 22888 18630
rect 22836 18566 22888 18572
rect 22756 18244 22968 18272
rect 22388 18154 22876 18170
rect 22376 18148 22888 18154
rect 22428 18142 22836 18148
rect 22376 18090 22428 18096
rect 22836 18090 22888 18096
rect 22940 17610 22968 18244
rect 22468 17604 22520 17610
rect 22468 17546 22520 17552
rect 22928 17604 22980 17610
rect 22928 17546 22980 17552
rect 22284 17128 22336 17134
rect 22284 17070 22336 17076
rect 22008 17060 22060 17066
rect 22008 17002 22060 17008
rect 22020 16794 22048 17002
rect 22376 16992 22428 16998
rect 22376 16934 22428 16940
rect 21916 16788 21968 16794
rect 21916 16730 21968 16736
rect 22008 16788 22060 16794
rect 22008 16730 22060 16736
rect 21548 16652 21600 16658
rect 21836 16646 21956 16674
rect 22388 16658 22416 16934
rect 21548 16594 21600 16600
rect 21456 16584 21508 16590
rect 21456 16526 21508 16532
rect 21468 16114 21496 16526
rect 21640 16516 21692 16522
rect 21640 16458 21692 16464
rect 21652 16114 21680 16458
rect 21456 16108 21508 16114
rect 21456 16050 21508 16056
rect 21640 16108 21692 16114
rect 21640 16050 21692 16056
rect 21732 16040 21784 16046
rect 21732 15982 21784 15988
rect 21824 16040 21876 16046
rect 21824 15982 21876 15988
rect 21744 15745 21772 15982
rect 21730 15736 21786 15745
rect 21730 15671 21786 15680
rect 21744 15502 21772 15671
rect 21836 15638 21864 15982
rect 21824 15632 21876 15638
rect 21824 15574 21876 15580
rect 21732 15496 21784 15502
rect 21732 15438 21784 15444
rect 21836 15162 21864 15574
rect 21824 15156 21876 15162
rect 21824 15098 21876 15104
rect 21928 15026 21956 16646
rect 22284 16652 22336 16658
rect 22284 16594 22336 16600
rect 22376 16652 22428 16658
rect 22376 16594 22428 16600
rect 22296 15978 22324 16594
rect 22388 16250 22416 16594
rect 22376 16244 22428 16250
rect 22376 16186 22428 16192
rect 22284 15972 22336 15978
rect 22284 15914 22336 15920
rect 22098 15736 22154 15745
rect 22008 15700 22060 15706
rect 22098 15671 22154 15680
rect 22008 15642 22060 15648
rect 22020 15366 22048 15642
rect 22112 15638 22140 15671
rect 22100 15632 22152 15638
rect 22100 15574 22152 15580
rect 22480 15570 22508 17546
rect 22928 17128 22980 17134
rect 22928 17070 22980 17076
rect 22940 16726 22968 17070
rect 22928 16720 22980 16726
rect 22928 16662 22980 16668
rect 22836 16652 22888 16658
rect 22836 16594 22888 16600
rect 22652 16584 22704 16590
rect 22652 16526 22704 16532
rect 22664 15978 22692 16526
rect 22652 15972 22704 15978
rect 22652 15914 22704 15920
rect 22664 15706 22692 15914
rect 22652 15700 22704 15706
rect 22652 15642 22704 15648
rect 22744 15632 22796 15638
rect 22664 15580 22744 15586
rect 22664 15574 22796 15580
rect 22468 15564 22520 15570
rect 22468 15506 22520 15512
rect 22664 15558 22784 15574
rect 22008 15360 22060 15366
rect 22008 15302 22060 15308
rect 21916 15020 21968 15026
rect 21916 14962 21968 14968
rect 21088 14476 21140 14482
rect 21088 14418 21140 14424
rect 21272 14476 21324 14482
rect 21272 14418 21324 14424
rect 20720 14272 20772 14278
rect 20720 14214 20772 14220
rect 20732 13938 20760 14214
rect 21100 14006 21128 14418
rect 21732 14408 21784 14414
rect 21732 14350 21784 14356
rect 21744 14074 21772 14350
rect 21364 14068 21416 14074
rect 21364 14010 21416 14016
rect 21732 14068 21784 14074
rect 21732 14010 21784 14016
rect 20996 14000 21048 14006
rect 20996 13942 21048 13948
rect 21088 14000 21140 14006
rect 21088 13942 21140 13948
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 20352 13864 20404 13870
rect 20352 13806 20404 13812
rect 20364 12986 20392 13806
rect 20546 13628 20854 13637
rect 20546 13626 20552 13628
rect 20608 13626 20632 13628
rect 20688 13626 20712 13628
rect 20768 13626 20792 13628
rect 20848 13626 20854 13628
rect 20608 13574 20610 13626
rect 20790 13574 20792 13626
rect 20546 13572 20552 13574
rect 20608 13572 20632 13574
rect 20688 13572 20712 13574
rect 20768 13572 20792 13574
rect 20848 13572 20854 13574
rect 20546 13563 20854 13572
rect 21008 13394 21036 13942
rect 21272 13796 21324 13802
rect 21272 13738 21324 13744
rect 21284 13530 21312 13738
rect 21272 13524 21324 13530
rect 21272 13466 21324 13472
rect 20996 13388 21048 13394
rect 20996 13330 21048 13336
rect 20720 13320 20772 13326
rect 20720 13262 20772 13268
rect 20352 12980 20404 12986
rect 20352 12922 20404 12928
rect 20732 12850 20760 13262
rect 20720 12844 20772 12850
rect 20720 12786 20772 12792
rect 20076 12640 20128 12646
rect 20076 12582 20128 12588
rect 19708 12368 19760 12374
rect 19708 12310 19760 12316
rect 20088 12238 20116 12582
rect 20546 12540 20854 12549
rect 20546 12538 20552 12540
rect 20608 12538 20632 12540
rect 20688 12538 20712 12540
rect 20768 12538 20792 12540
rect 20848 12538 20854 12540
rect 20608 12486 20610 12538
rect 20790 12486 20792 12538
rect 20546 12484 20552 12486
rect 20608 12484 20632 12486
rect 20688 12484 20712 12486
rect 20768 12484 20792 12486
rect 20848 12484 20854 12486
rect 20546 12475 20854 12484
rect 19708 12232 19760 12238
rect 19708 12174 19760 12180
rect 20076 12232 20128 12238
rect 20076 12174 20128 12180
rect 19156 12096 19208 12102
rect 19156 12038 19208 12044
rect 19168 11898 19196 12038
rect 19156 11892 19208 11898
rect 19156 11834 19208 11840
rect 19720 11694 19748 12174
rect 20996 11824 21048 11830
rect 20996 11766 21048 11772
rect 19064 11688 19116 11694
rect 19064 11630 19116 11636
rect 19708 11688 19760 11694
rect 19708 11630 19760 11636
rect 19984 11688 20036 11694
rect 19984 11630 20036 11636
rect 18880 11552 18932 11558
rect 18880 11494 18932 11500
rect 19616 11552 19668 11558
rect 19616 11494 19668 11500
rect 18420 11144 18472 11150
rect 18420 11086 18472 11092
rect 18432 10606 18460 11086
rect 18892 10810 18920 11494
rect 19628 11286 19656 11494
rect 19996 11354 20024 11630
rect 20352 11552 20404 11558
rect 20352 11494 20404 11500
rect 20904 11552 20956 11558
rect 20904 11494 20956 11500
rect 19984 11348 20036 11354
rect 19984 11290 20036 11296
rect 19616 11280 19668 11286
rect 19616 11222 19668 11228
rect 20076 11212 20128 11218
rect 20076 11154 20128 11160
rect 20088 10810 20116 11154
rect 18880 10804 18932 10810
rect 18880 10746 18932 10752
rect 20076 10804 20128 10810
rect 20076 10746 20128 10752
rect 18420 10600 18472 10606
rect 18420 10542 18472 10548
rect 18328 10260 18380 10266
rect 18328 10202 18380 10208
rect 18432 10198 18460 10542
rect 18512 10532 18564 10538
rect 18512 10474 18564 10480
rect 18420 10192 18472 10198
rect 18420 10134 18472 10140
rect 18144 10124 18196 10130
rect 18144 10066 18196 10072
rect 17776 10056 17828 10062
rect 17776 9998 17828 10004
rect 16396 9988 16448 9994
rect 16396 9930 16448 9936
rect 16304 9580 16356 9586
rect 16304 9522 16356 9528
rect 16408 9518 16436 9930
rect 17040 9920 17092 9926
rect 17040 9862 17092 9868
rect 15936 9512 15988 9518
rect 15856 9472 15936 9500
rect 15752 9376 15804 9382
rect 15752 9318 15804 9324
rect 15660 9036 15712 9042
rect 15580 8996 15660 9024
rect 15660 8978 15712 8984
rect 15764 8974 15792 9318
rect 15856 9042 15884 9472
rect 15936 9454 15988 9460
rect 16396 9512 16448 9518
rect 16396 9454 16448 9460
rect 16948 9444 17000 9450
rect 16948 9386 17000 9392
rect 15936 9376 15988 9382
rect 15936 9318 15988 9324
rect 15948 9042 15976 9318
rect 16304 9104 16356 9110
rect 16304 9046 16356 9052
rect 15844 9036 15896 9042
rect 15844 8978 15896 8984
rect 15936 9036 15988 9042
rect 15936 8978 15988 8984
rect 15752 8968 15804 8974
rect 15752 8910 15804 8916
rect 15108 8560 15160 8566
rect 15108 8502 15160 8508
rect 15120 7954 15148 8502
rect 15292 8424 15344 8430
rect 15384 8424 15436 8430
rect 15292 8366 15344 8372
rect 15382 8392 15384 8401
rect 15568 8424 15620 8430
rect 15436 8392 15438 8401
rect 15304 7954 15332 8366
rect 15568 8366 15620 8372
rect 15382 8327 15438 8336
rect 15580 8072 15608 8366
rect 15488 8044 15608 8072
rect 15108 7948 15160 7954
rect 15108 7890 15160 7896
rect 15292 7948 15344 7954
rect 15292 7890 15344 7896
rect 15016 7336 15068 7342
rect 15120 7324 15148 7890
rect 15068 7296 15148 7324
rect 15200 7336 15252 7342
rect 15016 7278 15068 7284
rect 15304 7324 15332 7890
rect 15488 7818 15516 8044
rect 15568 7948 15620 7954
rect 15568 7890 15620 7896
rect 15660 7948 15712 7954
rect 15660 7890 15712 7896
rect 15476 7812 15528 7818
rect 15476 7754 15528 7760
rect 15580 7342 15608 7890
rect 15672 7546 15700 7890
rect 16316 7546 16344 9046
rect 16764 8968 16816 8974
rect 16764 8910 16816 8916
rect 16488 8424 16540 8430
rect 16488 8366 16540 8372
rect 16396 8288 16448 8294
rect 16396 8230 16448 8236
rect 16408 7954 16436 8230
rect 16396 7948 16448 7954
rect 16396 7890 16448 7896
rect 16500 7546 16528 8366
rect 15660 7540 15712 7546
rect 15660 7482 15712 7488
rect 16304 7540 16356 7546
rect 16304 7482 16356 7488
rect 16488 7540 16540 7546
rect 16488 7482 16540 7488
rect 15252 7296 15332 7324
rect 15568 7336 15620 7342
rect 15200 7278 15252 7284
rect 15568 7278 15620 7284
rect 16212 7200 16264 7206
rect 16212 7142 16264 7148
rect 16224 7002 16252 7142
rect 16212 6996 16264 7002
rect 16212 6938 16264 6944
rect 16316 6458 16344 7482
rect 16672 7268 16724 7274
rect 16672 7210 16724 7216
rect 16684 6866 16712 7210
rect 16672 6860 16724 6866
rect 16672 6802 16724 6808
rect 16304 6452 16356 6458
rect 16304 6394 16356 6400
rect 15752 6384 15804 6390
rect 15752 6326 15804 6332
rect 15292 6180 15344 6186
rect 15292 6122 15344 6128
rect 15476 6180 15528 6186
rect 15476 6122 15528 6128
rect 15200 6112 15252 6118
rect 15200 6054 15252 6060
rect 15212 5370 15240 6054
rect 15200 5364 15252 5370
rect 15200 5306 15252 5312
rect 15304 5250 15332 6122
rect 15488 5914 15516 6122
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 15476 5908 15528 5914
rect 15476 5850 15528 5856
rect 15580 5846 15608 6054
rect 15568 5840 15620 5846
rect 15568 5782 15620 5788
rect 15476 5772 15528 5778
rect 15476 5714 15528 5720
rect 15488 5370 15516 5714
rect 15476 5364 15528 5370
rect 15476 5306 15528 5312
rect 15212 5222 15332 5250
rect 15580 5234 15608 5782
rect 15764 5710 15792 6326
rect 16580 6248 16632 6254
rect 16580 6190 16632 6196
rect 16028 6112 16080 6118
rect 16028 6054 16080 6060
rect 16488 6112 16540 6118
rect 16488 6054 16540 6060
rect 16040 5778 16068 6054
rect 16500 5914 16528 6054
rect 16488 5908 16540 5914
rect 16488 5850 16540 5856
rect 16028 5772 16080 5778
rect 16028 5714 16080 5720
rect 15752 5704 15804 5710
rect 15752 5646 15804 5652
rect 15764 5370 15792 5646
rect 16592 5574 16620 6190
rect 16304 5568 16356 5574
rect 16304 5510 16356 5516
rect 16580 5568 16632 5574
rect 16580 5510 16632 5516
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 15568 5228 15620 5234
rect 15212 5030 15240 5222
rect 15568 5170 15620 5176
rect 16316 5166 16344 5510
rect 16304 5160 16356 5166
rect 16304 5102 16356 5108
rect 15200 5024 15252 5030
rect 15200 4966 15252 4972
rect 16304 4480 16356 4486
rect 16304 4422 16356 4428
rect 16316 4146 16344 4422
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16776 4078 16804 8910
rect 16856 8832 16908 8838
rect 16856 8774 16908 8780
rect 15476 4072 15528 4078
rect 15476 4014 15528 4020
rect 15936 4072 15988 4078
rect 15936 4014 15988 4020
rect 16488 4072 16540 4078
rect 16488 4014 16540 4020
rect 16764 4072 16816 4078
rect 16764 4014 16816 4020
rect 15200 3936 15252 3942
rect 14936 3884 15200 3890
rect 14936 3878 15252 3884
rect 14936 3862 15240 3878
rect 15488 3738 15516 4014
rect 15948 3738 15976 4014
rect 16304 3936 16356 3942
rect 16304 3878 16356 3884
rect 15476 3732 15528 3738
rect 15476 3674 15528 3680
rect 15936 3732 15988 3738
rect 15936 3674 15988 3680
rect 15108 3664 15160 3670
rect 15108 3606 15160 3612
rect 14832 3188 14884 3194
rect 14832 3130 14884 3136
rect 14740 3120 14792 3126
rect 14740 3062 14792 3068
rect 14280 2984 14332 2990
rect 14280 2926 14332 2932
rect 14464 2984 14516 2990
rect 14464 2926 14516 2932
rect 14188 2848 14240 2854
rect 14188 2790 14240 2796
rect 13830 2748 14138 2757
rect 13830 2746 13836 2748
rect 13892 2746 13916 2748
rect 13972 2746 13996 2748
rect 14052 2746 14076 2748
rect 14132 2746 14138 2748
rect 13892 2694 13894 2746
rect 14074 2694 14076 2746
rect 13830 2692 13836 2694
rect 13892 2692 13916 2694
rect 13972 2692 13996 2694
rect 14052 2692 14076 2694
rect 14132 2692 14138 2694
rect 13830 2683 14138 2692
rect 14200 1986 14228 2790
rect 14292 2514 14320 2926
rect 14280 2508 14332 2514
rect 14280 2450 14332 2456
rect 14200 1958 14320 1986
rect 14476 1970 14504 2926
rect 14188 1896 14240 1902
rect 14188 1838 14240 1844
rect 13830 1660 14138 1669
rect 13830 1658 13836 1660
rect 13892 1658 13916 1660
rect 13972 1658 13996 1660
rect 14052 1658 14076 1660
rect 14132 1658 14138 1660
rect 13892 1606 13894 1658
rect 14074 1606 14076 1658
rect 13830 1604 13836 1606
rect 13892 1604 13916 1606
rect 13972 1604 13996 1606
rect 14052 1604 14076 1606
rect 14132 1604 14138 1606
rect 13830 1595 14138 1604
rect 13544 1420 13596 1426
rect 13544 1362 13596 1368
rect 13728 1420 13780 1426
rect 13728 1362 13780 1368
rect 13360 1352 13412 1358
rect 13360 1294 13412 1300
rect 13372 1018 13400 1294
rect 13728 1216 13780 1222
rect 13728 1158 13780 1164
rect 13360 1012 13412 1018
rect 13360 954 13412 960
rect 13176 808 13228 814
rect 13176 750 13228 756
rect 13360 808 13412 814
rect 13360 750 13412 756
rect 13372 400 13400 750
rect 13740 456 13768 1158
rect 14200 814 14228 1838
rect 14292 814 14320 1958
rect 14464 1964 14516 1970
rect 14464 1906 14516 1912
rect 14556 1896 14608 1902
rect 14556 1838 14608 1844
rect 14568 1426 14596 1838
rect 14844 1426 14872 3130
rect 15120 2961 15148 3606
rect 16316 3602 16344 3878
rect 16500 3738 16528 4014
rect 16488 3732 16540 3738
rect 16488 3674 16540 3680
rect 15384 3596 15436 3602
rect 15384 3538 15436 3544
rect 16304 3596 16356 3602
rect 16304 3538 16356 3544
rect 15396 3194 15424 3538
rect 16304 3460 16356 3466
rect 16304 3402 16356 3408
rect 15476 3392 15528 3398
rect 15476 3334 15528 3340
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 15488 3126 15516 3334
rect 15476 3120 15528 3126
rect 15382 3088 15438 3097
rect 15476 3062 15528 3068
rect 15382 3023 15384 3032
rect 15436 3023 15438 3032
rect 15384 2994 15436 3000
rect 15936 2984 15988 2990
rect 15106 2952 15162 2961
rect 15936 2926 15988 2932
rect 15106 2887 15108 2896
rect 15160 2887 15162 2896
rect 15108 2858 15160 2864
rect 15948 2650 15976 2926
rect 16120 2848 16172 2854
rect 16120 2790 16172 2796
rect 15936 2644 15988 2650
rect 15936 2586 15988 2592
rect 16132 2514 16160 2790
rect 16316 2514 16344 3402
rect 16396 3392 16448 3398
rect 16396 3334 16448 3340
rect 16408 3058 16436 3334
rect 16396 3052 16448 3058
rect 16396 2994 16448 3000
rect 16868 2990 16896 8774
rect 16960 8498 16988 9386
rect 17052 8974 17080 9862
rect 17188 9820 17496 9829
rect 17188 9818 17194 9820
rect 17250 9818 17274 9820
rect 17330 9818 17354 9820
rect 17410 9818 17434 9820
rect 17490 9818 17496 9820
rect 17250 9766 17252 9818
rect 17432 9766 17434 9818
rect 17188 9764 17194 9766
rect 17250 9764 17274 9766
rect 17330 9764 17354 9766
rect 17410 9764 17434 9766
rect 17490 9764 17496 9766
rect 17188 9755 17496 9764
rect 18156 9081 18184 10066
rect 18524 10062 18552 10474
rect 18892 10266 18920 10746
rect 19892 10532 19944 10538
rect 19892 10474 19944 10480
rect 18880 10260 18932 10266
rect 18880 10202 18932 10208
rect 18512 10056 18564 10062
rect 18512 9998 18564 10004
rect 18236 9716 18288 9722
rect 18236 9658 18288 9664
rect 18142 9072 18198 9081
rect 17592 9036 17644 9042
rect 18142 9007 18198 9016
rect 17592 8978 17644 8984
rect 17040 8968 17092 8974
rect 17040 8910 17092 8916
rect 16948 8492 17000 8498
rect 16948 8434 17000 8440
rect 17052 8022 17080 8910
rect 17188 8732 17496 8741
rect 17188 8730 17194 8732
rect 17250 8730 17274 8732
rect 17330 8730 17354 8732
rect 17410 8730 17434 8732
rect 17490 8730 17496 8732
rect 17250 8678 17252 8730
rect 17432 8678 17434 8730
rect 17188 8676 17194 8678
rect 17250 8676 17274 8678
rect 17330 8676 17354 8678
rect 17410 8676 17434 8678
rect 17490 8676 17496 8678
rect 17188 8667 17496 8676
rect 17604 8634 17632 8978
rect 17592 8628 17644 8634
rect 17592 8570 17644 8576
rect 17960 8560 18012 8566
rect 17880 8520 17960 8548
rect 17040 8016 17092 8022
rect 17040 7958 17092 7964
rect 17684 7880 17736 7886
rect 17684 7822 17736 7828
rect 17188 7644 17496 7653
rect 17188 7642 17194 7644
rect 17250 7642 17274 7644
rect 17330 7642 17354 7644
rect 17410 7642 17434 7644
rect 17490 7642 17496 7644
rect 17250 7590 17252 7642
rect 17432 7590 17434 7642
rect 17188 7588 17194 7590
rect 17250 7588 17274 7590
rect 17330 7588 17354 7590
rect 17410 7588 17434 7590
rect 17490 7588 17496 7590
rect 17188 7579 17496 7588
rect 16948 7336 17000 7342
rect 16948 7278 17000 7284
rect 17040 7336 17092 7342
rect 17040 7278 17092 7284
rect 17132 7336 17184 7342
rect 17132 7278 17184 7284
rect 16960 6866 16988 7278
rect 17052 6866 17080 7278
rect 16948 6860 17000 6866
rect 16948 6802 17000 6808
rect 17040 6860 17092 6866
rect 17040 6802 17092 6808
rect 17052 6254 17080 6802
rect 17144 6798 17172 7278
rect 17696 6934 17724 7822
rect 17776 7744 17828 7750
rect 17776 7686 17828 7692
rect 17788 7274 17816 7686
rect 17880 7478 17908 8520
rect 17960 8502 18012 8508
rect 18144 7812 18196 7818
rect 18144 7754 18196 7760
rect 17868 7472 17920 7478
rect 17868 7414 17920 7420
rect 17960 7472 18012 7478
rect 17960 7414 18012 7420
rect 17776 7268 17828 7274
rect 17776 7210 17828 7216
rect 17684 6928 17736 6934
rect 17684 6870 17736 6876
rect 17788 6866 17816 7210
rect 17972 6866 18000 7414
rect 18156 7342 18184 7754
rect 18248 7426 18276 9658
rect 18696 9512 18748 9518
rect 18696 9454 18748 9460
rect 19524 9512 19576 9518
rect 19524 9454 19576 9460
rect 18708 9110 18736 9454
rect 18788 9376 18840 9382
rect 18788 9318 18840 9324
rect 18696 9104 18748 9110
rect 18696 9046 18748 9052
rect 18708 8634 18736 9046
rect 18696 8628 18748 8634
rect 18696 8570 18748 8576
rect 18696 8424 18748 8430
rect 18696 8366 18748 8372
rect 18328 8356 18380 8362
rect 18328 8298 18380 8304
rect 18340 8090 18368 8298
rect 18328 8084 18380 8090
rect 18328 8026 18380 8032
rect 18420 7744 18472 7750
rect 18420 7686 18472 7692
rect 18432 7546 18460 7686
rect 18420 7540 18472 7546
rect 18420 7482 18472 7488
rect 18248 7398 18368 7426
rect 18144 7336 18196 7342
rect 18144 7278 18196 7284
rect 18236 7336 18288 7342
rect 18236 7278 18288 7284
rect 18248 7188 18276 7278
rect 18064 7160 18276 7188
rect 17776 6860 17828 6866
rect 17776 6802 17828 6808
rect 17960 6860 18012 6866
rect 17960 6802 18012 6808
rect 18064 6798 18092 7160
rect 17132 6792 17184 6798
rect 17132 6734 17184 6740
rect 17684 6792 17736 6798
rect 17684 6734 17736 6740
rect 18052 6792 18104 6798
rect 18052 6734 18104 6740
rect 18144 6792 18196 6798
rect 18144 6734 18196 6740
rect 17592 6724 17644 6730
rect 17592 6666 17644 6672
rect 17188 6556 17496 6565
rect 17188 6554 17194 6556
rect 17250 6554 17274 6556
rect 17330 6554 17354 6556
rect 17410 6554 17434 6556
rect 17490 6554 17496 6556
rect 17250 6502 17252 6554
rect 17432 6502 17434 6554
rect 17188 6500 17194 6502
rect 17250 6500 17274 6502
rect 17330 6500 17354 6502
rect 17410 6500 17434 6502
rect 17490 6500 17496 6502
rect 17188 6491 17496 6500
rect 17040 6248 17092 6254
rect 17040 6190 17092 6196
rect 17132 6248 17184 6254
rect 17132 6190 17184 6196
rect 17144 6100 17172 6190
rect 17604 6118 17632 6666
rect 17052 6072 17172 6100
rect 17224 6112 17276 6118
rect 17052 3942 17080 6072
rect 17224 6054 17276 6060
rect 17592 6112 17644 6118
rect 17592 6054 17644 6060
rect 17236 5846 17264 6054
rect 17224 5840 17276 5846
rect 17224 5782 17276 5788
rect 17188 5468 17496 5477
rect 17188 5466 17194 5468
rect 17250 5466 17274 5468
rect 17330 5466 17354 5468
rect 17410 5466 17434 5468
rect 17490 5466 17496 5468
rect 17250 5414 17252 5466
rect 17432 5414 17434 5466
rect 17188 5412 17194 5414
rect 17250 5412 17274 5414
rect 17330 5412 17354 5414
rect 17410 5412 17434 5414
rect 17490 5412 17496 5414
rect 17188 5403 17496 5412
rect 17188 4380 17496 4389
rect 17188 4378 17194 4380
rect 17250 4378 17274 4380
rect 17330 4378 17354 4380
rect 17410 4378 17434 4380
rect 17490 4378 17496 4380
rect 17250 4326 17252 4378
rect 17432 4326 17434 4378
rect 17188 4324 17194 4326
rect 17250 4324 17274 4326
rect 17330 4324 17354 4326
rect 17410 4324 17434 4326
rect 17490 4324 17496 4326
rect 17188 4315 17496 4324
rect 17408 4004 17460 4010
rect 17408 3946 17460 3952
rect 17040 3936 17092 3942
rect 17040 3878 17092 3884
rect 17420 3738 17448 3946
rect 17408 3732 17460 3738
rect 17408 3674 17460 3680
rect 17040 3664 17092 3670
rect 17040 3606 17092 3612
rect 16856 2984 16908 2990
rect 16856 2926 16908 2932
rect 15476 2508 15528 2514
rect 15476 2450 15528 2456
rect 16120 2508 16172 2514
rect 16120 2450 16172 2456
rect 16304 2508 16356 2514
rect 16304 2450 16356 2456
rect 15200 2304 15252 2310
rect 15200 2246 15252 2252
rect 15212 1970 15240 2246
rect 15200 1964 15252 1970
rect 15200 1906 15252 1912
rect 15488 1902 15516 2450
rect 16304 2304 16356 2310
rect 16304 2246 16356 2252
rect 16580 2304 16632 2310
rect 16580 2246 16632 2252
rect 15476 1896 15528 1902
rect 15476 1838 15528 1844
rect 16120 1896 16172 1902
rect 16120 1838 16172 1844
rect 14464 1420 14516 1426
rect 14464 1362 14516 1368
rect 14556 1420 14608 1426
rect 14556 1362 14608 1368
rect 14832 1420 14884 1426
rect 14832 1362 14884 1368
rect 15568 1420 15620 1426
rect 15568 1362 15620 1368
rect 14188 808 14240 814
rect 14188 750 14240 756
rect 14280 808 14332 814
rect 14280 750 14332 756
rect 13830 572 14138 581
rect 13830 570 13836 572
rect 13892 570 13916 572
rect 13972 570 13996 572
rect 14052 570 14076 572
rect 14132 570 14138 572
rect 13892 518 13894 570
rect 14074 518 14076 570
rect 13830 516 13836 518
rect 13892 516 13916 518
rect 13972 516 13996 518
rect 14052 516 14076 518
rect 14132 516 14138 518
rect 13830 507 14138 516
rect 13740 428 13952 456
rect 13924 400 13952 428
rect 14476 400 14504 1362
rect 15016 808 15068 814
rect 15016 750 15068 756
rect 15028 400 15056 750
rect 15580 400 15608 1362
rect 16132 400 16160 1838
rect 16316 1426 16344 2246
rect 16396 1896 16448 1902
rect 16396 1838 16448 1844
rect 16304 1420 16356 1426
rect 16304 1362 16356 1368
rect 16408 814 16436 1838
rect 16592 814 16620 2246
rect 17052 1494 17080 3606
rect 17188 3292 17496 3301
rect 17188 3290 17194 3292
rect 17250 3290 17274 3292
rect 17330 3290 17354 3292
rect 17410 3290 17434 3292
rect 17490 3290 17496 3292
rect 17250 3238 17252 3290
rect 17432 3238 17434 3290
rect 17188 3236 17194 3238
rect 17250 3236 17274 3238
rect 17330 3236 17354 3238
rect 17410 3236 17434 3238
rect 17490 3236 17496 3238
rect 17188 3227 17496 3236
rect 17696 3126 17724 6734
rect 17868 6248 17920 6254
rect 17868 6190 17920 6196
rect 17776 6180 17828 6186
rect 17776 6122 17828 6128
rect 17788 5846 17816 6122
rect 17880 5846 17908 6190
rect 17776 5840 17828 5846
rect 17776 5782 17828 5788
rect 17868 5840 17920 5846
rect 17868 5782 17920 5788
rect 17880 5302 17908 5782
rect 17960 5636 18012 5642
rect 17960 5578 18012 5584
rect 17868 5296 17920 5302
rect 17868 5238 17920 5244
rect 17972 4690 18000 5578
rect 18156 5370 18184 6734
rect 18144 5364 18196 5370
rect 18144 5306 18196 5312
rect 18340 5234 18368 7398
rect 18420 6860 18472 6866
rect 18420 6802 18472 6808
rect 18432 6662 18460 6802
rect 18420 6656 18472 6662
rect 18420 6598 18472 6604
rect 18328 5228 18380 5234
rect 18328 5170 18380 5176
rect 18144 5160 18196 5166
rect 18144 5102 18196 5108
rect 18052 5024 18104 5030
rect 18052 4966 18104 4972
rect 18064 4690 18092 4966
rect 17960 4684 18012 4690
rect 17960 4626 18012 4632
rect 18052 4684 18104 4690
rect 18052 4626 18104 4632
rect 17868 3936 17920 3942
rect 17868 3878 17920 3884
rect 17880 3670 17908 3878
rect 17868 3664 17920 3670
rect 17868 3606 17920 3612
rect 18156 3534 18184 5102
rect 18340 4146 18368 5170
rect 18708 4826 18736 8366
rect 18800 7886 18828 9318
rect 19064 8968 19116 8974
rect 19064 8910 19116 8916
rect 19248 8968 19300 8974
rect 19248 8910 19300 8916
rect 19432 8968 19484 8974
rect 19432 8910 19484 8916
rect 18880 8832 18932 8838
rect 18880 8774 18932 8780
rect 18892 8430 18920 8774
rect 19076 8430 19104 8910
rect 19260 8566 19288 8910
rect 19248 8560 19300 8566
rect 19248 8502 19300 8508
rect 19444 8498 19472 8910
rect 19536 8634 19564 9454
rect 19616 9376 19668 9382
rect 19616 9318 19668 9324
rect 19628 9110 19656 9318
rect 19616 9104 19668 9110
rect 19616 9046 19668 9052
rect 19524 8628 19576 8634
rect 19524 8570 19576 8576
rect 19432 8492 19484 8498
rect 19432 8434 19484 8440
rect 19628 8430 19656 9046
rect 19904 8974 19932 10474
rect 20088 10130 20116 10746
rect 20364 10606 20392 11494
rect 20546 11452 20854 11461
rect 20546 11450 20552 11452
rect 20608 11450 20632 11452
rect 20688 11450 20712 11452
rect 20768 11450 20792 11452
rect 20848 11450 20854 11452
rect 20608 11398 20610 11450
rect 20790 11398 20792 11450
rect 20546 11396 20552 11398
rect 20608 11396 20632 11398
rect 20688 11396 20712 11398
rect 20768 11396 20792 11398
rect 20848 11396 20854 11398
rect 20546 11387 20854 11396
rect 20444 11348 20496 11354
rect 20444 11290 20496 11296
rect 20456 11014 20484 11290
rect 20812 11280 20864 11286
rect 20916 11268 20944 11494
rect 20864 11240 20944 11268
rect 20812 11222 20864 11228
rect 20444 11008 20496 11014
rect 20444 10950 20496 10956
rect 20456 10742 20484 10950
rect 20444 10736 20496 10742
rect 20444 10678 20496 10684
rect 21008 10606 21036 11766
rect 21088 11756 21140 11762
rect 21088 11698 21140 11704
rect 21100 10810 21128 11698
rect 21088 10804 21140 10810
rect 21088 10746 21140 10752
rect 20352 10600 20404 10606
rect 20352 10542 20404 10548
rect 20996 10600 21048 10606
rect 20996 10542 21048 10548
rect 20546 10364 20854 10373
rect 20546 10362 20552 10364
rect 20608 10362 20632 10364
rect 20688 10362 20712 10364
rect 20768 10362 20792 10364
rect 20848 10362 20854 10364
rect 20608 10310 20610 10362
rect 20790 10310 20792 10362
rect 20546 10308 20552 10310
rect 20608 10308 20632 10310
rect 20688 10308 20712 10310
rect 20768 10308 20792 10310
rect 20848 10308 20854 10310
rect 20546 10299 20854 10308
rect 20076 10124 20128 10130
rect 20076 10066 20128 10072
rect 20996 9512 21048 9518
rect 20996 9454 21048 9460
rect 19984 9444 20036 9450
rect 19984 9386 20036 9392
rect 19996 9178 20024 9386
rect 20546 9276 20854 9285
rect 20546 9274 20552 9276
rect 20608 9274 20632 9276
rect 20688 9274 20712 9276
rect 20768 9274 20792 9276
rect 20848 9274 20854 9276
rect 20608 9222 20610 9274
rect 20790 9222 20792 9274
rect 20546 9220 20552 9222
rect 20608 9220 20632 9222
rect 20688 9220 20712 9222
rect 20768 9220 20792 9222
rect 20848 9220 20854 9222
rect 20546 9211 20854 9220
rect 19984 9172 20036 9178
rect 19984 9114 20036 9120
rect 21008 9110 21036 9454
rect 21376 9382 21404 14010
rect 21928 13870 21956 14962
rect 22100 14952 22152 14958
rect 22100 14894 22152 14900
rect 22112 14550 22140 14894
rect 22100 14544 22152 14550
rect 22100 14486 22152 14492
rect 22008 14340 22060 14346
rect 22008 14282 22060 14288
rect 21916 13864 21968 13870
rect 21916 13806 21968 13812
rect 21456 13388 21508 13394
rect 21456 13330 21508 13336
rect 21548 13388 21600 13394
rect 21548 13330 21600 13336
rect 21468 12782 21496 13330
rect 21456 12776 21508 12782
rect 21456 12718 21508 12724
rect 21560 11286 21588 13330
rect 21824 12776 21876 12782
rect 21824 12718 21876 12724
rect 21640 12300 21692 12306
rect 21640 12242 21692 12248
rect 21548 11280 21600 11286
rect 21548 11222 21600 11228
rect 21560 10198 21588 11222
rect 21652 11014 21680 12242
rect 21836 11898 21864 12718
rect 22020 12434 22048 14282
rect 22112 14074 22140 14486
rect 22100 14068 22152 14074
rect 22100 14010 22152 14016
rect 22112 13326 22140 14010
rect 22192 13796 22244 13802
rect 22192 13738 22244 13744
rect 22204 13530 22232 13738
rect 22192 13524 22244 13530
rect 22192 13466 22244 13472
rect 22480 13394 22508 15506
rect 22560 15360 22612 15366
rect 22560 15302 22612 15308
rect 22572 14890 22600 15302
rect 22560 14884 22612 14890
rect 22560 14826 22612 14832
rect 22664 14482 22692 15558
rect 22848 14958 22876 16594
rect 22940 15434 22968 16662
rect 23020 16652 23072 16658
rect 23020 16594 23072 16600
rect 23032 16250 23060 16594
rect 23020 16244 23072 16250
rect 23020 16186 23072 16192
rect 22928 15428 22980 15434
rect 22928 15370 22980 15376
rect 22836 14952 22888 14958
rect 22836 14894 22888 14900
rect 23020 14544 23072 14550
rect 23020 14486 23072 14492
rect 22652 14476 22704 14482
rect 22652 14418 22704 14424
rect 22468 13388 22520 13394
rect 22468 13330 22520 13336
rect 22100 13320 22152 13326
rect 22100 13262 22152 13268
rect 22664 12850 22692 14418
rect 22744 13456 22796 13462
rect 22744 13398 22796 13404
rect 22652 12844 22704 12850
rect 22652 12786 22704 12792
rect 22756 12714 22784 13398
rect 23032 13258 23060 14486
rect 23020 13252 23072 13258
rect 23020 13194 23072 13200
rect 23032 12986 23060 13194
rect 22836 12980 22888 12986
rect 22836 12922 22888 12928
rect 23020 12980 23072 12986
rect 23020 12922 23072 12928
rect 22744 12708 22796 12714
rect 22744 12650 22796 12656
rect 22652 12640 22704 12646
rect 22652 12582 22704 12588
rect 22664 12442 22692 12582
rect 21928 12406 22048 12434
rect 22652 12436 22704 12442
rect 21824 11892 21876 11898
rect 21824 11834 21876 11840
rect 21732 11688 21784 11694
rect 21732 11630 21784 11636
rect 21744 11354 21772 11630
rect 21732 11348 21784 11354
rect 21732 11290 21784 11296
rect 21640 11008 21692 11014
rect 21640 10950 21692 10956
rect 21548 10192 21600 10198
rect 21548 10134 21600 10140
rect 21928 9450 21956 12406
rect 22652 12378 22704 12384
rect 22468 12300 22520 12306
rect 22468 12242 22520 12248
rect 22100 12232 22152 12238
rect 22100 12174 22152 12180
rect 22112 11762 22140 12174
rect 22100 11756 22152 11762
rect 22100 11698 22152 11704
rect 22008 11620 22060 11626
rect 22008 11562 22060 11568
rect 22020 11354 22048 11562
rect 22008 11348 22060 11354
rect 22008 11290 22060 11296
rect 22008 11212 22060 11218
rect 22008 11154 22060 11160
rect 22020 10606 22048 11154
rect 22112 10674 22140 11698
rect 22284 11688 22336 11694
rect 22284 11630 22336 11636
rect 22376 11688 22428 11694
rect 22376 11630 22428 11636
rect 22192 11008 22244 11014
rect 22192 10950 22244 10956
rect 22100 10668 22152 10674
rect 22100 10610 22152 10616
rect 22008 10600 22060 10606
rect 22008 10542 22060 10548
rect 21916 9444 21968 9450
rect 21916 9386 21968 9392
rect 21364 9376 21416 9382
rect 21364 9318 21416 9324
rect 20996 9104 21048 9110
rect 20996 9046 21048 9052
rect 21272 9104 21324 9110
rect 21272 9046 21324 9052
rect 20168 9036 20220 9042
rect 20168 8978 20220 8984
rect 20444 9036 20496 9042
rect 20444 8978 20496 8984
rect 19892 8968 19944 8974
rect 19892 8910 19944 8916
rect 20076 8968 20128 8974
rect 20076 8910 20128 8916
rect 19892 8832 19944 8838
rect 19892 8774 19944 8780
rect 19904 8430 19932 8774
rect 20088 8430 20116 8910
rect 20180 8498 20208 8978
rect 20456 8634 20484 8978
rect 20812 8900 20864 8906
rect 20812 8842 20864 8848
rect 20444 8628 20496 8634
rect 20444 8570 20496 8576
rect 20168 8492 20220 8498
rect 20168 8434 20220 8440
rect 18880 8424 18932 8430
rect 18880 8366 18932 8372
rect 19064 8424 19116 8430
rect 19064 8366 19116 8372
rect 19616 8424 19668 8430
rect 19616 8366 19668 8372
rect 19892 8424 19944 8430
rect 19892 8366 19944 8372
rect 20076 8424 20128 8430
rect 20076 8366 20128 8372
rect 19616 7948 19668 7954
rect 19616 7890 19668 7896
rect 18788 7880 18840 7886
rect 18788 7822 18840 7828
rect 18800 7410 18828 7822
rect 19524 7812 19576 7818
rect 19524 7754 19576 7760
rect 18880 7744 18932 7750
rect 18880 7686 18932 7692
rect 18892 7546 18920 7686
rect 19536 7546 19564 7754
rect 18880 7540 18932 7546
rect 18880 7482 18932 7488
rect 19524 7540 19576 7546
rect 19524 7482 19576 7488
rect 18788 7404 18840 7410
rect 18788 7346 18840 7352
rect 19064 7268 19116 7274
rect 19064 7210 19116 7216
rect 19076 7002 19104 7210
rect 19536 7206 19564 7482
rect 19628 7478 19656 7890
rect 19708 7880 19760 7886
rect 19708 7822 19760 7828
rect 19616 7472 19668 7478
rect 19616 7414 19668 7420
rect 19524 7200 19576 7206
rect 19524 7142 19576 7148
rect 19628 7002 19656 7414
rect 19720 7342 19748 7822
rect 19708 7336 19760 7342
rect 19708 7278 19760 7284
rect 19720 7002 19748 7278
rect 19064 6996 19116 7002
rect 19064 6938 19116 6944
rect 19616 6996 19668 7002
rect 19616 6938 19668 6944
rect 19708 6996 19760 7002
rect 19708 6938 19760 6944
rect 19708 5704 19760 5710
rect 19708 5646 19760 5652
rect 18880 5568 18932 5574
rect 18880 5510 18932 5516
rect 19340 5568 19392 5574
rect 19340 5510 19392 5516
rect 18892 5234 18920 5510
rect 18880 5228 18932 5234
rect 18880 5170 18932 5176
rect 19156 5160 19208 5166
rect 19156 5102 19208 5108
rect 19168 4826 19196 5102
rect 18696 4820 18748 4826
rect 18696 4762 18748 4768
rect 19156 4820 19208 4826
rect 19156 4762 19208 4768
rect 19352 4758 19380 5510
rect 19720 5302 19748 5646
rect 19708 5296 19760 5302
rect 19708 5238 19760 5244
rect 19904 5030 19932 8366
rect 20088 7954 20116 8366
rect 20180 7970 20208 8434
rect 20824 8430 20852 8842
rect 20812 8424 20864 8430
rect 20864 8384 20944 8412
rect 20812 8366 20864 8372
rect 20546 8188 20854 8197
rect 20546 8186 20552 8188
rect 20608 8186 20632 8188
rect 20688 8186 20712 8188
rect 20768 8186 20792 8188
rect 20848 8186 20854 8188
rect 20608 8134 20610 8186
rect 20790 8134 20792 8186
rect 20546 8132 20552 8134
rect 20608 8132 20632 8134
rect 20688 8132 20712 8134
rect 20768 8132 20792 8134
rect 20848 8132 20854 8134
rect 20546 8123 20854 8132
rect 20916 8090 20944 8384
rect 20904 8084 20956 8090
rect 20904 8026 20956 8032
rect 20180 7954 20300 7970
rect 20076 7948 20128 7954
rect 20180 7948 20312 7954
rect 20180 7942 20260 7948
rect 20076 7890 20128 7896
rect 20260 7890 20312 7896
rect 20904 7948 20956 7954
rect 20904 7890 20956 7896
rect 19984 7880 20036 7886
rect 19984 7822 20036 7828
rect 19996 7342 20024 7822
rect 20088 7342 20116 7890
rect 20916 7818 20944 7890
rect 21284 7886 21312 9046
rect 21376 9042 21404 9318
rect 21364 9036 21416 9042
rect 21364 8978 21416 8984
rect 21824 9036 21876 9042
rect 21824 8978 21876 8984
rect 21640 8424 21692 8430
rect 21640 8366 21692 8372
rect 21732 8424 21784 8430
rect 21732 8366 21784 8372
rect 21364 8288 21416 8294
rect 21364 8230 21416 8236
rect 21548 8288 21600 8294
rect 21548 8230 21600 8236
rect 21376 7954 21404 8230
rect 21560 7954 21588 8230
rect 21364 7948 21416 7954
rect 21364 7890 21416 7896
rect 21548 7948 21600 7954
rect 21548 7890 21600 7896
rect 21272 7880 21324 7886
rect 21272 7822 21324 7828
rect 20904 7812 20956 7818
rect 20904 7754 20956 7760
rect 20916 7546 20944 7754
rect 20904 7540 20956 7546
rect 20904 7482 20956 7488
rect 19984 7336 20036 7342
rect 19984 7278 20036 7284
rect 20076 7336 20128 7342
rect 20076 7278 20128 7284
rect 21180 7268 21232 7274
rect 21180 7210 21232 7216
rect 20546 7100 20854 7109
rect 20546 7098 20552 7100
rect 20608 7098 20632 7100
rect 20688 7098 20712 7100
rect 20768 7098 20792 7100
rect 20848 7098 20854 7100
rect 20608 7046 20610 7098
rect 20790 7046 20792 7098
rect 20546 7044 20552 7046
rect 20608 7044 20632 7046
rect 20688 7044 20712 7046
rect 20768 7044 20792 7046
rect 20848 7044 20854 7046
rect 20546 7035 20854 7044
rect 21192 6934 21220 7210
rect 21180 6928 21232 6934
rect 21180 6870 21232 6876
rect 20260 6860 20312 6866
rect 20260 6802 20312 6808
rect 19984 5772 20036 5778
rect 19984 5714 20036 5720
rect 19892 5024 19944 5030
rect 19892 4966 19944 4972
rect 19340 4752 19392 4758
rect 19340 4694 19392 4700
rect 18972 4684 19024 4690
rect 18972 4626 19024 4632
rect 18984 4282 19012 4626
rect 18972 4276 19024 4282
rect 18972 4218 19024 4224
rect 19248 4208 19300 4214
rect 19248 4150 19300 4156
rect 18328 4140 18380 4146
rect 18328 4082 18380 4088
rect 18236 4072 18288 4078
rect 18696 4072 18748 4078
rect 18288 4020 18552 4026
rect 18236 4014 18552 4020
rect 18696 4014 18748 4020
rect 18788 4072 18840 4078
rect 18788 4014 18840 4020
rect 18972 4072 19024 4078
rect 18972 4014 19024 4020
rect 18248 4010 18552 4014
rect 18248 4004 18564 4010
rect 18248 3998 18512 4004
rect 17960 3528 18012 3534
rect 17960 3470 18012 3476
rect 18144 3528 18196 3534
rect 18144 3470 18196 3476
rect 17684 3120 17736 3126
rect 17684 3062 17736 3068
rect 17972 2514 18000 3470
rect 18248 3466 18276 3998
rect 18512 3946 18564 3952
rect 18328 3936 18380 3942
rect 18328 3878 18380 3884
rect 18340 3738 18368 3878
rect 18328 3732 18380 3738
rect 18328 3674 18380 3680
rect 18708 3670 18736 4014
rect 18696 3664 18748 3670
rect 18696 3606 18748 3612
rect 18800 3602 18828 4014
rect 18880 3732 18932 3738
rect 18880 3674 18932 3680
rect 18788 3596 18840 3602
rect 18788 3538 18840 3544
rect 18604 3528 18656 3534
rect 18604 3470 18656 3476
rect 18236 3460 18288 3466
rect 18236 3402 18288 3408
rect 18420 3188 18472 3194
rect 18420 3130 18472 3136
rect 18144 3052 18196 3058
rect 18144 2994 18196 3000
rect 18052 2848 18104 2854
rect 18052 2790 18104 2796
rect 18064 2582 18092 2790
rect 18156 2650 18184 2994
rect 18432 2922 18460 3130
rect 18420 2916 18472 2922
rect 18420 2858 18472 2864
rect 18144 2644 18196 2650
rect 18144 2586 18196 2592
rect 18052 2576 18104 2582
rect 18052 2518 18104 2524
rect 17960 2508 18012 2514
rect 17960 2450 18012 2456
rect 18064 2378 18092 2518
rect 18156 2514 18184 2586
rect 18616 2514 18644 3470
rect 18800 3194 18828 3538
rect 18788 3188 18840 3194
rect 18788 3130 18840 3136
rect 18800 2990 18828 3130
rect 18788 2984 18840 2990
rect 18788 2926 18840 2932
rect 18788 2848 18840 2854
rect 18788 2790 18840 2796
rect 18800 2514 18828 2790
rect 18144 2508 18196 2514
rect 18144 2450 18196 2456
rect 18604 2508 18656 2514
rect 18604 2450 18656 2456
rect 18788 2508 18840 2514
rect 18788 2450 18840 2456
rect 18892 2496 18920 3674
rect 18984 3602 19012 4014
rect 18972 3596 19024 3602
rect 18972 3538 19024 3544
rect 19156 3596 19208 3602
rect 19156 3538 19208 3544
rect 18984 3466 19012 3538
rect 18972 3460 19024 3466
rect 18972 3402 19024 3408
rect 18984 3058 19012 3402
rect 18972 3052 19024 3058
rect 18972 2994 19024 3000
rect 19168 2990 19196 3538
rect 19260 3534 19288 4150
rect 19996 3942 20024 5714
rect 20272 4826 20300 6802
rect 21284 6322 21312 7822
rect 21652 7546 21680 8366
rect 21744 7546 21772 8366
rect 21836 8362 21864 8978
rect 21824 8356 21876 8362
rect 21824 8298 21876 8304
rect 21928 8022 21956 9386
rect 22020 9110 22048 10542
rect 22100 9920 22152 9926
rect 22100 9862 22152 9868
rect 22112 9518 22140 9862
rect 22100 9512 22152 9518
rect 22100 9454 22152 9460
rect 22204 9382 22232 10950
rect 22296 10130 22324 11630
rect 22388 11234 22416 11630
rect 22480 11354 22508 12242
rect 22560 12096 22612 12102
rect 22560 12038 22612 12044
rect 22572 11694 22600 12038
rect 22560 11688 22612 11694
rect 22560 11630 22612 11636
rect 22848 11558 22876 12922
rect 23124 11830 23152 24686
rect 23388 24608 23440 24614
rect 23388 24550 23440 24556
rect 23400 24342 23428 24550
rect 23388 24336 23440 24342
rect 23388 24278 23440 24284
rect 23676 24274 23704 25094
rect 23768 24954 23796 25230
rect 24044 25158 24072 25978
rect 24320 25974 24348 26250
rect 24308 25968 24360 25974
rect 24308 25910 24360 25916
rect 24320 25498 24348 25910
rect 24308 25492 24360 25498
rect 24308 25434 24360 25440
rect 24320 25362 24348 25434
rect 24308 25356 24360 25362
rect 24308 25298 24360 25304
rect 24032 25152 24084 25158
rect 24032 25094 24084 25100
rect 23904 25052 24212 25061
rect 23904 25050 23910 25052
rect 23966 25050 23990 25052
rect 24046 25050 24070 25052
rect 24126 25050 24150 25052
rect 24206 25050 24212 25052
rect 23966 24998 23968 25050
rect 24148 24998 24150 25050
rect 23904 24996 23910 24998
rect 23966 24996 23990 24998
rect 24046 24996 24070 24998
rect 24126 24996 24150 24998
rect 24206 24996 24212 24998
rect 23904 24987 24212 24996
rect 23756 24948 23808 24954
rect 23756 24890 23808 24896
rect 24320 24834 24348 25298
rect 24504 24970 24532 29582
rect 24860 28688 24912 28694
rect 24860 28630 24912 28636
rect 24584 28076 24636 28082
rect 24584 28018 24636 28024
rect 24596 27334 24624 28018
rect 24584 27328 24636 27334
rect 24584 27270 24636 27276
rect 24676 26240 24728 26246
rect 24676 26182 24728 26188
rect 24688 26042 24716 26182
rect 24676 26036 24728 26042
rect 24676 25978 24728 25984
rect 24872 25945 24900 28630
rect 24858 25936 24914 25945
rect 24858 25871 24914 25880
rect 24676 25696 24728 25702
rect 24676 25638 24728 25644
rect 24688 25430 24716 25638
rect 24872 25430 24900 25871
rect 24676 25424 24728 25430
rect 24676 25366 24728 25372
rect 24860 25424 24912 25430
rect 24860 25366 24912 25372
rect 24504 24942 24624 24970
rect 24044 24806 24348 24834
rect 24492 24812 24544 24818
rect 24044 24682 24072 24806
rect 24492 24754 24544 24760
rect 24400 24744 24452 24750
rect 24400 24686 24452 24692
rect 23756 24676 23808 24682
rect 23756 24618 23808 24624
rect 24032 24676 24084 24682
rect 24032 24618 24084 24624
rect 23664 24268 23716 24274
rect 23664 24210 23716 24216
rect 23768 24206 23796 24618
rect 24308 24608 24360 24614
rect 24308 24550 24360 24556
rect 24320 24410 24348 24550
rect 24412 24410 24440 24686
rect 24308 24404 24360 24410
rect 24308 24346 24360 24352
rect 24400 24404 24452 24410
rect 24400 24346 24452 24352
rect 24504 24342 24532 24754
rect 24492 24336 24544 24342
rect 24492 24278 24544 24284
rect 23756 24200 23808 24206
rect 24504 24154 24532 24278
rect 23756 24142 23808 24148
rect 23296 24064 23348 24070
rect 23296 24006 23348 24012
rect 23308 23322 23336 24006
rect 23768 23866 23796 24142
rect 24412 24126 24532 24154
rect 23904 23964 24212 23973
rect 23904 23962 23910 23964
rect 23966 23962 23990 23964
rect 24046 23962 24070 23964
rect 24126 23962 24150 23964
rect 24206 23962 24212 23964
rect 23966 23910 23968 23962
rect 24148 23910 24150 23962
rect 23904 23908 23910 23910
rect 23966 23908 23990 23910
rect 24046 23908 24070 23910
rect 24126 23908 24150 23910
rect 24206 23908 24212 23910
rect 23904 23899 24212 23908
rect 24412 23866 24440 24126
rect 24492 24064 24544 24070
rect 24492 24006 24544 24012
rect 23756 23860 23808 23866
rect 23756 23802 23808 23808
rect 23848 23860 23900 23866
rect 23848 23802 23900 23808
rect 24400 23860 24452 23866
rect 24400 23802 24452 23808
rect 23296 23316 23348 23322
rect 23296 23258 23348 23264
rect 23860 23186 23888 23802
rect 23848 23180 23900 23186
rect 23848 23122 23900 23128
rect 24504 22982 24532 24006
rect 24596 23118 24624 24942
rect 24676 24744 24728 24750
rect 24676 24686 24728 24692
rect 24860 24744 24912 24750
rect 24860 24686 24912 24692
rect 24688 23322 24716 24686
rect 24768 24608 24820 24614
rect 24768 24550 24820 24556
rect 24780 23594 24808 24550
rect 24872 24342 24900 24686
rect 24860 24336 24912 24342
rect 24860 24278 24912 24284
rect 24768 23588 24820 23594
rect 24768 23530 24820 23536
rect 24676 23316 24728 23322
rect 24676 23258 24728 23264
rect 24584 23112 24636 23118
rect 24584 23054 24636 23060
rect 24492 22976 24544 22982
rect 24492 22918 24544 22924
rect 23904 22876 24212 22885
rect 23904 22874 23910 22876
rect 23966 22874 23990 22876
rect 24046 22874 24070 22876
rect 24126 22874 24150 22876
rect 24206 22874 24212 22876
rect 23966 22822 23968 22874
rect 24148 22822 24150 22874
rect 23904 22820 23910 22822
rect 23966 22820 23990 22822
rect 24046 22820 24070 22822
rect 24126 22820 24150 22822
rect 24206 22820 24212 22822
rect 23904 22811 24212 22820
rect 23204 22568 23256 22574
rect 23204 22510 23256 22516
rect 23480 22568 23532 22574
rect 23480 22510 23532 22516
rect 23216 22234 23244 22510
rect 23204 22228 23256 22234
rect 23204 22170 23256 22176
rect 23296 22160 23348 22166
rect 23296 22102 23348 22108
rect 23308 21350 23336 22102
rect 23492 21690 23520 22510
rect 23940 22432 23992 22438
rect 23940 22374 23992 22380
rect 24860 22432 24912 22438
rect 24860 22374 24912 22380
rect 23952 22098 23980 22374
rect 23940 22092 23992 22098
rect 23940 22034 23992 22040
rect 23904 21788 24212 21797
rect 23904 21786 23910 21788
rect 23966 21786 23990 21788
rect 24046 21786 24070 21788
rect 24126 21786 24150 21788
rect 24206 21786 24212 21788
rect 23966 21734 23968 21786
rect 24148 21734 24150 21786
rect 23904 21732 23910 21734
rect 23966 21732 23990 21734
rect 24046 21732 24070 21734
rect 24126 21732 24150 21734
rect 24206 21732 24212 21734
rect 23904 21723 24212 21732
rect 23480 21684 23532 21690
rect 23480 21626 23532 21632
rect 24872 21418 24900 22374
rect 24860 21412 24912 21418
rect 24860 21354 24912 21360
rect 23296 21344 23348 21350
rect 23296 21286 23348 21292
rect 23308 21078 23336 21286
rect 23296 21072 23348 21078
rect 23296 21014 23348 21020
rect 23480 21072 23532 21078
rect 23480 21014 23532 21020
rect 23204 21004 23256 21010
rect 23204 20946 23256 20952
rect 23216 20330 23244 20946
rect 23308 20874 23336 21014
rect 23296 20868 23348 20874
rect 23296 20810 23348 20816
rect 23204 20324 23256 20330
rect 23204 20266 23256 20272
rect 23204 20052 23256 20058
rect 23204 19994 23256 20000
rect 23216 19786 23244 19994
rect 23204 19780 23256 19786
rect 23204 19722 23256 19728
rect 23308 19310 23336 20810
rect 23492 20602 23520 21014
rect 23572 20800 23624 20806
rect 23572 20742 23624 20748
rect 23756 20800 23808 20806
rect 23756 20742 23808 20748
rect 23480 20596 23532 20602
rect 23480 20538 23532 20544
rect 23584 20262 23612 20742
rect 23768 20398 23796 20742
rect 23904 20700 24212 20709
rect 23904 20698 23910 20700
rect 23966 20698 23990 20700
rect 24046 20698 24070 20700
rect 24126 20698 24150 20700
rect 24206 20698 24212 20700
rect 23966 20646 23968 20698
rect 24148 20646 24150 20698
rect 23904 20644 23910 20646
rect 23966 20644 23990 20646
rect 24046 20644 24070 20646
rect 24126 20644 24150 20646
rect 24206 20644 24212 20646
rect 23904 20635 24212 20644
rect 23756 20392 23808 20398
rect 23756 20334 23808 20340
rect 23572 20256 23624 20262
rect 23572 20198 23624 20204
rect 23388 19984 23440 19990
rect 23388 19926 23440 19932
rect 23296 19304 23348 19310
rect 23296 19246 23348 19252
rect 23400 19242 23428 19926
rect 23584 19854 23612 20198
rect 23572 19848 23624 19854
rect 23572 19790 23624 19796
rect 23904 19612 24212 19621
rect 23904 19610 23910 19612
rect 23966 19610 23990 19612
rect 24046 19610 24070 19612
rect 24126 19610 24150 19612
rect 24206 19610 24212 19612
rect 23966 19558 23968 19610
rect 24148 19558 24150 19610
rect 23904 19556 23910 19558
rect 23966 19556 23990 19558
rect 24046 19556 24070 19558
rect 24126 19556 24150 19558
rect 24206 19556 24212 19558
rect 23904 19547 24212 19556
rect 23388 19236 23440 19242
rect 23388 19178 23440 19184
rect 23296 19168 23348 19174
rect 23296 19110 23348 19116
rect 24768 19168 24820 19174
rect 24768 19110 24820 19116
rect 23204 18828 23256 18834
rect 23204 18770 23256 18776
rect 23216 18290 23244 18770
rect 23308 18426 23336 19110
rect 23388 18896 23440 18902
rect 23388 18838 23440 18844
rect 23400 18426 23428 18838
rect 23904 18524 24212 18533
rect 23904 18522 23910 18524
rect 23966 18522 23990 18524
rect 24046 18522 24070 18524
rect 24126 18522 24150 18524
rect 24206 18522 24212 18524
rect 23966 18470 23968 18522
rect 24148 18470 24150 18522
rect 23904 18468 23910 18470
rect 23966 18468 23990 18470
rect 24046 18468 24070 18470
rect 24126 18468 24150 18470
rect 24206 18468 24212 18470
rect 23904 18459 24212 18468
rect 23296 18420 23348 18426
rect 23296 18362 23348 18368
rect 23388 18420 23440 18426
rect 23388 18362 23440 18368
rect 24400 18352 24452 18358
rect 24400 18294 24452 18300
rect 23204 18284 23256 18290
rect 23204 18226 23256 18232
rect 23216 17882 23244 18226
rect 24412 18222 24440 18294
rect 24780 18222 24808 19110
rect 24964 18698 24992 31600
rect 26436 30802 26464 31600
rect 27262 31036 27570 31045
rect 27262 31034 27268 31036
rect 27324 31034 27348 31036
rect 27404 31034 27428 31036
rect 27484 31034 27508 31036
rect 27564 31034 27570 31036
rect 27324 30982 27326 31034
rect 27506 30982 27508 31034
rect 27262 30980 27268 30982
rect 27324 30980 27348 30982
rect 27404 30980 27428 30982
rect 27484 30980 27508 30982
rect 27564 30980 27570 30982
rect 27262 30971 27570 30980
rect 26424 30796 26476 30802
rect 26424 30738 26476 30744
rect 25504 30184 25556 30190
rect 25504 30126 25556 30132
rect 25044 29776 25096 29782
rect 25044 29718 25096 29724
rect 25056 28558 25084 29718
rect 25412 29572 25464 29578
rect 25412 29514 25464 29520
rect 25424 28626 25452 29514
rect 25516 29102 25544 30126
rect 27262 29948 27570 29957
rect 27262 29946 27268 29948
rect 27324 29946 27348 29948
rect 27404 29946 27428 29948
rect 27484 29946 27508 29948
rect 27564 29946 27570 29948
rect 27324 29894 27326 29946
rect 27506 29894 27508 29946
rect 27262 29892 27268 29894
rect 27324 29892 27348 29894
rect 27404 29892 27428 29894
rect 27484 29892 27508 29894
rect 27564 29892 27570 29894
rect 27262 29883 27570 29892
rect 26976 29640 27028 29646
rect 26976 29582 27028 29588
rect 26988 29306 27016 29582
rect 26976 29300 27028 29306
rect 26976 29242 27028 29248
rect 25504 29096 25556 29102
rect 25504 29038 25556 29044
rect 26148 29096 26200 29102
rect 26148 29038 26200 29044
rect 25596 29028 25648 29034
rect 25596 28970 25648 28976
rect 25608 28762 25636 28970
rect 25596 28756 25648 28762
rect 25596 28698 25648 28704
rect 25412 28620 25464 28626
rect 25412 28562 25464 28568
rect 25044 28552 25096 28558
rect 25044 28494 25096 28500
rect 25056 27946 25084 28494
rect 25136 28008 25188 28014
rect 25136 27950 25188 27956
rect 25044 27940 25096 27946
rect 25044 27882 25096 27888
rect 25056 27606 25084 27882
rect 25044 27600 25096 27606
rect 25044 27542 25096 27548
rect 25056 27010 25084 27542
rect 25148 27402 25176 27950
rect 25320 27872 25372 27878
rect 25320 27814 25372 27820
rect 25332 27606 25360 27814
rect 25320 27600 25372 27606
rect 25320 27542 25372 27548
rect 26160 27538 26188 29038
rect 27262 28860 27570 28869
rect 27262 28858 27268 28860
rect 27324 28858 27348 28860
rect 27404 28858 27428 28860
rect 27484 28858 27508 28860
rect 27564 28858 27570 28860
rect 27324 28806 27326 28858
rect 27506 28806 27508 28858
rect 27262 28804 27268 28806
rect 27324 28804 27348 28806
rect 27404 28804 27428 28806
rect 27484 28804 27508 28806
rect 27564 28804 27570 28806
rect 27262 28795 27570 28804
rect 27262 27772 27570 27781
rect 27262 27770 27268 27772
rect 27324 27770 27348 27772
rect 27404 27770 27428 27772
rect 27484 27770 27508 27772
rect 27564 27770 27570 27772
rect 27324 27718 27326 27770
rect 27506 27718 27508 27770
rect 27262 27716 27268 27718
rect 27324 27716 27348 27718
rect 27404 27716 27428 27718
rect 27484 27716 27508 27718
rect 27564 27716 27570 27718
rect 27262 27707 27570 27716
rect 26148 27532 26200 27538
rect 26148 27474 26200 27480
rect 25136 27396 25188 27402
rect 25136 27338 25188 27344
rect 25056 26982 25176 27010
rect 25044 26920 25096 26926
rect 25044 26862 25096 26868
rect 25056 26518 25084 26862
rect 25148 26790 25176 26982
rect 26160 26926 26188 27474
rect 25320 26920 25372 26926
rect 25320 26862 25372 26868
rect 26148 26920 26200 26926
rect 26148 26862 26200 26868
rect 25136 26784 25188 26790
rect 25136 26726 25188 26732
rect 25044 26512 25096 26518
rect 25044 26454 25096 26460
rect 25044 26376 25096 26382
rect 25044 26318 25096 26324
rect 25056 26042 25084 26318
rect 25044 26036 25096 26042
rect 25044 25978 25096 25984
rect 25148 25838 25176 26726
rect 25332 25906 25360 26862
rect 25872 26852 25924 26858
rect 25872 26794 25924 26800
rect 25596 26784 25648 26790
rect 25596 26726 25648 26732
rect 25608 26450 25636 26726
rect 25884 26586 25912 26794
rect 27262 26684 27570 26693
rect 27262 26682 27268 26684
rect 27324 26682 27348 26684
rect 27404 26682 27428 26684
rect 27484 26682 27508 26684
rect 27564 26682 27570 26684
rect 27324 26630 27326 26682
rect 27506 26630 27508 26682
rect 27262 26628 27268 26630
rect 27324 26628 27348 26630
rect 27404 26628 27428 26630
rect 27484 26628 27508 26630
rect 27564 26628 27570 26630
rect 27262 26619 27570 26628
rect 25872 26580 25924 26586
rect 25872 26522 25924 26528
rect 25596 26444 25648 26450
rect 25596 26386 25648 26392
rect 25320 25900 25372 25906
rect 25320 25842 25372 25848
rect 25136 25832 25188 25838
rect 25136 25774 25188 25780
rect 25044 25764 25096 25770
rect 25044 25706 25096 25712
rect 25056 25362 25084 25706
rect 25148 25498 25176 25774
rect 25228 25764 25280 25770
rect 25228 25706 25280 25712
rect 25240 25498 25268 25706
rect 25136 25492 25188 25498
rect 25136 25434 25188 25440
rect 25228 25492 25280 25498
rect 25228 25434 25280 25440
rect 25044 25356 25096 25362
rect 25044 25298 25096 25304
rect 25148 24698 25176 25434
rect 25332 25276 25360 25842
rect 27262 25596 27570 25605
rect 27262 25594 27268 25596
rect 27324 25594 27348 25596
rect 27404 25594 27428 25596
rect 27484 25594 27508 25596
rect 27564 25594 27570 25596
rect 27324 25542 27326 25594
rect 27506 25542 27508 25594
rect 27262 25540 27268 25542
rect 27324 25540 27348 25542
rect 27404 25540 27428 25542
rect 27484 25540 27508 25542
rect 27564 25540 27570 25542
rect 27262 25531 27570 25540
rect 25872 25356 25924 25362
rect 25872 25298 25924 25304
rect 25412 25288 25464 25294
rect 25332 25248 25412 25276
rect 25412 25230 25464 25236
rect 25424 24750 25452 25230
rect 25320 24744 25372 24750
rect 25148 24670 25268 24698
rect 25320 24686 25372 24692
rect 25412 24744 25464 24750
rect 25412 24686 25464 24692
rect 25136 24608 25188 24614
rect 25136 24550 25188 24556
rect 25148 24274 25176 24550
rect 25240 24342 25268 24670
rect 25228 24336 25280 24342
rect 25228 24278 25280 24284
rect 25332 24274 25360 24686
rect 25136 24268 25188 24274
rect 25136 24210 25188 24216
rect 25320 24268 25372 24274
rect 25320 24210 25372 24216
rect 25148 23254 25176 24210
rect 25424 23662 25452 24686
rect 25780 24608 25832 24614
rect 25780 24550 25832 24556
rect 25596 24336 25648 24342
rect 25596 24278 25648 24284
rect 25608 23730 25636 24278
rect 25792 24070 25820 24550
rect 25780 24064 25832 24070
rect 25780 24006 25832 24012
rect 25596 23724 25648 23730
rect 25596 23666 25648 23672
rect 25412 23656 25464 23662
rect 25412 23598 25464 23604
rect 25136 23248 25188 23254
rect 25136 23190 25188 23196
rect 25044 23112 25096 23118
rect 25044 23054 25096 23060
rect 25056 22642 25084 23054
rect 25424 22642 25452 23598
rect 25608 23186 25636 23666
rect 25780 23520 25832 23526
rect 25780 23462 25832 23468
rect 25596 23180 25648 23186
rect 25596 23122 25648 23128
rect 25044 22636 25096 22642
rect 25044 22578 25096 22584
rect 25412 22636 25464 22642
rect 25412 22578 25464 22584
rect 25056 20942 25084 22578
rect 25424 22094 25452 22578
rect 25792 22574 25820 23462
rect 25780 22568 25832 22574
rect 25780 22510 25832 22516
rect 25424 22066 25636 22094
rect 25608 22030 25636 22066
rect 25596 22024 25648 22030
rect 25596 21966 25648 21972
rect 25608 21690 25636 21966
rect 25596 21684 25648 21690
rect 25596 21626 25648 21632
rect 25596 21412 25648 21418
rect 25596 21354 25648 21360
rect 25608 21146 25636 21354
rect 25596 21140 25648 21146
rect 25596 21082 25648 21088
rect 25044 20936 25096 20942
rect 25044 20878 25096 20884
rect 25884 20398 25912 25298
rect 26056 24676 26108 24682
rect 26056 24618 26108 24624
rect 26068 24410 26096 24618
rect 26884 24608 26936 24614
rect 26884 24550 26936 24556
rect 25964 24404 26016 24410
rect 25964 24346 26016 24352
rect 26056 24404 26108 24410
rect 26056 24346 26108 24352
rect 25976 23662 26004 24346
rect 26896 24274 26924 24550
rect 27262 24508 27570 24517
rect 27262 24506 27268 24508
rect 27324 24506 27348 24508
rect 27404 24506 27428 24508
rect 27484 24506 27508 24508
rect 27564 24506 27570 24508
rect 27324 24454 27326 24506
rect 27506 24454 27508 24506
rect 27262 24452 27268 24454
rect 27324 24452 27348 24454
rect 27404 24452 27428 24454
rect 27484 24452 27508 24454
rect 27564 24452 27570 24454
rect 27262 24443 27570 24452
rect 26884 24268 26936 24274
rect 26884 24210 26936 24216
rect 25964 23656 26016 23662
rect 25964 23598 26016 23604
rect 26700 23656 26752 23662
rect 26700 23598 26752 23604
rect 26712 23322 26740 23598
rect 27262 23420 27570 23429
rect 27262 23418 27268 23420
rect 27324 23418 27348 23420
rect 27404 23418 27428 23420
rect 27484 23418 27508 23420
rect 27564 23418 27570 23420
rect 27324 23366 27326 23418
rect 27506 23366 27508 23418
rect 27262 23364 27268 23366
rect 27324 23364 27348 23366
rect 27404 23364 27428 23366
rect 27484 23364 27508 23366
rect 27564 23364 27570 23366
rect 27262 23355 27570 23364
rect 26700 23316 26752 23322
rect 26700 23258 26752 23264
rect 26884 23112 26936 23118
rect 26884 23054 26936 23060
rect 26896 22778 26924 23054
rect 26884 22772 26936 22778
rect 26884 22714 26936 22720
rect 27262 22332 27570 22341
rect 27262 22330 27268 22332
rect 27324 22330 27348 22332
rect 27404 22330 27428 22332
rect 27484 22330 27508 22332
rect 27564 22330 27570 22332
rect 27324 22278 27326 22330
rect 27506 22278 27508 22330
rect 27262 22276 27268 22278
rect 27324 22276 27348 22278
rect 27404 22276 27428 22278
rect 27484 22276 27508 22278
rect 27564 22276 27570 22278
rect 27262 22267 27570 22276
rect 26976 21344 27028 21350
rect 26976 21286 27028 21292
rect 26988 21010 27016 21286
rect 27262 21244 27570 21253
rect 27262 21242 27268 21244
rect 27324 21242 27348 21244
rect 27404 21242 27428 21244
rect 27484 21242 27508 21244
rect 27564 21242 27570 21244
rect 27324 21190 27326 21242
rect 27506 21190 27508 21242
rect 27262 21188 27268 21190
rect 27324 21188 27348 21190
rect 27404 21188 27428 21190
rect 27484 21188 27508 21190
rect 27564 21188 27570 21190
rect 27262 21179 27570 21188
rect 26976 21004 27028 21010
rect 26976 20946 27028 20952
rect 25872 20392 25924 20398
rect 25872 20334 25924 20340
rect 27068 20324 27120 20330
rect 27068 20266 27120 20272
rect 27080 19854 27108 20266
rect 27262 20156 27570 20165
rect 27262 20154 27268 20156
rect 27324 20154 27348 20156
rect 27404 20154 27428 20156
rect 27484 20154 27508 20156
rect 27564 20154 27570 20156
rect 27324 20102 27326 20154
rect 27506 20102 27508 20154
rect 27262 20100 27268 20102
rect 27324 20100 27348 20102
rect 27404 20100 27428 20102
rect 27484 20100 27508 20102
rect 27564 20100 27570 20102
rect 27262 20091 27570 20100
rect 27068 19848 27120 19854
rect 27068 19790 27120 19796
rect 27080 19310 27108 19790
rect 25136 19304 25188 19310
rect 25136 19246 25188 19252
rect 27068 19304 27120 19310
rect 27068 19246 27120 19252
rect 24952 18692 25004 18698
rect 24952 18634 25004 18640
rect 24860 18352 24912 18358
rect 24860 18294 24912 18300
rect 24400 18216 24452 18222
rect 24400 18158 24452 18164
rect 24768 18216 24820 18222
rect 24768 18158 24820 18164
rect 23940 18080 23992 18086
rect 23940 18022 23992 18028
rect 23204 17876 23256 17882
rect 23204 17818 23256 17824
rect 23952 17746 23980 18022
rect 24412 17882 24440 18158
rect 24400 17876 24452 17882
rect 24400 17818 24452 17824
rect 24780 17814 24808 18158
rect 24872 17882 24900 18294
rect 25148 18154 25176 19246
rect 25780 19236 25832 19242
rect 25780 19178 25832 19184
rect 25792 18970 25820 19178
rect 25780 18964 25832 18970
rect 25780 18906 25832 18912
rect 25504 18828 25556 18834
rect 25504 18770 25556 18776
rect 25516 18426 25544 18770
rect 25504 18420 25556 18426
rect 25504 18362 25556 18368
rect 27080 18222 27108 19246
rect 27262 19068 27570 19077
rect 27262 19066 27268 19068
rect 27324 19066 27348 19068
rect 27404 19066 27428 19068
rect 27484 19066 27508 19068
rect 27564 19066 27570 19068
rect 27324 19014 27326 19066
rect 27506 19014 27508 19066
rect 27262 19012 27268 19014
rect 27324 19012 27348 19014
rect 27404 19012 27428 19014
rect 27484 19012 27508 19014
rect 27564 19012 27570 19014
rect 27262 19003 27570 19012
rect 27068 18216 27120 18222
rect 27068 18158 27120 18164
rect 25136 18148 25188 18154
rect 25136 18090 25188 18096
rect 25504 18148 25556 18154
rect 25504 18090 25556 18096
rect 26608 18148 26660 18154
rect 26608 18090 26660 18096
rect 24860 17876 24912 17882
rect 24860 17818 24912 17824
rect 24768 17808 24820 17814
rect 24768 17750 24820 17756
rect 23940 17740 23992 17746
rect 23940 17682 23992 17688
rect 24676 17740 24728 17746
rect 24676 17682 24728 17688
rect 24308 17536 24360 17542
rect 24308 17478 24360 17484
rect 23904 17436 24212 17445
rect 23904 17434 23910 17436
rect 23966 17434 23990 17436
rect 24046 17434 24070 17436
rect 24126 17434 24150 17436
rect 24206 17434 24212 17436
rect 23966 17382 23968 17434
rect 24148 17382 24150 17434
rect 23904 17380 23910 17382
rect 23966 17380 23990 17382
rect 24046 17380 24070 17382
rect 24126 17380 24150 17382
rect 24206 17380 24212 17382
rect 23904 17371 24212 17380
rect 23204 17128 23256 17134
rect 23204 17070 23256 17076
rect 24124 17128 24176 17134
rect 24124 17070 24176 17076
rect 23216 15706 23244 17070
rect 23572 17060 23624 17066
rect 23572 17002 23624 17008
rect 23584 16114 23612 17002
rect 24136 16794 24164 17070
rect 24124 16788 24176 16794
rect 24124 16730 24176 16736
rect 24320 16726 24348 17478
rect 24400 16992 24452 16998
rect 24400 16934 24452 16940
rect 24308 16720 24360 16726
rect 24308 16662 24360 16668
rect 23904 16348 24212 16357
rect 23904 16346 23910 16348
rect 23966 16346 23990 16348
rect 24046 16346 24070 16348
rect 24126 16346 24150 16348
rect 24206 16346 24212 16348
rect 23966 16294 23968 16346
rect 24148 16294 24150 16346
rect 23904 16292 23910 16294
rect 23966 16292 23990 16294
rect 24046 16292 24070 16294
rect 24126 16292 24150 16294
rect 24206 16292 24212 16294
rect 23904 16283 24212 16292
rect 23572 16108 23624 16114
rect 23572 16050 23624 16056
rect 24216 16040 24268 16046
rect 24320 16028 24348 16662
rect 24412 16658 24440 16934
rect 24688 16794 24716 17682
rect 24676 16788 24728 16794
rect 24676 16730 24728 16736
rect 24584 16720 24636 16726
rect 24584 16662 24636 16668
rect 24400 16652 24452 16658
rect 24400 16594 24452 16600
rect 24596 16046 24624 16662
rect 24872 16658 24900 17818
rect 24952 17604 25004 17610
rect 24952 17546 25004 17552
rect 25044 17604 25096 17610
rect 25044 17546 25096 17552
rect 24964 17066 24992 17546
rect 25056 17134 25084 17546
rect 25516 17542 25544 18090
rect 25780 18080 25832 18086
rect 25780 18022 25832 18028
rect 26148 18080 26200 18086
rect 26148 18022 26200 18028
rect 25792 17746 25820 18022
rect 26160 17746 26188 18022
rect 26620 17882 26648 18090
rect 26608 17876 26660 17882
rect 26608 17818 26660 17824
rect 27080 17814 27108 18158
rect 27262 17980 27570 17989
rect 27262 17978 27268 17980
rect 27324 17978 27348 17980
rect 27404 17978 27428 17980
rect 27484 17978 27508 17980
rect 27564 17978 27570 17980
rect 27324 17926 27326 17978
rect 27506 17926 27508 17978
rect 27262 17924 27268 17926
rect 27324 17924 27348 17926
rect 27404 17924 27428 17926
rect 27484 17924 27508 17926
rect 27564 17924 27570 17926
rect 27262 17915 27570 17924
rect 27068 17808 27120 17814
rect 27068 17750 27120 17756
rect 25688 17740 25740 17746
rect 25688 17682 25740 17688
rect 25780 17740 25832 17746
rect 25780 17682 25832 17688
rect 25964 17740 26016 17746
rect 25964 17682 26016 17688
rect 26148 17740 26200 17746
rect 26148 17682 26200 17688
rect 26424 17740 26476 17746
rect 26424 17682 26476 17688
rect 25700 17626 25728 17682
rect 25976 17626 26004 17682
rect 25700 17598 26004 17626
rect 26436 17542 26464 17682
rect 25504 17536 25556 17542
rect 25504 17478 25556 17484
rect 26424 17536 26476 17542
rect 26424 17478 26476 17484
rect 25044 17128 25096 17134
rect 25044 17070 25096 17076
rect 24952 17060 25004 17066
rect 24952 17002 25004 17008
rect 25320 16992 25372 16998
rect 25320 16934 25372 16940
rect 25332 16794 25360 16934
rect 25320 16788 25372 16794
rect 25320 16730 25372 16736
rect 24860 16652 24912 16658
rect 24860 16594 24912 16600
rect 25516 16454 25544 17478
rect 25688 17128 25740 17134
rect 25688 17070 25740 17076
rect 24860 16448 24912 16454
rect 24860 16390 24912 16396
rect 25504 16448 25556 16454
rect 25504 16390 25556 16396
rect 24872 16114 24900 16390
rect 24860 16108 24912 16114
rect 24860 16050 24912 16056
rect 25700 16046 25728 17070
rect 26056 17060 26108 17066
rect 26056 17002 26108 17008
rect 26068 16794 26096 17002
rect 27262 16892 27570 16901
rect 27262 16890 27268 16892
rect 27324 16890 27348 16892
rect 27404 16890 27428 16892
rect 27484 16890 27508 16892
rect 27564 16890 27570 16892
rect 27324 16838 27326 16890
rect 27506 16838 27508 16890
rect 27262 16836 27268 16838
rect 27324 16836 27348 16838
rect 27404 16836 27428 16838
rect 27484 16836 27508 16838
rect 27564 16836 27570 16838
rect 27262 16827 27570 16836
rect 26056 16788 26108 16794
rect 26056 16730 26108 16736
rect 24268 16000 24348 16028
rect 24492 16040 24544 16046
rect 24216 15982 24268 15988
rect 24492 15982 24544 15988
rect 24584 16040 24636 16046
rect 24584 15982 24636 15988
rect 24676 16040 24728 16046
rect 24676 15982 24728 15988
rect 25688 16040 25740 16046
rect 25688 15982 25740 15988
rect 24400 15904 24452 15910
rect 24400 15846 24452 15852
rect 23204 15700 23256 15706
rect 23204 15642 23256 15648
rect 24412 15570 24440 15846
rect 24504 15706 24532 15982
rect 24492 15700 24544 15706
rect 24492 15642 24544 15648
rect 24596 15570 24624 15982
rect 24688 15570 24716 15982
rect 24400 15564 24452 15570
rect 24400 15506 24452 15512
rect 24584 15564 24636 15570
rect 24584 15506 24636 15512
rect 24676 15564 24728 15570
rect 24676 15506 24728 15512
rect 24952 15564 25004 15570
rect 24952 15506 25004 15512
rect 23664 15496 23716 15502
rect 23664 15438 23716 15444
rect 23676 15162 23704 15438
rect 23904 15260 24212 15269
rect 23904 15258 23910 15260
rect 23966 15258 23990 15260
rect 24046 15258 24070 15260
rect 24126 15258 24150 15260
rect 24206 15258 24212 15260
rect 23966 15206 23968 15258
rect 24148 15206 24150 15258
rect 23904 15204 23910 15206
rect 23966 15204 23990 15206
rect 24046 15204 24070 15206
rect 24126 15204 24150 15206
rect 24206 15204 24212 15206
rect 23904 15195 24212 15204
rect 23664 15156 23716 15162
rect 23664 15098 23716 15104
rect 24964 14890 24992 15506
rect 25700 15026 25728 15982
rect 26240 15904 26292 15910
rect 26240 15846 26292 15852
rect 26252 15502 26280 15846
rect 27262 15804 27570 15813
rect 27262 15802 27268 15804
rect 27324 15802 27348 15804
rect 27404 15802 27428 15804
rect 27484 15802 27508 15804
rect 27564 15802 27570 15804
rect 27324 15750 27326 15802
rect 27506 15750 27508 15802
rect 27262 15748 27268 15750
rect 27324 15748 27348 15750
rect 27404 15748 27428 15750
rect 27484 15748 27508 15750
rect 27564 15748 27570 15750
rect 27262 15739 27570 15748
rect 26608 15564 26660 15570
rect 26608 15506 26660 15512
rect 26240 15496 26292 15502
rect 26240 15438 26292 15444
rect 26332 15156 26384 15162
rect 26332 15098 26384 15104
rect 25044 15020 25096 15026
rect 25044 14962 25096 14968
rect 25688 15020 25740 15026
rect 25688 14962 25740 14968
rect 23296 14884 23348 14890
rect 23296 14826 23348 14832
rect 24952 14884 25004 14890
rect 24952 14826 25004 14832
rect 23308 14482 23336 14826
rect 23388 14816 23440 14822
rect 23388 14758 23440 14764
rect 23296 14476 23348 14482
rect 23296 14418 23348 14424
rect 23400 14278 23428 14758
rect 25056 14618 25084 14962
rect 23756 14612 23808 14618
rect 23756 14554 23808 14560
rect 25044 14612 25096 14618
rect 25044 14554 25096 14560
rect 23480 14408 23532 14414
rect 23480 14350 23532 14356
rect 23388 14272 23440 14278
rect 23388 14214 23440 14220
rect 23204 14000 23256 14006
rect 23204 13942 23256 13948
rect 23216 12374 23244 13942
rect 23400 13870 23428 14214
rect 23388 13864 23440 13870
rect 23388 13806 23440 13812
rect 23296 13728 23348 13734
rect 23296 13670 23348 13676
rect 23308 13394 23336 13670
rect 23296 13388 23348 13394
rect 23296 13330 23348 13336
rect 23296 13252 23348 13258
rect 23296 13194 23348 13200
rect 23388 13252 23440 13258
rect 23388 13194 23440 13200
rect 23308 12850 23336 13194
rect 23296 12844 23348 12850
rect 23296 12786 23348 12792
rect 23308 12646 23336 12786
rect 23296 12640 23348 12646
rect 23296 12582 23348 12588
rect 23400 12442 23428 13194
rect 23492 12442 23520 14350
rect 23572 14340 23624 14346
rect 23768 14328 23796 14554
rect 24952 14408 25004 14414
rect 24952 14350 25004 14356
rect 23624 14300 23796 14328
rect 23572 14282 23624 14288
rect 23904 14172 24212 14181
rect 23904 14170 23910 14172
rect 23966 14170 23990 14172
rect 24046 14170 24070 14172
rect 24126 14170 24150 14172
rect 24206 14170 24212 14172
rect 23966 14118 23968 14170
rect 24148 14118 24150 14170
rect 23904 14116 23910 14118
rect 23966 14116 23990 14118
rect 24046 14116 24070 14118
rect 24126 14116 24150 14118
rect 24206 14116 24212 14118
rect 23904 14107 24212 14116
rect 23756 13864 23808 13870
rect 23756 13806 23808 13812
rect 24860 13864 24912 13870
rect 24860 13806 24912 13812
rect 23572 13728 23624 13734
rect 23572 13670 23624 13676
rect 23584 13462 23612 13670
rect 23572 13456 23624 13462
rect 23572 13398 23624 13404
rect 23768 12918 23796 13806
rect 24400 13796 24452 13802
rect 24400 13738 24452 13744
rect 24308 13184 24360 13190
rect 24308 13126 24360 13132
rect 23904 13084 24212 13093
rect 23904 13082 23910 13084
rect 23966 13082 23990 13084
rect 24046 13082 24070 13084
rect 24126 13082 24150 13084
rect 24206 13082 24212 13084
rect 23966 13030 23968 13082
rect 24148 13030 24150 13082
rect 23904 13028 23910 13030
rect 23966 13028 23990 13030
rect 24046 13028 24070 13030
rect 24126 13028 24150 13030
rect 24206 13028 24212 13030
rect 23904 13019 24212 13028
rect 23756 12912 23808 12918
rect 23756 12854 23808 12860
rect 23388 12436 23440 12442
rect 23388 12378 23440 12384
rect 23480 12436 23532 12442
rect 23480 12378 23532 12384
rect 24320 12374 24348 13126
rect 23204 12368 23256 12374
rect 23204 12310 23256 12316
rect 24308 12368 24360 12374
rect 24308 12310 24360 12316
rect 24412 12306 24440 13738
rect 24584 13728 24636 13734
rect 24584 13670 24636 13676
rect 24400 12300 24452 12306
rect 24400 12242 24452 12248
rect 24596 12170 24624 13670
rect 24872 13326 24900 13806
rect 24964 13462 24992 14350
rect 25056 13870 25084 14554
rect 25700 14550 25728 14962
rect 26344 14906 26372 15098
rect 26252 14878 26372 14906
rect 26424 14884 26476 14890
rect 25688 14544 25740 14550
rect 25688 14486 25740 14492
rect 25700 14346 25728 14486
rect 25688 14340 25740 14346
rect 25688 14282 25740 14288
rect 25044 13864 25096 13870
rect 25044 13806 25096 13812
rect 25596 13864 25648 13870
rect 25700 13852 25728 14282
rect 25780 14272 25832 14278
rect 25780 14214 25832 14220
rect 25792 13870 25820 14214
rect 25648 13824 25728 13852
rect 25780 13864 25832 13870
rect 25596 13806 25648 13812
rect 25780 13806 25832 13812
rect 25412 13524 25464 13530
rect 25412 13466 25464 13472
rect 24952 13456 25004 13462
rect 24952 13398 25004 13404
rect 24860 13320 24912 13326
rect 24860 13262 24912 13268
rect 24872 12986 24900 13262
rect 24952 13184 25004 13190
rect 24952 13126 25004 13132
rect 25044 13184 25096 13190
rect 25044 13126 25096 13132
rect 24860 12980 24912 12986
rect 24860 12922 24912 12928
rect 24964 12782 24992 13126
rect 24952 12776 25004 12782
rect 24952 12718 25004 12724
rect 25056 12442 25084 13126
rect 25228 12708 25280 12714
rect 25228 12650 25280 12656
rect 25240 12442 25268 12650
rect 25044 12436 25096 12442
rect 25044 12378 25096 12384
rect 25228 12436 25280 12442
rect 25228 12378 25280 12384
rect 25424 12374 25452 13466
rect 25608 12850 25636 13806
rect 25688 13456 25740 13462
rect 25688 13398 25740 13404
rect 25596 12844 25648 12850
rect 25596 12786 25648 12792
rect 25412 12368 25464 12374
rect 25412 12310 25464 12316
rect 24584 12164 24636 12170
rect 24584 12106 24636 12112
rect 23204 12096 23256 12102
rect 23204 12038 23256 12044
rect 23112 11824 23164 11830
rect 23112 11766 23164 11772
rect 23216 11626 23244 12038
rect 23904 11996 24212 12005
rect 23904 11994 23910 11996
rect 23966 11994 23990 11996
rect 24046 11994 24070 11996
rect 24126 11994 24150 11996
rect 24206 11994 24212 11996
rect 23966 11942 23968 11994
rect 24148 11942 24150 11994
rect 23904 11940 23910 11942
rect 23966 11940 23990 11942
rect 24046 11940 24070 11942
rect 24126 11940 24150 11942
rect 24206 11940 24212 11942
rect 23904 11931 24212 11940
rect 24768 11892 24820 11898
rect 24872 11886 25084 11914
rect 24872 11880 24900 11886
rect 24820 11852 24900 11880
rect 24768 11834 24820 11840
rect 24952 11688 25004 11694
rect 24780 11648 24952 11676
rect 23204 11620 23256 11626
rect 23204 11562 23256 11568
rect 23664 11620 23716 11626
rect 23664 11562 23716 11568
rect 22836 11552 22888 11558
rect 22836 11494 22888 11500
rect 23020 11552 23072 11558
rect 23020 11494 23072 11500
rect 22468 11348 22520 11354
rect 22468 11290 22520 11296
rect 23032 11286 23060 11494
rect 23216 11354 23244 11562
rect 23480 11552 23532 11558
rect 23532 11500 23612 11506
rect 23480 11494 23612 11500
rect 23492 11478 23612 11494
rect 23584 11354 23612 11478
rect 23204 11348 23256 11354
rect 23204 11290 23256 11296
rect 23480 11348 23532 11354
rect 23480 11290 23532 11296
rect 23572 11348 23624 11354
rect 23572 11290 23624 11296
rect 23020 11280 23072 11286
rect 22388 11206 22508 11234
rect 23020 11222 23072 11228
rect 22376 11144 22428 11150
rect 22376 11086 22428 11092
rect 22284 10124 22336 10130
rect 22284 10066 22336 10072
rect 22296 9722 22324 10066
rect 22284 9716 22336 9722
rect 22284 9658 22336 9664
rect 22388 9654 22416 11086
rect 22480 10674 22508 11206
rect 22468 10668 22520 10674
rect 22468 10610 22520 10616
rect 22836 10668 22888 10674
rect 22836 10610 22888 10616
rect 22848 10130 22876 10610
rect 23296 10600 23348 10606
rect 23296 10542 23348 10548
rect 23308 10266 23336 10542
rect 23492 10266 23520 11290
rect 23572 11076 23624 11082
rect 23572 11018 23624 11024
rect 23584 10606 23612 11018
rect 23676 11014 23704 11562
rect 24492 11552 24544 11558
rect 24492 11494 24544 11500
rect 24584 11552 24636 11558
rect 24584 11494 24636 11500
rect 23664 11008 23716 11014
rect 23664 10950 23716 10956
rect 23572 10600 23624 10606
rect 23572 10542 23624 10548
rect 23296 10260 23348 10266
rect 23296 10202 23348 10208
rect 23480 10260 23532 10266
rect 23480 10202 23532 10208
rect 22560 10124 22612 10130
rect 22560 10066 22612 10072
rect 22836 10124 22888 10130
rect 22836 10066 22888 10072
rect 23020 10124 23072 10130
rect 23020 10066 23072 10072
rect 23388 10124 23440 10130
rect 23388 10066 23440 10072
rect 22376 9648 22428 9654
rect 22376 9590 22428 9596
rect 22192 9376 22244 9382
rect 22192 9318 22244 9324
rect 22008 9104 22060 9110
rect 22008 9046 22060 9052
rect 22572 8634 22600 10066
rect 22652 9512 22704 9518
rect 22652 9454 22704 9460
rect 22664 9178 22692 9454
rect 22652 9172 22704 9178
rect 22652 9114 22704 9120
rect 22560 8628 22612 8634
rect 22560 8570 22612 8576
rect 23032 8090 23060 10066
rect 23400 8430 23428 10066
rect 23388 8424 23440 8430
rect 23388 8366 23440 8372
rect 23492 8378 23520 10202
rect 23584 9586 23612 10542
rect 23676 9722 23704 10950
rect 23904 10908 24212 10917
rect 23904 10906 23910 10908
rect 23966 10906 23990 10908
rect 24046 10906 24070 10908
rect 24126 10906 24150 10908
rect 24206 10906 24212 10908
rect 23966 10854 23968 10906
rect 24148 10854 24150 10906
rect 23904 10852 23910 10854
rect 23966 10852 23990 10854
rect 24046 10852 24070 10854
rect 24126 10852 24150 10854
rect 24206 10852 24212 10854
rect 23904 10843 24212 10852
rect 24308 10668 24360 10674
rect 24308 10610 24360 10616
rect 23848 10532 23900 10538
rect 23848 10474 23900 10480
rect 23860 9994 23888 10474
rect 24320 10130 24348 10610
rect 24504 10130 24532 11494
rect 24596 11354 24624 11494
rect 24584 11348 24636 11354
rect 24584 11290 24636 11296
rect 24596 10130 24624 11290
rect 24780 10674 24808 11648
rect 24952 11630 25004 11636
rect 24768 10668 24820 10674
rect 24768 10610 24820 10616
rect 24768 10532 24820 10538
rect 24768 10474 24820 10480
rect 24308 10124 24360 10130
rect 24308 10066 24360 10072
rect 24492 10124 24544 10130
rect 24492 10066 24544 10072
rect 24584 10124 24636 10130
rect 24584 10066 24636 10072
rect 23848 9988 23900 9994
rect 23848 9930 23900 9936
rect 23756 9920 23808 9926
rect 23756 9862 23808 9868
rect 23664 9716 23716 9722
rect 23664 9658 23716 9664
rect 23572 9580 23624 9586
rect 23572 9522 23624 9528
rect 23768 9042 23796 9862
rect 23904 9820 24212 9829
rect 23904 9818 23910 9820
rect 23966 9818 23990 9820
rect 24046 9818 24070 9820
rect 24126 9818 24150 9820
rect 24206 9818 24212 9820
rect 23966 9766 23968 9818
rect 24148 9766 24150 9818
rect 23904 9764 23910 9766
rect 23966 9764 23990 9766
rect 24046 9764 24070 9766
rect 24126 9764 24150 9766
rect 24206 9764 24212 9766
rect 23904 9755 24212 9764
rect 24320 9586 24348 10066
rect 24596 9994 24624 10066
rect 24584 9988 24636 9994
rect 24584 9930 24636 9936
rect 24124 9580 24176 9586
rect 24124 9522 24176 9528
rect 24308 9580 24360 9586
rect 24308 9522 24360 9528
rect 24136 9042 24164 9522
rect 24596 9178 24624 9930
rect 24676 9512 24728 9518
rect 24676 9454 24728 9460
rect 24688 9382 24716 9454
rect 24676 9376 24728 9382
rect 24676 9318 24728 9324
rect 24584 9172 24636 9178
rect 24584 9114 24636 9120
rect 23756 9036 23808 9042
rect 23756 8978 23808 8984
rect 24124 9036 24176 9042
rect 24124 8978 24176 8984
rect 24308 9036 24360 9042
rect 24308 8978 24360 8984
rect 24136 8838 24164 8978
rect 24124 8832 24176 8838
rect 24124 8774 24176 8780
rect 23904 8732 24212 8741
rect 23904 8730 23910 8732
rect 23966 8730 23990 8732
rect 24046 8730 24070 8732
rect 24126 8730 24150 8732
rect 24206 8730 24212 8732
rect 23966 8678 23968 8730
rect 24148 8678 24150 8730
rect 23904 8676 23910 8678
rect 23966 8676 23990 8678
rect 24046 8676 24070 8678
rect 24126 8676 24150 8678
rect 24206 8676 24212 8678
rect 23904 8667 24212 8676
rect 24032 8492 24084 8498
rect 24032 8434 24084 8440
rect 23492 8362 23612 8378
rect 23492 8356 23624 8362
rect 23492 8350 23572 8356
rect 23572 8298 23624 8304
rect 23480 8288 23532 8294
rect 23480 8230 23532 8236
rect 23020 8084 23072 8090
rect 23020 8026 23072 8032
rect 21916 8016 21968 8022
rect 21916 7958 21968 7964
rect 23492 7954 23520 8230
rect 23584 7954 23612 8298
rect 24044 8090 24072 8434
rect 24124 8356 24176 8362
rect 24124 8298 24176 8304
rect 24032 8084 24084 8090
rect 24032 8026 24084 8032
rect 24136 8022 24164 8298
rect 24320 8090 24348 8978
rect 24688 8974 24716 9318
rect 24676 8968 24728 8974
rect 24676 8910 24728 8916
rect 24400 8424 24452 8430
rect 24400 8366 24452 8372
rect 24308 8084 24360 8090
rect 24308 8026 24360 8032
rect 24124 8016 24176 8022
rect 24124 7958 24176 7964
rect 23388 7948 23440 7954
rect 23388 7890 23440 7896
rect 23480 7948 23532 7954
rect 23480 7890 23532 7896
rect 23572 7948 23624 7954
rect 23572 7890 23624 7896
rect 24032 7948 24084 7954
rect 24032 7890 24084 7896
rect 23400 7834 23428 7890
rect 24044 7834 24072 7890
rect 23400 7806 24072 7834
rect 21916 7744 21968 7750
rect 21916 7686 21968 7692
rect 21640 7540 21692 7546
rect 21640 7482 21692 7488
rect 21732 7540 21784 7546
rect 21732 7482 21784 7488
rect 21928 7410 21956 7686
rect 21916 7404 21968 7410
rect 21916 7346 21968 7352
rect 21928 7206 21956 7346
rect 22008 7336 22060 7342
rect 22008 7278 22060 7284
rect 23020 7336 23072 7342
rect 23020 7278 23072 7284
rect 23296 7336 23348 7342
rect 23296 7278 23348 7284
rect 23572 7336 23624 7342
rect 23572 7278 23624 7284
rect 21916 7200 21968 7206
rect 21916 7142 21968 7148
rect 22020 6934 22048 7278
rect 22560 7200 22612 7206
rect 22560 7142 22612 7148
rect 21456 6928 21508 6934
rect 21456 6870 21508 6876
rect 22008 6928 22060 6934
rect 22008 6870 22060 6876
rect 21272 6316 21324 6322
rect 21272 6258 21324 6264
rect 20546 6012 20854 6021
rect 20546 6010 20552 6012
rect 20608 6010 20632 6012
rect 20688 6010 20712 6012
rect 20768 6010 20792 6012
rect 20848 6010 20854 6012
rect 20608 5958 20610 6010
rect 20790 5958 20792 6010
rect 20546 5956 20552 5958
rect 20608 5956 20632 5958
rect 20688 5956 20712 5958
rect 20768 5956 20792 5958
rect 20848 5956 20854 5958
rect 20546 5947 20854 5956
rect 21468 5794 21496 6870
rect 22572 6730 22600 7142
rect 23032 6730 23060 7278
rect 23308 6866 23336 7278
rect 23584 6866 23612 7278
rect 23296 6860 23348 6866
rect 23296 6802 23348 6808
rect 23572 6860 23624 6866
rect 23572 6802 23624 6808
rect 22560 6724 22612 6730
rect 22560 6666 22612 6672
rect 23020 6724 23072 6730
rect 23020 6666 23072 6672
rect 21640 6656 21692 6662
rect 21640 6598 21692 6604
rect 21652 6254 21680 6598
rect 21640 6248 21692 6254
rect 21640 6190 21692 6196
rect 22928 6248 22980 6254
rect 22928 6190 22980 6196
rect 21824 5908 21876 5914
rect 21824 5850 21876 5856
rect 21548 5840 21600 5846
rect 21468 5788 21548 5794
rect 21468 5782 21600 5788
rect 21468 5766 21588 5782
rect 21732 5772 21784 5778
rect 21732 5714 21784 5720
rect 20904 5568 20956 5574
rect 20904 5510 20956 5516
rect 20916 5166 20944 5510
rect 21744 5370 21772 5714
rect 21836 5370 21864 5850
rect 21916 5840 21968 5846
rect 21916 5782 21968 5788
rect 21732 5364 21784 5370
rect 21732 5306 21784 5312
rect 21824 5364 21876 5370
rect 21824 5306 21876 5312
rect 21744 5166 21772 5306
rect 21928 5166 21956 5782
rect 22940 5778 22968 6190
rect 23032 5914 23060 6666
rect 23308 6458 23336 6802
rect 23296 6452 23348 6458
rect 23296 6394 23348 6400
rect 23584 6322 23612 6802
rect 23572 6316 23624 6322
rect 23572 6258 23624 6264
rect 23112 6112 23164 6118
rect 23112 6054 23164 6060
rect 23020 5908 23072 5914
rect 23020 5850 23072 5856
rect 23124 5778 23152 6054
rect 22928 5772 22980 5778
rect 22928 5714 22980 5720
rect 23112 5772 23164 5778
rect 23112 5714 23164 5720
rect 22560 5568 22612 5574
rect 22560 5510 22612 5516
rect 22572 5234 22600 5510
rect 22560 5228 22612 5234
rect 22560 5170 22612 5176
rect 20904 5160 20956 5166
rect 20904 5102 20956 5108
rect 21732 5160 21784 5166
rect 21732 5102 21784 5108
rect 21916 5160 21968 5166
rect 21916 5102 21968 5108
rect 22100 5160 22152 5166
rect 22100 5102 22152 5108
rect 20546 4924 20854 4933
rect 20546 4922 20552 4924
rect 20608 4922 20632 4924
rect 20688 4922 20712 4924
rect 20768 4922 20792 4924
rect 20848 4922 20854 4924
rect 20608 4870 20610 4922
rect 20790 4870 20792 4922
rect 20546 4868 20552 4870
rect 20608 4868 20632 4870
rect 20688 4868 20712 4870
rect 20768 4868 20792 4870
rect 20848 4868 20854 4870
rect 20546 4859 20854 4868
rect 20260 4820 20312 4826
rect 20260 4762 20312 4768
rect 20720 4684 20772 4690
rect 20720 4626 20772 4632
rect 21824 4684 21876 4690
rect 21824 4626 21876 4632
rect 20732 4146 20760 4626
rect 20720 4140 20772 4146
rect 20720 4082 20772 4088
rect 21364 4140 21416 4146
rect 21364 4082 21416 4088
rect 20168 4004 20220 4010
rect 20168 3946 20220 3952
rect 20444 4004 20496 4010
rect 20444 3946 20496 3952
rect 19984 3936 20036 3942
rect 19984 3878 20036 3884
rect 20180 3602 20208 3946
rect 20456 3738 20484 3946
rect 20546 3836 20854 3845
rect 20546 3834 20552 3836
rect 20608 3834 20632 3836
rect 20688 3834 20712 3836
rect 20768 3834 20792 3836
rect 20848 3834 20854 3836
rect 20608 3782 20610 3834
rect 20790 3782 20792 3834
rect 20546 3780 20552 3782
rect 20608 3780 20632 3782
rect 20688 3780 20712 3782
rect 20768 3780 20792 3782
rect 20848 3780 20854 3782
rect 20546 3771 20854 3780
rect 20444 3732 20496 3738
rect 20444 3674 20496 3680
rect 20168 3596 20220 3602
rect 20168 3538 20220 3544
rect 20720 3596 20772 3602
rect 20720 3538 20772 3544
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 20076 3188 20128 3194
rect 20076 3130 20128 3136
rect 19156 2984 19208 2990
rect 19156 2926 19208 2932
rect 20088 2650 20116 3130
rect 20180 2990 20208 3538
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 20640 3398 20668 3470
rect 20444 3392 20496 3398
rect 20444 3334 20496 3340
rect 20628 3392 20680 3398
rect 20628 3334 20680 3340
rect 20456 3058 20484 3334
rect 20732 3210 20760 3538
rect 21376 3398 21404 4082
rect 21836 3738 21864 4626
rect 22112 4622 22140 5102
rect 22940 4826 22968 5714
rect 23676 5302 23704 7806
rect 23904 7644 24212 7653
rect 23904 7642 23910 7644
rect 23966 7642 23990 7644
rect 24046 7642 24070 7644
rect 24126 7642 24150 7644
rect 24206 7642 24212 7644
rect 23966 7590 23968 7642
rect 24148 7590 24150 7642
rect 23904 7588 23910 7590
rect 23966 7588 23990 7590
rect 24046 7588 24070 7590
rect 24126 7588 24150 7590
rect 24206 7588 24212 7590
rect 23904 7579 24212 7588
rect 23756 7268 23808 7274
rect 23756 7210 23808 7216
rect 23768 6866 23796 7210
rect 23756 6860 23808 6866
rect 23756 6802 23808 6808
rect 23904 6556 24212 6565
rect 23904 6554 23910 6556
rect 23966 6554 23990 6556
rect 24046 6554 24070 6556
rect 24126 6554 24150 6556
rect 24206 6554 24212 6556
rect 23966 6502 23968 6554
rect 24148 6502 24150 6554
rect 23904 6500 23910 6502
rect 23966 6500 23990 6502
rect 24046 6500 24070 6502
rect 24126 6500 24150 6502
rect 24206 6500 24212 6502
rect 23904 6491 24212 6500
rect 24412 6458 24440 8366
rect 24780 8294 24808 10474
rect 24860 10464 24912 10470
rect 24860 10406 24912 10412
rect 24952 10464 25004 10470
rect 24952 10406 25004 10412
rect 24872 10198 24900 10406
rect 24860 10192 24912 10198
rect 24860 10134 24912 10140
rect 24964 9450 24992 10406
rect 25056 9518 25084 11886
rect 25608 11762 25636 12786
rect 25700 12306 25728 13398
rect 26252 13190 26280 14878
rect 26424 14826 26476 14832
rect 26240 13184 26292 13190
rect 26240 13126 26292 13132
rect 26252 12782 26280 13126
rect 26240 12776 26292 12782
rect 26240 12718 26292 12724
rect 26056 12640 26108 12646
rect 26056 12582 26108 12588
rect 26068 12306 26096 12582
rect 26436 12442 26464 14826
rect 26620 14482 26648 15506
rect 26976 15496 27028 15502
rect 26976 15438 27028 15444
rect 26792 15428 26844 15434
rect 26792 15370 26844 15376
rect 26700 15360 26752 15366
rect 26700 15302 26752 15308
rect 26608 14476 26660 14482
rect 26608 14418 26660 14424
rect 26620 13530 26648 14418
rect 26608 13524 26660 13530
rect 26608 13466 26660 13472
rect 26608 13388 26660 13394
rect 26608 13330 26660 13336
rect 26424 12436 26476 12442
rect 26424 12378 26476 12384
rect 25688 12300 25740 12306
rect 25688 12242 25740 12248
rect 26056 12300 26108 12306
rect 26056 12242 26108 12248
rect 25700 12170 25728 12242
rect 26148 12232 26200 12238
rect 26148 12174 26200 12180
rect 25688 12164 25740 12170
rect 25688 12106 25740 12112
rect 25700 11898 25728 12106
rect 25688 11892 25740 11898
rect 25688 11834 25740 11840
rect 25596 11756 25648 11762
rect 25596 11698 25648 11704
rect 25136 11688 25188 11694
rect 25136 11630 25188 11636
rect 25148 10198 25176 11630
rect 26160 11354 26188 12174
rect 26620 11898 26648 13330
rect 26712 12306 26740 15302
rect 26804 12434 26832 15370
rect 26988 15162 27016 15438
rect 26976 15156 27028 15162
rect 26976 15098 27028 15104
rect 26884 14816 26936 14822
rect 26884 14758 26936 14764
rect 26896 14482 26924 14758
rect 27262 14716 27570 14725
rect 27262 14714 27268 14716
rect 27324 14714 27348 14716
rect 27404 14714 27428 14716
rect 27484 14714 27508 14716
rect 27564 14714 27570 14716
rect 27324 14662 27326 14714
rect 27506 14662 27508 14714
rect 27262 14660 27268 14662
rect 27324 14660 27348 14662
rect 27404 14660 27428 14662
rect 27484 14660 27508 14662
rect 27564 14660 27570 14662
rect 27262 14651 27570 14660
rect 26884 14476 26936 14482
rect 26884 14418 26936 14424
rect 26976 14476 27028 14482
rect 26976 14418 27028 14424
rect 26884 13728 26936 13734
rect 26884 13670 26936 13676
rect 26896 13394 26924 13670
rect 26884 13388 26936 13394
rect 26884 13330 26936 13336
rect 26804 12406 26924 12434
rect 26896 12306 26924 12406
rect 26988 12374 27016 14418
rect 27262 13628 27570 13637
rect 27262 13626 27268 13628
rect 27324 13626 27348 13628
rect 27404 13626 27428 13628
rect 27484 13626 27508 13628
rect 27564 13626 27570 13628
rect 27324 13574 27326 13626
rect 27506 13574 27508 13626
rect 27262 13572 27268 13574
rect 27324 13572 27348 13574
rect 27404 13572 27428 13574
rect 27484 13572 27508 13574
rect 27564 13572 27570 13574
rect 27262 13563 27570 13572
rect 27068 13320 27120 13326
rect 27068 13262 27120 13268
rect 27080 12986 27108 13262
rect 27068 12980 27120 12986
rect 27068 12922 27120 12928
rect 26976 12368 27028 12374
rect 26976 12310 27028 12316
rect 26700 12300 26752 12306
rect 26700 12242 26752 12248
rect 26884 12300 26936 12306
rect 26884 12242 26936 12248
rect 26608 11892 26660 11898
rect 26608 11834 26660 11840
rect 26976 11892 27028 11898
rect 26976 11834 27028 11840
rect 26424 11688 26476 11694
rect 26424 11630 26476 11636
rect 26148 11348 26200 11354
rect 26148 11290 26200 11296
rect 25596 11144 25648 11150
rect 25596 11086 25648 11092
rect 26056 11144 26108 11150
rect 26056 11086 26108 11092
rect 25412 11008 25464 11014
rect 25412 10950 25464 10956
rect 25424 10810 25452 10950
rect 25412 10804 25464 10810
rect 25412 10746 25464 10752
rect 25608 10606 25636 11086
rect 25320 10600 25372 10606
rect 25320 10542 25372 10548
rect 25596 10600 25648 10606
rect 25596 10542 25648 10548
rect 25136 10192 25188 10198
rect 25136 10134 25188 10140
rect 25136 10056 25188 10062
rect 25136 9998 25188 10004
rect 25148 9722 25176 9998
rect 25136 9716 25188 9722
rect 25136 9658 25188 9664
rect 25044 9512 25096 9518
rect 25044 9454 25096 9460
rect 25136 9512 25188 9518
rect 25136 9454 25188 9460
rect 25228 9512 25280 9518
rect 25228 9454 25280 9460
rect 24952 9444 25004 9450
rect 24952 9386 25004 9392
rect 25148 9382 25176 9454
rect 25136 9376 25188 9382
rect 25136 9318 25188 9324
rect 25148 9178 25176 9318
rect 25136 9172 25188 9178
rect 25136 9114 25188 9120
rect 25240 9110 25268 9454
rect 24860 9104 24912 9110
rect 24860 9046 24912 9052
rect 25228 9104 25280 9110
rect 25228 9046 25280 9052
rect 24768 8288 24820 8294
rect 24768 8230 24820 8236
rect 24492 8016 24544 8022
rect 24492 7958 24544 7964
rect 24504 7002 24532 7958
rect 24780 7954 24808 8230
rect 24872 8090 24900 9046
rect 24952 8832 25004 8838
rect 24952 8774 25004 8780
rect 24964 8430 24992 8774
rect 24952 8424 25004 8430
rect 24952 8366 25004 8372
rect 25044 8356 25096 8362
rect 25044 8298 25096 8304
rect 24860 8084 24912 8090
rect 24860 8026 24912 8032
rect 24768 7948 24820 7954
rect 24768 7890 24820 7896
rect 24584 7336 24636 7342
rect 24584 7278 24636 7284
rect 24492 6996 24544 7002
rect 24492 6938 24544 6944
rect 24596 6458 24624 7278
rect 25056 7274 25084 8298
rect 25332 8294 25360 10542
rect 25504 10464 25556 10470
rect 25504 10406 25556 10412
rect 25516 9722 25544 10406
rect 25504 9716 25556 9722
rect 25504 9658 25556 9664
rect 25608 9518 25636 10542
rect 26068 9994 26096 11086
rect 26160 10266 26188 11290
rect 26436 10266 26464 11630
rect 26884 10804 26936 10810
rect 26884 10746 26936 10752
rect 26148 10260 26200 10266
rect 26148 10202 26200 10208
rect 26424 10260 26476 10266
rect 26424 10202 26476 10208
rect 26056 9988 26108 9994
rect 26056 9930 26108 9936
rect 25596 9512 25648 9518
rect 25596 9454 25648 9460
rect 26240 9512 26292 9518
rect 26240 9454 26292 9460
rect 25608 8430 25636 9454
rect 25780 9444 25832 9450
rect 25780 9386 25832 9392
rect 25792 9178 25820 9386
rect 26056 9376 26108 9382
rect 26056 9318 26108 9324
rect 25780 9172 25832 9178
rect 25780 9114 25832 9120
rect 25964 9172 26016 9178
rect 25964 9114 26016 9120
rect 25596 8424 25648 8430
rect 25596 8366 25648 8372
rect 25688 8356 25740 8362
rect 25688 8298 25740 8304
rect 25320 8288 25372 8294
rect 25320 8230 25372 8236
rect 25332 8022 25360 8230
rect 25700 8090 25728 8298
rect 25688 8084 25740 8090
rect 25688 8026 25740 8032
rect 25320 8016 25372 8022
rect 25320 7958 25372 7964
rect 25872 7948 25924 7954
rect 25872 7890 25924 7896
rect 25884 7546 25912 7890
rect 25872 7540 25924 7546
rect 25872 7482 25924 7488
rect 25044 7268 25096 7274
rect 25044 7210 25096 7216
rect 24768 6860 24820 6866
rect 24768 6802 24820 6808
rect 24780 6662 24808 6802
rect 24768 6656 24820 6662
rect 24768 6598 24820 6604
rect 24400 6452 24452 6458
rect 24400 6394 24452 6400
rect 24584 6452 24636 6458
rect 24584 6394 24636 6400
rect 24308 5636 24360 5642
rect 24308 5578 24360 5584
rect 23904 5468 24212 5477
rect 23904 5466 23910 5468
rect 23966 5466 23990 5468
rect 24046 5466 24070 5468
rect 24126 5466 24150 5468
rect 24206 5466 24212 5468
rect 23966 5414 23968 5466
rect 24148 5414 24150 5466
rect 23904 5412 23910 5414
rect 23966 5412 23990 5414
rect 24046 5412 24070 5414
rect 24126 5412 24150 5414
rect 24206 5412 24212 5414
rect 23904 5403 24212 5412
rect 24320 5370 24348 5578
rect 24308 5364 24360 5370
rect 24308 5306 24360 5312
rect 23664 5296 23716 5302
rect 23664 5238 23716 5244
rect 23204 5160 23256 5166
rect 23204 5102 23256 5108
rect 24412 5114 24440 6394
rect 24676 5840 24728 5846
rect 24676 5782 24728 5788
rect 24584 5568 24636 5574
rect 24584 5510 24636 5516
rect 24596 5166 24624 5510
rect 24688 5234 24716 5782
rect 24780 5574 24808 6598
rect 24768 5568 24820 5574
rect 24768 5510 24820 5516
rect 24676 5228 24728 5234
rect 24676 5170 24728 5176
rect 24584 5160 24636 5166
rect 23216 4826 23244 5102
rect 24412 5086 24532 5114
rect 24584 5102 24636 5108
rect 24400 5024 24452 5030
rect 24400 4966 24452 4972
rect 24412 4826 24440 4966
rect 22928 4820 22980 4826
rect 22928 4762 22980 4768
rect 23204 4820 23256 4826
rect 23204 4762 23256 4768
rect 24400 4820 24452 4826
rect 24400 4762 24452 4768
rect 23388 4684 23440 4690
rect 23388 4626 23440 4632
rect 22100 4616 22152 4622
rect 22100 4558 22152 4564
rect 23400 4282 23428 4626
rect 24504 4486 24532 5086
rect 24596 4826 24624 5102
rect 24584 4820 24636 4826
rect 24584 4762 24636 4768
rect 24780 4690 24808 5510
rect 25056 5234 25084 7210
rect 25320 6928 25372 6934
rect 25320 6870 25372 6876
rect 25136 6860 25188 6866
rect 25136 6802 25188 6808
rect 25228 6860 25280 6866
rect 25228 6802 25280 6808
rect 25148 6662 25176 6802
rect 25240 6730 25268 6802
rect 25228 6724 25280 6730
rect 25228 6666 25280 6672
rect 25136 6656 25188 6662
rect 25136 6598 25188 6604
rect 25136 6248 25188 6254
rect 25136 6190 25188 6196
rect 25044 5228 25096 5234
rect 25044 5170 25096 5176
rect 24768 4684 24820 4690
rect 24768 4626 24820 4632
rect 24492 4480 24544 4486
rect 24492 4422 24544 4428
rect 23904 4380 24212 4389
rect 23904 4378 23910 4380
rect 23966 4378 23990 4380
rect 24046 4378 24070 4380
rect 24126 4378 24150 4380
rect 24206 4378 24212 4380
rect 23966 4326 23968 4378
rect 24148 4326 24150 4378
rect 23904 4324 23910 4326
rect 23966 4324 23990 4326
rect 24046 4324 24070 4326
rect 24126 4324 24150 4326
rect 24206 4324 24212 4326
rect 23904 4315 24212 4324
rect 22376 4276 22428 4282
rect 22376 4218 22428 4224
rect 23388 4276 23440 4282
rect 23388 4218 23440 4224
rect 22192 4072 22244 4078
rect 22192 4014 22244 4020
rect 21824 3732 21876 3738
rect 21824 3674 21876 3680
rect 21640 3460 21692 3466
rect 21640 3402 21692 3408
rect 21364 3392 21416 3398
rect 21364 3334 21416 3340
rect 20640 3182 20760 3210
rect 20640 3126 20668 3182
rect 20628 3120 20680 3126
rect 20628 3062 20680 3068
rect 20444 3052 20496 3058
rect 20444 2994 20496 3000
rect 20168 2984 20220 2990
rect 20168 2926 20220 2932
rect 20352 2848 20404 2854
rect 20352 2790 20404 2796
rect 20076 2644 20128 2650
rect 20076 2586 20128 2592
rect 20088 2514 20116 2586
rect 20364 2514 20392 2790
rect 20456 2582 20484 2994
rect 21652 2990 21680 3402
rect 22100 3392 22152 3398
rect 22100 3334 22152 3340
rect 22112 3194 22140 3334
rect 21824 3188 21876 3194
rect 21824 3130 21876 3136
rect 21916 3188 21968 3194
rect 21916 3130 21968 3136
rect 22100 3188 22152 3194
rect 22100 3130 22152 3136
rect 21836 2990 21864 3130
rect 21640 2984 21692 2990
rect 21638 2952 21640 2961
rect 21824 2984 21876 2990
rect 21692 2952 21694 2961
rect 21824 2926 21876 2932
rect 21928 2922 21956 3130
rect 22008 3052 22060 3058
rect 22008 2994 22060 3000
rect 21638 2887 21694 2896
rect 21916 2916 21968 2922
rect 21916 2858 21968 2864
rect 20546 2748 20854 2757
rect 20546 2746 20552 2748
rect 20608 2746 20632 2748
rect 20688 2746 20712 2748
rect 20768 2746 20792 2748
rect 20848 2746 20854 2748
rect 20608 2694 20610 2746
rect 20790 2694 20792 2746
rect 20546 2692 20552 2694
rect 20608 2692 20632 2694
rect 20688 2692 20712 2694
rect 20768 2692 20792 2694
rect 20848 2692 20854 2694
rect 20546 2683 20854 2692
rect 20444 2576 20496 2582
rect 20444 2518 20496 2524
rect 22020 2514 22048 2994
rect 18972 2508 19024 2514
rect 18892 2468 18972 2496
rect 18052 2372 18104 2378
rect 18052 2314 18104 2320
rect 17684 2304 17736 2310
rect 17684 2246 17736 2252
rect 18512 2304 18564 2310
rect 18512 2246 18564 2252
rect 17188 2204 17496 2213
rect 17188 2202 17194 2204
rect 17250 2202 17274 2204
rect 17330 2202 17354 2204
rect 17410 2202 17434 2204
rect 17490 2202 17496 2204
rect 17250 2150 17252 2202
rect 17432 2150 17434 2202
rect 17188 2148 17194 2150
rect 17250 2148 17274 2150
rect 17330 2148 17354 2150
rect 17410 2148 17434 2150
rect 17490 2148 17496 2150
rect 17188 2139 17496 2148
rect 17316 1896 17368 1902
rect 17316 1838 17368 1844
rect 17592 1896 17644 1902
rect 17592 1838 17644 1844
rect 17040 1488 17092 1494
rect 17040 1430 17092 1436
rect 17328 1426 17356 1838
rect 16764 1420 16816 1426
rect 16684 1380 16764 1408
rect 16396 808 16448 814
rect 16396 750 16448 756
rect 16580 808 16632 814
rect 16580 750 16632 756
rect 16684 400 16712 1380
rect 16764 1362 16816 1368
rect 17316 1420 17368 1426
rect 17316 1362 17368 1368
rect 17188 1116 17496 1125
rect 17188 1114 17194 1116
rect 17250 1114 17274 1116
rect 17330 1114 17354 1116
rect 17410 1114 17434 1116
rect 17490 1114 17496 1116
rect 17250 1062 17252 1114
rect 17432 1062 17434 1114
rect 17188 1060 17194 1062
rect 17250 1060 17274 1062
rect 17330 1060 17354 1062
rect 17410 1060 17434 1062
rect 17490 1060 17496 1062
rect 17188 1051 17496 1060
rect 17604 814 17632 1838
rect 17696 814 17724 2246
rect 17868 1896 17920 1902
rect 17868 1838 17920 1844
rect 17776 1556 17828 1562
rect 17776 1498 17828 1504
rect 17224 808 17276 814
rect 17224 750 17276 756
rect 17592 808 17644 814
rect 17592 750 17644 756
rect 17684 808 17736 814
rect 17684 750 17736 756
rect 17236 400 17264 750
rect 17788 400 17816 1498
rect 17880 1494 17908 1838
rect 18524 1494 18552 2246
rect 18892 2106 18920 2468
rect 18972 2450 19024 2456
rect 20076 2508 20128 2514
rect 20076 2450 20128 2456
rect 20352 2508 20404 2514
rect 20720 2508 20772 2514
rect 20352 2450 20404 2456
rect 20640 2468 20720 2496
rect 18972 2304 19024 2310
rect 18972 2246 19024 2252
rect 19064 2304 19116 2310
rect 19064 2246 19116 2252
rect 19800 2304 19852 2310
rect 19800 2246 19852 2252
rect 20260 2304 20312 2310
rect 20260 2246 20312 2252
rect 18880 2100 18932 2106
rect 18880 2042 18932 2048
rect 18696 1896 18748 1902
rect 18696 1838 18748 1844
rect 17868 1488 17920 1494
rect 17868 1430 17920 1436
rect 18512 1488 18564 1494
rect 18512 1430 18564 1436
rect 18708 882 18736 1838
rect 18880 1420 18932 1426
rect 18880 1362 18932 1368
rect 18696 876 18748 882
rect 18696 818 18748 824
rect 18328 808 18380 814
rect 18328 750 18380 756
rect 18340 400 18368 750
rect 18892 400 18920 1362
rect 18984 814 19012 2246
rect 19076 1494 19104 2246
rect 19812 1902 19840 2246
rect 19248 1896 19300 1902
rect 19248 1838 19300 1844
rect 19800 1896 19852 1902
rect 19800 1838 19852 1844
rect 19064 1488 19116 1494
rect 19064 1430 19116 1436
rect 19260 1358 19288 1838
rect 20076 1420 20128 1426
rect 20076 1362 20128 1368
rect 19248 1352 19300 1358
rect 19248 1294 19300 1300
rect 19984 1216 20036 1222
rect 19984 1158 20036 1164
rect 19996 882 20024 1158
rect 19984 876 20036 882
rect 19984 818 20036 824
rect 18972 808 19024 814
rect 18972 750 19024 756
rect 19432 808 19484 814
rect 20088 762 20116 1362
rect 20272 814 20300 2246
rect 20640 2038 20668 2468
rect 20720 2450 20772 2456
rect 22008 2508 22060 2514
rect 22008 2450 22060 2456
rect 22204 2378 22232 4014
rect 22388 3942 22416 4218
rect 22928 4072 22980 4078
rect 22928 4014 22980 4020
rect 23204 4072 23256 4078
rect 23204 4014 23256 4020
rect 23756 4072 23808 4078
rect 23756 4014 23808 4020
rect 22376 3936 22428 3942
rect 22376 3878 22428 3884
rect 22560 3596 22612 3602
rect 22560 3538 22612 3544
rect 22572 3194 22600 3538
rect 22836 3528 22888 3534
rect 22836 3470 22888 3476
rect 22560 3188 22612 3194
rect 22560 3130 22612 3136
rect 22284 2508 22336 2514
rect 22284 2450 22336 2456
rect 22192 2372 22244 2378
rect 22192 2314 22244 2320
rect 21548 2304 21600 2310
rect 21548 2246 21600 2252
rect 20628 2032 20680 2038
rect 20628 1974 20680 1980
rect 20444 1896 20496 1902
rect 20444 1838 20496 1844
rect 21364 1896 21416 1902
rect 21364 1838 21416 1844
rect 19432 750 19484 756
rect 19444 400 19472 750
rect 19996 734 20116 762
rect 20260 808 20312 814
rect 20260 750 20312 756
rect 19996 400 20024 734
rect 20456 474 20484 1838
rect 20546 1660 20854 1669
rect 20546 1658 20552 1660
rect 20608 1658 20632 1660
rect 20688 1658 20712 1660
rect 20768 1658 20792 1660
rect 20848 1658 20854 1660
rect 20608 1606 20610 1658
rect 20790 1606 20792 1658
rect 20546 1604 20552 1606
rect 20608 1604 20632 1606
rect 20688 1604 20712 1606
rect 20768 1604 20792 1606
rect 20848 1604 20854 1606
rect 20546 1595 20854 1604
rect 21272 1352 21324 1358
rect 21272 1294 21324 1300
rect 21284 1018 21312 1294
rect 21376 1018 21404 1838
rect 21560 1426 21588 2246
rect 22204 1986 22232 2314
rect 22296 2106 22324 2450
rect 22284 2100 22336 2106
rect 22284 2042 22336 2048
rect 22376 2032 22428 2038
rect 22204 1958 22324 1986
rect 22376 1974 22428 1980
rect 22192 1896 22244 1902
rect 22192 1838 22244 1844
rect 21548 1420 21600 1426
rect 21548 1362 21600 1368
rect 21640 1420 21692 1426
rect 21640 1362 21692 1368
rect 21272 1012 21324 1018
rect 21272 954 21324 960
rect 21364 1012 21416 1018
rect 21364 954 21416 960
rect 21088 808 21140 814
rect 21088 750 21140 756
rect 20546 572 20854 581
rect 20546 570 20552 572
rect 20608 570 20632 572
rect 20688 570 20712 572
rect 20768 570 20792 572
rect 20848 570 20854 572
rect 20608 518 20610 570
rect 20790 518 20792 570
rect 20546 516 20552 518
rect 20608 516 20632 518
rect 20688 516 20712 518
rect 20768 516 20792 518
rect 20848 516 20854 518
rect 20546 507 20854 516
rect 20444 468 20496 474
rect 20628 468 20680 474
rect 20444 410 20496 416
rect 20548 428 20628 456
rect 20548 400 20576 428
rect 20628 410 20680 416
rect 21100 400 21128 750
rect 21652 400 21680 1362
rect 22204 400 22232 1838
rect 22296 1494 22324 1958
rect 22284 1488 22336 1494
rect 22284 1430 22336 1436
rect 22388 814 22416 1974
rect 22468 1896 22520 1902
rect 22468 1838 22520 1844
rect 22480 1426 22508 1838
rect 22468 1420 22520 1426
rect 22468 1362 22520 1368
rect 22572 814 22600 3130
rect 22848 3058 22876 3470
rect 22940 3398 22968 4014
rect 23112 3664 23164 3670
rect 23112 3606 23164 3612
rect 22928 3392 22980 3398
rect 22928 3334 22980 3340
rect 22940 3194 22968 3334
rect 22928 3188 22980 3194
rect 22928 3130 22980 3136
rect 22836 3052 22888 3058
rect 22836 2994 22888 3000
rect 22848 2774 22876 2994
rect 22940 2938 22968 3130
rect 23124 2961 23152 3606
rect 23216 3602 23244 4014
rect 23388 3936 23440 3942
rect 23388 3878 23440 3884
rect 23204 3596 23256 3602
rect 23204 3538 23256 3544
rect 23400 3194 23428 3878
rect 23664 3392 23716 3398
rect 23664 3334 23716 3340
rect 23388 3188 23440 3194
rect 23388 3130 23440 3136
rect 23676 2990 23704 3334
rect 23768 3176 23796 4014
rect 25148 3738 25176 6190
rect 25240 5914 25268 6666
rect 25332 6458 25360 6870
rect 25976 6866 26004 9114
rect 26068 8906 26096 9318
rect 26252 9042 26280 9454
rect 26896 9042 26924 10746
rect 26988 10130 27016 11834
rect 27080 11218 27108 12922
rect 27262 12540 27570 12549
rect 27262 12538 27268 12540
rect 27324 12538 27348 12540
rect 27404 12538 27428 12540
rect 27484 12538 27508 12540
rect 27564 12538 27570 12540
rect 27324 12486 27326 12538
rect 27506 12486 27508 12538
rect 27262 12484 27268 12486
rect 27324 12484 27348 12486
rect 27404 12484 27428 12486
rect 27484 12484 27508 12486
rect 27564 12484 27570 12486
rect 27262 12475 27570 12484
rect 27262 11452 27570 11461
rect 27262 11450 27268 11452
rect 27324 11450 27348 11452
rect 27404 11450 27428 11452
rect 27484 11450 27508 11452
rect 27564 11450 27570 11452
rect 27324 11398 27326 11450
rect 27506 11398 27508 11450
rect 27262 11396 27268 11398
rect 27324 11396 27348 11398
rect 27404 11396 27428 11398
rect 27484 11396 27508 11398
rect 27564 11396 27570 11398
rect 27262 11387 27570 11396
rect 27068 11212 27120 11218
rect 27068 11154 27120 11160
rect 27068 11008 27120 11014
rect 27068 10950 27120 10956
rect 26976 10124 27028 10130
rect 26976 10066 27028 10072
rect 27080 9654 27108 10950
rect 27262 10364 27570 10373
rect 27262 10362 27268 10364
rect 27324 10362 27348 10364
rect 27404 10362 27428 10364
rect 27484 10362 27508 10364
rect 27564 10362 27570 10364
rect 27324 10310 27326 10362
rect 27506 10310 27508 10362
rect 27262 10308 27268 10310
rect 27324 10308 27348 10310
rect 27404 10308 27428 10310
rect 27484 10308 27508 10310
rect 27564 10308 27570 10310
rect 27262 10299 27570 10308
rect 27068 9648 27120 9654
rect 27068 9590 27120 9596
rect 26148 9036 26200 9042
rect 26148 8978 26200 8984
rect 26240 9036 26292 9042
rect 26240 8978 26292 8984
rect 26884 9036 26936 9042
rect 26884 8978 26936 8984
rect 26056 8900 26108 8906
rect 26056 8842 26108 8848
rect 26068 8090 26096 8842
rect 26056 8084 26108 8090
rect 26056 8026 26108 8032
rect 26056 7200 26108 7206
rect 26056 7142 26108 7148
rect 25412 6860 25464 6866
rect 25412 6802 25464 6808
rect 25964 6860 26016 6866
rect 25964 6802 26016 6808
rect 25424 6458 25452 6802
rect 25688 6656 25740 6662
rect 25688 6598 25740 6604
rect 25320 6452 25372 6458
rect 25320 6394 25372 6400
rect 25412 6452 25464 6458
rect 25412 6394 25464 6400
rect 25700 6186 25728 6598
rect 25964 6316 26016 6322
rect 25964 6258 26016 6264
rect 25976 6186 26004 6258
rect 26068 6254 26096 7142
rect 26160 6866 26188 8978
rect 26252 7954 26280 8978
rect 26424 8832 26476 8838
rect 26424 8774 26476 8780
rect 26436 8090 26464 8774
rect 26884 8288 26936 8294
rect 26884 8230 26936 8236
rect 26424 8084 26476 8090
rect 26424 8026 26476 8032
rect 26240 7948 26292 7954
rect 26240 7890 26292 7896
rect 26436 7002 26464 8026
rect 26792 7880 26844 7886
rect 26792 7822 26844 7828
rect 26424 6996 26476 7002
rect 26424 6938 26476 6944
rect 26804 6866 26832 7822
rect 26896 7410 26924 8230
rect 27080 7954 27108 9590
rect 27262 9276 27570 9285
rect 27262 9274 27268 9276
rect 27324 9274 27348 9276
rect 27404 9274 27428 9276
rect 27484 9274 27508 9276
rect 27564 9274 27570 9276
rect 27324 9222 27326 9274
rect 27506 9222 27508 9274
rect 27262 9220 27268 9222
rect 27324 9220 27348 9222
rect 27404 9220 27428 9222
rect 27484 9220 27508 9222
rect 27564 9220 27570 9222
rect 27262 9211 27570 9220
rect 27262 8188 27570 8197
rect 27262 8186 27268 8188
rect 27324 8186 27348 8188
rect 27404 8186 27428 8188
rect 27484 8186 27508 8188
rect 27564 8186 27570 8188
rect 27324 8134 27326 8186
rect 27506 8134 27508 8186
rect 27262 8132 27268 8134
rect 27324 8132 27348 8134
rect 27404 8132 27428 8134
rect 27484 8132 27508 8134
rect 27564 8132 27570 8134
rect 27262 8123 27570 8132
rect 27068 7948 27120 7954
rect 27068 7890 27120 7896
rect 26884 7404 26936 7410
rect 26884 7346 26936 7352
rect 27262 7100 27570 7109
rect 27262 7098 27268 7100
rect 27324 7098 27348 7100
rect 27404 7098 27428 7100
rect 27484 7098 27508 7100
rect 27564 7098 27570 7100
rect 27324 7046 27326 7098
rect 27506 7046 27508 7098
rect 27262 7044 27268 7046
rect 27324 7044 27348 7046
rect 27404 7044 27428 7046
rect 27484 7044 27508 7046
rect 27564 7044 27570 7046
rect 27262 7035 27570 7044
rect 26148 6860 26200 6866
rect 26148 6802 26200 6808
rect 26792 6860 26844 6866
rect 26792 6802 26844 6808
rect 26056 6248 26108 6254
rect 26056 6190 26108 6196
rect 25688 6180 25740 6186
rect 25688 6122 25740 6128
rect 25964 6180 26016 6186
rect 25964 6122 26016 6128
rect 27262 6012 27570 6021
rect 27262 6010 27268 6012
rect 27324 6010 27348 6012
rect 27404 6010 27428 6012
rect 27484 6010 27508 6012
rect 27564 6010 27570 6012
rect 27324 5958 27326 6010
rect 27506 5958 27508 6010
rect 27262 5956 27268 5958
rect 27324 5956 27348 5958
rect 27404 5956 27428 5958
rect 27484 5956 27508 5958
rect 27564 5956 27570 5958
rect 27262 5947 27570 5956
rect 25228 5908 25280 5914
rect 25228 5850 25280 5856
rect 25228 5772 25280 5778
rect 25228 5714 25280 5720
rect 25412 5772 25464 5778
rect 25412 5714 25464 5720
rect 25688 5772 25740 5778
rect 25688 5714 25740 5720
rect 25240 4554 25268 5714
rect 25320 5568 25372 5574
rect 25320 5510 25372 5516
rect 25332 5166 25360 5510
rect 25320 5160 25372 5166
rect 25320 5102 25372 5108
rect 25424 4758 25452 5714
rect 25700 5030 25728 5714
rect 25688 5024 25740 5030
rect 25688 4966 25740 4972
rect 25700 4758 25728 4966
rect 27262 4924 27570 4933
rect 27262 4922 27268 4924
rect 27324 4922 27348 4924
rect 27404 4922 27428 4924
rect 27484 4922 27508 4924
rect 27564 4922 27570 4924
rect 27324 4870 27326 4922
rect 27506 4870 27508 4922
rect 27262 4868 27268 4870
rect 27324 4868 27348 4870
rect 27404 4868 27428 4870
rect 27484 4868 27508 4870
rect 27564 4868 27570 4870
rect 27262 4859 27570 4868
rect 25412 4752 25464 4758
rect 25412 4694 25464 4700
rect 25688 4752 25740 4758
rect 25688 4694 25740 4700
rect 25228 4548 25280 4554
rect 25228 4490 25280 4496
rect 25424 4282 25452 4694
rect 25412 4276 25464 4282
rect 25412 4218 25464 4224
rect 27262 3836 27570 3845
rect 27262 3834 27268 3836
rect 27324 3834 27348 3836
rect 27404 3834 27428 3836
rect 27484 3834 27508 3836
rect 27564 3834 27570 3836
rect 27324 3782 27326 3834
rect 27506 3782 27508 3834
rect 27262 3780 27268 3782
rect 27324 3780 27348 3782
rect 27404 3780 27428 3782
rect 27484 3780 27508 3782
rect 27564 3780 27570 3782
rect 27262 3771 27570 3780
rect 25136 3732 25188 3738
rect 25136 3674 25188 3680
rect 24768 3596 24820 3602
rect 24768 3538 24820 3544
rect 23904 3292 24212 3301
rect 23904 3290 23910 3292
rect 23966 3290 23990 3292
rect 24046 3290 24070 3292
rect 24126 3290 24150 3292
rect 24206 3290 24212 3292
rect 23966 3238 23968 3290
rect 24148 3238 24150 3290
rect 23904 3236 23910 3238
rect 23966 3236 23990 3238
rect 24046 3236 24070 3238
rect 24126 3236 24150 3238
rect 24206 3236 24212 3238
rect 23904 3227 24212 3236
rect 24780 3194 24808 3538
rect 25044 3392 25096 3398
rect 25044 3334 25096 3340
rect 23940 3188 23992 3194
rect 23768 3148 23940 3176
rect 23940 3130 23992 3136
rect 24308 3188 24360 3194
rect 24308 3130 24360 3136
rect 24768 3188 24820 3194
rect 24768 3130 24820 3136
rect 23664 2984 23716 2990
rect 23110 2952 23166 2961
rect 22940 2910 23060 2938
rect 22848 2746 22968 2774
rect 22940 1494 22968 2746
rect 23032 2310 23060 2910
rect 23664 2926 23716 2932
rect 24216 2984 24268 2990
rect 24216 2926 24268 2932
rect 23110 2887 23112 2896
rect 23164 2887 23166 2896
rect 23112 2858 23164 2864
rect 23124 2650 23152 2858
rect 23112 2644 23164 2650
rect 23112 2586 23164 2592
rect 24228 2378 24256 2926
rect 24320 2650 24348 3130
rect 25056 2990 25084 3334
rect 25320 3052 25372 3058
rect 25320 2994 25372 3000
rect 25044 2984 25096 2990
rect 25044 2926 25096 2932
rect 25136 2848 25188 2854
rect 25136 2790 25188 2796
rect 24308 2644 24360 2650
rect 24308 2586 24360 2592
rect 23664 2372 23716 2378
rect 23664 2314 23716 2320
rect 24216 2372 24268 2378
rect 24216 2314 24268 2320
rect 23020 2304 23072 2310
rect 23020 2246 23072 2252
rect 23572 1964 23624 1970
rect 23572 1906 23624 1912
rect 23388 1896 23440 1902
rect 23388 1838 23440 1844
rect 22928 1488 22980 1494
rect 22928 1430 22980 1436
rect 22836 1420 22888 1426
rect 22756 1380 22836 1408
rect 22376 808 22428 814
rect 22376 750 22428 756
rect 22560 808 22612 814
rect 22560 750 22612 756
rect 22756 400 22784 1380
rect 22836 1362 22888 1368
rect 23400 1358 23428 1838
rect 23388 1352 23440 1358
rect 23388 1294 23440 1300
rect 23584 1018 23612 1906
rect 23572 1012 23624 1018
rect 23572 954 23624 960
rect 23676 814 23704 2314
rect 23904 2204 24212 2213
rect 23904 2202 23910 2204
rect 23966 2202 23990 2204
rect 24046 2202 24070 2204
rect 24126 2202 24150 2204
rect 24206 2202 24212 2204
rect 23966 2150 23968 2202
rect 24148 2150 24150 2202
rect 23904 2148 23910 2150
rect 23966 2148 23990 2150
rect 24046 2148 24070 2150
rect 24126 2148 24150 2150
rect 24206 2148 24212 2150
rect 23904 2139 24212 2148
rect 24320 1902 24348 2586
rect 24860 1964 24912 1970
rect 24860 1906 24912 1912
rect 23756 1896 23808 1902
rect 23756 1838 23808 1844
rect 24308 1896 24360 1902
rect 24308 1838 24360 1844
rect 23768 882 23796 1838
rect 24872 1426 24900 1906
rect 24952 1896 25004 1902
rect 24952 1838 25004 1844
rect 24308 1420 24360 1426
rect 24308 1362 24360 1368
rect 24860 1420 24912 1426
rect 24860 1362 24912 1368
rect 23904 1116 24212 1125
rect 23904 1114 23910 1116
rect 23966 1114 23990 1116
rect 24046 1114 24070 1116
rect 24126 1114 24150 1116
rect 24206 1114 24212 1116
rect 23966 1062 23968 1114
rect 24148 1062 24150 1114
rect 23904 1060 23910 1062
rect 23966 1060 23990 1062
rect 24046 1060 24070 1062
rect 24126 1060 24150 1062
rect 24206 1060 24212 1062
rect 23904 1051 24212 1060
rect 23756 876 23808 882
rect 23756 818 23808 824
rect 23296 808 23348 814
rect 23296 750 23348 756
rect 23664 808 23716 814
rect 23664 750 23716 756
rect 23308 400 23336 750
rect 23860 462 23980 490
rect 23860 400 23888 462
rect 3528 326 3924 354
rect 3974 0 4030 400
rect 4526 0 4582 400
rect 5078 0 5134 400
rect 5630 0 5686 400
rect 6182 0 6238 400
rect 6734 0 6790 400
rect 7286 0 7342 400
rect 7838 0 7894 400
rect 8390 0 8446 400
rect 8942 0 8998 400
rect 9494 0 9550 400
rect 10046 0 10102 400
rect 10598 0 10654 400
rect 11150 0 11206 400
rect 11702 0 11758 400
rect 12254 0 12310 400
rect 12806 0 12862 400
rect 13358 0 13414 400
rect 13910 0 13966 400
rect 14462 0 14518 400
rect 15014 0 15070 400
rect 15566 0 15622 400
rect 16118 0 16174 400
rect 16670 0 16726 400
rect 17222 0 17278 400
rect 17774 0 17830 400
rect 18326 0 18382 400
rect 18878 0 18934 400
rect 19430 0 19486 400
rect 19982 0 20038 400
rect 20534 0 20590 400
rect 21086 0 21142 400
rect 21638 0 21694 400
rect 22190 0 22246 400
rect 22742 0 22798 400
rect 23294 0 23350 400
rect 23846 0 23902 400
rect 23952 354 23980 462
rect 24320 354 24348 1362
rect 24492 808 24544 814
rect 24412 768 24492 796
rect 24412 400 24440 768
rect 24492 750 24544 756
rect 24964 400 24992 1838
rect 25148 1426 25176 2790
rect 25228 1896 25280 1902
rect 25228 1838 25280 1844
rect 25136 1420 25188 1426
rect 25136 1362 25188 1368
rect 25240 814 25268 1838
rect 25332 814 25360 2994
rect 27262 2748 27570 2757
rect 27262 2746 27268 2748
rect 27324 2746 27348 2748
rect 27404 2746 27428 2748
rect 27484 2746 27508 2748
rect 27564 2746 27570 2748
rect 27324 2694 27326 2746
rect 27506 2694 27508 2746
rect 27262 2692 27268 2694
rect 27324 2692 27348 2694
rect 27404 2692 27428 2694
rect 27484 2692 27508 2694
rect 27564 2692 27570 2694
rect 27262 2683 27570 2692
rect 27262 1660 27570 1669
rect 27262 1658 27268 1660
rect 27324 1658 27348 1660
rect 27404 1658 27428 1660
rect 27484 1658 27508 1660
rect 27564 1658 27570 1660
rect 27324 1606 27326 1658
rect 27506 1606 27508 1658
rect 27262 1604 27268 1606
rect 27324 1604 27348 1606
rect 27404 1604 27428 1606
rect 27484 1604 27508 1606
rect 27564 1604 27570 1606
rect 27262 1595 27570 1604
rect 25504 1420 25556 1426
rect 25504 1362 25556 1368
rect 25228 808 25280 814
rect 25228 750 25280 756
rect 25320 808 25372 814
rect 25320 750 25372 756
rect 25516 400 25544 1362
rect 26056 808 26108 814
rect 26056 750 26108 756
rect 26068 400 26096 750
rect 27262 572 27570 581
rect 27262 570 27268 572
rect 27324 570 27348 572
rect 27404 570 27428 572
rect 27484 570 27508 572
rect 27564 570 27570 572
rect 27324 518 27326 570
rect 27506 518 27508 570
rect 27262 516 27268 518
rect 27324 516 27348 518
rect 27404 516 27428 518
rect 27484 516 27508 518
rect 27564 516 27570 518
rect 27262 507 27570 516
rect 23952 326 24348 354
rect 24398 0 24454 400
rect 24950 0 25006 400
rect 25502 0 25558 400
rect 26054 0 26110 400
<< via2 >>
rect 3762 30490 3818 30492
rect 3842 30490 3898 30492
rect 3922 30490 3978 30492
rect 4002 30490 4058 30492
rect 3762 30438 3808 30490
rect 3808 30438 3818 30490
rect 3842 30438 3872 30490
rect 3872 30438 3884 30490
rect 3884 30438 3898 30490
rect 3922 30438 3936 30490
rect 3936 30438 3948 30490
rect 3948 30438 3978 30490
rect 4002 30438 4012 30490
rect 4012 30438 4058 30490
rect 3762 30436 3818 30438
rect 3842 30436 3898 30438
rect 3922 30436 3978 30438
rect 4002 30436 4058 30438
rect 1674 15564 1730 15600
rect 1674 15544 1676 15564
rect 1676 15544 1728 15564
rect 1728 15544 1730 15564
rect 3762 29402 3818 29404
rect 3842 29402 3898 29404
rect 3922 29402 3978 29404
rect 4002 29402 4058 29404
rect 3762 29350 3808 29402
rect 3808 29350 3818 29402
rect 3842 29350 3872 29402
rect 3872 29350 3884 29402
rect 3884 29350 3898 29402
rect 3922 29350 3936 29402
rect 3936 29350 3948 29402
rect 3948 29350 3978 29402
rect 4002 29350 4012 29402
rect 4012 29350 4058 29402
rect 3762 29348 3818 29350
rect 3842 29348 3898 29350
rect 3922 29348 3978 29350
rect 4002 29348 4058 29350
rect 7120 31034 7176 31036
rect 7200 31034 7256 31036
rect 7280 31034 7336 31036
rect 7360 31034 7416 31036
rect 7120 30982 7166 31034
rect 7166 30982 7176 31034
rect 7200 30982 7230 31034
rect 7230 30982 7242 31034
rect 7242 30982 7256 31034
rect 7280 30982 7294 31034
rect 7294 30982 7306 31034
rect 7306 30982 7336 31034
rect 7360 30982 7370 31034
rect 7370 30982 7416 31034
rect 7120 30980 7176 30982
rect 7200 30980 7256 30982
rect 7280 30980 7336 30982
rect 7360 30980 7416 30982
rect 3762 28314 3818 28316
rect 3842 28314 3898 28316
rect 3922 28314 3978 28316
rect 4002 28314 4058 28316
rect 3762 28262 3808 28314
rect 3808 28262 3818 28314
rect 3842 28262 3872 28314
rect 3872 28262 3884 28314
rect 3884 28262 3898 28314
rect 3922 28262 3936 28314
rect 3936 28262 3948 28314
rect 3948 28262 3978 28314
rect 4002 28262 4012 28314
rect 4012 28262 4058 28314
rect 3762 28260 3818 28262
rect 3842 28260 3898 28262
rect 3922 28260 3978 28262
rect 4002 28260 4058 28262
rect 3762 27226 3818 27228
rect 3842 27226 3898 27228
rect 3922 27226 3978 27228
rect 4002 27226 4058 27228
rect 3762 27174 3808 27226
rect 3808 27174 3818 27226
rect 3842 27174 3872 27226
rect 3872 27174 3884 27226
rect 3884 27174 3898 27226
rect 3922 27174 3936 27226
rect 3936 27174 3948 27226
rect 3948 27174 3978 27226
rect 4002 27174 4012 27226
rect 4012 27174 4058 27226
rect 3762 27172 3818 27174
rect 3842 27172 3898 27174
rect 3922 27172 3978 27174
rect 4002 27172 4058 27174
rect 3762 26138 3818 26140
rect 3842 26138 3898 26140
rect 3922 26138 3978 26140
rect 4002 26138 4058 26140
rect 3762 26086 3808 26138
rect 3808 26086 3818 26138
rect 3842 26086 3872 26138
rect 3872 26086 3884 26138
rect 3884 26086 3898 26138
rect 3922 26086 3936 26138
rect 3936 26086 3948 26138
rect 3948 26086 3978 26138
rect 4002 26086 4012 26138
rect 4012 26086 4058 26138
rect 3762 26084 3818 26086
rect 3842 26084 3898 26086
rect 3922 26084 3978 26086
rect 4002 26084 4058 26086
rect 3762 25050 3818 25052
rect 3842 25050 3898 25052
rect 3922 25050 3978 25052
rect 4002 25050 4058 25052
rect 3762 24998 3808 25050
rect 3808 24998 3818 25050
rect 3842 24998 3872 25050
rect 3872 24998 3884 25050
rect 3884 24998 3898 25050
rect 3922 24998 3936 25050
rect 3936 24998 3948 25050
rect 3948 24998 3978 25050
rect 4002 24998 4012 25050
rect 4012 24998 4058 25050
rect 3762 24996 3818 24998
rect 3842 24996 3898 24998
rect 3922 24996 3978 24998
rect 4002 24996 4058 24998
rect 3762 23962 3818 23964
rect 3842 23962 3898 23964
rect 3922 23962 3978 23964
rect 4002 23962 4058 23964
rect 3762 23910 3808 23962
rect 3808 23910 3818 23962
rect 3842 23910 3872 23962
rect 3872 23910 3884 23962
rect 3884 23910 3898 23962
rect 3922 23910 3936 23962
rect 3936 23910 3948 23962
rect 3948 23910 3978 23962
rect 4002 23910 4012 23962
rect 4012 23910 4058 23962
rect 3762 23908 3818 23910
rect 3842 23908 3898 23910
rect 3922 23908 3978 23910
rect 4002 23908 4058 23910
rect 3790 23604 3792 23624
rect 3792 23604 3844 23624
rect 3844 23604 3846 23624
rect 3790 23568 3846 23604
rect 3762 22874 3818 22876
rect 3842 22874 3898 22876
rect 3922 22874 3978 22876
rect 4002 22874 4058 22876
rect 3762 22822 3808 22874
rect 3808 22822 3818 22874
rect 3842 22822 3872 22874
rect 3872 22822 3884 22874
rect 3884 22822 3898 22874
rect 3922 22822 3936 22874
rect 3936 22822 3948 22874
rect 3948 22822 3978 22874
rect 4002 22822 4012 22874
rect 4012 22822 4058 22874
rect 3762 22820 3818 22822
rect 3842 22820 3898 22822
rect 3922 22820 3978 22822
rect 4002 22820 4058 22822
rect 5906 26288 5962 26344
rect 4986 23604 4988 23624
rect 4988 23604 5040 23624
rect 5040 23604 5042 23624
rect 4986 23568 5042 23604
rect 2318 10004 2320 10024
rect 2320 10004 2372 10024
rect 2372 10004 2374 10024
rect 2318 9968 2374 10004
rect 3762 21786 3818 21788
rect 3842 21786 3898 21788
rect 3922 21786 3978 21788
rect 4002 21786 4058 21788
rect 3762 21734 3808 21786
rect 3808 21734 3818 21786
rect 3842 21734 3872 21786
rect 3872 21734 3884 21786
rect 3884 21734 3898 21786
rect 3922 21734 3936 21786
rect 3936 21734 3948 21786
rect 3948 21734 3978 21786
rect 4002 21734 4012 21786
rect 4012 21734 4058 21786
rect 3762 21732 3818 21734
rect 3842 21732 3898 21734
rect 3922 21732 3978 21734
rect 4002 21732 4058 21734
rect 3762 20698 3818 20700
rect 3842 20698 3898 20700
rect 3922 20698 3978 20700
rect 4002 20698 4058 20700
rect 3762 20646 3808 20698
rect 3808 20646 3818 20698
rect 3842 20646 3872 20698
rect 3872 20646 3884 20698
rect 3884 20646 3898 20698
rect 3922 20646 3936 20698
rect 3936 20646 3948 20698
rect 3948 20646 3978 20698
rect 4002 20646 4012 20698
rect 4012 20646 4058 20698
rect 3762 20644 3818 20646
rect 3842 20644 3898 20646
rect 3922 20644 3978 20646
rect 4002 20644 4058 20646
rect 3762 19610 3818 19612
rect 3842 19610 3898 19612
rect 3922 19610 3978 19612
rect 4002 19610 4058 19612
rect 3762 19558 3808 19610
rect 3808 19558 3818 19610
rect 3842 19558 3872 19610
rect 3872 19558 3884 19610
rect 3884 19558 3898 19610
rect 3922 19558 3936 19610
rect 3936 19558 3948 19610
rect 3948 19558 3978 19610
rect 4002 19558 4012 19610
rect 4012 19558 4058 19610
rect 3762 19556 3818 19558
rect 3842 19556 3898 19558
rect 3922 19556 3978 19558
rect 4002 19556 4058 19558
rect 5354 21972 5356 21992
rect 5356 21972 5408 21992
rect 5408 21972 5410 21992
rect 5354 21936 5410 21972
rect 3762 18522 3818 18524
rect 3842 18522 3898 18524
rect 3922 18522 3978 18524
rect 4002 18522 4058 18524
rect 3762 18470 3808 18522
rect 3808 18470 3818 18522
rect 3842 18470 3872 18522
rect 3872 18470 3884 18522
rect 3884 18470 3898 18522
rect 3922 18470 3936 18522
rect 3936 18470 3948 18522
rect 3948 18470 3978 18522
rect 4002 18470 4012 18522
rect 4012 18470 4058 18522
rect 3762 18468 3818 18470
rect 3842 18468 3898 18470
rect 3922 18468 3978 18470
rect 4002 18468 4058 18470
rect 3762 17434 3818 17436
rect 3842 17434 3898 17436
rect 3922 17434 3978 17436
rect 4002 17434 4058 17436
rect 3762 17382 3808 17434
rect 3808 17382 3818 17434
rect 3842 17382 3872 17434
rect 3872 17382 3884 17434
rect 3884 17382 3898 17434
rect 3922 17382 3936 17434
rect 3936 17382 3948 17434
rect 3948 17382 3978 17434
rect 4002 17382 4012 17434
rect 4012 17382 4058 17434
rect 3762 17380 3818 17382
rect 3842 17380 3898 17382
rect 3922 17380 3978 17382
rect 4002 17380 4058 17382
rect 3762 16346 3818 16348
rect 3842 16346 3898 16348
rect 3922 16346 3978 16348
rect 4002 16346 4058 16348
rect 3762 16294 3808 16346
rect 3808 16294 3818 16346
rect 3842 16294 3872 16346
rect 3872 16294 3884 16346
rect 3884 16294 3898 16346
rect 3922 16294 3936 16346
rect 3936 16294 3948 16346
rect 3948 16294 3978 16346
rect 4002 16294 4012 16346
rect 4012 16294 4058 16346
rect 3762 16292 3818 16294
rect 3842 16292 3898 16294
rect 3922 16292 3978 16294
rect 4002 16292 4058 16294
rect 6182 23180 6238 23216
rect 6182 23160 6184 23180
rect 6184 23160 6236 23180
rect 6236 23160 6238 23180
rect 7120 29946 7176 29948
rect 7200 29946 7256 29948
rect 7280 29946 7336 29948
rect 7360 29946 7416 29948
rect 7120 29894 7166 29946
rect 7166 29894 7176 29946
rect 7200 29894 7230 29946
rect 7230 29894 7242 29946
rect 7242 29894 7256 29946
rect 7280 29894 7294 29946
rect 7294 29894 7306 29946
rect 7306 29894 7336 29946
rect 7360 29894 7370 29946
rect 7370 29894 7416 29946
rect 7120 29892 7176 29894
rect 7200 29892 7256 29894
rect 7280 29892 7336 29894
rect 7360 29892 7416 29894
rect 7120 28858 7176 28860
rect 7200 28858 7256 28860
rect 7280 28858 7336 28860
rect 7360 28858 7416 28860
rect 7120 28806 7166 28858
rect 7166 28806 7176 28858
rect 7200 28806 7230 28858
rect 7230 28806 7242 28858
rect 7242 28806 7256 28858
rect 7280 28806 7294 28858
rect 7294 28806 7306 28858
rect 7306 28806 7336 28858
rect 7360 28806 7370 28858
rect 7370 28806 7416 28858
rect 7120 28804 7176 28806
rect 7200 28804 7256 28806
rect 7280 28804 7336 28806
rect 7360 28804 7416 28806
rect 7120 27770 7176 27772
rect 7200 27770 7256 27772
rect 7280 27770 7336 27772
rect 7360 27770 7416 27772
rect 7120 27718 7166 27770
rect 7166 27718 7176 27770
rect 7200 27718 7230 27770
rect 7230 27718 7242 27770
rect 7242 27718 7256 27770
rect 7280 27718 7294 27770
rect 7294 27718 7306 27770
rect 7306 27718 7336 27770
rect 7360 27718 7370 27770
rect 7370 27718 7416 27770
rect 7120 27716 7176 27718
rect 7200 27716 7256 27718
rect 7280 27716 7336 27718
rect 7360 27716 7416 27718
rect 6734 26288 6790 26344
rect 10478 30490 10534 30492
rect 10558 30490 10614 30492
rect 10638 30490 10694 30492
rect 10718 30490 10774 30492
rect 10478 30438 10524 30490
rect 10524 30438 10534 30490
rect 10558 30438 10588 30490
rect 10588 30438 10600 30490
rect 10600 30438 10614 30490
rect 10638 30438 10652 30490
rect 10652 30438 10664 30490
rect 10664 30438 10694 30490
rect 10718 30438 10728 30490
rect 10728 30438 10774 30490
rect 10478 30436 10534 30438
rect 10558 30436 10614 30438
rect 10638 30436 10694 30438
rect 10718 30436 10774 30438
rect 7120 26682 7176 26684
rect 7200 26682 7256 26684
rect 7280 26682 7336 26684
rect 7360 26682 7416 26684
rect 7120 26630 7166 26682
rect 7166 26630 7176 26682
rect 7200 26630 7230 26682
rect 7230 26630 7242 26682
rect 7242 26630 7256 26682
rect 7280 26630 7294 26682
rect 7294 26630 7306 26682
rect 7306 26630 7336 26682
rect 7360 26630 7370 26682
rect 7370 26630 7416 26682
rect 7120 26628 7176 26630
rect 7200 26628 7256 26630
rect 7280 26628 7336 26630
rect 7360 26628 7416 26630
rect 10478 29402 10534 29404
rect 10558 29402 10614 29404
rect 10638 29402 10694 29404
rect 10718 29402 10774 29404
rect 10478 29350 10524 29402
rect 10524 29350 10534 29402
rect 10558 29350 10588 29402
rect 10588 29350 10600 29402
rect 10600 29350 10614 29402
rect 10638 29350 10652 29402
rect 10652 29350 10664 29402
rect 10664 29350 10694 29402
rect 10718 29350 10728 29402
rect 10728 29350 10774 29402
rect 10478 29348 10534 29350
rect 10558 29348 10614 29350
rect 10638 29348 10694 29350
rect 10718 29348 10774 29350
rect 10478 28314 10534 28316
rect 10558 28314 10614 28316
rect 10638 28314 10694 28316
rect 10718 28314 10774 28316
rect 10478 28262 10524 28314
rect 10524 28262 10534 28314
rect 10558 28262 10588 28314
rect 10588 28262 10600 28314
rect 10600 28262 10614 28314
rect 10638 28262 10652 28314
rect 10652 28262 10664 28314
rect 10664 28262 10694 28314
rect 10718 28262 10728 28314
rect 10728 28262 10774 28314
rect 10478 28260 10534 28262
rect 10558 28260 10614 28262
rect 10638 28260 10694 28262
rect 10718 28260 10774 28262
rect 13836 31034 13892 31036
rect 13916 31034 13972 31036
rect 13996 31034 14052 31036
rect 14076 31034 14132 31036
rect 13836 30982 13882 31034
rect 13882 30982 13892 31034
rect 13916 30982 13946 31034
rect 13946 30982 13958 31034
rect 13958 30982 13972 31034
rect 13996 30982 14010 31034
rect 14010 30982 14022 31034
rect 14022 30982 14052 31034
rect 14076 30982 14086 31034
rect 14086 30982 14132 31034
rect 13836 30980 13892 30982
rect 13916 30980 13972 30982
rect 13996 30980 14052 30982
rect 14076 30980 14132 30982
rect 20552 31034 20608 31036
rect 20632 31034 20688 31036
rect 20712 31034 20768 31036
rect 20792 31034 20848 31036
rect 20552 30982 20598 31034
rect 20598 30982 20608 31034
rect 20632 30982 20662 31034
rect 20662 30982 20674 31034
rect 20674 30982 20688 31034
rect 20712 30982 20726 31034
rect 20726 30982 20738 31034
rect 20738 30982 20768 31034
rect 20792 30982 20802 31034
rect 20802 30982 20848 31034
rect 20552 30980 20608 30982
rect 20632 30980 20688 30982
rect 20712 30980 20768 30982
rect 20792 30980 20848 30982
rect 17682 30796 17738 30832
rect 17682 30776 17684 30796
rect 17684 30776 17736 30796
rect 17736 30776 17738 30796
rect 19062 30796 19118 30832
rect 19062 30776 19064 30796
rect 19064 30776 19116 30796
rect 19116 30776 19118 30796
rect 7120 25594 7176 25596
rect 7200 25594 7256 25596
rect 7280 25594 7336 25596
rect 7360 25594 7416 25596
rect 7120 25542 7166 25594
rect 7166 25542 7176 25594
rect 7200 25542 7230 25594
rect 7230 25542 7242 25594
rect 7242 25542 7256 25594
rect 7280 25542 7294 25594
rect 7294 25542 7306 25594
rect 7306 25542 7336 25594
rect 7360 25542 7370 25594
rect 7370 25542 7416 25594
rect 7120 25540 7176 25542
rect 7200 25540 7256 25542
rect 7280 25540 7336 25542
rect 7360 25540 7416 25542
rect 6642 23296 6698 23352
rect 7120 24506 7176 24508
rect 7200 24506 7256 24508
rect 7280 24506 7336 24508
rect 7360 24506 7416 24508
rect 7120 24454 7166 24506
rect 7166 24454 7176 24506
rect 7200 24454 7230 24506
rect 7230 24454 7242 24506
rect 7242 24454 7256 24506
rect 7280 24454 7294 24506
rect 7294 24454 7306 24506
rect 7306 24454 7336 24506
rect 7360 24454 7370 24506
rect 7370 24454 7416 24506
rect 7120 24452 7176 24454
rect 7200 24452 7256 24454
rect 7280 24452 7336 24454
rect 7360 24452 7416 24454
rect 7120 23418 7176 23420
rect 7200 23418 7256 23420
rect 7280 23418 7336 23420
rect 7360 23418 7416 23420
rect 7120 23366 7166 23418
rect 7166 23366 7176 23418
rect 7200 23366 7230 23418
rect 7230 23366 7242 23418
rect 7242 23366 7256 23418
rect 7280 23366 7294 23418
rect 7294 23366 7306 23418
rect 7306 23366 7336 23418
rect 7360 23366 7370 23418
rect 7370 23366 7416 23418
rect 7120 23364 7176 23366
rect 7200 23364 7256 23366
rect 7280 23364 7336 23366
rect 7360 23364 7416 23366
rect 3762 15258 3818 15260
rect 3842 15258 3898 15260
rect 3922 15258 3978 15260
rect 4002 15258 4058 15260
rect 3762 15206 3808 15258
rect 3808 15206 3818 15258
rect 3842 15206 3872 15258
rect 3872 15206 3884 15258
rect 3884 15206 3898 15258
rect 3922 15206 3936 15258
rect 3936 15206 3948 15258
rect 3948 15206 3978 15258
rect 4002 15206 4012 15258
rect 4012 15206 4058 15258
rect 3762 15204 3818 15206
rect 3842 15204 3898 15206
rect 3922 15204 3978 15206
rect 4002 15204 4058 15206
rect 3762 14170 3818 14172
rect 3842 14170 3898 14172
rect 3922 14170 3978 14172
rect 4002 14170 4058 14172
rect 3762 14118 3808 14170
rect 3808 14118 3818 14170
rect 3842 14118 3872 14170
rect 3872 14118 3884 14170
rect 3884 14118 3898 14170
rect 3922 14118 3936 14170
rect 3936 14118 3948 14170
rect 3948 14118 3978 14170
rect 4002 14118 4012 14170
rect 4012 14118 4058 14170
rect 3762 14116 3818 14118
rect 3842 14116 3898 14118
rect 3922 14116 3978 14118
rect 4002 14116 4058 14118
rect 3762 13082 3818 13084
rect 3842 13082 3898 13084
rect 3922 13082 3978 13084
rect 4002 13082 4058 13084
rect 3762 13030 3808 13082
rect 3808 13030 3818 13082
rect 3842 13030 3872 13082
rect 3872 13030 3884 13082
rect 3884 13030 3898 13082
rect 3922 13030 3936 13082
rect 3936 13030 3948 13082
rect 3948 13030 3978 13082
rect 4002 13030 4012 13082
rect 4012 13030 4058 13082
rect 3762 13028 3818 13030
rect 3842 13028 3898 13030
rect 3922 13028 3978 13030
rect 4002 13028 4058 13030
rect 3762 11994 3818 11996
rect 3842 11994 3898 11996
rect 3922 11994 3978 11996
rect 4002 11994 4058 11996
rect 3762 11942 3808 11994
rect 3808 11942 3818 11994
rect 3842 11942 3872 11994
rect 3872 11942 3884 11994
rect 3884 11942 3898 11994
rect 3922 11942 3936 11994
rect 3936 11942 3948 11994
rect 3948 11942 3978 11994
rect 4002 11942 4012 11994
rect 4012 11942 4058 11994
rect 3762 11940 3818 11942
rect 3842 11940 3898 11942
rect 3922 11940 3978 11942
rect 4002 11940 4058 11942
rect 3762 10906 3818 10908
rect 3842 10906 3898 10908
rect 3922 10906 3978 10908
rect 4002 10906 4058 10908
rect 3762 10854 3808 10906
rect 3808 10854 3818 10906
rect 3842 10854 3872 10906
rect 3872 10854 3884 10906
rect 3884 10854 3898 10906
rect 3922 10854 3936 10906
rect 3936 10854 3948 10906
rect 3948 10854 3978 10906
rect 4002 10854 4012 10906
rect 4012 10854 4058 10906
rect 3762 10852 3818 10854
rect 3842 10852 3898 10854
rect 3922 10852 3978 10854
rect 4002 10852 4058 10854
rect 2870 10140 2872 10160
rect 2872 10140 2924 10160
rect 2924 10140 2926 10160
rect 2870 10104 2926 10140
rect 3146 9968 3202 10024
rect 4250 10104 4306 10160
rect 3762 9818 3818 9820
rect 3842 9818 3898 9820
rect 3922 9818 3978 9820
rect 4002 9818 4058 9820
rect 3762 9766 3808 9818
rect 3808 9766 3818 9818
rect 3842 9766 3872 9818
rect 3872 9766 3884 9818
rect 3884 9766 3898 9818
rect 3922 9766 3936 9818
rect 3936 9766 3948 9818
rect 3948 9766 3978 9818
rect 4002 9766 4012 9818
rect 4012 9766 4058 9818
rect 3762 9764 3818 9766
rect 3842 9764 3898 9766
rect 3922 9764 3978 9766
rect 4002 9764 4058 9766
rect 3762 8730 3818 8732
rect 3842 8730 3898 8732
rect 3922 8730 3978 8732
rect 4002 8730 4058 8732
rect 3762 8678 3808 8730
rect 3808 8678 3818 8730
rect 3842 8678 3872 8730
rect 3872 8678 3884 8730
rect 3884 8678 3898 8730
rect 3922 8678 3936 8730
rect 3936 8678 3948 8730
rect 3948 8678 3978 8730
rect 4002 8678 4012 8730
rect 4012 8678 4058 8730
rect 3762 8676 3818 8678
rect 3842 8676 3898 8678
rect 3922 8676 3978 8678
rect 4002 8676 4058 8678
rect 3762 7642 3818 7644
rect 3842 7642 3898 7644
rect 3922 7642 3978 7644
rect 4002 7642 4058 7644
rect 3762 7590 3808 7642
rect 3808 7590 3818 7642
rect 3842 7590 3872 7642
rect 3872 7590 3884 7642
rect 3884 7590 3898 7642
rect 3922 7590 3936 7642
rect 3936 7590 3948 7642
rect 3948 7590 3978 7642
rect 4002 7590 4012 7642
rect 4012 7590 4058 7642
rect 3762 7588 3818 7590
rect 3842 7588 3898 7590
rect 3922 7588 3978 7590
rect 4002 7588 4058 7590
rect 7120 22330 7176 22332
rect 7200 22330 7256 22332
rect 7280 22330 7336 22332
rect 7360 22330 7416 22332
rect 7120 22278 7166 22330
rect 7166 22278 7176 22330
rect 7200 22278 7230 22330
rect 7230 22278 7242 22330
rect 7242 22278 7256 22330
rect 7280 22278 7294 22330
rect 7294 22278 7306 22330
rect 7306 22278 7336 22330
rect 7360 22278 7370 22330
rect 7370 22278 7416 22330
rect 7120 22276 7176 22278
rect 7200 22276 7256 22278
rect 7280 22276 7336 22278
rect 7360 22276 7416 22278
rect 7746 23160 7802 23216
rect 7120 21242 7176 21244
rect 7200 21242 7256 21244
rect 7280 21242 7336 21244
rect 7360 21242 7416 21244
rect 7120 21190 7166 21242
rect 7166 21190 7176 21242
rect 7200 21190 7230 21242
rect 7230 21190 7242 21242
rect 7242 21190 7256 21242
rect 7280 21190 7294 21242
rect 7294 21190 7306 21242
rect 7306 21190 7336 21242
rect 7360 21190 7370 21242
rect 7370 21190 7416 21242
rect 7120 21188 7176 21190
rect 7200 21188 7256 21190
rect 7280 21188 7336 21190
rect 7360 21188 7416 21190
rect 7120 20154 7176 20156
rect 7200 20154 7256 20156
rect 7280 20154 7336 20156
rect 7360 20154 7416 20156
rect 7120 20102 7166 20154
rect 7166 20102 7176 20154
rect 7200 20102 7230 20154
rect 7230 20102 7242 20154
rect 7242 20102 7256 20154
rect 7280 20102 7294 20154
rect 7294 20102 7306 20154
rect 7306 20102 7336 20154
rect 7360 20102 7370 20154
rect 7370 20102 7416 20154
rect 7120 20100 7176 20102
rect 7200 20100 7256 20102
rect 7280 20100 7336 20102
rect 7360 20100 7416 20102
rect 7120 19066 7176 19068
rect 7200 19066 7256 19068
rect 7280 19066 7336 19068
rect 7360 19066 7416 19068
rect 7120 19014 7166 19066
rect 7166 19014 7176 19066
rect 7200 19014 7230 19066
rect 7230 19014 7242 19066
rect 7242 19014 7256 19066
rect 7280 19014 7294 19066
rect 7294 19014 7306 19066
rect 7306 19014 7336 19066
rect 7360 19014 7370 19066
rect 7370 19014 7416 19066
rect 7120 19012 7176 19014
rect 7200 19012 7256 19014
rect 7280 19012 7336 19014
rect 7360 19012 7416 19014
rect 7120 17978 7176 17980
rect 7200 17978 7256 17980
rect 7280 17978 7336 17980
rect 7360 17978 7416 17980
rect 7120 17926 7166 17978
rect 7166 17926 7176 17978
rect 7200 17926 7230 17978
rect 7230 17926 7242 17978
rect 7242 17926 7256 17978
rect 7280 17926 7294 17978
rect 7294 17926 7306 17978
rect 7306 17926 7336 17978
rect 7360 17926 7370 17978
rect 7370 17926 7416 17978
rect 7120 17924 7176 17926
rect 7200 17924 7256 17926
rect 7280 17924 7336 17926
rect 7360 17924 7416 17926
rect 7120 16890 7176 16892
rect 7200 16890 7256 16892
rect 7280 16890 7336 16892
rect 7360 16890 7416 16892
rect 7120 16838 7166 16890
rect 7166 16838 7176 16890
rect 7200 16838 7230 16890
rect 7230 16838 7242 16890
rect 7242 16838 7256 16890
rect 7280 16838 7294 16890
rect 7294 16838 7306 16890
rect 7306 16838 7336 16890
rect 7360 16838 7370 16890
rect 7370 16838 7416 16890
rect 7120 16836 7176 16838
rect 7200 16836 7256 16838
rect 7280 16836 7336 16838
rect 7360 16836 7416 16838
rect 10478 27226 10534 27228
rect 10558 27226 10614 27228
rect 10638 27226 10694 27228
rect 10718 27226 10774 27228
rect 10478 27174 10524 27226
rect 10524 27174 10534 27226
rect 10558 27174 10588 27226
rect 10588 27174 10600 27226
rect 10600 27174 10614 27226
rect 10638 27174 10652 27226
rect 10652 27174 10664 27226
rect 10664 27174 10694 27226
rect 10718 27174 10728 27226
rect 10728 27174 10774 27226
rect 10478 27172 10534 27174
rect 10558 27172 10614 27174
rect 10638 27172 10694 27174
rect 10718 27172 10774 27174
rect 10478 26138 10534 26140
rect 10558 26138 10614 26140
rect 10638 26138 10694 26140
rect 10718 26138 10774 26140
rect 10478 26086 10524 26138
rect 10524 26086 10534 26138
rect 10558 26086 10588 26138
rect 10588 26086 10600 26138
rect 10600 26086 10614 26138
rect 10638 26086 10652 26138
rect 10652 26086 10664 26138
rect 10664 26086 10694 26138
rect 10718 26086 10728 26138
rect 10728 26086 10774 26138
rect 10478 26084 10534 26086
rect 10558 26084 10614 26086
rect 10638 26084 10694 26086
rect 10718 26084 10774 26086
rect 10478 25050 10534 25052
rect 10558 25050 10614 25052
rect 10638 25050 10694 25052
rect 10718 25050 10774 25052
rect 10478 24998 10524 25050
rect 10524 24998 10534 25050
rect 10558 24998 10588 25050
rect 10588 24998 10600 25050
rect 10600 24998 10614 25050
rect 10638 24998 10652 25050
rect 10652 24998 10664 25050
rect 10664 24998 10694 25050
rect 10718 24998 10728 25050
rect 10728 24998 10774 25050
rect 10478 24996 10534 24998
rect 10558 24996 10614 24998
rect 10638 24996 10694 24998
rect 10718 24996 10774 24998
rect 10478 23962 10534 23964
rect 10558 23962 10614 23964
rect 10638 23962 10694 23964
rect 10718 23962 10774 23964
rect 10478 23910 10524 23962
rect 10524 23910 10534 23962
rect 10558 23910 10588 23962
rect 10588 23910 10600 23962
rect 10600 23910 10614 23962
rect 10638 23910 10652 23962
rect 10652 23910 10664 23962
rect 10664 23910 10694 23962
rect 10718 23910 10728 23962
rect 10728 23910 10774 23962
rect 10478 23908 10534 23910
rect 10558 23908 10614 23910
rect 10638 23908 10694 23910
rect 10718 23908 10774 23910
rect 10322 23180 10378 23216
rect 10322 23160 10324 23180
rect 10324 23160 10376 23180
rect 10376 23160 10378 23180
rect 9678 21004 9734 21040
rect 9678 20984 9680 21004
rect 9680 20984 9732 21004
rect 9732 20984 9734 21004
rect 9678 20440 9734 20496
rect 7120 15802 7176 15804
rect 7200 15802 7256 15804
rect 7280 15802 7336 15804
rect 7360 15802 7416 15804
rect 7120 15750 7166 15802
rect 7166 15750 7176 15802
rect 7200 15750 7230 15802
rect 7230 15750 7242 15802
rect 7242 15750 7256 15802
rect 7280 15750 7294 15802
rect 7294 15750 7306 15802
rect 7306 15750 7336 15802
rect 7360 15750 7370 15802
rect 7370 15750 7416 15802
rect 7120 15748 7176 15750
rect 7200 15748 7256 15750
rect 7280 15748 7336 15750
rect 7360 15748 7416 15750
rect 7120 14714 7176 14716
rect 7200 14714 7256 14716
rect 7280 14714 7336 14716
rect 7360 14714 7416 14716
rect 7120 14662 7166 14714
rect 7166 14662 7176 14714
rect 7200 14662 7230 14714
rect 7230 14662 7242 14714
rect 7242 14662 7256 14714
rect 7280 14662 7294 14714
rect 7294 14662 7306 14714
rect 7306 14662 7336 14714
rect 7360 14662 7370 14714
rect 7370 14662 7416 14714
rect 7120 14660 7176 14662
rect 7200 14660 7256 14662
rect 7280 14660 7336 14662
rect 7360 14660 7416 14662
rect 7120 13626 7176 13628
rect 7200 13626 7256 13628
rect 7280 13626 7336 13628
rect 7360 13626 7416 13628
rect 7120 13574 7166 13626
rect 7166 13574 7176 13626
rect 7200 13574 7230 13626
rect 7230 13574 7242 13626
rect 7242 13574 7256 13626
rect 7280 13574 7294 13626
rect 7294 13574 7306 13626
rect 7306 13574 7336 13626
rect 7360 13574 7370 13626
rect 7370 13574 7416 13626
rect 7120 13572 7176 13574
rect 7200 13572 7256 13574
rect 7280 13572 7336 13574
rect 7360 13572 7416 13574
rect 7120 12538 7176 12540
rect 7200 12538 7256 12540
rect 7280 12538 7336 12540
rect 7360 12538 7416 12540
rect 7120 12486 7166 12538
rect 7166 12486 7176 12538
rect 7200 12486 7230 12538
rect 7230 12486 7242 12538
rect 7242 12486 7256 12538
rect 7280 12486 7294 12538
rect 7294 12486 7306 12538
rect 7306 12486 7336 12538
rect 7360 12486 7370 12538
rect 7370 12486 7416 12538
rect 7120 12484 7176 12486
rect 7200 12484 7256 12486
rect 7280 12484 7336 12486
rect 7360 12484 7416 12486
rect 7120 11450 7176 11452
rect 7200 11450 7256 11452
rect 7280 11450 7336 11452
rect 7360 11450 7416 11452
rect 7120 11398 7166 11450
rect 7166 11398 7176 11450
rect 7200 11398 7230 11450
rect 7230 11398 7242 11450
rect 7242 11398 7256 11450
rect 7280 11398 7294 11450
rect 7294 11398 7306 11450
rect 7306 11398 7336 11450
rect 7360 11398 7370 11450
rect 7370 11398 7416 11450
rect 7120 11396 7176 11398
rect 7200 11396 7256 11398
rect 7280 11396 7336 11398
rect 7360 11396 7416 11398
rect 9494 16632 9550 16688
rect 7120 10362 7176 10364
rect 7200 10362 7256 10364
rect 7280 10362 7336 10364
rect 7360 10362 7416 10364
rect 7120 10310 7166 10362
rect 7166 10310 7176 10362
rect 7200 10310 7230 10362
rect 7230 10310 7242 10362
rect 7242 10310 7256 10362
rect 7280 10310 7294 10362
rect 7294 10310 7306 10362
rect 7306 10310 7336 10362
rect 7360 10310 7370 10362
rect 7370 10310 7416 10362
rect 7120 10308 7176 10310
rect 7200 10308 7256 10310
rect 7280 10308 7336 10310
rect 7360 10308 7416 10310
rect 7120 9274 7176 9276
rect 7200 9274 7256 9276
rect 7280 9274 7336 9276
rect 7360 9274 7416 9276
rect 7120 9222 7166 9274
rect 7166 9222 7176 9274
rect 7200 9222 7230 9274
rect 7230 9222 7242 9274
rect 7242 9222 7256 9274
rect 7280 9222 7294 9274
rect 7294 9222 7306 9274
rect 7306 9222 7336 9274
rect 7360 9222 7370 9274
rect 7370 9222 7416 9274
rect 7120 9220 7176 9222
rect 7200 9220 7256 9222
rect 7280 9220 7336 9222
rect 7360 9220 7416 9222
rect 7120 8186 7176 8188
rect 7200 8186 7256 8188
rect 7280 8186 7336 8188
rect 7360 8186 7416 8188
rect 7120 8134 7166 8186
rect 7166 8134 7176 8186
rect 7200 8134 7230 8186
rect 7230 8134 7242 8186
rect 7242 8134 7256 8186
rect 7280 8134 7294 8186
rect 7294 8134 7306 8186
rect 7306 8134 7336 8186
rect 7360 8134 7370 8186
rect 7370 8134 7416 8186
rect 7120 8132 7176 8134
rect 7200 8132 7256 8134
rect 7280 8132 7336 8134
rect 7360 8132 7416 8134
rect 3762 6554 3818 6556
rect 3842 6554 3898 6556
rect 3922 6554 3978 6556
rect 4002 6554 4058 6556
rect 3762 6502 3808 6554
rect 3808 6502 3818 6554
rect 3842 6502 3872 6554
rect 3872 6502 3884 6554
rect 3884 6502 3898 6554
rect 3922 6502 3936 6554
rect 3936 6502 3948 6554
rect 3948 6502 3978 6554
rect 4002 6502 4012 6554
rect 4012 6502 4058 6554
rect 3762 6500 3818 6502
rect 3842 6500 3898 6502
rect 3922 6500 3978 6502
rect 4002 6500 4058 6502
rect 3762 5466 3818 5468
rect 3842 5466 3898 5468
rect 3922 5466 3978 5468
rect 4002 5466 4058 5468
rect 3762 5414 3808 5466
rect 3808 5414 3818 5466
rect 3842 5414 3872 5466
rect 3872 5414 3884 5466
rect 3884 5414 3898 5466
rect 3922 5414 3936 5466
rect 3936 5414 3948 5466
rect 3948 5414 3978 5466
rect 4002 5414 4012 5466
rect 4012 5414 4058 5466
rect 3762 5412 3818 5414
rect 3842 5412 3898 5414
rect 3922 5412 3978 5414
rect 4002 5412 4058 5414
rect 7120 7098 7176 7100
rect 7200 7098 7256 7100
rect 7280 7098 7336 7100
rect 7360 7098 7416 7100
rect 7120 7046 7166 7098
rect 7166 7046 7176 7098
rect 7200 7046 7230 7098
rect 7230 7046 7242 7098
rect 7242 7046 7256 7098
rect 7280 7046 7294 7098
rect 7294 7046 7306 7098
rect 7306 7046 7336 7098
rect 7360 7046 7370 7098
rect 7370 7046 7416 7098
rect 7120 7044 7176 7046
rect 7200 7044 7256 7046
rect 7280 7044 7336 7046
rect 7360 7044 7416 7046
rect 3762 4378 3818 4380
rect 3842 4378 3898 4380
rect 3922 4378 3978 4380
rect 4002 4378 4058 4380
rect 3762 4326 3808 4378
rect 3808 4326 3818 4378
rect 3842 4326 3872 4378
rect 3872 4326 3884 4378
rect 3884 4326 3898 4378
rect 3922 4326 3936 4378
rect 3936 4326 3948 4378
rect 3948 4326 3978 4378
rect 4002 4326 4012 4378
rect 4012 4326 4058 4378
rect 3762 4324 3818 4326
rect 3842 4324 3898 4326
rect 3922 4324 3978 4326
rect 4002 4324 4058 4326
rect 7120 6010 7176 6012
rect 7200 6010 7256 6012
rect 7280 6010 7336 6012
rect 7360 6010 7416 6012
rect 7120 5958 7166 6010
rect 7166 5958 7176 6010
rect 7200 5958 7230 6010
rect 7230 5958 7242 6010
rect 7242 5958 7256 6010
rect 7280 5958 7294 6010
rect 7294 5958 7306 6010
rect 7306 5958 7336 6010
rect 7360 5958 7370 6010
rect 7370 5958 7416 6010
rect 7120 5956 7176 5958
rect 7200 5956 7256 5958
rect 7280 5956 7336 5958
rect 7360 5956 7416 5958
rect 3762 3290 3818 3292
rect 3842 3290 3898 3292
rect 3922 3290 3978 3292
rect 4002 3290 4058 3292
rect 3762 3238 3808 3290
rect 3808 3238 3818 3290
rect 3842 3238 3872 3290
rect 3872 3238 3884 3290
rect 3884 3238 3898 3290
rect 3922 3238 3936 3290
rect 3936 3238 3948 3290
rect 3948 3238 3978 3290
rect 4002 3238 4012 3290
rect 4012 3238 4058 3290
rect 3762 3236 3818 3238
rect 3842 3236 3898 3238
rect 3922 3236 3978 3238
rect 4002 3236 4058 3238
rect 3762 2202 3818 2204
rect 3842 2202 3898 2204
rect 3922 2202 3978 2204
rect 4002 2202 4058 2204
rect 3762 2150 3808 2202
rect 3808 2150 3818 2202
rect 3842 2150 3872 2202
rect 3872 2150 3884 2202
rect 3884 2150 3898 2202
rect 3922 2150 3936 2202
rect 3936 2150 3948 2202
rect 3948 2150 3978 2202
rect 4002 2150 4012 2202
rect 4012 2150 4058 2202
rect 3762 2148 3818 2150
rect 3842 2148 3898 2150
rect 3922 2148 3978 2150
rect 4002 2148 4058 2150
rect 3762 1114 3818 1116
rect 3842 1114 3898 1116
rect 3922 1114 3978 1116
rect 4002 1114 4058 1116
rect 3762 1062 3808 1114
rect 3808 1062 3818 1114
rect 3842 1062 3872 1114
rect 3872 1062 3884 1114
rect 3884 1062 3898 1114
rect 3922 1062 3936 1114
rect 3936 1062 3948 1114
rect 3948 1062 3978 1114
rect 4002 1062 4012 1114
rect 4012 1062 4058 1114
rect 3762 1060 3818 1062
rect 3842 1060 3898 1062
rect 3922 1060 3978 1062
rect 4002 1060 4058 1062
rect 10046 20984 10102 21040
rect 10478 22874 10534 22876
rect 10558 22874 10614 22876
rect 10638 22874 10694 22876
rect 10718 22874 10774 22876
rect 10478 22822 10524 22874
rect 10524 22822 10534 22874
rect 10558 22822 10588 22874
rect 10588 22822 10600 22874
rect 10600 22822 10614 22874
rect 10638 22822 10652 22874
rect 10652 22822 10664 22874
rect 10664 22822 10694 22874
rect 10718 22822 10728 22874
rect 10728 22822 10774 22874
rect 10478 22820 10534 22822
rect 10558 22820 10614 22822
rect 10638 22820 10694 22822
rect 10718 22820 10774 22822
rect 10478 21786 10534 21788
rect 10558 21786 10614 21788
rect 10638 21786 10694 21788
rect 10718 21786 10774 21788
rect 10478 21734 10524 21786
rect 10524 21734 10534 21786
rect 10558 21734 10588 21786
rect 10588 21734 10600 21786
rect 10600 21734 10614 21786
rect 10638 21734 10652 21786
rect 10652 21734 10664 21786
rect 10664 21734 10694 21786
rect 10718 21734 10728 21786
rect 10728 21734 10774 21786
rect 10478 21732 10534 21734
rect 10558 21732 10614 21734
rect 10638 21732 10694 21734
rect 10718 21732 10774 21734
rect 10046 17876 10102 17912
rect 10046 17856 10048 17876
rect 10048 17856 10100 17876
rect 10100 17856 10102 17876
rect 10478 20698 10534 20700
rect 10558 20698 10614 20700
rect 10638 20698 10694 20700
rect 10718 20698 10774 20700
rect 10478 20646 10524 20698
rect 10524 20646 10534 20698
rect 10558 20646 10588 20698
rect 10588 20646 10600 20698
rect 10600 20646 10614 20698
rect 10638 20646 10652 20698
rect 10652 20646 10664 20698
rect 10664 20646 10694 20698
rect 10718 20646 10728 20698
rect 10728 20646 10774 20698
rect 10478 20644 10534 20646
rect 10558 20644 10614 20646
rect 10638 20644 10694 20646
rect 10718 20644 10774 20646
rect 11242 22072 11298 22128
rect 11058 21936 11114 21992
rect 12530 23568 12586 23624
rect 13836 29946 13892 29948
rect 13916 29946 13972 29948
rect 13996 29946 14052 29948
rect 14076 29946 14132 29948
rect 13836 29894 13882 29946
rect 13882 29894 13892 29946
rect 13916 29894 13946 29946
rect 13946 29894 13958 29946
rect 13958 29894 13972 29946
rect 13996 29894 14010 29946
rect 14010 29894 14022 29946
rect 14022 29894 14052 29946
rect 14076 29894 14086 29946
rect 14086 29894 14132 29946
rect 13836 29892 13892 29894
rect 13916 29892 13972 29894
rect 13996 29892 14052 29894
rect 14076 29892 14132 29894
rect 13836 28858 13892 28860
rect 13916 28858 13972 28860
rect 13996 28858 14052 28860
rect 14076 28858 14132 28860
rect 13836 28806 13882 28858
rect 13882 28806 13892 28858
rect 13916 28806 13946 28858
rect 13946 28806 13958 28858
rect 13958 28806 13972 28858
rect 13996 28806 14010 28858
rect 14010 28806 14022 28858
rect 14022 28806 14052 28858
rect 14076 28806 14086 28858
rect 14086 28806 14132 28858
rect 13836 28804 13892 28806
rect 13916 28804 13972 28806
rect 13996 28804 14052 28806
rect 14076 28804 14132 28806
rect 13836 27770 13892 27772
rect 13916 27770 13972 27772
rect 13996 27770 14052 27772
rect 14076 27770 14132 27772
rect 13836 27718 13882 27770
rect 13882 27718 13892 27770
rect 13916 27718 13946 27770
rect 13946 27718 13958 27770
rect 13958 27718 13972 27770
rect 13996 27718 14010 27770
rect 14010 27718 14022 27770
rect 14022 27718 14052 27770
rect 14076 27718 14086 27770
rect 14086 27718 14132 27770
rect 13836 27716 13892 27718
rect 13916 27716 13972 27718
rect 13996 27716 14052 27718
rect 14076 27716 14132 27718
rect 13836 26682 13892 26684
rect 13916 26682 13972 26684
rect 13996 26682 14052 26684
rect 14076 26682 14132 26684
rect 13836 26630 13882 26682
rect 13882 26630 13892 26682
rect 13916 26630 13946 26682
rect 13946 26630 13958 26682
rect 13958 26630 13972 26682
rect 13996 26630 14010 26682
rect 14010 26630 14022 26682
rect 14022 26630 14052 26682
rect 14076 26630 14086 26682
rect 14086 26630 14132 26682
rect 13836 26628 13892 26630
rect 13916 26628 13972 26630
rect 13996 26628 14052 26630
rect 14076 26628 14132 26630
rect 14186 26424 14242 26480
rect 17194 30490 17250 30492
rect 17274 30490 17330 30492
rect 17354 30490 17410 30492
rect 17434 30490 17490 30492
rect 17194 30438 17240 30490
rect 17240 30438 17250 30490
rect 17274 30438 17304 30490
rect 17304 30438 17316 30490
rect 17316 30438 17330 30490
rect 17354 30438 17368 30490
rect 17368 30438 17380 30490
rect 17380 30438 17410 30490
rect 17434 30438 17444 30490
rect 17444 30438 17490 30490
rect 17194 30436 17250 30438
rect 17274 30436 17330 30438
rect 17354 30436 17410 30438
rect 17434 30436 17490 30438
rect 13836 25594 13892 25596
rect 13916 25594 13972 25596
rect 13996 25594 14052 25596
rect 14076 25594 14132 25596
rect 13836 25542 13882 25594
rect 13882 25542 13892 25594
rect 13916 25542 13946 25594
rect 13946 25542 13958 25594
rect 13958 25542 13972 25594
rect 13996 25542 14010 25594
rect 14010 25542 14022 25594
rect 14022 25542 14052 25594
rect 14076 25542 14086 25594
rect 14086 25542 14132 25594
rect 13836 25540 13892 25542
rect 13916 25540 13972 25542
rect 13996 25540 14052 25542
rect 14076 25540 14132 25542
rect 11978 20440 12034 20496
rect 10478 19610 10534 19612
rect 10558 19610 10614 19612
rect 10638 19610 10694 19612
rect 10718 19610 10774 19612
rect 10478 19558 10524 19610
rect 10524 19558 10534 19610
rect 10558 19558 10588 19610
rect 10588 19558 10600 19610
rect 10600 19558 10614 19610
rect 10638 19558 10652 19610
rect 10652 19558 10664 19610
rect 10664 19558 10694 19610
rect 10718 19558 10728 19610
rect 10728 19558 10774 19610
rect 10478 19556 10534 19558
rect 10558 19556 10614 19558
rect 10638 19556 10694 19558
rect 10718 19556 10774 19558
rect 10478 18522 10534 18524
rect 10558 18522 10614 18524
rect 10638 18522 10694 18524
rect 10718 18522 10774 18524
rect 10478 18470 10524 18522
rect 10524 18470 10534 18522
rect 10558 18470 10588 18522
rect 10588 18470 10600 18522
rect 10600 18470 10614 18522
rect 10638 18470 10652 18522
rect 10652 18470 10664 18522
rect 10664 18470 10694 18522
rect 10718 18470 10728 18522
rect 10728 18470 10774 18522
rect 10478 18468 10534 18470
rect 10558 18468 10614 18470
rect 10638 18468 10694 18470
rect 10718 18468 10774 18470
rect 10478 17434 10534 17436
rect 10558 17434 10614 17436
rect 10638 17434 10694 17436
rect 10718 17434 10774 17436
rect 10478 17382 10524 17434
rect 10524 17382 10534 17434
rect 10558 17382 10588 17434
rect 10588 17382 10600 17434
rect 10600 17382 10614 17434
rect 10638 17382 10652 17434
rect 10652 17382 10664 17434
rect 10664 17382 10694 17434
rect 10718 17382 10728 17434
rect 10728 17382 10774 17434
rect 10478 17380 10534 17382
rect 10558 17380 10614 17382
rect 10638 17380 10694 17382
rect 10718 17380 10774 17382
rect 10478 16346 10534 16348
rect 10558 16346 10614 16348
rect 10638 16346 10694 16348
rect 10718 16346 10774 16348
rect 10478 16294 10524 16346
rect 10524 16294 10534 16346
rect 10558 16294 10588 16346
rect 10588 16294 10600 16346
rect 10600 16294 10614 16346
rect 10638 16294 10652 16346
rect 10652 16294 10664 16346
rect 10664 16294 10694 16346
rect 10718 16294 10728 16346
rect 10728 16294 10774 16346
rect 10478 16292 10534 16294
rect 10558 16292 10614 16294
rect 10638 16292 10694 16294
rect 10718 16292 10774 16294
rect 10478 15258 10534 15260
rect 10558 15258 10614 15260
rect 10638 15258 10694 15260
rect 10718 15258 10774 15260
rect 10478 15206 10524 15258
rect 10524 15206 10534 15258
rect 10558 15206 10588 15258
rect 10588 15206 10600 15258
rect 10600 15206 10614 15258
rect 10638 15206 10652 15258
rect 10652 15206 10664 15258
rect 10664 15206 10694 15258
rect 10718 15206 10728 15258
rect 10728 15206 10774 15258
rect 10478 15204 10534 15206
rect 10558 15204 10614 15206
rect 10638 15204 10694 15206
rect 10718 15204 10774 15206
rect 10478 14170 10534 14172
rect 10558 14170 10614 14172
rect 10638 14170 10694 14172
rect 10718 14170 10774 14172
rect 10478 14118 10524 14170
rect 10524 14118 10534 14170
rect 10558 14118 10588 14170
rect 10588 14118 10600 14170
rect 10600 14118 10614 14170
rect 10638 14118 10652 14170
rect 10652 14118 10664 14170
rect 10664 14118 10694 14170
rect 10718 14118 10728 14170
rect 10728 14118 10774 14170
rect 10478 14116 10534 14118
rect 10558 14116 10614 14118
rect 10638 14116 10694 14118
rect 10718 14116 10774 14118
rect 13836 24506 13892 24508
rect 13916 24506 13972 24508
rect 13996 24506 14052 24508
rect 14076 24506 14132 24508
rect 13836 24454 13882 24506
rect 13882 24454 13892 24506
rect 13916 24454 13946 24506
rect 13946 24454 13958 24506
rect 13958 24454 13972 24506
rect 13996 24454 14010 24506
rect 14010 24454 14022 24506
rect 14022 24454 14052 24506
rect 14076 24454 14086 24506
rect 14086 24454 14132 24506
rect 13836 24452 13892 24454
rect 13916 24452 13972 24454
rect 13996 24452 14052 24454
rect 14076 24452 14132 24454
rect 15382 26288 15438 26344
rect 13266 23568 13322 23624
rect 11242 15136 11298 15192
rect 13836 23418 13892 23420
rect 13916 23418 13972 23420
rect 13996 23418 14052 23420
rect 14076 23418 14132 23420
rect 13836 23366 13882 23418
rect 13882 23366 13892 23418
rect 13916 23366 13946 23418
rect 13946 23366 13958 23418
rect 13958 23366 13972 23418
rect 13996 23366 14010 23418
rect 14010 23366 14022 23418
rect 14022 23366 14052 23418
rect 14076 23366 14086 23418
rect 14086 23366 14132 23418
rect 13836 23364 13892 23366
rect 13916 23364 13972 23366
rect 13996 23364 14052 23366
rect 14076 23364 14132 23366
rect 13836 22330 13892 22332
rect 13916 22330 13972 22332
rect 13996 22330 14052 22332
rect 14076 22330 14132 22332
rect 13836 22278 13882 22330
rect 13882 22278 13892 22330
rect 13916 22278 13946 22330
rect 13946 22278 13958 22330
rect 13958 22278 13972 22330
rect 13996 22278 14010 22330
rect 14010 22278 14022 22330
rect 14022 22278 14052 22330
rect 14076 22278 14086 22330
rect 14086 22278 14132 22330
rect 13836 22276 13892 22278
rect 13916 22276 13972 22278
rect 13996 22276 14052 22278
rect 14076 22276 14132 22278
rect 13450 21392 13506 21448
rect 13836 21242 13892 21244
rect 13916 21242 13972 21244
rect 13996 21242 14052 21244
rect 14076 21242 14132 21244
rect 13836 21190 13882 21242
rect 13882 21190 13892 21242
rect 13916 21190 13946 21242
rect 13946 21190 13958 21242
rect 13958 21190 13972 21242
rect 13996 21190 14010 21242
rect 14010 21190 14022 21242
rect 14022 21190 14052 21242
rect 14076 21190 14086 21242
rect 14086 21190 14132 21242
rect 13836 21188 13892 21190
rect 13916 21188 13972 21190
rect 13996 21188 14052 21190
rect 14076 21188 14132 21190
rect 7120 4922 7176 4924
rect 7200 4922 7256 4924
rect 7280 4922 7336 4924
rect 7360 4922 7416 4924
rect 7120 4870 7166 4922
rect 7166 4870 7176 4922
rect 7200 4870 7230 4922
rect 7230 4870 7242 4922
rect 7242 4870 7256 4922
rect 7280 4870 7294 4922
rect 7294 4870 7306 4922
rect 7306 4870 7336 4922
rect 7360 4870 7370 4922
rect 7370 4870 7416 4922
rect 7120 4868 7176 4870
rect 7200 4868 7256 4870
rect 7280 4868 7336 4870
rect 7360 4868 7416 4870
rect 7120 3834 7176 3836
rect 7200 3834 7256 3836
rect 7280 3834 7336 3836
rect 7360 3834 7416 3836
rect 7120 3782 7166 3834
rect 7166 3782 7176 3834
rect 7200 3782 7230 3834
rect 7230 3782 7242 3834
rect 7242 3782 7256 3834
rect 7280 3782 7294 3834
rect 7294 3782 7306 3834
rect 7306 3782 7336 3834
rect 7360 3782 7370 3834
rect 7370 3782 7416 3834
rect 7120 3780 7176 3782
rect 7200 3780 7256 3782
rect 7280 3780 7336 3782
rect 7360 3780 7416 3782
rect 7120 2746 7176 2748
rect 7200 2746 7256 2748
rect 7280 2746 7336 2748
rect 7360 2746 7416 2748
rect 7120 2694 7166 2746
rect 7166 2694 7176 2746
rect 7200 2694 7230 2746
rect 7230 2694 7242 2746
rect 7242 2694 7256 2746
rect 7280 2694 7294 2746
rect 7294 2694 7306 2746
rect 7306 2694 7336 2746
rect 7360 2694 7370 2746
rect 7370 2694 7416 2746
rect 7120 2692 7176 2694
rect 7200 2692 7256 2694
rect 7280 2692 7336 2694
rect 7360 2692 7416 2694
rect 10478 13082 10534 13084
rect 10558 13082 10614 13084
rect 10638 13082 10694 13084
rect 10718 13082 10774 13084
rect 10478 13030 10524 13082
rect 10524 13030 10534 13082
rect 10558 13030 10588 13082
rect 10588 13030 10600 13082
rect 10600 13030 10614 13082
rect 10638 13030 10652 13082
rect 10652 13030 10664 13082
rect 10664 13030 10694 13082
rect 10718 13030 10728 13082
rect 10728 13030 10774 13082
rect 10478 13028 10534 13030
rect 10558 13028 10614 13030
rect 10638 13028 10694 13030
rect 10718 13028 10774 13030
rect 10478 11994 10534 11996
rect 10558 11994 10614 11996
rect 10638 11994 10694 11996
rect 10718 11994 10774 11996
rect 10478 11942 10524 11994
rect 10524 11942 10534 11994
rect 10558 11942 10588 11994
rect 10588 11942 10600 11994
rect 10600 11942 10614 11994
rect 10638 11942 10652 11994
rect 10652 11942 10664 11994
rect 10664 11942 10694 11994
rect 10718 11942 10728 11994
rect 10728 11942 10774 11994
rect 10478 11940 10534 11942
rect 10558 11940 10614 11942
rect 10638 11940 10694 11942
rect 10718 11940 10774 11942
rect 10478 10906 10534 10908
rect 10558 10906 10614 10908
rect 10638 10906 10694 10908
rect 10718 10906 10774 10908
rect 10478 10854 10524 10906
rect 10524 10854 10534 10906
rect 10558 10854 10588 10906
rect 10588 10854 10600 10906
rect 10600 10854 10614 10906
rect 10638 10854 10652 10906
rect 10652 10854 10664 10906
rect 10664 10854 10694 10906
rect 10718 10854 10728 10906
rect 10728 10854 10774 10906
rect 10478 10852 10534 10854
rect 10558 10852 10614 10854
rect 10638 10852 10694 10854
rect 10718 10852 10774 10854
rect 13836 20154 13892 20156
rect 13916 20154 13972 20156
rect 13996 20154 14052 20156
rect 14076 20154 14132 20156
rect 13836 20102 13882 20154
rect 13882 20102 13892 20154
rect 13916 20102 13946 20154
rect 13946 20102 13958 20154
rect 13958 20102 13972 20154
rect 13996 20102 14010 20154
rect 14010 20102 14022 20154
rect 14022 20102 14052 20154
rect 14076 20102 14086 20154
rect 14086 20102 14132 20154
rect 13836 20100 13892 20102
rect 13916 20100 13972 20102
rect 13996 20100 14052 20102
rect 14076 20100 14132 20102
rect 14186 19352 14242 19408
rect 13836 19066 13892 19068
rect 13916 19066 13972 19068
rect 13996 19066 14052 19068
rect 14076 19066 14132 19068
rect 13836 19014 13882 19066
rect 13882 19014 13892 19066
rect 13916 19014 13946 19066
rect 13946 19014 13958 19066
rect 13958 19014 13972 19066
rect 13996 19014 14010 19066
rect 14010 19014 14022 19066
rect 14022 19014 14052 19066
rect 14076 19014 14086 19066
rect 14086 19014 14132 19066
rect 13836 19012 13892 19014
rect 13916 19012 13972 19014
rect 13996 19012 14052 19014
rect 14076 19012 14132 19014
rect 13836 17978 13892 17980
rect 13916 17978 13972 17980
rect 13996 17978 14052 17980
rect 14076 17978 14132 17980
rect 13836 17926 13882 17978
rect 13882 17926 13892 17978
rect 13916 17926 13946 17978
rect 13946 17926 13958 17978
rect 13958 17926 13972 17978
rect 13996 17926 14010 17978
rect 14010 17926 14022 17978
rect 14022 17926 14052 17978
rect 14076 17926 14086 17978
rect 14086 17926 14132 17978
rect 13836 17924 13892 17926
rect 13916 17924 13972 17926
rect 13996 17924 14052 17926
rect 14076 17924 14132 17926
rect 13836 16890 13892 16892
rect 13916 16890 13972 16892
rect 13996 16890 14052 16892
rect 14076 16890 14132 16892
rect 13836 16838 13882 16890
rect 13882 16838 13892 16890
rect 13916 16838 13946 16890
rect 13946 16838 13958 16890
rect 13958 16838 13972 16890
rect 13996 16838 14010 16890
rect 14010 16838 14022 16890
rect 14022 16838 14052 16890
rect 14076 16838 14086 16890
rect 14086 16838 14132 16890
rect 13836 16836 13892 16838
rect 13916 16836 13972 16838
rect 13996 16836 14052 16838
rect 14076 16836 14132 16838
rect 16670 26288 16726 26344
rect 16670 25916 16672 25936
rect 16672 25916 16724 25936
rect 16724 25916 16726 25936
rect 16670 25880 16726 25916
rect 17194 29402 17250 29404
rect 17274 29402 17330 29404
rect 17354 29402 17410 29404
rect 17434 29402 17490 29404
rect 17194 29350 17240 29402
rect 17240 29350 17250 29402
rect 17274 29350 17304 29402
rect 17304 29350 17316 29402
rect 17316 29350 17330 29402
rect 17354 29350 17368 29402
rect 17368 29350 17380 29402
rect 17380 29350 17410 29402
rect 17434 29350 17444 29402
rect 17444 29350 17490 29402
rect 17194 29348 17250 29350
rect 17274 29348 17330 29350
rect 17354 29348 17410 29350
rect 17434 29348 17490 29350
rect 17194 28314 17250 28316
rect 17274 28314 17330 28316
rect 17354 28314 17410 28316
rect 17434 28314 17490 28316
rect 17194 28262 17240 28314
rect 17240 28262 17250 28314
rect 17274 28262 17304 28314
rect 17304 28262 17316 28314
rect 17316 28262 17330 28314
rect 17354 28262 17368 28314
rect 17368 28262 17380 28314
rect 17380 28262 17410 28314
rect 17434 28262 17444 28314
rect 17444 28262 17490 28314
rect 17194 28260 17250 28262
rect 17274 28260 17330 28262
rect 17354 28260 17410 28262
rect 17434 28260 17490 28262
rect 15382 23160 15438 23216
rect 15106 18164 15108 18184
rect 15108 18164 15160 18184
rect 15160 18164 15162 18184
rect 15106 18128 15162 18164
rect 15842 23024 15898 23080
rect 15658 19760 15714 19816
rect 13836 15802 13892 15804
rect 13916 15802 13972 15804
rect 13996 15802 14052 15804
rect 14076 15802 14132 15804
rect 13836 15750 13882 15802
rect 13882 15750 13892 15802
rect 13916 15750 13946 15802
rect 13946 15750 13958 15802
rect 13958 15750 13972 15802
rect 13996 15750 14010 15802
rect 14010 15750 14022 15802
rect 14022 15750 14052 15802
rect 14076 15750 14086 15802
rect 14086 15750 14132 15802
rect 13836 15748 13892 15750
rect 13916 15748 13972 15750
rect 13996 15748 14052 15750
rect 14076 15748 14132 15750
rect 15934 16652 15990 16688
rect 15934 16632 15936 16652
rect 15936 16632 15988 16652
rect 15988 16632 15990 16652
rect 13836 14714 13892 14716
rect 13916 14714 13972 14716
rect 13996 14714 14052 14716
rect 14076 14714 14132 14716
rect 13836 14662 13882 14714
rect 13882 14662 13892 14714
rect 13916 14662 13946 14714
rect 13946 14662 13958 14714
rect 13958 14662 13972 14714
rect 13996 14662 14010 14714
rect 14010 14662 14022 14714
rect 14022 14662 14052 14714
rect 14076 14662 14086 14714
rect 14086 14662 14132 14714
rect 13836 14660 13892 14662
rect 13916 14660 13972 14662
rect 13996 14660 14052 14662
rect 14076 14660 14132 14662
rect 10478 9818 10534 9820
rect 10558 9818 10614 9820
rect 10638 9818 10694 9820
rect 10718 9818 10774 9820
rect 10478 9766 10524 9818
rect 10524 9766 10534 9818
rect 10558 9766 10588 9818
rect 10588 9766 10600 9818
rect 10600 9766 10614 9818
rect 10638 9766 10652 9818
rect 10652 9766 10664 9818
rect 10664 9766 10694 9818
rect 10718 9766 10728 9818
rect 10728 9766 10774 9818
rect 10478 9764 10534 9766
rect 10558 9764 10614 9766
rect 10638 9764 10694 9766
rect 10718 9764 10774 9766
rect 10478 8730 10534 8732
rect 10558 8730 10614 8732
rect 10638 8730 10694 8732
rect 10718 8730 10774 8732
rect 10478 8678 10524 8730
rect 10524 8678 10534 8730
rect 10558 8678 10588 8730
rect 10588 8678 10600 8730
rect 10600 8678 10614 8730
rect 10638 8678 10652 8730
rect 10652 8678 10664 8730
rect 10664 8678 10694 8730
rect 10718 8678 10728 8730
rect 10728 8678 10774 8730
rect 10478 8676 10534 8678
rect 10558 8676 10614 8678
rect 10638 8676 10694 8678
rect 10718 8676 10774 8678
rect 10478 7642 10534 7644
rect 10558 7642 10614 7644
rect 10638 7642 10694 7644
rect 10718 7642 10774 7644
rect 10478 7590 10524 7642
rect 10524 7590 10534 7642
rect 10558 7590 10588 7642
rect 10588 7590 10600 7642
rect 10600 7590 10614 7642
rect 10638 7590 10652 7642
rect 10652 7590 10664 7642
rect 10664 7590 10694 7642
rect 10718 7590 10728 7642
rect 10728 7590 10774 7642
rect 10478 7588 10534 7590
rect 10558 7588 10614 7590
rect 10638 7588 10694 7590
rect 10718 7588 10774 7590
rect 10478 6554 10534 6556
rect 10558 6554 10614 6556
rect 10638 6554 10694 6556
rect 10718 6554 10774 6556
rect 10478 6502 10524 6554
rect 10524 6502 10534 6554
rect 10558 6502 10588 6554
rect 10588 6502 10600 6554
rect 10600 6502 10614 6554
rect 10638 6502 10652 6554
rect 10652 6502 10664 6554
rect 10664 6502 10694 6554
rect 10718 6502 10728 6554
rect 10728 6502 10774 6554
rect 10478 6500 10534 6502
rect 10558 6500 10614 6502
rect 10638 6500 10694 6502
rect 10718 6500 10774 6502
rect 10478 5466 10534 5468
rect 10558 5466 10614 5468
rect 10638 5466 10694 5468
rect 10718 5466 10774 5468
rect 10478 5414 10524 5466
rect 10524 5414 10534 5466
rect 10558 5414 10588 5466
rect 10588 5414 10600 5466
rect 10600 5414 10614 5466
rect 10638 5414 10652 5466
rect 10652 5414 10664 5466
rect 10664 5414 10694 5466
rect 10718 5414 10728 5466
rect 10728 5414 10774 5466
rect 10478 5412 10534 5414
rect 10558 5412 10614 5414
rect 10638 5412 10694 5414
rect 10718 5412 10774 5414
rect 10478 4378 10534 4380
rect 10558 4378 10614 4380
rect 10638 4378 10694 4380
rect 10718 4378 10774 4380
rect 10478 4326 10524 4378
rect 10524 4326 10534 4378
rect 10558 4326 10588 4378
rect 10588 4326 10600 4378
rect 10600 4326 10614 4378
rect 10638 4326 10652 4378
rect 10652 4326 10664 4378
rect 10664 4326 10694 4378
rect 10718 4326 10728 4378
rect 10728 4326 10774 4378
rect 10478 4324 10534 4326
rect 10558 4324 10614 4326
rect 10638 4324 10694 4326
rect 10718 4324 10774 4326
rect 12162 10548 12164 10568
rect 12164 10548 12216 10568
rect 12216 10548 12218 10568
rect 12162 10512 12218 10548
rect 12438 10512 12494 10568
rect 12346 9968 12402 10024
rect 12070 9596 12072 9616
rect 12072 9596 12124 9616
rect 12124 9596 12126 9616
rect 12070 9560 12126 9596
rect 12622 9968 12678 10024
rect 13726 13912 13782 13968
rect 12622 9016 12678 9072
rect 13836 13626 13892 13628
rect 13916 13626 13972 13628
rect 13996 13626 14052 13628
rect 14076 13626 14132 13628
rect 13836 13574 13882 13626
rect 13882 13574 13892 13626
rect 13916 13574 13946 13626
rect 13946 13574 13958 13626
rect 13958 13574 13972 13626
rect 13996 13574 14010 13626
rect 14010 13574 14022 13626
rect 14022 13574 14052 13626
rect 14076 13574 14086 13626
rect 14086 13574 14132 13626
rect 13836 13572 13892 13574
rect 13916 13572 13972 13574
rect 13996 13572 14052 13574
rect 14076 13572 14132 13574
rect 13836 12538 13892 12540
rect 13916 12538 13972 12540
rect 13996 12538 14052 12540
rect 14076 12538 14132 12540
rect 13836 12486 13882 12538
rect 13882 12486 13892 12538
rect 13916 12486 13946 12538
rect 13946 12486 13958 12538
rect 13958 12486 13972 12538
rect 13996 12486 14010 12538
rect 14010 12486 14022 12538
rect 14022 12486 14052 12538
rect 14076 12486 14086 12538
rect 14086 12486 14132 12538
rect 13836 12484 13892 12486
rect 13916 12484 13972 12486
rect 13996 12484 14052 12486
rect 14076 12484 14132 12486
rect 13836 11450 13892 11452
rect 13916 11450 13972 11452
rect 13996 11450 14052 11452
rect 14076 11450 14132 11452
rect 13836 11398 13882 11450
rect 13882 11398 13892 11450
rect 13916 11398 13946 11450
rect 13946 11398 13958 11450
rect 13958 11398 13972 11450
rect 13996 11398 14010 11450
rect 14010 11398 14022 11450
rect 14022 11398 14052 11450
rect 14076 11398 14086 11450
rect 14086 11398 14132 11450
rect 13836 11396 13892 11398
rect 13916 11396 13972 11398
rect 13996 11396 14052 11398
rect 14076 11396 14132 11398
rect 16210 22072 16266 22128
rect 16210 21428 16212 21448
rect 16212 21428 16264 21448
rect 16264 21428 16266 21448
rect 16210 21392 16266 21428
rect 16118 18148 16174 18184
rect 16118 18128 16120 18148
rect 16120 18128 16172 18148
rect 16172 18128 16174 18148
rect 17194 27226 17250 27228
rect 17274 27226 17330 27228
rect 17354 27226 17410 27228
rect 17434 27226 17490 27228
rect 17194 27174 17240 27226
rect 17240 27174 17250 27226
rect 17274 27174 17304 27226
rect 17304 27174 17316 27226
rect 17316 27174 17330 27226
rect 17354 27174 17368 27226
rect 17368 27174 17380 27226
rect 17380 27174 17410 27226
rect 17434 27174 17444 27226
rect 17444 27174 17490 27226
rect 17194 27172 17250 27174
rect 17274 27172 17330 27174
rect 17354 27172 17410 27174
rect 17434 27172 17490 27174
rect 17194 26138 17250 26140
rect 17274 26138 17330 26140
rect 17354 26138 17410 26140
rect 17434 26138 17490 26140
rect 17194 26086 17240 26138
rect 17240 26086 17250 26138
rect 17274 26086 17304 26138
rect 17304 26086 17316 26138
rect 17316 26086 17330 26138
rect 17354 26086 17368 26138
rect 17368 26086 17380 26138
rect 17380 26086 17410 26138
rect 17434 26086 17444 26138
rect 17444 26086 17490 26138
rect 17194 26084 17250 26086
rect 17274 26084 17330 26086
rect 17354 26084 17410 26086
rect 17434 26084 17490 26086
rect 17590 25880 17646 25936
rect 17774 27376 17830 27432
rect 17958 26424 18014 26480
rect 18234 26696 18290 26752
rect 18510 26696 18566 26752
rect 17194 25050 17250 25052
rect 17274 25050 17330 25052
rect 17354 25050 17410 25052
rect 17434 25050 17490 25052
rect 17194 24998 17240 25050
rect 17240 24998 17250 25050
rect 17274 24998 17304 25050
rect 17304 24998 17316 25050
rect 17316 24998 17330 25050
rect 17354 24998 17368 25050
rect 17368 24998 17380 25050
rect 17380 24998 17410 25050
rect 17434 24998 17444 25050
rect 17444 24998 17490 25050
rect 17194 24996 17250 24998
rect 17274 24996 17330 24998
rect 17354 24996 17410 24998
rect 17434 24996 17490 24998
rect 17194 23962 17250 23964
rect 17274 23962 17330 23964
rect 17354 23962 17410 23964
rect 17434 23962 17490 23964
rect 17194 23910 17240 23962
rect 17240 23910 17250 23962
rect 17274 23910 17304 23962
rect 17304 23910 17316 23962
rect 17316 23910 17330 23962
rect 17354 23910 17368 23962
rect 17368 23910 17380 23962
rect 17380 23910 17410 23962
rect 17434 23910 17444 23962
rect 17444 23910 17490 23962
rect 17194 23908 17250 23910
rect 17274 23908 17330 23910
rect 17354 23908 17410 23910
rect 17434 23908 17490 23910
rect 17958 25608 18014 25664
rect 17194 22874 17250 22876
rect 17274 22874 17330 22876
rect 17354 22874 17410 22876
rect 17434 22874 17490 22876
rect 17194 22822 17240 22874
rect 17240 22822 17250 22874
rect 17274 22822 17304 22874
rect 17304 22822 17316 22874
rect 17316 22822 17330 22874
rect 17354 22822 17368 22874
rect 17368 22822 17380 22874
rect 17380 22822 17410 22874
rect 17434 22822 17444 22874
rect 17444 22822 17490 22874
rect 17194 22820 17250 22822
rect 17274 22820 17330 22822
rect 17354 22820 17410 22822
rect 17434 22820 17490 22822
rect 18142 22072 18198 22128
rect 17774 21956 17830 21992
rect 17774 21936 17776 21956
rect 17776 21936 17828 21956
rect 17828 21936 17830 21956
rect 17194 21786 17250 21788
rect 17274 21786 17330 21788
rect 17354 21786 17410 21788
rect 17434 21786 17490 21788
rect 17194 21734 17240 21786
rect 17240 21734 17250 21786
rect 17274 21734 17304 21786
rect 17304 21734 17316 21786
rect 17316 21734 17330 21786
rect 17354 21734 17368 21786
rect 17368 21734 17380 21786
rect 17380 21734 17410 21786
rect 17434 21734 17444 21786
rect 17444 21734 17490 21786
rect 17194 21732 17250 21734
rect 17274 21732 17330 21734
rect 17354 21732 17410 21734
rect 17434 21732 17490 21734
rect 17038 21004 17094 21040
rect 17038 20984 17040 21004
rect 17040 20984 17092 21004
rect 17092 20984 17094 21004
rect 17194 20698 17250 20700
rect 17274 20698 17330 20700
rect 17354 20698 17410 20700
rect 17434 20698 17490 20700
rect 17194 20646 17240 20698
rect 17240 20646 17250 20698
rect 17274 20646 17304 20698
rect 17304 20646 17316 20698
rect 17316 20646 17330 20698
rect 17354 20646 17368 20698
rect 17368 20646 17380 20698
rect 17380 20646 17410 20698
rect 17434 20646 17444 20698
rect 17444 20646 17490 20698
rect 17194 20644 17250 20646
rect 17274 20644 17330 20646
rect 17354 20644 17410 20646
rect 17434 20644 17490 20646
rect 16762 19216 16818 19272
rect 14002 10648 14058 10704
rect 13836 10362 13892 10364
rect 13916 10362 13972 10364
rect 13996 10362 14052 10364
rect 14076 10362 14132 10364
rect 13836 10310 13882 10362
rect 13882 10310 13892 10362
rect 13916 10310 13946 10362
rect 13946 10310 13958 10362
rect 13958 10310 13972 10362
rect 13996 10310 14010 10362
rect 14010 10310 14022 10362
rect 14022 10310 14052 10362
rect 14076 10310 14086 10362
rect 14086 10310 14132 10362
rect 13836 10308 13892 10310
rect 13916 10308 13972 10310
rect 13996 10308 14052 10310
rect 14076 10308 14132 10310
rect 14186 9560 14242 9616
rect 13836 9274 13892 9276
rect 13916 9274 13972 9276
rect 13996 9274 14052 9276
rect 14076 9274 14132 9276
rect 13836 9222 13882 9274
rect 13882 9222 13892 9274
rect 13916 9222 13946 9274
rect 13946 9222 13958 9274
rect 13958 9222 13972 9274
rect 13996 9222 14010 9274
rect 14010 9222 14022 9274
rect 14022 9222 14052 9274
rect 14076 9222 14086 9274
rect 14086 9222 14132 9274
rect 13836 9220 13892 9222
rect 13916 9220 13972 9222
rect 13996 9220 14052 9222
rect 14076 9220 14132 9222
rect 14186 9036 14242 9072
rect 14186 9016 14188 9036
rect 14188 9016 14240 9036
rect 14240 9016 14242 9036
rect 13836 8186 13892 8188
rect 13916 8186 13972 8188
rect 13996 8186 14052 8188
rect 14076 8186 14132 8188
rect 13836 8134 13882 8186
rect 13882 8134 13892 8186
rect 13916 8134 13946 8186
rect 13946 8134 13958 8186
rect 13958 8134 13972 8186
rect 13996 8134 14010 8186
rect 14010 8134 14022 8186
rect 14022 8134 14052 8186
rect 14076 8134 14086 8186
rect 14086 8134 14132 8186
rect 13836 8132 13892 8134
rect 13916 8132 13972 8134
rect 13996 8132 14052 8134
rect 14076 8132 14132 8134
rect 13836 7098 13892 7100
rect 13916 7098 13972 7100
rect 13996 7098 14052 7100
rect 14076 7098 14132 7100
rect 13836 7046 13882 7098
rect 13882 7046 13892 7098
rect 13916 7046 13946 7098
rect 13946 7046 13958 7098
rect 13958 7046 13972 7098
rect 13996 7046 14010 7098
rect 14010 7046 14022 7098
rect 14022 7046 14052 7098
rect 14076 7046 14086 7098
rect 14086 7046 14132 7098
rect 13836 7044 13892 7046
rect 13916 7044 13972 7046
rect 13996 7044 14052 7046
rect 14076 7044 14132 7046
rect 13836 6010 13892 6012
rect 13916 6010 13972 6012
rect 13996 6010 14052 6012
rect 14076 6010 14132 6012
rect 13836 5958 13882 6010
rect 13882 5958 13892 6010
rect 13916 5958 13946 6010
rect 13946 5958 13958 6010
rect 13958 5958 13972 6010
rect 13996 5958 14010 6010
rect 14010 5958 14022 6010
rect 14022 5958 14052 6010
rect 14076 5958 14086 6010
rect 14086 5958 14132 6010
rect 13836 5956 13892 5958
rect 13916 5956 13972 5958
rect 13996 5956 14052 5958
rect 14076 5956 14132 5958
rect 14830 8372 14832 8392
rect 14832 8372 14884 8392
rect 14884 8372 14886 8392
rect 14830 8336 14886 8372
rect 10478 3290 10534 3292
rect 10558 3290 10614 3292
rect 10638 3290 10694 3292
rect 10718 3290 10774 3292
rect 10478 3238 10524 3290
rect 10524 3238 10534 3290
rect 10558 3238 10588 3290
rect 10588 3238 10600 3290
rect 10600 3238 10614 3290
rect 10638 3238 10652 3290
rect 10652 3238 10664 3290
rect 10664 3238 10694 3290
rect 10718 3238 10728 3290
rect 10728 3238 10774 3290
rect 10478 3236 10534 3238
rect 10558 3236 10614 3238
rect 10638 3236 10694 3238
rect 10718 3236 10774 3238
rect 7120 1658 7176 1660
rect 7200 1658 7256 1660
rect 7280 1658 7336 1660
rect 7360 1658 7416 1660
rect 7120 1606 7166 1658
rect 7166 1606 7176 1658
rect 7200 1606 7230 1658
rect 7230 1606 7242 1658
rect 7242 1606 7256 1658
rect 7280 1606 7294 1658
rect 7294 1606 7306 1658
rect 7306 1606 7336 1658
rect 7360 1606 7370 1658
rect 7370 1606 7416 1658
rect 7120 1604 7176 1606
rect 7200 1604 7256 1606
rect 7280 1604 7336 1606
rect 7360 1604 7416 1606
rect 7120 570 7176 572
rect 7200 570 7256 572
rect 7280 570 7336 572
rect 7360 570 7416 572
rect 7120 518 7166 570
rect 7166 518 7176 570
rect 7200 518 7230 570
rect 7230 518 7242 570
rect 7242 518 7256 570
rect 7280 518 7294 570
rect 7294 518 7306 570
rect 7306 518 7336 570
rect 7360 518 7370 570
rect 7370 518 7416 570
rect 7120 516 7176 518
rect 7200 516 7256 518
rect 7280 516 7336 518
rect 7360 516 7416 518
rect 10478 2202 10534 2204
rect 10558 2202 10614 2204
rect 10638 2202 10694 2204
rect 10718 2202 10774 2204
rect 10478 2150 10524 2202
rect 10524 2150 10534 2202
rect 10558 2150 10588 2202
rect 10588 2150 10600 2202
rect 10600 2150 10614 2202
rect 10638 2150 10652 2202
rect 10652 2150 10664 2202
rect 10664 2150 10694 2202
rect 10718 2150 10728 2202
rect 10728 2150 10774 2202
rect 10478 2148 10534 2150
rect 10558 2148 10614 2150
rect 10638 2148 10694 2150
rect 10718 2148 10774 2150
rect 13836 4922 13892 4924
rect 13916 4922 13972 4924
rect 13996 4922 14052 4924
rect 14076 4922 14132 4924
rect 13836 4870 13882 4922
rect 13882 4870 13892 4922
rect 13916 4870 13946 4922
rect 13946 4870 13958 4922
rect 13958 4870 13972 4922
rect 13996 4870 14010 4922
rect 14010 4870 14022 4922
rect 14022 4870 14052 4922
rect 14076 4870 14086 4922
rect 14086 4870 14132 4922
rect 13836 4868 13892 4870
rect 13916 4868 13972 4870
rect 13996 4868 14052 4870
rect 14076 4868 14132 4870
rect 13836 3834 13892 3836
rect 13916 3834 13972 3836
rect 13996 3834 14052 3836
rect 14076 3834 14132 3836
rect 13836 3782 13882 3834
rect 13882 3782 13892 3834
rect 13916 3782 13946 3834
rect 13946 3782 13958 3834
rect 13958 3782 13972 3834
rect 13996 3782 14010 3834
rect 14010 3782 14022 3834
rect 14022 3782 14052 3834
rect 14076 3782 14086 3834
rect 14086 3782 14132 3834
rect 13836 3780 13892 3782
rect 13916 3780 13972 3782
rect 13996 3780 14052 3782
rect 14076 3780 14132 3782
rect 13542 3032 13598 3088
rect 11334 2932 11336 2952
rect 11336 2932 11388 2952
rect 11388 2932 11390 2952
rect 11334 2896 11390 2932
rect 10478 1114 10534 1116
rect 10558 1114 10614 1116
rect 10638 1114 10694 1116
rect 10718 1114 10774 1116
rect 10478 1062 10524 1114
rect 10524 1062 10534 1114
rect 10558 1062 10588 1114
rect 10588 1062 10600 1114
rect 10600 1062 10614 1114
rect 10638 1062 10652 1114
rect 10652 1062 10664 1114
rect 10664 1062 10694 1114
rect 10718 1062 10728 1114
rect 10728 1062 10774 1114
rect 10478 1060 10534 1062
rect 10558 1060 10614 1062
rect 10638 1060 10694 1062
rect 10718 1060 10774 1062
rect 13910 2916 13966 2952
rect 13910 2896 13912 2916
rect 13912 2896 13964 2916
rect 13964 2896 13966 2916
rect 17194 19610 17250 19612
rect 17274 19610 17330 19612
rect 17354 19610 17410 19612
rect 17434 19610 17490 19612
rect 17194 19558 17240 19610
rect 17240 19558 17250 19610
rect 17274 19558 17304 19610
rect 17304 19558 17316 19610
rect 17316 19558 17330 19610
rect 17354 19558 17368 19610
rect 17368 19558 17380 19610
rect 17380 19558 17410 19610
rect 17434 19558 17444 19610
rect 17444 19558 17490 19610
rect 17194 19556 17250 19558
rect 17274 19556 17330 19558
rect 17354 19556 17410 19558
rect 17434 19556 17490 19558
rect 17222 19236 17278 19272
rect 17222 19216 17224 19236
rect 17224 19216 17276 19236
rect 17276 19216 17278 19236
rect 17590 19236 17646 19272
rect 17590 19216 17592 19236
rect 17592 19216 17644 19236
rect 17644 19216 17646 19236
rect 17194 18522 17250 18524
rect 17274 18522 17330 18524
rect 17354 18522 17410 18524
rect 17434 18522 17490 18524
rect 17194 18470 17240 18522
rect 17240 18470 17250 18522
rect 17274 18470 17304 18522
rect 17304 18470 17316 18522
rect 17316 18470 17330 18522
rect 17354 18470 17368 18522
rect 17368 18470 17380 18522
rect 17380 18470 17410 18522
rect 17434 18470 17444 18522
rect 17444 18470 17490 18522
rect 17194 18468 17250 18470
rect 17274 18468 17330 18470
rect 17354 18468 17410 18470
rect 17434 18468 17490 18470
rect 17682 18264 17738 18320
rect 18234 20440 18290 20496
rect 17194 17434 17250 17436
rect 17274 17434 17330 17436
rect 17354 17434 17410 17436
rect 17434 17434 17490 17436
rect 17194 17382 17240 17434
rect 17240 17382 17250 17434
rect 17274 17382 17304 17434
rect 17304 17382 17316 17434
rect 17316 17382 17330 17434
rect 17354 17382 17368 17434
rect 17368 17382 17380 17434
rect 17380 17382 17410 17434
rect 17434 17382 17444 17434
rect 17444 17382 17490 17434
rect 17194 17380 17250 17382
rect 17274 17380 17330 17382
rect 17354 17380 17410 17382
rect 17434 17380 17490 17382
rect 17194 16346 17250 16348
rect 17274 16346 17330 16348
rect 17354 16346 17410 16348
rect 17434 16346 17490 16348
rect 17194 16294 17240 16346
rect 17240 16294 17250 16346
rect 17274 16294 17304 16346
rect 17304 16294 17316 16346
rect 17316 16294 17330 16346
rect 17354 16294 17368 16346
rect 17368 16294 17380 16346
rect 17380 16294 17410 16346
rect 17434 16294 17444 16346
rect 17444 16294 17490 16346
rect 17194 16292 17250 16294
rect 17274 16292 17330 16294
rect 17354 16292 17410 16294
rect 17434 16292 17490 16294
rect 17194 15258 17250 15260
rect 17274 15258 17330 15260
rect 17354 15258 17410 15260
rect 17434 15258 17490 15260
rect 17194 15206 17240 15258
rect 17240 15206 17250 15258
rect 17274 15206 17304 15258
rect 17304 15206 17316 15258
rect 17316 15206 17330 15258
rect 17354 15206 17368 15258
rect 17368 15206 17380 15258
rect 17380 15206 17410 15258
rect 17434 15206 17444 15258
rect 17444 15206 17490 15258
rect 17194 15204 17250 15206
rect 17274 15204 17330 15206
rect 17354 15204 17410 15206
rect 17434 15204 17490 15206
rect 17194 14170 17250 14172
rect 17274 14170 17330 14172
rect 17354 14170 17410 14172
rect 17434 14170 17490 14172
rect 17194 14118 17240 14170
rect 17240 14118 17250 14170
rect 17274 14118 17304 14170
rect 17304 14118 17316 14170
rect 17316 14118 17330 14170
rect 17354 14118 17368 14170
rect 17368 14118 17380 14170
rect 17380 14118 17410 14170
rect 17434 14118 17444 14170
rect 17444 14118 17490 14170
rect 17194 14116 17250 14118
rect 17274 14116 17330 14118
rect 17354 14116 17410 14118
rect 17434 14116 17490 14118
rect 17194 13082 17250 13084
rect 17274 13082 17330 13084
rect 17354 13082 17410 13084
rect 17434 13082 17490 13084
rect 17194 13030 17240 13082
rect 17240 13030 17250 13082
rect 17274 13030 17304 13082
rect 17304 13030 17316 13082
rect 17316 13030 17330 13082
rect 17354 13030 17368 13082
rect 17368 13030 17380 13082
rect 17380 13030 17410 13082
rect 17434 13030 17444 13082
rect 17444 13030 17490 13082
rect 17194 13028 17250 13030
rect 17274 13028 17330 13030
rect 17354 13028 17410 13030
rect 17434 13028 17490 13030
rect 17194 11994 17250 11996
rect 17274 11994 17330 11996
rect 17354 11994 17410 11996
rect 17434 11994 17490 11996
rect 17194 11942 17240 11994
rect 17240 11942 17250 11994
rect 17274 11942 17304 11994
rect 17304 11942 17316 11994
rect 17316 11942 17330 11994
rect 17354 11942 17368 11994
rect 17368 11942 17380 11994
rect 17380 11942 17410 11994
rect 17434 11942 17444 11994
rect 17444 11942 17490 11994
rect 17194 11940 17250 11942
rect 17274 11940 17330 11942
rect 17354 11940 17410 11942
rect 17434 11940 17490 11942
rect 17194 10906 17250 10908
rect 17274 10906 17330 10908
rect 17354 10906 17410 10908
rect 17434 10906 17490 10908
rect 17194 10854 17240 10906
rect 17240 10854 17250 10906
rect 17274 10854 17304 10906
rect 17304 10854 17316 10906
rect 17316 10854 17330 10906
rect 17354 10854 17368 10906
rect 17368 10854 17380 10906
rect 17380 10854 17410 10906
rect 17434 10854 17444 10906
rect 17444 10854 17490 10906
rect 17194 10852 17250 10854
rect 17274 10852 17330 10854
rect 17354 10852 17410 10854
rect 17434 10852 17490 10854
rect 20552 29946 20608 29948
rect 20632 29946 20688 29948
rect 20712 29946 20768 29948
rect 20792 29946 20848 29948
rect 20552 29894 20598 29946
rect 20598 29894 20608 29946
rect 20632 29894 20662 29946
rect 20662 29894 20674 29946
rect 20674 29894 20688 29946
rect 20712 29894 20726 29946
rect 20726 29894 20738 29946
rect 20738 29894 20768 29946
rect 20792 29894 20802 29946
rect 20802 29894 20848 29946
rect 20552 29892 20608 29894
rect 20632 29892 20688 29894
rect 20712 29892 20768 29894
rect 20792 29892 20848 29894
rect 20552 28858 20608 28860
rect 20632 28858 20688 28860
rect 20712 28858 20768 28860
rect 20792 28858 20848 28860
rect 20552 28806 20598 28858
rect 20598 28806 20608 28858
rect 20632 28806 20662 28858
rect 20662 28806 20674 28858
rect 20674 28806 20688 28858
rect 20712 28806 20726 28858
rect 20726 28806 20738 28858
rect 20738 28806 20768 28858
rect 20792 28806 20802 28858
rect 20802 28806 20848 28858
rect 20552 28804 20608 28806
rect 20632 28804 20688 28806
rect 20712 28804 20768 28806
rect 20792 28804 20848 28806
rect 20552 27770 20608 27772
rect 20632 27770 20688 27772
rect 20712 27770 20768 27772
rect 20792 27770 20848 27772
rect 20552 27718 20598 27770
rect 20598 27718 20608 27770
rect 20632 27718 20662 27770
rect 20662 27718 20674 27770
rect 20674 27718 20688 27770
rect 20712 27718 20726 27770
rect 20726 27718 20738 27770
rect 20738 27718 20768 27770
rect 20792 27718 20802 27770
rect 20802 27718 20848 27770
rect 20552 27716 20608 27718
rect 20632 27716 20688 27718
rect 20712 27716 20768 27718
rect 20792 27716 20848 27718
rect 20552 26682 20608 26684
rect 20632 26682 20688 26684
rect 20712 26682 20768 26684
rect 20792 26682 20848 26684
rect 20552 26630 20598 26682
rect 20598 26630 20608 26682
rect 20632 26630 20662 26682
rect 20662 26630 20674 26682
rect 20674 26630 20688 26682
rect 20712 26630 20726 26682
rect 20726 26630 20738 26682
rect 20738 26630 20768 26682
rect 20792 26630 20802 26682
rect 20802 26630 20848 26682
rect 20552 26628 20608 26630
rect 20632 26628 20688 26630
rect 20712 26628 20768 26630
rect 20792 26628 20848 26630
rect 20552 25594 20608 25596
rect 20632 25594 20688 25596
rect 20712 25594 20768 25596
rect 20792 25594 20848 25596
rect 20552 25542 20598 25594
rect 20598 25542 20608 25594
rect 20632 25542 20662 25594
rect 20662 25542 20674 25594
rect 20674 25542 20688 25594
rect 20712 25542 20726 25594
rect 20726 25542 20738 25594
rect 20738 25542 20768 25594
rect 20792 25542 20802 25594
rect 20802 25542 20848 25594
rect 20552 25540 20608 25542
rect 20632 25540 20688 25542
rect 20712 25540 20768 25542
rect 20792 25540 20848 25542
rect 22282 29008 22338 29064
rect 20552 24506 20608 24508
rect 20632 24506 20688 24508
rect 20712 24506 20768 24508
rect 20792 24506 20848 24508
rect 20552 24454 20598 24506
rect 20598 24454 20608 24506
rect 20632 24454 20662 24506
rect 20662 24454 20674 24506
rect 20674 24454 20688 24506
rect 20712 24454 20726 24506
rect 20726 24454 20738 24506
rect 20738 24454 20768 24506
rect 20792 24454 20802 24506
rect 20802 24454 20848 24506
rect 20552 24452 20608 24454
rect 20632 24452 20688 24454
rect 20712 24452 20768 24454
rect 20792 24452 20848 24454
rect 23294 29180 23296 29200
rect 23296 29180 23348 29200
rect 23348 29180 23350 29200
rect 23294 29144 23350 29180
rect 23910 30490 23966 30492
rect 23990 30490 24046 30492
rect 24070 30490 24126 30492
rect 24150 30490 24206 30492
rect 23910 30438 23956 30490
rect 23956 30438 23966 30490
rect 23990 30438 24020 30490
rect 24020 30438 24032 30490
rect 24032 30438 24046 30490
rect 24070 30438 24084 30490
rect 24084 30438 24096 30490
rect 24096 30438 24126 30490
rect 24150 30438 24160 30490
rect 24160 30438 24206 30490
rect 23910 30436 23966 30438
rect 23990 30436 24046 30438
rect 24070 30436 24126 30438
rect 24150 30436 24206 30438
rect 23570 29144 23626 29200
rect 23910 29402 23966 29404
rect 23990 29402 24046 29404
rect 24070 29402 24126 29404
rect 24150 29402 24206 29404
rect 23910 29350 23956 29402
rect 23956 29350 23966 29402
rect 23990 29350 24020 29402
rect 24020 29350 24032 29402
rect 24032 29350 24046 29402
rect 24070 29350 24084 29402
rect 24084 29350 24096 29402
rect 24096 29350 24126 29402
rect 24150 29350 24160 29402
rect 24160 29350 24206 29402
rect 23910 29348 23966 29350
rect 23990 29348 24046 29350
rect 24070 29348 24126 29350
rect 24150 29348 24206 29350
rect 24030 29008 24086 29064
rect 23910 28314 23966 28316
rect 23990 28314 24046 28316
rect 24070 28314 24126 28316
rect 24150 28314 24206 28316
rect 23910 28262 23956 28314
rect 23956 28262 23966 28314
rect 23990 28262 24020 28314
rect 24020 28262 24032 28314
rect 24032 28262 24046 28314
rect 24070 28262 24084 28314
rect 24084 28262 24096 28314
rect 24096 28262 24126 28314
rect 24150 28262 24160 28314
rect 24160 28262 24206 28314
rect 23910 28260 23966 28262
rect 23990 28260 24046 28262
rect 24070 28260 24126 28262
rect 24150 28260 24206 28262
rect 23910 27226 23966 27228
rect 23990 27226 24046 27228
rect 24070 27226 24126 27228
rect 24150 27226 24206 27228
rect 23910 27174 23956 27226
rect 23956 27174 23966 27226
rect 23990 27174 24020 27226
rect 24020 27174 24032 27226
rect 24032 27174 24046 27226
rect 24070 27174 24084 27226
rect 24084 27174 24096 27226
rect 24096 27174 24126 27226
rect 24150 27174 24160 27226
rect 24160 27174 24206 27226
rect 23910 27172 23966 27174
rect 23990 27172 24046 27174
rect 24070 27172 24126 27174
rect 24150 27172 24206 27174
rect 23910 26138 23966 26140
rect 23990 26138 24046 26140
rect 24070 26138 24126 26140
rect 24150 26138 24206 26140
rect 23910 26086 23956 26138
rect 23956 26086 23966 26138
rect 23990 26086 24020 26138
rect 24020 26086 24032 26138
rect 24032 26086 24046 26138
rect 24070 26086 24084 26138
rect 24084 26086 24096 26138
rect 24096 26086 24126 26138
rect 24150 26086 24160 26138
rect 24160 26086 24206 26138
rect 23910 26084 23966 26086
rect 23990 26084 24046 26086
rect 24070 26084 24126 26086
rect 24150 26084 24206 26086
rect 20552 23418 20608 23420
rect 20632 23418 20688 23420
rect 20712 23418 20768 23420
rect 20792 23418 20848 23420
rect 20552 23366 20598 23418
rect 20598 23366 20608 23418
rect 20632 23366 20662 23418
rect 20662 23366 20674 23418
rect 20674 23366 20688 23418
rect 20712 23366 20726 23418
rect 20726 23366 20738 23418
rect 20738 23366 20768 23418
rect 20792 23366 20802 23418
rect 20802 23366 20848 23418
rect 20552 23364 20608 23366
rect 20632 23364 20688 23366
rect 20712 23364 20768 23366
rect 20792 23364 20848 23366
rect 20552 22330 20608 22332
rect 20632 22330 20688 22332
rect 20712 22330 20768 22332
rect 20792 22330 20848 22332
rect 20552 22278 20598 22330
rect 20598 22278 20608 22330
rect 20632 22278 20662 22330
rect 20662 22278 20674 22330
rect 20674 22278 20688 22330
rect 20712 22278 20726 22330
rect 20726 22278 20738 22330
rect 20738 22278 20768 22330
rect 20792 22278 20802 22330
rect 20802 22278 20848 22330
rect 20552 22276 20608 22278
rect 20632 22276 20688 22278
rect 20712 22276 20768 22278
rect 20792 22276 20848 22278
rect 20552 21242 20608 21244
rect 20632 21242 20688 21244
rect 20712 21242 20768 21244
rect 20792 21242 20848 21244
rect 20552 21190 20598 21242
rect 20598 21190 20608 21242
rect 20632 21190 20662 21242
rect 20662 21190 20674 21242
rect 20674 21190 20688 21242
rect 20712 21190 20726 21242
rect 20726 21190 20738 21242
rect 20738 21190 20768 21242
rect 20792 21190 20802 21242
rect 20802 21190 20848 21242
rect 20552 21188 20608 21190
rect 20632 21188 20688 21190
rect 20712 21188 20768 21190
rect 20792 21188 20848 21190
rect 20552 20154 20608 20156
rect 20632 20154 20688 20156
rect 20712 20154 20768 20156
rect 20792 20154 20848 20156
rect 20552 20102 20598 20154
rect 20598 20102 20608 20154
rect 20632 20102 20662 20154
rect 20662 20102 20674 20154
rect 20674 20102 20688 20154
rect 20712 20102 20726 20154
rect 20726 20102 20738 20154
rect 20738 20102 20768 20154
rect 20792 20102 20802 20154
rect 20802 20102 20848 20154
rect 20552 20100 20608 20102
rect 20632 20100 20688 20102
rect 20712 20100 20768 20102
rect 20792 20100 20848 20102
rect 20552 19066 20608 19068
rect 20632 19066 20688 19068
rect 20712 19066 20768 19068
rect 20792 19066 20848 19068
rect 20552 19014 20598 19066
rect 20598 19014 20608 19066
rect 20632 19014 20662 19066
rect 20662 19014 20674 19066
rect 20674 19014 20688 19066
rect 20712 19014 20726 19066
rect 20726 19014 20738 19066
rect 20738 19014 20768 19066
rect 20792 19014 20802 19066
rect 20802 19014 20848 19066
rect 20552 19012 20608 19014
rect 20632 19012 20688 19014
rect 20712 19012 20768 19014
rect 20792 19012 20848 19014
rect 20552 17978 20608 17980
rect 20632 17978 20688 17980
rect 20712 17978 20768 17980
rect 20792 17978 20848 17980
rect 20552 17926 20598 17978
rect 20598 17926 20608 17978
rect 20632 17926 20662 17978
rect 20662 17926 20674 17978
rect 20674 17926 20688 17978
rect 20712 17926 20726 17978
rect 20726 17926 20738 17978
rect 20738 17926 20768 17978
rect 20792 17926 20802 17978
rect 20802 17926 20848 17978
rect 20552 17924 20608 17926
rect 20632 17924 20688 17926
rect 20712 17924 20768 17926
rect 20792 17924 20848 17926
rect 17774 10784 17830 10840
rect 17222 10512 17278 10568
rect 18234 10784 18290 10840
rect 20552 16890 20608 16892
rect 20632 16890 20688 16892
rect 20712 16890 20768 16892
rect 20792 16890 20848 16892
rect 20552 16838 20598 16890
rect 20598 16838 20608 16890
rect 20632 16838 20662 16890
rect 20662 16838 20674 16890
rect 20674 16838 20688 16890
rect 20712 16838 20726 16890
rect 20726 16838 20738 16890
rect 20738 16838 20768 16890
rect 20792 16838 20802 16890
rect 20802 16838 20848 16890
rect 20552 16836 20608 16838
rect 20632 16836 20688 16838
rect 20712 16836 20768 16838
rect 20792 16836 20848 16838
rect 20552 15802 20608 15804
rect 20632 15802 20688 15804
rect 20712 15802 20768 15804
rect 20792 15802 20848 15804
rect 20552 15750 20598 15802
rect 20598 15750 20608 15802
rect 20632 15750 20662 15802
rect 20662 15750 20674 15802
rect 20674 15750 20688 15802
rect 20712 15750 20726 15802
rect 20726 15750 20738 15802
rect 20738 15750 20768 15802
rect 20792 15750 20802 15802
rect 20802 15750 20848 15802
rect 20552 15748 20608 15750
rect 20632 15748 20688 15750
rect 20712 15748 20768 15750
rect 20792 15748 20848 15750
rect 20552 14714 20608 14716
rect 20632 14714 20688 14716
rect 20712 14714 20768 14716
rect 20792 14714 20848 14716
rect 20552 14662 20598 14714
rect 20598 14662 20608 14714
rect 20632 14662 20662 14714
rect 20662 14662 20674 14714
rect 20674 14662 20688 14714
rect 20712 14662 20726 14714
rect 20726 14662 20738 14714
rect 20738 14662 20768 14714
rect 20792 14662 20802 14714
rect 20802 14662 20848 14714
rect 20552 14660 20608 14662
rect 20632 14660 20688 14662
rect 20712 14660 20768 14662
rect 20792 14660 20848 14662
rect 21730 15680 21786 15736
rect 22098 15680 22154 15736
rect 20552 13626 20608 13628
rect 20632 13626 20688 13628
rect 20712 13626 20768 13628
rect 20792 13626 20848 13628
rect 20552 13574 20598 13626
rect 20598 13574 20608 13626
rect 20632 13574 20662 13626
rect 20662 13574 20674 13626
rect 20674 13574 20688 13626
rect 20712 13574 20726 13626
rect 20726 13574 20738 13626
rect 20738 13574 20768 13626
rect 20792 13574 20802 13626
rect 20802 13574 20848 13626
rect 20552 13572 20608 13574
rect 20632 13572 20688 13574
rect 20712 13572 20768 13574
rect 20792 13572 20848 13574
rect 20552 12538 20608 12540
rect 20632 12538 20688 12540
rect 20712 12538 20768 12540
rect 20792 12538 20848 12540
rect 20552 12486 20598 12538
rect 20598 12486 20608 12538
rect 20632 12486 20662 12538
rect 20662 12486 20674 12538
rect 20674 12486 20688 12538
rect 20712 12486 20726 12538
rect 20726 12486 20738 12538
rect 20738 12486 20768 12538
rect 20792 12486 20802 12538
rect 20802 12486 20848 12538
rect 20552 12484 20608 12486
rect 20632 12484 20688 12486
rect 20712 12484 20768 12486
rect 20792 12484 20848 12486
rect 15382 8372 15384 8392
rect 15384 8372 15436 8392
rect 15436 8372 15438 8392
rect 15382 8336 15438 8372
rect 13836 2746 13892 2748
rect 13916 2746 13972 2748
rect 13996 2746 14052 2748
rect 14076 2746 14132 2748
rect 13836 2694 13882 2746
rect 13882 2694 13892 2746
rect 13916 2694 13946 2746
rect 13946 2694 13958 2746
rect 13958 2694 13972 2746
rect 13996 2694 14010 2746
rect 14010 2694 14022 2746
rect 14022 2694 14052 2746
rect 14076 2694 14086 2746
rect 14086 2694 14132 2746
rect 13836 2692 13892 2694
rect 13916 2692 13972 2694
rect 13996 2692 14052 2694
rect 14076 2692 14132 2694
rect 13836 1658 13892 1660
rect 13916 1658 13972 1660
rect 13996 1658 14052 1660
rect 14076 1658 14132 1660
rect 13836 1606 13882 1658
rect 13882 1606 13892 1658
rect 13916 1606 13946 1658
rect 13946 1606 13958 1658
rect 13958 1606 13972 1658
rect 13996 1606 14010 1658
rect 14010 1606 14022 1658
rect 14022 1606 14052 1658
rect 14076 1606 14086 1658
rect 14086 1606 14132 1658
rect 13836 1604 13892 1606
rect 13916 1604 13972 1606
rect 13996 1604 14052 1606
rect 14076 1604 14132 1606
rect 15382 3052 15438 3088
rect 15382 3032 15384 3052
rect 15384 3032 15436 3052
rect 15436 3032 15438 3052
rect 15106 2916 15162 2952
rect 15106 2896 15108 2916
rect 15108 2896 15160 2916
rect 15160 2896 15162 2916
rect 17194 9818 17250 9820
rect 17274 9818 17330 9820
rect 17354 9818 17410 9820
rect 17434 9818 17490 9820
rect 17194 9766 17240 9818
rect 17240 9766 17250 9818
rect 17274 9766 17304 9818
rect 17304 9766 17316 9818
rect 17316 9766 17330 9818
rect 17354 9766 17368 9818
rect 17368 9766 17380 9818
rect 17380 9766 17410 9818
rect 17434 9766 17444 9818
rect 17444 9766 17490 9818
rect 17194 9764 17250 9766
rect 17274 9764 17330 9766
rect 17354 9764 17410 9766
rect 17434 9764 17490 9766
rect 18142 9016 18198 9072
rect 17194 8730 17250 8732
rect 17274 8730 17330 8732
rect 17354 8730 17410 8732
rect 17434 8730 17490 8732
rect 17194 8678 17240 8730
rect 17240 8678 17250 8730
rect 17274 8678 17304 8730
rect 17304 8678 17316 8730
rect 17316 8678 17330 8730
rect 17354 8678 17368 8730
rect 17368 8678 17380 8730
rect 17380 8678 17410 8730
rect 17434 8678 17444 8730
rect 17444 8678 17490 8730
rect 17194 8676 17250 8678
rect 17274 8676 17330 8678
rect 17354 8676 17410 8678
rect 17434 8676 17490 8678
rect 17194 7642 17250 7644
rect 17274 7642 17330 7644
rect 17354 7642 17410 7644
rect 17434 7642 17490 7644
rect 17194 7590 17240 7642
rect 17240 7590 17250 7642
rect 17274 7590 17304 7642
rect 17304 7590 17316 7642
rect 17316 7590 17330 7642
rect 17354 7590 17368 7642
rect 17368 7590 17380 7642
rect 17380 7590 17410 7642
rect 17434 7590 17444 7642
rect 17444 7590 17490 7642
rect 17194 7588 17250 7590
rect 17274 7588 17330 7590
rect 17354 7588 17410 7590
rect 17434 7588 17490 7590
rect 17194 6554 17250 6556
rect 17274 6554 17330 6556
rect 17354 6554 17410 6556
rect 17434 6554 17490 6556
rect 17194 6502 17240 6554
rect 17240 6502 17250 6554
rect 17274 6502 17304 6554
rect 17304 6502 17316 6554
rect 17316 6502 17330 6554
rect 17354 6502 17368 6554
rect 17368 6502 17380 6554
rect 17380 6502 17410 6554
rect 17434 6502 17444 6554
rect 17444 6502 17490 6554
rect 17194 6500 17250 6502
rect 17274 6500 17330 6502
rect 17354 6500 17410 6502
rect 17434 6500 17490 6502
rect 17194 5466 17250 5468
rect 17274 5466 17330 5468
rect 17354 5466 17410 5468
rect 17434 5466 17490 5468
rect 17194 5414 17240 5466
rect 17240 5414 17250 5466
rect 17274 5414 17304 5466
rect 17304 5414 17316 5466
rect 17316 5414 17330 5466
rect 17354 5414 17368 5466
rect 17368 5414 17380 5466
rect 17380 5414 17410 5466
rect 17434 5414 17444 5466
rect 17444 5414 17490 5466
rect 17194 5412 17250 5414
rect 17274 5412 17330 5414
rect 17354 5412 17410 5414
rect 17434 5412 17490 5414
rect 17194 4378 17250 4380
rect 17274 4378 17330 4380
rect 17354 4378 17410 4380
rect 17434 4378 17490 4380
rect 17194 4326 17240 4378
rect 17240 4326 17250 4378
rect 17274 4326 17304 4378
rect 17304 4326 17316 4378
rect 17316 4326 17330 4378
rect 17354 4326 17368 4378
rect 17368 4326 17380 4378
rect 17380 4326 17410 4378
rect 17434 4326 17444 4378
rect 17444 4326 17490 4378
rect 17194 4324 17250 4326
rect 17274 4324 17330 4326
rect 17354 4324 17410 4326
rect 17434 4324 17490 4326
rect 13836 570 13892 572
rect 13916 570 13972 572
rect 13996 570 14052 572
rect 14076 570 14132 572
rect 13836 518 13882 570
rect 13882 518 13892 570
rect 13916 518 13946 570
rect 13946 518 13958 570
rect 13958 518 13972 570
rect 13996 518 14010 570
rect 14010 518 14022 570
rect 14022 518 14052 570
rect 14076 518 14086 570
rect 14086 518 14132 570
rect 13836 516 13892 518
rect 13916 516 13972 518
rect 13996 516 14052 518
rect 14076 516 14132 518
rect 17194 3290 17250 3292
rect 17274 3290 17330 3292
rect 17354 3290 17410 3292
rect 17434 3290 17490 3292
rect 17194 3238 17240 3290
rect 17240 3238 17250 3290
rect 17274 3238 17304 3290
rect 17304 3238 17316 3290
rect 17316 3238 17330 3290
rect 17354 3238 17368 3290
rect 17368 3238 17380 3290
rect 17380 3238 17410 3290
rect 17434 3238 17444 3290
rect 17444 3238 17490 3290
rect 17194 3236 17250 3238
rect 17274 3236 17330 3238
rect 17354 3236 17410 3238
rect 17434 3236 17490 3238
rect 20552 11450 20608 11452
rect 20632 11450 20688 11452
rect 20712 11450 20768 11452
rect 20792 11450 20848 11452
rect 20552 11398 20598 11450
rect 20598 11398 20608 11450
rect 20632 11398 20662 11450
rect 20662 11398 20674 11450
rect 20674 11398 20688 11450
rect 20712 11398 20726 11450
rect 20726 11398 20738 11450
rect 20738 11398 20768 11450
rect 20792 11398 20802 11450
rect 20802 11398 20848 11450
rect 20552 11396 20608 11398
rect 20632 11396 20688 11398
rect 20712 11396 20768 11398
rect 20792 11396 20848 11398
rect 20552 10362 20608 10364
rect 20632 10362 20688 10364
rect 20712 10362 20768 10364
rect 20792 10362 20848 10364
rect 20552 10310 20598 10362
rect 20598 10310 20608 10362
rect 20632 10310 20662 10362
rect 20662 10310 20674 10362
rect 20674 10310 20688 10362
rect 20712 10310 20726 10362
rect 20726 10310 20738 10362
rect 20738 10310 20768 10362
rect 20792 10310 20802 10362
rect 20802 10310 20848 10362
rect 20552 10308 20608 10310
rect 20632 10308 20688 10310
rect 20712 10308 20768 10310
rect 20792 10308 20848 10310
rect 20552 9274 20608 9276
rect 20632 9274 20688 9276
rect 20712 9274 20768 9276
rect 20792 9274 20848 9276
rect 20552 9222 20598 9274
rect 20598 9222 20608 9274
rect 20632 9222 20662 9274
rect 20662 9222 20674 9274
rect 20674 9222 20688 9274
rect 20712 9222 20726 9274
rect 20726 9222 20738 9274
rect 20738 9222 20768 9274
rect 20792 9222 20802 9274
rect 20802 9222 20848 9274
rect 20552 9220 20608 9222
rect 20632 9220 20688 9222
rect 20712 9220 20768 9222
rect 20792 9220 20848 9222
rect 20552 8186 20608 8188
rect 20632 8186 20688 8188
rect 20712 8186 20768 8188
rect 20792 8186 20848 8188
rect 20552 8134 20598 8186
rect 20598 8134 20608 8186
rect 20632 8134 20662 8186
rect 20662 8134 20674 8186
rect 20674 8134 20688 8186
rect 20712 8134 20726 8186
rect 20726 8134 20738 8186
rect 20738 8134 20768 8186
rect 20792 8134 20802 8186
rect 20802 8134 20848 8186
rect 20552 8132 20608 8134
rect 20632 8132 20688 8134
rect 20712 8132 20768 8134
rect 20792 8132 20848 8134
rect 20552 7098 20608 7100
rect 20632 7098 20688 7100
rect 20712 7098 20768 7100
rect 20792 7098 20848 7100
rect 20552 7046 20598 7098
rect 20598 7046 20608 7098
rect 20632 7046 20662 7098
rect 20662 7046 20674 7098
rect 20674 7046 20688 7098
rect 20712 7046 20726 7098
rect 20726 7046 20738 7098
rect 20738 7046 20768 7098
rect 20792 7046 20802 7098
rect 20802 7046 20848 7098
rect 20552 7044 20608 7046
rect 20632 7044 20688 7046
rect 20712 7044 20768 7046
rect 20792 7044 20848 7046
rect 23910 25050 23966 25052
rect 23990 25050 24046 25052
rect 24070 25050 24126 25052
rect 24150 25050 24206 25052
rect 23910 24998 23956 25050
rect 23956 24998 23966 25050
rect 23990 24998 24020 25050
rect 24020 24998 24032 25050
rect 24032 24998 24046 25050
rect 24070 24998 24084 25050
rect 24084 24998 24096 25050
rect 24096 24998 24126 25050
rect 24150 24998 24160 25050
rect 24160 24998 24206 25050
rect 23910 24996 23966 24998
rect 23990 24996 24046 24998
rect 24070 24996 24126 24998
rect 24150 24996 24206 24998
rect 24858 25880 24914 25936
rect 23910 23962 23966 23964
rect 23990 23962 24046 23964
rect 24070 23962 24126 23964
rect 24150 23962 24206 23964
rect 23910 23910 23956 23962
rect 23956 23910 23966 23962
rect 23990 23910 24020 23962
rect 24020 23910 24032 23962
rect 24032 23910 24046 23962
rect 24070 23910 24084 23962
rect 24084 23910 24096 23962
rect 24096 23910 24126 23962
rect 24150 23910 24160 23962
rect 24160 23910 24206 23962
rect 23910 23908 23966 23910
rect 23990 23908 24046 23910
rect 24070 23908 24126 23910
rect 24150 23908 24206 23910
rect 23910 22874 23966 22876
rect 23990 22874 24046 22876
rect 24070 22874 24126 22876
rect 24150 22874 24206 22876
rect 23910 22822 23956 22874
rect 23956 22822 23966 22874
rect 23990 22822 24020 22874
rect 24020 22822 24032 22874
rect 24032 22822 24046 22874
rect 24070 22822 24084 22874
rect 24084 22822 24096 22874
rect 24096 22822 24126 22874
rect 24150 22822 24160 22874
rect 24160 22822 24206 22874
rect 23910 22820 23966 22822
rect 23990 22820 24046 22822
rect 24070 22820 24126 22822
rect 24150 22820 24206 22822
rect 23910 21786 23966 21788
rect 23990 21786 24046 21788
rect 24070 21786 24126 21788
rect 24150 21786 24206 21788
rect 23910 21734 23956 21786
rect 23956 21734 23966 21786
rect 23990 21734 24020 21786
rect 24020 21734 24032 21786
rect 24032 21734 24046 21786
rect 24070 21734 24084 21786
rect 24084 21734 24096 21786
rect 24096 21734 24126 21786
rect 24150 21734 24160 21786
rect 24160 21734 24206 21786
rect 23910 21732 23966 21734
rect 23990 21732 24046 21734
rect 24070 21732 24126 21734
rect 24150 21732 24206 21734
rect 23910 20698 23966 20700
rect 23990 20698 24046 20700
rect 24070 20698 24126 20700
rect 24150 20698 24206 20700
rect 23910 20646 23956 20698
rect 23956 20646 23966 20698
rect 23990 20646 24020 20698
rect 24020 20646 24032 20698
rect 24032 20646 24046 20698
rect 24070 20646 24084 20698
rect 24084 20646 24096 20698
rect 24096 20646 24126 20698
rect 24150 20646 24160 20698
rect 24160 20646 24206 20698
rect 23910 20644 23966 20646
rect 23990 20644 24046 20646
rect 24070 20644 24126 20646
rect 24150 20644 24206 20646
rect 23910 19610 23966 19612
rect 23990 19610 24046 19612
rect 24070 19610 24126 19612
rect 24150 19610 24206 19612
rect 23910 19558 23956 19610
rect 23956 19558 23966 19610
rect 23990 19558 24020 19610
rect 24020 19558 24032 19610
rect 24032 19558 24046 19610
rect 24070 19558 24084 19610
rect 24084 19558 24096 19610
rect 24096 19558 24126 19610
rect 24150 19558 24160 19610
rect 24160 19558 24206 19610
rect 23910 19556 23966 19558
rect 23990 19556 24046 19558
rect 24070 19556 24126 19558
rect 24150 19556 24206 19558
rect 23910 18522 23966 18524
rect 23990 18522 24046 18524
rect 24070 18522 24126 18524
rect 24150 18522 24206 18524
rect 23910 18470 23956 18522
rect 23956 18470 23966 18522
rect 23990 18470 24020 18522
rect 24020 18470 24032 18522
rect 24032 18470 24046 18522
rect 24070 18470 24084 18522
rect 24084 18470 24096 18522
rect 24096 18470 24126 18522
rect 24150 18470 24160 18522
rect 24160 18470 24206 18522
rect 23910 18468 23966 18470
rect 23990 18468 24046 18470
rect 24070 18468 24126 18470
rect 24150 18468 24206 18470
rect 27268 31034 27324 31036
rect 27348 31034 27404 31036
rect 27428 31034 27484 31036
rect 27508 31034 27564 31036
rect 27268 30982 27314 31034
rect 27314 30982 27324 31034
rect 27348 30982 27378 31034
rect 27378 30982 27390 31034
rect 27390 30982 27404 31034
rect 27428 30982 27442 31034
rect 27442 30982 27454 31034
rect 27454 30982 27484 31034
rect 27508 30982 27518 31034
rect 27518 30982 27564 31034
rect 27268 30980 27324 30982
rect 27348 30980 27404 30982
rect 27428 30980 27484 30982
rect 27508 30980 27564 30982
rect 27268 29946 27324 29948
rect 27348 29946 27404 29948
rect 27428 29946 27484 29948
rect 27508 29946 27564 29948
rect 27268 29894 27314 29946
rect 27314 29894 27324 29946
rect 27348 29894 27378 29946
rect 27378 29894 27390 29946
rect 27390 29894 27404 29946
rect 27428 29894 27442 29946
rect 27442 29894 27454 29946
rect 27454 29894 27484 29946
rect 27508 29894 27518 29946
rect 27518 29894 27564 29946
rect 27268 29892 27324 29894
rect 27348 29892 27404 29894
rect 27428 29892 27484 29894
rect 27508 29892 27564 29894
rect 27268 28858 27324 28860
rect 27348 28858 27404 28860
rect 27428 28858 27484 28860
rect 27508 28858 27564 28860
rect 27268 28806 27314 28858
rect 27314 28806 27324 28858
rect 27348 28806 27378 28858
rect 27378 28806 27390 28858
rect 27390 28806 27404 28858
rect 27428 28806 27442 28858
rect 27442 28806 27454 28858
rect 27454 28806 27484 28858
rect 27508 28806 27518 28858
rect 27518 28806 27564 28858
rect 27268 28804 27324 28806
rect 27348 28804 27404 28806
rect 27428 28804 27484 28806
rect 27508 28804 27564 28806
rect 27268 27770 27324 27772
rect 27348 27770 27404 27772
rect 27428 27770 27484 27772
rect 27508 27770 27564 27772
rect 27268 27718 27314 27770
rect 27314 27718 27324 27770
rect 27348 27718 27378 27770
rect 27378 27718 27390 27770
rect 27390 27718 27404 27770
rect 27428 27718 27442 27770
rect 27442 27718 27454 27770
rect 27454 27718 27484 27770
rect 27508 27718 27518 27770
rect 27518 27718 27564 27770
rect 27268 27716 27324 27718
rect 27348 27716 27404 27718
rect 27428 27716 27484 27718
rect 27508 27716 27564 27718
rect 27268 26682 27324 26684
rect 27348 26682 27404 26684
rect 27428 26682 27484 26684
rect 27508 26682 27564 26684
rect 27268 26630 27314 26682
rect 27314 26630 27324 26682
rect 27348 26630 27378 26682
rect 27378 26630 27390 26682
rect 27390 26630 27404 26682
rect 27428 26630 27442 26682
rect 27442 26630 27454 26682
rect 27454 26630 27484 26682
rect 27508 26630 27518 26682
rect 27518 26630 27564 26682
rect 27268 26628 27324 26630
rect 27348 26628 27404 26630
rect 27428 26628 27484 26630
rect 27508 26628 27564 26630
rect 27268 25594 27324 25596
rect 27348 25594 27404 25596
rect 27428 25594 27484 25596
rect 27508 25594 27564 25596
rect 27268 25542 27314 25594
rect 27314 25542 27324 25594
rect 27348 25542 27378 25594
rect 27378 25542 27390 25594
rect 27390 25542 27404 25594
rect 27428 25542 27442 25594
rect 27442 25542 27454 25594
rect 27454 25542 27484 25594
rect 27508 25542 27518 25594
rect 27518 25542 27564 25594
rect 27268 25540 27324 25542
rect 27348 25540 27404 25542
rect 27428 25540 27484 25542
rect 27508 25540 27564 25542
rect 27268 24506 27324 24508
rect 27348 24506 27404 24508
rect 27428 24506 27484 24508
rect 27508 24506 27564 24508
rect 27268 24454 27314 24506
rect 27314 24454 27324 24506
rect 27348 24454 27378 24506
rect 27378 24454 27390 24506
rect 27390 24454 27404 24506
rect 27428 24454 27442 24506
rect 27442 24454 27454 24506
rect 27454 24454 27484 24506
rect 27508 24454 27518 24506
rect 27518 24454 27564 24506
rect 27268 24452 27324 24454
rect 27348 24452 27404 24454
rect 27428 24452 27484 24454
rect 27508 24452 27564 24454
rect 27268 23418 27324 23420
rect 27348 23418 27404 23420
rect 27428 23418 27484 23420
rect 27508 23418 27564 23420
rect 27268 23366 27314 23418
rect 27314 23366 27324 23418
rect 27348 23366 27378 23418
rect 27378 23366 27390 23418
rect 27390 23366 27404 23418
rect 27428 23366 27442 23418
rect 27442 23366 27454 23418
rect 27454 23366 27484 23418
rect 27508 23366 27518 23418
rect 27518 23366 27564 23418
rect 27268 23364 27324 23366
rect 27348 23364 27404 23366
rect 27428 23364 27484 23366
rect 27508 23364 27564 23366
rect 27268 22330 27324 22332
rect 27348 22330 27404 22332
rect 27428 22330 27484 22332
rect 27508 22330 27564 22332
rect 27268 22278 27314 22330
rect 27314 22278 27324 22330
rect 27348 22278 27378 22330
rect 27378 22278 27390 22330
rect 27390 22278 27404 22330
rect 27428 22278 27442 22330
rect 27442 22278 27454 22330
rect 27454 22278 27484 22330
rect 27508 22278 27518 22330
rect 27518 22278 27564 22330
rect 27268 22276 27324 22278
rect 27348 22276 27404 22278
rect 27428 22276 27484 22278
rect 27508 22276 27564 22278
rect 27268 21242 27324 21244
rect 27348 21242 27404 21244
rect 27428 21242 27484 21244
rect 27508 21242 27564 21244
rect 27268 21190 27314 21242
rect 27314 21190 27324 21242
rect 27348 21190 27378 21242
rect 27378 21190 27390 21242
rect 27390 21190 27404 21242
rect 27428 21190 27442 21242
rect 27442 21190 27454 21242
rect 27454 21190 27484 21242
rect 27508 21190 27518 21242
rect 27518 21190 27564 21242
rect 27268 21188 27324 21190
rect 27348 21188 27404 21190
rect 27428 21188 27484 21190
rect 27508 21188 27564 21190
rect 27268 20154 27324 20156
rect 27348 20154 27404 20156
rect 27428 20154 27484 20156
rect 27508 20154 27564 20156
rect 27268 20102 27314 20154
rect 27314 20102 27324 20154
rect 27348 20102 27378 20154
rect 27378 20102 27390 20154
rect 27390 20102 27404 20154
rect 27428 20102 27442 20154
rect 27442 20102 27454 20154
rect 27454 20102 27484 20154
rect 27508 20102 27518 20154
rect 27518 20102 27564 20154
rect 27268 20100 27324 20102
rect 27348 20100 27404 20102
rect 27428 20100 27484 20102
rect 27508 20100 27564 20102
rect 27268 19066 27324 19068
rect 27348 19066 27404 19068
rect 27428 19066 27484 19068
rect 27508 19066 27564 19068
rect 27268 19014 27314 19066
rect 27314 19014 27324 19066
rect 27348 19014 27378 19066
rect 27378 19014 27390 19066
rect 27390 19014 27404 19066
rect 27428 19014 27442 19066
rect 27442 19014 27454 19066
rect 27454 19014 27484 19066
rect 27508 19014 27518 19066
rect 27518 19014 27564 19066
rect 27268 19012 27324 19014
rect 27348 19012 27404 19014
rect 27428 19012 27484 19014
rect 27508 19012 27564 19014
rect 23910 17434 23966 17436
rect 23990 17434 24046 17436
rect 24070 17434 24126 17436
rect 24150 17434 24206 17436
rect 23910 17382 23956 17434
rect 23956 17382 23966 17434
rect 23990 17382 24020 17434
rect 24020 17382 24032 17434
rect 24032 17382 24046 17434
rect 24070 17382 24084 17434
rect 24084 17382 24096 17434
rect 24096 17382 24126 17434
rect 24150 17382 24160 17434
rect 24160 17382 24206 17434
rect 23910 17380 23966 17382
rect 23990 17380 24046 17382
rect 24070 17380 24126 17382
rect 24150 17380 24206 17382
rect 23910 16346 23966 16348
rect 23990 16346 24046 16348
rect 24070 16346 24126 16348
rect 24150 16346 24206 16348
rect 23910 16294 23956 16346
rect 23956 16294 23966 16346
rect 23990 16294 24020 16346
rect 24020 16294 24032 16346
rect 24032 16294 24046 16346
rect 24070 16294 24084 16346
rect 24084 16294 24096 16346
rect 24096 16294 24126 16346
rect 24150 16294 24160 16346
rect 24160 16294 24206 16346
rect 23910 16292 23966 16294
rect 23990 16292 24046 16294
rect 24070 16292 24126 16294
rect 24150 16292 24206 16294
rect 27268 17978 27324 17980
rect 27348 17978 27404 17980
rect 27428 17978 27484 17980
rect 27508 17978 27564 17980
rect 27268 17926 27314 17978
rect 27314 17926 27324 17978
rect 27348 17926 27378 17978
rect 27378 17926 27390 17978
rect 27390 17926 27404 17978
rect 27428 17926 27442 17978
rect 27442 17926 27454 17978
rect 27454 17926 27484 17978
rect 27508 17926 27518 17978
rect 27518 17926 27564 17978
rect 27268 17924 27324 17926
rect 27348 17924 27404 17926
rect 27428 17924 27484 17926
rect 27508 17924 27564 17926
rect 27268 16890 27324 16892
rect 27348 16890 27404 16892
rect 27428 16890 27484 16892
rect 27508 16890 27564 16892
rect 27268 16838 27314 16890
rect 27314 16838 27324 16890
rect 27348 16838 27378 16890
rect 27378 16838 27390 16890
rect 27390 16838 27404 16890
rect 27428 16838 27442 16890
rect 27442 16838 27454 16890
rect 27454 16838 27484 16890
rect 27508 16838 27518 16890
rect 27518 16838 27564 16890
rect 27268 16836 27324 16838
rect 27348 16836 27404 16838
rect 27428 16836 27484 16838
rect 27508 16836 27564 16838
rect 23910 15258 23966 15260
rect 23990 15258 24046 15260
rect 24070 15258 24126 15260
rect 24150 15258 24206 15260
rect 23910 15206 23956 15258
rect 23956 15206 23966 15258
rect 23990 15206 24020 15258
rect 24020 15206 24032 15258
rect 24032 15206 24046 15258
rect 24070 15206 24084 15258
rect 24084 15206 24096 15258
rect 24096 15206 24126 15258
rect 24150 15206 24160 15258
rect 24160 15206 24206 15258
rect 23910 15204 23966 15206
rect 23990 15204 24046 15206
rect 24070 15204 24126 15206
rect 24150 15204 24206 15206
rect 27268 15802 27324 15804
rect 27348 15802 27404 15804
rect 27428 15802 27484 15804
rect 27508 15802 27564 15804
rect 27268 15750 27314 15802
rect 27314 15750 27324 15802
rect 27348 15750 27378 15802
rect 27378 15750 27390 15802
rect 27390 15750 27404 15802
rect 27428 15750 27442 15802
rect 27442 15750 27454 15802
rect 27454 15750 27484 15802
rect 27508 15750 27518 15802
rect 27518 15750 27564 15802
rect 27268 15748 27324 15750
rect 27348 15748 27404 15750
rect 27428 15748 27484 15750
rect 27508 15748 27564 15750
rect 23910 14170 23966 14172
rect 23990 14170 24046 14172
rect 24070 14170 24126 14172
rect 24150 14170 24206 14172
rect 23910 14118 23956 14170
rect 23956 14118 23966 14170
rect 23990 14118 24020 14170
rect 24020 14118 24032 14170
rect 24032 14118 24046 14170
rect 24070 14118 24084 14170
rect 24084 14118 24096 14170
rect 24096 14118 24126 14170
rect 24150 14118 24160 14170
rect 24160 14118 24206 14170
rect 23910 14116 23966 14118
rect 23990 14116 24046 14118
rect 24070 14116 24126 14118
rect 24150 14116 24206 14118
rect 23910 13082 23966 13084
rect 23990 13082 24046 13084
rect 24070 13082 24126 13084
rect 24150 13082 24206 13084
rect 23910 13030 23956 13082
rect 23956 13030 23966 13082
rect 23990 13030 24020 13082
rect 24020 13030 24032 13082
rect 24032 13030 24046 13082
rect 24070 13030 24084 13082
rect 24084 13030 24096 13082
rect 24096 13030 24126 13082
rect 24150 13030 24160 13082
rect 24160 13030 24206 13082
rect 23910 13028 23966 13030
rect 23990 13028 24046 13030
rect 24070 13028 24126 13030
rect 24150 13028 24206 13030
rect 23910 11994 23966 11996
rect 23990 11994 24046 11996
rect 24070 11994 24126 11996
rect 24150 11994 24206 11996
rect 23910 11942 23956 11994
rect 23956 11942 23966 11994
rect 23990 11942 24020 11994
rect 24020 11942 24032 11994
rect 24032 11942 24046 11994
rect 24070 11942 24084 11994
rect 24084 11942 24096 11994
rect 24096 11942 24126 11994
rect 24150 11942 24160 11994
rect 24160 11942 24206 11994
rect 23910 11940 23966 11942
rect 23990 11940 24046 11942
rect 24070 11940 24126 11942
rect 24150 11940 24206 11942
rect 23910 10906 23966 10908
rect 23990 10906 24046 10908
rect 24070 10906 24126 10908
rect 24150 10906 24206 10908
rect 23910 10854 23956 10906
rect 23956 10854 23966 10906
rect 23990 10854 24020 10906
rect 24020 10854 24032 10906
rect 24032 10854 24046 10906
rect 24070 10854 24084 10906
rect 24084 10854 24096 10906
rect 24096 10854 24126 10906
rect 24150 10854 24160 10906
rect 24160 10854 24206 10906
rect 23910 10852 23966 10854
rect 23990 10852 24046 10854
rect 24070 10852 24126 10854
rect 24150 10852 24206 10854
rect 23910 9818 23966 9820
rect 23990 9818 24046 9820
rect 24070 9818 24126 9820
rect 24150 9818 24206 9820
rect 23910 9766 23956 9818
rect 23956 9766 23966 9818
rect 23990 9766 24020 9818
rect 24020 9766 24032 9818
rect 24032 9766 24046 9818
rect 24070 9766 24084 9818
rect 24084 9766 24096 9818
rect 24096 9766 24126 9818
rect 24150 9766 24160 9818
rect 24160 9766 24206 9818
rect 23910 9764 23966 9766
rect 23990 9764 24046 9766
rect 24070 9764 24126 9766
rect 24150 9764 24206 9766
rect 23910 8730 23966 8732
rect 23990 8730 24046 8732
rect 24070 8730 24126 8732
rect 24150 8730 24206 8732
rect 23910 8678 23956 8730
rect 23956 8678 23966 8730
rect 23990 8678 24020 8730
rect 24020 8678 24032 8730
rect 24032 8678 24046 8730
rect 24070 8678 24084 8730
rect 24084 8678 24096 8730
rect 24096 8678 24126 8730
rect 24150 8678 24160 8730
rect 24160 8678 24206 8730
rect 23910 8676 23966 8678
rect 23990 8676 24046 8678
rect 24070 8676 24126 8678
rect 24150 8676 24206 8678
rect 20552 6010 20608 6012
rect 20632 6010 20688 6012
rect 20712 6010 20768 6012
rect 20792 6010 20848 6012
rect 20552 5958 20598 6010
rect 20598 5958 20608 6010
rect 20632 5958 20662 6010
rect 20662 5958 20674 6010
rect 20674 5958 20688 6010
rect 20712 5958 20726 6010
rect 20726 5958 20738 6010
rect 20738 5958 20768 6010
rect 20792 5958 20802 6010
rect 20802 5958 20848 6010
rect 20552 5956 20608 5958
rect 20632 5956 20688 5958
rect 20712 5956 20768 5958
rect 20792 5956 20848 5958
rect 20552 4922 20608 4924
rect 20632 4922 20688 4924
rect 20712 4922 20768 4924
rect 20792 4922 20848 4924
rect 20552 4870 20598 4922
rect 20598 4870 20608 4922
rect 20632 4870 20662 4922
rect 20662 4870 20674 4922
rect 20674 4870 20688 4922
rect 20712 4870 20726 4922
rect 20726 4870 20738 4922
rect 20738 4870 20768 4922
rect 20792 4870 20802 4922
rect 20802 4870 20848 4922
rect 20552 4868 20608 4870
rect 20632 4868 20688 4870
rect 20712 4868 20768 4870
rect 20792 4868 20848 4870
rect 20552 3834 20608 3836
rect 20632 3834 20688 3836
rect 20712 3834 20768 3836
rect 20792 3834 20848 3836
rect 20552 3782 20598 3834
rect 20598 3782 20608 3834
rect 20632 3782 20662 3834
rect 20662 3782 20674 3834
rect 20674 3782 20688 3834
rect 20712 3782 20726 3834
rect 20726 3782 20738 3834
rect 20738 3782 20768 3834
rect 20792 3782 20802 3834
rect 20802 3782 20848 3834
rect 20552 3780 20608 3782
rect 20632 3780 20688 3782
rect 20712 3780 20768 3782
rect 20792 3780 20848 3782
rect 23910 7642 23966 7644
rect 23990 7642 24046 7644
rect 24070 7642 24126 7644
rect 24150 7642 24206 7644
rect 23910 7590 23956 7642
rect 23956 7590 23966 7642
rect 23990 7590 24020 7642
rect 24020 7590 24032 7642
rect 24032 7590 24046 7642
rect 24070 7590 24084 7642
rect 24084 7590 24096 7642
rect 24096 7590 24126 7642
rect 24150 7590 24160 7642
rect 24160 7590 24206 7642
rect 23910 7588 23966 7590
rect 23990 7588 24046 7590
rect 24070 7588 24126 7590
rect 24150 7588 24206 7590
rect 23910 6554 23966 6556
rect 23990 6554 24046 6556
rect 24070 6554 24126 6556
rect 24150 6554 24206 6556
rect 23910 6502 23956 6554
rect 23956 6502 23966 6554
rect 23990 6502 24020 6554
rect 24020 6502 24032 6554
rect 24032 6502 24046 6554
rect 24070 6502 24084 6554
rect 24084 6502 24096 6554
rect 24096 6502 24126 6554
rect 24150 6502 24160 6554
rect 24160 6502 24206 6554
rect 23910 6500 23966 6502
rect 23990 6500 24046 6502
rect 24070 6500 24126 6502
rect 24150 6500 24206 6502
rect 27268 14714 27324 14716
rect 27348 14714 27404 14716
rect 27428 14714 27484 14716
rect 27508 14714 27564 14716
rect 27268 14662 27314 14714
rect 27314 14662 27324 14714
rect 27348 14662 27378 14714
rect 27378 14662 27390 14714
rect 27390 14662 27404 14714
rect 27428 14662 27442 14714
rect 27442 14662 27454 14714
rect 27454 14662 27484 14714
rect 27508 14662 27518 14714
rect 27518 14662 27564 14714
rect 27268 14660 27324 14662
rect 27348 14660 27404 14662
rect 27428 14660 27484 14662
rect 27508 14660 27564 14662
rect 27268 13626 27324 13628
rect 27348 13626 27404 13628
rect 27428 13626 27484 13628
rect 27508 13626 27564 13628
rect 27268 13574 27314 13626
rect 27314 13574 27324 13626
rect 27348 13574 27378 13626
rect 27378 13574 27390 13626
rect 27390 13574 27404 13626
rect 27428 13574 27442 13626
rect 27442 13574 27454 13626
rect 27454 13574 27484 13626
rect 27508 13574 27518 13626
rect 27518 13574 27564 13626
rect 27268 13572 27324 13574
rect 27348 13572 27404 13574
rect 27428 13572 27484 13574
rect 27508 13572 27564 13574
rect 23910 5466 23966 5468
rect 23990 5466 24046 5468
rect 24070 5466 24126 5468
rect 24150 5466 24206 5468
rect 23910 5414 23956 5466
rect 23956 5414 23966 5466
rect 23990 5414 24020 5466
rect 24020 5414 24032 5466
rect 24032 5414 24046 5466
rect 24070 5414 24084 5466
rect 24084 5414 24096 5466
rect 24096 5414 24126 5466
rect 24150 5414 24160 5466
rect 24160 5414 24206 5466
rect 23910 5412 23966 5414
rect 23990 5412 24046 5414
rect 24070 5412 24126 5414
rect 24150 5412 24206 5414
rect 23910 4378 23966 4380
rect 23990 4378 24046 4380
rect 24070 4378 24126 4380
rect 24150 4378 24206 4380
rect 23910 4326 23956 4378
rect 23956 4326 23966 4378
rect 23990 4326 24020 4378
rect 24020 4326 24032 4378
rect 24032 4326 24046 4378
rect 24070 4326 24084 4378
rect 24084 4326 24096 4378
rect 24096 4326 24126 4378
rect 24150 4326 24160 4378
rect 24160 4326 24206 4378
rect 23910 4324 23966 4326
rect 23990 4324 24046 4326
rect 24070 4324 24126 4326
rect 24150 4324 24206 4326
rect 21638 2932 21640 2952
rect 21640 2932 21692 2952
rect 21692 2932 21694 2952
rect 21638 2896 21694 2932
rect 20552 2746 20608 2748
rect 20632 2746 20688 2748
rect 20712 2746 20768 2748
rect 20792 2746 20848 2748
rect 20552 2694 20598 2746
rect 20598 2694 20608 2746
rect 20632 2694 20662 2746
rect 20662 2694 20674 2746
rect 20674 2694 20688 2746
rect 20712 2694 20726 2746
rect 20726 2694 20738 2746
rect 20738 2694 20768 2746
rect 20792 2694 20802 2746
rect 20802 2694 20848 2746
rect 20552 2692 20608 2694
rect 20632 2692 20688 2694
rect 20712 2692 20768 2694
rect 20792 2692 20848 2694
rect 17194 2202 17250 2204
rect 17274 2202 17330 2204
rect 17354 2202 17410 2204
rect 17434 2202 17490 2204
rect 17194 2150 17240 2202
rect 17240 2150 17250 2202
rect 17274 2150 17304 2202
rect 17304 2150 17316 2202
rect 17316 2150 17330 2202
rect 17354 2150 17368 2202
rect 17368 2150 17380 2202
rect 17380 2150 17410 2202
rect 17434 2150 17444 2202
rect 17444 2150 17490 2202
rect 17194 2148 17250 2150
rect 17274 2148 17330 2150
rect 17354 2148 17410 2150
rect 17434 2148 17490 2150
rect 17194 1114 17250 1116
rect 17274 1114 17330 1116
rect 17354 1114 17410 1116
rect 17434 1114 17490 1116
rect 17194 1062 17240 1114
rect 17240 1062 17250 1114
rect 17274 1062 17304 1114
rect 17304 1062 17316 1114
rect 17316 1062 17330 1114
rect 17354 1062 17368 1114
rect 17368 1062 17380 1114
rect 17380 1062 17410 1114
rect 17434 1062 17444 1114
rect 17444 1062 17490 1114
rect 17194 1060 17250 1062
rect 17274 1060 17330 1062
rect 17354 1060 17410 1062
rect 17434 1060 17490 1062
rect 20552 1658 20608 1660
rect 20632 1658 20688 1660
rect 20712 1658 20768 1660
rect 20792 1658 20848 1660
rect 20552 1606 20598 1658
rect 20598 1606 20608 1658
rect 20632 1606 20662 1658
rect 20662 1606 20674 1658
rect 20674 1606 20688 1658
rect 20712 1606 20726 1658
rect 20726 1606 20738 1658
rect 20738 1606 20768 1658
rect 20792 1606 20802 1658
rect 20802 1606 20848 1658
rect 20552 1604 20608 1606
rect 20632 1604 20688 1606
rect 20712 1604 20768 1606
rect 20792 1604 20848 1606
rect 20552 570 20608 572
rect 20632 570 20688 572
rect 20712 570 20768 572
rect 20792 570 20848 572
rect 20552 518 20598 570
rect 20598 518 20608 570
rect 20632 518 20662 570
rect 20662 518 20674 570
rect 20674 518 20688 570
rect 20712 518 20726 570
rect 20726 518 20738 570
rect 20738 518 20768 570
rect 20792 518 20802 570
rect 20802 518 20848 570
rect 20552 516 20608 518
rect 20632 516 20688 518
rect 20712 516 20768 518
rect 20792 516 20848 518
rect 27268 12538 27324 12540
rect 27348 12538 27404 12540
rect 27428 12538 27484 12540
rect 27508 12538 27564 12540
rect 27268 12486 27314 12538
rect 27314 12486 27324 12538
rect 27348 12486 27378 12538
rect 27378 12486 27390 12538
rect 27390 12486 27404 12538
rect 27428 12486 27442 12538
rect 27442 12486 27454 12538
rect 27454 12486 27484 12538
rect 27508 12486 27518 12538
rect 27518 12486 27564 12538
rect 27268 12484 27324 12486
rect 27348 12484 27404 12486
rect 27428 12484 27484 12486
rect 27508 12484 27564 12486
rect 27268 11450 27324 11452
rect 27348 11450 27404 11452
rect 27428 11450 27484 11452
rect 27508 11450 27564 11452
rect 27268 11398 27314 11450
rect 27314 11398 27324 11450
rect 27348 11398 27378 11450
rect 27378 11398 27390 11450
rect 27390 11398 27404 11450
rect 27428 11398 27442 11450
rect 27442 11398 27454 11450
rect 27454 11398 27484 11450
rect 27508 11398 27518 11450
rect 27518 11398 27564 11450
rect 27268 11396 27324 11398
rect 27348 11396 27404 11398
rect 27428 11396 27484 11398
rect 27508 11396 27564 11398
rect 27268 10362 27324 10364
rect 27348 10362 27404 10364
rect 27428 10362 27484 10364
rect 27508 10362 27564 10364
rect 27268 10310 27314 10362
rect 27314 10310 27324 10362
rect 27348 10310 27378 10362
rect 27378 10310 27390 10362
rect 27390 10310 27404 10362
rect 27428 10310 27442 10362
rect 27442 10310 27454 10362
rect 27454 10310 27484 10362
rect 27508 10310 27518 10362
rect 27518 10310 27564 10362
rect 27268 10308 27324 10310
rect 27348 10308 27404 10310
rect 27428 10308 27484 10310
rect 27508 10308 27564 10310
rect 27268 9274 27324 9276
rect 27348 9274 27404 9276
rect 27428 9274 27484 9276
rect 27508 9274 27564 9276
rect 27268 9222 27314 9274
rect 27314 9222 27324 9274
rect 27348 9222 27378 9274
rect 27378 9222 27390 9274
rect 27390 9222 27404 9274
rect 27428 9222 27442 9274
rect 27442 9222 27454 9274
rect 27454 9222 27484 9274
rect 27508 9222 27518 9274
rect 27518 9222 27564 9274
rect 27268 9220 27324 9222
rect 27348 9220 27404 9222
rect 27428 9220 27484 9222
rect 27508 9220 27564 9222
rect 27268 8186 27324 8188
rect 27348 8186 27404 8188
rect 27428 8186 27484 8188
rect 27508 8186 27564 8188
rect 27268 8134 27314 8186
rect 27314 8134 27324 8186
rect 27348 8134 27378 8186
rect 27378 8134 27390 8186
rect 27390 8134 27404 8186
rect 27428 8134 27442 8186
rect 27442 8134 27454 8186
rect 27454 8134 27484 8186
rect 27508 8134 27518 8186
rect 27518 8134 27564 8186
rect 27268 8132 27324 8134
rect 27348 8132 27404 8134
rect 27428 8132 27484 8134
rect 27508 8132 27564 8134
rect 27268 7098 27324 7100
rect 27348 7098 27404 7100
rect 27428 7098 27484 7100
rect 27508 7098 27564 7100
rect 27268 7046 27314 7098
rect 27314 7046 27324 7098
rect 27348 7046 27378 7098
rect 27378 7046 27390 7098
rect 27390 7046 27404 7098
rect 27428 7046 27442 7098
rect 27442 7046 27454 7098
rect 27454 7046 27484 7098
rect 27508 7046 27518 7098
rect 27518 7046 27564 7098
rect 27268 7044 27324 7046
rect 27348 7044 27404 7046
rect 27428 7044 27484 7046
rect 27508 7044 27564 7046
rect 27268 6010 27324 6012
rect 27348 6010 27404 6012
rect 27428 6010 27484 6012
rect 27508 6010 27564 6012
rect 27268 5958 27314 6010
rect 27314 5958 27324 6010
rect 27348 5958 27378 6010
rect 27378 5958 27390 6010
rect 27390 5958 27404 6010
rect 27428 5958 27442 6010
rect 27442 5958 27454 6010
rect 27454 5958 27484 6010
rect 27508 5958 27518 6010
rect 27518 5958 27564 6010
rect 27268 5956 27324 5958
rect 27348 5956 27404 5958
rect 27428 5956 27484 5958
rect 27508 5956 27564 5958
rect 27268 4922 27324 4924
rect 27348 4922 27404 4924
rect 27428 4922 27484 4924
rect 27508 4922 27564 4924
rect 27268 4870 27314 4922
rect 27314 4870 27324 4922
rect 27348 4870 27378 4922
rect 27378 4870 27390 4922
rect 27390 4870 27404 4922
rect 27428 4870 27442 4922
rect 27442 4870 27454 4922
rect 27454 4870 27484 4922
rect 27508 4870 27518 4922
rect 27518 4870 27564 4922
rect 27268 4868 27324 4870
rect 27348 4868 27404 4870
rect 27428 4868 27484 4870
rect 27508 4868 27564 4870
rect 27268 3834 27324 3836
rect 27348 3834 27404 3836
rect 27428 3834 27484 3836
rect 27508 3834 27564 3836
rect 27268 3782 27314 3834
rect 27314 3782 27324 3834
rect 27348 3782 27378 3834
rect 27378 3782 27390 3834
rect 27390 3782 27404 3834
rect 27428 3782 27442 3834
rect 27442 3782 27454 3834
rect 27454 3782 27484 3834
rect 27508 3782 27518 3834
rect 27518 3782 27564 3834
rect 27268 3780 27324 3782
rect 27348 3780 27404 3782
rect 27428 3780 27484 3782
rect 27508 3780 27564 3782
rect 23910 3290 23966 3292
rect 23990 3290 24046 3292
rect 24070 3290 24126 3292
rect 24150 3290 24206 3292
rect 23910 3238 23956 3290
rect 23956 3238 23966 3290
rect 23990 3238 24020 3290
rect 24020 3238 24032 3290
rect 24032 3238 24046 3290
rect 24070 3238 24084 3290
rect 24084 3238 24096 3290
rect 24096 3238 24126 3290
rect 24150 3238 24160 3290
rect 24160 3238 24206 3290
rect 23910 3236 23966 3238
rect 23990 3236 24046 3238
rect 24070 3236 24126 3238
rect 24150 3236 24206 3238
rect 23110 2916 23166 2952
rect 23110 2896 23112 2916
rect 23112 2896 23164 2916
rect 23164 2896 23166 2916
rect 23910 2202 23966 2204
rect 23990 2202 24046 2204
rect 24070 2202 24126 2204
rect 24150 2202 24206 2204
rect 23910 2150 23956 2202
rect 23956 2150 23966 2202
rect 23990 2150 24020 2202
rect 24020 2150 24032 2202
rect 24032 2150 24046 2202
rect 24070 2150 24084 2202
rect 24084 2150 24096 2202
rect 24096 2150 24126 2202
rect 24150 2150 24160 2202
rect 24160 2150 24206 2202
rect 23910 2148 23966 2150
rect 23990 2148 24046 2150
rect 24070 2148 24126 2150
rect 24150 2148 24206 2150
rect 23910 1114 23966 1116
rect 23990 1114 24046 1116
rect 24070 1114 24126 1116
rect 24150 1114 24206 1116
rect 23910 1062 23956 1114
rect 23956 1062 23966 1114
rect 23990 1062 24020 1114
rect 24020 1062 24032 1114
rect 24032 1062 24046 1114
rect 24070 1062 24084 1114
rect 24084 1062 24096 1114
rect 24096 1062 24126 1114
rect 24150 1062 24160 1114
rect 24160 1062 24206 1114
rect 23910 1060 23966 1062
rect 23990 1060 24046 1062
rect 24070 1060 24126 1062
rect 24150 1060 24206 1062
rect 27268 2746 27324 2748
rect 27348 2746 27404 2748
rect 27428 2746 27484 2748
rect 27508 2746 27564 2748
rect 27268 2694 27314 2746
rect 27314 2694 27324 2746
rect 27348 2694 27378 2746
rect 27378 2694 27390 2746
rect 27390 2694 27404 2746
rect 27428 2694 27442 2746
rect 27442 2694 27454 2746
rect 27454 2694 27484 2746
rect 27508 2694 27518 2746
rect 27518 2694 27564 2746
rect 27268 2692 27324 2694
rect 27348 2692 27404 2694
rect 27428 2692 27484 2694
rect 27508 2692 27564 2694
rect 27268 1658 27324 1660
rect 27348 1658 27404 1660
rect 27428 1658 27484 1660
rect 27508 1658 27564 1660
rect 27268 1606 27314 1658
rect 27314 1606 27324 1658
rect 27348 1606 27378 1658
rect 27378 1606 27390 1658
rect 27390 1606 27404 1658
rect 27428 1606 27442 1658
rect 27442 1606 27454 1658
rect 27454 1606 27484 1658
rect 27508 1606 27518 1658
rect 27518 1606 27564 1658
rect 27268 1604 27324 1606
rect 27348 1604 27404 1606
rect 27428 1604 27484 1606
rect 27508 1604 27564 1606
rect 27268 570 27324 572
rect 27348 570 27404 572
rect 27428 570 27484 572
rect 27508 570 27564 572
rect 27268 518 27314 570
rect 27314 518 27324 570
rect 27348 518 27378 570
rect 27378 518 27390 570
rect 27390 518 27404 570
rect 27428 518 27442 570
rect 27442 518 27454 570
rect 27454 518 27484 570
rect 27508 518 27518 570
rect 27518 518 27564 570
rect 27268 516 27324 518
rect 27348 516 27404 518
rect 27428 516 27484 518
rect 27508 516 27564 518
<< metal3 >>
rect 7110 31040 7426 31041
rect 7110 30976 7116 31040
rect 7180 30976 7196 31040
rect 7260 30976 7276 31040
rect 7340 30976 7356 31040
rect 7420 30976 7426 31040
rect 7110 30975 7426 30976
rect 13826 31040 14142 31041
rect 13826 30976 13832 31040
rect 13896 30976 13912 31040
rect 13976 30976 13992 31040
rect 14056 30976 14072 31040
rect 14136 30976 14142 31040
rect 13826 30975 14142 30976
rect 20542 31040 20858 31041
rect 20542 30976 20548 31040
rect 20612 30976 20628 31040
rect 20692 30976 20708 31040
rect 20772 30976 20788 31040
rect 20852 30976 20858 31040
rect 20542 30975 20858 30976
rect 27258 31040 27574 31041
rect 27258 30976 27264 31040
rect 27328 30976 27344 31040
rect 27408 30976 27424 31040
rect 27488 30976 27504 31040
rect 27568 30976 27574 31040
rect 27258 30975 27574 30976
rect 17677 30834 17743 30837
rect 19057 30834 19123 30837
rect 17677 30832 19123 30834
rect 17677 30776 17682 30832
rect 17738 30776 19062 30832
rect 19118 30776 19123 30832
rect 17677 30774 19123 30776
rect 17677 30771 17743 30774
rect 19057 30771 19123 30774
rect 3752 30496 4068 30497
rect 3752 30432 3758 30496
rect 3822 30432 3838 30496
rect 3902 30432 3918 30496
rect 3982 30432 3998 30496
rect 4062 30432 4068 30496
rect 3752 30431 4068 30432
rect 10468 30496 10784 30497
rect 10468 30432 10474 30496
rect 10538 30432 10554 30496
rect 10618 30432 10634 30496
rect 10698 30432 10714 30496
rect 10778 30432 10784 30496
rect 10468 30431 10784 30432
rect 17184 30496 17500 30497
rect 17184 30432 17190 30496
rect 17254 30432 17270 30496
rect 17334 30432 17350 30496
rect 17414 30432 17430 30496
rect 17494 30432 17500 30496
rect 17184 30431 17500 30432
rect 23900 30496 24216 30497
rect 23900 30432 23906 30496
rect 23970 30432 23986 30496
rect 24050 30432 24066 30496
rect 24130 30432 24146 30496
rect 24210 30432 24216 30496
rect 23900 30431 24216 30432
rect 7110 29952 7426 29953
rect 7110 29888 7116 29952
rect 7180 29888 7196 29952
rect 7260 29888 7276 29952
rect 7340 29888 7356 29952
rect 7420 29888 7426 29952
rect 7110 29887 7426 29888
rect 13826 29952 14142 29953
rect 13826 29888 13832 29952
rect 13896 29888 13912 29952
rect 13976 29888 13992 29952
rect 14056 29888 14072 29952
rect 14136 29888 14142 29952
rect 13826 29887 14142 29888
rect 20542 29952 20858 29953
rect 20542 29888 20548 29952
rect 20612 29888 20628 29952
rect 20692 29888 20708 29952
rect 20772 29888 20788 29952
rect 20852 29888 20858 29952
rect 20542 29887 20858 29888
rect 27258 29952 27574 29953
rect 27258 29888 27264 29952
rect 27328 29888 27344 29952
rect 27408 29888 27424 29952
rect 27488 29888 27504 29952
rect 27568 29888 27574 29952
rect 27258 29887 27574 29888
rect 3752 29408 4068 29409
rect 3752 29344 3758 29408
rect 3822 29344 3838 29408
rect 3902 29344 3918 29408
rect 3982 29344 3998 29408
rect 4062 29344 4068 29408
rect 3752 29343 4068 29344
rect 10468 29408 10784 29409
rect 10468 29344 10474 29408
rect 10538 29344 10554 29408
rect 10618 29344 10634 29408
rect 10698 29344 10714 29408
rect 10778 29344 10784 29408
rect 10468 29343 10784 29344
rect 17184 29408 17500 29409
rect 17184 29344 17190 29408
rect 17254 29344 17270 29408
rect 17334 29344 17350 29408
rect 17414 29344 17430 29408
rect 17494 29344 17500 29408
rect 17184 29343 17500 29344
rect 23900 29408 24216 29409
rect 23900 29344 23906 29408
rect 23970 29344 23986 29408
rect 24050 29344 24066 29408
rect 24130 29344 24146 29408
rect 24210 29344 24216 29408
rect 23900 29343 24216 29344
rect 23289 29202 23355 29205
rect 23565 29202 23631 29205
rect 23289 29200 23631 29202
rect 23289 29144 23294 29200
rect 23350 29144 23570 29200
rect 23626 29144 23631 29200
rect 23289 29142 23631 29144
rect 23289 29139 23355 29142
rect 23565 29139 23631 29142
rect 22277 29066 22343 29069
rect 24025 29066 24091 29069
rect 22277 29064 24091 29066
rect 22277 29008 22282 29064
rect 22338 29008 24030 29064
rect 24086 29008 24091 29064
rect 22277 29006 24091 29008
rect 22277 29003 22343 29006
rect 24025 29003 24091 29006
rect 7110 28864 7426 28865
rect 7110 28800 7116 28864
rect 7180 28800 7196 28864
rect 7260 28800 7276 28864
rect 7340 28800 7356 28864
rect 7420 28800 7426 28864
rect 7110 28799 7426 28800
rect 13826 28864 14142 28865
rect 13826 28800 13832 28864
rect 13896 28800 13912 28864
rect 13976 28800 13992 28864
rect 14056 28800 14072 28864
rect 14136 28800 14142 28864
rect 13826 28799 14142 28800
rect 20542 28864 20858 28865
rect 20542 28800 20548 28864
rect 20612 28800 20628 28864
rect 20692 28800 20708 28864
rect 20772 28800 20788 28864
rect 20852 28800 20858 28864
rect 20542 28799 20858 28800
rect 27258 28864 27574 28865
rect 27258 28800 27264 28864
rect 27328 28800 27344 28864
rect 27408 28800 27424 28864
rect 27488 28800 27504 28864
rect 27568 28800 27574 28864
rect 27258 28799 27574 28800
rect 3752 28320 4068 28321
rect 3752 28256 3758 28320
rect 3822 28256 3838 28320
rect 3902 28256 3918 28320
rect 3982 28256 3998 28320
rect 4062 28256 4068 28320
rect 3752 28255 4068 28256
rect 10468 28320 10784 28321
rect 10468 28256 10474 28320
rect 10538 28256 10554 28320
rect 10618 28256 10634 28320
rect 10698 28256 10714 28320
rect 10778 28256 10784 28320
rect 10468 28255 10784 28256
rect 17184 28320 17500 28321
rect 17184 28256 17190 28320
rect 17254 28256 17270 28320
rect 17334 28256 17350 28320
rect 17414 28256 17430 28320
rect 17494 28256 17500 28320
rect 17184 28255 17500 28256
rect 23900 28320 24216 28321
rect 23900 28256 23906 28320
rect 23970 28256 23986 28320
rect 24050 28256 24066 28320
rect 24130 28256 24146 28320
rect 24210 28256 24216 28320
rect 23900 28255 24216 28256
rect 7110 27776 7426 27777
rect 7110 27712 7116 27776
rect 7180 27712 7196 27776
rect 7260 27712 7276 27776
rect 7340 27712 7356 27776
rect 7420 27712 7426 27776
rect 7110 27711 7426 27712
rect 13826 27776 14142 27777
rect 13826 27712 13832 27776
rect 13896 27712 13912 27776
rect 13976 27712 13992 27776
rect 14056 27712 14072 27776
rect 14136 27712 14142 27776
rect 13826 27711 14142 27712
rect 20542 27776 20858 27777
rect 20542 27712 20548 27776
rect 20612 27712 20628 27776
rect 20692 27712 20708 27776
rect 20772 27712 20788 27776
rect 20852 27712 20858 27776
rect 20542 27711 20858 27712
rect 27258 27776 27574 27777
rect 27258 27712 27264 27776
rect 27328 27712 27344 27776
rect 27408 27712 27424 27776
rect 27488 27712 27504 27776
rect 27568 27712 27574 27776
rect 27258 27711 27574 27712
rect 17769 27436 17835 27437
rect 17718 27372 17724 27436
rect 17788 27434 17835 27436
rect 17788 27432 17880 27434
rect 17830 27376 17880 27432
rect 17788 27374 17880 27376
rect 17788 27372 17835 27374
rect 17769 27371 17835 27372
rect 3752 27232 4068 27233
rect 3752 27168 3758 27232
rect 3822 27168 3838 27232
rect 3902 27168 3918 27232
rect 3982 27168 3998 27232
rect 4062 27168 4068 27232
rect 3752 27167 4068 27168
rect 10468 27232 10784 27233
rect 10468 27168 10474 27232
rect 10538 27168 10554 27232
rect 10618 27168 10634 27232
rect 10698 27168 10714 27232
rect 10778 27168 10784 27232
rect 10468 27167 10784 27168
rect 17184 27232 17500 27233
rect 17184 27168 17190 27232
rect 17254 27168 17270 27232
rect 17334 27168 17350 27232
rect 17414 27168 17430 27232
rect 17494 27168 17500 27232
rect 17184 27167 17500 27168
rect 23900 27232 24216 27233
rect 23900 27168 23906 27232
rect 23970 27168 23986 27232
rect 24050 27168 24066 27232
rect 24130 27168 24146 27232
rect 24210 27168 24216 27232
rect 23900 27167 24216 27168
rect 18229 26754 18295 26757
rect 18505 26754 18571 26757
rect 18229 26752 18571 26754
rect 18229 26696 18234 26752
rect 18290 26696 18510 26752
rect 18566 26696 18571 26752
rect 18229 26694 18571 26696
rect 18229 26691 18295 26694
rect 18505 26691 18571 26694
rect 7110 26688 7426 26689
rect 7110 26624 7116 26688
rect 7180 26624 7196 26688
rect 7260 26624 7276 26688
rect 7340 26624 7356 26688
rect 7420 26624 7426 26688
rect 7110 26623 7426 26624
rect 13826 26688 14142 26689
rect 13826 26624 13832 26688
rect 13896 26624 13912 26688
rect 13976 26624 13992 26688
rect 14056 26624 14072 26688
rect 14136 26624 14142 26688
rect 13826 26623 14142 26624
rect 20542 26688 20858 26689
rect 20542 26624 20548 26688
rect 20612 26624 20628 26688
rect 20692 26624 20708 26688
rect 20772 26624 20788 26688
rect 20852 26624 20858 26688
rect 20542 26623 20858 26624
rect 27258 26688 27574 26689
rect 27258 26624 27264 26688
rect 27328 26624 27344 26688
rect 27408 26624 27424 26688
rect 27488 26624 27504 26688
rect 27568 26624 27574 26688
rect 27258 26623 27574 26624
rect 14181 26482 14247 26485
rect 17953 26482 18019 26485
rect 14181 26480 18019 26482
rect 14181 26424 14186 26480
rect 14242 26424 17958 26480
rect 18014 26424 18019 26480
rect 14181 26422 18019 26424
rect 14181 26419 14247 26422
rect 17953 26419 18019 26422
rect 5901 26346 5967 26349
rect 6729 26346 6795 26349
rect 15377 26346 15443 26349
rect 16665 26346 16731 26349
rect 5901 26344 16731 26346
rect 5901 26288 5906 26344
rect 5962 26288 6734 26344
rect 6790 26288 15382 26344
rect 15438 26288 16670 26344
rect 16726 26288 16731 26344
rect 5901 26286 16731 26288
rect 5901 26283 5967 26286
rect 6729 26283 6795 26286
rect 15377 26283 15443 26286
rect 16665 26283 16731 26286
rect 3752 26144 4068 26145
rect 3752 26080 3758 26144
rect 3822 26080 3838 26144
rect 3902 26080 3918 26144
rect 3982 26080 3998 26144
rect 4062 26080 4068 26144
rect 3752 26079 4068 26080
rect 10468 26144 10784 26145
rect 10468 26080 10474 26144
rect 10538 26080 10554 26144
rect 10618 26080 10634 26144
rect 10698 26080 10714 26144
rect 10778 26080 10784 26144
rect 10468 26079 10784 26080
rect 17184 26144 17500 26145
rect 17184 26080 17190 26144
rect 17254 26080 17270 26144
rect 17334 26080 17350 26144
rect 17414 26080 17430 26144
rect 17494 26080 17500 26144
rect 17184 26079 17500 26080
rect 23900 26144 24216 26145
rect 23900 26080 23906 26144
rect 23970 26080 23986 26144
rect 24050 26080 24066 26144
rect 24130 26080 24146 26144
rect 24210 26080 24216 26144
rect 23900 26079 24216 26080
rect 16665 25940 16731 25941
rect 16614 25938 16620 25940
rect 16574 25878 16620 25938
rect 16684 25938 16731 25940
rect 17585 25938 17651 25941
rect 16684 25936 17651 25938
rect 16726 25880 17590 25936
rect 17646 25880 17651 25936
rect 16614 25876 16620 25878
rect 16684 25878 17651 25880
rect 16684 25876 16731 25878
rect 16665 25875 16731 25876
rect 17585 25875 17651 25878
rect 17718 25876 17724 25940
rect 17788 25938 17794 25940
rect 24853 25938 24919 25941
rect 17788 25936 24919 25938
rect 17788 25880 24858 25936
rect 24914 25880 24919 25936
rect 17788 25878 24919 25880
rect 17788 25876 17794 25878
rect 24853 25875 24919 25878
rect 17953 25668 18019 25669
rect 17902 25604 17908 25668
rect 17972 25666 18019 25668
rect 17972 25664 18064 25666
rect 18014 25608 18064 25664
rect 17972 25606 18064 25608
rect 17972 25604 18019 25606
rect 17953 25603 18019 25604
rect 7110 25600 7426 25601
rect 7110 25536 7116 25600
rect 7180 25536 7196 25600
rect 7260 25536 7276 25600
rect 7340 25536 7356 25600
rect 7420 25536 7426 25600
rect 7110 25535 7426 25536
rect 13826 25600 14142 25601
rect 13826 25536 13832 25600
rect 13896 25536 13912 25600
rect 13976 25536 13992 25600
rect 14056 25536 14072 25600
rect 14136 25536 14142 25600
rect 13826 25535 14142 25536
rect 20542 25600 20858 25601
rect 20542 25536 20548 25600
rect 20612 25536 20628 25600
rect 20692 25536 20708 25600
rect 20772 25536 20788 25600
rect 20852 25536 20858 25600
rect 20542 25535 20858 25536
rect 27258 25600 27574 25601
rect 27258 25536 27264 25600
rect 27328 25536 27344 25600
rect 27408 25536 27424 25600
rect 27488 25536 27504 25600
rect 27568 25536 27574 25600
rect 27258 25535 27574 25536
rect 3752 25056 4068 25057
rect 3752 24992 3758 25056
rect 3822 24992 3838 25056
rect 3902 24992 3918 25056
rect 3982 24992 3998 25056
rect 4062 24992 4068 25056
rect 3752 24991 4068 24992
rect 10468 25056 10784 25057
rect 10468 24992 10474 25056
rect 10538 24992 10554 25056
rect 10618 24992 10634 25056
rect 10698 24992 10714 25056
rect 10778 24992 10784 25056
rect 10468 24991 10784 24992
rect 17184 25056 17500 25057
rect 17184 24992 17190 25056
rect 17254 24992 17270 25056
rect 17334 24992 17350 25056
rect 17414 24992 17430 25056
rect 17494 24992 17500 25056
rect 17184 24991 17500 24992
rect 23900 25056 24216 25057
rect 23900 24992 23906 25056
rect 23970 24992 23986 25056
rect 24050 24992 24066 25056
rect 24130 24992 24146 25056
rect 24210 24992 24216 25056
rect 23900 24991 24216 24992
rect 7110 24512 7426 24513
rect 7110 24448 7116 24512
rect 7180 24448 7196 24512
rect 7260 24448 7276 24512
rect 7340 24448 7356 24512
rect 7420 24448 7426 24512
rect 7110 24447 7426 24448
rect 13826 24512 14142 24513
rect 13826 24448 13832 24512
rect 13896 24448 13912 24512
rect 13976 24448 13992 24512
rect 14056 24448 14072 24512
rect 14136 24448 14142 24512
rect 13826 24447 14142 24448
rect 20542 24512 20858 24513
rect 20542 24448 20548 24512
rect 20612 24448 20628 24512
rect 20692 24448 20708 24512
rect 20772 24448 20788 24512
rect 20852 24448 20858 24512
rect 20542 24447 20858 24448
rect 27258 24512 27574 24513
rect 27258 24448 27264 24512
rect 27328 24448 27344 24512
rect 27408 24448 27424 24512
rect 27488 24448 27504 24512
rect 27568 24448 27574 24512
rect 27258 24447 27574 24448
rect 3752 23968 4068 23969
rect 3752 23904 3758 23968
rect 3822 23904 3838 23968
rect 3902 23904 3918 23968
rect 3982 23904 3998 23968
rect 4062 23904 4068 23968
rect 3752 23903 4068 23904
rect 10468 23968 10784 23969
rect 10468 23904 10474 23968
rect 10538 23904 10554 23968
rect 10618 23904 10634 23968
rect 10698 23904 10714 23968
rect 10778 23904 10784 23968
rect 10468 23903 10784 23904
rect 17184 23968 17500 23969
rect 17184 23904 17190 23968
rect 17254 23904 17270 23968
rect 17334 23904 17350 23968
rect 17414 23904 17430 23968
rect 17494 23904 17500 23968
rect 17184 23903 17500 23904
rect 23900 23968 24216 23969
rect 23900 23904 23906 23968
rect 23970 23904 23986 23968
rect 24050 23904 24066 23968
rect 24130 23904 24146 23968
rect 24210 23904 24216 23968
rect 23900 23903 24216 23904
rect 3785 23626 3851 23629
rect 4981 23626 5047 23629
rect 3785 23624 5047 23626
rect 3785 23568 3790 23624
rect 3846 23568 4986 23624
rect 5042 23568 5047 23624
rect 3785 23566 5047 23568
rect 3785 23563 3851 23566
rect 4981 23563 5047 23566
rect 12525 23626 12591 23629
rect 13261 23626 13327 23629
rect 17902 23626 17908 23628
rect 12525 23624 17908 23626
rect 12525 23568 12530 23624
rect 12586 23568 13266 23624
rect 13322 23568 17908 23624
rect 12525 23566 17908 23568
rect 12525 23563 12591 23566
rect 13261 23563 13327 23566
rect 17902 23564 17908 23566
rect 17972 23564 17978 23628
rect 7110 23424 7426 23425
rect 7110 23360 7116 23424
rect 7180 23360 7196 23424
rect 7260 23360 7276 23424
rect 7340 23360 7356 23424
rect 7420 23360 7426 23424
rect 7110 23359 7426 23360
rect 13826 23424 14142 23425
rect 13826 23360 13832 23424
rect 13896 23360 13912 23424
rect 13976 23360 13992 23424
rect 14056 23360 14072 23424
rect 14136 23360 14142 23424
rect 13826 23359 14142 23360
rect 20542 23424 20858 23425
rect 20542 23360 20548 23424
rect 20612 23360 20628 23424
rect 20692 23360 20708 23424
rect 20772 23360 20788 23424
rect 20852 23360 20858 23424
rect 20542 23359 20858 23360
rect 27258 23424 27574 23425
rect 27258 23360 27264 23424
rect 27328 23360 27344 23424
rect 27408 23360 27424 23424
rect 27488 23360 27504 23424
rect 27568 23360 27574 23424
rect 27258 23359 27574 23360
rect 6637 23354 6703 23357
rect 6637 23352 6746 23354
rect 6637 23296 6642 23352
rect 6698 23296 6746 23352
rect 6637 23291 6746 23296
rect 6177 23218 6243 23221
rect 6686 23218 6746 23291
rect 7606 23294 12450 23354
rect 7606 23218 7666 23294
rect 6177 23216 7666 23218
rect 6177 23160 6182 23216
rect 6238 23160 7666 23216
rect 6177 23158 7666 23160
rect 7741 23218 7807 23221
rect 10317 23218 10383 23221
rect 12390 23218 12450 23294
rect 15377 23218 15443 23221
rect 7741 23216 10426 23218
rect 7741 23160 7746 23216
rect 7802 23160 10322 23216
rect 10378 23160 10426 23216
rect 7741 23158 10426 23160
rect 12390 23216 15443 23218
rect 12390 23160 15382 23216
rect 15438 23160 15443 23216
rect 12390 23158 15443 23160
rect 6177 23155 6243 23158
rect 7741 23155 7807 23158
rect 10317 23155 10426 23158
rect 15377 23155 15443 23158
rect 10366 23082 10426 23155
rect 15837 23082 15903 23085
rect 10366 23080 15903 23082
rect 10366 23024 15842 23080
rect 15898 23024 15903 23080
rect 10366 23022 15903 23024
rect 15837 23019 15903 23022
rect 3752 22880 4068 22881
rect 3752 22816 3758 22880
rect 3822 22816 3838 22880
rect 3902 22816 3918 22880
rect 3982 22816 3998 22880
rect 4062 22816 4068 22880
rect 3752 22815 4068 22816
rect 10468 22880 10784 22881
rect 10468 22816 10474 22880
rect 10538 22816 10554 22880
rect 10618 22816 10634 22880
rect 10698 22816 10714 22880
rect 10778 22816 10784 22880
rect 10468 22815 10784 22816
rect 17184 22880 17500 22881
rect 17184 22816 17190 22880
rect 17254 22816 17270 22880
rect 17334 22816 17350 22880
rect 17414 22816 17430 22880
rect 17494 22816 17500 22880
rect 17184 22815 17500 22816
rect 23900 22880 24216 22881
rect 23900 22816 23906 22880
rect 23970 22816 23986 22880
rect 24050 22816 24066 22880
rect 24130 22816 24146 22880
rect 24210 22816 24216 22880
rect 23900 22815 24216 22816
rect 7110 22336 7426 22337
rect 7110 22272 7116 22336
rect 7180 22272 7196 22336
rect 7260 22272 7276 22336
rect 7340 22272 7356 22336
rect 7420 22272 7426 22336
rect 7110 22271 7426 22272
rect 13826 22336 14142 22337
rect 13826 22272 13832 22336
rect 13896 22272 13912 22336
rect 13976 22272 13992 22336
rect 14056 22272 14072 22336
rect 14136 22272 14142 22336
rect 13826 22271 14142 22272
rect 20542 22336 20858 22337
rect 20542 22272 20548 22336
rect 20612 22272 20628 22336
rect 20692 22272 20708 22336
rect 20772 22272 20788 22336
rect 20852 22272 20858 22336
rect 20542 22271 20858 22272
rect 27258 22336 27574 22337
rect 27258 22272 27264 22336
rect 27328 22272 27344 22336
rect 27408 22272 27424 22336
rect 27488 22272 27504 22336
rect 27568 22272 27574 22336
rect 27258 22271 27574 22272
rect 11094 22068 11100 22132
rect 11164 22130 11170 22132
rect 11237 22130 11303 22133
rect 16205 22130 16271 22133
rect 18137 22130 18203 22133
rect 11164 22128 18203 22130
rect 11164 22072 11242 22128
rect 11298 22072 16210 22128
rect 16266 22072 18142 22128
rect 18198 22072 18203 22128
rect 11164 22070 18203 22072
rect 11164 22068 11170 22070
rect 11237 22067 11303 22070
rect 16205 22067 16271 22070
rect 18137 22067 18203 22070
rect 5206 21932 5212 21996
rect 5276 21994 5282 21996
rect 5349 21994 5415 21997
rect 5276 21992 5415 21994
rect 5276 21936 5354 21992
rect 5410 21936 5415 21992
rect 5276 21934 5415 21936
rect 5276 21932 5282 21934
rect 5349 21931 5415 21934
rect 11053 21994 11119 21997
rect 11278 21994 11284 21996
rect 11053 21992 11284 21994
rect 11053 21936 11058 21992
rect 11114 21936 11284 21992
rect 11053 21934 11284 21936
rect 11053 21931 11119 21934
rect 11278 21932 11284 21934
rect 11348 21994 11354 21996
rect 17769 21994 17835 21997
rect 11348 21992 17835 21994
rect 11348 21936 17774 21992
rect 17830 21936 17835 21992
rect 11348 21934 17835 21936
rect 11348 21932 11354 21934
rect 17769 21931 17835 21934
rect 3752 21792 4068 21793
rect 3752 21728 3758 21792
rect 3822 21728 3838 21792
rect 3902 21728 3918 21792
rect 3982 21728 3998 21792
rect 4062 21728 4068 21792
rect 3752 21727 4068 21728
rect 10468 21792 10784 21793
rect 10468 21728 10474 21792
rect 10538 21728 10554 21792
rect 10618 21728 10634 21792
rect 10698 21728 10714 21792
rect 10778 21728 10784 21792
rect 10468 21727 10784 21728
rect 17184 21792 17500 21793
rect 17184 21728 17190 21792
rect 17254 21728 17270 21792
rect 17334 21728 17350 21792
rect 17414 21728 17430 21792
rect 17494 21728 17500 21792
rect 17184 21727 17500 21728
rect 23900 21792 24216 21793
rect 23900 21728 23906 21792
rect 23970 21728 23986 21792
rect 24050 21728 24066 21792
rect 24130 21728 24146 21792
rect 24210 21728 24216 21792
rect 23900 21727 24216 21728
rect 13445 21450 13511 21453
rect 16205 21450 16271 21453
rect 13445 21448 16271 21450
rect 13445 21392 13450 21448
rect 13506 21392 16210 21448
rect 16266 21392 16271 21448
rect 13445 21390 16271 21392
rect 13445 21387 13511 21390
rect 16205 21387 16271 21390
rect 7110 21248 7426 21249
rect 7110 21184 7116 21248
rect 7180 21184 7196 21248
rect 7260 21184 7276 21248
rect 7340 21184 7356 21248
rect 7420 21184 7426 21248
rect 7110 21183 7426 21184
rect 13826 21248 14142 21249
rect 13826 21184 13832 21248
rect 13896 21184 13912 21248
rect 13976 21184 13992 21248
rect 14056 21184 14072 21248
rect 14136 21184 14142 21248
rect 13826 21183 14142 21184
rect 20542 21248 20858 21249
rect 20542 21184 20548 21248
rect 20612 21184 20628 21248
rect 20692 21184 20708 21248
rect 20772 21184 20788 21248
rect 20852 21184 20858 21248
rect 20542 21183 20858 21184
rect 27258 21248 27574 21249
rect 27258 21184 27264 21248
rect 27328 21184 27344 21248
rect 27408 21184 27424 21248
rect 27488 21184 27504 21248
rect 27568 21184 27574 21248
rect 27258 21183 27574 21184
rect 9673 21042 9739 21045
rect 10041 21042 10107 21045
rect 17033 21042 17099 21045
rect 9673 21040 17099 21042
rect 9673 20984 9678 21040
rect 9734 20984 10046 21040
rect 10102 20984 17038 21040
rect 17094 20984 17099 21040
rect 9673 20982 17099 20984
rect 9673 20979 9739 20982
rect 10041 20979 10107 20982
rect 17033 20979 17099 20982
rect 3752 20704 4068 20705
rect 3752 20640 3758 20704
rect 3822 20640 3838 20704
rect 3902 20640 3918 20704
rect 3982 20640 3998 20704
rect 4062 20640 4068 20704
rect 3752 20639 4068 20640
rect 10468 20704 10784 20705
rect 10468 20640 10474 20704
rect 10538 20640 10554 20704
rect 10618 20640 10634 20704
rect 10698 20640 10714 20704
rect 10778 20640 10784 20704
rect 10468 20639 10784 20640
rect 17184 20704 17500 20705
rect 17184 20640 17190 20704
rect 17254 20640 17270 20704
rect 17334 20640 17350 20704
rect 17414 20640 17430 20704
rect 17494 20640 17500 20704
rect 17184 20639 17500 20640
rect 23900 20704 24216 20705
rect 23900 20640 23906 20704
rect 23970 20640 23986 20704
rect 24050 20640 24066 20704
rect 24130 20640 24146 20704
rect 24210 20640 24216 20704
rect 23900 20639 24216 20640
rect 9673 20498 9739 20501
rect 11973 20498 12039 20501
rect 18229 20498 18295 20501
rect 9673 20496 18295 20498
rect 9673 20440 9678 20496
rect 9734 20440 11978 20496
rect 12034 20440 18234 20496
rect 18290 20440 18295 20496
rect 9673 20438 18295 20440
rect 9673 20435 9739 20438
rect 11973 20435 12039 20438
rect 18229 20435 18295 20438
rect 7110 20160 7426 20161
rect 7110 20096 7116 20160
rect 7180 20096 7196 20160
rect 7260 20096 7276 20160
rect 7340 20096 7356 20160
rect 7420 20096 7426 20160
rect 7110 20095 7426 20096
rect 13826 20160 14142 20161
rect 13826 20096 13832 20160
rect 13896 20096 13912 20160
rect 13976 20096 13992 20160
rect 14056 20096 14072 20160
rect 14136 20096 14142 20160
rect 13826 20095 14142 20096
rect 20542 20160 20858 20161
rect 20542 20096 20548 20160
rect 20612 20096 20628 20160
rect 20692 20096 20708 20160
rect 20772 20096 20788 20160
rect 20852 20096 20858 20160
rect 20542 20095 20858 20096
rect 27258 20160 27574 20161
rect 27258 20096 27264 20160
rect 27328 20096 27344 20160
rect 27408 20096 27424 20160
rect 27488 20096 27504 20160
rect 27568 20096 27574 20160
rect 27258 20095 27574 20096
rect 15653 19818 15719 19821
rect 16062 19818 16068 19820
rect 15653 19816 16068 19818
rect 15653 19760 15658 19816
rect 15714 19760 16068 19816
rect 15653 19758 16068 19760
rect 15653 19755 15719 19758
rect 16062 19756 16068 19758
rect 16132 19756 16138 19820
rect 3752 19616 4068 19617
rect 3752 19552 3758 19616
rect 3822 19552 3838 19616
rect 3902 19552 3918 19616
rect 3982 19552 3998 19616
rect 4062 19552 4068 19616
rect 3752 19551 4068 19552
rect 10468 19616 10784 19617
rect 10468 19552 10474 19616
rect 10538 19552 10554 19616
rect 10618 19552 10634 19616
rect 10698 19552 10714 19616
rect 10778 19552 10784 19616
rect 10468 19551 10784 19552
rect 17184 19616 17500 19617
rect 17184 19552 17190 19616
rect 17254 19552 17270 19616
rect 17334 19552 17350 19616
rect 17414 19552 17430 19616
rect 17494 19552 17500 19616
rect 17184 19551 17500 19552
rect 23900 19616 24216 19617
rect 23900 19552 23906 19616
rect 23970 19552 23986 19616
rect 24050 19552 24066 19616
rect 24130 19552 24146 19616
rect 24210 19552 24216 19616
rect 23900 19551 24216 19552
rect 12566 19348 12572 19412
rect 12636 19410 12642 19412
rect 14181 19410 14247 19413
rect 12636 19408 14247 19410
rect 12636 19352 14186 19408
rect 14242 19352 14247 19408
rect 12636 19350 14247 19352
rect 12636 19348 12642 19350
rect 14181 19347 14247 19350
rect 16614 19212 16620 19276
rect 16684 19274 16690 19276
rect 16757 19274 16823 19277
rect 17217 19274 17283 19277
rect 16684 19272 17283 19274
rect 16684 19216 16762 19272
rect 16818 19216 17222 19272
rect 17278 19216 17283 19272
rect 16684 19214 17283 19216
rect 16684 19212 16690 19214
rect 16757 19211 16823 19214
rect 17217 19211 17283 19214
rect 17585 19274 17651 19277
rect 17718 19274 17724 19276
rect 17585 19272 17724 19274
rect 17585 19216 17590 19272
rect 17646 19216 17724 19272
rect 17585 19214 17724 19216
rect 17585 19211 17651 19214
rect 17718 19212 17724 19214
rect 17788 19212 17794 19276
rect 7110 19072 7426 19073
rect 7110 19008 7116 19072
rect 7180 19008 7196 19072
rect 7260 19008 7276 19072
rect 7340 19008 7356 19072
rect 7420 19008 7426 19072
rect 7110 19007 7426 19008
rect 13826 19072 14142 19073
rect 13826 19008 13832 19072
rect 13896 19008 13912 19072
rect 13976 19008 13992 19072
rect 14056 19008 14072 19072
rect 14136 19008 14142 19072
rect 13826 19007 14142 19008
rect 20542 19072 20858 19073
rect 20542 19008 20548 19072
rect 20612 19008 20628 19072
rect 20692 19008 20708 19072
rect 20772 19008 20788 19072
rect 20852 19008 20858 19072
rect 20542 19007 20858 19008
rect 27258 19072 27574 19073
rect 27258 19008 27264 19072
rect 27328 19008 27344 19072
rect 27408 19008 27424 19072
rect 27488 19008 27504 19072
rect 27568 19008 27574 19072
rect 27258 19007 27574 19008
rect 3752 18528 4068 18529
rect 3752 18464 3758 18528
rect 3822 18464 3838 18528
rect 3902 18464 3918 18528
rect 3982 18464 3998 18528
rect 4062 18464 4068 18528
rect 3752 18463 4068 18464
rect 10468 18528 10784 18529
rect 10468 18464 10474 18528
rect 10538 18464 10554 18528
rect 10618 18464 10634 18528
rect 10698 18464 10714 18528
rect 10778 18464 10784 18528
rect 10468 18463 10784 18464
rect 17184 18528 17500 18529
rect 17184 18464 17190 18528
rect 17254 18464 17270 18528
rect 17334 18464 17350 18528
rect 17414 18464 17430 18528
rect 17494 18464 17500 18528
rect 17184 18463 17500 18464
rect 23900 18528 24216 18529
rect 23900 18464 23906 18528
rect 23970 18464 23986 18528
rect 24050 18464 24066 18528
rect 24130 18464 24146 18528
rect 24210 18464 24216 18528
rect 23900 18463 24216 18464
rect 17677 18322 17743 18325
rect 17902 18322 17908 18324
rect 17677 18320 17908 18322
rect 17677 18264 17682 18320
rect 17738 18264 17908 18320
rect 17677 18262 17908 18264
rect 17677 18259 17743 18262
rect 17902 18260 17908 18262
rect 17972 18260 17978 18324
rect 15101 18186 15167 18189
rect 16113 18186 16179 18189
rect 15101 18184 16179 18186
rect 15101 18128 15106 18184
rect 15162 18128 16118 18184
rect 16174 18128 16179 18184
rect 15101 18126 16179 18128
rect 15101 18123 15167 18126
rect 16113 18123 16179 18126
rect 7110 17984 7426 17985
rect 7110 17920 7116 17984
rect 7180 17920 7196 17984
rect 7260 17920 7276 17984
rect 7340 17920 7356 17984
rect 7420 17920 7426 17984
rect 7110 17919 7426 17920
rect 13826 17984 14142 17985
rect 13826 17920 13832 17984
rect 13896 17920 13912 17984
rect 13976 17920 13992 17984
rect 14056 17920 14072 17984
rect 14136 17920 14142 17984
rect 13826 17919 14142 17920
rect 20542 17984 20858 17985
rect 20542 17920 20548 17984
rect 20612 17920 20628 17984
rect 20692 17920 20708 17984
rect 20772 17920 20788 17984
rect 20852 17920 20858 17984
rect 20542 17919 20858 17920
rect 27258 17984 27574 17985
rect 27258 17920 27264 17984
rect 27328 17920 27344 17984
rect 27408 17920 27424 17984
rect 27488 17920 27504 17984
rect 27568 17920 27574 17984
rect 27258 17919 27574 17920
rect 10041 17914 10107 17917
rect 11094 17914 11100 17916
rect 10041 17912 11100 17914
rect 10041 17856 10046 17912
rect 10102 17856 11100 17912
rect 10041 17854 11100 17856
rect 10041 17851 10107 17854
rect 11094 17852 11100 17854
rect 11164 17852 11170 17916
rect 3752 17440 4068 17441
rect 3752 17376 3758 17440
rect 3822 17376 3838 17440
rect 3902 17376 3918 17440
rect 3982 17376 3998 17440
rect 4062 17376 4068 17440
rect 3752 17375 4068 17376
rect 10468 17440 10784 17441
rect 10468 17376 10474 17440
rect 10538 17376 10554 17440
rect 10618 17376 10634 17440
rect 10698 17376 10714 17440
rect 10778 17376 10784 17440
rect 10468 17375 10784 17376
rect 17184 17440 17500 17441
rect 17184 17376 17190 17440
rect 17254 17376 17270 17440
rect 17334 17376 17350 17440
rect 17414 17376 17430 17440
rect 17494 17376 17500 17440
rect 17184 17375 17500 17376
rect 23900 17440 24216 17441
rect 23900 17376 23906 17440
rect 23970 17376 23986 17440
rect 24050 17376 24066 17440
rect 24130 17376 24146 17440
rect 24210 17376 24216 17440
rect 23900 17375 24216 17376
rect 7110 16896 7426 16897
rect 7110 16832 7116 16896
rect 7180 16832 7196 16896
rect 7260 16832 7276 16896
rect 7340 16832 7356 16896
rect 7420 16832 7426 16896
rect 7110 16831 7426 16832
rect 13826 16896 14142 16897
rect 13826 16832 13832 16896
rect 13896 16832 13912 16896
rect 13976 16832 13992 16896
rect 14056 16832 14072 16896
rect 14136 16832 14142 16896
rect 13826 16831 14142 16832
rect 20542 16896 20858 16897
rect 20542 16832 20548 16896
rect 20612 16832 20628 16896
rect 20692 16832 20708 16896
rect 20772 16832 20788 16896
rect 20852 16832 20858 16896
rect 20542 16831 20858 16832
rect 27258 16896 27574 16897
rect 27258 16832 27264 16896
rect 27328 16832 27344 16896
rect 27408 16832 27424 16896
rect 27488 16832 27504 16896
rect 27568 16832 27574 16896
rect 27258 16831 27574 16832
rect 9489 16690 9555 16693
rect 12566 16690 12572 16692
rect 9489 16688 12572 16690
rect 9489 16632 9494 16688
rect 9550 16632 12572 16688
rect 9489 16630 12572 16632
rect 9489 16627 9555 16630
rect 12566 16628 12572 16630
rect 12636 16628 12642 16692
rect 15929 16690 15995 16693
rect 16062 16690 16068 16692
rect 15929 16688 16068 16690
rect 15929 16632 15934 16688
rect 15990 16632 16068 16688
rect 15929 16630 16068 16632
rect 15929 16627 15995 16630
rect 16062 16628 16068 16630
rect 16132 16628 16138 16692
rect 3752 16352 4068 16353
rect 3752 16288 3758 16352
rect 3822 16288 3838 16352
rect 3902 16288 3918 16352
rect 3982 16288 3998 16352
rect 4062 16288 4068 16352
rect 3752 16287 4068 16288
rect 10468 16352 10784 16353
rect 10468 16288 10474 16352
rect 10538 16288 10554 16352
rect 10618 16288 10634 16352
rect 10698 16288 10714 16352
rect 10778 16288 10784 16352
rect 10468 16287 10784 16288
rect 17184 16352 17500 16353
rect 17184 16288 17190 16352
rect 17254 16288 17270 16352
rect 17334 16288 17350 16352
rect 17414 16288 17430 16352
rect 17494 16288 17500 16352
rect 17184 16287 17500 16288
rect 23900 16352 24216 16353
rect 23900 16288 23906 16352
rect 23970 16288 23986 16352
rect 24050 16288 24066 16352
rect 24130 16288 24146 16352
rect 24210 16288 24216 16352
rect 23900 16287 24216 16288
rect 7110 15808 7426 15809
rect 7110 15744 7116 15808
rect 7180 15744 7196 15808
rect 7260 15744 7276 15808
rect 7340 15744 7356 15808
rect 7420 15744 7426 15808
rect 7110 15743 7426 15744
rect 13826 15808 14142 15809
rect 13826 15744 13832 15808
rect 13896 15744 13912 15808
rect 13976 15744 13992 15808
rect 14056 15744 14072 15808
rect 14136 15744 14142 15808
rect 13826 15743 14142 15744
rect 20542 15808 20858 15809
rect 20542 15744 20548 15808
rect 20612 15744 20628 15808
rect 20692 15744 20708 15808
rect 20772 15744 20788 15808
rect 20852 15744 20858 15808
rect 20542 15743 20858 15744
rect 27258 15808 27574 15809
rect 27258 15744 27264 15808
rect 27328 15744 27344 15808
rect 27408 15744 27424 15808
rect 27488 15744 27504 15808
rect 27568 15744 27574 15808
rect 27258 15743 27574 15744
rect 21725 15738 21791 15741
rect 22093 15738 22159 15741
rect 21725 15736 22159 15738
rect 21725 15680 21730 15736
rect 21786 15680 22098 15736
rect 22154 15680 22159 15736
rect 21725 15678 22159 15680
rect 21725 15675 21791 15678
rect 22093 15675 22159 15678
rect 1669 15602 1735 15605
rect 5206 15602 5212 15604
rect 1669 15600 5212 15602
rect 1669 15544 1674 15600
rect 1730 15544 5212 15600
rect 1669 15542 5212 15544
rect 1669 15539 1735 15542
rect 5206 15540 5212 15542
rect 5276 15540 5282 15604
rect 3752 15264 4068 15265
rect 3752 15200 3758 15264
rect 3822 15200 3838 15264
rect 3902 15200 3918 15264
rect 3982 15200 3998 15264
rect 4062 15200 4068 15264
rect 3752 15199 4068 15200
rect 10468 15264 10784 15265
rect 10468 15200 10474 15264
rect 10538 15200 10554 15264
rect 10618 15200 10634 15264
rect 10698 15200 10714 15264
rect 10778 15200 10784 15264
rect 10468 15199 10784 15200
rect 17184 15264 17500 15265
rect 17184 15200 17190 15264
rect 17254 15200 17270 15264
rect 17334 15200 17350 15264
rect 17414 15200 17430 15264
rect 17494 15200 17500 15264
rect 17184 15199 17500 15200
rect 23900 15264 24216 15265
rect 23900 15200 23906 15264
rect 23970 15200 23986 15264
rect 24050 15200 24066 15264
rect 24130 15200 24146 15264
rect 24210 15200 24216 15264
rect 23900 15199 24216 15200
rect 11237 15196 11303 15197
rect 11237 15192 11284 15196
rect 11348 15194 11354 15196
rect 11237 15136 11242 15192
rect 11237 15132 11284 15136
rect 11348 15134 11394 15194
rect 11348 15132 11354 15134
rect 11237 15131 11303 15132
rect 7110 14720 7426 14721
rect 7110 14656 7116 14720
rect 7180 14656 7196 14720
rect 7260 14656 7276 14720
rect 7340 14656 7356 14720
rect 7420 14656 7426 14720
rect 7110 14655 7426 14656
rect 13826 14720 14142 14721
rect 13826 14656 13832 14720
rect 13896 14656 13912 14720
rect 13976 14656 13992 14720
rect 14056 14656 14072 14720
rect 14136 14656 14142 14720
rect 13826 14655 14142 14656
rect 20542 14720 20858 14721
rect 20542 14656 20548 14720
rect 20612 14656 20628 14720
rect 20692 14656 20708 14720
rect 20772 14656 20788 14720
rect 20852 14656 20858 14720
rect 20542 14655 20858 14656
rect 27258 14720 27574 14721
rect 27258 14656 27264 14720
rect 27328 14656 27344 14720
rect 27408 14656 27424 14720
rect 27488 14656 27504 14720
rect 27568 14656 27574 14720
rect 27258 14655 27574 14656
rect 3752 14176 4068 14177
rect 3752 14112 3758 14176
rect 3822 14112 3838 14176
rect 3902 14112 3918 14176
rect 3982 14112 3998 14176
rect 4062 14112 4068 14176
rect 3752 14111 4068 14112
rect 10468 14176 10784 14177
rect 10468 14112 10474 14176
rect 10538 14112 10554 14176
rect 10618 14112 10634 14176
rect 10698 14112 10714 14176
rect 10778 14112 10784 14176
rect 10468 14111 10784 14112
rect 17184 14176 17500 14177
rect 17184 14112 17190 14176
rect 17254 14112 17270 14176
rect 17334 14112 17350 14176
rect 17414 14112 17430 14176
rect 17494 14112 17500 14176
rect 17184 14111 17500 14112
rect 23900 14176 24216 14177
rect 23900 14112 23906 14176
rect 23970 14112 23986 14176
rect 24050 14112 24066 14176
rect 24130 14112 24146 14176
rect 24210 14112 24216 14176
rect 23900 14111 24216 14112
rect 12566 13908 12572 13972
rect 12636 13970 12642 13972
rect 13721 13970 13787 13973
rect 12636 13968 13787 13970
rect 12636 13912 13726 13968
rect 13782 13912 13787 13968
rect 12636 13910 13787 13912
rect 12636 13908 12642 13910
rect 13721 13907 13787 13910
rect 7110 13632 7426 13633
rect 7110 13568 7116 13632
rect 7180 13568 7196 13632
rect 7260 13568 7276 13632
rect 7340 13568 7356 13632
rect 7420 13568 7426 13632
rect 7110 13567 7426 13568
rect 13826 13632 14142 13633
rect 13826 13568 13832 13632
rect 13896 13568 13912 13632
rect 13976 13568 13992 13632
rect 14056 13568 14072 13632
rect 14136 13568 14142 13632
rect 13826 13567 14142 13568
rect 20542 13632 20858 13633
rect 20542 13568 20548 13632
rect 20612 13568 20628 13632
rect 20692 13568 20708 13632
rect 20772 13568 20788 13632
rect 20852 13568 20858 13632
rect 20542 13567 20858 13568
rect 27258 13632 27574 13633
rect 27258 13568 27264 13632
rect 27328 13568 27344 13632
rect 27408 13568 27424 13632
rect 27488 13568 27504 13632
rect 27568 13568 27574 13632
rect 27258 13567 27574 13568
rect 3752 13088 4068 13089
rect 3752 13024 3758 13088
rect 3822 13024 3838 13088
rect 3902 13024 3918 13088
rect 3982 13024 3998 13088
rect 4062 13024 4068 13088
rect 3752 13023 4068 13024
rect 10468 13088 10784 13089
rect 10468 13024 10474 13088
rect 10538 13024 10554 13088
rect 10618 13024 10634 13088
rect 10698 13024 10714 13088
rect 10778 13024 10784 13088
rect 10468 13023 10784 13024
rect 17184 13088 17500 13089
rect 17184 13024 17190 13088
rect 17254 13024 17270 13088
rect 17334 13024 17350 13088
rect 17414 13024 17430 13088
rect 17494 13024 17500 13088
rect 17184 13023 17500 13024
rect 23900 13088 24216 13089
rect 23900 13024 23906 13088
rect 23970 13024 23986 13088
rect 24050 13024 24066 13088
rect 24130 13024 24146 13088
rect 24210 13024 24216 13088
rect 23900 13023 24216 13024
rect 7110 12544 7426 12545
rect 7110 12480 7116 12544
rect 7180 12480 7196 12544
rect 7260 12480 7276 12544
rect 7340 12480 7356 12544
rect 7420 12480 7426 12544
rect 7110 12479 7426 12480
rect 13826 12544 14142 12545
rect 13826 12480 13832 12544
rect 13896 12480 13912 12544
rect 13976 12480 13992 12544
rect 14056 12480 14072 12544
rect 14136 12480 14142 12544
rect 13826 12479 14142 12480
rect 20542 12544 20858 12545
rect 20542 12480 20548 12544
rect 20612 12480 20628 12544
rect 20692 12480 20708 12544
rect 20772 12480 20788 12544
rect 20852 12480 20858 12544
rect 20542 12479 20858 12480
rect 27258 12544 27574 12545
rect 27258 12480 27264 12544
rect 27328 12480 27344 12544
rect 27408 12480 27424 12544
rect 27488 12480 27504 12544
rect 27568 12480 27574 12544
rect 27258 12479 27574 12480
rect 3752 12000 4068 12001
rect 3752 11936 3758 12000
rect 3822 11936 3838 12000
rect 3902 11936 3918 12000
rect 3982 11936 3998 12000
rect 4062 11936 4068 12000
rect 3752 11935 4068 11936
rect 10468 12000 10784 12001
rect 10468 11936 10474 12000
rect 10538 11936 10554 12000
rect 10618 11936 10634 12000
rect 10698 11936 10714 12000
rect 10778 11936 10784 12000
rect 10468 11935 10784 11936
rect 17184 12000 17500 12001
rect 17184 11936 17190 12000
rect 17254 11936 17270 12000
rect 17334 11936 17350 12000
rect 17414 11936 17430 12000
rect 17494 11936 17500 12000
rect 17184 11935 17500 11936
rect 23900 12000 24216 12001
rect 23900 11936 23906 12000
rect 23970 11936 23986 12000
rect 24050 11936 24066 12000
rect 24130 11936 24146 12000
rect 24210 11936 24216 12000
rect 23900 11935 24216 11936
rect 7110 11456 7426 11457
rect 7110 11392 7116 11456
rect 7180 11392 7196 11456
rect 7260 11392 7276 11456
rect 7340 11392 7356 11456
rect 7420 11392 7426 11456
rect 7110 11391 7426 11392
rect 13826 11456 14142 11457
rect 13826 11392 13832 11456
rect 13896 11392 13912 11456
rect 13976 11392 13992 11456
rect 14056 11392 14072 11456
rect 14136 11392 14142 11456
rect 13826 11391 14142 11392
rect 20542 11456 20858 11457
rect 20542 11392 20548 11456
rect 20612 11392 20628 11456
rect 20692 11392 20708 11456
rect 20772 11392 20788 11456
rect 20852 11392 20858 11456
rect 20542 11391 20858 11392
rect 27258 11456 27574 11457
rect 27258 11392 27264 11456
rect 27328 11392 27344 11456
rect 27408 11392 27424 11456
rect 27488 11392 27504 11456
rect 27568 11392 27574 11456
rect 27258 11391 27574 11392
rect 3752 10912 4068 10913
rect 3752 10848 3758 10912
rect 3822 10848 3838 10912
rect 3902 10848 3918 10912
rect 3982 10848 3998 10912
rect 4062 10848 4068 10912
rect 3752 10847 4068 10848
rect 10468 10912 10784 10913
rect 10468 10848 10474 10912
rect 10538 10848 10554 10912
rect 10618 10848 10634 10912
rect 10698 10848 10714 10912
rect 10778 10848 10784 10912
rect 10468 10847 10784 10848
rect 17184 10912 17500 10913
rect 17184 10848 17190 10912
rect 17254 10848 17270 10912
rect 17334 10848 17350 10912
rect 17414 10848 17430 10912
rect 17494 10848 17500 10912
rect 17184 10847 17500 10848
rect 23900 10912 24216 10913
rect 23900 10848 23906 10912
rect 23970 10848 23986 10912
rect 24050 10848 24066 10912
rect 24130 10848 24146 10912
rect 24210 10848 24216 10912
rect 23900 10847 24216 10848
rect 17769 10842 17835 10845
rect 18229 10842 18295 10845
rect 17726 10840 18295 10842
rect 17726 10784 17774 10840
rect 17830 10784 18234 10840
rect 18290 10784 18295 10840
rect 17726 10782 18295 10784
rect 17726 10779 17835 10782
rect 18229 10779 18295 10782
rect 13997 10706 14063 10709
rect 17726 10706 17786 10779
rect 13997 10704 17786 10706
rect 13997 10648 14002 10704
rect 14058 10648 17786 10704
rect 13997 10646 17786 10648
rect 13997 10643 14063 10646
rect 12157 10570 12223 10573
rect 12433 10570 12499 10573
rect 17217 10570 17283 10573
rect 12157 10568 17283 10570
rect 12157 10512 12162 10568
rect 12218 10512 12438 10568
rect 12494 10512 17222 10568
rect 17278 10512 17283 10568
rect 12157 10510 17283 10512
rect 12157 10507 12223 10510
rect 12433 10507 12499 10510
rect 17217 10507 17283 10510
rect 7110 10368 7426 10369
rect 7110 10304 7116 10368
rect 7180 10304 7196 10368
rect 7260 10304 7276 10368
rect 7340 10304 7356 10368
rect 7420 10304 7426 10368
rect 7110 10303 7426 10304
rect 13826 10368 14142 10369
rect 13826 10304 13832 10368
rect 13896 10304 13912 10368
rect 13976 10304 13992 10368
rect 14056 10304 14072 10368
rect 14136 10304 14142 10368
rect 13826 10303 14142 10304
rect 20542 10368 20858 10369
rect 20542 10304 20548 10368
rect 20612 10304 20628 10368
rect 20692 10304 20708 10368
rect 20772 10304 20788 10368
rect 20852 10304 20858 10368
rect 20542 10303 20858 10304
rect 27258 10368 27574 10369
rect 27258 10304 27264 10368
rect 27328 10304 27344 10368
rect 27408 10304 27424 10368
rect 27488 10304 27504 10368
rect 27568 10304 27574 10368
rect 27258 10303 27574 10304
rect 2865 10162 2931 10165
rect 4245 10162 4311 10165
rect 2865 10160 4311 10162
rect 2865 10104 2870 10160
rect 2926 10104 4250 10160
rect 4306 10104 4311 10160
rect 2865 10102 4311 10104
rect 2865 10099 2931 10102
rect 4245 10099 4311 10102
rect 2313 10026 2379 10029
rect 3141 10026 3207 10029
rect 2313 10024 3207 10026
rect 2313 9968 2318 10024
rect 2374 9968 3146 10024
rect 3202 9968 3207 10024
rect 2313 9966 3207 9968
rect 2313 9963 2379 9966
rect 3141 9963 3207 9966
rect 12341 10026 12407 10029
rect 12617 10026 12683 10029
rect 12341 10024 12683 10026
rect 12341 9968 12346 10024
rect 12402 9968 12622 10024
rect 12678 9968 12683 10024
rect 12341 9966 12683 9968
rect 12341 9963 12407 9966
rect 12617 9963 12683 9966
rect 3752 9824 4068 9825
rect 3752 9760 3758 9824
rect 3822 9760 3838 9824
rect 3902 9760 3918 9824
rect 3982 9760 3998 9824
rect 4062 9760 4068 9824
rect 3752 9759 4068 9760
rect 10468 9824 10784 9825
rect 10468 9760 10474 9824
rect 10538 9760 10554 9824
rect 10618 9760 10634 9824
rect 10698 9760 10714 9824
rect 10778 9760 10784 9824
rect 10468 9759 10784 9760
rect 17184 9824 17500 9825
rect 17184 9760 17190 9824
rect 17254 9760 17270 9824
rect 17334 9760 17350 9824
rect 17414 9760 17430 9824
rect 17494 9760 17500 9824
rect 17184 9759 17500 9760
rect 23900 9824 24216 9825
rect 23900 9760 23906 9824
rect 23970 9760 23986 9824
rect 24050 9760 24066 9824
rect 24130 9760 24146 9824
rect 24210 9760 24216 9824
rect 23900 9759 24216 9760
rect 12065 9618 12131 9621
rect 14181 9618 14247 9621
rect 12065 9616 14247 9618
rect 12065 9560 12070 9616
rect 12126 9560 14186 9616
rect 14242 9560 14247 9616
rect 12065 9558 14247 9560
rect 12065 9555 12131 9558
rect 14181 9555 14247 9558
rect 7110 9280 7426 9281
rect 7110 9216 7116 9280
rect 7180 9216 7196 9280
rect 7260 9216 7276 9280
rect 7340 9216 7356 9280
rect 7420 9216 7426 9280
rect 7110 9215 7426 9216
rect 13826 9280 14142 9281
rect 13826 9216 13832 9280
rect 13896 9216 13912 9280
rect 13976 9216 13992 9280
rect 14056 9216 14072 9280
rect 14136 9216 14142 9280
rect 13826 9215 14142 9216
rect 20542 9280 20858 9281
rect 20542 9216 20548 9280
rect 20612 9216 20628 9280
rect 20692 9216 20708 9280
rect 20772 9216 20788 9280
rect 20852 9216 20858 9280
rect 20542 9215 20858 9216
rect 27258 9280 27574 9281
rect 27258 9216 27264 9280
rect 27328 9216 27344 9280
rect 27408 9216 27424 9280
rect 27488 9216 27504 9280
rect 27568 9216 27574 9280
rect 27258 9215 27574 9216
rect 12617 9074 12683 9077
rect 14181 9074 14247 9077
rect 18137 9074 18203 9077
rect 12617 9072 18203 9074
rect 12617 9016 12622 9072
rect 12678 9016 14186 9072
rect 14242 9016 18142 9072
rect 18198 9016 18203 9072
rect 12617 9014 18203 9016
rect 12617 9011 12683 9014
rect 14181 9011 14247 9014
rect 18137 9011 18203 9014
rect 3752 8736 4068 8737
rect 3752 8672 3758 8736
rect 3822 8672 3838 8736
rect 3902 8672 3918 8736
rect 3982 8672 3998 8736
rect 4062 8672 4068 8736
rect 3752 8671 4068 8672
rect 10468 8736 10784 8737
rect 10468 8672 10474 8736
rect 10538 8672 10554 8736
rect 10618 8672 10634 8736
rect 10698 8672 10714 8736
rect 10778 8672 10784 8736
rect 10468 8671 10784 8672
rect 17184 8736 17500 8737
rect 17184 8672 17190 8736
rect 17254 8672 17270 8736
rect 17334 8672 17350 8736
rect 17414 8672 17430 8736
rect 17494 8672 17500 8736
rect 17184 8671 17500 8672
rect 23900 8736 24216 8737
rect 23900 8672 23906 8736
rect 23970 8672 23986 8736
rect 24050 8672 24066 8736
rect 24130 8672 24146 8736
rect 24210 8672 24216 8736
rect 23900 8671 24216 8672
rect 14825 8394 14891 8397
rect 15377 8394 15443 8397
rect 14825 8392 15443 8394
rect 14825 8336 14830 8392
rect 14886 8336 15382 8392
rect 15438 8336 15443 8392
rect 14825 8334 15443 8336
rect 14825 8331 14891 8334
rect 15377 8331 15443 8334
rect 7110 8192 7426 8193
rect 7110 8128 7116 8192
rect 7180 8128 7196 8192
rect 7260 8128 7276 8192
rect 7340 8128 7356 8192
rect 7420 8128 7426 8192
rect 7110 8127 7426 8128
rect 13826 8192 14142 8193
rect 13826 8128 13832 8192
rect 13896 8128 13912 8192
rect 13976 8128 13992 8192
rect 14056 8128 14072 8192
rect 14136 8128 14142 8192
rect 13826 8127 14142 8128
rect 20542 8192 20858 8193
rect 20542 8128 20548 8192
rect 20612 8128 20628 8192
rect 20692 8128 20708 8192
rect 20772 8128 20788 8192
rect 20852 8128 20858 8192
rect 20542 8127 20858 8128
rect 27258 8192 27574 8193
rect 27258 8128 27264 8192
rect 27328 8128 27344 8192
rect 27408 8128 27424 8192
rect 27488 8128 27504 8192
rect 27568 8128 27574 8192
rect 27258 8127 27574 8128
rect 3752 7648 4068 7649
rect 3752 7584 3758 7648
rect 3822 7584 3838 7648
rect 3902 7584 3918 7648
rect 3982 7584 3998 7648
rect 4062 7584 4068 7648
rect 3752 7583 4068 7584
rect 10468 7648 10784 7649
rect 10468 7584 10474 7648
rect 10538 7584 10554 7648
rect 10618 7584 10634 7648
rect 10698 7584 10714 7648
rect 10778 7584 10784 7648
rect 10468 7583 10784 7584
rect 17184 7648 17500 7649
rect 17184 7584 17190 7648
rect 17254 7584 17270 7648
rect 17334 7584 17350 7648
rect 17414 7584 17430 7648
rect 17494 7584 17500 7648
rect 17184 7583 17500 7584
rect 23900 7648 24216 7649
rect 23900 7584 23906 7648
rect 23970 7584 23986 7648
rect 24050 7584 24066 7648
rect 24130 7584 24146 7648
rect 24210 7584 24216 7648
rect 23900 7583 24216 7584
rect 7110 7104 7426 7105
rect 7110 7040 7116 7104
rect 7180 7040 7196 7104
rect 7260 7040 7276 7104
rect 7340 7040 7356 7104
rect 7420 7040 7426 7104
rect 7110 7039 7426 7040
rect 13826 7104 14142 7105
rect 13826 7040 13832 7104
rect 13896 7040 13912 7104
rect 13976 7040 13992 7104
rect 14056 7040 14072 7104
rect 14136 7040 14142 7104
rect 13826 7039 14142 7040
rect 20542 7104 20858 7105
rect 20542 7040 20548 7104
rect 20612 7040 20628 7104
rect 20692 7040 20708 7104
rect 20772 7040 20788 7104
rect 20852 7040 20858 7104
rect 20542 7039 20858 7040
rect 27258 7104 27574 7105
rect 27258 7040 27264 7104
rect 27328 7040 27344 7104
rect 27408 7040 27424 7104
rect 27488 7040 27504 7104
rect 27568 7040 27574 7104
rect 27258 7039 27574 7040
rect 3752 6560 4068 6561
rect 3752 6496 3758 6560
rect 3822 6496 3838 6560
rect 3902 6496 3918 6560
rect 3982 6496 3998 6560
rect 4062 6496 4068 6560
rect 3752 6495 4068 6496
rect 10468 6560 10784 6561
rect 10468 6496 10474 6560
rect 10538 6496 10554 6560
rect 10618 6496 10634 6560
rect 10698 6496 10714 6560
rect 10778 6496 10784 6560
rect 10468 6495 10784 6496
rect 17184 6560 17500 6561
rect 17184 6496 17190 6560
rect 17254 6496 17270 6560
rect 17334 6496 17350 6560
rect 17414 6496 17430 6560
rect 17494 6496 17500 6560
rect 17184 6495 17500 6496
rect 23900 6560 24216 6561
rect 23900 6496 23906 6560
rect 23970 6496 23986 6560
rect 24050 6496 24066 6560
rect 24130 6496 24146 6560
rect 24210 6496 24216 6560
rect 23900 6495 24216 6496
rect 7110 6016 7426 6017
rect 7110 5952 7116 6016
rect 7180 5952 7196 6016
rect 7260 5952 7276 6016
rect 7340 5952 7356 6016
rect 7420 5952 7426 6016
rect 7110 5951 7426 5952
rect 13826 6016 14142 6017
rect 13826 5952 13832 6016
rect 13896 5952 13912 6016
rect 13976 5952 13992 6016
rect 14056 5952 14072 6016
rect 14136 5952 14142 6016
rect 13826 5951 14142 5952
rect 20542 6016 20858 6017
rect 20542 5952 20548 6016
rect 20612 5952 20628 6016
rect 20692 5952 20708 6016
rect 20772 5952 20788 6016
rect 20852 5952 20858 6016
rect 20542 5951 20858 5952
rect 27258 6016 27574 6017
rect 27258 5952 27264 6016
rect 27328 5952 27344 6016
rect 27408 5952 27424 6016
rect 27488 5952 27504 6016
rect 27568 5952 27574 6016
rect 27258 5951 27574 5952
rect 3752 5472 4068 5473
rect 3752 5408 3758 5472
rect 3822 5408 3838 5472
rect 3902 5408 3918 5472
rect 3982 5408 3998 5472
rect 4062 5408 4068 5472
rect 3752 5407 4068 5408
rect 10468 5472 10784 5473
rect 10468 5408 10474 5472
rect 10538 5408 10554 5472
rect 10618 5408 10634 5472
rect 10698 5408 10714 5472
rect 10778 5408 10784 5472
rect 10468 5407 10784 5408
rect 17184 5472 17500 5473
rect 17184 5408 17190 5472
rect 17254 5408 17270 5472
rect 17334 5408 17350 5472
rect 17414 5408 17430 5472
rect 17494 5408 17500 5472
rect 17184 5407 17500 5408
rect 23900 5472 24216 5473
rect 23900 5408 23906 5472
rect 23970 5408 23986 5472
rect 24050 5408 24066 5472
rect 24130 5408 24146 5472
rect 24210 5408 24216 5472
rect 23900 5407 24216 5408
rect 7110 4928 7426 4929
rect 7110 4864 7116 4928
rect 7180 4864 7196 4928
rect 7260 4864 7276 4928
rect 7340 4864 7356 4928
rect 7420 4864 7426 4928
rect 7110 4863 7426 4864
rect 13826 4928 14142 4929
rect 13826 4864 13832 4928
rect 13896 4864 13912 4928
rect 13976 4864 13992 4928
rect 14056 4864 14072 4928
rect 14136 4864 14142 4928
rect 13826 4863 14142 4864
rect 20542 4928 20858 4929
rect 20542 4864 20548 4928
rect 20612 4864 20628 4928
rect 20692 4864 20708 4928
rect 20772 4864 20788 4928
rect 20852 4864 20858 4928
rect 20542 4863 20858 4864
rect 27258 4928 27574 4929
rect 27258 4864 27264 4928
rect 27328 4864 27344 4928
rect 27408 4864 27424 4928
rect 27488 4864 27504 4928
rect 27568 4864 27574 4928
rect 27258 4863 27574 4864
rect 3752 4384 4068 4385
rect 3752 4320 3758 4384
rect 3822 4320 3838 4384
rect 3902 4320 3918 4384
rect 3982 4320 3998 4384
rect 4062 4320 4068 4384
rect 3752 4319 4068 4320
rect 10468 4384 10784 4385
rect 10468 4320 10474 4384
rect 10538 4320 10554 4384
rect 10618 4320 10634 4384
rect 10698 4320 10714 4384
rect 10778 4320 10784 4384
rect 10468 4319 10784 4320
rect 17184 4384 17500 4385
rect 17184 4320 17190 4384
rect 17254 4320 17270 4384
rect 17334 4320 17350 4384
rect 17414 4320 17430 4384
rect 17494 4320 17500 4384
rect 17184 4319 17500 4320
rect 23900 4384 24216 4385
rect 23900 4320 23906 4384
rect 23970 4320 23986 4384
rect 24050 4320 24066 4384
rect 24130 4320 24146 4384
rect 24210 4320 24216 4384
rect 23900 4319 24216 4320
rect 7110 3840 7426 3841
rect 7110 3776 7116 3840
rect 7180 3776 7196 3840
rect 7260 3776 7276 3840
rect 7340 3776 7356 3840
rect 7420 3776 7426 3840
rect 7110 3775 7426 3776
rect 13826 3840 14142 3841
rect 13826 3776 13832 3840
rect 13896 3776 13912 3840
rect 13976 3776 13992 3840
rect 14056 3776 14072 3840
rect 14136 3776 14142 3840
rect 13826 3775 14142 3776
rect 20542 3840 20858 3841
rect 20542 3776 20548 3840
rect 20612 3776 20628 3840
rect 20692 3776 20708 3840
rect 20772 3776 20788 3840
rect 20852 3776 20858 3840
rect 20542 3775 20858 3776
rect 27258 3840 27574 3841
rect 27258 3776 27264 3840
rect 27328 3776 27344 3840
rect 27408 3776 27424 3840
rect 27488 3776 27504 3840
rect 27568 3776 27574 3840
rect 27258 3775 27574 3776
rect 3752 3296 4068 3297
rect 3752 3232 3758 3296
rect 3822 3232 3838 3296
rect 3902 3232 3918 3296
rect 3982 3232 3998 3296
rect 4062 3232 4068 3296
rect 3752 3231 4068 3232
rect 10468 3296 10784 3297
rect 10468 3232 10474 3296
rect 10538 3232 10554 3296
rect 10618 3232 10634 3296
rect 10698 3232 10714 3296
rect 10778 3232 10784 3296
rect 10468 3231 10784 3232
rect 17184 3296 17500 3297
rect 17184 3232 17190 3296
rect 17254 3232 17270 3296
rect 17334 3232 17350 3296
rect 17414 3232 17430 3296
rect 17494 3232 17500 3296
rect 17184 3231 17500 3232
rect 23900 3296 24216 3297
rect 23900 3232 23906 3296
rect 23970 3232 23986 3296
rect 24050 3232 24066 3296
rect 24130 3232 24146 3296
rect 24210 3232 24216 3296
rect 23900 3231 24216 3232
rect 13537 3090 13603 3093
rect 15377 3090 15443 3093
rect 13537 3088 15443 3090
rect 13537 3032 13542 3088
rect 13598 3032 15382 3088
rect 15438 3032 15443 3088
rect 13537 3030 15443 3032
rect 13537 3027 13603 3030
rect 15377 3027 15443 3030
rect 11329 2954 11395 2957
rect 13905 2954 13971 2957
rect 15101 2954 15167 2957
rect 11329 2952 15167 2954
rect 11329 2896 11334 2952
rect 11390 2896 13910 2952
rect 13966 2896 15106 2952
rect 15162 2896 15167 2952
rect 11329 2894 15167 2896
rect 11329 2891 11395 2894
rect 13905 2891 13971 2894
rect 15101 2891 15167 2894
rect 21633 2954 21699 2957
rect 23105 2954 23171 2957
rect 21633 2952 23171 2954
rect 21633 2896 21638 2952
rect 21694 2896 23110 2952
rect 23166 2896 23171 2952
rect 21633 2894 23171 2896
rect 21633 2891 21699 2894
rect 23105 2891 23171 2894
rect 7110 2752 7426 2753
rect 7110 2688 7116 2752
rect 7180 2688 7196 2752
rect 7260 2688 7276 2752
rect 7340 2688 7356 2752
rect 7420 2688 7426 2752
rect 7110 2687 7426 2688
rect 13826 2752 14142 2753
rect 13826 2688 13832 2752
rect 13896 2688 13912 2752
rect 13976 2688 13992 2752
rect 14056 2688 14072 2752
rect 14136 2688 14142 2752
rect 13826 2687 14142 2688
rect 20542 2752 20858 2753
rect 20542 2688 20548 2752
rect 20612 2688 20628 2752
rect 20692 2688 20708 2752
rect 20772 2688 20788 2752
rect 20852 2688 20858 2752
rect 20542 2687 20858 2688
rect 27258 2752 27574 2753
rect 27258 2688 27264 2752
rect 27328 2688 27344 2752
rect 27408 2688 27424 2752
rect 27488 2688 27504 2752
rect 27568 2688 27574 2752
rect 27258 2687 27574 2688
rect 3752 2208 4068 2209
rect 3752 2144 3758 2208
rect 3822 2144 3838 2208
rect 3902 2144 3918 2208
rect 3982 2144 3998 2208
rect 4062 2144 4068 2208
rect 3752 2143 4068 2144
rect 10468 2208 10784 2209
rect 10468 2144 10474 2208
rect 10538 2144 10554 2208
rect 10618 2144 10634 2208
rect 10698 2144 10714 2208
rect 10778 2144 10784 2208
rect 10468 2143 10784 2144
rect 17184 2208 17500 2209
rect 17184 2144 17190 2208
rect 17254 2144 17270 2208
rect 17334 2144 17350 2208
rect 17414 2144 17430 2208
rect 17494 2144 17500 2208
rect 17184 2143 17500 2144
rect 23900 2208 24216 2209
rect 23900 2144 23906 2208
rect 23970 2144 23986 2208
rect 24050 2144 24066 2208
rect 24130 2144 24146 2208
rect 24210 2144 24216 2208
rect 23900 2143 24216 2144
rect 7110 1664 7426 1665
rect 7110 1600 7116 1664
rect 7180 1600 7196 1664
rect 7260 1600 7276 1664
rect 7340 1600 7356 1664
rect 7420 1600 7426 1664
rect 7110 1599 7426 1600
rect 13826 1664 14142 1665
rect 13826 1600 13832 1664
rect 13896 1600 13912 1664
rect 13976 1600 13992 1664
rect 14056 1600 14072 1664
rect 14136 1600 14142 1664
rect 13826 1599 14142 1600
rect 20542 1664 20858 1665
rect 20542 1600 20548 1664
rect 20612 1600 20628 1664
rect 20692 1600 20708 1664
rect 20772 1600 20788 1664
rect 20852 1600 20858 1664
rect 20542 1599 20858 1600
rect 27258 1664 27574 1665
rect 27258 1600 27264 1664
rect 27328 1600 27344 1664
rect 27408 1600 27424 1664
rect 27488 1600 27504 1664
rect 27568 1600 27574 1664
rect 27258 1599 27574 1600
rect 3752 1120 4068 1121
rect 3752 1056 3758 1120
rect 3822 1056 3838 1120
rect 3902 1056 3918 1120
rect 3982 1056 3998 1120
rect 4062 1056 4068 1120
rect 3752 1055 4068 1056
rect 10468 1120 10784 1121
rect 10468 1056 10474 1120
rect 10538 1056 10554 1120
rect 10618 1056 10634 1120
rect 10698 1056 10714 1120
rect 10778 1056 10784 1120
rect 10468 1055 10784 1056
rect 17184 1120 17500 1121
rect 17184 1056 17190 1120
rect 17254 1056 17270 1120
rect 17334 1056 17350 1120
rect 17414 1056 17430 1120
rect 17494 1056 17500 1120
rect 17184 1055 17500 1056
rect 23900 1120 24216 1121
rect 23900 1056 23906 1120
rect 23970 1056 23986 1120
rect 24050 1056 24066 1120
rect 24130 1056 24146 1120
rect 24210 1056 24216 1120
rect 23900 1055 24216 1056
rect 7110 576 7426 577
rect 7110 512 7116 576
rect 7180 512 7196 576
rect 7260 512 7276 576
rect 7340 512 7356 576
rect 7420 512 7426 576
rect 7110 511 7426 512
rect 13826 576 14142 577
rect 13826 512 13832 576
rect 13896 512 13912 576
rect 13976 512 13992 576
rect 14056 512 14072 576
rect 14136 512 14142 576
rect 13826 511 14142 512
rect 20542 576 20858 577
rect 20542 512 20548 576
rect 20612 512 20628 576
rect 20692 512 20708 576
rect 20772 512 20788 576
rect 20852 512 20858 576
rect 20542 511 20858 512
rect 27258 576 27574 577
rect 27258 512 27264 576
rect 27328 512 27344 576
rect 27408 512 27424 576
rect 27488 512 27504 576
rect 27568 512 27574 576
rect 27258 511 27574 512
<< via3 >>
rect 7116 31036 7180 31040
rect 7116 30980 7120 31036
rect 7120 30980 7176 31036
rect 7176 30980 7180 31036
rect 7116 30976 7180 30980
rect 7196 31036 7260 31040
rect 7196 30980 7200 31036
rect 7200 30980 7256 31036
rect 7256 30980 7260 31036
rect 7196 30976 7260 30980
rect 7276 31036 7340 31040
rect 7276 30980 7280 31036
rect 7280 30980 7336 31036
rect 7336 30980 7340 31036
rect 7276 30976 7340 30980
rect 7356 31036 7420 31040
rect 7356 30980 7360 31036
rect 7360 30980 7416 31036
rect 7416 30980 7420 31036
rect 7356 30976 7420 30980
rect 13832 31036 13896 31040
rect 13832 30980 13836 31036
rect 13836 30980 13892 31036
rect 13892 30980 13896 31036
rect 13832 30976 13896 30980
rect 13912 31036 13976 31040
rect 13912 30980 13916 31036
rect 13916 30980 13972 31036
rect 13972 30980 13976 31036
rect 13912 30976 13976 30980
rect 13992 31036 14056 31040
rect 13992 30980 13996 31036
rect 13996 30980 14052 31036
rect 14052 30980 14056 31036
rect 13992 30976 14056 30980
rect 14072 31036 14136 31040
rect 14072 30980 14076 31036
rect 14076 30980 14132 31036
rect 14132 30980 14136 31036
rect 14072 30976 14136 30980
rect 20548 31036 20612 31040
rect 20548 30980 20552 31036
rect 20552 30980 20608 31036
rect 20608 30980 20612 31036
rect 20548 30976 20612 30980
rect 20628 31036 20692 31040
rect 20628 30980 20632 31036
rect 20632 30980 20688 31036
rect 20688 30980 20692 31036
rect 20628 30976 20692 30980
rect 20708 31036 20772 31040
rect 20708 30980 20712 31036
rect 20712 30980 20768 31036
rect 20768 30980 20772 31036
rect 20708 30976 20772 30980
rect 20788 31036 20852 31040
rect 20788 30980 20792 31036
rect 20792 30980 20848 31036
rect 20848 30980 20852 31036
rect 20788 30976 20852 30980
rect 27264 31036 27328 31040
rect 27264 30980 27268 31036
rect 27268 30980 27324 31036
rect 27324 30980 27328 31036
rect 27264 30976 27328 30980
rect 27344 31036 27408 31040
rect 27344 30980 27348 31036
rect 27348 30980 27404 31036
rect 27404 30980 27408 31036
rect 27344 30976 27408 30980
rect 27424 31036 27488 31040
rect 27424 30980 27428 31036
rect 27428 30980 27484 31036
rect 27484 30980 27488 31036
rect 27424 30976 27488 30980
rect 27504 31036 27568 31040
rect 27504 30980 27508 31036
rect 27508 30980 27564 31036
rect 27564 30980 27568 31036
rect 27504 30976 27568 30980
rect 3758 30492 3822 30496
rect 3758 30436 3762 30492
rect 3762 30436 3818 30492
rect 3818 30436 3822 30492
rect 3758 30432 3822 30436
rect 3838 30492 3902 30496
rect 3838 30436 3842 30492
rect 3842 30436 3898 30492
rect 3898 30436 3902 30492
rect 3838 30432 3902 30436
rect 3918 30492 3982 30496
rect 3918 30436 3922 30492
rect 3922 30436 3978 30492
rect 3978 30436 3982 30492
rect 3918 30432 3982 30436
rect 3998 30492 4062 30496
rect 3998 30436 4002 30492
rect 4002 30436 4058 30492
rect 4058 30436 4062 30492
rect 3998 30432 4062 30436
rect 10474 30492 10538 30496
rect 10474 30436 10478 30492
rect 10478 30436 10534 30492
rect 10534 30436 10538 30492
rect 10474 30432 10538 30436
rect 10554 30492 10618 30496
rect 10554 30436 10558 30492
rect 10558 30436 10614 30492
rect 10614 30436 10618 30492
rect 10554 30432 10618 30436
rect 10634 30492 10698 30496
rect 10634 30436 10638 30492
rect 10638 30436 10694 30492
rect 10694 30436 10698 30492
rect 10634 30432 10698 30436
rect 10714 30492 10778 30496
rect 10714 30436 10718 30492
rect 10718 30436 10774 30492
rect 10774 30436 10778 30492
rect 10714 30432 10778 30436
rect 17190 30492 17254 30496
rect 17190 30436 17194 30492
rect 17194 30436 17250 30492
rect 17250 30436 17254 30492
rect 17190 30432 17254 30436
rect 17270 30492 17334 30496
rect 17270 30436 17274 30492
rect 17274 30436 17330 30492
rect 17330 30436 17334 30492
rect 17270 30432 17334 30436
rect 17350 30492 17414 30496
rect 17350 30436 17354 30492
rect 17354 30436 17410 30492
rect 17410 30436 17414 30492
rect 17350 30432 17414 30436
rect 17430 30492 17494 30496
rect 17430 30436 17434 30492
rect 17434 30436 17490 30492
rect 17490 30436 17494 30492
rect 17430 30432 17494 30436
rect 23906 30492 23970 30496
rect 23906 30436 23910 30492
rect 23910 30436 23966 30492
rect 23966 30436 23970 30492
rect 23906 30432 23970 30436
rect 23986 30492 24050 30496
rect 23986 30436 23990 30492
rect 23990 30436 24046 30492
rect 24046 30436 24050 30492
rect 23986 30432 24050 30436
rect 24066 30492 24130 30496
rect 24066 30436 24070 30492
rect 24070 30436 24126 30492
rect 24126 30436 24130 30492
rect 24066 30432 24130 30436
rect 24146 30492 24210 30496
rect 24146 30436 24150 30492
rect 24150 30436 24206 30492
rect 24206 30436 24210 30492
rect 24146 30432 24210 30436
rect 7116 29948 7180 29952
rect 7116 29892 7120 29948
rect 7120 29892 7176 29948
rect 7176 29892 7180 29948
rect 7116 29888 7180 29892
rect 7196 29948 7260 29952
rect 7196 29892 7200 29948
rect 7200 29892 7256 29948
rect 7256 29892 7260 29948
rect 7196 29888 7260 29892
rect 7276 29948 7340 29952
rect 7276 29892 7280 29948
rect 7280 29892 7336 29948
rect 7336 29892 7340 29948
rect 7276 29888 7340 29892
rect 7356 29948 7420 29952
rect 7356 29892 7360 29948
rect 7360 29892 7416 29948
rect 7416 29892 7420 29948
rect 7356 29888 7420 29892
rect 13832 29948 13896 29952
rect 13832 29892 13836 29948
rect 13836 29892 13892 29948
rect 13892 29892 13896 29948
rect 13832 29888 13896 29892
rect 13912 29948 13976 29952
rect 13912 29892 13916 29948
rect 13916 29892 13972 29948
rect 13972 29892 13976 29948
rect 13912 29888 13976 29892
rect 13992 29948 14056 29952
rect 13992 29892 13996 29948
rect 13996 29892 14052 29948
rect 14052 29892 14056 29948
rect 13992 29888 14056 29892
rect 14072 29948 14136 29952
rect 14072 29892 14076 29948
rect 14076 29892 14132 29948
rect 14132 29892 14136 29948
rect 14072 29888 14136 29892
rect 20548 29948 20612 29952
rect 20548 29892 20552 29948
rect 20552 29892 20608 29948
rect 20608 29892 20612 29948
rect 20548 29888 20612 29892
rect 20628 29948 20692 29952
rect 20628 29892 20632 29948
rect 20632 29892 20688 29948
rect 20688 29892 20692 29948
rect 20628 29888 20692 29892
rect 20708 29948 20772 29952
rect 20708 29892 20712 29948
rect 20712 29892 20768 29948
rect 20768 29892 20772 29948
rect 20708 29888 20772 29892
rect 20788 29948 20852 29952
rect 20788 29892 20792 29948
rect 20792 29892 20848 29948
rect 20848 29892 20852 29948
rect 20788 29888 20852 29892
rect 27264 29948 27328 29952
rect 27264 29892 27268 29948
rect 27268 29892 27324 29948
rect 27324 29892 27328 29948
rect 27264 29888 27328 29892
rect 27344 29948 27408 29952
rect 27344 29892 27348 29948
rect 27348 29892 27404 29948
rect 27404 29892 27408 29948
rect 27344 29888 27408 29892
rect 27424 29948 27488 29952
rect 27424 29892 27428 29948
rect 27428 29892 27484 29948
rect 27484 29892 27488 29948
rect 27424 29888 27488 29892
rect 27504 29948 27568 29952
rect 27504 29892 27508 29948
rect 27508 29892 27564 29948
rect 27564 29892 27568 29948
rect 27504 29888 27568 29892
rect 3758 29404 3822 29408
rect 3758 29348 3762 29404
rect 3762 29348 3818 29404
rect 3818 29348 3822 29404
rect 3758 29344 3822 29348
rect 3838 29404 3902 29408
rect 3838 29348 3842 29404
rect 3842 29348 3898 29404
rect 3898 29348 3902 29404
rect 3838 29344 3902 29348
rect 3918 29404 3982 29408
rect 3918 29348 3922 29404
rect 3922 29348 3978 29404
rect 3978 29348 3982 29404
rect 3918 29344 3982 29348
rect 3998 29404 4062 29408
rect 3998 29348 4002 29404
rect 4002 29348 4058 29404
rect 4058 29348 4062 29404
rect 3998 29344 4062 29348
rect 10474 29404 10538 29408
rect 10474 29348 10478 29404
rect 10478 29348 10534 29404
rect 10534 29348 10538 29404
rect 10474 29344 10538 29348
rect 10554 29404 10618 29408
rect 10554 29348 10558 29404
rect 10558 29348 10614 29404
rect 10614 29348 10618 29404
rect 10554 29344 10618 29348
rect 10634 29404 10698 29408
rect 10634 29348 10638 29404
rect 10638 29348 10694 29404
rect 10694 29348 10698 29404
rect 10634 29344 10698 29348
rect 10714 29404 10778 29408
rect 10714 29348 10718 29404
rect 10718 29348 10774 29404
rect 10774 29348 10778 29404
rect 10714 29344 10778 29348
rect 17190 29404 17254 29408
rect 17190 29348 17194 29404
rect 17194 29348 17250 29404
rect 17250 29348 17254 29404
rect 17190 29344 17254 29348
rect 17270 29404 17334 29408
rect 17270 29348 17274 29404
rect 17274 29348 17330 29404
rect 17330 29348 17334 29404
rect 17270 29344 17334 29348
rect 17350 29404 17414 29408
rect 17350 29348 17354 29404
rect 17354 29348 17410 29404
rect 17410 29348 17414 29404
rect 17350 29344 17414 29348
rect 17430 29404 17494 29408
rect 17430 29348 17434 29404
rect 17434 29348 17490 29404
rect 17490 29348 17494 29404
rect 17430 29344 17494 29348
rect 23906 29404 23970 29408
rect 23906 29348 23910 29404
rect 23910 29348 23966 29404
rect 23966 29348 23970 29404
rect 23906 29344 23970 29348
rect 23986 29404 24050 29408
rect 23986 29348 23990 29404
rect 23990 29348 24046 29404
rect 24046 29348 24050 29404
rect 23986 29344 24050 29348
rect 24066 29404 24130 29408
rect 24066 29348 24070 29404
rect 24070 29348 24126 29404
rect 24126 29348 24130 29404
rect 24066 29344 24130 29348
rect 24146 29404 24210 29408
rect 24146 29348 24150 29404
rect 24150 29348 24206 29404
rect 24206 29348 24210 29404
rect 24146 29344 24210 29348
rect 7116 28860 7180 28864
rect 7116 28804 7120 28860
rect 7120 28804 7176 28860
rect 7176 28804 7180 28860
rect 7116 28800 7180 28804
rect 7196 28860 7260 28864
rect 7196 28804 7200 28860
rect 7200 28804 7256 28860
rect 7256 28804 7260 28860
rect 7196 28800 7260 28804
rect 7276 28860 7340 28864
rect 7276 28804 7280 28860
rect 7280 28804 7336 28860
rect 7336 28804 7340 28860
rect 7276 28800 7340 28804
rect 7356 28860 7420 28864
rect 7356 28804 7360 28860
rect 7360 28804 7416 28860
rect 7416 28804 7420 28860
rect 7356 28800 7420 28804
rect 13832 28860 13896 28864
rect 13832 28804 13836 28860
rect 13836 28804 13892 28860
rect 13892 28804 13896 28860
rect 13832 28800 13896 28804
rect 13912 28860 13976 28864
rect 13912 28804 13916 28860
rect 13916 28804 13972 28860
rect 13972 28804 13976 28860
rect 13912 28800 13976 28804
rect 13992 28860 14056 28864
rect 13992 28804 13996 28860
rect 13996 28804 14052 28860
rect 14052 28804 14056 28860
rect 13992 28800 14056 28804
rect 14072 28860 14136 28864
rect 14072 28804 14076 28860
rect 14076 28804 14132 28860
rect 14132 28804 14136 28860
rect 14072 28800 14136 28804
rect 20548 28860 20612 28864
rect 20548 28804 20552 28860
rect 20552 28804 20608 28860
rect 20608 28804 20612 28860
rect 20548 28800 20612 28804
rect 20628 28860 20692 28864
rect 20628 28804 20632 28860
rect 20632 28804 20688 28860
rect 20688 28804 20692 28860
rect 20628 28800 20692 28804
rect 20708 28860 20772 28864
rect 20708 28804 20712 28860
rect 20712 28804 20768 28860
rect 20768 28804 20772 28860
rect 20708 28800 20772 28804
rect 20788 28860 20852 28864
rect 20788 28804 20792 28860
rect 20792 28804 20848 28860
rect 20848 28804 20852 28860
rect 20788 28800 20852 28804
rect 27264 28860 27328 28864
rect 27264 28804 27268 28860
rect 27268 28804 27324 28860
rect 27324 28804 27328 28860
rect 27264 28800 27328 28804
rect 27344 28860 27408 28864
rect 27344 28804 27348 28860
rect 27348 28804 27404 28860
rect 27404 28804 27408 28860
rect 27344 28800 27408 28804
rect 27424 28860 27488 28864
rect 27424 28804 27428 28860
rect 27428 28804 27484 28860
rect 27484 28804 27488 28860
rect 27424 28800 27488 28804
rect 27504 28860 27568 28864
rect 27504 28804 27508 28860
rect 27508 28804 27564 28860
rect 27564 28804 27568 28860
rect 27504 28800 27568 28804
rect 3758 28316 3822 28320
rect 3758 28260 3762 28316
rect 3762 28260 3818 28316
rect 3818 28260 3822 28316
rect 3758 28256 3822 28260
rect 3838 28316 3902 28320
rect 3838 28260 3842 28316
rect 3842 28260 3898 28316
rect 3898 28260 3902 28316
rect 3838 28256 3902 28260
rect 3918 28316 3982 28320
rect 3918 28260 3922 28316
rect 3922 28260 3978 28316
rect 3978 28260 3982 28316
rect 3918 28256 3982 28260
rect 3998 28316 4062 28320
rect 3998 28260 4002 28316
rect 4002 28260 4058 28316
rect 4058 28260 4062 28316
rect 3998 28256 4062 28260
rect 10474 28316 10538 28320
rect 10474 28260 10478 28316
rect 10478 28260 10534 28316
rect 10534 28260 10538 28316
rect 10474 28256 10538 28260
rect 10554 28316 10618 28320
rect 10554 28260 10558 28316
rect 10558 28260 10614 28316
rect 10614 28260 10618 28316
rect 10554 28256 10618 28260
rect 10634 28316 10698 28320
rect 10634 28260 10638 28316
rect 10638 28260 10694 28316
rect 10694 28260 10698 28316
rect 10634 28256 10698 28260
rect 10714 28316 10778 28320
rect 10714 28260 10718 28316
rect 10718 28260 10774 28316
rect 10774 28260 10778 28316
rect 10714 28256 10778 28260
rect 17190 28316 17254 28320
rect 17190 28260 17194 28316
rect 17194 28260 17250 28316
rect 17250 28260 17254 28316
rect 17190 28256 17254 28260
rect 17270 28316 17334 28320
rect 17270 28260 17274 28316
rect 17274 28260 17330 28316
rect 17330 28260 17334 28316
rect 17270 28256 17334 28260
rect 17350 28316 17414 28320
rect 17350 28260 17354 28316
rect 17354 28260 17410 28316
rect 17410 28260 17414 28316
rect 17350 28256 17414 28260
rect 17430 28316 17494 28320
rect 17430 28260 17434 28316
rect 17434 28260 17490 28316
rect 17490 28260 17494 28316
rect 17430 28256 17494 28260
rect 23906 28316 23970 28320
rect 23906 28260 23910 28316
rect 23910 28260 23966 28316
rect 23966 28260 23970 28316
rect 23906 28256 23970 28260
rect 23986 28316 24050 28320
rect 23986 28260 23990 28316
rect 23990 28260 24046 28316
rect 24046 28260 24050 28316
rect 23986 28256 24050 28260
rect 24066 28316 24130 28320
rect 24066 28260 24070 28316
rect 24070 28260 24126 28316
rect 24126 28260 24130 28316
rect 24066 28256 24130 28260
rect 24146 28316 24210 28320
rect 24146 28260 24150 28316
rect 24150 28260 24206 28316
rect 24206 28260 24210 28316
rect 24146 28256 24210 28260
rect 7116 27772 7180 27776
rect 7116 27716 7120 27772
rect 7120 27716 7176 27772
rect 7176 27716 7180 27772
rect 7116 27712 7180 27716
rect 7196 27772 7260 27776
rect 7196 27716 7200 27772
rect 7200 27716 7256 27772
rect 7256 27716 7260 27772
rect 7196 27712 7260 27716
rect 7276 27772 7340 27776
rect 7276 27716 7280 27772
rect 7280 27716 7336 27772
rect 7336 27716 7340 27772
rect 7276 27712 7340 27716
rect 7356 27772 7420 27776
rect 7356 27716 7360 27772
rect 7360 27716 7416 27772
rect 7416 27716 7420 27772
rect 7356 27712 7420 27716
rect 13832 27772 13896 27776
rect 13832 27716 13836 27772
rect 13836 27716 13892 27772
rect 13892 27716 13896 27772
rect 13832 27712 13896 27716
rect 13912 27772 13976 27776
rect 13912 27716 13916 27772
rect 13916 27716 13972 27772
rect 13972 27716 13976 27772
rect 13912 27712 13976 27716
rect 13992 27772 14056 27776
rect 13992 27716 13996 27772
rect 13996 27716 14052 27772
rect 14052 27716 14056 27772
rect 13992 27712 14056 27716
rect 14072 27772 14136 27776
rect 14072 27716 14076 27772
rect 14076 27716 14132 27772
rect 14132 27716 14136 27772
rect 14072 27712 14136 27716
rect 20548 27772 20612 27776
rect 20548 27716 20552 27772
rect 20552 27716 20608 27772
rect 20608 27716 20612 27772
rect 20548 27712 20612 27716
rect 20628 27772 20692 27776
rect 20628 27716 20632 27772
rect 20632 27716 20688 27772
rect 20688 27716 20692 27772
rect 20628 27712 20692 27716
rect 20708 27772 20772 27776
rect 20708 27716 20712 27772
rect 20712 27716 20768 27772
rect 20768 27716 20772 27772
rect 20708 27712 20772 27716
rect 20788 27772 20852 27776
rect 20788 27716 20792 27772
rect 20792 27716 20848 27772
rect 20848 27716 20852 27772
rect 20788 27712 20852 27716
rect 27264 27772 27328 27776
rect 27264 27716 27268 27772
rect 27268 27716 27324 27772
rect 27324 27716 27328 27772
rect 27264 27712 27328 27716
rect 27344 27772 27408 27776
rect 27344 27716 27348 27772
rect 27348 27716 27404 27772
rect 27404 27716 27408 27772
rect 27344 27712 27408 27716
rect 27424 27772 27488 27776
rect 27424 27716 27428 27772
rect 27428 27716 27484 27772
rect 27484 27716 27488 27772
rect 27424 27712 27488 27716
rect 27504 27772 27568 27776
rect 27504 27716 27508 27772
rect 27508 27716 27564 27772
rect 27564 27716 27568 27772
rect 27504 27712 27568 27716
rect 17724 27432 17788 27436
rect 17724 27376 17774 27432
rect 17774 27376 17788 27432
rect 17724 27372 17788 27376
rect 3758 27228 3822 27232
rect 3758 27172 3762 27228
rect 3762 27172 3818 27228
rect 3818 27172 3822 27228
rect 3758 27168 3822 27172
rect 3838 27228 3902 27232
rect 3838 27172 3842 27228
rect 3842 27172 3898 27228
rect 3898 27172 3902 27228
rect 3838 27168 3902 27172
rect 3918 27228 3982 27232
rect 3918 27172 3922 27228
rect 3922 27172 3978 27228
rect 3978 27172 3982 27228
rect 3918 27168 3982 27172
rect 3998 27228 4062 27232
rect 3998 27172 4002 27228
rect 4002 27172 4058 27228
rect 4058 27172 4062 27228
rect 3998 27168 4062 27172
rect 10474 27228 10538 27232
rect 10474 27172 10478 27228
rect 10478 27172 10534 27228
rect 10534 27172 10538 27228
rect 10474 27168 10538 27172
rect 10554 27228 10618 27232
rect 10554 27172 10558 27228
rect 10558 27172 10614 27228
rect 10614 27172 10618 27228
rect 10554 27168 10618 27172
rect 10634 27228 10698 27232
rect 10634 27172 10638 27228
rect 10638 27172 10694 27228
rect 10694 27172 10698 27228
rect 10634 27168 10698 27172
rect 10714 27228 10778 27232
rect 10714 27172 10718 27228
rect 10718 27172 10774 27228
rect 10774 27172 10778 27228
rect 10714 27168 10778 27172
rect 17190 27228 17254 27232
rect 17190 27172 17194 27228
rect 17194 27172 17250 27228
rect 17250 27172 17254 27228
rect 17190 27168 17254 27172
rect 17270 27228 17334 27232
rect 17270 27172 17274 27228
rect 17274 27172 17330 27228
rect 17330 27172 17334 27228
rect 17270 27168 17334 27172
rect 17350 27228 17414 27232
rect 17350 27172 17354 27228
rect 17354 27172 17410 27228
rect 17410 27172 17414 27228
rect 17350 27168 17414 27172
rect 17430 27228 17494 27232
rect 17430 27172 17434 27228
rect 17434 27172 17490 27228
rect 17490 27172 17494 27228
rect 17430 27168 17494 27172
rect 23906 27228 23970 27232
rect 23906 27172 23910 27228
rect 23910 27172 23966 27228
rect 23966 27172 23970 27228
rect 23906 27168 23970 27172
rect 23986 27228 24050 27232
rect 23986 27172 23990 27228
rect 23990 27172 24046 27228
rect 24046 27172 24050 27228
rect 23986 27168 24050 27172
rect 24066 27228 24130 27232
rect 24066 27172 24070 27228
rect 24070 27172 24126 27228
rect 24126 27172 24130 27228
rect 24066 27168 24130 27172
rect 24146 27228 24210 27232
rect 24146 27172 24150 27228
rect 24150 27172 24206 27228
rect 24206 27172 24210 27228
rect 24146 27168 24210 27172
rect 7116 26684 7180 26688
rect 7116 26628 7120 26684
rect 7120 26628 7176 26684
rect 7176 26628 7180 26684
rect 7116 26624 7180 26628
rect 7196 26684 7260 26688
rect 7196 26628 7200 26684
rect 7200 26628 7256 26684
rect 7256 26628 7260 26684
rect 7196 26624 7260 26628
rect 7276 26684 7340 26688
rect 7276 26628 7280 26684
rect 7280 26628 7336 26684
rect 7336 26628 7340 26684
rect 7276 26624 7340 26628
rect 7356 26684 7420 26688
rect 7356 26628 7360 26684
rect 7360 26628 7416 26684
rect 7416 26628 7420 26684
rect 7356 26624 7420 26628
rect 13832 26684 13896 26688
rect 13832 26628 13836 26684
rect 13836 26628 13892 26684
rect 13892 26628 13896 26684
rect 13832 26624 13896 26628
rect 13912 26684 13976 26688
rect 13912 26628 13916 26684
rect 13916 26628 13972 26684
rect 13972 26628 13976 26684
rect 13912 26624 13976 26628
rect 13992 26684 14056 26688
rect 13992 26628 13996 26684
rect 13996 26628 14052 26684
rect 14052 26628 14056 26684
rect 13992 26624 14056 26628
rect 14072 26684 14136 26688
rect 14072 26628 14076 26684
rect 14076 26628 14132 26684
rect 14132 26628 14136 26684
rect 14072 26624 14136 26628
rect 20548 26684 20612 26688
rect 20548 26628 20552 26684
rect 20552 26628 20608 26684
rect 20608 26628 20612 26684
rect 20548 26624 20612 26628
rect 20628 26684 20692 26688
rect 20628 26628 20632 26684
rect 20632 26628 20688 26684
rect 20688 26628 20692 26684
rect 20628 26624 20692 26628
rect 20708 26684 20772 26688
rect 20708 26628 20712 26684
rect 20712 26628 20768 26684
rect 20768 26628 20772 26684
rect 20708 26624 20772 26628
rect 20788 26684 20852 26688
rect 20788 26628 20792 26684
rect 20792 26628 20848 26684
rect 20848 26628 20852 26684
rect 20788 26624 20852 26628
rect 27264 26684 27328 26688
rect 27264 26628 27268 26684
rect 27268 26628 27324 26684
rect 27324 26628 27328 26684
rect 27264 26624 27328 26628
rect 27344 26684 27408 26688
rect 27344 26628 27348 26684
rect 27348 26628 27404 26684
rect 27404 26628 27408 26684
rect 27344 26624 27408 26628
rect 27424 26684 27488 26688
rect 27424 26628 27428 26684
rect 27428 26628 27484 26684
rect 27484 26628 27488 26684
rect 27424 26624 27488 26628
rect 27504 26684 27568 26688
rect 27504 26628 27508 26684
rect 27508 26628 27564 26684
rect 27564 26628 27568 26684
rect 27504 26624 27568 26628
rect 3758 26140 3822 26144
rect 3758 26084 3762 26140
rect 3762 26084 3818 26140
rect 3818 26084 3822 26140
rect 3758 26080 3822 26084
rect 3838 26140 3902 26144
rect 3838 26084 3842 26140
rect 3842 26084 3898 26140
rect 3898 26084 3902 26140
rect 3838 26080 3902 26084
rect 3918 26140 3982 26144
rect 3918 26084 3922 26140
rect 3922 26084 3978 26140
rect 3978 26084 3982 26140
rect 3918 26080 3982 26084
rect 3998 26140 4062 26144
rect 3998 26084 4002 26140
rect 4002 26084 4058 26140
rect 4058 26084 4062 26140
rect 3998 26080 4062 26084
rect 10474 26140 10538 26144
rect 10474 26084 10478 26140
rect 10478 26084 10534 26140
rect 10534 26084 10538 26140
rect 10474 26080 10538 26084
rect 10554 26140 10618 26144
rect 10554 26084 10558 26140
rect 10558 26084 10614 26140
rect 10614 26084 10618 26140
rect 10554 26080 10618 26084
rect 10634 26140 10698 26144
rect 10634 26084 10638 26140
rect 10638 26084 10694 26140
rect 10694 26084 10698 26140
rect 10634 26080 10698 26084
rect 10714 26140 10778 26144
rect 10714 26084 10718 26140
rect 10718 26084 10774 26140
rect 10774 26084 10778 26140
rect 10714 26080 10778 26084
rect 17190 26140 17254 26144
rect 17190 26084 17194 26140
rect 17194 26084 17250 26140
rect 17250 26084 17254 26140
rect 17190 26080 17254 26084
rect 17270 26140 17334 26144
rect 17270 26084 17274 26140
rect 17274 26084 17330 26140
rect 17330 26084 17334 26140
rect 17270 26080 17334 26084
rect 17350 26140 17414 26144
rect 17350 26084 17354 26140
rect 17354 26084 17410 26140
rect 17410 26084 17414 26140
rect 17350 26080 17414 26084
rect 17430 26140 17494 26144
rect 17430 26084 17434 26140
rect 17434 26084 17490 26140
rect 17490 26084 17494 26140
rect 17430 26080 17494 26084
rect 23906 26140 23970 26144
rect 23906 26084 23910 26140
rect 23910 26084 23966 26140
rect 23966 26084 23970 26140
rect 23906 26080 23970 26084
rect 23986 26140 24050 26144
rect 23986 26084 23990 26140
rect 23990 26084 24046 26140
rect 24046 26084 24050 26140
rect 23986 26080 24050 26084
rect 24066 26140 24130 26144
rect 24066 26084 24070 26140
rect 24070 26084 24126 26140
rect 24126 26084 24130 26140
rect 24066 26080 24130 26084
rect 24146 26140 24210 26144
rect 24146 26084 24150 26140
rect 24150 26084 24206 26140
rect 24206 26084 24210 26140
rect 24146 26080 24210 26084
rect 16620 25936 16684 25940
rect 16620 25880 16670 25936
rect 16670 25880 16684 25936
rect 16620 25876 16684 25880
rect 17724 25876 17788 25940
rect 17908 25664 17972 25668
rect 17908 25608 17958 25664
rect 17958 25608 17972 25664
rect 17908 25604 17972 25608
rect 7116 25596 7180 25600
rect 7116 25540 7120 25596
rect 7120 25540 7176 25596
rect 7176 25540 7180 25596
rect 7116 25536 7180 25540
rect 7196 25596 7260 25600
rect 7196 25540 7200 25596
rect 7200 25540 7256 25596
rect 7256 25540 7260 25596
rect 7196 25536 7260 25540
rect 7276 25596 7340 25600
rect 7276 25540 7280 25596
rect 7280 25540 7336 25596
rect 7336 25540 7340 25596
rect 7276 25536 7340 25540
rect 7356 25596 7420 25600
rect 7356 25540 7360 25596
rect 7360 25540 7416 25596
rect 7416 25540 7420 25596
rect 7356 25536 7420 25540
rect 13832 25596 13896 25600
rect 13832 25540 13836 25596
rect 13836 25540 13892 25596
rect 13892 25540 13896 25596
rect 13832 25536 13896 25540
rect 13912 25596 13976 25600
rect 13912 25540 13916 25596
rect 13916 25540 13972 25596
rect 13972 25540 13976 25596
rect 13912 25536 13976 25540
rect 13992 25596 14056 25600
rect 13992 25540 13996 25596
rect 13996 25540 14052 25596
rect 14052 25540 14056 25596
rect 13992 25536 14056 25540
rect 14072 25596 14136 25600
rect 14072 25540 14076 25596
rect 14076 25540 14132 25596
rect 14132 25540 14136 25596
rect 14072 25536 14136 25540
rect 20548 25596 20612 25600
rect 20548 25540 20552 25596
rect 20552 25540 20608 25596
rect 20608 25540 20612 25596
rect 20548 25536 20612 25540
rect 20628 25596 20692 25600
rect 20628 25540 20632 25596
rect 20632 25540 20688 25596
rect 20688 25540 20692 25596
rect 20628 25536 20692 25540
rect 20708 25596 20772 25600
rect 20708 25540 20712 25596
rect 20712 25540 20768 25596
rect 20768 25540 20772 25596
rect 20708 25536 20772 25540
rect 20788 25596 20852 25600
rect 20788 25540 20792 25596
rect 20792 25540 20848 25596
rect 20848 25540 20852 25596
rect 20788 25536 20852 25540
rect 27264 25596 27328 25600
rect 27264 25540 27268 25596
rect 27268 25540 27324 25596
rect 27324 25540 27328 25596
rect 27264 25536 27328 25540
rect 27344 25596 27408 25600
rect 27344 25540 27348 25596
rect 27348 25540 27404 25596
rect 27404 25540 27408 25596
rect 27344 25536 27408 25540
rect 27424 25596 27488 25600
rect 27424 25540 27428 25596
rect 27428 25540 27484 25596
rect 27484 25540 27488 25596
rect 27424 25536 27488 25540
rect 27504 25596 27568 25600
rect 27504 25540 27508 25596
rect 27508 25540 27564 25596
rect 27564 25540 27568 25596
rect 27504 25536 27568 25540
rect 3758 25052 3822 25056
rect 3758 24996 3762 25052
rect 3762 24996 3818 25052
rect 3818 24996 3822 25052
rect 3758 24992 3822 24996
rect 3838 25052 3902 25056
rect 3838 24996 3842 25052
rect 3842 24996 3898 25052
rect 3898 24996 3902 25052
rect 3838 24992 3902 24996
rect 3918 25052 3982 25056
rect 3918 24996 3922 25052
rect 3922 24996 3978 25052
rect 3978 24996 3982 25052
rect 3918 24992 3982 24996
rect 3998 25052 4062 25056
rect 3998 24996 4002 25052
rect 4002 24996 4058 25052
rect 4058 24996 4062 25052
rect 3998 24992 4062 24996
rect 10474 25052 10538 25056
rect 10474 24996 10478 25052
rect 10478 24996 10534 25052
rect 10534 24996 10538 25052
rect 10474 24992 10538 24996
rect 10554 25052 10618 25056
rect 10554 24996 10558 25052
rect 10558 24996 10614 25052
rect 10614 24996 10618 25052
rect 10554 24992 10618 24996
rect 10634 25052 10698 25056
rect 10634 24996 10638 25052
rect 10638 24996 10694 25052
rect 10694 24996 10698 25052
rect 10634 24992 10698 24996
rect 10714 25052 10778 25056
rect 10714 24996 10718 25052
rect 10718 24996 10774 25052
rect 10774 24996 10778 25052
rect 10714 24992 10778 24996
rect 17190 25052 17254 25056
rect 17190 24996 17194 25052
rect 17194 24996 17250 25052
rect 17250 24996 17254 25052
rect 17190 24992 17254 24996
rect 17270 25052 17334 25056
rect 17270 24996 17274 25052
rect 17274 24996 17330 25052
rect 17330 24996 17334 25052
rect 17270 24992 17334 24996
rect 17350 25052 17414 25056
rect 17350 24996 17354 25052
rect 17354 24996 17410 25052
rect 17410 24996 17414 25052
rect 17350 24992 17414 24996
rect 17430 25052 17494 25056
rect 17430 24996 17434 25052
rect 17434 24996 17490 25052
rect 17490 24996 17494 25052
rect 17430 24992 17494 24996
rect 23906 25052 23970 25056
rect 23906 24996 23910 25052
rect 23910 24996 23966 25052
rect 23966 24996 23970 25052
rect 23906 24992 23970 24996
rect 23986 25052 24050 25056
rect 23986 24996 23990 25052
rect 23990 24996 24046 25052
rect 24046 24996 24050 25052
rect 23986 24992 24050 24996
rect 24066 25052 24130 25056
rect 24066 24996 24070 25052
rect 24070 24996 24126 25052
rect 24126 24996 24130 25052
rect 24066 24992 24130 24996
rect 24146 25052 24210 25056
rect 24146 24996 24150 25052
rect 24150 24996 24206 25052
rect 24206 24996 24210 25052
rect 24146 24992 24210 24996
rect 7116 24508 7180 24512
rect 7116 24452 7120 24508
rect 7120 24452 7176 24508
rect 7176 24452 7180 24508
rect 7116 24448 7180 24452
rect 7196 24508 7260 24512
rect 7196 24452 7200 24508
rect 7200 24452 7256 24508
rect 7256 24452 7260 24508
rect 7196 24448 7260 24452
rect 7276 24508 7340 24512
rect 7276 24452 7280 24508
rect 7280 24452 7336 24508
rect 7336 24452 7340 24508
rect 7276 24448 7340 24452
rect 7356 24508 7420 24512
rect 7356 24452 7360 24508
rect 7360 24452 7416 24508
rect 7416 24452 7420 24508
rect 7356 24448 7420 24452
rect 13832 24508 13896 24512
rect 13832 24452 13836 24508
rect 13836 24452 13892 24508
rect 13892 24452 13896 24508
rect 13832 24448 13896 24452
rect 13912 24508 13976 24512
rect 13912 24452 13916 24508
rect 13916 24452 13972 24508
rect 13972 24452 13976 24508
rect 13912 24448 13976 24452
rect 13992 24508 14056 24512
rect 13992 24452 13996 24508
rect 13996 24452 14052 24508
rect 14052 24452 14056 24508
rect 13992 24448 14056 24452
rect 14072 24508 14136 24512
rect 14072 24452 14076 24508
rect 14076 24452 14132 24508
rect 14132 24452 14136 24508
rect 14072 24448 14136 24452
rect 20548 24508 20612 24512
rect 20548 24452 20552 24508
rect 20552 24452 20608 24508
rect 20608 24452 20612 24508
rect 20548 24448 20612 24452
rect 20628 24508 20692 24512
rect 20628 24452 20632 24508
rect 20632 24452 20688 24508
rect 20688 24452 20692 24508
rect 20628 24448 20692 24452
rect 20708 24508 20772 24512
rect 20708 24452 20712 24508
rect 20712 24452 20768 24508
rect 20768 24452 20772 24508
rect 20708 24448 20772 24452
rect 20788 24508 20852 24512
rect 20788 24452 20792 24508
rect 20792 24452 20848 24508
rect 20848 24452 20852 24508
rect 20788 24448 20852 24452
rect 27264 24508 27328 24512
rect 27264 24452 27268 24508
rect 27268 24452 27324 24508
rect 27324 24452 27328 24508
rect 27264 24448 27328 24452
rect 27344 24508 27408 24512
rect 27344 24452 27348 24508
rect 27348 24452 27404 24508
rect 27404 24452 27408 24508
rect 27344 24448 27408 24452
rect 27424 24508 27488 24512
rect 27424 24452 27428 24508
rect 27428 24452 27484 24508
rect 27484 24452 27488 24508
rect 27424 24448 27488 24452
rect 27504 24508 27568 24512
rect 27504 24452 27508 24508
rect 27508 24452 27564 24508
rect 27564 24452 27568 24508
rect 27504 24448 27568 24452
rect 3758 23964 3822 23968
rect 3758 23908 3762 23964
rect 3762 23908 3818 23964
rect 3818 23908 3822 23964
rect 3758 23904 3822 23908
rect 3838 23964 3902 23968
rect 3838 23908 3842 23964
rect 3842 23908 3898 23964
rect 3898 23908 3902 23964
rect 3838 23904 3902 23908
rect 3918 23964 3982 23968
rect 3918 23908 3922 23964
rect 3922 23908 3978 23964
rect 3978 23908 3982 23964
rect 3918 23904 3982 23908
rect 3998 23964 4062 23968
rect 3998 23908 4002 23964
rect 4002 23908 4058 23964
rect 4058 23908 4062 23964
rect 3998 23904 4062 23908
rect 10474 23964 10538 23968
rect 10474 23908 10478 23964
rect 10478 23908 10534 23964
rect 10534 23908 10538 23964
rect 10474 23904 10538 23908
rect 10554 23964 10618 23968
rect 10554 23908 10558 23964
rect 10558 23908 10614 23964
rect 10614 23908 10618 23964
rect 10554 23904 10618 23908
rect 10634 23964 10698 23968
rect 10634 23908 10638 23964
rect 10638 23908 10694 23964
rect 10694 23908 10698 23964
rect 10634 23904 10698 23908
rect 10714 23964 10778 23968
rect 10714 23908 10718 23964
rect 10718 23908 10774 23964
rect 10774 23908 10778 23964
rect 10714 23904 10778 23908
rect 17190 23964 17254 23968
rect 17190 23908 17194 23964
rect 17194 23908 17250 23964
rect 17250 23908 17254 23964
rect 17190 23904 17254 23908
rect 17270 23964 17334 23968
rect 17270 23908 17274 23964
rect 17274 23908 17330 23964
rect 17330 23908 17334 23964
rect 17270 23904 17334 23908
rect 17350 23964 17414 23968
rect 17350 23908 17354 23964
rect 17354 23908 17410 23964
rect 17410 23908 17414 23964
rect 17350 23904 17414 23908
rect 17430 23964 17494 23968
rect 17430 23908 17434 23964
rect 17434 23908 17490 23964
rect 17490 23908 17494 23964
rect 17430 23904 17494 23908
rect 23906 23964 23970 23968
rect 23906 23908 23910 23964
rect 23910 23908 23966 23964
rect 23966 23908 23970 23964
rect 23906 23904 23970 23908
rect 23986 23964 24050 23968
rect 23986 23908 23990 23964
rect 23990 23908 24046 23964
rect 24046 23908 24050 23964
rect 23986 23904 24050 23908
rect 24066 23964 24130 23968
rect 24066 23908 24070 23964
rect 24070 23908 24126 23964
rect 24126 23908 24130 23964
rect 24066 23904 24130 23908
rect 24146 23964 24210 23968
rect 24146 23908 24150 23964
rect 24150 23908 24206 23964
rect 24206 23908 24210 23964
rect 24146 23904 24210 23908
rect 17908 23564 17972 23628
rect 7116 23420 7180 23424
rect 7116 23364 7120 23420
rect 7120 23364 7176 23420
rect 7176 23364 7180 23420
rect 7116 23360 7180 23364
rect 7196 23420 7260 23424
rect 7196 23364 7200 23420
rect 7200 23364 7256 23420
rect 7256 23364 7260 23420
rect 7196 23360 7260 23364
rect 7276 23420 7340 23424
rect 7276 23364 7280 23420
rect 7280 23364 7336 23420
rect 7336 23364 7340 23420
rect 7276 23360 7340 23364
rect 7356 23420 7420 23424
rect 7356 23364 7360 23420
rect 7360 23364 7416 23420
rect 7416 23364 7420 23420
rect 7356 23360 7420 23364
rect 13832 23420 13896 23424
rect 13832 23364 13836 23420
rect 13836 23364 13892 23420
rect 13892 23364 13896 23420
rect 13832 23360 13896 23364
rect 13912 23420 13976 23424
rect 13912 23364 13916 23420
rect 13916 23364 13972 23420
rect 13972 23364 13976 23420
rect 13912 23360 13976 23364
rect 13992 23420 14056 23424
rect 13992 23364 13996 23420
rect 13996 23364 14052 23420
rect 14052 23364 14056 23420
rect 13992 23360 14056 23364
rect 14072 23420 14136 23424
rect 14072 23364 14076 23420
rect 14076 23364 14132 23420
rect 14132 23364 14136 23420
rect 14072 23360 14136 23364
rect 20548 23420 20612 23424
rect 20548 23364 20552 23420
rect 20552 23364 20608 23420
rect 20608 23364 20612 23420
rect 20548 23360 20612 23364
rect 20628 23420 20692 23424
rect 20628 23364 20632 23420
rect 20632 23364 20688 23420
rect 20688 23364 20692 23420
rect 20628 23360 20692 23364
rect 20708 23420 20772 23424
rect 20708 23364 20712 23420
rect 20712 23364 20768 23420
rect 20768 23364 20772 23420
rect 20708 23360 20772 23364
rect 20788 23420 20852 23424
rect 20788 23364 20792 23420
rect 20792 23364 20848 23420
rect 20848 23364 20852 23420
rect 20788 23360 20852 23364
rect 27264 23420 27328 23424
rect 27264 23364 27268 23420
rect 27268 23364 27324 23420
rect 27324 23364 27328 23420
rect 27264 23360 27328 23364
rect 27344 23420 27408 23424
rect 27344 23364 27348 23420
rect 27348 23364 27404 23420
rect 27404 23364 27408 23420
rect 27344 23360 27408 23364
rect 27424 23420 27488 23424
rect 27424 23364 27428 23420
rect 27428 23364 27484 23420
rect 27484 23364 27488 23420
rect 27424 23360 27488 23364
rect 27504 23420 27568 23424
rect 27504 23364 27508 23420
rect 27508 23364 27564 23420
rect 27564 23364 27568 23420
rect 27504 23360 27568 23364
rect 3758 22876 3822 22880
rect 3758 22820 3762 22876
rect 3762 22820 3818 22876
rect 3818 22820 3822 22876
rect 3758 22816 3822 22820
rect 3838 22876 3902 22880
rect 3838 22820 3842 22876
rect 3842 22820 3898 22876
rect 3898 22820 3902 22876
rect 3838 22816 3902 22820
rect 3918 22876 3982 22880
rect 3918 22820 3922 22876
rect 3922 22820 3978 22876
rect 3978 22820 3982 22876
rect 3918 22816 3982 22820
rect 3998 22876 4062 22880
rect 3998 22820 4002 22876
rect 4002 22820 4058 22876
rect 4058 22820 4062 22876
rect 3998 22816 4062 22820
rect 10474 22876 10538 22880
rect 10474 22820 10478 22876
rect 10478 22820 10534 22876
rect 10534 22820 10538 22876
rect 10474 22816 10538 22820
rect 10554 22876 10618 22880
rect 10554 22820 10558 22876
rect 10558 22820 10614 22876
rect 10614 22820 10618 22876
rect 10554 22816 10618 22820
rect 10634 22876 10698 22880
rect 10634 22820 10638 22876
rect 10638 22820 10694 22876
rect 10694 22820 10698 22876
rect 10634 22816 10698 22820
rect 10714 22876 10778 22880
rect 10714 22820 10718 22876
rect 10718 22820 10774 22876
rect 10774 22820 10778 22876
rect 10714 22816 10778 22820
rect 17190 22876 17254 22880
rect 17190 22820 17194 22876
rect 17194 22820 17250 22876
rect 17250 22820 17254 22876
rect 17190 22816 17254 22820
rect 17270 22876 17334 22880
rect 17270 22820 17274 22876
rect 17274 22820 17330 22876
rect 17330 22820 17334 22876
rect 17270 22816 17334 22820
rect 17350 22876 17414 22880
rect 17350 22820 17354 22876
rect 17354 22820 17410 22876
rect 17410 22820 17414 22876
rect 17350 22816 17414 22820
rect 17430 22876 17494 22880
rect 17430 22820 17434 22876
rect 17434 22820 17490 22876
rect 17490 22820 17494 22876
rect 17430 22816 17494 22820
rect 23906 22876 23970 22880
rect 23906 22820 23910 22876
rect 23910 22820 23966 22876
rect 23966 22820 23970 22876
rect 23906 22816 23970 22820
rect 23986 22876 24050 22880
rect 23986 22820 23990 22876
rect 23990 22820 24046 22876
rect 24046 22820 24050 22876
rect 23986 22816 24050 22820
rect 24066 22876 24130 22880
rect 24066 22820 24070 22876
rect 24070 22820 24126 22876
rect 24126 22820 24130 22876
rect 24066 22816 24130 22820
rect 24146 22876 24210 22880
rect 24146 22820 24150 22876
rect 24150 22820 24206 22876
rect 24206 22820 24210 22876
rect 24146 22816 24210 22820
rect 7116 22332 7180 22336
rect 7116 22276 7120 22332
rect 7120 22276 7176 22332
rect 7176 22276 7180 22332
rect 7116 22272 7180 22276
rect 7196 22332 7260 22336
rect 7196 22276 7200 22332
rect 7200 22276 7256 22332
rect 7256 22276 7260 22332
rect 7196 22272 7260 22276
rect 7276 22332 7340 22336
rect 7276 22276 7280 22332
rect 7280 22276 7336 22332
rect 7336 22276 7340 22332
rect 7276 22272 7340 22276
rect 7356 22332 7420 22336
rect 7356 22276 7360 22332
rect 7360 22276 7416 22332
rect 7416 22276 7420 22332
rect 7356 22272 7420 22276
rect 13832 22332 13896 22336
rect 13832 22276 13836 22332
rect 13836 22276 13892 22332
rect 13892 22276 13896 22332
rect 13832 22272 13896 22276
rect 13912 22332 13976 22336
rect 13912 22276 13916 22332
rect 13916 22276 13972 22332
rect 13972 22276 13976 22332
rect 13912 22272 13976 22276
rect 13992 22332 14056 22336
rect 13992 22276 13996 22332
rect 13996 22276 14052 22332
rect 14052 22276 14056 22332
rect 13992 22272 14056 22276
rect 14072 22332 14136 22336
rect 14072 22276 14076 22332
rect 14076 22276 14132 22332
rect 14132 22276 14136 22332
rect 14072 22272 14136 22276
rect 20548 22332 20612 22336
rect 20548 22276 20552 22332
rect 20552 22276 20608 22332
rect 20608 22276 20612 22332
rect 20548 22272 20612 22276
rect 20628 22332 20692 22336
rect 20628 22276 20632 22332
rect 20632 22276 20688 22332
rect 20688 22276 20692 22332
rect 20628 22272 20692 22276
rect 20708 22332 20772 22336
rect 20708 22276 20712 22332
rect 20712 22276 20768 22332
rect 20768 22276 20772 22332
rect 20708 22272 20772 22276
rect 20788 22332 20852 22336
rect 20788 22276 20792 22332
rect 20792 22276 20848 22332
rect 20848 22276 20852 22332
rect 20788 22272 20852 22276
rect 27264 22332 27328 22336
rect 27264 22276 27268 22332
rect 27268 22276 27324 22332
rect 27324 22276 27328 22332
rect 27264 22272 27328 22276
rect 27344 22332 27408 22336
rect 27344 22276 27348 22332
rect 27348 22276 27404 22332
rect 27404 22276 27408 22332
rect 27344 22272 27408 22276
rect 27424 22332 27488 22336
rect 27424 22276 27428 22332
rect 27428 22276 27484 22332
rect 27484 22276 27488 22332
rect 27424 22272 27488 22276
rect 27504 22332 27568 22336
rect 27504 22276 27508 22332
rect 27508 22276 27564 22332
rect 27564 22276 27568 22332
rect 27504 22272 27568 22276
rect 11100 22068 11164 22132
rect 5212 21932 5276 21996
rect 11284 21932 11348 21996
rect 3758 21788 3822 21792
rect 3758 21732 3762 21788
rect 3762 21732 3818 21788
rect 3818 21732 3822 21788
rect 3758 21728 3822 21732
rect 3838 21788 3902 21792
rect 3838 21732 3842 21788
rect 3842 21732 3898 21788
rect 3898 21732 3902 21788
rect 3838 21728 3902 21732
rect 3918 21788 3982 21792
rect 3918 21732 3922 21788
rect 3922 21732 3978 21788
rect 3978 21732 3982 21788
rect 3918 21728 3982 21732
rect 3998 21788 4062 21792
rect 3998 21732 4002 21788
rect 4002 21732 4058 21788
rect 4058 21732 4062 21788
rect 3998 21728 4062 21732
rect 10474 21788 10538 21792
rect 10474 21732 10478 21788
rect 10478 21732 10534 21788
rect 10534 21732 10538 21788
rect 10474 21728 10538 21732
rect 10554 21788 10618 21792
rect 10554 21732 10558 21788
rect 10558 21732 10614 21788
rect 10614 21732 10618 21788
rect 10554 21728 10618 21732
rect 10634 21788 10698 21792
rect 10634 21732 10638 21788
rect 10638 21732 10694 21788
rect 10694 21732 10698 21788
rect 10634 21728 10698 21732
rect 10714 21788 10778 21792
rect 10714 21732 10718 21788
rect 10718 21732 10774 21788
rect 10774 21732 10778 21788
rect 10714 21728 10778 21732
rect 17190 21788 17254 21792
rect 17190 21732 17194 21788
rect 17194 21732 17250 21788
rect 17250 21732 17254 21788
rect 17190 21728 17254 21732
rect 17270 21788 17334 21792
rect 17270 21732 17274 21788
rect 17274 21732 17330 21788
rect 17330 21732 17334 21788
rect 17270 21728 17334 21732
rect 17350 21788 17414 21792
rect 17350 21732 17354 21788
rect 17354 21732 17410 21788
rect 17410 21732 17414 21788
rect 17350 21728 17414 21732
rect 17430 21788 17494 21792
rect 17430 21732 17434 21788
rect 17434 21732 17490 21788
rect 17490 21732 17494 21788
rect 17430 21728 17494 21732
rect 23906 21788 23970 21792
rect 23906 21732 23910 21788
rect 23910 21732 23966 21788
rect 23966 21732 23970 21788
rect 23906 21728 23970 21732
rect 23986 21788 24050 21792
rect 23986 21732 23990 21788
rect 23990 21732 24046 21788
rect 24046 21732 24050 21788
rect 23986 21728 24050 21732
rect 24066 21788 24130 21792
rect 24066 21732 24070 21788
rect 24070 21732 24126 21788
rect 24126 21732 24130 21788
rect 24066 21728 24130 21732
rect 24146 21788 24210 21792
rect 24146 21732 24150 21788
rect 24150 21732 24206 21788
rect 24206 21732 24210 21788
rect 24146 21728 24210 21732
rect 7116 21244 7180 21248
rect 7116 21188 7120 21244
rect 7120 21188 7176 21244
rect 7176 21188 7180 21244
rect 7116 21184 7180 21188
rect 7196 21244 7260 21248
rect 7196 21188 7200 21244
rect 7200 21188 7256 21244
rect 7256 21188 7260 21244
rect 7196 21184 7260 21188
rect 7276 21244 7340 21248
rect 7276 21188 7280 21244
rect 7280 21188 7336 21244
rect 7336 21188 7340 21244
rect 7276 21184 7340 21188
rect 7356 21244 7420 21248
rect 7356 21188 7360 21244
rect 7360 21188 7416 21244
rect 7416 21188 7420 21244
rect 7356 21184 7420 21188
rect 13832 21244 13896 21248
rect 13832 21188 13836 21244
rect 13836 21188 13892 21244
rect 13892 21188 13896 21244
rect 13832 21184 13896 21188
rect 13912 21244 13976 21248
rect 13912 21188 13916 21244
rect 13916 21188 13972 21244
rect 13972 21188 13976 21244
rect 13912 21184 13976 21188
rect 13992 21244 14056 21248
rect 13992 21188 13996 21244
rect 13996 21188 14052 21244
rect 14052 21188 14056 21244
rect 13992 21184 14056 21188
rect 14072 21244 14136 21248
rect 14072 21188 14076 21244
rect 14076 21188 14132 21244
rect 14132 21188 14136 21244
rect 14072 21184 14136 21188
rect 20548 21244 20612 21248
rect 20548 21188 20552 21244
rect 20552 21188 20608 21244
rect 20608 21188 20612 21244
rect 20548 21184 20612 21188
rect 20628 21244 20692 21248
rect 20628 21188 20632 21244
rect 20632 21188 20688 21244
rect 20688 21188 20692 21244
rect 20628 21184 20692 21188
rect 20708 21244 20772 21248
rect 20708 21188 20712 21244
rect 20712 21188 20768 21244
rect 20768 21188 20772 21244
rect 20708 21184 20772 21188
rect 20788 21244 20852 21248
rect 20788 21188 20792 21244
rect 20792 21188 20848 21244
rect 20848 21188 20852 21244
rect 20788 21184 20852 21188
rect 27264 21244 27328 21248
rect 27264 21188 27268 21244
rect 27268 21188 27324 21244
rect 27324 21188 27328 21244
rect 27264 21184 27328 21188
rect 27344 21244 27408 21248
rect 27344 21188 27348 21244
rect 27348 21188 27404 21244
rect 27404 21188 27408 21244
rect 27344 21184 27408 21188
rect 27424 21244 27488 21248
rect 27424 21188 27428 21244
rect 27428 21188 27484 21244
rect 27484 21188 27488 21244
rect 27424 21184 27488 21188
rect 27504 21244 27568 21248
rect 27504 21188 27508 21244
rect 27508 21188 27564 21244
rect 27564 21188 27568 21244
rect 27504 21184 27568 21188
rect 3758 20700 3822 20704
rect 3758 20644 3762 20700
rect 3762 20644 3818 20700
rect 3818 20644 3822 20700
rect 3758 20640 3822 20644
rect 3838 20700 3902 20704
rect 3838 20644 3842 20700
rect 3842 20644 3898 20700
rect 3898 20644 3902 20700
rect 3838 20640 3902 20644
rect 3918 20700 3982 20704
rect 3918 20644 3922 20700
rect 3922 20644 3978 20700
rect 3978 20644 3982 20700
rect 3918 20640 3982 20644
rect 3998 20700 4062 20704
rect 3998 20644 4002 20700
rect 4002 20644 4058 20700
rect 4058 20644 4062 20700
rect 3998 20640 4062 20644
rect 10474 20700 10538 20704
rect 10474 20644 10478 20700
rect 10478 20644 10534 20700
rect 10534 20644 10538 20700
rect 10474 20640 10538 20644
rect 10554 20700 10618 20704
rect 10554 20644 10558 20700
rect 10558 20644 10614 20700
rect 10614 20644 10618 20700
rect 10554 20640 10618 20644
rect 10634 20700 10698 20704
rect 10634 20644 10638 20700
rect 10638 20644 10694 20700
rect 10694 20644 10698 20700
rect 10634 20640 10698 20644
rect 10714 20700 10778 20704
rect 10714 20644 10718 20700
rect 10718 20644 10774 20700
rect 10774 20644 10778 20700
rect 10714 20640 10778 20644
rect 17190 20700 17254 20704
rect 17190 20644 17194 20700
rect 17194 20644 17250 20700
rect 17250 20644 17254 20700
rect 17190 20640 17254 20644
rect 17270 20700 17334 20704
rect 17270 20644 17274 20700
rect 17274 20644 17330 20700
rect 17330 20644 17334 20700
rect 17270 20640 17334 20644
rect 17350 20700 17414 20704
rect 17350 20644 17354 20700
rect 17354 20644 17410 20700
rect 17410 20644 17414 20700
rect 17350 20640 17414 20644
rect 17430 20700 17494 20704
rect 17430 20644 17434 20700
rect 17434 20644 17490 20700
rect 17490 20644 17494 20700
rect 17430 20640 17494 20644
rect 23906 20700 23970 20704
rect 23906 20644 23910 20700
rect 23910 20644 23966 20700
rect 23966 20644 23970 20700
rect 23906 20640 23970 20644
rect 23986 20700 24050 20704
rect 23986 20644 23990 20700
rect 23990 20644 24046 20700
rect 24046 20644 24050 20700
rect 23986 20640 24050 20644
rect 24066 20700 24130 20704
rect 24066 20644 24070 20700
rect 24070 20644 24126 20700
rect 24126 20644 24130 20700
rect 24066 20640 24130 20644
rect 24146 20700 24210 20704
rect 24146 20644 24150 20700
rect 24150 20644 24206 20700
rect 24206 20644 24210 20700
rect 24146 20640 24210 20644
rect 7116 20156 7180 20160
rect 7116 20100 7120 20156
rect 7120 20100 7176 20156
rect 7176 20100 7180 20156
rect 7116 20096 7180 20100
rect 7196 20156 7260 20160
rect 7196 20100 7200 20156
rect 7200 20100 7256 20156
rect 7256 20100 7260 20156
rect 7196 20096 7260 20100
rect 7276 20156 7340 20160
rect 7276 20100 7280 20156
rect 7280 20100 7336 20156
rect 7336 20100 7340 20156
rect 7276 20096 7340 20100
rect 7356 20156 7420 20160
rect 7356 20100 7360 20156
rect 7360 20100 7416 20156
rect 7416 20100 7420 20156
rect 7356 20096 7420 20100
rect 13832 20156 13896 20160
rect 13832 20100 13836 20156
rect 13836 20100 13892 20156
rect 13892 20100 13896 20156
rect 13832 20096 13896 20100
rect 13912 20156 13976 20160
rect 13912 20100 13916 20156
rect 13916 20100 13972 20156
rect 13972 20100 13976 20156
rect 13912 20096 13976 20100
rect 13992 20156 14056 20160
rect 13992 20100 13996 20156
rect 13996 20100 14052 20156
rect 14052 20100 14056 20156
rect 13992 20096 14056 20100
rect 14072 20156 14136 20160
rect 14072 20100 14076 20156
rect 14076 20100 14132 20156
rect 14132 20100 14136 20156
rect 14072 20096 14136 20100
rect 20548 20156 20612 20160
rect 20548 20100 20552 20156
rect 20552 20100 20608 20156
rect 20608 20100 20612 20156
rect 20548 20096 20612 20100
rect 20628 20156 20692 20160
rect 20628 20100 20632 20156
rect 20632 20100 20688 20156
rect 20688 20100 20692 20156
rect 20628 20096 20692 20100
rect 20708 20156 20772 20160
rect 20708 20100 20712 20156
rect 20712 20100 20768 20156
rect 20768 20100 20772 20156
rect 20708 20096 20772 20100
rect 20788 20156 20852 20160
rect 20788 20100 20792 20156
rect 20792 20100 20848 20156
rect 20848 20100 20852 20156
rect 20788 20096 20852 20100
rect 27264 20156 27328 20160
rect 27264 20100 27268 20156
rect 27268 20100 27324 20156
rect 27324 20100 27328 20156
rect 27264 20096 27328 20100
rect 27344 20156 27408 20160
rect 27344 20100 27348 20156
rect 27348 20100 27404 20156
rect 27404 20100 27408 20156
rect 27344 20096 27408 20100
rect 27424 20156 27488 20160
rect 27424 20100 27428 20156
rect 27428 20100 27484 20156
rect 27484 20100 27488 20156
rect 27424 20096 27488 20100
rect 27504 20156 27568 20160
rect 27504 20100 27508 20156
rect 27508 20100 27564 20156
rect 27564 20100 27568 20156
rect 27504 20096 27568 20100
rect 16068 19756 16132 19820
rect 3758 19612 3822 19616
rect 3758 19556 3762 19612
rect 3762 19556 3818 19612
rect 3818 19556 3822 19612
rect 3758 19552 3822 19556
rect 3838 19612 3902 19616
rect 3838 19556 3842 19612
rect 3842 19556 3898 19612
rect 3898 19556 3902 19612
rect 3838 19552 3902 19556
rect 3918 19612 3982 19616
rect 3918 19556 3922 19612
rect 3922 19556 3978 19612
rect 3978 19556 3982 19612
rect 3918 19552 3982 19556
rect 3998 19612 4062 19616
rect 3998 19556 4002 19612
rect 4002 19556 4058 19612
rect 4058 19556 4062 19612
rect 3998 19552 4062 19556
rect 10474 19612 10538 19616
rect 10474 19556 10478 19612
rect 10478 19556 10534 19612
rect 10534 19556 10538 19612
rect 10474 19552 10538 19556
rect 10554 19612 10618 19616
rect 10554 19556 10558 19612
rect 10558 19556 10614 19612
rect 10614 19556 10618 19612
rect 10554 19552 10618 19556
rect 10634 19612 10698 19616
rect 10634 19556 10638 19612
rect 10638 19556 10694 19612
rect 10694 19556 10698 19612
rect 10634 19552 10698 19556
rect 10714 19612 10778 19616
rect 10714 19556 10718 19612
rect 10718 19556 10774 19612
rect 10774 19556 10778 19612
rect 10714 19552 10778 19556
rect 17190 19612 17254 19616
rect 17190 19556 17194 19612
rect 17194 19556 17250 19612
rect 17250 19556 17254 19612
rect 17190 19552 17254 19556
rect 17270 19612 17334 19616
rect 17270 19556 17274 19612
rect 17274 19556 17330 19612
rect 17330 19556 17334 19612
rect 17270 19552 17334 19556
rect 17350 19612 17414 19616
rect 17350 19556 17354 19612
rect 17354 19556 17410 19612
rect 17410 19556 17414 19612
rect 17350 19552 17414 19556
rect 17430 19612 17494 19616
rect 17430 19556 17434 19612
rect 17434 19556 17490 19612
rect 17490 19556 17494 19612
rect 17430 19552 17494 19556
rect 23906 19612 23970 19616
rect 23906 19556 23910 19612
rect 23910 19556 23966 19612
rect 23966 19556 23970 19612
rect 23906 19552 23970 19556
rect 23986 19612 24050 19616
rect 23986 19556 23990 19612
rect 23990 19556 24046 19612
rect 24046 19556 24050 19612
rect 23986 19552 24050 19556
rect 24066 19612 24130 19616
rect 24066 19556 24070 19612
rect 24070 19556 24126 19612
rect 24126 19556 24130 19612
rect 24066 19552 24130 19556
rect 24146 19612 24210 19616
rect 24146 19556 24150 19612
rect 24150 19556 24206 19612
rect 24206 19556 24210 19612
rect 24146 19552 24210 19556
rect 12572 19348 12636 19412
rect 16620 19212 16684 19276
rect 17724 19212 17788 19276
rect 7116 19068 7180 19072
rect 7116 19012 7120 19068
rect 7120 19012 7176 19068
rect 7176 19012 7180 19068
rect 7116 19008 7180 19012
rect 7196 19068 7260 19072
rect 7196 19012 7200 19068
rect 7200 19012 7256 19068
rect 7256 19012 7260 19068
rect 7196 19008 7260 19012
rect 7276 19068 7340 19072
rect 7276 19012 7280 19068
rect 7280 19012 7336 19068
rect 7336 19012 7340 19068
rect 7276 19008 7340 19012
rect 7356 19068 7420 19072
rect 7356 19012 7360 19068
rect 7360 19012 7416 19068
rect 7416 19012 7420 19068
rect 7356 19008 7420 19012
rect 13832 19068 13896 19072
rect 13832 19012 13836 19068
rect 13836 19012 13892 19068
rect 13892 19012 13896 19068
rect 13832 19008 13896 19012
rect 13912 19068 13976 19072
rect 13912 19012 13916 19068
rect 13916 19012 13972 19068
rect 13972 19012 13976 19068
rect 13912 19008 13976 19012
rect 13992 19068 14056 19072
rect 13992 19012 13996 19068
rect 13996 19012 14052 19068
rect 14052 19012 14056 19068
rect 13992 19008 14056 19012
rect 14072 19068 14136 19072
rect 14072 19012 14076 19068
rect 14076 19012 14132 19068
rect 14132 19012 14136 19068
rect 14072 19008 14136 19012
rect 20548 19068 20612 19072
rect 20548 19012 20552 19068
rect 20552 19012 20608 19068
rect 20608 19012 20612 19068
rect 20548 19008 20612 19012
rect 20628 19068 20692 19072
rect 20628 19012 20632 19068
rect 20632 19012 20688 19068
rect 20688 19012 20692 19068
rect 20628 19008 20692 19012
rect 20708 19068 20772 19072
rect 20708 19012 20712 19068
rect 20712 19012 20768 19068
rect 20768 19012 20772 19068
rect 20708 19008 20772 19012
rect 20788 19068 20852 19072
rect 20788 19012 20792 19068
rect 20792 19012 20848 19068
rect 20848 19012 20852 19068
rect 20788 19008 20852 19012
rect 27264 19068 27328 19072
rect 27264 19012 27268 19068
rect 27268 19012 27324 19068
rect 27324 19012 27328 19068
rect 27264 19008 27328 19012
rect 27344 19068 27408 19072
rect 27344 19012 27348 19068
rect 27348 19012 27404 19068
rect 27404 19012 27408 19068
rect 27344 19008 27408 19012
rect 27424 19068 27488 19072
rect 27424 19012 27428 19068
rect 27428 19012 27484 19068
rect 27484 19012 27488 19068
rect 27424 19008 27488 19012
rect 27504 19068 27568 19072
rect 27504 19012 27508 19068
rect 27508 19012 27564 19068
rect 27564 19012 27568 19068
rect 27504 19008 27568 19012
rect 3758 18524 3822 18528
rect 3758 18468 3762 18524
rect 3762 18468 3818 18524
rect 3818 18468 3822 18524
rect 3758 18464 3822 18468
rect 3838 18524 3902 18528
rect 3838 18468 3842 18524
rect 3842 18468 3898 18524
rect 3898 18468 3902 18524
rect 3838 18464 3902 18468
rect 3918 18524 3982 18528
rect 3918 18468 3922 18524
rect 3922 18468 3978 18524
rect 3978 18468 3982 18524
rect 3918 18464 3982 18468
rect 3998 18524 4062 18528
rect 3998 18468 4002 18524
rect 4002 18468 4058 18524
rect 4058 18468 4062 18524
rect 3998 18464 4062 18468
rect 10474 18524 10538 18528
rect 10474 18468 10478 18524
rect 10478 18468 10534 18524
rect 10534 18468 10538 18524
rect 10474 18464 10538 18468
rect 10554 18524 10618 18528
rect 10554 18468 10558 18524
rect 10558 18468 10614 18524
rect 10614 18468 10618 18524
rect 10554 18464 10618 18468
rect 10634 18524 10698 18528
rect 10634 18468 10638 18524
rect 10638 18468 10694 18524
rect 10694 18468 10698 18524
rect 10634 18464 10698 18468
rect 10714 18524 10778 18528
rect 10714 18468 10718 18524
rect 10718 18468 10774 18524
rect 10774 18468 10778 18524
rect 10714 18464 10778 18468
rect 17190 18524 17254 18528
rect 17190 18468 17194 18524
rect 17194 18468 17250 18524
rect 17250 18468 17254 18524
rect 17190 18464 17254 18468
rect 17270 18524 17334 18528
rect 17270 18468 17274 18524
rect 17274 18468 17330 18524
rect 17330 18468 17334 18524
rect 17270 18464 17334 18468
rect 17350 18524 17414 18528
rect 17350 18468 17354 18524
rect 17354 18468 17410 18524
rect 17410 18468 17414 18524
rect 17350 18464 17414 18468
rect 17430 18524 17494 18528
rect 17430 18468 17434 18524
rect 17434 18468 17490 18524
rect 17490 18468 17494 18524
rect 17430 18464 17494 18468
rect 23906 18524 23970 18528
rect 23906 18468 23910 18524
rect 23910 18468 23966 18524
rect 23966 18468 23970 18524
rect 23906 18464 23970 18468
rect 23986 18524 24050 18528
rect 23986 18468 23990 18524
rect 23990 18468 24046 18524
rect 24046 18468 24050 18524
rect 23986 18464 24050 18468
rect 24066 18524 24130 18528
rect 24066 18468 24070 18524
rect 24070 18468 24126 18524
rect 24126 18468 24130 18524
rect 24066 18464 24130 18468
rect 24146 18524 24210 18528
rect 24146 18468 24150 18524
rect 24150 18468 24206 18524
rect 24206 18468 24210 18524
rect 24146 18464 24210 18468
rect 17908 18260 17972 18324
rect 7116 17980 7180 17984
rect 7116 17924 7120 17980
rect 7120 17924 7176 17980
rect 7176 17924 7180 17980
rect 7116 17920 7180 17924
rect 7196 17980 7260 17984
rect 7196 17924 7200 17980
rect 7200 17924 7256 17980
rect 7256 17924 7260 17980
rect 7196 17920 7260 17924
rect 7276 17980 7340 17984
rect 7276 17924 7280 17980
rect 7280 17924 7336 17980
rect 7336 17924 7340 17980
rect 7276 17920 7340 17924
rect 7356 17980 7420 17984
rect 7356 17924 7360 17980
rect 7360 17924 7416 17980
rect 7416 17924 7420 17980
rect 7356 17920 7420 17924
rect 13832 17980 13896 17984
rect 13832 17924 13836 17980
rect 13836 17924 13892 17980
rect 13892 17924 13896 17980
rect 13832 17920 13896 17924
rect 13912 17980 13976 17984
rect 13912 17924 13916 17980
rect 13916 17924 13972 17980
rect 13972 17924 13976 17980
rect 13912 17920 13976 17924
rect 13992 17980 14056 17984
rect 13992 17924 13996 17980
rect 13996 17924 14052 17980
rect 14052 17924 14056 17980
rect 13992 17920 14056 17924
rect 14072 17980 14136 17984
rect 14072 17924 14076 17980
rect 14076 17924 14132 17980
rect 14132 17924 14136 17980
rect 14072 17920 14136 17924
rect 20548 17980 20612 17984
rect 20548 17924 20552 17980
rect 20552 17924 20608 17980
rect 20608 17924 20612 17980
rect 20548 17920 20612 17924
rect 20628 17980 20692 17984
rect 20628 17924 20632 17980
rect 20632 17924 20688 17980
rect 20688 17924 20692 17980
rect 20628 17920 20692 17924
rect 20708 17980 20772 17984
rect 20708 17924 20712 17980
rect 20712 17924 20768 17980
rect 20768 17924 20772 17980
rect 20708 17920 20772 17924
rect 20788 17980 20852 17984
rect 20788 17924 20792 17980
rect 20792 17924 20848 17980
rect 20848 17924 20852 17980
rect 20788 17920 20852 17924
rect 27264 17980 27328 17984
rect 27264 17924 27268 17980
rect 27268 17924 27324 17980
rect 27324 17924 27328 17980
rect 27264 17920 27328 17924
rect 27344 17980 27408 17984
rect 27344 17924 27348 17980
rect 27348 17924 27404 17980
rect 27404 17924 27408 17980
rect 27344 17920 27408 17924
rect 27424 17980 27488 17984
rect 27424 17924 27428 17980
rect 27428 17924 27484 17980
rect 27484 17924 27488 17980
rect 27424 17920 27488 17924
rect 27504 17980 27568 17984
rect 27504 17924 27508 17980
rect 27508 17924 27564 17980
rect 27564 17924 27568 17980
rect 27504 17920 27568 17924
rect 11100 17852 11164 17916
rect 3758 17436 3822 17440
rect 3758 17380 3762 17436
rect 3762 17380 3818 17436
rect 3818 17380 3822 17436
rect 3758 17376 3822 17380
rect 3838 17436 3902 17440
rect 3838 17380 3842 17436
rect 3842 17380 3898 17436
rect 3898 17380 3902 17436
rect 3838 17376 3902 17380
rect 3918 17436 3982 17440
rect 3918 17380 3922 17436
rect 3922 17380 3978 17436
rect 3978 17380 3982 17436
rect 3918 17376 3982 17380
rect 3998 17436 4062 17440
rect 3998 17380 4002 17436
rect 4002 17380 4058 17436
rect 4058 17380 4062 17436
rect 3998 17376 4062 17380
rect 10474 17436 10538 17440
rect 10474 17380 10478 17436
rect 10478 17380 10534 17436
rect 10534 17380 10538 17436
rect 10474 17376 10538 17380
rect 10554 17436 10618 17440
rect 10554 17380 10558 17436
rect 10558 17380 10614 17436
rect 10614 17380 10618 17436
rect 10554 17376 10618 17380
rect 10634 17436 10698 17440
rect 10634 17380 10638 17436
rect 10638 17380 10694 17436
rect 10694 17380 10698 17436
rect 10634 17376 10698 17380
rect 10714 17436 10778 17440
rect 10714 17380 10718 17436
rect 10718 17380 10774 17436
rect 10774 17380 10778 17436
rect 10714 17376 10778 17380
rect 17190 17436 17254 17440
rect 17190 17380 17194 17436
rect 17194 17380 17250 17436
rect 17250 17380 17254 17436
rect 17190 17376 17254 17380
rect 17270 17436 17334 17440
rect 17270 17380 17274 17436
rect 17274 17380 17330 17436
rect 17330 17380 17334 17436
rect 17270 17376 17334 17380
rect 17350 17436 17414 17440
rect 17350 17380 17354 17436
rect 17354 17380 17410 17436
rect 17410 17380 17414 17436
rect 17350 17376 17414 17380
rect 17430 17436 17494 17440
rect 17430 17380 17434 17436
rect 17434 17380 17490 17436
rect 17490 17380 17494 17436
rect 17430 17376 17494 17380
rect 23906 17436 23970 17440
rect 23906 17380 23910 17436
rect 23910 17380 23966 17436
rect 23966 17380 23970 17436
rect 23906 17376 23970 17380
rect 23986 17436 24050 17440
rect 23986 17380 23990 17436
rect 23990 17380 24046 17436
rect 24046 17380 24050 17436
rect 23986 17376 24050 17380
rect 24066 17436 24130 17440
rect 24066 17380 24070 17436
rect 24070 17380 24126 17436
rect 24126 17380 24130 17436
rect 24066 17376 24130 17380
rect 24146 17436 24210 17440
rect 24146 17380 24150 17436
rect 24150 17380 24206 17436
rect 24206 17380 24210 17436
rect 24146 17376 24210 17380
rect 7116 16892 7180 16896
rect 7116 16836 7120 16892
rect 7120 16836 7176 16892
rect 7176 16836 7180 16892
rect 7116 16832 7180 16836
rect 7196 16892 7260 16896
rect 7196 16836 7200 16892
rect 7200 16836 7256 16892
rect 7256 16836 7260 16892
rect 7196 16832 7260 16836
rect 7276 16892 7340 16896
rect 7276 16836 7280 16892
rect 7280 16836 7336 16892
rect 7336 16836 7340 16892
rect 7276 16832 7340 16836
rect 7356 16892 7420 16896
rect 7356 16836 7360 16892
rect 7360 16836 7416 16892
rect 7416 16836 7420 16892
rect 7356 16832 7420 16836
rect 13832 16892 13896 16896
rect 13832 16836 13836 16892
rect 13836 16836 13892 16892
rect 13892 16836 13896 16892
rect 13832 16832 13896 16836
rect 13912 16892 13976 16896
rect 13912 16836 13916 16892
rect 13916 16836 13972 16892
rect 13972 16836 13976 16892
rect 13912 16832 13976 16836
rect 13992 16892 14056 16896
rect 13992 16836 13996 16892
rect 13996 16836 14052 16892
rect 14052 16836 14056 16892
rect 13992 16832 14056 16836
rect 14072 16892 14136 16896
rect 14072 16836 14076 16892
rect 14076 16836 14132 16892
rect 14132 16836 14136 16892
rect 14072 16832 14136 16836
rect 20548 16892 20612 16896
rect 20548 16836 20552 16892
rect 20552 16836 20608 16892
rect 20608 16836 20612 16892
rect 20548 16832 20612 16836
rect 20628 16892 20692 16896
rect 20628 16836 20632 16892
rect 20632 16836 20688 16892
rect 20688 16836 20692 16892
rect 20628 16832 20692 16836
rect 20708 16892 20772 16896
rect 20708 16836 20712 16892
rect 20712 16836 20768 16892
rect 20768 16836 20772 16892
rect 20708 16832 20772 16836
rect 20788 16892 20852 16896
rect 20788 16836 20792 16892
rect 20792 16836 20848 16892
rect 20848 16836 20852 16892
rect 20788 16832 20852 16836
rect 27264 16892 27328 16896
rect 27264 16836 27268 16892
rect 27268 16836 27324 16892
rect 27324 16836 27328 16892
rect 27264 16832 27328 16836
rect 27344 16892 27408 16896
rect 27344 16836 27348 16892
rect 27348 16836 27404 16892
rect 27404 16836 27408 16892
rect 27344 16832 27408 16836
rect 27424 16892 27488 16896
rect 27424 16836 27428 16892
rect 27428 16836 27484 16892
rect 27484 16836 27488 16892
rect 27424 16832 27488 16836
rect 27504 16892 27568 16896
rect 27504 16836 27508 16892
rect 27508 16836 27564 16892
rect 27564 16836 27568 16892
rect 27504 16832 27568 16836
rect 12572 16628 12636 16692
rect 16068 16628 16132 16692
rect 3758 16348 3822 16352
rect 3758 16292 3762 16348
rect 3762 16292 3818 16348
rect 3818 16292 3822 16348
rect 3758 16288 3822 16292
rect 3838 16348 3902 16352
rect 3838 16292 3842 16348
rect 3842 16292 3898 16348
rect 3898 16292 3902 16348
rect 3838 16288 3902 16292
rect 3918 16348 3982 16352
rect 3918 16292 3922 16348
rect 3922 16292 3978 16348
rect 3978 16292 3982 16348
rect 3918 16288 3982 16292
rect 3998 16348 4062 16352
rect 3998 16292 4002 16348
rect 4002 16292 4058 16348
rect 4058 16292 4062 16348
rect 3998 16288 4062 16292
rect 10474 16348 10538 16352
rect 10474 16292 10478 16348
rect 10478 16292 10534 16348
rect 10534 16292 10538 16348
rect 10474 16288 10538 16292
rect 10554 16348 10618 16352
rect 10554 16292 10558 16348
rect 10558 16292 10614 16348
rect 10614 16292 10618 16348
rect 10554 16288 10618 16292
rect 10634 16348 10698 16352
rect 10634 16292 10638 16348
rect 10638 16292 10694 16348
rect 10694 16292 10698 16348
rect 10634 16288 10698 16292
rect 10714 16348 10778 16352
rect 10714 16292 10718 16348
rect 10718 16292 10774 16348
rect 10774 16292 10778 16348
rect 10714 16288 10778 16292
rect 17190 16348 17254 16352
rect 17190 16292 17194 16348
rect 17194 16292 17250 16348
rect 17250 16292 17254 16348
rect 17190 16288 17254 16292
rect 17270 16348 17334 16352
rect 17270 16292 17274 16348
rect 17274 16292 17330 16348
rect 17330 16292 17334 16348
rect 17270 16288 17334 16292
rect 17350 16348 17414 16352
rect 17350 16292 17354 16348
rect 17354 16292 17410 16348
rect 17410 16292 17414 16348
rect 17350 16288 17414 16292
rect 17430 16348 17494 16352
rect 17430 16292 17434 16348
rect 17434 16292 17490 16348
rect 17490 16292 17494 16348
rect 17430 16288 17494 16292
rect 23906 16348 23970 16352
rect 23906 16292 23910 16348
rect 23910 16292 23966 16348
rect 23966 16292 23970 16348
rect 23906 16288 23970 16292
rect 23986 16348 24050 16352
rect 23986 16292 23990 16348
rect 23990 16292 24046 16348
rect 24046 16292 24050 16348
rect 23986 16288 24050 16292
rect 24066 16348 24130 16352
rect 24066 16292 24070 16348
rect 24070 16292 24126 16348
rect 24126 16292 24130 16348
rect 24066 16288 24130 16292
rect 24146 16348 24210 16352
rect 24146 16292 24150 16348
rect 24150 16292 24206 16348
rect 24206 16292 24210 16348
rect 24146 16288 24210 16292
rect 7116 15804 7180 15808
rect 7116 15748 7120 15804
rect 7120 15748 7176 15804
rect 7176 15748 7180 15804
rect 7116 15744 7180 15748
rect 7196 15804 7260 15808
rect 7196 15748 7200 15804
rect 7200 15748 7256 15804
rect 7256 15748 7260 15804
rect 7196 15744 7260 15748
rect 7276 15804 7340 15808
rect 7276 15748 7280 15804
rect 7280 15748 7336 15804
rect 7336 15748 7340 15804
rect 7276 15744 7340 15748
rect 7356 15804 7420 15808
rect 7356 15748 7360 15804
rect 7360 15748 7416 15804
rect 7416 15748 7420 15804
rect 7356 15744 7420 15748
rect 13832 15804 13896 15808
rect 13832 15748 13836 15804
rect 13836 15748 13892 15804
rect 13892 15748 13896 15804
rect 13832 15744 13896 15748
rect 13912 15804 13976 15808
rect 13912 15748 13916 15804
rect 13916 15748 13972 15804
rect 13972 15748 13976 15804
rect 13912 15744 13976 15748
rect 13992 15804 14056 15808
rect 13992 15748 13996 15804
rect 13996 15748 14052 15804
rect 14052 15748 14056 15804
rect 13992 15744 14056 15748
rect 14072 15804 14136 15808
rect 14072 15748 14076 15804
rect 14076 15748 14132 15804
rect 14132 15748 14136 15804
rect 14072 15744 14136 15748
rect 20548 15804 20612 15808
rect 20548 15748 20552 15804
rect 20552 15748 20608 15804
rect 20608 15748 20612 15804
rect 20548 15744 20612 15748
rect 20628 15804 20692 15808
rect 20628 15748 20632 15804
rect 20632 15748 20688 15804
rect 20688 15748 20692 15804
rect 20628 15744 20692 15748
rect 20708 15804 20772 15808
rect 20708 15748 20712 15804
rect 20712 15748 20768 15804
rect 20768 15748 20772 15804
rect 20708 15744 20772 15748
rect 20788 15804 20852 15808
rect 20788 15748 20792 15804
rect 20792 15748 20848 15804
rect 20848 15748 20852 15804
rect 20788 15744 20852 15748
rect 27264 15804 27328 15808
rect 27264 15748 27268 15804
rect 27268 15748 27324 15804
rect 27324 15748 27328 15804
rect 27264 15744 27328 15748
rect 27344 15804 27408 15808
rect 27344 15748 27348 15804
rect 27348 15748 27404 15804
rect 27404 15748 27408 15804
rect 27344 15744 27408 15748
rect 27424 15804 27488 15808
rect 27424 15748 27428 15804
rect 27428 15748 27484 15804
rect 27484 15748 27488 15804
rect 27424 15744 27488 15748
rect 27504 15804 27568 15808
rect 27504 15748 27508 15804
rect 27508 15748 27564 15804
rect 27564 15748 27568 15804
rect 27504 15744 27568 15748
rect 5212 15540 5276 15604
rect 3758 15260 3822 15264
rect 3758 15204 3762 15260
rect 3762 15204 3818 15260
rect 3818 15204 3822 15260
rect 3758 15200 3822 15204
rect 3838 15260 3902 15264
rect 3838 15204 3842 15260
rect 3842 15204 3898 15260
rect 3898 15204 3902 15260
rect 3838 15200 3902 15204
rect 3918 15260 3982 15264
rect 3918 15204 3922 15260
rect 3922 15204 3978 15260
rect 3978 15204 3982 15260
rect 3918 15200 3982 15204
rect 3998 15260 4062 15264
rect 3998 15204 4002 15260
rect 4002 15204 4058 15260
rect 4058 15204 4062 15260
rect 3998 15200 4062 15204
rect 10474 15260 10538 15264
rect 10474 15204 10478 15260
rect 10478 15204 10534 15260
rect 10534 15204 10538 15260
rect 10474 15200 10538 15204
rect 10554 15260 10618 15264
rect 10554 15204 10558 15260
rect 10558 15204 10614 15260
rect 10614 15204 10618 15260
rect 10554 15200 10618 15204
rect 10634 15260 10698 15264
rect 10634 15204 10638 15260
rect 10638 15204 10694 15260
rect 10694 15204 10698 15260
rect 10634 15200 10698 15204
rect 10714 15260 10778 15264
rect 10714 15204 10718 15260
rect 10718 15204 10774 15260
rect 10774 15204 10778 15260
rect 10714 15200 10778 15204
rect 17190 15260 17254 15264
rect 17190 15204 17194 15260
rect 17194 15204 17250 15260
rect 17250 15204 17254 15260
rect 17190 15200 17254 15204
rect 17270 15260 17334 15264
rect 17270 15204 17274 15260
rect 17274 15204 17330 15260
rect 17330 15204 17334 15260
rect 17270 15200 17334 15204
rect 17350 15260 17414 15264
rect 17350 15204 17354 15260
rect 17354 15204 17410 15260
rect 17410 15204 17414 15260
rect 17350 15200 17414 15204
rect 17430 15260 17494 15264
rect 17430 15204 17434 15260
rect 17434 15204 17490 15260
rect 17490 15204 17494 15260
rect 17430 15200 17494 15204
rect 23906 15260 23970 15264
rect 23906 15204 23910 15260
rect 23910 15204 23966 15260
rect 23966 15204 23970 15260
rect 23906 15200 23970 15204
rect 23986 15260 24050 15264
rect 23986 15204 23990 15260
rect 23990 15204 24046 15260
rect 24046 15204 24050 15260
rect 23986 15200 24050 15204
rect 24066 15260 24130 15264
rect 24066 15204 24070 15260
rect 24070 15204 24126 15260
rect 24126 15204 24130 15260
rect 24066 15200 24130 15204
rect 24146 15260 24210 15264
rect 24146 15204 24150 15260
rect 24150 15204 24206 15260
rect 24206 15204 24210 15260
rect 24146 15200 24210 15204
rect 11284 15192 11348 15196
rect 11284 15136 11298 15192
rect 11298 15136 11348 15192
rect 11284 15132 11348 15136
rect 7116 14716 7180 14720
rect 7116 14660 7120 14716
rect 7120 14660 7176 14716
rect 7176 14660 7180 14716
rect 7116 14656 7180 14660
rect 7196 14716 7260 14720
rect 7196 14660 7200 14716
rect 7200 14660 7256 14716
rect 7256 14660 7260 14716
rect 7196 14656 7260 14660
rect 7276 14716 7340 14720
rect 7276 14660 7280 14716
rect 7280 14660 7336 14716
rect 7336 14660 7340 14716
rect 7276 14656 7340 14660
rect 7356 14716 7420 14720
rect 7356 14660 7360 14716
rect 7360 14660 7416 14716
rect 7416 14660 7420 14716
rect 7356 14656 7420 14660
rect 13832 14716 13896 14720
rect 13832 14660 13836 14716
rect 13836 14660 13892 14716
rect 13892 14660 13896 14716
rect 13832 14656 13896 14660
rect 13912 14716 13976 14720
rect 13912 14660 13916 14716
rect 13916 14660 13972 14716
rect 13972 14660 13976 14716
rect 13912 14656 13976 14660
rect 13992 14716 14056 14720
rect 13992 14660 13996 14716
rect 13996 14660 14052 14716
rect 14052 14660 14056 14716
rect 13992 14656 14056 14660
rect 14072 14716 14136 14720
rect 14072 14660 14076 14716
rect 14076 14660 14132 14716
rect 14132 14660 14136 14716
rect 14072 14656 14136 14660
rect 20548 14716 20612 14720
rect 20548 14660 20552 14716
rect 20552 14660 20608 14716
rect 20608 14660 20612 14716
rect 20548 14656 20612 14660
rect 20628 14716 20692 14720
rect 20628 14660 20632 14716
rect 20632 14660 20688 14716
rect 20688 14660 20692 14716
rect 20628 14656 20692 14660
rect 20708 14716 20772 14720
rect 20708 14660 20712 14716
rect 20712 14660 20768 14716
rect 20768 14660 20772 14716
rect 20708 14656 20772 14660
rect 20788 14716 20852 14720
rect 20788 14660 20792 14716
rect 20792 14660 20848 14716
rect 20848 14660 20852 14716
rect 20788 14656 20852 14660
rect 27264 14716 27328 14720
rect 27264 14660 27268 14716
rect 27268 14660 27324 14716
rect 27324 14660 27328 14716
rect 27264 14656 27328 14660
rect 27344 14716 27408 14720
rect 27344 14660 27348 14716
rect 27348 14660 27404 14716
rect 27404 14660 27408 14716
rect 27344 14656 27408 14660
rect 27424 14716 27488 14720
rect 27424 14660 27428 14716
rect 27428 14660 27484 14716
rect 27484 14660 27488 14716
rect 27424 14656 27488 14660
rect 27504 14716 27568 14720
rect 27504 14660 27508 14716
rect 27508 14660 27564 14716
rect 27564 14660 27568 14716
rect 27504 14656 27568 14660
rect 3758 14172 3822 14176
rect 3758 14116 3762 14172
rect 3762 14116 3818 14172
rect 3818 14116 3822 14172
rect 3758 14112 3822 14116
rect 3838 14172 3902 14176
rect 3838 14116 3842 14172
rect 3842 14116 3898 14172
rect 3898 14116 3902 14172
rect 3838 14112 3902 14116
rect 3918 14172 3982 14176
rect 3918 14116 3922 14172
rect 3922 14116 3978 14172
rect 3978 14116 3982 14172
rect 3918 14112 3982 14116
rect 3998 14172 4062 14176
rect 3998 14116 4002 14172
rect 4002 14116 4058 14172
rect 4058 14116 4062 14172
rect 3998 14112 4062 14116
rect 10474 14172 10538 14176
rect 10474 14116 10478 14172
rect 10478 14116 10534 14172
rect 10534 14116 10538 14172
rect 10474 14112 10538 14116
rect 10554 14172 10618 14176
rect 10554 14116 10558 14172
rect 10558 14116 10614 14172
rect 10614 14116 10618 14172
rect 10554 14112 10618 14116
rect 10634 14172 10698 14176
rect 10634 14116 10638 14172
rect 10638 14116 10694 14172
rect 10694 14116 10698 14172
rect 10634 14112 10698 14116
rect 10714 14172 10778 14176
rect 10714 14116 10718 14172
rect 10718 14116 10774 14172
rect 10774 14116 10778 14172
rect 10714 14112 10778 14116
rect 17190 14172 17254 14176
rect 17190 14116 17194 14172
rect 17194 14116 17250 14172
rect 17250 14116 17254 14172
rect 17190 14112 17254 14116
rect 17270 14172 17334 14176
rect 17270 14116 17274 14172
rect 17274 14116 17330 14172
rect 17330 14116 17334 14172
rect 17270 14112 17334 14116
rect 17350 14172 17414 14176
rect 17350 14116 17354 14172
rect 17354 14116 17410 14172
rect 17410 14116 17414 14172
rect 17350 14112 17414 14116
rect 17430 14172 17494 14176
rect 17430 14116 17434 14172
rect 17434 14116 17490 14172
rect 17490 14116 17494 14172
rect 17430 14112 17494 14116
rect 23906 14172 23970 14176
rect 23906 14116 23910 14172
rect 23910 14116 23966 14172
rect 23966 14116 23970 14172
rect 23906 14112 23970 14116
rect 23986 14172 24050 14176
rect 23986 14116 23990 14172
rect 23990 14116 24046 14172
rect 24046 14116 24050 14172
rect 23986 14112 24050 14116
rect 24066 14172 24130 14176
rect 24066 14116 24070 14172
rect 24070 14116 24126 14172
rect 24126 14116 24130 14172
rect 24066 14112 24130 14116
rect 24146 14172 24210 14176
rect 24146 14116 24150 14172
rect 24150 14116 24206 14172
rect 24206 14116 24210 14172
rect 24146 14112 24210 14116
rect 12572 13908 12636 13972
rect 7116 13628 7180 13632
rect 7116 13572 7120 13628
rect 7120 13572 7176 13628
rect 7176 13572 7180 13628
rect 7116 13568 7180 13572
rect 7196 13628 7260 13632
rect 7196 13572 7200 13628
rect 7200 13572 7256 13628
rect 7256 13572 7260 13628
rect 7196 13568 7260 13572
rect 7276 13628 7340 13632
rect 7276 13572 7280 13628
rect 7280 13572 7336 13628
rect 7336 13572 7340 13628
rect 7276 13568 7340 13572
rect 7356 13628 7420 13632
rect 7356 13572 7360 13628
rect 7360 13572 7416 13628
rect 7416 13572 7420 13628
rect 7356 13568 7420 13572
rect 13832 13628 13896 13632
rect 13832 13572 13836 13628
rect 13836 13572 13892 13628
rect 13892 13572 13896 13628
rect 13832 13568 13896 13572
rect 13912 13628 13976 13632
rect 13912 13572 13916 13628
rect 13916 13572 13972 13628
rect 13972 13572 13976 13628
rect 13912 13568 13976 13572
rect 13992 13628 14056 13632
rect 13992 13572 13996 13628
rect 13996 13572 14052 13628
rect 14052 13572 14056 13628
rect 13992 13568 14056 13572
rect 14072 13628 14136 13632
rect 14072 13572 14076 13628
rect 14076 13572 14132 13628
rect 14132 13572 14136 13628
rect 14072 13568 14136 13572
rect 20548 13628 20612 13632
rect 20548 13572 20552 13628
rect 20552 13572 20608 13628
rect 20608 13572 20612 13628
rect 20548 13568 20612 13572
rect 20628 13628 20692 13632
rect 20628 13572 20632 13628
rect 20632 13572 20688 13628
rect 20688 13572 20692 13628
rect 20628 13568 20692 13572
rect 20708 13628 20772 13632
rect 20708 13572 20712 13628
rect 20712 13572 20768 13628
rect 20768 13572 20772 13628
rect 20708 13568 20772 13572
rect 20788 13628 20852 13632
rect 20788 13572 20792 13628
rect 20792 13572 20848 13628
rect 20848 13572 20852 13628
rect 20788 13568 20852 13572
rect 27264 13628 27328 13632
rect 27264 13572 27268 13628
rect 27268 13572 27324 13628
rect 27324 13572 27328 13628
rect 27264 13568 27328 13572
rect 27344 13628 27408 13632
rect 27344 13572 27348 13628
rect 27348 13572 27404 13628
rect 27404 13572 27408 13628
rect 27344 13568 27408 13572
rect 27424 13628 27488 13632
rect 27424 13572 27428 13628
rect 27428 13572 27484 13628
rect 27484 13572 27488 13628
rect 27424 13568 27488 13572
rect 27504 13628 27568 13632
rect 27504 13572 27508 13628
rect 27508 13572 27564 13628
rect 27564 13572 27568 13628
rect 27504 13568 27568 13572
rect 3758 13084 3822 13088
rect 3758 13028 3762 13084
rect 3762 13028 3818 13084
rect 3818 13028 3822 13084
rect 3758 13024 3822 13028
rect 3838 13084 3902 13088
rect 3838 13028 3842 13084
rect 3842 13028 3898 13084
rect 3898 13028 3902 13084
rect 3838 13024 3902 13028
rect 3918 13084 3982 13088
rect 3918 13028 3922 13084
rect 3922 13028 3978 13084
rect 3978 13028 3982 13084
rect 3918 13024 3982 13028
rect 3998 13084 4062 13088
rect 3998 13028 4002 13084
rect 4002 13028 4058 13084
rect 4058 13028 4062 13084
rect 3998 13024 4062 13028
rect 10474 13084 10538 13088
rect 10474 13028 10478 13084
rect 10478 13028 10534 13084
rect 10534 13028 10538 13084
rect 10474 13024 10538 13028
rect 10554 13084 10618 13088
rect 10554 13028 10558 13084
rect 10558 13028 10614 13084
rect 10614 13028 10618 13084
rect 10554 13024 10618 13028
rect 10634 13084 10698 13088
rect 10634 13028 10638 13084
rect 10638 13028 10694 13084
rect 10694 13028 10698 13084
rect 10634 13024 10698 13028
rect 10714 13084 10778 13088
rect 10714 13028 10718 13084
rect 10718 13028 10774 13084
rect 10774 13028 10778 13084
rect 10714 13024 10778 13028
rect 17190 13084 17254 13088
rect 17190 13028 17194 13084
rect 17194 13028 17250 13084
rect 17250 13028 17254 13084
rect 17190 13024 17254 13028
rect 17270 13084 17334 13088
rect 17270 13028 17274 13084
rect 17274 13028 17330 13084
rect 17330 13028 17334 13084
rect 17270 13024 17334 13028
rect 17350 13084 17414 13088
rect 17350 13028 17354 13084
rect 17354 13028 17410 13084
rect 17410 13028 17414 13084
rect 17350 13024 17414 13028
rect 17430 13084 17494 13088
rect 17430 13028 17434 13084
rect 17434 13028 17490 13084
rect 17490 13028 17494 13084
rect 17430 13024 17494 13028
rect 23906 13084 23970 13088
rect 23906 13028 23910 13084
rect 23910 13028 23966 13084
rect 23966 13028 23970 13084
rect 23906 13024 23970 13028
rect 23986 13084 24050 13088
rect 23986 13028 23990 13084
rect 23990 13028 24046 13084
rect 24046 13028 24050 13084
rect 23986 13024 24050 13028
rect 24066 13084 24130 13088
rect 24066 13028 24070 13084
rect 24070 13028 24126 13084
rect 24126 13028 24130 13084
rect 24066 13024 24130 13028
rect 24146 13084 24210 13088
rect 24146 13028 24150 13084
rect 24150 13028 24206 13084
rect 24206 13028 24210 13084
rect 24146 13024 24210 13028
rect 7116 12540 7180 12544
rect 7116 12484 7120 12540
rect 7120 12484 7176 12540
rect 7176 12484 7180 12540
rect 7116 12480 7180 12484
rect 7196 12540 7260 12544
rect 7196 12484 7200 12540
rect 7200 12484 7256 12540
rect 7256 12484 7260 12540
rect 7196 12480 7260 12484
rect 7276 12540 7340 12544
rect 7276 12484 7280 12540
rect 7280 12484 7336 12540
rect 7336 12484 7340 12540
rect 7276 12480 7340 12484
rect 7356 12540 7420 12544
rect 7356 12484 7360 12540
rect 7360 12484 7416 12540
rect 7416 12484 7420 12540
rect 7356 12480 7420 12484
rect 13832 12540 13896 12544
rect 13832 12484 13836 12540
rect 13836 12484 13892 12540
rect 13892 12484 13896 12540
rect 13832 12480 13896 12484
rect 13912 12540 13976 12544
rect 13912 12484 13916 12540
rect 13916 12484 13972 12540
rect 13972 12484 13976 12540
rect 13912 12480 13976 12484
rect 13992 12540 14056 12544
rect 13992 12484 13996 12540
rect 13996 12484 14052 12540
rect 14052 12484 14056 12540
rect 13992 12480 14056 12484
rect 14072 12540 14136 12544
rect 14072 12484 14076 12540
rect 14076 12484 14132 12540
rect 14132 12484 14136 12540
rect 14072 12480 14136 12484
rect 20548 12540 20612 12544
rect 20548 12484 20552 12540
rect 20552 12484 20608 12540
rect 20608 12484 20612 12540
rect 20548 12480 20612 12484
rect 20628 12540 20692 12544
rect 20628 12484 20632 12540
rect 20632 12484 20688 12540
rect 20688 12484 20692 12540
rect 20628 12480 20692 12484
rect 20708 12540 20772 12544
rect 20708 12484 20712 12540
rect 20712 12484 20768 12540
rect 20768 12484 20772 12540
rect 20708 12480 20772 12484
rect 20788 12540 20852 12544
rect 20788 12484 20792 12540
rect 20792 12484 20848 12540
rect 20848 12484 20852 12540
rect 20788 12480 20852 12484
rect 27264 12540 27328 12544
rect 27264 12484 27268 12540
rect 27268 12484 27324 12540
rect 27324 12484 27328 12540
rect 27264 12480 27328 12484
rect 27344 12540 27408 12544
rect 27344 12484 27348 12540
rect 27348 12484 27404 12540
rect 27404 12484 27408 12540
rect 27344 12480 27408 12484
rect 27424 12540 27488 12544
rect 27424 12484 27428 12540
rect 27428 12484 27484 12540
rect 27484 12484 27488 12540
rect 27424 12480 27488 12484
rect 27504 12540 27568 12544
rect 27504 12484 27508 12540
rect 27508 12484 27564 12540
rect 27564 12484 27568 12540
rect 27504 12480 27568 12484
rect 3758 11996 3822 12000
rect 3758 11940 3762 11996
rect 3762 11940 3818 11996
rect 3818 11940 3822 11996
rect 3758 11936 3822 11940
rect 3838 11996 3902 12000
rect 3838 11940 3842 11996
rect 3842 11940 3898 11996
rect 3898 11940 3902 11996
rect 3838 11936 3902 11940
rect 3918 11996 3982 12000
rect 3918 11940 3922 11996
rect 3922 11940 3978 11996
rect 3978 11940 3982 11996
rect 3918 11936 3982 11940
rect 3998 11996 4062 12000
rect 3998 11940 4002 11996
rect 4002 11940 4058 11996
rect 4058 11940 4062 11996
rect 3998 11936 4062 11940
rect 10474 11996 10538 12000
rect 10474 11940 10478 11996
rect 10478 11940 10534 11996
rect 10534 11940 10538 11996
rect 10474 11936 10538 11940
rect 10554 11996 10618 12000
rect 10554 11940 10558 11996
rect 10558 11940 10614 11996
rect 10614 11940 10618 11996
rect 10554 11936 10618 11940
rect 10634 11996 10698 12000
rect 10634 11940 10638 11996
rect 10638 11940 10694 11996
rect 10694 11940 10698 11996
rect 10634 11936 10698 11940
rect 10714 11996 10778 12000
rect 10714 11940 10718 11996
rect 10718 11940 10774 11996
rect 10774 11940 10778 11996
rect 10714 11936 10778 11940
rect 17190 11996 17254 12000
rect 17190 11940 17194 11996
rect 17194 11940 17250 11996
rect 17250 11940 17254 11996
rect 17190 11936 17254 11940
rect 17270 11996 17334 12000
rect 17270 11940 17274 11996
rect 17274 11940 17330 11996
rect 17330 11940 17334 11996
rect 17270 11936 17334 11940
rect 17350 11996 17414 12000
rect 17350 11940 17354 11996
rect 17354 11940 17410 11996
rect 17410 11940 17414 11996
rect 17350 11936 17414 11940
rect 17430 11996 17494 12000
rect 17430 11940 17434 11996
rect 17434 11940 17490 11996
rect 17490 11940 17494 11996
rect 17430 11936 17494 11940
rect 23906 11996 23970 12000
rect 23906 11940 23910 11996
rect 23910 11940 23966 11996
rect 23966 11940 23970 11996
rect 23906 11936 23970 11940
rect 23986 11996 24050 12000
rect 23986 11940 23990 11996
rect 23990 11940 24046 11996
rect 24046 11940 24050 11996
rect 23986 11936 24050 11940
rect 24066 11996 24130 12000
rect 24066 11940 24070 11996
rect 24070 11940 24126 11996
rect 24126 11940 24130 11996
rect 24066 11936 24130 11940
rect 24146 11996 24210 12000
rect 24146 11940 24150 11996
rect 24150 11940 24206 11996
rect 24206 11940 24210 11996
rect 24146 11936 24210 11940
rect 7116 11452 7180 11456
rect 7116 11396 7120 11452
rect 7120 11396 7176 11452
rect 7176 11396 7180 11452
rect 7116 11392 7180 11396
rect 7196 11452 7260 11456
rect 7196 11396 7200 11452
rect 7200 11396 7256 11452
rect 7256 11396 7260 11452
rect 7196 11392 7260 11396
rect 7276 11452 7340 11456
rect 7276 11396 7280 11452
rect 7280 11396 7336 11452
rect 7336 11396 7340 11452
rect 7276 11392 7340 11396
rect 7356 11452 7420 11456
rect 7356 11396 7360 11452
rect 7360 11396 7416 11452
rect 7416 11396 7420 11452
rect 7356 11392 7420 11396
rect 13832 11452 13896 11456
rect 13832 11396 13836 11452
rect 13836 11396 13892 11452
rect 13892 11396 13896 11452
rect 13832 11392 13896 11396
rect 13912 11452 13976 11456
rect 13912 11396 13916 11452
rect 13916 11396 13972 11452
rect 13972 11396 13976 11452
rect 13912 11392 13976 11396
rect 13992 11452 14056 11456
rect 13992 11396 13996 11452
rect 13996 11396 14052 11452
rect 14052 11396 14056 11452
rect 13992 11392 14056 11396
rect 14072 11452 14136 11456
rect 14072 11396 14076 11452
rect 14076 11396 14132 11452
rect 14132 11396 14136 11452
rect 14072 11392 14136 11396
rect 20548 11452 20612 11456
rect 20548 11396 20552 11452
rect 20552 11396 20608 11452
rect 20608 11396 20612 11452
rect 20548 11392 20612 11396
rect 20628 11452 20692 11456
rect 20628 11396 20632 11452
rect 20632 11396 20688 11452
rect 20688 11396 20692 11452
rect 20628 11392 20692 11396
rect 20708 11452 20772 11456
rect 20708 11396 20712 11452
rect 20712 11396 20768 11452
rect 20768 11396 20772 11452
rect 20708 11392 20772 11396
rect 20788 11452 20852 11456
rect 20788 11396 20792 11452
rect 20792 11396 20848 11452
rect 20848 11396 20852 11452
rect 20788 11392 20852 11396
rect 27264 11452 27328 11456
rect 27264 11396 27268 11452
rect 27268 11396 27324 11452
rect 27324 11396 27328 11452
rect 27264 11392 27328 11396
rect 27344 11452 27408 11456
rect 27344 11396 27348 11452
rect 27348 11396 27404 11452
rect 27404 11396 27408 11452
rect 27344 11392 27408 11396
rect 27424 11452 27488 11456
rect 27424 11396 27428 11452
rect 27428 11396 27484 11452
rect 27484 11396 27488 11452
rect 27424 11392 27488 11396
rect 27504 11452 27568 11456
rect 27504 11396 27508 11452
rect 27508 11396 27564 11452
rect 27564 11396 27568 11452
rect 27504 11392 27568 11396
rect 3758 10908 3822 10912
rect 3758 10852 3762 10908
rect 3762 10852 3818 10908
rect 3818 10852 3822 10908
rect 3758 10848 3822 10852
rect 3838 10908 3902 10912
rect 3838 10852 3842 10908
rect 3842 10852 3898 10908
rect 3898 10852 3902 10908
rect 3838 10848 3902 10852
rect 3918 10908 3982 10912
rect 3918 10852 3922 10908
rect 3922 10852 3978 10908
rect 3978 10852 3982 10908
rect 3918 10848 3982 10852
rect 3998 10908 4062 10912
rect 3998 10852 4002 10908
rect 4002 10852 4058 10908
rect 4058 10852 4062 10908
rect 3998 10848 4062 10852
rect 10474 10908 10538 10912
rect 10474 10852 10478 10908
rect 10478 10852 10534 10908
rect 10534 10852 10538 10908
rect 10474 10848 10538 10852
rect 10554 10908 10618 10912
rect 10554 10852 10558 10908
rect 10558 10852 10614 10908
rect 10614 10852 10618 10908
rect 10554 10848 10618 10852
rect 10634 10908 10698 10912
rect 10634 10852 10638 10908
rect 10638 10852 10694 10908
rect 10694 10852 10698 10908
rect 10634 10848 10698 10852
rect 10714 10908 10778 10912
rect 10714 10852 10718 10908
rect 10718 10852 10774 10908
rect 10774 10852 10778 10908
rect 10714 10848 10778 10852
rect 17190 10908 17254 10912
rect 17190 10852 17194 10908
rect 17194 10852 17250 10908
rect 17250 10852 17254 10908
rect 17190 10848 17254 10852
rect 17270 10908 17334 10912
rect 17270 10852 17274 10908
rect 17274 10852 17330 10908
rect 17330 10852 17334 10908
rect 17270 10848 17334 10852
rect 17350 10908 17414 10912
rect 17350 10852 17354 10908
rect 17354 10852 17410 10908
rect 17410 10852 17414 10908
rect 17350 10848 17414 10852
rect 17430 10908 17494 10912
rect 17430 10852 17434 10908
rect 17434 10852 17490 10908
rect 17490 10852 17494 10908
rect 17430 10848 17494 10852
rect 23906 10908 23970 10912
rect 23906 10852 23910 10908
rect 23910 10852 23966 10908
rect 23966 10852 23970 10908
rect 23906 10848 23970 10852
rect 23986 10908 24050 10912
rect 23986 10852 23990 10908
rect 23990 10852 24046 10908
rect 24046 10852 24050 10908
rect 23986 10848 24050 10852
rect 24066 10908 24130 10912
rect 24066 10852 24070 10908
rect 24070 10852 24126 10908
rect 24126 10852 24130 10908
rect 24066 10848 24130 10852
rect 24146 10908 24210 10912
rect 24146 10852 24150 10908
rect 24150 10852 24206 10908
rect 24206 10852 24210 10908
rect 24146 10848 24210 10852
rect 7116 10364 7180 10368
rect 7116 10308 7120 10364
rect 7120 10308 7176 10364
rect 7176 10308 7180 10364
rect 7116 10304 7180 10308
rect 7196 10364 7260 10368
rect 7196 10308 7200 10364
rect 7200 10308 7256 10364
rect 7256 10308 7260 10364
rect 7196 10304 7260 10308
rect 7276 10364 7340 10368
rect 7276 10308 7280 10364
rect 7280 10308 7336 10364
rect 7336 10308 7340 10364
rect 7276 10304 7340 10308
rect 7356 10364 7420 10368
rect 7356 10308 7360 10364
rect 7360 10308 7416 10364
rect 7416 10308 7420 10364
rect 7356 10304 7420 10308
rect 13832 10364 13896 10368
rect 13832 10308 13836 10364
rect 13836 10308 13892 10364
rect 13892 10308 13896 10364
rect 13832 10304 13896 10308
rect 13912 10364 13976 10368
rect 13912 10308 13916 10364
rect 13916 10308 13972 10364
rect 13972 10308 13976 10364
rect 13912 10304 13976 10308
rect 13992 10364 14056 10368
rect 13992 10308 13996 10364
rect 13996 10308 14052 10364
rect 14052 10308 14056 10364
rect 13992 10304 14056 10308
rect 14072 10364 14136 10368
rect 14072 10308 14076 10364
rect 14076 10308 14132 10364
rect 14132 10308 14136 10364
rect 14072 10304 14136 10308
rect 20548 10364 20612 10368
rect 20548 10308 20552 10364
rect 20552 10308 20608 10364
rect 20608 10308 20612 10364
rect 20548 10304 20612 10308
rect 20628 10364 20692 10368
rect 20628 10308 20632 10364
rect 20632 10308 20688 10364
rect 20688 10308 20692 10364
rect 20628 10304 20692 10308
rect 20708 10364 20772 10368
rect 20708 10308 20712 10364
rect 20712 10308 20768 10364
rect 20768 10308 20772 10364
rect 20708 10304 20772 10308
rect 20788 10364 20852 10368
rect 20788 10308 20792 10364
rect 20792 10308 20848 10364
rect 20848 10308 20852 10364
rect 20788 10304 20852 10308
rect 27264 10364 27328 10368
rect 27264 10308 27268 10364
rect 27268 10308 27324 10364
rect 27324 10308 27328 10364
rect 27264 10304 27328 10308
rect 27344 10364 27408 10368
rect 27344 10308 27348 10364
rect 27348 10308 27404 10364
rect 27404 10308 27408 10364
rect 27344 10304 27408 10308
rect 27424 10364 27488 10368
rect 27424 10308 27428 10364
rect 27428 10308 27484 10364
rect 27484 10308 27488 10364
rect 27424 10304 27488 10308
rect 27504 10364 27568 10368
rect 27504 10308 27508 10364
rect 27508 10308 27564 10364
rect 27564 10308 27568 10364
rect 27504 10304 27568 10308
rect 3758 9820 3822 9824
rect 3758 9764 3762 9820
rect 3762 9764 3818 9820
rect 3818 9764 3822 9820
rect 3758 9760 3822 9764
rect 3838 9820 3902 9824
rect 3838 9764 3842 9820
rect 3842 9764 3898 9820
rect 3898 9764 3902 9820
rect 3838 9760 3902 9764
rect 3918 9820 3982 9824
rect 3918 9764 3922 9820
rect 3922 9764 3978 9820
rect 3978 9764 3982 9820
rect 3918 9760 3982 9764
rect 3998 9820 4062 9824
rect 3998 9764 4002 9820
rect 4002 9764 4058 9820
rect 4058 9764 4062 9820
rect 3998 9760 4062 9764
rect 10474 9820 10538 9824
rect 10474 9764 10478 9820
rect 10478 9764 10534 9820
rect 10534 9764 10538 9820
rect 10474 9760 10538 9764
rect 10554 9820 10618 9824
rect 10554 9764 10558 9820
rect 10558 9764 10614 9820
rect 10614 9764 10618 9820
rect 10554 9760 10618 9764
rect 10634 9820 10698 9824
rect 10634 9764 10638 9820
rect 10638 9764 10694 9820
rect 10694 9764 10698 9820
rect 10634 9760 10698 9764
rect 10714 9820 10778 9824
rect 10714 9764 10718 9820
rect 10718 9764 10774 9820
rect 10774 9764 10778 9820
rect 10714 9760 10778 9764
rect 17190 9820 17254 9824
rect 17190 9764 17194 9820
rect 17194 9764 17250 9820
rect 17250 9764 17254 9820
rect 17190 9760 17254 9764
rect 17270 9820 17334 9824
rect 17270 9764 17274 9820
rect 17274 9764 17330 9820
rect 17330 9764 17334 9820
rect 17270 9760 17334 9764
rect 17350 9820 17414 9824
rect 17350 9764 17354 9820
rect 17354 9764 17410 9820
rect 17410 9764 17414 9820
rect 17350 9760 17414 9764
rect 17430 9820 17494 9824
rect 17430 9764 17434 9820
rect 17434 9764 17490 9820
rect 17490 9764 17494 9820
rect 17430 9760 17494 9764
rect 23906 9820 23970 9824
rect 23906 9764 23910 9820
rect 23910 9764 23966 9820
rect 23966 9764 23970 9820
rect 23906 9760 23970 9764
rect 23986 9820 24050 9824
rect 23986 9764 23990 9820
rect 23990 9764 24046 9820
rect 24046 9764 24050 9820
rect 23986 9760 24050 9764
rect 24066 9820 24130 9824
rect 24066 9764 24070 9820
rect 24070 9764 24126 9820
rect 24126 9764 24130 9820
rect 24066 9760 24130 9764
rect 24146 9820 24210 9824
rect 24146 9764 24150 9820
rect 24150 9764 24206 9820
rect 24206 9764 24210 9820
rect 24146 9760 24210 9764
rect 7116 9276 7180 9280
rect 7116 9220 7120 9276
rect 7120 9220 7176 9276
rect 7176 9220 7180 9276
rect 7116 9216 7180 9220
rect 7196 9276 7260 9280
rect 7196 9220 7200 9276
rect 7200 9220 7256 9276
rect 7256 9220 7260 9276
rect 7196 9216 7260 9220
rect 7276 9276 7340 9280
rect 7276 9220 7280 9276
rect 7280 9220 7336 9276
rect 7336 9220 7340 9276
rect 7276 9216 7340 9220
rect 7356 9276 7420 9280
rect 7356 9220 7360 9276
rect 7360 9220 7416 9276
rect 7416 9220 7420 9276
rect 7356 9216 7420 9220
rect 13832 9276 13896 9280
rect 13832 9220 13836 9276
rect 13836 9220 13892 9276
rect 13892 9220 13896 9276
rect 13832 9216 13896 9220
rect 13912 9276 13976 9280
rect 13912 9220 13916 9276
rect 13916 9220 13972 9276
rect 13972 9220 13976 9276
rect 13912 9216 13976 9220
rect 13992 9276 14056 9280
rect 13992 9220 13996 9276
rect 13996 9220 14052 9276
rect 14052 9220 14056 9276
rect 13992 9216 14056 9220
rect 14072 9276 14136 9280
rect 14072 9220 14076 9276
rect 14076 9220 14132 9276
rect 14132 9220 14136 9276
rect 14072 9216 14136 9220
rect 20548 9276 20612 9280
rect 20548 9220 20552 9276
rect 20552 9220 20608 9276
rect 20608 9220 20612 9276
rect 20548 9216 20612 9220
rect 20628 9276 20692 9280
rect 20628 9220 20632 9276
rect 20632 9220 20688 9276
rect 20688 9220 20692 9276
rect 20628 9216 20692 9220
rect 20708 9276 20772 9280
rect 20708 9220 20712 9276
rect 20712 9220 20768 9276
rect 20768 9220 20772 9276
rect 20708 9216 20772 9220
rect 20788 9276 20852 9280
rect 20788 9220 20792 9276
rect 20792 9220 20848 9276
rect 20848 9220 20852 9276
rect 20788 9216 20852 9220
rect 27264 9276 27328 9280
rect 27264 9220 27268 9276
rect 27268 9220 27324 9276
rect 27324 9220 27328 9276
rect 27264 9216 27328 9220
rect 27344 9276 27408 9280
rect 27344 9220 27348 9276
rect 27348 9220 27404 9276
rect 27404 9220 27408 9276
rect 27344 9216 27408 9220
rect 27424 9276 27488 9280
rect 27424 9220 27428 9276
rect 27428 9220 27484 9276
rect 27484 9220 27488 9276
rect 27424 9216 27488 9220
rect 27504 9276 27568 9280
rect 27504 9220 27508 9276
rect 27508 9220 27564 9276
rect 27564 9220 27568 9276
rect 27504 9216 27568 9220
rect 3758 8732 3822 8736
rect 3758 8676 3762 8732
rect 3762 8676 3818 8732
rect 3818 8676 3822 8732
rect 3758 8672 3822 8676
rect 3838 8732 3902 8736
rect 3838 8676 3842 8732
rect 3842 8676 3898 8732
rect 3898 8676 3902 8732
rect 3838 8672 3902 8676
rect 3918 8732 3982 8736
rect 3918 8676 3922 8732
rect 3922 8676 3978 8732
rect 3978 8676 3982 8732
rect 3918 8672 3982 8676
rect 3998 8732 4062 8736
rect 3998 8676 4002 8732
rect 4002 8676 4058 8732
rect 4058 8676 4062 8732
rect 3998 8672 4062 8676
rect 10474 8732 10538 8736
rect 10474 8676 10478 8732
rect 10478 8676 10534 8732
rect 10534 8676 10538 8732
rect 10474 8672 10538 8676
rect 10554 8732 10618 8736
rect 10554 8676 10558 8732
rect 10558 8676 10614 8732
rect 10614 8676 10618 8732
rect 10554 8672 10618 8676
rect 10634 8732 10698 8736
rect 10634 8676 10638 8732
rect 10638 8676 10694 8732
rect 10694 8676 10698 8732
rect 10634 8672 10698 8676
rect 10714 8732 10778 8736
rect 10714 8676 10718 8732
rect 10718 8676 10774 8732
rect 10774 8676 10778 8732
rect 10714 8672 10778 8676
rect 17190 8732 17254 8736
rect 17190 8676 17194 8732
rect 17194 8676 17250 8732
rect 17250 8676 17254 8732
rect 17190 8672 17254 8676
rect 17270 8732 17334 8736
rect 17270 8676 17274 8732
rect 17274 8676 17330 8732
rect 17330 8676 17334 8732
rect 17270 8672 17334 8676
rect 17350 8732 17414 8736
rect 17350 8676 17354 8732
rect 17354 8676 17410 8732
rect 17410 8676 17414 8732
rect 17350 8672 17414 8676
rect 17430 8732 17494 8736
rect 17430 8676 17434 8732
rect 17434 8676 17490 8732
rect 17490 8676 17494 8732
rect 17430 8672 17494 8676
rect 23906 8732 23970 8736
rect 23906 8676 23910 8732
rect 23910 8676 23966 8732
rect 23966 8676 23970 8732
rect 23906 8672 23970 8676
rect 23986 8732 24050 8736
rect 23986 8676 23990 8732
rect 23990 8676 24046 8732
rect 24046 8676 24050 8732
rect 23986 8672 24050 8676
rect 24066 8732 24130 8736
rect 24066 8676 24070 8732
rect 24070 8676 24126 8732
rect 24126 8676 24130 8732
rect 24066 8672 24130 8676
rect 24146 8732 24210 8736
rect 24146 8676 24150 8732
rect 24150 8676 24206 8732
rect 24206 8676 24210 8732
rect 24146 8672 24210 8676
rect 7116 8188 7180 8192
rect 7116 8132 7120 8188
rect 7120 8132 7176 8188
rect 7176 8132 7180 8188
rect 7116 8128 7180 8132
rect 7196 8188 7260 8192
rect 7196 8132 7200 8188
rect 7200 8132 7256 8188
rect 7256 8132 7260 8188
rect 7196 8128 7260 8132
rect 7276 8188 7340 8192
rect 7276 8132 7280 8188
rect 7280 8132 7336 8188
rect 7336 8132 7340 8188
rect 7276 8128 7340 8132
rect 7356 8188 7420 8192
rect 7356 8132 7360 8188
rect 7360 8132 7416 8188
rect 7416 8132 7420 8188
rect 7356 8128 7420 8132
rect 13832 8188 13896 8192
rect 13832 8132 13836 8188
rect 13836 8132 13892 8188
rect 13892 8132 13896 8188
rect 13832 8128 13896 8132
rect 13912 8188 13976 8192
rect 13912 8132 13916 8188
rect 13916 8132 13972 8188
rect 13972 8132 13976 8188
rect 13912 8128 13976 8132
rect 13992 8188 14056 8192
rect 13992 8132 13996 8188
rect 13996 8132 14052 8188
rect 14052 8132 14056 8188
rect 13992 8128 14056 8132
rect 14072 8188 14136 8192
rect 14072 8132 14076 8188
rect 14076 8132 14132 8188
rect 14132 8132 14136 8188
rect 14072 8128 14136 8132
rect 20548 8188 20612 8192
rect 20548 8132 20552 8188
rect 20552 8132 20608 8188
rect 20608 8132 20612 8188
rect 20548 8128 20612 8132
rect 20628 8188 20692 8192
rect 20628 8132 20632 8188
rect 20632 8132 20688 8188
rect 20688 8132 20692 8188
rect 20628 8128 20692 8132
rect 20708 8188 20772 8192
rect 20708 8132 20712 8188
rect 20712 8132 20768 8188
rect 20768 8132 20772 8188
rect 20708 8128 20772 8132
rect 20788 8188 20852 8192
rect 20788 8132 20792 8188
rect 20792 8132 20848 8188
rect 20848 8132 20852 8188
rect 20788 8128 20852 8132
rect 27264 8188 27328 8192
rect 27264 8132 27268 8188
rect 27268 8132 27324 8188
rect 27324 8132 27328 8188
rect 27264 8128 27328 8132
rect 27344 8188 27408 8192
rect 27344 8132 27348 8188
rect 27348 8132 27404 8188
rect 27404 8132 27408 8188
rect 27344 8128 27408 8132
rect 27424 8188 27488 8192
rect 27424 8132 27428 8188
rect 27428 8132 27484 8188
rect 27484 8132 27488 8188
rect 27424 8128 27488 8132
rect 27504 8188 27568 8192
rect 27504 8132 27508 8188
rect 27508 8132 27564 8188
rect 27564 8132 27568 8188
rect 27504 8128 27568 8132
rect 3758 7644 3822 7648
rect 3758 7588 3762 7644
rect 3762 7588 3818 7644
rect 3818 7588 3822 7644
rect 3758 7584 3822 7588
rect 3838 7644 3902 7648
rect 3838 7588 3842 7644
rect 3842 7588 3898 7644
rect 3898 7588 3902 7644
rect 3838 7584 3902 7588
rect 3918 7644 3982 7648
rect 3918 7588 3922 7644
rect 3922 7588 3978 7644
rect 3978 7588 3982 7644
rect 3918 7584 3982 7588
rect 3998 7644 4062 7648
rect 3998 7588 4002 7644
rect 4002 7588 4058 7644
rect 4058 7588 4062 7644
rect 3998 7584 4062 7588
rect 10474 7644 10538 7648
rect 10474 7588 10478 7644
rect 10478 7588 10534 7644
rect 10534 7588 10538 7644
rect 10474 7584 10538 7588
rect 10554 7644 10618 7648
rect 10554 7588 10558 7644
rect 10558 7588 10614 7644
rect 10614 7588 10618 7644
rect 10554 7584 10618 7588
rect 10634 7644 10698 7648
rect 10634 7588 10638 7644
rect 10638 7588 10694 7644
rect 10694 7588 10698 7644
rect 10634 7584 10698 7588
rect 10714 7644 10778 7648
rect 10714 7588 10718 7644
rect 10718 7588 10774 7644
rect 10774 7588 10778 7644
rect 10714 7584 10778 7588
rect 17190 7644 17254 7648
rect 17190 7588 17194 7644
rect 17194 7588 17250 7644
rect 17250 7588 17254 7644
rect 17190 7584 17254 7588
rect 17270 7644 17334 7648
rect 17270 7588 17274 7644
rect 17274 7588 17330 7644
rect 17330 7588 17334 7644
rect 17270 7584 17334 7588
rect 17350 7644 17414 7648
rect 17350 7588 17354 7644
rect 17354 7588 17410 7644
rect 17410 7588 17414 7644
rect 17350 7584 17414 7588
rect 17430 7644 17494 7648
rect 17430 7588 17434 7644
rect 17434 7588 17490 7644
rect 17490 7588 17494 7644
rect 17430 7584 17494 7588
rect 23906 7644 23970 7648
rect 23906 7588 23910 7644
rect 23910 7588 23966 7644
rect 23966 7588 23970 7644
rect 23906 7584 23970 7588
rect 23986 7644 24050 7648
rect 23986 7588 23990 7644
rect 23990 7588 24046 7644
rect 24046 7588 24050 7644
rect 23986 7584 24050 7588
rect 24066 7644 24130 7648
rect 24066 7588 24070 7644
rect 24070 7588 24126 7644
rect 24126 7588 24130 7644
rect 24066 7584 24130 7588
rect 24146 7644 24210 7648
rect 24146 7588 24150 7644
rect 24150 7588 24206 7644
rect 24206 7588 24210 7644
rect 24146 7584 24210 7588
rect 7116 7100 7180 7104
rect 7116 7044 7120 7100
rect 7120 7044 7176 7100
rect 7176 7044 7180 7100
rect 7116 7040 7180 7044
rect 7196 7100 7260 7104
rect 7196 7044 7200 7100
rect 7200 7044 7256 7100
rect 7256 7044 7260 7100
rect 7196 7040 7260 7044
rect 7276 7100 7340 7104
rect 7276 7044 7280 7100
rect 7280 7044 7336 7100
rect 7336 7044 7340 7100
rect 7276 7040 7340 7044
rect 7356 7100 7420 7104
rect 7356 7044 7360 7100
rect 7360 7044 7416 7100
rect 7416 7044 7420 7100
rect 7356 7040 7420 7044
rect 13832 7100 13896 7104
rect 13832 7044 13836 7100
rect 13836 7044 13892 7100
rect 13892 7044 13896 7100
rect 13832 7040 13896 7044
rect 13912 7100 13976 7104
rect 13912 7044 13916 7100
rect 13916 7044 13972 7100
rect 13972 7044 13976 7100
rect 13912 7040 13976 7044
rect 13992 7100 14056 7104
rect 13992 7044 13996 7100
rect 13996 7044 14052 7100
rect 14052 7044 14056 7100
rect 13992 7040 14056 7044
rect 14072 7100 14136 7104
rect 14072 7044 14076 7100
rect 14076 7044 14132 7100
rect 14132 7044 14136 7100
rect 14072 7040 14136 7044
rect 20548 7100 20612 7104
rect 20548 7044 20552 7100
rect 20552 7044 20608 7100
rect 20608 7044 20612 7100
rect 20548 7040 20612 7044
rect 20628 7100 20692 7104
rect 20628 7044 20632 7100
rect 20632 7044 20688 7100
rect 20688 7044 20692 7100
rect 20628 7040 20692 7044
rect 20708 7100 20772 7104
rect 20708 7044 20712 7100
rect 20712 7044 20768 7100
rect 20768 7044 20772 7100
rect 20708 7040 20772 7044
rect 20788 7100 20852 7104
rect 20788 7044 20792 7100
rect 20792 7044 20848 7100
rect 20848 7044 20852 7100
rect 20788 7040 20852 7044
rect 27264 7100 27328 7104
rect 27264 7044 27268 7100
rect 27268 7044 27324 7100
rect 27324 7044 27328 7100
rect 27264 7040 27328 7044
rect 27344 7100 27408 7104
rect 27344 7044 27348 7100
rect 27348 7044 27404 7100
rect 27404 7044 27408 7100
rect 27344 7040 27408 7044
rect 27424 7100 27488 7104
rect 27424 7044 27428 7100
rect 27428 7044 27484 7100
rect 27484 7044 27488 7100
rect 27424 7040 27488 7044
rect 27504 7100 27568 7104
rect 27504 7044 27508 7100
rect 27508 7044 27564 7100
rect 27564 7044 27568 7100
rect 27504 7040 27568 7044
rect 3758 6556 3822 6560
rect 3758 6500 3762 6556
rect 3762 6500 3818 6556
rect 3818 6500 3822 6556
rect 3758 6496 3822 6500
rect 3838 6556 3902 6560
rect 3838 6500 3842 6556
rect 3842 6500 3898 6556
rect 3898 6500 3902 6556
rect 3838 6496 3902 6500
rect 3918 6556 3982 6560
rect 3918 6500 3922 6556
rect 3922 6500 3978 6556
rect 3978 6500 3982 6556
rect 3918 6496 3982 6500
rect 3998 6556 4062 6560
rect 3998 6500 4002 6556
rect 4002 6500 4058 6556
rect 4058 6500 4062 6556
rect 3998 6496 4062 6500
rect 10474 6556 10538 6560
rect 10474 6500 10478 6556
rect 10478 6500 10534 6556
rect 10534 6500 10538 6556
rect 10474 6496 10538 6500
rect 10554 6556 10618 6560
rect 10554 6500 10558 6556
rect 10558 6500 10614 6556
rect 10614 6500 10618 6556
rect 10554 6496 10618 6500
rect 10634 6556 10698 6560
rect 10634 6500 10638 6556
rect 10638 6500 10694 6556
rect 10694 6500 10698 6556
rect 10634 6496 10698 6500
rect 10714 6556 10778 6560
rect 10714 6500 10718 6556
rect 10718 6500 10774 6556
rect 10774 6500 10778 6556
rect 10714 6496 10778 6500
rect 17190 6556 17254 6560
rect 17190 6500 17194 6556
rect 17194 6500 17250 6556
rect 17250 6500 17254 6556
rect 17190 6496 17254 6500
rect 17270 6556 17334 6560
rect 17270 6500 17274 6556
rect 17274 6500 17330 6556
rect 17330 6500 17334 6556
rect 17270 6496 17334 6500
rect 17350 6556 17414 6560
rect 17350 6500 17354 6556
rect 17354 6500 17410 6556
rect 17410 6500 17414 6556
rect 17350 6496 17414 6500
rect 17430 6556 17494 6560
rect 17430 6500 17434 6556
rect 17434 6500 17490 6556
rect 17490 6500 17494 6556
rect 17430 6496 17494 6500
rect 23906 6556 23970 6560
rect 23906 6500 23910 6556
rect 23910 6500 23966 6556
rect 23966 6500 23970 6556
rect 23906 6496 23970 6500
rect 23986 6556 24050 6560
rect 23986 6500 23990 6556
rect 23990 6500 24046 6556
rect 24046 6500 24050 6556
rect 23986 6496 24050 6500
rect 24066 6556 24130 6560
rect 24066 6500 24070 6556
rect 24070 6500 24126 6556
rect 24126 6500 24130 6556
rect 24066 6496 24130 6500
rect 24146 6556 24210 6560
rect 24146 6500 24150 6556
rect 24150 6500 24206 6556
rect 24206 6500 24210 6556
rect 24146 6496 24210 6500
rect 7116 6012 7180 6016
rect 7116 5956 7120 6012
rect 7120 5956 7176 6012
rect 7176 5956 7180 6012
rect 7116 5952 7180 5956
rect 7196 6012 7260 6016
rect 7196 5956 7200 6012
rect 7200 5956 7256 6012
rect 7256 5956 7260 6012
rect 7196 5952 7260 5956
rect 7276 6012 7340 6016
rect 7276 5956 7280 6012
rect 7280 5956 7336 6012
rect 7336 5956 7340 6012
rect 7276 5952 7340 5956
rect 7356 6012 7420 6016
rect 7356 5956 7360 6012
rect 7360 5956 7416 6012
rect 7416 5956 7420 6012
rect 7356 5952 7420 5956
rect 13832 6012 13896 6016
rect 13832 5956 13836 6012
rect 13836 5956 13892 6012
rect 13892 5956 13896 6012
rect 13832 5952 13896 5956
rect 13912 6012 13976 6016
rect 13912 5956 13916 6012
rect 13916 5956 13972 6012
rect 13972 5956 13976 6012
rect 13912 5952 13976 5956
rect 13992 6012 14056 6016
rect 13992 5956 13996 6012
rect 13996 5956 14052 6012
rect 14052 5956 14056 6012
rect 13992 5952 14056 5956
rect 14072 6012 14136 6016
rect 14072 5956 14076 6012
rect 14076 5956 14132 6012
rect 14132 5956 14136 6012
rect 14072 5952 14136 5956
rect 20548 6012 20612 6016
rect 20548 5956 20552 6012
rect 20552 5956 20608 6012
rect 20608 5956 20612 6012
rect 20548 5952 20612 5956
rect 20628 6012 20692 6016
rect 20628 5956 20632 6012
rect 20632 5956 20688 6012
rect 20688 5956 20692 6012
rect 20628 5952 20692 5956
rect 20708 6012 20772 6016
rect 20708 5956 20712 6012
rect 20712 5956 20768 6012
rect 20768 5956 20772 6012
rect 20708 5952 20772 5956
rect 20788 6012 20852 6016
rect 20788 5956 20792 6012
rect 20792 5956 20848 6012
rect 20848 5956 20852 6012
rect 20788 5952 20852 5956
rect 27264 6012 27328 6016
rect 27264 5956 27268 6012
rect 27268 5956 27324 6012
rect 27324 5956 27328 6012
rect 27264 5952 27328 5956
rect 27344 6012 27408 6016
rect 27344 5956 27348 6012
rect 27348 5956 27404 6012
rect 27404 5956 27408 6012
rect 27344 5952 27408 5956
rect 27424 6012 27488 6016
rect 27424 5956 27428 6012
rect 27428 5956 27484 6012
rect 27484 5956 27488 6012
rect 27424 5952 27488 5956
rect 27504 6012 27568 6016
rect 27504 5956 27508 6012
rect 27508 5956 27564 6012
rect 27564 5956 27568 6012
rect 27504 5952 27568 5956
rect 3758 5468 3822 5472
rect 3758 5412 3762 5468
rect 3762 5412 3818 5468
rect 3818 5412 3822 5468
rect 3758 5408 3822 5412
rect 3838 5468 3902 5472
rect 3838 5412 3842 5468
rect 3842 5412 3898 5468
rect 3898 5412 3902 5468
rect 3838 5408 3902 5412
rect 3918 5468 3982 5472
rect 3918 5412 3922 5468
rect 3922 5412 3978 5468
rect 3978 5412 3982 5468
rect 3918 5408 3982 5412
rect 3998 5468 4062 5472
rect 3998 5412 4002 5468
rect 4002 5412 4058 5468
rect 4058 5412 4062 5468
rect 3998 5408 4062 5412
rect 10474 5468 10538 5472
rect 10474 5412 10478 5468
rect 10478 5412 10534 5468
rect 10534 5412 10538 5468
rect 10474 5408 10538 5412
rect 10554 5468 10618 5472
rect 10554 5412 10558 5468
rect 10558 5412 10614 5468
rect 10614 5412 10618 5468
rect 10554 5408 10618 5412
rect 10634 5468 10698 5472
rect 10634 5412 10638 5468
rect 10638 5412 10694 5468
rect 10694 5412 10698 5468
rect 10634 5408 10698 5412
rect 10714 5468 10778 5472
rect 10714 5412 10718 5468
rect 10718 5412 10774 5468
rect 10774 5412 10778 5468
rect 10714 5408 10778 5412
rect 17190 5468 17254 5472
rect 17190 5412 17194 5468
rect 17194 5412 17250 5468
rect 17250 5412 17254 5468
rect 17190 5408 17254 5412
rect 17270 5468 17334 5472
rect 17270 5412 17274 5468
rect 17274 5412 17330 5468
rect 17330 5412 17334 5468
rect 17270 5408 17334 5412
rect 17350 5468 17414 5472
rect 17350 5412 17354 5468
rect 17354 5412 17410 5468
rect 17410 5412 17414 5468
rect 17350 5408 17414 5412
rect 17430 5468 17494 5472
rect 17430 5412 17434 5468
rect 17434 5412 17490 5468
rect 17490 5412 17494 5468
rect 17430 5408 17494 5412
rect 23906 5468 23970 5472
rect 23906 5412 23910 5468
rect 23910 5412 23966 5468
rect 23966 5412 23970 5468
rect 23906 5408 23970 5412
rect 23986 5468 24050 5472
rect 23986 5412 23990 5468
rect 23990 5412 24046 5468
rect 24046 5412 24050 5468
rect 23986 5408 24050 5412
rect 24066 5468 24130 5472
rect 24066 5412 24070 5468
rect 24070 5412 24126 5468
rect 24126 5412 24130 5468
rect 24066 5408 24130 5412
rect 24146 5468 24210 5472
rect 24146 5412 24150 5468
rect 24150 5412 24206 5468
rect 24206 5412 24210 5468
rect 24146 5408 24210 5412
rect 7116 4924 7180 4928
rect 7116 4868 7120 4924
rect 7120 4868 7176 4924
rect 7176 4868 7180 4924
rect 7116 4864 7180 4868
rect 7196 4924 7260 4928
rect 7196 4868 7200 4924
rect 7200 4868 7256 4924
rect 7256 4868 7260 4924
rect 7196 4864 7260 4868
rect 7276 4924 7340 4928
rect 7276 4868 7280 4924
rect 7280 4868 7336 4924
rect 7336 4868 7340 4924
rect 7276 4864 7340 4868
rect 7356 4924 7420 4928
rect 7356 4868 7360 4924
rect 7360 4868 7416 4924
rect 7416 4868 7420 4924
rect 7356 4864 7420 4868
rect 13832 4924 13896 4928
rect 13832 4868 13836 4924
rect 13836 4868 13892 4924
rect 13892 4868 13896 4924
rect 13832 4864 13896 4868
rect 13912 4924 13976 4928
rect 13912 4868 13916 4924
rect 13916 4868 13972 4924
rect 13972 4868 13976 4924
rect 13912 4864 13976 4868
rect 13992 4924 14056 4928
rect 13992 4868 13996 4924
rect 13996 4868 14052 4924
rect 14052 4868 14056 4924
rect 13992 4864 14056 4868
rect 14072 4924 14136 4928
rect 14072 4868 14076 4924
rect 14076 4868 14132 4924
rect 14132 4868 14136 4924
rect 14072 4864 14136 4868
rect 20548 4924 20612 4928
rect 20548 4868 20552 4924
rect 20552 4868 20608 4924
rect 20608 4868 20612 4924
rect 20548 4864 20612 4868
rect 20628 4924 20692 4928
rect 20628 4868 20632 4924
rect 20632 4868 20688 4924
rect 20688 4868 20692 4924
rect 20628 4864 20692 4868
rect 20708 4924 20772 4928
rect 20708 4868 20712 4924
rect 20712 4868 20768 4924
rect 20768 4868 20772 4924
rect 20708 4864 20772 4868
rect 20788 4924 20852 4928
rect 20788 4868 20792 4924
rect 20792 4868 20848 4924
rect 20848 4868 20852 4924
rect 20788 4864 20852 4868
rect 27264 4924 27328 4928
rect 27264 4868 27268 4924
rect 27268 4868 27324 4924
rect 27324 4868 27328 4924
rect 27264 4864 27328 4868
rect 27344 4924 27408 4928
rect 27344 4868 27348 4924
rect 27348 4868 27404 4924
rect 27404 4868 27408 4924
rect 27344 4864 27408 4868
rect 27424 4924 27488 4928
rect 27424 4868 27428 4924
rect 27428 4868 27484 4924
rect 27484 4868 27488 4924
rect 27424 4864 27488 4868
rect 27504 4924 27568 4928
rect 27504 4868 27508 4924
rect 27508 4868 27564 4924
rect 27564 4868 27568 4924
rect 27504 4864 27568 4868
rect 3758 4380 3822 4384
rect 3758 4324 3762 4380
rect 3762 4324 3818 4380
rect 3818 4324 3822 4380
rect 3758 4320 3822 4324
rect 3838 4380 3902 4384
rect 3838 4324 3842 4380
rect 3842 4324 3898 4380
rect 3898 4324 3902 4380
rect 3838 4320 3902 4324
rect 3918 4380 3982 4384
rect 3918 4324 3922 4380
rect 3922 4324 3978 4380
rect 3978 4324 3982 4380
rect 3918 4320 3982 4324
rect 3998 4380 4062 4384
rect 3998 4324 4002 4380
rect 4002 4324 4058 4380
rect 4058 4324 4062 4380
rect 3998 4320 4062 4324
rect 10474 4380 10538 4384
rect 10474 4324 10478 4380
rect 10478 4324 10534 4380
rect 10534 4324 10538 4380
rect 10474 4320 10538 4324
rect 10554 4380 10618 4384
rect 10554 4324 10558 4380
rect 10558 4324 10614 4380
rect 10614 4324 10618 4380
rect 10554 4320 10618 4324
rect 10634 4380 10698 4384
rect 10634 4324 10638 4380
rect 10638 4324 10694 4380
rect 10694 4324 10698 4380
rect 10634 4320 10698 4324
rect 10714 4380 10778 4384
rect 10714 4324 10718 4380
rect 10718 4324 10774 4380
rect 10774 4324 10778 4380
rect 10714 4320 10778 4324
rect 17190 4380 17254 4384
rect 17190 4324 17194 4380
rect 17194 4324 17250 4380
rect 17250 4324 17254 4380
rect 17190 4320 17254 4324
rect 17270 4380 17334 4384
rect 17270 4324 17274 4380
rect 17274 4324 17330 4380
rect 17330 4324 17334 4380
rect 17270 4320 17334 4324
rect 17350 4380 17414 4384
rect 17350 4324 17354 4380
rect 17354 4324 17410 4380
rect 17410 4324 17414 4380
rect 17350 4320 17414 4324
rect 17430 4380 17494 4384
rect 17430 4324 17434 4380
rect 17434 4324 17490 4380
rect 17490 4324 17494 4380
rect 17430 4320 17494 4324
rect 23906 4380 23970 4384
rect 23906 4324 23910 4380
rect 23910 4324 23966 4380
rect 23966 4324 23970 4380
rect 23906 4320 23970 4324
rect 23986 4380 24050 4384
rect 23986 4324 23990 4380
rect 23990 4324 24046 4380
rect 24046 4324 24050 4380
rect 23986 4320 24050 4324
rect 24066 4380 24130 4384
rect 24066 4324 24070 4380
rect 24070 4324 24126 4380
rect 24126 4324 24130 4380
rect 24066 4320 24130 4324
rect 24146 4380 24210 4384
rect 24146 4324 24150 4380
rect 24150 4324 24206 4380
rect 24206 4324 24210 4380
rect 24146 4320 24210 4324
rect 7116 3836 7180 3840
rect 7116 3780 7120 3836
rect 7120 3780 7176 3836
rect 7176 3780 7180 3836
rect 7116 3776 7180 3780
rect 7196 3836 7260 3840
rect 7196 3780 7200 3836
rect 7200 3780 7256 3836
rect 7256 3780 7260 3836
rect 7196 3776 7260 3780
rect 7276 3836 7340 3840
rect 7276 3780 7280 3836
rect 7280 3780 7336 3836
rect 7336 3780 7340 3836
rect 7276 3776 7340 3780
rect 7356 3836 7420 3840
rect 7356 3780 7360 3836
rect 7360 3780 7416 3836
rect 7416 3780 7420 3836
rect 7356 3776 7420 3780
rect 13832 3836 13896 3840
rect 13832 3780 13836 3836
rect 13836 3780 13892 3836
rect 13892 3780 13896 3836
rect 13832 3776 13896 3780
rect 13912 3836 13976 3840
rect 13912 3780 13916 3836
rect 13916 3780 13972 3836
rect 13972 3780 13976 3836
rect 13912 3776 13976 3780
rect 13992 3836 14056 3840
rect 13992 3780 13996 3836
rect 13996 3780 14052 3836
rect 14052 3780 14056 3836
rect 13992 3776 14056 3780
rect 14072 3836 14136 3840
rect 14072 3780 14076 3836
rect 14076 3780 14132 3836
rect 14132 3780 14136 3836
rect 14072 3776 14136 3780
rect 20548 3836 20612 3840
rect 20548 3780 20552 3836
rect 20552 3780 20608 3836
rect 20608 3780 20612 3836
rect 20548 3776 20612 3780
rect 20628 3836 20692 3840
rect 20628 3780 20632 3836
rect 20632 3780 20688 3836
rect 20688 3780 20692 3836
rect 20628 3776 20692 3780
rect 20708 3836 20772 3840
rect 20708 3780 20712 3836
rect 20712 3780 20768 3836
rect 20768 3780 20772 3836
rect 20708 3776 20772 3780
rect 20788 3836 20852 3840
rect 20788 3780 20792 3836
rect 20792 3780 20848 3836
rect 20848 3780 20852 3836
rect 20788 3776 20852 3780
rect 27264 3836 27328 3840
rect 27264 3780 27268 3836
rect 27268 3780 27324 3836
rect 27324 3780 27328 3836
rect 27264 3776 27328 3780
rect 27344 3836 27408 3840
rect 27344 3780 27348 3836
rect 27348 3780 27404 3836
rect 27404 3780 27408 3836
rect 27344 3776 27408 3780
rect 27424 3836 27488 3840
rect 27424 3780 27428 3836
rect 27428 3780 27484 3836
rect 27484 3780 27488 3836
rect 27424 3776 27488 3780
rect 27504 3836 27568 3840
rect 27504 3780 27508 3836
rect 27508 3780 27564 3836
rect 27564 3780 27568 3836
rect 27504 3776 27568 3780
rect 3758 3292 3822 3296
rect 3758 3236 3762 3292
rect 3762 3236 3818 3292
rect 3818 3236 3822 3292
rect 3758 3232 3822 3236
rect 3838 3292 3902 3296
rect 3838 3236 3842 3292
rect 3842 3236 3898 3292
rect 3898 3236 3902 3292
rect 3838 3232 3902 3236
rect 3918 3292 3982 3296
rect 3918 3236 3922 3292
rect 3922 3236 3978 3292
rect 3978 3236 3982 3292
rect 3918 3232 3982 3236
rect 3998 3292 4062 3296
rect 3998 3236 4002 3292
rect 4002 3236 4058 3292
rect 4058 3236 4062 3292
rect 3998 3232 4062 3236
rect 10474 3292 10538 3296
rect 10474 3236 10478 3292
rect 10478 3236 10534 3292
rect 10534 3236 10538 3292
rect 10474 3232 10538 3236
rect 10554 3292 10618 3296
rect 10554 3236 10558 3292
rect 10558 3236 10614 3292
rect 10614 3236 10618 3292
rect 10554 3232 10618 3236
rect 10634 3292 10698 3296
rect 10634 3236 10638 3292
rect 10638 3236 10694 3292
rect 10694 3236 10698 3292
rect 10634 3232 10698 3236
rect 10714 3292 10778 3296
rect 10714 3236 10718 3292
rect 10718 3236 10774 3292
rect 10774 3236 10778 3292
rect 10714 3232 10778 3236
rect 17190 3292 17254 3296
rect 17190 3236 17194 3292
rect 17194 3236 17250 3292
rect 17250 3236 17254 3292
rect 17190 3232 17254 3236
rect 17270 3292 17334 3296
rect 17270 3236 17274 3292
rect 17274 3236 17330 3292
rect 17330 3236 17334 3292
rect 17270 3232 17334 3236
rect 17350 3292 17414 3296
rect 17350 3236 17354 3292
rect 17354 3236 17410 3292
rect 17410 3236 17414 3292
rect 17350 3232 17414 3236
rect 17430 3292 17494 3296
rect 17430 3236 17434 3292
rect 17434 3236 17490 3292
rect 17490 3236 17494 3292
rect 17430 3232 17494 3236
rect 23906 3292 23970 3296
rect 23906 3236 23910 3292
rect 23910 3236 23966 3292
rect 23966 3236 23970 3292
rect 23906 3232 23970 3236
rect 23986 3292 24050 3296
rect 23986 3236 23990 3292
rect 23990 3236 24046 3292
rect 24046 3236 24050 3292
rect 23986 3232 24050 3236
rect 24066 3292 24130 3296
rect 24066 3236 24070 3292
rect 24070 3236 24126 3292
rect 24126 3236 24130 3292
rect 24066 3232 24130 3236
rect 24146 3292 24210 3296
rect 24146 3236 24150 3292
rect 24150 3236 24206 3292
rect 24206 3236 24210 3292
rect 24146 3232 24210 3236
rect 7116 2748 7180 2752
rect 7116 2692 7120 2748
rect 7120 2692 7176 2748
rect 7176 2692 7180 2748
rect 7116 2688 7180 2692
rect 7196 2748 7260 2752
rect 7196 2692 7200 2748
rect 7200 2692 7256 2748
rect 7256 2692 7260 2748
rect 7196 2688 7260 2692
rect 7276 2748 7340 2752
rect 7276 2692 7280 2748
rect 7280 2692 7336 2748
rect 7336 2692 7340 2748
rect 7276 2688 7340 2692
rect 7356 2748 7420 2752
rect 7356 2692 7360 2748
rect 7360 2692 7416 2748
rect 7416 2692 7420 2748
rect 7356 2688 7420 2692
rect 13832 2748 13896 2752
rect 13832 2692 13836 2748
rect 13836 2692 13892 2748
rect 13892 2692 13896 2748
rect 13832 2688 13896 2692
rect 13912 2748 13976 2752
rect 13912 2692 13916 2748
rect 13916 2692 13972 2748
rect 13972 2692 13976 2748
rect 13912 2688 13976 2692
rect 13992 2748 14056 2752
rect 13992 2692 13996 2748
rect 13996 2692 14052 2748
rect 14052 2692 14056 2748
rect 13992 2688 14056 2692
rect 14072 2748 14136 2752
rect 14072 2692 14076 2748
rect 14076 2692 14132 2748
rect 14132 2692 14136 2748
rect 14072 2688 14136 2692
rect 20548 2748 20612 2752
rect 20548 2692 20552 2748
rect 20552 2692 20608 2748
rect 20608 2692 20612 2748
rect 20548 2688 20612 2692
rect 20628 2748 20692 2752
rect 20628 2692 20632 2748
rect 20632 2692 20688 2748
rect 20688 2692 20692 2748
rect 20628 2688 20692 2692
rect 20708 2748 20772 2752
rect 20708 2692 20712 2748
rect 20712 2692 20768 2748
rect 20768 2692 20772 2748
rect 20708 2688 20772 2692
rect 20788 2748 20852 2752
rect 20788 2692 20792 2748
rect 20792 2692 20848 2748
rect 20848 2692 20852 2748
rect 20788 2688 20852 2692
rect 27264 2748 27328 2752
rect 27264 2692 27268 2748
rect 27268 2692 27324 2748
rect 27324 2692 27328 2748
rect 27264 2688 27328 2692
rect 27344 2748 27408 2752
rect 27344 2692 27348 2748
rect 27348 2692 27404 2748
rect 27404 2692 27408 2748
rect 27344 2688 27408 2692
rect 27424 2748 27488 2752
rect 27424 2692 27428 2748
rect 27428 2692 27484 2748
rect 27484 2692 27488 2748
rect 27424 2688 27488 2692
rect 27504 2748 27568 2752
rect 27504 2692 27508 2748
rect 27508 2692 27564 2748
rect 27564 2692 27568 2748
rect 27504 2688 27568 2692
rect 3758 2204 3822 2208
rect 3758 2148 3762 2204
rect 3762 2148 3818 2204
rect 3818 2148 3822 2204
rect 3758 2144 3822 2148
rect 3838 2204 3902 2208
rect 3838 2148 3842 2204
rect 3842 2148 3898 2204
rect 3898 2148 3902 2204
rect 3838 2144 3902 2148
rect 3918 2204 3982 2208
rect 3918 2148 3922 2204
rect 3922 2148 3978 2204
rect 3978 2148 3982 2204
rect 3918 2144 3982 2148
rect 3998 2204 4062 2208
rect 3998 2148 4002 2204
rect 4002 2148 4058 2204
rect 4058 2148 4062 2204
rect 3998 2144 4062 2148
rect 10474 2204 10538 2208
rect 10474 2148 10478 2204
rect 10478 2148 10534 2204
rect 10534 2148 10538 2204
rect 10474 2144 10538 2148
rect 10554 2204 10618 2208
rect 10554 2148 10558 2204
rect 10558 2148 10614 2204
rect 10614 2148 10618 2204
rect 10554 2144 10618 2148
rect 10634 2204 10698 2208
rect 10634 2148 10638 2204
rect 10638 2148 10694 2204
rect 10694 2148 10698 2204
rect 10634 2144 10698 2148
rect 10714 2204 10778 2208
rect 10714 2148 10718 2204
rect 10718 2148 10774 2204
rect 10774 2148 10778 2204
rect 10714 2144 10778 2148
rect 17190 2204 17254 2208
rect 17190 2148 17194 2204
rect 17194 2148 17250 2204
rect 17250 2148 17254 2204
rect 17190 2144 17254 2148
rect 17270 2204 17334 2208
rect 17270 2148 17274 2204
rect 17274 2148 17330 2204
rect 17330 2148 17334 2204
rect 17270 2144 17334 2148
rect 17350 2204 17414 2208
rect 17350 2148 17354 2204
rect 17354 2148 17410 2204
rect 17410 2148 17414 2204
rect 17350 2144 17414 2148
rect 17430 2204 17494 2208
rect 17430 2148 17434 2204
rect 17434 2148 17490 2204
rect 17490 2148 17494 2204
rect 17430 2144 17494 2148
rect 23906 2204 23970 2208
rect 23906 2148 23910 2204
rect 23910 2148 23966 2204
rect 23966 2148 23970 2204
rect 23906 2144 23970 2148
rect 23986 2204 24050 2208
rect 23986 2148 23990 2204
rect 23990 2148 24046 2204
rect 24046 2148 24050 2204
rect 23986 2144 24050 2148
rect 24066 2204 24130 2208
rect 24066 2148 24070 2204
rect 24070 2148 24126 2204
rect 24126 2148 24130 2204
rect 24066 2144 24130 2148
rect 24146 2204 24210 2208
rect 24146 2148 24150 2204
rect 24150 2148 24206 2204
rect 24206 2148 24210 2204
rect 24146 2144 24210 2148
rect 7116 1660 7180 1664
rect 7116 1604 7120 1660
rect 7120 1604 7176 1660
rect 7176 1604 7180 1660
rect 7116 1600 7180 1604
rect 7196 1660 7260 1664
rect 7196 1604 7200 1660
rect 7200 1604 7256 1660
rect 7256 1604 7260 1660
rect 7196 1600 7260 1604
rect 7276 1660 7340 1664
rect 7276 1604 7280 1660
rect 7280 1604 7336 1660
rect 7336 1604 7340 1660
rect 7276 1600 7340 1604
rect 7356 1660 7420 1664
rect 7356 1604 7360 1660
rect 7360 1604 7416 1660
rect 7416 1604 7420 1660
rect 7356 1600 7420 1604
rect 13832 1660 13896 1664
rect 13832 1604 13836 1660
rect 13836 1604 13892 1660
rect 13892 1604 13896 1660
rect 13832 1600 13896 1604
rect 13912 1660 13976 1664
rect 13912 1604 13916 1660
rect 13916 1604 13972 1660
rect 13972 1604 13976 1660
rect 13912 1600 13976 1604
rect 13992 1660 14056 1664
rect 13992 1604 13996 1660
rect 13996 1604 14052 1660
rect 14052 1604 14056 1660
rect 13992 1600 14056 1604
rect 14072 1660 14136 1664
rect 14072 1604 14076 1660
rect 14076 1604 14132 1660
rect 14132 1604 14136 1660
rect 14072 1600 14136 1604
rect 20548 1660 20612 1664
rect 20548 1604 20552 1660
rect 20552 1604 20608 1660
rect 20608 1604 20612 1660
rect 20548 1600 20612 1604
rect 20628 1660 20692 1664
rect 20628 1604 20632 1660
rect 20632 1604 20688 1660
rect 20688 1604 20692 1660
rect 20628 1600 20692 1604
rect 20708 1660 20772 1664
rect 20708 1604 20712 1660
rect 20712 1604 20768 1660
rect 20768 1604 20772 1660
rect 20708 1600 20772 1604
rect 20788 1660 20852 1664
rect 20788 1604 20792 1660
rect 20792 1604 20848 1660
rect 20848 1604 20852 1660
rect 20788 1600 20852 1604
rect 27264 1660 27328 1664
rect 27264 1604 27268 1660
rect 27268 1604 27324 1660
rect 27324 1604 27328 1660
rect 27264 1600 27328 1604
rect 27344 1660 27408 1664
rect 27344 1604 27348 1660
rect 27348 1604 27404 1660
rect 27404 1604 27408 1660
rect 27344 1600 27408 1604
rect 27424 1660 27488 1664
rect 27424 1604 27428 1660
rect 27428 1604 27484 1660
rect 27484 1604 27488 1660
rect 27424 1600 27488 1604
rect 27504 1660 27568 1664
rect 27504 1604 27508 1660
rect 27508 1604 27564 1660
rect 27564 1604 27568 1660
rect 27504 1600 27568 1604
rect 3758 1116 3822 1120
rect 3758 1060 3762 1116
rect 3762 1060 3818 1116
rect 3818 1060 3822 1116
rect 3758 1056 3822 1060
rect 3838 1116 3902 1120
rect 3838 1060 3842 1116
rect 3842 1060 3898 1116
rect 3898 1060 3902 1116
rect 3838 1056 3902 1060
rect 3918 1116 3982 1120
rect 3918 1060 3922 1116
rect 3922 1060 3978 1116
rect 3978 1060 3982 1116
rect 3918 1056 3982 1060
rect 3998 1116 4062 1120
rect 3998 1060 4002 1116
rect 4002 1060 4058 1116
rect 4058 1060 4062 1116
rect 3998 1056 4062 1060
rect 10474 1116 10538 1120
rect 10474 1060 10478 1116
rect 10478 1060 10534 1116
rect 10534 1060 10538 1116
rect 10474 1056 10538 1060
rect 10554 1116 10618 1120
rect 10554 1060 10558 1116
rect 10558 1060 10614 1116
rect 10614 1060 10618 1116
rect 10554 1056 10618 1060
rect 10634 1116 10698 1120
rect 10634 1060 10638 1116
rect 10638 1060 10694 1116
rect 10694 1060 10698 1116
rect 10634 1056 10698 1060
rect 10714 1116 10778 1120
rect 10714 1060 10718 1116
rect 10718 1060 10774 1116
rect 10774 1060 10778 1116
rect 10714 1056 10778 1060
rect 17190 1116 17254 1120
rect 17190 1060 17194 1116
rect 17194 1060 17250 1116
rect 17250 1060 17254 1116
rect 17190 1056 17254 1060
rect 17270 1116 17334 1120
rect 17270 1060 17274 1116
rect 17274 1060 17330 1116
rect 17330 1060 17334 1116
rect 17270 1056 17334 1060
rect 17350 1116 17414 1120
rect 17350 1060 17354 1116
rect 17354 1060 17410 1116
rect 17410 1060 17414 1116
rect 17350 1056 17414 1060
rect 17430 1116 17494 1120
rect 17430 1060 17434 1116
rect 17434 1060 17490 1116
rect 17490 1060 17494 1116
rect 17430 1056 17494 1060
rect 23906 1116 23970 1120
rect 23906 1060 23910 1116
rect 23910 1060 23966 1116
rect 23966 1060 23970 1116
rect 23906 1056 23970 1060
rect 23986 1116 24050 1120
rect 23986 1060 23990 1116
rect 23990 1060 24046 1116
rect 24046 1060 24050 1116
rect 23986 1056 24050 1060
rect 24066 1116 24130 1120
rect 24066 1060 24070 1116
rect 24070 1060 24126 1116
rect 24126 1060 24130 1116
rect 24066 1056 24130 1060
rect 24146 1116 24210 1120
rect 24146 1060 24150 1116
rect 24150 1060 24206 1116
rect 24206 1060 24210 1116
rect 24146 1056 24210 1060
rect 7116 572 7180 576
rect 7116 516 7120 572
rect 7120 516 7176 572
rect 7176 516 7180 572
rect 7116 512 7180 516
rect 7196 572 7260 576
rect 7196 516 7200 572
rect 7200 516 7256 572
rect 7256 516 7260 572
rect 7196 512 7260 516
rect 7276 572 7340 576
rect 7276 516 7280 572
rect 7280 516 7336 572
rect 7336 516 7340 572
rect 7276 512 7340 516
rect 7356 572 7420 576
rect 7356 516 7360 572
rect 7360 516 7416 572
rect 7416 516 7420 572
rect 7356 512 7420 516
rect 13832 572 13896 576
rect 13832 516 13836 572
rect 13836 516 13892 572
rect 13892 516 13896 572
rect 13832 512 13896 516
rect 13912 572 13976 576
rect 13912 516 13916 572
rect 13916 516 13972 572
rect 13972 516 13976 572
rect 13912 512 13976 516
rect 13992 572 14056 576
rect 13992 516 13996 572
rect 13996 516 14052 572
rect 14052 516 14056 572
rect 13992 512 14056 516
rect 14072 572 14136 576
rect 14072 516 14076 572
rect 14076 516 14132 572
rect 14132 516 14136 572
rect 14072 512 14136 516
rect 20548 572 20612 576
rect 20548 516 20552 572
rect 20552 516 20608 572
rect 20608 516 20612 572
rect 20548 512 20612 516
rect 20628 572 20692 576
rect 20628 516 20632 572
rect 20632 516 20688 572
rect 20688 516 20692 572
rect 20628 512 20692 516
rect 20708 572 20772 576
rect 20708 516 20712 572
rect 20712 516 20768 572
rect 20768 516 20772 572
rect 20708 512 20772 516
rect 20788 572 20852 576
rect 20788 516 20792 572
rect 20792 516 20848 572
rect 20848 516 20852 572
rect 20788 512 20852 516
rect 27264 572 27328 576
rect 27264 516 27268 572
rect 27268 516 27324 572
rect 27324 516 27328 572
rect 27264 512 27328 516
rect 27344 572 27408 576
rect 27344 516 27348 572
rect 27348 516 27404 572
rect 27404 516 27408 572
rect 27344 512 27408 516
rect 27424 572 27488 576
rect 27424 516 27428 572
rect 27428 516 27484 572
rect 27484 516 27488 572
rect 27424 512 27488 516
rect 27504 572 27568 576
rect 27504 516 27508 572
rect 27508 516 27564 572
rect 27564 516 27568 572
rect 27504 512 27568 516
<< metal4 >>
rect 3750 30496 4070 31056
rect 3750 30432 3758 30496
rect 3822 30432 3838 30496
rect 3902 30432 3918 30496
rect 3982 30432 3998 30496
rect 4062 30432 4070 30496
rect 3750 29408 4070 30432
rect 3750 29344 3758 29408
rect 3822 29344 3838 29408
rect 3902 29344 3918 29408
rect 3982 29344 3998 29408
rect 4062 29344 4070 29408
rect 3750 28320 4070 29344
rect 3750 28256 3758 28320
rect 3822 28256 3838 28320
rect 3902 28256 3918 28320
rect 3982 28256 3998 28320
rect 4062 28256 4070 28320
rect 3750 27232 4070 28256
rect 3750 27168 3758 27232
rect 3822 27168 3838 27232
rect 3902 27168 3918 27232
rect 3982 27168 3998 27232
rect 4062 27168 4070 27232
rect 3750 26144 4070 27168
rect 3750 26080 3758 26144
rect 3822 26080 3838 26144
rect 3902 26080 3918 26144
rect 3982 26080 3998 26144
rect 4062 26080 4070 26144
rect 3750 25056 4070 26080
rect 3750 24992 3758 25056
rect 3822 24992 3838 25056
rect 3902 24992 3918 25056
rect 3982 24992 3998 25056
rect 4062 24992 4070 25056
rect 3750 23968 4070 24992
rect 3750 23904 3758 23968
rect 3822 23904 3838 23968
rect 3902 23904 3918 23968
rect 3982 23904 3998 23968
rect 4062 23904 4070 23968
rect 3750 22880 4070 23904
rect 3750 22816 3758 22880
rect 3822 22816 3838 22880
rect 3902 22816 3918 22880
rect 3982 22816 3998 22880
rect 4062 22816 4070 22880
rect 3750 21792 4070 22816
rect 7108 31040 7428 31056
rect 7108 30976 7116 31040
rect 7180 30976 7196 31040
rect 7260 30976 7276 31040
rect 7340 30976 7356 31040
rect 7420 30976 7428 31040
rect 7108 29952 7428 30976
rect 7108 29888 7116 29952
rect 7180 29888 7196 29952
rect 7260 29888 7276 29952
rect 7340 29888 7356 29952
rect 7420 29888 7428 29952
rect 7108 28864 7428 29888
rect 7108 28800 7116 28864
rect 7180 28800 7196 28864
rect 7260 28800 7276 28864
rect 7340 28800 7356 28864
rect 7420 28800 7428 28864
rect 7108 27776 7428 28800
rect 7108 27712 7116 27776
rect 7180 27712 7196 27776
rect 7260 27712 7276 27776
rect 7340 27712 7356 27776
rect 7420 27712 7428 27776
rect 7108 26688 7428 27712
rect 7108 26624 7116 26688
rect 7180 26624 7196 26688
rect 7260 26624 7276 26688
rect 7340 26624 7356 26688
rect 7420 26624 7428 26688
rect 7108 25600 7428 26624
rect 7108 25536 7116 25600
rect 7180 25536 7196 25600
rect 7260 25536 7276 25600
rect 7340 25536 7356 25600
rect 7420 25536 7428 25600
rect 7108 24512 7428 25536
rect 7108 24448 7116 24512
rect 7180 24448 7196 24512
rect 7260 24448 7276 24512
rect 7340 24448 7356 24512
rect 7420 24448 7428 24512
rect 7108 23424 7428 24448
rect 7108 23360 7116 23424
rect 7180 23360 7196 23424
rect 7260 23360 7276 23424
rect 7340 23360 7356 23424
rect 7420 23360 7428 23424
rect 7108 22336 7428 23360
rect 7108 22272 7116 22336
rect 7180 22272 7196 22336
rect 7260 22272 7276 22336
rect 7340 22272 7356 22336
rect 7420 22272 7428 22336
rect 5211 21996 5277 21997
rect 5211 21932 5212 21996
rect 5276 21932 5277 21996
rect 5211 21931 5277 21932
rect 3750 21728 3758 21792
rect 3822 21728 3838 21792
rect 3902 21728 3918 21792
rect 3982 21728 3998 21792
rect 4062 21728 4070 21792
rect 3750 20704 4070 21728
rect 3750 20640 3758 20704
rect 3822 20640 3838 20704
rect 3902 20640 3918 20704
rect 3982 20640 3998 20704
rect 4062 20640 4070 20704
rect 3750 19616 4070 20640
rect 3750 19552 3758 19616
rect 3822 19552 3838 19616
rect 3902 19552 3918 19616
rect 3982 19552 3998 19616
rect 4062 19552 4070 19616
rect 3750 18528 4070 19552
rect 3750 18464 3758 18528
rect 3822 18464 3838 18528
rect 3902 18464 3918 18528
rect 3982 18464 3998 18528
rect 4062 18464 4070 18528
rect 3750 17440 4070 18464
rect 3750 17376 3758 17440
rect 3822 17376 3838 17440
rect 3902 17376 3918 17440
rect 3982 17376 3998 17440
rect 4062 17376 4070 17440
rect 3750 16352 4070 17376
rect 3750 16288 3758 16352
rect 3822 16288 3838 16352
rect 3902 16288 3918 16352
rect 3982 16288 3998 16352
rect 4062 16288 4070 16352
rect 3750 15264 4070 16288
rect 5214 15605 5274 21931
rect 7108 21248 7428 22272
rect 7108 21184 7116 21248
rect 7180 21184 7196 21248
rect 7260 21184 7276 21248
rect 7340 21184 7356 21248
rect 7420 21184 7428 21248
rect 7108 20160 7428 21184
rect 7108 20096 7116 20160
rect 7180 20096 7196 20160
rect 7260 20096 7276 20160
rect 7340 20096 7356 20160
rect 7420 20096 7428 20160
rect 7108 19072 7428 20096
rect 7108 19008 7116 19072
rect 7180 19008 7196 19072
rect 7260 19008 7276 19072
rect 7340 19008 7356 19072
rect 7420 19008 7428 19072
rect 7108 17984 7428 19008
rect 7108 17920 7116 17984
rect 7180 17920 7196 17984
rect 7260 17920 7276 17984
rect 7340 17920 7356 17984
rect 7420 17920 7428 17984
rect 7108 16896 7428 17920
rect 7108 16832 7116 16896
rect 7180 16832 7196 16896
rect 7260 16832 7276 16896
rect 7340 16832 7356 16896
rect 7420 16832 7428 16896
rect 7108 15808 7428 16832
rect 7108 15744 7116 15808
rect 7180 15744 7196 15808
rect 7260 15744 7276 15808
rect 7340 15744 7356 15808
rect 7420 15744 7428 15808
rect 5211 15604 5277 15605
rect 5211 15540 5212 15604
rect 5276 15540 5277 15604
rect 5211 15539 5277 15540
rect 3750 15200 3758 15264
rect 3822 15200 3838 15264
rect 3902 15200 3918 15264
rect 3982 15200 3998 15264
rect 4062 15200 4070 15264
rect 3750 14176 4070 15200
rect 3750 14112 3758 14176
rect 3822 14112 3838 14176
rect 3902 14112 3918 14176
rect 3982 14112 3998 14176
rect 4062 14112 4070 14176
rect 3750 13088 4070 14112
rect 3750 13024 3758 13088
rect 3822 13024 3838 13088
rect 3902 13024 3918 13088
rect 3982 13024 3998 13088
rect 4062 13024 4070 13088
rect 3750 12000 4070 13024
rect 3750 11936 3758 12000
rect 3822 11936 3838 12000
rect 3902 11936 3918 12000
rect 3982 11936 3998 12000
rect 4062 11936 4070 12000
rect 3750 10912 4070 11936
rect 3750 10848 3758 10912
rect 3822 10848 3838 10912
rect 3902 10848 3918 10912
rect 3982 10848 3998 10912
rect 4062 10848 4070 10912
rect 3750 9824 4070 10848
rect 3750 9760 3758 9824
rect 3822 9760 3838 9824
rect 3902 9760 3918 9824
rect 3982 9760 3998 9824
rect 4062 9760 4070 9824
rect 3750 8736 4070 9760
rect 3750 8672 3758 8736
rect 3822 8672 3838 8736
rect 3902 8672 3918 8736
rect 3982 8672 3998 8736
rect 4062 8672 4070 8736
rect 3750 7648 4070 8672
rect 3750 7584 3758 7648
rect 3822 7584 3838 7648
rect 3902 7584 3918 7648
rect 3982 7584 3998 7648
rect 4062 7584 4070 7648
rect 3750 6560 4070 7584
rect 3750 6496 3758 6560
rect 3822 6496 3838 6560
rect 3902 6496 3918 6560
rect 3982 6496 3998 6560
rect 4062 6496 4070 6560
rect 3750 5472 4070 6496
rect 3750 5408 3758 5472
rect 3822 5408 3838 5472
rect 3902 5408 3918 5472
rect 3982 5408 3998 5472
rect 4062 5408 4070 5472
rect 3750 4384 4070 5408
rect 3750 4320 3758 4384
rect 3822 4320 3838 4384
rect 3902 4320 3918 4384
rect 3982 4320 3998 4384
rect 4062 4320 4070 4384
rect 3750 3296 4070 4320
rect 3750 3232 3758 3296
rect 3822 3232 3838 3296
rect 3902 3232 3918 3296
rect 3982 3232 3998 3296
rect 4062 3232 4070 3296
rect 3750 2208 4070 3232
rect 3750 2144 3758 2208
rect 3822 2144 3838 2208
rect 3902 2144 3918 2208
rect 3982 2144 3998 2208
rect 4062 2144 4070 2208
rect 3750 1120 4070 2144
rect 3750 1056 3758 1120
rect 3822 1056 3838 1120
rect 3902 1056 3918 1120
rect 3982 1056 3998 1120
rect 4062 1056 4070 1120
rect 3750 496 4070 1056
rect 7108 14720 7428 15744
rect 7108 14656 7116 14720
rect 7180 14656 7196 14720
rect 7260 14656 7276 14720
rect 7340 14656 7356 14720
rect 7420 14656 7428 14720
rect 7108 13632 7428 14656
rect 7108 13568 7116 13632
rect 7180 13568 7196 13632
rect 7260 13568 7276 13632
rect 7340 13568 7356 13632
rect 7420 13568 7428 13632
rect 7108 12544 7428 13568
rect 7108 12480 7116 12544
rect 7180 12480 7196 12544
rect 7260 12480 7276 12544
rect 7340 12480 7356 12544
rect 7420 12480 7428 12544
rect 7108 11456 7428 12480
rect 7108 11392 7116 11456
rect 7180 11392 7196 11456
rect 7260 11392 7276 11456
rect 7340 11392 7356 11456
rect 7420 11392 7428 11456
rect 7108 10368 7428 11392
rect 7108 10304 7116 10368
rect 7180 10304 7196 10368
rect 7260 10304 7276 10368
rect 7340 10304 7356 10368
rect 7420 10304 7428 10368
rect 7108 9280 7428 10304
rect 7108 9216 7116 9280
rect 7180 9216 7196 9280
rect 7260 9216 7276 9280
rect 7340 9216 7356 9280
rect 7420 9216 7428 9280
rect 7108 8192 7428 9216
rect 7108 8128 7116 8192
rect 7180 8128 7196 8192
rect 7260 8128 7276 8192
rect 7340 8128 7356 8192
rect 7420 8128 7428 8192
rect 7108 7104 7428 8128
rect 7108 7040 7116 7104
rect 7180 7040 7196 7104
rect 7260 7040 7276 7104
rect 7340 7040 7356 7104
rect 7420 7040 7428 7104
rect 7108 6016 7428 7040
rect 7108 5952 7116 6016
rect 7180 5952 7196 6016
rect 7260 5952 7276 6016
rect 7340 5952 7356 6016
rect 7420 5952 7428 6016
rect 7108 4928 7428 5952
rect 7108 4864 7116 4928
rect 7180 4864 7196 4928
rect 7260 4864 7276 4928
rect 7340 4864 7356 4928
rect 7420 4864 7428 4928
rect 7108 3840 7428 4864
rect 7108 3776 7116 3840
rect 7180 3776 7196 3840
rect 7260 3776 7276 3840
rect 7340 3776 7356 3840
rect 7420 3776 7428 3840
rect 7108 2752 7428 3776
rect 7108 2688 7116 2752
rect 7180 2688 7196 2752
rect 7260 2688 7276 2752
rect 7340 2688 7356 2752
rect 7420 2688 7428 2752
rect 7108 1664 7428 2688
rect 7108 1600 7116 1664
rect 7180 1600 7196 1664
rect 7260 1600 7276 1664
rect 7340 1600 7356 1664
rect 7420 1600 7428 1664
rect 7108 576 7428 1600
rect 7108 512 7116 576
rect 7180 512 7196 576
rect 7260 512 7276 576
rect 7340 512 7356 576
rect 7420 512 7428 576
rect 7108 496 7428 512
rect 10466 30496 10786 31056
rect 10466 30432 10474 30496
rect 10538 30432 10554 30496
rect 10618 30432 10634 30496
rect 10698 30432 10714 30496
rect 10778 30432 10786 30496
rect 10466 29408 10786 30432
rect 10466 29344 10474 29408
rect 10538 29344 10554 29408
rect 10618 29344 10634 29408
rect 10698 29344 10714 29408
rect 10778 29344 10786 29408
rect 10466 28320 10786 29344
rect 10466 28256 10474 28320
rect 10538 28256 10554 28320
rect 10618 28256 10634 28320
rect 10698 28256 10714 28320
rect 10778 28256 10786 28320
rect 10466 27232 10786 28256
rect 10466 27168 10474 27232
rect 10538 27168 10554 27232
rect 10618 27168 10634 27232
rect 10698 27168 10714 27232
rect 10778 27168 10786 27232
rect 10466 26144 10786 27168
rect 10466 26080 10474 26144
rect 10538 26080 10554 26144
rect 10618 26080 10634 26144
rect 10698 26080 10714 26144
rect 10778 26080 10786 26144
rect 10466 25056 10786 26080
rect 10466 24992 10474 25056
rect 10538 24992 10554 25056
rect 10618 24992 10634 25056
rect 10698 24992 10714 25056
rect 10778 24992 10786 25056
rect 10466 23968 10786 24992
rect 10466 23904 10474 23968
rect 10538 23904 10554 23968
rect 10618 23904 10634 23968
rect 10698 23904 10714 23968
rect 10778 23904 10786 23968
rect 10466 22880 10786 23904
rect 10466 22816 10474 22880
rect 10538 22816 10554 22880
rect 10618 22816 10634 22880
rect 10698 22816 10714 22880
rect 10778 22816 10786 22880
rect 10466 21792 10786 22816
rect 13824 31040 14144 31056
rect 13824 30976 13832 31040
rect 13896 30976 13912 31040
rect 13976 30976 13992 31040
rect 14056 30976 14072 31040
rect 14136 30976 14144 31040
rect 13824 29952 14144 30976
rect 13824 29888 13832 29952
rect 13896 29888 13912 29952
rect 13976 29888 13992 29952
rect 14056 29888 14072 29952
rect 14136 29888 14144 29952
rect 13824 28864 14144 29888
rect 13824 28800 13832 28864
rect 13896 28800 13912 28864
rect 13976 28800 13992 28864
rect 14056 28800 14072 28864
rect 14136 28800 14144 28864
rect 13824 27776 14144 28800
rect 13824 27712 13832 27776
rect 13896 27712 13912 27776
rect 13976 27712 13992 27776
rect 14056 27712 14072 27776
rect 14136 27712 14144 27776
rect 13824 26688 14144 27712
rect 13824 26624 13832 26688
rect 13896 26624 13912 26688
rect 13976 26624 13992 26688
rect 14056 26624 14072 26688
rect 14136 26624 14144 26688
rect 13824 25600 14144 26624
rect 17182 30496 17502 31056
rect 17182 30432 17190 30496
rect 17254 30432 17270 30496
rect 17334 30432 17350 30496
rect 17414 30432 17430 30496
rect 17494 30432 17502 30496
rect 17182 29408 17502 30432
rect 17182 29344 17190 29408
rect 17254 29344 17270 29408
rect 17334 29344 17350 29408
rect 17414 29344 17430 29408
rect 17494 29344 17502 29408
rect 17182 28320 17502 29344
rect 17182 28256 17190 28320
rect 17254 28256 17270 28320
rect 17334 28256 17350 28320
rect 17414 28256 17430 28320
rect 17494 28256 17502 28320
rect 17182 27232 17502 28256
rect 20540 31040 20860 31056
rect 20540 30976 20548 31040
rect 20612 30976 20628 31040
rect 20692 30976 20708 31040
rect 20772 30976 20788 31040
rect 20852 30976 20860 31040
rect 20540 29952 20860 30976
rect 20540 29888 20548 29952
rect 20612 29888 20628 29952
rect 20692 29888 20708 29952
rect 20772 29888 20788 29952
rect 20852 29888 20860 29952
rect 20540 28864 20860 29888
rect 20540 28800 20548 28864
rect 20612 28800 20628 28864
rect 20692 28800 20708 28864
rect 20772 28800 20788 28864
rect 20852 28800 20860 28864
rect 20540 27776 20860 28800
rect 20540 27712 20548 27776
rect 20612 27712 20628 27776
rect 20692 27712 20708 27776
rect 20772 27712 20788 27776
rect 20852 27712 20860 27776
rect 17723 27436 17789 27437
rect 17723 27372 17724 27436
rect 17788 27372 17789 27436
rect 17723 27371 17789 27372
rect 17182 27168 17190 27232
rect 17254 27168 17270 27232
rect 17334 27168 17350 27232
rect 17414 27168 17430 27232
rect 17494 27168 17502 27232
rect 17182 26144 17502 27168
rect 17182 26080 17190 26144
rect 17254 26080 17270 26144
rect 17334 26080 17350 26144
rect 17414 26080 17430 26144
rect 17494 26080 17502 26144
rect 16619 25940 16685 25941
rect 16619 25876 16620 25940
rect 16684 25876 16685 25940
rect 16619 25875 16685 25876
rect 13824 25536 13832 25600
rect 13896 25536 13912 25600
rect 13976 25536 13992 25600
rect 14056 25536 14072 25600
rect 14136 25536 14144 25600
rect 13824 24512 14144 25536
rect 13824 24448 13832 24512
rect 13896 24448 13912 24512
rect 13976 24448 13992 24512
rect 14056 24448 14072 24512
rect 14136 24448 14144 24512
rect 13824 23424 14144 24448
rect 13824 23360 13832 23424
rect 13896 23360 13912 23424
rect 13976 23360 13992 23424
rect 14056 23360 14072 23424
rect 14136 23360 14144 23424
rect 13824 22336 14144 23360
rect 13824 22272 13832 22336
rect 13896 22272 13912 22336
rect 13976 22272 13992 22336
rect 14056 22272 14072 22336
rect 14136 22272 14144 22336
rect 11099 22132 11165 22133
rect 11099 22068 11100 22132
rect 11164 22068 11165 22132
rect 11099 22067 11165 22068
rect 10466 21728 10474 21792
rect 10538 21728 10554 21792
rect 10618 21728 10634 21792
rect 10698 21728 10714 21792
rect 10778 21728 10786 21792
rect 10466 20704 10786 21728
rect 10466 20640 10474 20704
rect 10538 20640 10554 20704
rect 10618 20640 10634 20704
rect 10698 20640 10714 20704
rect 10778 20640 10786 20704
rect 10466 19616 10786 20640
rect 10466 19552 10474 19616
rect 10538 19552 10554 19616
rect 10618 19552 10634 19616
rect 10698 19552 10714 19616
rect 10778 19552 10786 19616
rect 10466 18528 10786 19552
rect 10466 18464 10474 18528
rect 10538 18464 10554 18528
rect 10618 18464 10634 18528
rect 10698 18464 10714 18528
rect 10778 18464 10786 18528
rect 10466 17440 10786 18464
rect 11102 17917 11162 22067
rect 11283 21996 11349 21997
rect 11283 21932 11284 21996
rect 11348 21932 11349 21996
rect 11283 21931 11349 21932
rect 11099 17916 11165 17917
rect 11099 17852 11100 17916
rect 11164 17852 11165 17916
rect 11099 17851 11165 17852
rect 10466 17376 10474 17440
rect 10538 17376 10554 17440
rect 10618 17376 10634 17440
rect 10698 17376 10714 17440
rect 10778 17376 10786 17440
rect 10466 16352 10786 17376
rect 10466 16288 10474 16352
rect 10538 16288 10554 16352
rect 10618 16288 10634 16352
rect 10698 16288 10714 16352
rect 10778 16288 10786 16352
rect 10466 15264 10786 16288
rect 10466 15200 10474 15264
rect 10538 15200 10554 15264
rect 10618 15200 10634 15264
rect 10698 15200 10714 15264
rect 10778 15200 10786 15264
rect 10466 14176 10786 15200
rect 11286 15197 11346 21931
rect 13824 21248 14144 22272
rect 13824 21184 13832 21248
rect 13896 21184 13912 21248
rect 13976 21184 13992 21248
rect 14056 21184 14072 21248
rect 14136 21184 14144 21248
rect 13824 20160 14144 21184
rect 13824 20096 13832 20160
rect 13896 20096 13912 20160
rect 13976 20096 13992 20160
rect 14056 20096 14072 20160
rect 14136 20096 14144 20160
rect 12571 19412 12637 19413
rect 12571 19348 12572 19412
rect 12636 19348 12637 19412
rect 12571 19347 12637 19348
rect 12574 16693 12634 19347
rect 13824 19072 14144 20096
rect 16067 19820 16133 19821
rect 16067 19756 16068 19820
rect 16132 19756 16133 19820
rect 16067 19755 16133 19756
rect 13824 19008 13832 19072
rect 13896 19008 13912 19072
rect 13976 19008 13992 19072
rect 14056 19008 14072 19072
rect 14136 19008 14144 19072
rect 13824 17984 14144 19008
rect 13824 17920 13832 17984
rect 13896 17920 13912 17984
rect 13976 17920 13992 17984
rect 14056 17920 14072 17984
rect 14136 17920 14144 17984
rect 13824 16896 14144 17920
rect 13824 16832 13832 16896
rect 13896 16832 13912 16896
rect 13976 16832 13992 16896
rect 14056 16832 14072 16896
rect 14136 16832 14144 16896
rect 12571 16692 12637 16693
rect 12571 16628 12572 16692
rect 12636 16628 12637 16692
rect 12571 16627 12637 16628
rect 11283 15196 11349 15197
rect 11283 15132 11284 15196
rect 11348 15132 11349 15196
rect 11283 15131 11349 15132
rect 10466 14112 10474 14176
rect 10538 14112 10554 14176
rect 10618 14112 10634 14176
rect 10698 14112 10714 14176
rect 10778 14112 10786 14176
rect 10466 13088 10786 14112
rect 12574 13973 12634 16627
rect 13824 15808 14144 16832
rect 16070 16693 16130 19755
rect 16622 19277 16682 25875
rect 17182 25056 17502 26080
rect 17726 25941 17786 27371
rect 20540 26688 20860 27712
rect 20540 26624 20548 26688
rect 20612 26624 20628 26688
rect 20692 26624 20708 26688
rect 20772 26624 20788 26688
rect 20852 26624 20860 26688
rect 17723 25940 17789 25941
rect 17723 25876 17724 25940
rect 17788 25876 17789 25940
rect 17723 25875 17789 25876
rect 17182 24992 17190 25056
rect 17254 24992 17270 25056
rect 17334 24992 17350 25056
rect 17414 24992 17430 25056
rect 17494 24992 17502 25056
rect 17182 23968 17502 24992
rect 17182 23904 17190 23968
rect 17254 23904 17270 23968
rect 17334 23904 17350 23968
rect 17414 23904 17430 23968
rect 17494 23904 17502 23968
rect 17182 22880 17502 23904
rect 17182 22816 17190 22880
rect 17254 22816 17270 22880
rect 17334 22816 17350 22880
rect 17414 22816 17430 22880
rect 17494 22816 17502 22880
rect 17182 21792 17502 22816
rect 17182 21728 17190 21792
rect 17254 21728 17270 21792
rect 17334 21728 17350 21792
rect 17414 21728 17430 21792
rect 17494 21728 17502 21792
rect 17182 20704 17502 21728
rect 17182 20640 17190 20704
rect 17254 20640 17270 20704
rect 17334 20640 17350 20704
rect 17414 20640 17430 20704
rect 17494 20640 17502 20704
rect 17182 19616 17502 20640
rect 17182 19552 17190 19616
rect 17254 19552 17270 19616
rect 17334 19552 17350 19616
rect 17414 19552 17430 19616
rect 17494 19552 17502 19616
rect 16619 19276 16685 19277
rect 16619 19212 16620 19276
rect 16684 19212 16685 19276
rect 16619 19211 16685 19212
rect 17182 18528 17502 19552
rect 17726 19277 17786 25875
rect 17907 25668 17973 25669
rect 17907 25604 17908 25668
rect 17972 25604 17973 25668
rect 17907 25603 17973 25604
rect 17910 23629 17970 25603
rect 20540 25600 20860 26624
rect 20540 25536 20548 25600
rect 20612 25536 20628 25600
rect 20692 25536 20708 25600
rect 20772 25536 20788 25600
rect 20852 25536 20860 25600
rect 20540 24512 20860 25536
rect 20540 24448 20548 24512
rect 20612 24448 20628 24512
rect 20692 24448 20708 24512
rect 20772 24448 20788 24512
rect 20852 24448 20860 24512
rect 17907 23628 17973 23629
rect 17907 23564 17908 23628
rect 17972 23564 17973 23628
rect 17907 23563 17973 23564
rect 17723 19276 17789 19277
rect 17723 19212 17724 19276
rect 17788 19212 17789 19276
rect 17723 19211 17789 19212
rect 17182 18464 17190 18528
rect 17254 18464 17270 18528
rect 17334 18464 17350 18528
rect 17414 18464 17430 18528
rect 17494 18464 17502 18528
rect 17182 17440 17502 18464
rect 17910 18325 17970 23563
rect 20540 23424 20860 24448
rect 20540 23360 20548 23424
rect 20612 23360 20628 23424
rect 20692 23360 20708 23424
rect 20772 23360 20788 23424
rect 20852 23360 20860 23424
rect 20540 22336 20860 23360
rect 20540 22272 20548 22336
rect 20612 22272 20628 22336
rect 20692 22272 20708 22336
rect 20772 22272 20788 22336
rect 20852 22272 20860 22336
rect 20540 21248 20860 22272
rect 20540 21184 20548 21248
rect 20612 21184 20628 21248
rect 20692 21184 20708 21248
rect 20772 21184 20788 21248
rect 20852 21184 20860 21248
rect 20540 20160 20860 21184
rect 20540 20096 20548 20160
rect 20612 20096 20628 20160
rect 20692 20096 20708 20160
rect 20772 20096 20788 20160
rect 20852 20096 20860 20160
rect 20540 19072 20860 20096
rect 20540 19008 20548 19072
rect 20612 19008 20628 19072
rect 20692 19008 20708 19072
rect 20772 19008 20788 19072
rect 20852 19008 20860 19072
rect 17907 18324 17973 18325
rect 17907 18260 17908 18324
rect 17972 18260 17973 18324
rect 17907 18259 17973 18260
rect 17182 17376 17190 17440
rect 17254 17376 17270 17440
rect 17334 17376 17350 17440
rect 17414 17376 17430 17440
rect 17494 17376 17502 17440
rect 16067 16692 16133 16693
rect 16067 16628 16068 16692
rect 16132 16628 16133 16692
rect 16067 16627 16133 16628
rect 13824 15744 13832 15808
rect 13896 15744 13912 15808
rect 13976 15744 13992 15808
rect 14056 15744 14072 15808
rect 14136 15744 14144 15808
rect 13824 14720 14144 15744
rect 13824 14656 13832 14720
rect 13896 14656 13912 14720
rect 13976 14656 13992 14720
rect 14056 14656 14072 14720
rect 14136 14656 14144 14720
rect 12571 13972 12637 13973
rect 12571 13908 12572 13972
rect 12636 13908 12637 13972
rect 12571 13907 12637 13908
rect 10466 13024 10474 13088
rect 10538 13024 10554 13088
rect 10618 13024 10634 13088
rect 10698 13024 10714 13088
rect 10778 13024 10786 13088
rect 10466 12000 10786 13024
rect 10466 11936 10474 12000
rect 10538 11936 10554 12000
rect 10618 11936 10634 12000
rect 10698 11936 10714 12000
rect 10778 11936 10786 12000
rect 10466 10912 10786 11936
rect 10466 10848 10474 10912
rect 10538 10848 10554 10912
rect 10618 10848 10634 10912
rect 10698 10848 10714 10912
rect 10778 10848 10786 10912
rect 10466 9824 10786 10848
rect 10466 9760 10474 9824
rect 10538 9760 10554 9824
rect 10618 9760 10634 9824
rect 10698 9760 10714 9824
rect 10778 9760 10786 9824
rect 10466 8736 10786 9760
rect 10466 8672 10474 8736
rect 10538 8672 10554 8736
rect 10618 8672 10634 8736
rect 10698 8672 10714 8736
rect 10778 8672 10786 8736
rect 10466 7648 10786 8672
rect 10466 7584 10474 7648
rect 10538 7584 10554 7648
rect 10618 7584 10634 7648
rect 10698 7584 10714 7648
rect 10778 7584 10786 7648
rect 10466 6560 10786 7584
rect 10466 6496 10474 6560
rect 10538 6496 10554 6560
rect 10618 6496 10634 6560
rect 10698 6496 10714 6560
rect 10778 6496 10786 6560
rect 10466 5472 10786 6496
rect 10466 5408 10474 5472
rect 10538 5408 10554 5472
rect 10618 5408 10634 5472
rect 10698 5408 10714 5472
rect 10778 5408 10786 5472
rect 10466 4384 10786 5408
rect 10466 4320 10474 4384
rect 10538 4320 10554 4384
rect 10618 4320 10634 4384
rect 10698 4320 10714 4384
rect 10778 4320 10786 4384
rect 10466 3296 10786 4320
rect 10466 3232 10474 3296
rect 10538 3232 10554 3296
rect 10618 3232 10634 3296
rect 10698 3232 10714 3296
rect 10778 3232 10786 3296
rect 10466 2208 10786 3232
rect 10466 2144 10474 2208
rect 10538 2144 10554 2208
rect 10618 2144 10634 2208
rect 10698 2144 10714 2208
rect 10778 2144 10786 2208
rect 10466 1120 10786 2144
rect 10466 1056 10474 1120
rect 10538 1056 10554 1120
rect 10618 1056 10634 1120
rect 10698 1056 10714 1120
rect 10778 1056 10786 1120
rect 10466 496 10786 1056
rect 13824 13632 14144 14656
rect 13824 13568 13832 13632
rect 13896 13568 13912 13632
rect 13976 13568 13992 13632
rect 14056 13568 14072 13632
rect 14136 13568 14144 13632
rect 13824 12544 14144 13568
rect 13824 12480 13832 12544
rect 13896 12480 13912 12544
rect 13976 12480 13992 12544
rect 14056 12480 14072 12544
rect 14136 12480 14144 12544
rect 13824 11456 14144 12480
rect 13824 11392 13832 11456
rect 13896 11392 13912 11456
rect 13976 11392 13992 11456
rect 14056 11392 14072 11456
rect 14136 11392 14144 11456
rect 13824 10368 14144 11392
rect 13824 10304 13832 10368
rect 13896 10304 13912 10368
rect 13976 10304 13992 10368
rect 14056 10304 14072 10368
rect 14136 10304 14144 10368
rect 13824 9280 14144 10304
rect 13824 9216 13832 9280
rect 13896 9216 13912 9280
rect 13976 9216 13992 9280
rect 14056 9216 14072 9280
rect 14136 9216 14144 9280
rect 13824 8192 14144 9216
rect 13824 8128 13832 8192
rect 13896 8128 13912 8192
rect 13976 8128 13992 8192
rect 14056 8128 14072 8192
rect 14136 8128 14144 8192
rect 13824 7104 14144 8128
rect 13824 7040 13832 7104
rect 13896 7040 13912 7104
rect 13976 7040 13992 7104
rect 14056 7040 14072 7104
rect 14136 7040 14144 7104
rect 13824 6016 14144 7040
rect 13824 5952 13832 6016
rect 13896 5952 13912 6016
rect 13976 5952 13992 6016
rect 14056 5952 14072 6016
rect 14136 5952 14144 6016
rect 13824 4928 14144 5952
rect 13824 4864 13832 4928
rect 13896 4864 13912 4928
rect 13976 4864 13992 4928
rect 14056 4864 14072 4928
rect 14136 4864 14144 4928
rect 13824 3840 14144 4864
rect 13824 3776 13832 3840
rect 13896 3776 13912 3840
rect 13976 3776 13992 3840
rect 14056 3776 14072 3840
rect 14136 3776 14144 3840
rect 13824 2752 14144 3776
rect 13824 2688 13832 2752
rect 13896 2688 13912 2752
rect 13976 2688 13992 2752
rect 14056 2688 14072 2752
rect 14136 2688 14144 2752
rect 13824 1664 14144 2688
rect 13824 1600 13832 1664
rect 13896 1600 13912 1664
rect 13976 1600 13992 1664
rect 14056 1600 14072 1664
rect 14136 1600 14144 1664
rect 13824 576 14144 1600
rect 13824 512 13832 576
rect 13896 512 13912 576
rect 13976 512 13992 576
rect 14056 512 14072 576
rect 14136 512 14144 576
rect 13824 496 14144 512
rect 17182 16352 17502 17376
rect 17182 16288 17190 16352
rect 17254 16288 17270 16352
rect 17334 16288 17350 16352
rect 17414 16288 17430 16352
rect 17494 16288 17502 16352
rect 17182 15264 17502 16288
rect 17182 15200 17190 15264
rect 17254 15200 17270 15264
rect 17334 15200 17350 15264
rect 17414 15200 17430 15264
rect 17494 15200 17502 15264
rect 17182 14176 17502 15200
rect 17182 14112 17190 14176
rect 17254 14112 17270 14176
rect 17334 14112 17350 14176
rect 17414 14112 17430 14176
rect 17494 14112 17502 14176
rect 17182 13088 17502 14112
rect 17182 13024 17190 13088
rect 17254 13024 17270 13088
rect 17334 13024 17350 13088
rect 17414 13024 17430 13088
rect 17494 13024 17502 13088
rect 17182 12000 17502 13024
rect 17182 11936 17190 12000
rect 17254 11936 17270 12000
rect 17334 11936 17350 12000
rect 17414 11936 17430 12000
rect 17494 11936 17502 12000
rect 17182 10912 17502 11936
rect 17182 10848 17190 10912
rect 17254 10848 17270 10912
rect 17334 10848 17350 10912
rect 17414 10848 17430 10912
rect 17494 10848 17502 10912
rect 17182 9824 17502 10848
rect 17182 9760 17190 9824
rect 17254 9760 17270 9824
rect 17334 9760 17350 9824
rect 17414 9760 17430 9824
rect 17494 9760 17502 9824
rect 17182 8736 17502 9760
rect 17182 8672 17190 8736
rect 17254 8672 17270 8736
rect 17334 8672 17350 8736
rect 17414 8672 17430 8736
rect 17494 8672 17502 8736
rect 17182 7648 17502 8672
rect 17182 7584 17190 7648
rect 17254 7584 17270 7648
rect 17334 7584 17350 7648
rect 17414 7584 17430 7648
rect 17494 7584 17502 7648
rect 17182 6560 17502 7584
rect 17182 6496 17190 6560
rect 17254 6496 17270 6560
rect 17334 6496 17350 6560
rect 17414 6496 17430 6560
rect 17494 6496 17502 6560
rect 17182 5472 17502 6496
rect 17182 5408 17190 5472
rect 17254 5408 17270 5472
rect 17334 5408 17350 5472
rect 17414 5408 17430 5472
rect 17494 5408 17502 5472
rect 17182 4384 17502 5408
rect 17182 4320 17190 4384
rect 17254 4320 17270 4384
rect 17334 4320 17350 4384
rect 17414 4320 17430 4384
rect 17494 4320 17502 4384
rect 17182 3296 17502 4320
rect 17182 3232 17190 3296
rect 17254 3232 17270 3296
rect 17334 3232 17350 3296
rect 17414 3232 17430 3296
rect 17494 3232 17502 3296
rect 17182 2208 17502 3232
rect 17182 2144 17190 2208
rect 17254 2144 17270 2208
rect 17334 2144 17350 2208
rect 17414 2144 17430 2208
rect 17494 2144 17502 2208
rect 17182 1120 17502 2144
rect 17182 1056 17190 1120
rect 17254 1056 17270 1120
rect 17334 1056 17350 1120
rect 17414 1056 17430 1120
rect 17494 1056 17502 1120
rect 17182 496 17502 1056
rect 20540 17984 20860 19008
rect 20540 17920 20548 17984
rect 20612 17920 20628 17984
rect 20692 17920 20708 17984
rect 20772 17920 20788 17984
rect 20852 17920 20860 17984
rect 20540 16896 20860 17920
rect 20540 16832 20548 16896
rect 20612 16832 20628 16896
rect 20692 16832 20708 16896
rect 20772 16832 20788 16896
rect 20852 16832 20860 16896
rect 20540 15808 20860 16832
rect 20540 15744 20548 15808
rect 20612 15744 20628 15808
rect 20692 15744 20708 15808
rect 20772 15744 20788 15808
rect 20852 15744 20860 15808
rect 20540 14720 20860 15744
rect 20540 14656 20548 14720
rect 20612 14656 20628 14720
rect 20692 14656 20708 14720
rect 20772 14656 20788 14720
rect 20852 14656 20860 14720
rect 20540 13632 20860 14656
rect 20540 13568 20548 13632
rect 20612 13568 20628 13632
rect 20692 13568 20708 13632
rect 20772 13568 20788 13632
rect 20852 13568 20860 13632
rect 20540 12544 20860 13568
rect 20540 12480 20548 12544
rect 20612 12480 20628 12544
rect 20692 12480 20708 12544
rect 20772 12480 20788 12544
rect 20852 12480 20860 12544
rect 20540 11456 20860 12480
rect 20540 11392 20548 11456
rect 20612 11392 20628 11456
rect 20692 11392 20708 11456
rect 20772 11392 20788 11456
rect 20852 11392 20860 11456
rect 20540 10368 20860 11392
rect 20540 10304 20548 10368
rect 20612 10304 20628 10368
rect 20692 10304 20708 10368
rect 20772 10304 20788 10368
rect 20852 10304 20860 10368
rect 20540 9280 20860 10304
rect 20540 9216 20548 9280
rect 20612 9216 20628 9280
rect 20692 9216 20708 9280
rect 20772 9216 20788 9280
rect 20852 9216 20860 9280
rect 20540 8192 20860 9216
rect 20540 8128 20548 8192
rect 20612 8128 20628 8192
rect 20692 8128 20708 8192
rect 20772 8128 20788 8192
rect 20852 8128 20860 8192
rect 20540 7104 20860 8128
rect 20540 7040 20548 7104
rect 20612 7040 20628 7104
rect 20692 7040 20708 7104
rect 20772 7040 20788 7104
rect 20852 7040 20860 7104
rect 20540 6016 20860 7040
rect 20540 5952 20548 6016
rect 20612 5952 20628 6016
rect 20692 5952 20708 6016
rect 20772 5952 20788 6016
rect 20852 5952 20860 6016
rect 20540 4928 20860 5952
rect 20540 4864 20548 4928
rect 20612 4864 20628 4928
rect 20692 4864 20708 4928
rect 20772 4864 20788 4928
rect 20852 4864 20860 4928
rect 20540 3840 20860 4864
rect 20540 3776 20548 3840
rect 20612 3776 20628 3840
rect 20692 3776 20708 3840
rect 20772 3776 20788 3840
rect 20852 3776 20860 3840
rect 20540 2752 20860 3776
rect 20540 2688 20548 2752
rect 20612 2688 20628 2752
rect 20692 2688 20708 2752
rect 20772 2688 20788 2752
rect 20852 2688 20860 2752
rect 20540 1664 20860 2688
rect 20540 1600 20548 1664
rect 20612 1600 20628 1664
rect 20692 1600 20708 1664
rect 20772 1600 20788 1664
rect 20852 1600 20860 1664
rect 20540 576 20860 1600
rect 20540 512 20548 576
rect 20612 512 20628 576
rect 20692 512 20708 576
rect 20772 512 20788 576
rect 20852 512 20860 576
rect 20540 496 20860 512
rect 23898 30496 24218 31056
rect 23898 30432 23906 30496
rect 23970 30432 23986 30496
rect 24050 30432 24066 30496
rect 24130 30432 24146 30496
rect 24210 30432 24218 30496
rect 23898 29408 24218 30432
rect 23898 29344 23906 29408
rect 23970 29344 23986 29408
rect 24050 29344 24066 29408
rect 24130 29344 24146 29408
rect 24210 29344 24218 29408
rect 23898 28320 24218 29344
rect 23898 28256 23906 28320
rect 23970 28256 23986 28320
rect 24050 28256 24066 28320
rect 24130 28256 24146 28320
rect 24210 28256 24218 28320
rect 23898 27232 24218 28256
rect 23898 27168 23906 27232
rect 23970 27168 23986 27232
rect 24050 27168 24066 27232
rect 24130 27168 24146 27232
rect 24210 27168 24218 27232
rect 23898 26144 24218 27168
rect 23898 26080 23906 26144
rect 23970 26080 23986 26144
rect 24050 26080 24066 26144
rect 24130 26080 24146 26144
rect 24210 26080 24218 26144
rect 23898 25056 24218 26080
rect 23898 24992 23906 25056
rect 23970 24992 23986 25056
rect 24050 24992 24066 25056
rect 24130 24992 24146 25056
rect 24210 24992 24218 25056
rect 23898 23968 24218 24992
rect 23898 23904 23906 23968
rect 23970 23904 23986 23968
rect 24050 23904 24066 23968
rect 24130 23904 24146 23968
rect 24210 23904 24218 23968
rect 23898 22880 24218 23904
rect 23898 22816 23906 22880
rect 23970 22816 23986 22880
rect 24050 22816 24066 22880
rect 24130 22816 24146 22880
rect 24210 22816 24218 22880
rect 23898 21792 24218 22816
rect 23898 21728 23906 21792
rect 23970 21728 23986 21792
rect 24050 21728 24066 21792
rect 24130 21728 24146 21792
rect 24210 21728 24218 21792
rect 23898 20704 24218 21728
rect 23898 20640 23906 20704
rect 23970 20640 23986 20704
rect 24050 20640 24066 20704
rect 24130 20640 24146 20704
rect 24210 20640 24218 20704
rect 23898 19616 24218 20640
rect 23898 19552 23906 19616
rect 23970 19552 23986 19616
rect 24050 19552 24066 19616
rect 24130 19552 24146 19616
rect 24210 19552 24218 19616
rect 23898 18528 24218 19552
rect 23898 18464 23906 18528
rect 23970 18464 23986 18528
rect 24050 18464 24066 18528
rect 24130 18464 24146 18528
rect 24210 18464 24218 18528
rect 23898 17440 24218 18464
rect 23898 17376 23906 17440
rect 23970 17376 23986 17440
rect 24050 17376 24066 17440
rect 24130 17376 24146 17440
rect 24210 17376 24218 17440
rect 23898 16352 24218 17376
rect 23898 16288 23906 16352
rect 23970 16288 23986 16352
rect 24050 16288 24066 16352
rect 24130 16288 24146 16352
rect 24210 16288 24218 16352
rect 23898 15264 24218 16288
rect 23898 15200 23906 15264
rect 23970 15200 23986 15264
rect 24050 15200 24066 15264
rect 24130 15200 24146 15264
rect 24210 15200 24218 15264
rect 23898 14176 24218 15200
rect 23898 14112 23906 14176
rect 23970 14112 23986 14176
rect 24050 14112 24066 14176
rect 24130 14112 24146 14176
rect 24210 14112 24218 14176
rect 23898 13088 24218 14112
rect 23898 13024 23906 13088
rect 23970 13024 23986 13088
rect 24050 13024 24066 13088
rect 24130 13024 24146 13088
rect 24210 13024 24218 13088
rect 23898 12000 24218 13024
rect 23898 11936 23906 12000
rect 23970 11936 23986 12000
rect 24050 11936 24066 12000
rect 24130 11936 24146 12000
rect 24210 11936 24218 12000
rect 23898 10912 24218 11936
rect 23898 10848 23906 10912
rect 23970 10848 23986 10912
rect 24050 10848 24066 10912
rect 24130 10848 24146 10912
rect 24210 10848 24218 10912
rect 23898 9824 24218 10848
rect 23898 9760 23906 9824
rect 23970 9760 23986 9824
rect 24050 9760 24066 9824
rect 24130 9760 24146 9824
rect 24210 9760 24218 9824
rect 23898 8736 24218 9760
rect 23898 8672 23906 8736
rect 23970 8672 23986 8736
rect 24050 8672 24066 8736
rect 24130 8672 24146 8736
rect 24210 8672 24218 8736
rect 23898 7648 24218 8672
rect 23898 7584 23906 7648
rect 23970 7584 23986 7648
rect 24050 7584 24066 7648
rect 24130 7584 24146 7648
rect 24210 7584 24218 7648
rect 23898 6560 24218 7584
rect 23898 6496 23906 6560
rect 23970 6496 23986 6560
rect 24050 6496 24066 6560
rect 24130 6496 24146 6560
rect 24210 6496 24218 6560
rect 23898 5472 24218 6496
rect 23898 5408 23906 5472
rect 23970 5408 23986 5472
rect 24050 5408 24066 5472
rect 24130 5408 24146 5472
rect 24210 5408 24218 5472
rect 23898 4384 24218 5408
rect 23898 4320 23906 4384
rect 23970 4320 23986 4384
rect 24050 4320 24066 4384
rect 24130 4320 24146 4384
rect 24210 4320 24218 4384
rect 23898 3296 24218 4320
rect 23898 3232 23906 3296
rect 23970 3232 23986 3296
rect 24050 3232 24066 3296
rect 24130 3232 24146 3296
rect 24210 3232 24218 3296
rect 23898 2208 24218 3232
rect 23898 2144 23906 2208
rect 23970 2144 23986 2208
rect 24050 2144 24066 2208
rect 24130 2144 24146 2208
rect 24210 2144 24218 2208
rect 23898 1120 24218 2144
rect 23898 1056 23906 1120
rect 23970 1056 23986 1120
rect 24050 1056 24066 1120
rect 24130 1056 24146 1120
rect 24210 1056 24218 1120
rect 23898 496 24218 1056
rect 27256 31040 27576 31056
rect 27256 30976 27264 31040
rect 27328 30976 27344 31040
rect 27408 30976 27424 31040
rect 27488 30976 27504 31040
rect 27568 30976 27576 31040
rect 27256 29952 27576 30976
rect 27256 29888 27264 29952
rect 27328 29888 27344 29952
rect 27408 29888 27424 29952
rect 27488 29888 27504 29952
rect 27568 29888 27576 29952
rect 27256 28864 27576 29888
rect 27256 28800 27264 28864
rect 27328 28800 27344 28864
rect 27408 28800 27424 28864
rect 27488 28800 27504 28864
rect 27568 28800 27576 28864
rect 27256 27776 27576 28800
rect 27256 27712 27264 27776
rect 27328 27712 27344 27776
rect 27408 27712 27424 27776
rect 27488 27712 27504 27776
rect 27568 27712 27576 27776
rect 27256 26688 27576 27712
rect 27256 26624 27264 26688
rect 27328 26624 27344 26688
rect 27408 26624 27424 26688
rect 27488 26624 27504 26688
rect 27568 26624 27576 26688
rect 27256 25600 27576 26624
rect 27256 25536 27264 25600
rect 27328 25536 27344 25600
rect 27408 25536 27424 25600
rect 27488 25536 27504 25600
rect 27568 25536 27576 25600
rect 27256 24512 27576 25536
rect 27256 24448 27264 24512
rect 27328 24448 27344 24512
rect 27408 24448 27424 24512
rect 27488 24448 27504 24512
rect 27568 24448 27576 24512
rect 27256 23424 27576 24448
rect 27256 23360 27264 23424
rect 27328 23360 27344 23424
rect 27408 23360 27424 23424
rect 27488 23360 27504 23424
rect 27568 23360 27576 23424
rect 27256 22336 27576 23360
rect 27256 22272 27264 22336
rect 27328 22272 27344 22336
rect 27408 22272 27424 22336
rect 27488 22272 27504 22336
rect 27568 22272 27576 22336
rect 27256 21248 27576 22272
rect 27256 21184 27264 21248
rect 27328 21184 27344 21248
rect 27408 21184 27424 21248
rect 27488 21184 27504 21248
rect 27568 21184 27576 21248
rect 27256 20160 27576 21184
rect 27256 20096 27264 20160
rect 27328 20096 27344 20160
rect 27408 20096 27424 20160
rect 27488 20096 27504 20160
rect 27568 20096 27576 20160
rect 27256 19072 27576 20096
rect 27256 19008 27264 19072
rect 27328 19008 27344 19072
rect 27408 19008 27424 19072
rect 27488 19008 27504 19072
rect 27568 19008 27576 19072
rect 27256 17984 27576 19008
rect 27256 17920 27264 17984
rect 27328 17920 27344 17984
rect 27408 17920 27424 17984
rect 27488 17920 27504 17984
rect 27568 17920 27576 17984
rect 27256 16896 27576 17920
rect 27256 16832 27264 16896
rect 27328 16832 27344 16896
rect 27408 16832 27424 16896
rect 27488 16832 27504 16896
rect 27568 16832 27576 16896
rect 27256 15808 27576 16832
rect 27256 15744 27264 15808
rect 27328 15744 27344 15808
rect 27408 15744 27424 15808
rect 27488 15744 27504 15808
rect 27568 15744 27576 15808
rect 27256 14720 27576 15744
rect 27256 14656 27264 14720
rect 27328 14656 27344 14720
rect 27408 14656 27424 14720
rect 27488 14656 27504 14720
rect 27568 14656 27576 14720
rect 27256 13632 27576 14656
rect 27256 13568 27264 13632
rect 27328 13568 27344 13632
rect 27408 13568 27424 13632
rect 27488 13568 27504 13632
rect 27568 13568 27576 13632
rect 27256 12544 27576 13568
rect 27256 12480 27264 12544
rect 27328 12480 27344 12544
rect 27408 12480 27424 12544
rect 27488 12480 27504 12544
rect 27568 12480 27576 12544
rect 27256 11456 27576 12480
rect 27256 11392 27264 11456
rect 27328 11392 27344 11456
rect 27408 11392 27424 11456
rect 27488 11392 27504 11456
rect 27568 11392 27576 11456
rect 27256 10368 27576 11392
rect 27256 10304 27264 10368
rect 27328 10304 27344 10368
rect 27408 10304 27424 10368
rect 27488 10304 27504 10368
rect 27568 10304 27576 10368
rect 27256 9280 27576 10304
rect 27256 9216 27264 9280
rect 27328 9216 27344 9280
rect 27408 9216 27424 9280
rect 27488 9216 27504 9280
rect 27568 9216 27576 9280
rect 27256 8192 27576 9216
rect 27256 8128 27264 8192
rect 27328 8128 27344 8192
rect 27408 8128 27424 8192
rect 27488 8128 27504 8192
rect 27568 8128 27576 8192
rect 27256 7104 27576 8128
rect 27256 7040 27264 7104
rect 27328 7040 27344 7104
rect 27408 7040 27424 7104
rect 27488 7040 27504 7104
rect 27568 7040 27576 7104
rect 27256 6016 27576 7040
rect 27256 5952 27264 6016
rect 27328 5952 27344 6016
rect 27408 5952 27424 6016
rect 27488 5952 27504 6016
rect 27568 5952 27576 6016
rect 27256 4928 27576 5952
rect 27256 4864 27264 4928
rect 27328 4864 27344 4928
rect 27408 4864 27424 4928
rect 27488 4864 27504 4928
rect 27568 4864 27576 4928
rect 27256 3840 27576 4864
rect 27256 3776 27264 3840
rect 27328 3776 27344 3840
rect 27408 3776 27424 3840
rect 27488 3776 27504 3840
rect 27568 3776 27576 3840
rect 27256 2752 27576 3776
rect 27256 2688 27264 2752
rect 27328 2688 27344 2752
rect 27408 2688 27424 2752
rect 27488 2688 27504 2752
rect 27568 2688 27576 2752
rect 27256 1664 27576 2688
rect 27256 1600 27264 1664
rect 27328 1600 27344 1664
rect 27408 1600 27424 1664
rect 27488 1600 27504 1664
rect 27568 1600 27576 1664
rect 27256 576 27576 1600
rect 27256 512 27264 576
rect 27328 512 27344 576
rect 27408 512 27424 576
rect 27488 512 27504 576
rect 27568 512 27576 576
rect 27256 496 27576 512
use sky130_fd_sc_hd__and4_1  _1052_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3036 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1053_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2116 0 1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1054_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2392 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1055_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2300 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1056_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2944 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1057_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2760 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1058_
timestamp 1704896540
transform -1 0 2392 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1059_
timestamp 1704896540
transform -1 0 2116 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1060_
timestamp 1704896540
transform 1 0 1012 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1061_
timestamp 1704896540
transform -1 0 3128 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1062_
timestamp 1704896540
transform 1 0 1748 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1063_
timestamp 1704896540
transform 1 0 2024 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1064_
timestamp 1704896540
transform -1 0 3036 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1065_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2300 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1066_
timestamp 1704896540
transform -1 0 2760 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1067_
timestamp 1704896540
transform -1 0 1932 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1068_
timestamp 1704896540
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1069_
timestamp 1704896540
transform -1 0 1840 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1070_
timestamp 1704896540
transform 1 0 2300 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1071_
timestamp 1704896540
transform -1 0 2300 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1072_
timestamp 1704896540
transform 1 0 1196 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1073_
timestamp 1704896540
transform 1 0 2024 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1074_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2944 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1075_
timestamp 1704896540
transform 1 0 2484 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1076_
timestamp 1704896540
transform -1 0 4324 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1077_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2116 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _1078_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4048 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _1079_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6716 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1080_
timestamp 1704896540
transform 1 0 7728 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1081_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6164 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1082_
timestamp 1704896540
transform 1 0 5796 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1083_
timestamp 1704896540
transform 1 0 6348 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1084_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6440 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1085_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6532 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1086_
timestamp 1704896540
transform -1 0 7452 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1087_
timestamp 1704896540
transform -1 0 7084 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1088_
timestamp 1704896540
transform -1 0 5704 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1089_
timestamp 1704896540
transform -1 0 6624 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1090_
timestamp 1704896540
transform 1 0 6900 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1091_
timestamp 1704896540
transform -1 0 5612 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1092_
timestamp 1704896540
transform 1 0 4876 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1093_
timestamp 1704896540
transform 1 0 5612 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _1094_
timestamp 1704896540
transform 1 0 6164 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1095_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 17572 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1096_
timestamp 1704896540
transform -1 0 18400 0 1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1097_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 19320 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1098_
timestamp 1704896540
transform -1 0 19320 0 1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1099_
timestamp 1704896540
transform 1 0 18676 0 -1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1100_
timestamp 1704896540
transform -1 0 18124 0 -1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1101_
timestamp 1704896540
transform 1 0 17204 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1102_
timestamp 1704896540
transform 1 0 17940 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1103_
timestamp 1704896540
transform -1 0 18308 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1104_
timestamp 1704896540
transform 1 0 18032 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1105_
timestamp 1704896540
transform 1 0 7084 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1106_
timestamp 1704896540
transform 1 0 7452 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1107_
timestamp 1704896540
transform 1 0 7544 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1108_
timestamp 1704896540
transform -1 0 8096 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1109_
timestamp 1704896540
transform 1 0 8372 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1110_
timestamp 1704896540
transform -1 0 8280 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1111_
timestamp 1704896540
transform -1 0 8096 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1112_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8004 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _1113_
timestamp 1704896540
transform 1 0 6256 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1114_
timestamp 1704896540
transform -1 0 7360 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1115_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7268 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1116_
timestamp 1704896540
transform 1 0 6624 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1117_
timestamp 1704896540
transform -1 0 6164 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1118_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6164 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1119_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5980 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1120_
timestamp 1704896540
transform 1 0 5520 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1121_
timestamp 1704896540
transform 1 0 5796 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1122_
timestamp 1704896540
transform 1 0 5060 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1123_
timestamp 1704896540
transform -1 0 4876 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1124_
timestamp 1704896540
transform -1 0 5520 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1125_
timestamp 1704896540
transform 1 0 4508 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_1  _1126_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5060 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1127_
timestamp 1704896540
transform 1 0 4048 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1128_
timestamp 1704896540
transform 1 0 4232 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1129_
timestamp 1704896540
transform -1 0 4508 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1130_
timestamp 1704896540
transform 1 0 3220 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1131_
timestamp 1704896540
transform 1 0 3036 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1132_
timestamp 1704896540
transform -1 0 3220 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1133_
timestamp 1704896540
transform -1 0 3128 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1134_
timestamp 1704896540
transform 1 0 3220 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1135_
timestamp 1704896540
transform -1 0 4140 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1136_
timestamp 1704896540
transform 1 0 2392 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1137_
timestamp 1704896540
transform -1 0 2300 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1138_
timestamp 1704896540
transform 1 0 2300 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1139_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2484 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1140_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3312 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1141_
timestamp 1704896540
transform 1 0 3220 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1142_
timestamp 1704896540
transform 1 0 2484 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1143_
timestamp 1704896540
transform 1 0 2576 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1144_
timestamp 1704896540
transform 1 0 1932 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1145_
timestamp 1704896540
transform -1 0 3680 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1146_
timestamp 1704896540
transform 1 0 2944 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _1147_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2484 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1148_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3128 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1149_
timestamp 1704896540
transform -1 0 2944 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1150_
timestamp 1704896540
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1151_
timestamp 1704896540
transform -1 0 4232 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1152_
timestamp 1704896540
transform -1 0 4692 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1153_
timestamp 1704896540
transform -1 0 4232 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1154_
timestamp 1704896540
transform -1 0 2760 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1155_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3036 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1156_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2576 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1157_
timestamp 1704896540
transform 1 0 3220 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1158_
timestamp 1704896540
transform -1 0 3588 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1159_
timestamp 1704896540
transform -1 0 15548 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1160_
timestamp 1704896540
transform -1 0 15824 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1161_
timestamp 1704896540
transform 1 0 15088 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1162_
timestamp 1704896540
transform 1 0 15548 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1163_
timestamp 1704896540
transform 1 0 17848 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1164_
timestamp 1704896540
transform -1 0 17480 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1165_
timestamp 1704896540
transform -1 0 17848 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1166_
timestamp 1704896540
transform -1 0 17204 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _1167_
timestamp 1704896540
transform -1 0 16652 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1168_
timestamp 1704896540
transform -1 0 16468 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1169_
timestamp 1704896540
transform -1 0 17388 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1170_
timestamp 1704896540
transform -1 0 17848 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1171_
timestamp 1704896540
transform -1 0 18492 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1172_
timestamp 1704896540
transform 1 0 16652 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1173_
timestamp 1704896540
transform 1 0 16468 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1174_
timestamp 1704896540
transform 1 0 15824 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1175_
timestamp 1704896540
transform 1 0 16284 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1176_
timestamp 1704896540
transform 1 0 14904 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1177_
timestamp 1704896540
transform -1 0 15640 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1178_
timestamp 1704896540
transform -1 0 15824 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1179_
timestamp 1704896540
transform 1 0 14812 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_2  _1180_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 15088 0 -1 8160
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1181_
timestamp 1704896540
transform 1 0 13984 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1182_
timestamp 1704896540
transform 1 0 14076 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1183_
timestamp 1704896540
transform 1 0 13800 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1184_
timestamp 1704896540
transform -1 0 13432 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1185_
timestamp 1704896540
transform 1 0 13524 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1186_
timestamp 1704896540
transform -1 0 13616 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1187_
timestamp 1704896540
transform 1 0 12420 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1188_
timestamp 1704896540
transform -1 0 14076 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1189_
timestamp 1704896540
transform -1 0 13340 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1190_
timestamp 1704896540
transform -1 0 12604 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1191_
timestamp 1704896540
transform -1 0 11960 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1192_
timestamp 1704896540
transform 1 0 12420 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1193_
timestamp 1704896540
transform -1 0 12420 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1194_
timestamp 1704896540
transform 1 0 12328 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1195_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11592 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1196_
timestamp 1704896540
transform -1 0 10488 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1197_
timestamp 1704896540
transform -1 0 10764 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1198_
timestamp 1704896540
transform 1 0 11960 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1199_
timestamp 1704896540
transform 1 0 9384 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_2  _1200_
timestamp 1704896540
transform 1 0 10028 0 1 5984
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1201_
timestamp 1704896540
transform 1 0 8924 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1202_
timestamp 1704896540
transform 1 0 9016 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1203_
timestamp 1704896540
transform -1 0 10488 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1204_
timestamp 1704896540
transform 1 0 10948 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1205_
timestamp 1704896540
transform -1 0 10764 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1206_
timestamp 1704896540
transform 1 0 9292 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1207_
timestamp 1704896540
transform 1 0 9936 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1208_
timestamp 1704896540
transform -1 0 9200 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1209_
timestamp 1704896540
transform -1 0 8648 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _1210_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9752 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1211_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9660 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1212_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6900 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1213_
timestamp 1704896540
transform -1 0 19780 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_2  _1214_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 18860 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1215_
timestamp 1704896540
transform 1 0 9384 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1216_
timestamp 1704896540
transform 1 0 8372 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1217_
timestamp 1704896540
transform 1 0 7084 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1218_
timestamp 1704896540
transform -1 0 9384 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_2  _1219_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8464 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1220_
timestamp 1704896540
transform 1 0 6440 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1221_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7268 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _1222_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8372 0 1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _1223_
timestamp 1704896540
transform -1 0 9936 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1224_
timestamp 1704896540
transform 1 0 7636 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1225_
timestamp 1704896540
transform 1 0 7084 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1226_
timestamp 1704896540
transform -1 0 9752 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_2  _1227_
timestamp 1704896540
transform 1 0 8648 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1228_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7544 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1229_
timestamp 1704896540
transform 1 0 2760 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1230_
timestamp 1704896540
transform -1 0 6256 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1231_
timestamp 1704896540
transform 1 0 6900 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1232_
timestamp 1704896540
transform 1 0 6256 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_2  _1233_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8740 0 1 9248
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1234_
timestamp 1704896540
transform 1 0 8832 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1235_
timestamp 1704896540
transform -1 0 7728 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1236_
timestamp 1704896540
transform -1 0 8096 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1237_
timestamp 1704896540
transform 1 0 8188 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1238_
timestamp 1704896540
transform -1 0 8096 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1239_
timestamp 1704896540
transform 1 0 7544 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1240_
timestamp 1704896540
transform -1 0 8832 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1241_
timestamp 1704896540
transform -1 0 3588 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_2  _1242_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6072 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1243_
timestamp 1704896540
transform 1 0 3588 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1244_
timestamp 1704896540
transform -1 0 5060 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _1245_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6716 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1246_
timestamp 1704896540
transform 1 0 4508 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1247_
timestamp 1704896540
transform 1 0 6072 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1248_
timestamp 1704896540
transform -1 0 5704 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1249_
timestamp 1704896540
transform 1 0 4508 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1250_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4048 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1251_
timestamp 1704896540
transform -1 0 4968 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1252_
timestamp 1704896540
transform -1 0 6348 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1253_
timestamp 1704896540
transform 1 0 5152 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1254_
timestamp 1704896540
transform -1 0 4600 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1255_
timestamp 1704896540
transform -1 0 4416 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1256_
timestamp 1704896540
transform 1 0 4600 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1257_
timestamp 1704896540
transform 1 0 4968 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1258_
timestamp 1704896540
transform 1 0 6900 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1259_
timestamp 1704896540
transform 1 0 6716 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1260_
timestamp 1704896540
transform -1 0 6900 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1261_
timestamp 1704896540
transform -1 0 3128 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1262_
timestamp 1704896540
transform -1 0 6440 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1263_
timestamp 1704896540
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1264_
timestamp 1704896540
transform -1 0 5520 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1265_
timestamp 1704896540
transform -1 0 7820 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1266_
timestamp 1704896540
transform -1 0 7544 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1267_
timestamp 1704896540
transform -1 0 4876 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1268_
timestamp 1704896540
transform 1 0 4324 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1269_
timestamp 1704896540
transform -1 0 3772 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1270_
timestamp 1704896540
transform -1 0 3496 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1271_
timestamp 1704896540
transform -1 0 3772 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1272_
timestamp 1704896540
transform -1 0 17756 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1273_
timestamp 1704896540
transform 1 0 17204 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1274_
timestamp 1704896540
transform 1 0 12972 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_2  _1275_
timestamp 1704896540
transform 1 0 12604 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1276_
timestamp 1704896540
transform 1 0 13064 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1277_
timestamp 1704896540
transform 1 0 11960 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1278_
timestamp 1704896540
transform 1 0 11868 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1279_
timestamp 1704896540
transform 1 0 12604 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1280_
timestamp 1704896540
transform 1 0 12880 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_2  _1281_
timestamp 1704896540
transform 1 0 12420 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1282_
timestamp 1704896540
transform 1 0 13064 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_2  _1283_
timestamp 1704896540
transform 1 0 11592 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1284_
timestamp 1704896540
transform -1 0 10028 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1285_
timestamp 1704896540
transform 1 0 10212 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1286_
timestamp 1704896540
transform 1 0 11040 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1287_
timestamp 1704896540
transform 1 0 12236 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1288_
timestamp 1704896540
transform 1 0 11316 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1289_
timestamp 1704896540
transform -1 0 12236 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _1290_
timestamp 1704896540
transform 1 0 10580 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1291_
timestamp 1704896540
transform 1 0 14720 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1292_
timestamp 1704896540
transform -1 0 16008 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1293_
timestamp 1704896540
transform 1 0 11868 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1294_
timestamp 1704896540
transform -1 0 15272 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1295_
timestamp 1704896540
transform 1 0 15272 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1296_
timestamp 1704896540
transform 1 0 15824 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1297_
timestamp 1704896540
transform -1 0 16560 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1298_
timestamp 1704896540
transform 1 0 12420 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _1299_
timestamp 1704896540
transform -1 0 12144 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1300_
timestamp 1704896540
transform 1 0 12420 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _1301_
timestamp 1704896540
transform 1 0 15364 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1302_
timestamp 1704896540
transform -1 0 16376 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1303_
timestamp 1704896540
transform 1 0 10948 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _1304_
timestamp 1704896540
transform -1 0 14260 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1305_
timestamp 1704896540
transform -1 0 14168 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1306_
timestamp 1704896540
transform 1 0 15548 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1307_
timestamp 1704896540
transform -1 0 16376 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1308_
timestamp 1704896540
transform -1 0 10580 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1309_
timestamp 1704896540
transform -1 0 13432 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1310_
timestamp 1704896540
transform -1 0 12880 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1311_
timestamp 1704896540
transform 1 0 14260 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1312_
timestamp 1704896540
transform 1 0 12788 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1313_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 13432 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1314_
timestamp 1704896540
transform -1 0 14352 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1315_
timestamp 1704896540
transform 1 0 13156 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1316_
timestamp 1704896540
transform -1 0 13800 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1317_
timestamp 1704896540
transform -1 0 14076 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1318_
timestamp 1704896540
transform -1 0 13432 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1319_
timestamp 1704896540
transform -1 0 11684 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1320_
timestamp 1704896540
transform -1 0 10856 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1321_
timestamp 1704896540
transform 1 0 10488 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1322_
timestamp 1704896540
transform 1 0 15272 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1323_
timestamp 1704896540
transform -1 0 16652 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1324_
timestamp 1704896540
transform 1 0 12788 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1325_
timestamp 1704896540
transform 1 0 13064 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1326_
timestamp 1704896540
transform -1 0 11868 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1327_
timestamp 1704896540
transform -1 0 11592 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1328_
timestamp 1704896540
transform -1 0 11224 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1329_
timestamp 1704896540
transform -1 0 10212 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1330_
timestamp 1704896540
transform 1 0 9660 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1331_
timestamp 1704896540
transform -1 0 18584 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1332_
timestamp 1704896540
transform 1 0 17388 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1333_
timestamp 1704896540
transform -1 0 16468 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_2  _1334_
timestamp 1704896540
transform 1 0 15456 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1335_
timestamp 1704896540
transform 1 0 16100 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1336_
timestamp 1704896540
transform 1 0 14444 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1337_
timestamp 1704896540
transform 1 0 17388 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1338_
timestamp 1704896540
transform 1 0 17756 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1339_
timestamp 1704896540
transform 1 0 16468 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_2  _1340_
timestamp 1704896540
transform 1 0 15272 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1341_
timestamp 1704896540
transform 1 0 16100 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_2  _1342_
timestamp 1704896540
transform 1 0 15272 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1343_
timestamp 1704896540
transform -1 0 18492 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1344_
timestamp 1704896540
transform 1 0 17664 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1345_
timestamp 1704896540
transform -1 0 18952 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1346_
timestamp 1704896540
transform 1 0 18124 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1347_
timestamp 1704896540
transform 1 0 19596 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1348_
timestamp 1704896540
transform 1 0 18952 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _1349_
timestamp 1704896540
transform 1 0 18676 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1350_
timestamp 1704896540
transform 1 0 22632 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1351_
timestamp 1704896540
transform -1 0 23736 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1352_
timestamp 1704896540
transform 1 0 19504 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1353_
timestamp 1704896540
transform -1 0 23276 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1354_
timestamp 1704896540
transform 1 0 23276 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1355_
timestamp 1704896540
transform 1 0 23828 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1356_
timestamp 1704896540
transform -1 0 23736 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1357_
timestamp 1704896540
transform 1 0 19596 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _1358_
timestamp 1704896540
transform 1 0 20056 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1359_
timestamp 1704896540
transform 1 0 20516 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _1360_
timestamp 1704896540
transform 1 0 22632 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1361_
timestamp 1704896540
transform -1 0 23828 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1362_
timestamp 1704896540
transform 1 0 18768 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _1363_
timestamp 1704896540
transform 1 0 21620 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1364_
timestamp 1704896540
transform -1 0 22448 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1365_
timestamp 1704896540
transform 1 0 24288 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1366_
timestamp 1704896540
transform 1 0 24748 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1367_
timestamp 1704896540
transform 1 0 17480 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1368_
timestamp 1704896540
transform -1 0 22356 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1369_
timestamp 1704896540
transform -1 0 20884 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1370_
timestamp 1704896540
transform 1 0 22356 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1371_
timestamp 1704896540
transform 1 0 20700 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1372_
timestamp 1704896540
transform 1 0 21344 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1373_
timestamp 1704896540
transform -1 0 22080 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1374_
timestamp 1704896540
transform 1 0 21528 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1375_
timestamp 1704896540
transform -1 0 22172 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1376_
timestamp 1704896540
transform 1 0 22172 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1377_
timestamp 1704896540
transform 1 0 23184 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1378_
timestamp 1704896540
transform 1 0 17940 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1379_
timestamp 1704896540
transform -1 0 19228 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1380_
timestamp 1704896540
transform 1 0 17940 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1381_
timestamp 1704896540
transform 1 0 23736 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1382_
timestamp 1704896540
transform -1 0 25300 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1383_
timestamp 1704896540
transform -1 0 21160 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1384_
timestamp 1704896540
transform -1 0 20884 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1385_
timestamp 1704896540
transform -1 0 20332 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1386_
timestamp 1704896540
transform -1 0 20056 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1387_
timestamp 1704896540
transform -1 0 19136 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1388_
timestamp 1704896540
transform -1 0 18860 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1389_
timestamp 1704896540
transform -1 0 18216 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_2  _1390_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11592 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1391_
timestamp 1704896540
transform 1 0 11868 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1392_
timestamp 1704896540
transform 1 0 12328 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_2  _1393_
timestamp 1704896540
transform 1 0 14904 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1394_
timestamp 1704896540
transform 1 0 11776 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1395_
timestamp 1704896540
transform 1 0 17112 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1396_
timestamp 1704896540
transform 1 0 16100 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1397_
timestamp 1704896540
transform -1 0 20792 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_2  _1398_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12604 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _1399_
timestamp 1704896540
transform 1 0 17112 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1400_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 19504 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1401_
timestamp 1704896540
transform -1 0 19320 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1402_
timestamp 1704896540
transform -1 0 20608 0 1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1403_
timestamp 1704896540
transform 1 0 19596 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1404_
timestamp 1704896540
transform -1 0 19688 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1405_
timestamp 1704896540
transform -1 0 19320 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1406_
timestamp 1704896540
transform 1 0 18400 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1407_
timestamp 1704896540
transform -1 0 18584 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1408_
timestamp 1704896540
transform -1 0 18032 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1409_
timestamp 1704896540
transform 1 0 17020 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1410_
timestamp 1704896540
transform -1 0 16744 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1411_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 16468 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_2  _1412_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 13892 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1413_
timestamp 1704896540
transform 1 0 12788 0 1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1414_
timestamp 1704896540
transform -1 0 11316 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _1415_
timestamp 1704896540
transform 1 0 13984 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1416_
timestamp 1704896540
transform -1 0 10212 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1417_
timestamp 1704896540
transform 1 0 9016 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1418_
timestamp 1704896540
transform -1 0 17388 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1419_
timestamp 1704896540
transform 1 0 8372 0 -1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1420_
timestamp 1704896540
transform 1 0 8832 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1421_
timestamp 1704896540
transform 1 0 18032 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1422_
timestamp 1704896540
transform 1 0 7820 0 1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1423_
timestamp 1704896540
transform 1 0 9292 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1424_
timestamp 1704896540
transform 1 0 15916 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1425_
timestamp 1704896540
transform -1 0 10580 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1426_
timestamp 1704896540
transform 1 0 9936 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1427_
timestamp 1704896540
transform 1 0 16744 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1428_
timestamp 1704896540
transform -1 0 10856 0 -1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1429_
timestamp 1704896540
transform -1 0 9936 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1430_
timestamp 1704896540
transform -1 0 13064 0 -1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1431_
timestamp 1704896540
transform 1 0 11868 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1432_
timestamp 1704896540
transform -1 0 12052 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1433_
timestamp 1704896540
transform -1 0 13984 0 1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1434_
timestamp 1704896540
transform 1 0 11776 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1435_
timestamp 1704896540
transform -1 0 14812 0 1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1436_
timestamp 1704896540
transform 1 0 12604 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_4  _1437_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 13432 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_1  _1438_
timestamp 1704896540
transform 1 0 12880 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1439_
timestamp 1704896540
transform -1 0 14444 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1440_
timestamp 1704896540
transform 1 0 12972 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1441_
timestamp 1704896540
transform -1 0 13616 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1442_
timestamp 1704896540
transform -1 0 12972 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1443_
timestamp 1704896540
transform 1 0 12236 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1444_
timestamp 1704896540
transform -1 0 14076 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1445_
timestamp 1704896540
transform 1 0 12604 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1446_
timestamp 1704896540
transform -1 0 13248 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1447_
timestamp 1704896540
transform 1 0 12420 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1448_
timestamp 1704896540
transform -1 0 13984 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1449_
timestamp 1704896540
transform -1 0 13524 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1450_
timestamp 1704896540
transform -1 0 17296 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1451_
timestamp 1704896540
transform -1 0 17940 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1452_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5704 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1453_
timestamp 1704896540
transform 1 0 17756 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1454_
timestamp 1704896540
transform 1 0 17940 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1455_
timestamp 1704896540
transform -1 0 18124 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1456_
timestamp 1704896540
transform 1 0 18584 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1457_
timestamp 1704896540
transform -1 0 20056 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1458_
timestamp 1704896540
transform -1 0 15456 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1459_
timestamp 1704896540
transform 1 0 8372 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1460_
timestamp 1704896540
transform 1 0 21712 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1461_
timestamp 1704896540
transform 1 0 21712 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1462_
timestamp 1704896540
transform -1 0 21712 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1463_
timestamp 1704896540
transform 1 0 20884 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1464_
timestamp 1704896540
transform -1 0 25576 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1465_
timestamp 1704896540
transform -1 0 25760 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1466_
timestamp 1704896540
transform 1 0 24288 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1467_
timestamp 1704896540
transform -1 0 20976 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _1468_
timestamp 1704896540
transform 1 0 24196 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _1469_
timestamp 1704896540
transform 1 0 24012 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1470_
timestamp 1704896540
transform -1 0 25484 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1471_
timestamp 1704896540
transform -1 0 25208 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1472_
timestamp 1704896540
transform -1 0 26220 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1473_
timestamp 1704896540
transform -1 0 25484 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1474_
timestamp 1704896540
transform 1 0 24380 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1475_
timestamp 1704896540
transform -1 0 25760 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1476_
timestamp 1704896540
transform 1 0 24012 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1477_
timestamp 1704896540
transform -1 0 24656 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1478_
timestamp 1704896540
transform 1 0 23184 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1479_
timestamp 1704896540
transform -1 0 23184 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1480_
timestamp 1704896540
transform -1 0 24288 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1481_
timestamp 1704896540
transform 1 0 23000 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_2  _1482_
timestamp 1704896540
transform 1 0 23000 0 -1 7072
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1483_
timestamp 1704896540
transform 1 0 21344 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1484_
timestamp 1704896540
transform -1 0 21712 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1485_
timestamp 1704896540
transform 1 0 22724 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1486_
timestamp 1704896540
transform -1 0 24288 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1487_
timestamp 1704896540
transform -1 0 24012 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1488_
timestamp 1704896540
transform -1 0 21712 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _1489_
timestamp 1704896540
transform -1 0 6348 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1490_
timestamp 1704896540
transform 1 0 21712 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1491_
timestamp 1704896540
transform -1 0 21804 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1492_
timestamp 1704896540
transform 1 0 19596 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1493_
timestamp 1704896540
transform -1 0 21068 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1494_
timestamp 1704896540
transform -1 0 21528 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1495_
timestamp 1704896540
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1496_
timestamp 1704896540
transform 1 0 20056 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1497_
timestamp 1704896540
transform 1 0 20516 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1498_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 19964 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1499_
timestamp 1704896540
transform -1 0 20056 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1500_
timestamp 1704896540
transform 1 0 20056 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1501_
timestamp 1704896540
transform 1 0 20148 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1502_
timestamp 1704896540
transform 1 0 19320 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_2  _1503_
timestamp 1704896540
transform 1 0 19412 0 1 7072
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1504_
timestamp 1704896540
transform -1 0 19136 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1505_
timestamp 1704896540
transform -1 0 18124 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1506_
timestamp 1704896540
transform -1 0 18952 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1507_
timestamp 1704896540
transform 1 0 19136 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1508_
timestamp 1704896540
transform -1 0 18952 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1509_
timestamp 1704896540
transform 1 0 18584 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1510_
timestamp 1704896540
transform 1 0 17664 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1511_
timestamp 1704896540
transform -1 0 18400 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1512_
timestamp 1704896540
transform 1 0 17480 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _1513_
timestamp 1704896540
transform 1 0 19320 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1514_
timestamp 1704896540
transform 1 0 11040 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1515_
timestamp 1704896540
transform -1 0 16744 0 -1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _1516_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 14352 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1517_
timestamp 1704896540
transform -1 0 13340 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1518_
timestamp 1704896540
transform 1 0 12972 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1519_
timestamp 1704896540
transform 1 0 13984 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1520_
timestamp 1704896540
transform 1 0 13524 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1521_
timestamp 1704896540
transform 1 0 12880 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1522_
timestamp 1704896540
transform -1 0 13800 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1523_
timestamp 1704896540
transform 1 0 10856 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1524_
timestamp 1704896540
transform 1 0 10212 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1525_
timestamp 1704896540
transform -1 0 11224 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1526_
timestamp 1704896540
transform 1 0 11040 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1527_
timestamp 1704896540
transform 1 0 10120 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1528_
timestamp 1704896540
transform 1 0 10580 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1529_
timestamp 1704896540
transform 1 0 12144 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1530_
timestamp 1704896540
transform 1 0 11408 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1531_
timestamp 1704896540
transform 1 0 1656 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1532_
timestamp 1704896540
transform 1 0 1656 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1533_
timestamp 1704896540
transform 1 0 1380 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1534_
timestamp 1704896540
transform 1 0 2668 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1535_
timestamp 1704896540
transform 1 0 2944 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1536_
timestamp 1704896540
transform 1 0 2300 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1537_
timestamp 1704896540
transform -1 0 3772 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1538_
timestamp 1704896540
transform 1 0 1932 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1539_
timestamp 1704896540
transform 1 0 1380 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1540_
timestamp 1704896540
transform -1 0 3680 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1541_
timestamp 1704896540
transform 1 0 3220 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1542_
timestamp 1704896540
transform -1 0 3036 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1543_
timestamp 1704896540
transform 1 0 2576 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1544_
timestamp 1704896540
transform -1 0 5336 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1545_
timestamp 1704896540
transform 1 0 8740 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1546_
timestamp 1704896540
transform 1 0 6808 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1547_
timestamp 1704896540
transform -1 0 4140 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1548_
timestamp 1704896540
transform 1 0 4140 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1549_
timestamp 1704896540
transform 1 0 4048 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1550_
timestamp 1704896540
transform 1 0 11040 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1551_
timestamp 1704896540
transform -1 0 11776 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1552_
timestamp 1704896540
transform 1 0 11500 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1553_
timestamp 1704896540
transform 1 0 11316 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1554_
timestamp 1704896540
transform 1 0 11684 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1555_
timestamp 1704896540
transform 1 0 10948 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1556_
timestamp 1704896540
transform 1 0 10212 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1557_
timestamp 1704896540
transform 1 0 10120 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1558_
timestamp 1704896540
transform 1 0 9568 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1559_
timestamp 1704896540
transform 1 0 9200 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1560_
timestamp 1704896540
transform 1 0 11224 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1561_
timestamp 1704896540
transform 1 0 11040 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1562_
timestamp 1704896540
transform -1 0 10396 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1563_
timestamp 1704896540
transform 1 0 15548 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1564_
timestamp 1704896540
transform 1 0 16100 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1565_
timestamp 1704896540
transform -1 0 9752 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1566_
timestamp 1704896540
transform -1 0 9752 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1567_
timestamp 1704896540
transform -1 0 7452 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1568_
timestamp 1704896540
transform 1 0 5336 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1569_
timestamp 1704896540
transform -1 0 8832 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1570_
timestamp 1704896540
transform -1 0 8004 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1571_
timestamp 1704896540
transform 1 0 8464 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1572_
timestamp 1704896540
transform -1 0 9108 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1573_
timestamp 1704896540
transform -1 0 8188 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1574_
timestamp 1704896540
transform 1 0 6716 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1575_
timestamp 1704896540
transform 1 0 6900 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1576_
timestamp 1704896540
transform 1 0 7636 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1577_
timestamp 1704896540
transform -1 0 6900 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1578_
timestamp 1704896540
transform 1 0 6256 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1579_
timestamp 1704896540
transform 1 0 7268 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1580_
timestamp 1704896540
transform 1 0 7268 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1581_
timestamp 1704896540
transform 1 0 8556 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1582_
timestamp 1704896540
transform 1 0 8556 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_4  _1583_
timestamp 1704896540
transform 1 0 11684 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_1  _1584_
timestamp 1704896540
transform -1 0 13432 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1585_
timestamp 1704896540
transform -1 0 8280 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1586_
timestamp 1704896540
transform 1 0 13708 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1587_
timestamp 1704896540
transform -1 0 15456 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1588_
timestamp 1704896540
transform 1 0 13892 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1589_
timestamp 1704896540
transform -1 0 14628 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1590_
timestamp 1704896540
transform 1 0 13616 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1591_
timestamp 1704896540
transform -1 0 15732 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1592_
timestamp 1704896540
transform 1 0 14720 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1593_
timestamp 1704896540
transform -1 0 14628 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1594_
timestamp 1704896540
transform 1 0 13800 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1595_
timestamp 1704896540
transform 1 0 14260 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1596_
timestamp 1704896540
transform 1 0 15364 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1597_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 14904 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1598_
timestamp 1704896540
transform 1 0 13524 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1599_
timestamp 1704896540
transform -1 0 7360 0 -1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1600_
timestamp 1704896540
transform 1 0 6164 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1601_
timestamp 1704896540
transform -1 0 7636 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1602_
timestamp 1704896540
transform -1 0 8188 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1603_
timestamp 1704896540
transform -1 0 6808 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1604_
timestamp 1704896540
transform 1 0 6808 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1605_
timestamp 1704896540
transform -1 0 7084 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1606_
timestamp 1704896540
transform -1 0 6532 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1607_
timestamp 1704896540
transform 1 0 7084 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1608_
timestamp 1704896540
transform 1 0 12512 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1609_
timestamp 1704896540
transform -1 0 12512 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1610_
timestamp 1704896540
transform -1 0 12144 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1611_
timestamp 1704896540
transform 1 0 11316 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1612_
timestamp 1704896540
transform -1 0 12512 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1613_
timestamp 1704896540
transform 1 0 11500 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1614_
timestamp 1704896540
transform -1 0 14996 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1615_
timestamp 1704896540
transform -1 0 13156 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1616_
timestamp 1704896540
transform 1 0 12144 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1617_
timestamp 1704896540
transform -1 0 13064 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1618_
timestamp 1704896540
transform 1 0 11500 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1619_
timestamp 1704896540
transform -1 0 13156 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1620_
timestamp 1704896540
transform 1 0 12144 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1621_
timestamp 1704896540
transform 1 0 21160 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1622_
timestamp 1704896540
transform 1 0 20148 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1623_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 20424 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1624_
timestamp 1704896540
transform -1 0 21160 0 1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1625_
timestamp 1704896540
transform -1 0 20516 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1626_
timestamp 1704896540
transform 1 0 20884 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1627_
timestamp 1704896540
transform -1 0 23368 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1628_
timestamp 1704896540
transform 1 0 22172 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1629_
timestamp 1704896540
transform -1 0 21528 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1630_
timestamp 1704896540
transform 1 0 21528 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_1  _1631_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 21804 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1632_
timestamp 1704896540
transform 1 0 20056 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1633_
timestamp 1704896540
transform -1 0 23092 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1634_
timestamp 1704896540
transform 1 0 20148 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _1635_
timestamp 1704896540
transform -1 0 21804 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1636_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 20332 0 1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1637_
timestamp 1704896540
transform 1 0 21804 0 -1 29920
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1638_
timestamp 1704896540
transform -1 0 21160 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1639_
timestamp 1704896540
transform 1 0 21252 0 1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1640_
timestamp 1704896540
transform -1 0 23920 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1641_
timestamp 1704896540
transform -1 0 22264 0 1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1642_
timestamp 1704896540
transform -1 0 23092 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1643_
timestamp 1704896540
transform -1 0 21712 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__o32ai_1  _1644_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 21252 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1645_
timestamp 1704896540
transform -1 0 23920 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1646_
timestamp 1704896540
transform 1 0 24288 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1647_
timestamp 1704896540
transform -1 0 26772 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1648_
timestamp 1704896540
transform -1 0 26956 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1649_
timestamp 1704896540
transform -1 0 22540 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1650_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 22080 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1651_
timestamp 1704896540
transform 1 0 21252 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1652_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 21344 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1653_
timestamp 1704896540
transform 1 0 21620 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1654_
timestamp 1704896540
transform -1 0 22724 0 -1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _1655_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 22448 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1656_
timestamp 1704896540
transform 1 0 21160 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1657_
timestamp 1704896540
transform -1 0 21344 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1658_
timestamp 1704896540
transform 1 0 5796 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _1659_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3128 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1660_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4784 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1661_
timestamp 1704896540
transform 1 0 5520 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_4  _1662_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7360 0 -1 29920
box -38 -48 1602 592
use sky130_fd_sc_hd__a21bo_1  _1663_
timestamp 1704896540
transform 1 0 21344 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1664_
timestamp 1704896540
transform -1 0 22724 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1665_
timestamp 1704896540
transform 1 0 20148 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1666_
timestamp 1704896540
transform -1 0 21068 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1667_
timestamp 1704896540
transform 1 0 22724 0 -1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1668_
timestamp 1704896540
transform 1 0 24564 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1669_
timestamp 1704896540
transform 1 0 6348 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1670_
timestamp 1704896540
transform 1 0 5888 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1671_
timestamp 1704896540
transform 1 0 24564 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1672_
timestamp 1704896540
transform 1 0 25392 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1673_
timestamp 1704896540
transform 1 0 22356 0 1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1674_
timestamp 1704896540
transform 1 0 23092 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1675_
timestamp 1704896540
transform -1 0 23552 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1676_
timestamp 1704896540
transform 1 0 22724 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1677_
timestamp 1704896540
transform 1 0 22264 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1678_
timestamp 1704896540
transform 1 0 23368 0 -1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1679_
timestamp 1704896540
transform 1 0 23552 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1680_
timestamp 1704896540
transform -1 0 24104 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1681_
timestamp 1704896540
transform -1 0 23644 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1682_
timestamp 1704896540
transform 1 0 23276 0 1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1683_
timestamp 1704896540
transform -1 0 24748 0 1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1684_
timestamp 1704896540
transform -1 0 24288 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1685_
timestamp 1704896540
transform -1 0 24288 0 1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1686_
timestamp 1704896540
transform -1 0 23276 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1687_
timestamp 1704896540
transform 1 0 24196 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1688_
timestamp 1704896540
transform -1 0 25392 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1689_
timestamp 1704896540
transform 1 0 24288 0 1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1690_
timestamp 1704896540
transform 1 0 23828 0 1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1691_
timestamp 1704896540
transform 1 0 24748 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1692_
timestamp 1704896540
transform -1 0 25852 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1693_
timestamp 1704896540
transform -1 0 24288 0 -1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1694_
timestamp 1704896540
transform -1 0 25116 0 -1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1695_
timestamp 1704896540
transform 1 0 24288 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1696_
timestamp 1704896540
transform -1 0 25300 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1697_
timestamp 1704896540
transform -1 0 24104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1698_
timestamp 1704896540
transform -1 0 23828 0 -1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1699_
timestamp 1704896540
transform -1 0 24288 0 1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1700_
timestamp 1704896540
transform -1 0 23368 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1701_
timestamp 1704896540
transform 1 0 23828 0 1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1702_
timestamp 1704896540
transform 1 0 23000 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1703_
timestamp 1704896540
transform 1 0 23368 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1704_
timestamp 1704896540
transform -1 0 24932 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1705_
timestamp 1704896540
transform 1 0 24840 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1706_
timestamp 1704896540
transform 1 0 24288 0 -1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1707_
timestamp 1704896540
transform -1 0 24840 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1708_
timestamp 1704896540
transform 1 0 25116 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1709_
timestamp 1704896540
transform 1 0 25116 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1710_
timestamp 1704896540
transform 1 0 25576 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1711_
timestamp 1704896540
transform 1 0 26036 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1712_
timestamp 1704896540
transform 1 0 25484 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1713_
timestamp 1704896540
transform -1 0 18492 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1714_
timestamp 1704896540
transform -1 0 16836 0 1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1715_
timestamp 1704896540
transform -1 0 17388 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1716_
timestamp 1704896540
transform 1 0 15640 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1717_
timestamp 1704896540
transform -1 0 15732 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1718_
timestamp 1704896540
transform -1 0 14996 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1719_
timestamp 1704896540
transform 1 0 14628 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1720_
timestamp 1704896540
transform -1 0 12144 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1721_
timestamp 1704896540
transform 1 0 10948 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1722_
timestamp 1704896540
transform 1 0 11224 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1723_
timestamp 1704896540
transform -1 0 9200 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1724_
timestamp 1704896540
transform 1 0 8464 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1725_
timestamp 1704896540
transform 1 0 8556 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1726_
timestamp 1704896540
transform -1 0 9660 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1727_
timestamp 1704896540
transform 1 0 9016 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1728_
timestamp 1704896540
transform -1 0 10764 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1729_
timestamp 1704896540
transform 1 0 9936 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1730_
timestamp 1704896540
transform -1 0 10948 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1731_
timestamp 1704896540
transform -1 0 10304 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1732_
timestamp 1704896540
transform -1 0 13248 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1733_
timestamp 1704896540
transform 1 0 11960 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1734_
timestamp 1704896540
transform -1 0 11868 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1735_
timestamp 1704896540
transform -1 0 13800 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1736_
timestamp 1704896540
transform 1 0 12696 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1737_
timestamp 1704896540
transform -1 0 14168 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1738_
timestamp 1704896540
transform -1 0 13248 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1739_
timestamp 1704896540
transform -1 0 18032 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1740_
timestamp 1704896540
transform 1 0 15364 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1741_
timestamp 1704896540
transform -1 0 14628 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _1742_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 16100 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1743_
timestamp 1704896540
transform -1 0 16008 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1744_
timestamp 1704896540
transform 1 0 15456 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1745_
timestamp 1704896540
transform 1 0 15456 0 1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1746_
timestamp 1704896540
transform 1 0 15456 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1747_
timestamp 1704896540
transform -1 0 7268 0 -1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1748_
timestamp 1704896540
transform 1 0 6348 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1749_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8740 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1750_
timestamp 1704896540
transform -1 0 8188 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1751_
timestamp 1704896540
transform -1 0 8372 0 -1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1752_
timestamp 1704896540
transform 1 0 6900 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1753_
timestamp 1704896540
transform 1 0 9016 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1754_
timestamp 1704896540
transform 1 0 8372 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1755_
timestamp 1704896540
transform -1 0 9016 0 1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1756_
timestamp 1704896540
transform 1 0 8648 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1757_
timestamp 1704896540
transform -1 0 10856 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1758_
timestamp 1704896540
transform -1 0 10580 0 -1 29920
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1759_
timestamp 1704896540
transform -1 0 10396 0 -1 31008
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1760_
timestamp 1704896540
transform -1 0 9476 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1761_
timestamp 1704896540
transform -1 0 10672 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1762_
timestamp 1704896540
transform 1 0 10028 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1763_
timestamp 1704896540
transform -1 0 10580 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1764_
timestamp 1704896540
transform 1 0 9384 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1765_
timestamp 1704896540
transform -1 0 11224 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1766_
timestamp 1704896540
transform 1 0 10948 0 1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1767_
timestamp 1704896540
transform 1 0 11224 0 -1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1768_
timestamp 1704896540
transform 1 0 11592 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1769_
timestamp 1704896540
transform -1 0 13432 0 1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1770_
timestamp 1704896540
transform 1 0 12972 0 1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1771_
timestamp 1704896540
transform 1 0 12880 0 -1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1772_
timestamp 1704896540
transform 1 0 13524 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1773_
timestamp 1704896540
transform 1 0 13524 0 1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1774_
timestamp 1704896540
transform 1 0 14444 0 -1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1775_
timestamp 1704896540
transform 1 0 13800 0 -1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1776_
timestamp 1704896540
transform -1 0 14536 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1777_
timestamp 1704896540
transform -1 0 15916 0 -1 29920
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1778_
timestamp 1704896540
transform 1 0 14352 0 -1 29920
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1779_
timestamp 1704896540
transform 1 0 14812 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1780_
timestamp 1704896540
transform 1 0 15364 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1781_
timestamp 1704896540
transform 1 0 14996 0 -1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1782_
timestamp 1704896540
transform 1 0 15272 0 1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1783_
timestamp 1704896540
transform -1 0 16744 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1784_
timestamp 1704896540
transform -1 0 16008 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1785_
timestamp 1704896540
transform 1 0 16560 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1786_
timestamp 1704896540
transform 1 0 16100 0 -1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1787_
timestamp 1704896540
transform 1 0 16100 0 1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1788_
timestamp 1704896540
transform -1 0 17112 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1789_
timestamp 1704896540
transform 1 0 16100 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1790_
timestamp 1704896540
transform 1 0 16836 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1791_
timestamp 1704896540
transform 1 0 17296 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1792_
timestamp 1704896540
transform -1 0 19044 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1793_
timestamp 1704896540
transform -1 0 18584 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1794_
timestamp 1704896540
transform 1 0 16008 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1795_
timestamp 1704896540
transform 1 0 17940 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1796_
timestamp 1704896540
transform -1 0 19136 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1797_
timestamp 1704896540
transform 1 0 16928 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1798_
timestamp 1704896540
transform -1 0 19412 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1799_
timestamp 1704896540
transform -1 0 19320 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1800_
timestamp 1704896540
transform -1 0 18400 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1801_
timestamp 1704896540
transform 1 0 16928 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1802_
timestamp 1704896540
transform -1 0 19872 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1803_
timestamp 1704896540
transform 1 0 18032 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1804_
timestamp 1704896540
transform -1 0 24472 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1805_
timestamp 1704896540
transform 1 0 21988 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1806_
timestamp 1704896540
transform 1 0 21252 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1807_
timestamp 1704896540
transform 1 0 20700 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1808_
timestamp 1704896540
transform 1 0 21068 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1809_
timestamp 1704896540
transform 1 0 21344 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1810_
timestamp 1704896540
transform -1 0 22724 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1811_
timestamp 1704896540
transform -1 0 24932 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1812_
timestamp 1704896540
transform -1 0 24380 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1813_
timestamp 1704896540
transform 1 0 20700 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1814_
timestamp 1704896540
transform -1 0 23276 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1815_
timestamp 1704896540
transform -1 0 23920 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1816_
timestamp 1704896540
transform -1 0 22724 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1817_
timestamp 1704896540
transform 1 0 22172 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1818_
timestamp 1704896540
transform 1 0 20516 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1819_
timestamp 1704896540
transform -1 0 22356 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1820_
timestamp 1704896540
transform -1 0 21804 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1821_
timestamp 1704896540
transform 1 0 21068 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1822_
timestamp 1704896540
transform -1 0 22632 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1823_
timestamp 1704896540
transform -1 0 22264 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1824_
timestamp 1704896540
transform 1 0 21252 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1825_
timestamp 1704896540
transform -1 0 22816 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1826_
timestamp 1704896540
transform -1 0 22540 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1827_
timestamp 1704896540
transform -1 0 23276 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1828_
timestamp 1704896540
transform -1 0 24104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1829_
timestamp 1704896540
transform -1 0 21988 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1830_
timestamp 1704896540
transform -1 0 21988 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1831_
timestamp 1704896540
transform 1 0 21344 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1832_
timestamp 1704896540
transform -1 0 22632 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1833_
timestamp 1704896540
transform -1 0 21804 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _1834_
timestamp 1704896540
transform 1 0 21988 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1835_
timestamp 1704896540
transform -1 0 20424 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1836_
timestamp 1704896540
transform -1 0 21528 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1837_
timestamp 1704896540
transform 1 0 19964 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1838_
timestamp 1704896540
transform 1 0 20792 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1839_
timestamp 1704896540
transform 1 0 22540 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1840_
timestamp 1704896540
transform 1 0 23276 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1841_
timestamp 1704896540
transform 1 0 24656 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1842_
timestamp 1704896540
transform 1 0 25392 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1843_
timestamp 1704896540
transform 1 0 21804 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1844_
timestamp 1704896540
transform -1 0 23184 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1845_
timestamp 1704896540
transform 1 0 22816 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1846_
timestamp 1704896540
transform -1 0 23460 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1847_
timestamp 1704896540
transform 1 0 22172 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1848_
timestamp 1704896540
transform -1 0 22632 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1849_
timestamp 1704896540
transform 1 0 22724 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1850_
timestamp 1704896540
transform -1 0 24104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1851_
timestamp 1704896540
transform 1 0 23460 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1852_
timestamp 1704896540
transform 1 0 23000 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1853_
timestamp 1704896540
transform 1 0 23276 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1854_
timestamp 1704896540
transform -1 0 24196 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1855_
timestamp 1704896540
transform -1 0 23000 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1856_
timestamp 1704896540
transform -1 0 22540 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1857_
timestamp 1704896540
transform 1 0 23000 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1858_
timestamp 1704896540
transform -1 0 24196 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1859_
timestamp 1704896540
transform 1 0 23184 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1860_
timestamp 1704896540
transform -1 0 22540 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1861_
timestamp 1704896540
transform -1 0 23184 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1862_
timestamp 1704896540
transform -1 0 24104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1863_
timestamp 1704896540
transform 1 0 24656 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1864_
timestamp 1704896540
transform 1 0 24380 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1865_
timestamp 1704896540
transform 1 0 25116 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1866_
timestamp 1704896540
transform -1 0 25852 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1867_
timestamp 1704896540
transform 1 0 25760 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1868_
timestamp 1704896540
transform -1 0 26312 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1869_
timestamp 1704896540
transform 1 0 25116 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1870_
timestamp 1704896540
transform -1 0 26680 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1871_
timestamp 1704896540
transform -1 0 24932 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1872_
timestamp 1704896540
transform 1 0 25024 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1873_
timestamp 1704896540
transform 1 0 24932 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1874_
timestamp 1704896540
transform -1 0 26128 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1875_
timestamp 1704896540
transform 1 0 24564 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1876_
timestamp 1704896540
transform -1 0 25024 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1877_
timestamp 1704896540
transform 1 0 23828 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1878_
timestamp 1704896540
transform -1 0 24472 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _1879_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 22540 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__a21boi_1  _1880_
timestamp 1704896540
transform 1 0 22724 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1881_
timestamp 1704896540
transform -1 0 11224 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1882_
timestamp 1704896540
transform -1 0 11592 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1883_
timestamp 1704896540
transform -1 0 11408 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1884_
timestamp 1704896540
transform 1 0 10120 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1885_
timestamp 1704896540
transform 1 0 9568 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1886_
timestamp 1704896540
transform -1 0 10488 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1887_
timestamp 1704896540
transform 1 0 8740 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1888_
timestamp 1704896540
transform 1 0 9384 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1889_
timestamp 1704896540
transform -1 0 10948 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1890_
timestamp 1704896540
transform -1 0 10488 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1891_
timestamp 1704896540
transform 1 0 9016 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1892_
timestamp 1704896540
transform 1 0 10948 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1893_
timestamp 1704896540
transform -1 0 11776 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1894_
timestamp 1704896540
transform 1 0 4692 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1895_
timestamp 1704896540
transform 1 0 5060 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1896_
timestamp 1704896540
transform 1 0 15180 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1897_
timestamp 1704896540
transform 1 0 15456 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1898_
timestamp 1704896540
transform 1 0 14076 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1899_
timestamp 1704896540
transform 1 0 14444 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1900_
timestamp 1704896540
transform -1 0 13432 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1901_
timestamp 1704896540
transform 1 0 14904 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1902_
timestamp 1704896540
transform 1 0 13616 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1903_
timestamp 1704896540
transform -1 0 13984 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1904_
timestamp 1704896540
transform 1 0 14996 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1905_
timestamp 1704896540
transform -1 0 14904 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1906_
timestamp 1704896540
transform 1 0 14536 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1907_
timestamp 1704896540
transform 1 0 14720 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1908_
timestamp 1704896540
transform 1 0 15548 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1909_
timestamp 1704896540
transform 1 0 15364 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1910_
timestamp 1704896540
transform -1 0 16744 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1911_
timestamp 1704896540
transform 1 0 16192 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1912_
timestamp 1704896540
transform 1 0 15548 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1913_
timestamp 1704896540
transform 1 0 14996 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1914_
timestamp 1704896540
transform -1 0 15456 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1915_
timestamp 1704896540
transform -1 0 14260 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1916_
timestamp 1704896540
transform -1 0 16100 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1917_
timestamp 1704896540
transform 1 0 16008 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1918_
timestamp 1704896540
transform 1 0 15364 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1919_
timestamp 1704896540
transform -1 0 16744 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1920_
timestamp 1704896540
transform 1 0 15732 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1921_
timestamp 1704896540
transform 1 0 16100 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1922_
timestamp 1704896540
transform 1 0 16560 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1923_
timestamp 1704896540
transform -1 0 17296 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1924_
timestamp 1704896540
transform 1 0 15180 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1925_
timestamp 1704896540
transform 1 0 17848 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1926_
timestamp 1704896540
transform -1 0 18584 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1927_
timestamp 1704896540
transform 1 0 16836 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1928_
timestamp 1704896540
transform 1 0 21252 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1929_
timestamp 1704896540
transform 1 0 22264 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1930_
timestamp 1704896540
transform -1 0 24932 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _1931_
timestamp 1704896540
transform 1 0 20608 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1932_
timestamp 1704896540
transform 1 0 23460 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1933_
timestamp 1704896540
transform 1 0 21620 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1934_
timestamp 1704896540
transform 1 0 21712 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1935_
timestamp 1704896540
transform 1 0 22816 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1936_
timestamp 1704896540
transform 1 0 23184 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1937_
timestamp 1704896540
transform -1 0 25024 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1938_
timestamp 1704896540
transform -1 0 23000 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1939_
timestamp 1704896540
transform -1 0 23092 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1940_
timestamp 1704896540
transform -1 0 23644 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1941_
timestamp 1704896540
transform 1 0 22080 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1942_
timestamp 1704896540
transform -1 0 23736 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1943_
timestamp 1704896540
transform -1 0 23552 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1944_
timestamp 1704896540
transform 1 0 24380 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1945_
timestamp 1704896540
transform -1 0 24840 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1946_
timestamp 1704896540
transform 1 0 26404 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1947_
timestamp 1704896540
transform 1 0 25576 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1948_
timestamp 1704896540
transform 1 0 25760 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1949_
timestamp 1704896540
transform 1 0 25576 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1950_
timestamp 1704896540
transform 1 0 21896 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1951_
timestamp 1704896540
transform -1 0 25576 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1952_
timestamp 1704896540
transform -1 0 26220 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1953_
timestamp 1704896540
transform -1 0 25668 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1954_
timestamp 1704896540
transform 1 0 21528 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1955_
timestamp 1704896540
transform 1 0 25300 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1956_
timestamp 1704896540
transform 1 0 25116 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1957_
timestamp 1704896540
transform 1 0 26404 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1958_
timestamp 1704896540
transform 1 0 24932 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1959_
timestamp 1704896540
transform 1 0 26404 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1960_
timestamp 1704896540
transform -1 0 24288 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1961_
timestamp 1704896540
transform -1 0 23644 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1962_
timestamp 1704896540
transform 1 0 23000 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1963_
timestamp 1704896540
transform -1 0 24196 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1964_
timestamp 1704896540
transform -1 0 23736 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1965_
timestamp 1704896540
transform 1 0 22724 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1966_
timestamp 1704896540
transform -1 0 26220 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1967_
timestamp 1704896540
transform -1 0 25116 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1968_
timestamp 1704896540
transform -1 0 25484 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1969_
timestamp 1704896540
transform -1 0 23736 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1970_
timestamp 1704896540
transform -1 0 21896 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1971_
timestamp 1704896540
transform 1 0 21896 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _1972_
timestamp 1704896540
transform 1 0 21528 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__o2111a_1  _1973_
timestamp 1704896540
transform 1 0 22172 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1974_
timestamp 1704896540
transform 1 0 16928 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1975_
timestamp 1704896540
transform 1 0 17572 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1976_
timestamp 1704896540
transform -1 0 20884 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1977_
timestamp 1704896540
transform -1 0 18032 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1978_
timestamp 1704896540
transform 1 0 18400 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1979_
timestamp 1704896540
transform -1 0 21620 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1980_
timestamp 1704896540
transform -1 0 17572 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1981_
timestamp 1704896540
transform -1 0 21896 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1982_
timestamp 1704896540
transform -1 0 18032 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1983_
timestamp 1704896540
transform -1 0 20056 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1984_
timestamp 1704896540
transform -1 0 7452 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1985_
timestamp 1704896540
transform -1 0 7820 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _1986_
timestamp 1704896540
transform 1 0 6440 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1987_
timestamp 1704896540
transform -1 0 11316 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1988_
timestamp 1704896540
transform 1 0 9292 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1989_
timestamp 1704896540
transform -1 0 9016 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1990_
timestamp 1704896540
transform 1 0 8648 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1991_
timestamp 1704896540
transform 1 0 9016 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1992_
timestamp 1704896540
transform -1 0 8556 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1993_
timestamp 1704896540
transform -1 0 15456 0 1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1994_
timestamp 1704896540
transform -1 0 17112 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1995_
timestamp 1704896540
transform 1 0 14352 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1996_
timestamp 1704896540
transform 1 0 13892 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1997_
timestamp 1704896540
transform -1 0 15548 0 1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1998_
timestamp 1704896540
transform 1 0 14628 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1999_
timestamp 1704896540
transform 1 0 14812 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2000_
timestamp 1704896540
transform -1 0 17848 0 1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _2001_
timestamp 1704896540
transform 1 0 16100 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2002_
timestamp 1704896540
transform -1 0 15916 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2003_
timestamp 1704896540
transform 1 0 15548 0 -1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _2004_
timestamp 1704896540
transform 1 0 16100 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2005_
timestamp 1704896540
transform 1 0 15272 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2006_
timestamp 1704896540
transform -1 0 6440 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _2007_
timestamp 1704896540
transform -1 0 6348 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _2008_
timestamp 1704896540
transform 1 0 4968 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _2009_
timestamp 1704896540
transform 1 0 4416 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_1  _2010_
timestamp 1704896540
transform 1 0 5152 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2011_
timestamp 1704896540
transform 1 0 6440 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2012_
timestamp 1704896540
transform 1 0 4600 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2013_
timestamp 1704896540
transform 1 0 4876 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _2014_
timestamp 1704896540
transform 1 0 4876 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2015_
timestamp 1704896540
transform 1 0 5428 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2016_
timestamp 1704896540
transform -1 0 6072 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2017_
timestamp 1704896540
transform -1 0 6348 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2018_
timestamp 1704896540
transform -1 0 3496 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2019_
timestamp 1704896540
transform 1 0 3312 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2020_
timestamp 1704896540
transform 1 0 3588 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _2021_
timestamp 1704896540
transform 1 0 3680 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _2022_
timestamp 1704896540
transform 1 0 3588 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2023_
timestamp 1704896540
transform -1 0 3312 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2024_
timestamp 1704896540
transform 1 0 3036 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2025_
timestamp 1704896540
transform -1 0 5520 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2026_
timestamp 1704896540
transform -1 0 5152 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _2027_
timestamp 1704896540
transform 1 0 3956 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2028_
timestamp 1704896540
transform 1 0 4324 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _2029_
timestamp 1704896540
transform -1 0 5336 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__o211ai_1  _2030_
timestamp 1704896540
transform 1 0 4600 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _2031_
timestamp 1704896540
transform 1 0 4048 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _2032_
timestamp 1704896540
transform -1 0 6164 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2033_
timestamp 1704896540
transform 1 0 5520 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _2034_
timestamp 1704896540
transform 1 0 5796 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _2035_
timestamp 1704896540
transform -1 0 6348 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _2036_
timestamp 1704896540
transform 1 0 4692 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _2037_
timestamp 1704896540
transform 1 0 3956 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _2038_
timestamp 1704896540
transform 1 0 5060 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2039_
timestamp 1704896540
transform 1 0 5152 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _2040_
timestamp 1704896540
transform -1 0 5060 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2041_
timestamp 1704896540
transform 1 0 3220 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _2042_
timestamp 1704896540
transform -1 0 4876 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _2043_
timestamp 1704896540
transform 1 0 2484 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _2044_
timestamp 1704896540
transform 1 0 3220 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__o2111ai_1  _2045_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3956 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2046_
timestamp 1704896540
transform 1 0 3404 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2047_
timestamp 1704896540
transform 1 0 4324 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2048_
timestamp 1704896540
transform -1 0 2944 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2049_
timestamp 1704896540
transform 1 0 2852 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2050_
timestamp 1704896540
transform 1 0 3036 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2051_
timestamp 1704896540
transform 1 0 4968 0 1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _2052_
timestamp 1704896540
transform 1 0 4692 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2053_
timestamp 1704896540
transform -1 0 4324 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2054_
timestamp 1704896540
transform -1 0 4876 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2055_
timestamp 1704896540
transform 1 0 4324 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2056_
timestamp 1704896540
transform 1 0 4692 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__nor4b_1  _2057_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4876 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2058_
timestamp 1704896540
transform 1 0 4876 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2059_
timestamp 1704896540
transform -1 0 5060 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _2060_
timestamp 1704896540
transform -1 0 5980 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _2061_
timestamp 1704896540
transform -1 0 6440 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2062_
timestamp 1704896540
transform -1 0 5520 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _2063_
timestamp 1704896540
transform -1 0 5428 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _2064_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4784 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2065_
timestamp 1704896540
transform 1 0 1748 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _2066_
timestamp 1704896540
transform -1 0 6440 0 -1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2067_
timestamp 1704896540
transform -1 0 4048 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _2068_
timestamp 1704896540
transform -1 0 6440 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2069_
timestamp 1704896540
transform 1 0 4968 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2070_
timestamp 1704896540
transform -1 0 4876 0 -1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2071_
timestamp 1704896540
transform -1 0 4416 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _2072_
timestamp 1704896540
transform 1 0 5060 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2073_
timestamp 1704896540
transform 1 0 4508 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _2074_
timestamp 1704896540
transform 1 0 3588 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _2075_
timestamp 1704896540
transform 1 0 3864 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2076_
timestamp 1704896540
transform -1 0 3404 0 -1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2077_
timestamp 1704896540
transform -1 0 3036 0 1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _2078_
timestamp 1704896540
transform 1 0 2300 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _2079_
timestamp 1704896540
transform -1 0 3496 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2080_
timestamp 1704896540
transform -1 0 2760 0 -1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2081_
timestamp 1704896540
transform -1 0 3220 0 -1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _2082_
timestamp 1704896540
transform -1 0 2944 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _2083_
timestamp 1704896540
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2084_
timestamp 1704896540
transform 1 0 2576 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2085_
timestamp 1704896540
transform 1 0 2300 0 -1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _2086_
timestamp 1704896540
transform 1 0 2392 0 1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2087_
timestamp 1704896540
transform -1 0 3128 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2088_
timestamp 1704896540
transform -1 0 2484 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2089_
timestamp 1704896540
transform -1 0 2024 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2090_
timestamp 1704896540
transform -1 0 2576 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2091_
timestamp 1704896540
transform -1 0 2116 0 1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2092_
timestamp 1704896540
transform 1 0 1012 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2093_
timestamp 1704896540
transform -1 0 3036 0 1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2094_
timestamp 1704896540
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _2095_
timestamp 1704896540
transform -1 0 2024 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _2096_
timestamp 1704896540
transform -1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2097_
timestamp 1704896540
transform -1 0 2944 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2098_
timestamp 1704896540
transform -1 0 2024 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _2099_
timestamp 1704896540
transform -1 0 1656 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2100_
timestamp 1704896540
transform 1 0 920 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2101_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9844 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2102_
timestamp 1704896540
transform 1 0 19320 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2103_
timestamp 1704896540
transform 1 0 19688 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2104_
timestamp 1704896540
transform 1 0 18676 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2105_
timestamp 1704896540
transform 1 0 16744 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2106_
timestamp 1704896540
transform 1 0 8464 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2107_
timestamp 1704896540
transform 1 0 8372 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2108_
timestamp 1704896540
transform 1 0 8648 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2109_
timestamp 1704896540
transform 1 0 9476 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2110_
timestamp 1704896540
transform 1 0 10120 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2111_
timestamp 1704896540
transform 1 0 11132 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2112_
timestamp 1704896540
transform 1 0 11316 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2113_
timestamp 1704896540
transform 1 0 11960 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2114_
timestamp 1704896540
transform 1 0 13524 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2115_
timestamp 1704896540
transform 1 0 11500 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2116_
timestamp 1704896540
transform 1 0 12144 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2117_
timestamp 1704896540
transform 1 0 11868 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2118_
timestamp 1704896540
transform 1 0 13524 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2119_
timestamp 1704896540
transform 1 0 18860 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2120_
timestamp 1704896540
transform 1 0 17296 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2121_
timestamp 1704896540
transform 1 0 19228 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2122_
timestamp 1704896540
transform 1 0 19228 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2123_
timestamp 1704896540
transform 1 0 20240 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2124_
timestamp 1704896540
transform 1 0 25024 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2125_
timestamp 1704896540
transform 1 0 24656 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2126_
timestamp 1704896540
transform 1 0 21712 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2127_
timestamp 1704896540
transform 1 0 21252 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2128_
timestamp 1704896540
transform -1 0 20608 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2129_
timestamp 1704896540
transform 1 0 18124 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2130_
timestamp 1704896540
transform 1 0 17020 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2131_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2392 0 -1 29920
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2132_
timestamp 1704896540
transform 1 0 13340 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2133_
timestamp 1704896540
transform 1 0 13340 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2134_
timestamp 1704896540
transform -1 0 11592 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2135_
timestamp 1704896540
transform 1 0 9936 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2136_
timestamp 1704896540
transform 1 0 11316 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2137_
timestamp 1704896540
transform 1 0 1932 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2138_
timestamp 1704896540
transform 1 0 828 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2139_
timestamp 1704896540
transform -1 0 4692 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2140_
timestamp 1704896540
transform 1 0 828 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2141_
timestamp 1704896540
transform 1 0 2300 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2142_
timestamp 1704896540
transform 1 0 4140 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2143_
timestamp 1704896540
transform 1 0 3680 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2144_
timestamp 1704896540
transform -1 0 10856 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2145_
timestamp 1704896540
transform 1 0 10212 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2146_
timestamp 1704896540
transform 1 0 8740 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2147_
timestamp 1704896540
transform 1 0 10396 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2148_
timestamp 1704896540
transform 1 0 5612 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2149_
timestamp 1704896540
transform -1 0 8464 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2150_
timestamp 1704896540
transform -1 0 9844 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2151_
timestamp 1704896540
transform 1 0 5888 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2152_
timestamp 1704896540
transform -1 0 8280 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2153_
timestamp 1704896540
transform 1 0 6072 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2154_
timestamp 1704896540
transform -1 0 7912 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2155_
timestamp 1704896540
transform -1 0 9384 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2156_
timestamp 1704896540
transform 1 0 13524 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2157_
timestamp 1704896540
transform 1 0 13156 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2158_
timestamp 1704896540
transform 1 0 14260 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2159_
timestamp 1704896540
transform 1 0 13524 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2160_
timestamp 1704896540
transform 1 0 14720 0 1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2161_
timestamp 1704896540
transform 1 0 6624 0 -1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2162_
timestamp 1704896540
transform -1 0 7820 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2163_
timestamp 1704896540
transform 1 0 7452 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2164_
timestamp 1704896540
transform -1 0 7176 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2165_
timestamp 1704896540
transform -1 0 9200 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2166_
timestamp 1704896540
transform 1 0 5428 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2167_
timestamp 1704896540
transform 1 0 5520 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2168_
timestamp 1704896540
transform -1 0 8924 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2169_
timestamp 1704896540
transform 1 0 10948 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2170_
timestamp 1704896540
transform 1 0 11040 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2171_
timestamp 1704896540
transform 1 0 11776 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2172_
timestamp 1704896540
transform 1 0 11132 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2173_
timestamp 1704896540
transform 1 0 12052 0 -1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2174_
timestamp 1704896540
transform -1 0 21160 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2175_
timestamp 1704896540
transform 1 0 25484 0 1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2176_
timestamp 1704896540
transform 1 0 22264 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2177_
timestamp 1704896540
transform -1 0 25576 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2178_
timestamp 1704896540
transform 1 0 24012 0 1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2179_
timestamp 1704896540
transform -1 0 26312 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2180_
timestamp 1704896540
transform 1 0 25576 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2181_
timestamp 1704896540
transform -1 0 26404 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2182_
timestamp 1704896540
transform -1 0 23736 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2183_
timestamp 1704896540
transform 1 0 22264 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2184_
timestamp 1704896540
transform -1 0 25484 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2185_
timestamp 1704896540
transform 1 0 25668 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2186_
timestamp 1704896540
transform 1 0 25484 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2187_
timestamp 1704896540
transform 1 0 15180 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2188_
timestamp 1704896540
transform 1 0 6624 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2189_
timestamp 1704896540
transform 1 0 6440 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2190_
timestamp 1704896540
transform 1 0 8004 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2191_
timestamp 1704896540
transform 1 0 9476 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2192_
timestamp 1704896540
transform 1 0 8924 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2193_
timestamp 1704896540
transform 1 0 11316 0 1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2194_
timestamp 1704896540
transform 1 0 12696 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2195_
timestamp 1704896540
transform -1 0 15456 0 1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2196_
timestamp 1704896540
transform -1 0 15364 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2197_
timestamp 1704896540
transform -1 0 17480 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2198_
timestamp 1704896540
transform 1 0 16744 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2199_
timestamp 1704896540
transform 1 0 16284 0 1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2200_
timestamp 1704896540
transform 1 0 18676 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2201_
timestamp 1704896540
transform -1 0 17848 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2202_
timestamp 1704896540
transform 1 0 16376 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2203_
timestamp 1704896540
transform 1 0 18676 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2204_
timestamp 1704896540
transform 1 0 16468 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2205_
timestamp 1704896540
transform -1 0 19044 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2206_
timestamp 1704896540
transform -1 0 20792 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2207_
timestamp 1704896540
transform 1 0 25300 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2208_
timestamp 1704896540
transform -1 0 24748 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2209_
timestamp 1704896540
transform -1 0 25300 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2210_
timestamp 1704896540
transform -1 0 25668 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2211_
timestamp 1704896540
transform -1 0 25668 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2212_
timestamp 1704896540
transform -1 0 24288 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2213_
timestamp 1704896540
transform -1 0 27048 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2214_
timestamp 1704896540
transform -1 0 27140 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2215_
timestamp 1704896540
transform 1 0 25668 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2216_
timestamp 1704896540
transform 1 0 25024 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2217_
timestamp 1704896540
transform 1 0 22264 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2218_
timestamp 1704896540
transform 1 0 22724 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2219_
timestamp 1704896540
transform 1 0 9384 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2220_
timestamp 1704896540
transform -1 0 11040 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2221_
timestamp 1704896540
transform 1 0 7912 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2222_
timestamp 1704896540
transform -1 0 11132 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2223_
timestamp 1704896540
transform -1 0 9568 0 -1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2224_
timestamp 1704896540
transform 1 0 4784 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2225_
timestamp 1704896540
transform -1 0 17388 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2226_
timestamp 1704896540
transform 1 0 14260 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2227_
timestamp 1704896540
transform -1 0 17572 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2228_
timestamp 1704896540
transform -1 0 17756 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2229_
timestamp 1704896540
transform 1 0 13708 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2230_
timestamp 1704896540
transform 1 0 15640 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2231_
timestamp 1704896540
transform -1 0 22080 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2232_
timestamp 1704896540
transform -1 0 25484 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2233_
timestamp 1704896540
transform 1 0 22540 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2234_
timestamp 1704896540
transform 1 0 20976 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2235_
timestamp 1704896540
transform -1 0 24104 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2236_
timestamp 1704896540
transform -1 0 25300 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2237_
timestamp 1704896540
transform 1 0 25576 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2238_
timestamp 1704896540
transform 1 0 25668 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2239_
timestamp 1704896540
transform 1 0 25484 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2240_
timestamp 1704896540
transform 1 0 25668 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2241_
timestamp 1704896540
transform 1 0 25668 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2242_
timestamp 1704896540
transform 1 0 25668 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2243_
timestamp 1704896540
transform 1 0 25484 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2244_
timestamp 1704896540
transform 1 0 23644 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2245_
timestamp 1704896540
transform -1 0 25300 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2246_
timestamp 1704896540
transform 1 0 21804 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2247_
timestamp 1704896540
transform 1 0 20700 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2248_
timestamp 1704896540
transform 1 0 18768 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2249_
timestamp 1704896540
transform 1 0 17112 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2250_
timestamp 1704896540
transform 1 0 19044 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2251_
timestamp 1704896540
transform 1 0 19136 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2252_
timestamp 1704896540
transform 1 0 17296 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2253_
timestamp 1704896540
transform 1 0 19136 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2254_
timestamp 1704896540
transform 1 0 17572 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2255_
timestamp 1704896540
transform 1 0 18952 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2256_
timestamp 1704896540
transform 1 0 8372 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2257_
timestamp 1704896540
transform 1 0 13524 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2258_
timestamp 1704896540
transform 1 0 14168 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2259_
timestamp 1704896540
transform 1 0 15916 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2260_
timestamp 1704896540
transform 1 0 15180 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2261_
timestamp 1704896540
transform 1 0 3496 0 1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2262_
timestamp 1704896540
transform 1 0 4784 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2263_
timestamp 1704896540
transform 1 0 3496 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2264_
timestamp 1704896540
transform -1 0 3956 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2265_
timestamp 1704896540
transform 1 0 828 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2266_
timestamp 1704896540
transform 1 0 2760 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2267_
timestamp 1704896540
transform 1 0 828 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2268_
timestamp 1704896540
transform 1 0 828 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2269_
timestamp 1704896540
transform 1 0 828 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2270_
timestamp 1704896540
transform 1 0 3220 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2271_
timestamp 1704896540
transform 1 0 828 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2272_
timestamp 1704896540
transform -1 0 3956 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2273_
timestamp 1704896540
transform 1 0 828 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2274_
timestamp 1704896540
transform 1 0 828 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2275_
timestamp 1704896540
transform -1 0 4692 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2276_
timestamp 1704896540
transform 1 0 2668 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2277_
timestamp 1704896540
transform 1 0 3588 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2278_
timestamp 1704896540
transform 1 0 6256 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2279_
timestamp 1704896540
transform 1 0 6440 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2280_
timestamp 1704896540
transform 1 0 5796 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2281_
timestamp 1704896540
transform 1 0 4232 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2282_
timestamp 1704896540
transform -1 0 7360 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dlxtn_2  _2283_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8096 0 -1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2283__61 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8648 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2284__62
timestamp 1704896540
transform -1 0 8188 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2284_
timestamp 1704896540
transform 1 0 7912 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2285__63
timestamp 1704896540
transform -1 0 7728 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2285_
timestamp 1704896540
transform 1 0 6716 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_2  _2286_
timestamp 1704896540
transform 1 0 6716 0 1 544
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2286__64
timestamp 1704896540
transform 1 0 6440 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2287_
timestamp 1704896540
transform 1 0 6256 0 1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2287__65
timestamp 1704896540
transform -1 0 7268 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2288__66
timestamp 1704896540
transform -1 0 6348 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2288_
timestamp 1704896540
transform 1 0 5060 0 1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_2  _2289_
timestamp 1704896540
transform -1 0 6992 0 -1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2289__67
timestamp 1704896540
transform 1 0 5796 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2290_
timestamp 1704896540
transform 1 0 4508 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2290__68
timestamp 1704896540
transform -1 0 5704 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2291__69
timestamp 1704896540
transform 1 0 4048 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2291_
timestamp 1704896540
transform 1 0 4232 0 1 544
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_2  _2292_
timestamp 1704896540
transform 1 0 3312 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2292__70
timestamp 1704896540
transform -1 0 3680 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2293__71
timestamp 1704896540
transform -1 0 3956 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2293_
timestamp 1704896540
transform -1 0 3312 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2294__72
timestamp 1704896540
transform 1 0 2024 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2294_
timestamp 1704896540
transform 1 0 2300 0 -1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_2  _2295_
timestamp 1704896540
transform 1 0 1932 0 1 544
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2295__73
timestamp 1704896540
transform -1 0 2392 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2296__74
timestamp 1704896540
transform -1 0 1656 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2296_
timestamp 1704896540
transform 1 0 920 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2297__75
timestamp 1704896540
transform -1 0 1288 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2297_
timestamp 1704896540
transform 1 0 920 0 1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_1  _2298_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5980 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2298__76
timestamp 1704896540
transform -1 0 6624 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2299__77
timestamp 1704896540
transform -1 0 8740 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _2299_
timestamp 1704896540
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _2300_
timestamp 1704896540
transform 1 0 4600 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2300__78
timestamp 1704896540
transform -1 0 5152 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2301__79
timestamp 1704896540
transform 1 0 3864 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _2301_
timestamp 1704896540
transform 1 0 4140 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _2302_
timestamp 1704896540
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2302__80
timestamp 1704896540
transform 1 0 2484 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2303__81
timestamp 1704896540
transform -1 0 1472 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _2303_
timestamp 1704896540
transform 1 0 1104 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2304__82
timestamp 1704896540
transform 1 0 1288 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _2304_
timestamp 1704896540
transform 1 0 1564 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2305__83
timestamp 1704896540
transform 1 0 4140 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _2305_
timestamp 1704896540
transform -1 0 4600 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2306__38
timestamp 1704896540
transform 1 0 16652 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2306_
timestamp 1704896540
transform 1 0 17296 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_2  _2307_
timestamp 1704896540
transform 1 0 16192 0 1 544
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2307__39
timestamp 1704896540
transform -1 0 16652 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2308__40
timestamp 1704896540
transform 1 0 15732 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2308_
timestamp 1704896540
transform 1 0 16100 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2309__41
timestamp 1704896540
transform -1 0 15548 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2309_
timestamp 1704896540
transform 1 0 15180 0 1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_2  _2310_
timestamp 1704896540
transform 1 0 14536 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2310__42
timestamp 1704896540
transform -1 0 14812 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2311__43
timestamp 1704896540
transform -1 0 14352 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2311_
timestamp 1704896540
transform 1 0 13984 0 1 544
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_2  _2312_
timestamp 1704896540
transform 1 0 13340 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2312__44
timestamp 1704896540
transform -1 0 13892 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2313_
timestamp 1704896540
transform -1 0 13340 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2313__45
timestamp 1704896540
transform -1 0 13800 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2314__46
timestamp 1704896540
transform -1 0 12604 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2314_
timestamp 1704896540
transform 1 0 12236 0 1 544
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2315__47
timestamp 1704896540
transform 1 0 11316 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2315_
timestamp 1704896540
transform 1 0 11592 0 1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2316__48
timestamp 1704896540
transform -1 0 11316 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2316_
timestamp 1704896540
transform 1 0 10948 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_2  _2317_
timestamp 1704896540
transform 1 0 10948 0 1 544
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2317__49
timestamp 1704896540
transform 1 0 10672 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2318__50
timestamp 1704896540
transform 1 0 9384 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2318_
timestamp 1704896540
transform 1 0 9660 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2319__51
timestamp 1704896540
transform 1 0 9108 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2319_
timestamp 1704896540
transform 1 0 9384 0 1 544
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2320__52
timestamp 1704896540
transform -1 0 9292 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2320_
timestamp 1704896540
transform 1 0 9016 0 1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_1  _2321_
timestamp 1704896540
transform 1 0 12328 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2321__53
timestamp 1704896540
transform -1 0 12696 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _2322_
timestamp 1704896540
transform 1 0 16284 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2322__54
timestamp 1704896540
transform -1 0 16652 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2323__55
timestamp 1704896540
transform -1 0 16836 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _2323_
timestamp 1704896540
transform 1 0 16376 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2324__56
timestamp 1704896540
transform 1 0 13892 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _2324_
timestamp 1704896540
transform 1 0 14168 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2325__57
timestamp 1704896540
transform -1 0 13708 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _2325_
timestamp 1704896540
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2326__58
timestamp 1704896540
transform 1 0 10304 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _2326_
timestamp 1704896540
transform 1 0 10580 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _2327_
timestamp 1704896540
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2327__59
timestamp 1704896540
transform -1 0 9936 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2328__60
timestamp 1704896540
transform -1 0 9660 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _2328_
timestamp 1704896540
transform 1 0 9384 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2329__15
timestamp 1704896540
transform -1 0 25668 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2329_
timestamp 1704896540
transform 1 0 25024 0 1 544
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2330__16
timestamp 1704896540
transform -1 0 25392 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2330_
timestamp 1704896540
transform 1 0 24840 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_2  _2331_
timestamp 1704896540
transform 1 0 23920 0 1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2331__17
timestamp 1704896540
transform 1 0 23460 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2332__18
timestamp 1704896540
transform 1 0 23460 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2332_
timestamp 1704896540
transform 1 0 23828 0 1 544
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_2  _2333_
timestamp 1704896540
transform 1 0 23644 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2333__19
timestamp 1704896540
transform 1 0 22908 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2334_
timestamp 1704896540
transform 1 0 22172 0 1 544
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2334__20
timestamp 1704896540
transform -1 0 22908 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2335__21
timestamp 1704896540
transform -1 0 22632 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2335_
timestamp 1704896540
transform 1 0 22448 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_2  _2336_
timestamp 1704896540
transform 1 0 21160 0 1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2336__22
timestamp 1704896540
transform -1 0 21804 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2337__23
timestamp 1704896540
transform -1 0 21528 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2337_
timestamp 1704896540
transform 1 0 21252 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2338__24
timestamp 1704896540
transform -1 0 21160 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2338_
timestamp 1704896540
transform 1 0 19964 0 1 544
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2339__25
timestamp 1704896540
transform 1 0 19228 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2339_
timestamp 1704896540
transform 1 0 19504 0 1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_2  _2340_
timestamp 1704896540
transform 1 0 19688 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2340__26
timestamp 1704896540
transform 1 0 18952 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2341_
timestamp 1704896540
transform 1 0 18676 0 1 544
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2341__27
timestamp 1704896540
transform -1 0 18952 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2342_
timestamp 1704896540
transform 1 0 18492 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2342__28
timestamp 1704896540
transform 1 0 17664 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2343_
timestamp 1704896540
transform 1 0 17388 0 1 544
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2343__29
timestamp 1704896540
transform -1 0 17664 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2344_
timestamp 1704896540
transform 1 0 18676 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2345_
timestamp 1704896540
transform 1 0 18768 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2346_
timestamp 1704896540
transform 1 0 18860 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2347_
timestamp 1704896540
transform 1 0 17296 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2348_
timestamp 1704896540
transform 1 0 17848 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2349_
timestamp 1704896540
transform 1 0 19320 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2350_
timestamp 1704896540
transform 1 0 17756 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2351_
timestamp 1704896540
transform 1 0 18676 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _2352__30
timestamp 1704896540
transform -1 0 20240 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _2352_
timestamp 1704896540
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _2353_
timestamp 1704896540
transform 1 0 24288 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2353__31
timestamp 1704896540
transform 1 0 24012 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2354__32
timestamp 1704896540
transform 1 0 24196 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _2354_
timestamp 1704896540
transform 1 0 24472 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2355__33
timestamp 1704896540
transform -1 0 22448 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _2355_
timestamp 1704896540
transform 1 0 22080 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _2356_
timestamp 1704896540
transform 1 0 22540 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2356__34
timestamp 1704896540
transform -1 0 22816 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2357__35
timestamp 1704896540
transform -1 0 19228 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _2357_
timestamp 1704896540
transform 1 0 18860 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2358__36
timestamp 1704896540
transform -1 0 19596 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _2358_
timestamp 1704896540
transform 1 0 19228 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _2359_
timestamp 1704896540
transform 1 0 17756 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2359__37
timestamp 1704896540
transform -1 0 18584 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2360_
timestamp 1704896540
transform 1 0 19044 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2361_
timestamp 1704896540
transform -1 0 8556 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2362_
timestamp 1704896540
transform 1 0 6900 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2363_
timestamp 1704896540
transform 1 0 4876 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2364_
timestamp 1704896540
transform 1 0 3404 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2365_
timestamp 1704896540
transform 1 0 1656 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2366_
timestamp 1704896540
transform 1 0 828 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2367_
timestamp 1704896540
transform 1 0 828 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2368_
timestamp 1704896540
transform 1 0 2760 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2369_
timestamp 1704896540
transform 1 0 3220 0 1 29920
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2370_
timestamp 1704896540
transform -1 0 15824 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2371_
timestamp 1704896540
transform 1 0 16192 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2372_
timestamp 1704896540
transform 1 0 16100 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2373_
timestamp 1704896540
transform 1 0 13616 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2374_
timestamp 1704896540
transform -1 0 14996 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2375_
timestamp 1704896540
transform 1 0 10948 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2376_
timestamp 1704896540
transform 1 0 8556 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2377_
timestamp 1704896540
transform 1 0 9200 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2378_
timestamp 1704896540
transform -1 0 3128 0 1 29920
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11408 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1704896540
transform 1 0 2576 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 15732 0 -1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1704896540
transform -1 0 11132 0 1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1704896540
transform 1 0 19228 0 -1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9200 0 1 17952
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_1_clk
timestamp 1704896540
transform -1 0 6992 0 -1 21216
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_2_clk
timestamp 1704896540
transform -1 0 2668 0 -1 21216
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_3_clk
timestamp 1704896540
transform 1 0 3220 0 1 25568
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_4_clk
timestamp 1704896540
transform -1 0 5428 0 -1 29920
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_5_clk
timestamp 1704896540
transform 1 0 8924 0 1 27744
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_6_clk
timestamp 1704896540
transform 1 0 10856 0 1 25568
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_7_clk
timestamp 1704896540
transform 1 0 13892 0 -1 22304
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_8_clk
timestamp 1704896540
transform -1 0 17848 0 -1 27744
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_9_clk
timestamp 1704896540
transform -1 0 22264 0 -1 28832
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_10_clk
timestamp 1704896540
transform 1 0 25300 0 -1 25568
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_11_clk
timestamp 1704896540
transform 1 0 25944 0 1 20128
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_12_clk
timestamp 1704896540
transform 1 0 17572 0 1 19040
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_13_clk
timestamp 1704896540
transform 1 0 21252 0 -1 14688
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_14_clk
timestamp 1704896540
transform 1 0 25300 0 -1 14688
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_15_clk
timestamp 1704896540
transform 1 0 23828 0 1 9248
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_16_clk
timestamp 1704896540
transform -1 0 18584 0 -1 8160
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_17_clk
timestamp 1704896540
transform 1 0 13708 0 1 13600
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_18_clk
timestamp 1704896540
transform 1 0 10488 0 1 8160
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_19_clk
timestamp 1704896540
transform -1 0 4232 0 -1 8160
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_20_clk
timestamp 1704896540
transform 1 0 3680 0 -1 14688
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 828 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1288 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_12 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1656 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_29
timestamp 1704896540
transform 1 0 3220 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_37
timestamp 1704896540
transform 1 0 3956 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5796 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_65
timestamp 1704896540
transform 1 0 6532 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 1704896540
transform 1 0 8188 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8372 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_91
timestamp 1704896540
transform 1 0 8924 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_95
timestamp 1704896540
transform 1 0 9292 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1704896540
transform 1 0 10580 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_126
timestamp 1704896540
transform 1 0 12144 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_141
timestamp 1704896540
transform 1 0 13524 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_145
timestamp 1704896540
transform 1 0 13892 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_159
timestamp 1704896540
transform 1 0 15180 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_167
timestamp 1704896540
transform 1 0 15916 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_169
timestamp 1704896540
transform 1 0 16100 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_210
timestamp 1704896540
transform 1 0 19872 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_231 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 21804 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_248
timestamp 1704896540
transform 1 0 23368 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_279
timestamp 1704896540
transform 1 0 26220 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_281
timestamp 1704896540
transform 1 0 26404 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_3
timestamp 1704896540
transform 1 0 828 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_63
timestamp 1704896540
transform 1 0 6348 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_277
timestamp 1704896540
transform 1 0 26036 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_281
timestamp 1704896540
transform 1 0 26404 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_3
timestamp 1704896540
transform 1 0 828 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_20
timestamp 1704896540
transform 1 0 2392 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1704896540
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_35
timestamp 1704896540
transform 1 0 3772 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_47
timestamp 1704896540
transform 1 0 4876 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_78
timestamp 1704896540
transform 1 0 7728 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_85
timestamp 1704896540
transform 1 0 8372 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_91
timestamp 1704896540
transform 1 0 8924 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_105
timestamp 1704896540
transform 1 0 10212 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_109
timestamp 1704896540
transform 1 0 10580 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_113
timestamp 1704896540
transform 1 0 10948 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1704896540
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_144
timestamp 1704896540
transform 1 0 13800 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_150
timestamp 1704896540
transform 1 0 14352 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_155
timestamp 1704896540
transform 1 0 14812 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_178
timestamp 1704896540
transform 1 0 16928 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_182
timestamp 1704896540
transform 1 0 17296 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1704896540
transform 1 0 17940 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1704896540
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_219
timestamp 1704896540
transform 1 0 20700 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_246
timestamp 1704896540
transform 1 0 23184 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_253
timestamp 1704896540
transform 1 0 23828 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_273 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 25668 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_285
timestamp 1704896540
transform 1 0 26772 0 1 1632
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1704896540
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_15
timestamp 1704896540
transform 1 0 1932 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_35
timestamp 1704896540
transform 1 0 3772 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_49
timestamp 1704896540
transform 1 0 5060 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_95
timestamp 1704896540
transform 1 0 9292 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_108
timestamp 1704896540
transform 1 0 10488 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_116
timestamp 1704896540
transform 1 0 11224 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_123
timestamp 1704896540
transform 1 0 11868 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_127
timestamp 1704896540
transform 1 0 12236 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_131
timestamp 1704896540
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_143
timestamp 1704896540
transform 1 0 13708 0 -1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_148
timestamp 1704896540
transform 1 0 14168 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_175
timestamp 1704896540
transform 1 0 16652 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_183
timestamp 1704896540
transform 1 0 17388 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_192
timestamp 1704896540
transform 1 0 18216 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_202
timestamp 1704896540
transform 1 0 19136 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_208
timestamp 1704896540
transform 1 0 19688 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_215
timestamp 1704896540
transform 1 0 20332 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_221
timestamp 1704896540
transform 1 0 20884 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_225
timestamp 1704896540
transform 1 0 21252 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_231
timestamp 1704896540
transform 1 0 21804 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_238
timestamp 1704896540
transform 1 0 22448 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_247
timestamp 1704896540
transform 1 0 23276 0 -1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_253
timestamp 1704896540
transform 1 0 23828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_265
timestamp 1704896540
transform 1 0 24932 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_277
timestamp 1704896540
transform 1 0 26036 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_281
timestamp 1704896540
transform 1 0 26404 0 -1 2720
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1704896540
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1704896540
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1704896540
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_29
timestamp 1704896540
transform 1 0 3220 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_33
timestamp 1704896540
transform 1 0 3588 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_37
timestamp 1704896540
transform 1 0 3956 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_60
timestamp 1704896540
transform 1 0 6072 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_70
timestamp 1704896540
transform 1 0 6992 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_78
timestamp 1704896540
transform 1 0 7728 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_82
timestamp 1704896540
transform 1 0 8096 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_88
timestamp 1704896540
transform 1 0 8648 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_96
timestamp 1704896540
transform 1 0 9384 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_114
timestamp 1704896540
transform 1 0 11040 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_118
timestamp 1704896540
transform 1 0 11408 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_126
timestamp 1704896540
transform 1 0 12144 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_136
timestamp 1704896540
transform 1 0 13064 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_152
timestamp 1704896540
transform 1 0 14536 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_168
timestamp 1704896540
transform 1 0 16008 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1704896540
transform 1 0 18492 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_202
timestamp 1704896540
transform 1 0 19136 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_206
timestamp 1704896540
transform 1 0 19504 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_212
timestamp 1704896540
transform 1 0 20056 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_216
timestamp 1704896540
transform 1 0 20424 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_221
timestamp 1704896540
transform 1 0 20884 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_247
timestamp 1704896540
transform 1 0 23276 0 1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_269
timestamp 1704896540
transform 1 0 25300 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_281
timestamp 1704896540
transform 1 0 26404 0 1 2720
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1704896540
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1704896540
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_27
timestamp 1704896540
transform 1 0 3036 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_42
timestamp 1704896540
transform 1 0 4416 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_49
timestamp 1704896540
transform 1 0 5060 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1704896540
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_57
timestamp 1704896540
transform 1 0 5796 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_63
timestamp 1704896540
transform 1 0 6348 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_72
timestamp 1704896540
transform 1 0 7176 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_78
timestamp 1704896540
transform 1 0 7728 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_82
timestamp 1704896540
transform 1 0 8096 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_86
timestamp 1704896540
transform 1 0 8464 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_92
timestamp 1704896540
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1704896540
transform 1 0 10212 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1704896540
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_116
timestamp 1704896540
transform 1 0 11224 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_122
timestamp 1704896540
transform 1 0 11776 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_134
timestamp 1704896540
transform 1 0 12880 0 -1 3808
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_146
timestamp 1704896540
transform 1 0 13984 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_158
timestamp 1704896540
transform 1 0 15088 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_169
timestamp 1704896540
transform 1 0 16100 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_177
timestamp 1704896540
transform 1 0 16836 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_185
timestamp 1704896540
transform 1 0 17572 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_195
timestamp 1704896540
transform 1 0 18492 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_201
timestamp 1704896540
transform 1 0 19044 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_205
timestamp 1704896540
transform 1 0 19412 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_222
timestamp 1704896540
transform 1 0 20976 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_225
timestamp 1704896540
transform 1 0 21252 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_232
timestamp 1704896540
transform 1 0 21896 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_244
timestamp 1704896540
transform 1 0 23000 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_272
timestamp 1704896540
transform 1 0 25576 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_281
timestamp 1704896540
transform 1 0 26404 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_3
timestamp 1704896540
transform 1 0 828 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_7
timestamp 1704896540
transform 1 0 1196 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_23
timestamp 1704896540
transform 1 0 2668 0 1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_44
timestamp 1704896540
transform 1 0 4600 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_56
timestamp 1704896540
transform 1 0 5704 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_63
timestamp 1704896540
transform 1 0 6348 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1704896540
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_93
timestamp 1704896540
transform 1 0 9108 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_111
timestamp 1704896540
transform 1 0 10764 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_121
timestamp 1704896540
transform 1 0 11684 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_129
timestamp 1704896540
transform 1 0 12420 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_134
timestamp 1704896540
transform 1 0 12880 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_141
timestamp 1704896540
transform 1 0 13524 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_150
timestamp 1704896540
transform 1 0 14352 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_156
timestamp 1704896540
transform 1 0 14904 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_165
timestamp 1704896540
transform 1 0 15732 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_188
timestamp 1704896540
transform 1 0 17848 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_210
timestamp 1704896540
transform 1 0 19872 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_221
timestamp 1704896540
transform 1 0 20884 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_227
timestamp 1704896540
transform 1 0 21436 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_231
timestamp 1704896540
transform 1 0 21804 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_240
timestamp 1704896540
transform 1 0 22632 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_247
timestamp 1704896540
transform 1 0 23276 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_253
timestamp 1704896540
transform 1 0 23828 0 1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_270
timestamp 1704896540
transform 1 0 25392 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_282
timestamp 1704896540
transform 1 0 26496 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_288
timestamp 1704896540
transform 1 0 27048 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_3
timestamp 1704896540
transform 1 0 828 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_18
timestamp 1704896540
transform 1 0 2208 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_24
timestamp 1704896540
transform 1 0 2760 0 -1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_29
timestamp 1704896540
transform 1 0 3220 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_41
timestamp 1704896540
transform 1 0 4324 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1704896540
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1704896540
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_73
timestamp 1704896540
transform 1 0 7268 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_89
timestamp 1704896540
transform 1 0 8740 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_95
timestamp 1704896540
transform 1 0 9292 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_102
timestamp 1704896540
transform 1 0 9936 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_108
timestamp 1704896540
transform 1 0 10488 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_113
timestamp 1704896540
transform 1 0 10948 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_135
timestamp 1704896540
transform 1 0 12972 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_143
timestamp 1704896540
transform 1 0 13708 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_160
timestamp 1704896540
transform 1 0 15272 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_169
timestamp 1704896540
transform 1 0 16100 0 -1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_175
timestamp 1704896540
transform 1 0 16652 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_199
timestamp 1704896540
transform 1 0 18860 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_215
timestamp 1704896540
transform 1 0 20332 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1704896540
transform 1 0 21068 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_225
timestamp 1704896540
transform 1 0 21252 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_249
timestamp 1704896540
transform 1 0 23460 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_262
timestamp 1704896540
transform 1 0 24656 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_266
timestamp 1704896540
transform 1 0 25024 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_272
timestamp 1704896540
transform 1 0 25576 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_281
timestamp 1704896540
transform 1 0 26404 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_3
timestamp 1704896540
transform 1 0 828 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_34
timestamp 1704896540
transform 1 0 3680 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_54
timestamp 1704896540
transform 1 0 5520 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_58
timestamp 1704896540
transform 1 0 5888 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_72
timestamp 1704896540
transform 1 0 7176 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_78
timestamp 1704896540
transform 1 0 7728 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_82
timestamp 1704896540
transform 1 0 8096 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_85
timestamp 1704896540
transform 1 0 8372 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_91
timestamp 1704896540
transform 1 0 8924 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_95
timestamp 1704896540
transform 1 0 9292 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_103
timestamp 1704896540
transform 1 0 10028 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_121
timestamp 1704896540
transform 1 0 11684 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_153
timestamp 1704896540
transform 1 0 14628 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_157
timestamp 1704896540
transform 1 0 14996 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_166
timestamp 1704896540
transform 1 0 15824 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_186
timestamp 1704896540
transform 1 0 17664 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_192
timestamp 1704896540
transform 1 0 18216 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_197
timestamp 1704896540
transform 1 0 18676 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_233
timestamp 1704896540
transform 1 0 21988 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_238
timestamp 1704896540
transform 1 0 22448 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1704896540
transform 1 0 23644 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_253
timestamp 1704896540
transform 1 0 23828 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_265
timestamp 1704896540
transform 1 0 24932 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_282
timestamp 1704896540
transform 1 0 26496 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_288
timestamp 1704896540
transform 1 0 27048 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_3
timestamp 1704896540
transform 1 0 828 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_10
timestamp 1704896540
transform 1 0 1472 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_18
timestamp 1704896540
transform 1 0 2208 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_23
timestamp 1704896540
transform 1 0 2668 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_30
timestamp 1704896540
transform 1 0 3312 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_57
timestamp 1704896540
transform 1 0 5796 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1704896540
transform 1 0 10764 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1704896540
transform 1 0 10948 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_125
timestamp 1704896540
transform 1 0 12052 0 -1 5984
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_132
timestamp 1704896540
transform 1 0 12696 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_149
timestamp 1704896540
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_166
timestamp 1704896540
transform 1 0 15824 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_169
timestamp 1704896540
transform 1 0 16100 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_196
timestamp 1704896540
transform 1 0 18584 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_203
timestamp 1704896540
transform 1 0 19228 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_207
timestamp 1704896540
transform 1 0 19596 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_220
timestamp 1704896540
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_235
timestamp 1704896540
transform 1 0 22172 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_242
timestamp 1704896540
transform 1 0 22816 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_246
timestamp 1704896540
transform 1 0 23184 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_274
timestamp 1704896540
transform 1 0 25760 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_281
timestamp 1704896540
transform 1 0 26404 0 -1 5984
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1704896540
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_15
timestamp 1704896540
transform 1 0 1932 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_23
timestamp 1704896540
transform 1 0 2668 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_42
timestamp 1704896540
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_50
timestamp 1704896540
transform 1 0 5152 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_61
timestamp 1704896540
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_66
timestamp 1704896540
transform 1 0 6624 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_70
timestamp 1704896540
transform 1 0 6992 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_81
timestamp 1704896540
transform 1 0 8004 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_85
timestamp 1704896540
transform 1 0 8372 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_113
timestamp 1704896540
transform 1 0 10948 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_131
timestamp 1704896540
transform 1 0 12604 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_157
timestamp 1704896540
transform 1 0 14996 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_166
timestamp 1704896540
transform 1 0 15824 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_175
timestamp 1704896540
transform 1 0 16652 0 1 5984
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_184
timestamp 1704896540
transform 1 0 17480 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1704896540
transform 1 0 18676 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1704896540
transform 1 0 19780 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_221
timestamp 1704896540
transform 1 0 20884 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1704896540
transform 1 0 23644 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_253
timestamp 1704896540
transform 1 0 23828 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_262
timestamp 1704896540
transform 1 0 24656 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_271
timestamp 1704896540
transform 1 0 25484 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_279
timestamp 1704896540
transform 1 0 26220 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_287
timestamp 1704896540
transform 1 0 26956 0 1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1704896540
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_15
timestamp 1704896540
transform 1 0 1932 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_34
timestamp 1704896540
transform 1 0 3680 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_54
timestamp 1704896540
transform 1 0 5520 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_57
timestamp 1704896540
transform 1 0 5796 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_71
timestamp 1704896540
transform 1 0 7084 0 -1 7072
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_82
timestamp 1704896540
transform 1 0 8096 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_94
timestamp 1704896540
transform 1 0 9200 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_106
timestamp 1704896540
transform 1 0 10304 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_134
timestamp 1704896540
transform 1 0 12880 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_139
timestamp 1704896540
transform 1 0 13340 0 -1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_144
timestamp 1704896540
transform 1 0 13800 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_156
timestamp 1704896540
transform 1 0 14904 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_169
timestamp 1704896540
transform 1 0 16100 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_215
timestamp 1704896540
transform 1 0 20332 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1704896540
transform 1 0 21068 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_225
timestamp 1704896540
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_231
timestamp 1704896540
transform 1 0 21804 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_243
timestamp 1704896540
transform 1 0 22908 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_254
timestamp 1704896540
transform 1 0 23920 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_258
timestamp 1704896540
transform 1 0 24288 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1704896540
transform 1 0 26220 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_286
timestamp 1704896540
transform 1 0 26864 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_19
timestamp 1704896540
transform 1 0 2300 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1704896540
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_36
timestamp 1704896540
transform 1 0 3864 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_50
timestamp 1704896540
transform 1 0 5152 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_69
timestamp 1704896540
transform 1 0 6900 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_90
timestamp 1704896540
transform 1 0 8832 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_94
timestamp 1704896540
transform 1 0 9200 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_111
timestamp 1704896540
transform 1 0 10764 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_119
timestamp 1704896540
transform 1 0 11500 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_135
timestamp 1704896540
transform 1 0 12972 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1704896540
transform 1 0 13340 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_150
timestamp 1704896540
transform 1 0 14352 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_154
timestamp 1704896540
transform 1 0 14720 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_162
timestamp 1704896540
transform 1 0 15456 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_173
timestamp 1704896540
transform 1 0 16468 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_183
timestamp 1704896540
transform 1 0 17388 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1704896540
transform 1 0 18492 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_202
timestamp 1704896540
transform 1 0 19136 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_215
timestamp 1704896540
transform 1 0 20332 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_223
timestamp 1704896540
transform 1 0 21068 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_237
timestamp 1704896540
transform 1 0 22356 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_243
timestamp 1704896540
transform 1 0 22908 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1704896540
transform 1 0 23644 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_253
timestamp 1704896540
transform 1 0 23828 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_278
timestamp 1704896540
transform 1 0 26128 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_288
timestamp 1704896540
transform 1 0 27048 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1704896540
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_15
timestamp 1704896540
transform 1 0 1932 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_24
timestamp 1704896540
transform 1 0 2760 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_28
timestamp 1704896540
transform 1 0 3128 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_43
timestamp 1704896540
transform 1 0 4508 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1704896540
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_60
timestamp 1704896540
transform 1 0 6072 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_110
timestamp 1704896540
transform 1 0 10672 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_118
timestamp 1704896540
transform 1 0 11408 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_203
timestamp 1704896540
transform 1 0 19228 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_211
timestamp 1704896540
transform 1 0 19964 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_246
timestamp 1704896540
transform 1 0 23184 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_258
timestamp 1704896540
transform 1 0 24288 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_3
timestamp 1704896540
transform 1 0 828 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_9
timestamp 1704896540
transform 1 0 1380 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_29
timestamp 1704896540
transform 1 0 3220 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_63
timestamp 1704896540
transform 1 0 6348 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_74
timestamp 1704896540
transform 1 0 7360 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_82
timestamp 1704896540
transform 1 0 8096 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_85
timestamp 1704896540
transform 1 0 8372 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_119
timestamp 1704896540
transform 1 0 11500 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_137
timestamp 1704896540
transform 1 0 13156 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_141
timestamp 1704896540
transform 1 0 13524 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_145
timestamp 1704896540
transform 1 0 13892 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_151
timestamp 1704896540
transform 1 0 14444 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_155
timestamp 1704896540
transform 1 0 14812 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_164
timestamp 1704896540
transform 1 0 15640 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_170
timestamp 1704896540
transform 1 0 16192 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_174
timestamp 1704896540
transform 1 0 16560 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_182
timestamp 1704896540
transform 1 0 17296 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_187
timestamp 1704896540
transform 1 0 17756 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_194
timestamp 1704896540
transform 1 0 18400 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_200
timestamp 1704896540
transform 1 0 18952 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_210
timestamp 1704896540
transform 1 0 19872 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_221
timestamp 1704896540
transform 1 0 20884 0 1 8160
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_231
timestamp 1704896540
transform 1 0 21804 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_243
timestamp 1704896540
transform 1 0 22908 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 1704896540
transform 1 0 23644 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_269
timestamp 1704896540
transform 1 0 25300 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_288
timestamp 1704896540
transform 1 0 27048 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_19
timestamp 1704896540
transform 1 0 2300 0 -1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_34
timestamp 1704896540
transform 1 0 3680 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_46
timestamp 1704896540
transform 1 0 4784 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_54
timestamp 1704896540
transform 1 0 5520 0 -1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1704896540
transform 1 0 5796 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_69
timestamp 1704896540
transform 1 0 6900 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_78
timestamp 1704896540
transform 1 0 7728 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_94
timestamp 1704896540
transform 1 0 9200 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_102
timestamp 1704896540
transform 1 0 9936 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_108
timestamp 1704896540
transform 1 0 10488 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_137
timestamp 1704896540
transform 1 0 13156 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_151
timestamp 1704896540
transform 1 0 14444 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_159
timestamp 1704896540
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_169
timestamp 1704896540
transform 1 0 16100 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_177
timestamp 1704896540
transform 1 0 16836 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_195
timestamp 1704896540
transform 1 0 18492 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 1704896540
transform 1 0 21068 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_225
timestamp 1704896540
transform 1 0 21252 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_229
timestamp 1704896540
transform 1 0 21620 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_234
timestamp 1704896540
transform 1 0 22080 0 -1 9248
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1704896540
transform 1 0 828 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_20
timestamp 1704896540
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_32
timestamp 1704896540
transform 1 0 3496 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_36
timestamp 1704896540
transform 1 0 3864 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_45
timestamp 1704896540
transform 1 0 4692 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_50
timestamp 1704896540
transform 1 0 5152 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_74
timestamp 1704896540
transform 1 0 7360 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_85
timestamp 1704896540
transform 1 0 8372 0 1 9248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_102
timestamp 1704896540
transform 1 0 9936 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_114
timestamp 1704896540
transform 1 0 11040 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_123
timestamp 1704896540
transform 1 0 11868 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1704896540
transform 1 0 13340 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_176
timestamp 1704896540
transform 1 0 16744 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_188
timestamp 1704896540
transform 1 0 17848 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_200
timestamp 1704896540
transform 1 0 18952 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_218
timestamp 1704896540
transform 1 0 20608 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_272
timestamp 1704896540
transform 1 0 25576 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1704896540
transform 1 0 828 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_15
timestamp 1704896540
transform 1 0 1932 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_57
timestamp 1704896540
transform 1 0 5796 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_83
timestamp 1704896540
transform 1 0 8188 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_92
timestamp 1704896540
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_118
timestamp 1704896540
transform 1 0 11408 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_130
timestamp 1704896540
transform 1 0 12512 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_134
timestamp 1704896540
transform 1 0 12880 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_138
timestamp 1704896540
transform 1 0 13248 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_150
timestamp 1704896540
transform 1 0 14352 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_166
timestamp 1704896540
transform 1 0 15824 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_188
timestamp 1704896540
transform 1 0 17848 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_201
timestamp 1704896540
transform 1 0 19044 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_213
timestamp 1704896540
transform 1 0 20148 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_221
timestamp 1704896540
transform 1 0 20884 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_225
timestamp 1704896540
transform 1 0 21252 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 1704896540
transform 1 0 26220 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1704896540
transform 1 0 828 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_15
timestamp 1704896540
transform 1 0 1932 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1704896540
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_33
timestamp 1704896540
transform 1 0 3588 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_48
timestamp 1704896540
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_67
timestamp 1704896540
transform 1 0 6716 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_76
timestamp 1704896540
transform 1 0 7544 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_85
timestamp 1704896540
transform 1 0 8372 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_99
timestamp 1704896540
transform 1 0 9660 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_103
timestamp 1704896540
transform 1 0 10028 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_110
timestamp 1704896540
transform 1 0 10672 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1704896540
transform 1 0 13340 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_141
timestamp 1704896540
transform 1 0 13524 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_153
timestamp 1704896540
transform 1 0 14628 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_159
timestamp 1704896540
transform 1 0 15180 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 1704896540
transform 1 0 18492 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_217
timestamp 1704896540
transform 1 0 20516 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_250
timestamp 1704896540
transform 1 0 23552 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_253
timestamp 1704896540
transform 1 0 23828 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_287
timestamp 1704896540
transform 1 0 26956 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_3
timestamp 1704896540
transform 1 0 828 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_15
timestamp 1704896540
transform 1 0 1932 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_19
timestamp 1704896540
transform 1 0 2300 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1704896540
transform 1 0 3036 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1704896540
transform 1 0 4140 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1704896540
transform 1 0 5244 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1704896540
transform 1 0 5612 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_57
timestamp 1704896540
transform 1 0 5796 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_66
timestamp 1704896540
transform 1 0 6624 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_78
timestamp 1704896540
transform 1 0 7728 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_90
timestamp 1704896540
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_100
timestamp 1704896540
transform 1 0 9752 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_108
timestamp 1704896540
transform 1 0 10488 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_113
timestamp 1704896540
transform 1 0 10948 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_130
timestamp 1704896540
transform 1 0 12512 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_136
timestamp 1704896540
transform 1 0 13064 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1704896540
transform 1 0 15916 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_172
timestamp 1704896540
transform 1 0 16376 0 -1 11424
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_187
timestamp 1704896540
transform 1 0 17756 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_225
timestamp 1704896540
transform 1 0 21252 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 1704896540
transform 1 0 26220 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_3
timestamp 1704896540
transform 1 0 828 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_7
timestamp 1704896540
transform 1 0 1196 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_24
timestamp 1704896540
transform 1 0 2760 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_50
timestamp 1704896540
transform 1 0 5152 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_56
timestamp 1704896540
transform 1 0 5704 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_79
timestamp 1704896540
transform 1 0 7820 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1704896540
transform 1 0 8188 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_114
timestamp 1704896540
transform 1 0 11040 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_137
timestamp 1704896540
transform 1 0 13156 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_141
timestamp 1704896540
transform 1 0 13524 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_171
timestamp 1704896540
transform 1 0 16284 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_194
timestamp 1704896540
transform 1 0 18400 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_197
timestamp 1704896540
transform 1 0 18676 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_205
timestamp 1704896540
transform 1 0 19412 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_209
timestamp 1704896540
transform 1 0 19780 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_223
timestamp 1704896540
transform 1 0 21068 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_227
timestamp 1704896540
transform 1 0 21436 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_245
timestamp 1704896540
transform 1 0 23092 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 1704896540
transform 1 0 23644 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_35
timestamp 1704896540
transform 1 0 3772 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_46
timestamp 1704896540
transform 1 0 4784 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1704896540
transform 1 0 5612 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1704896540
transform 1 0 10764 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_142
timestamp 1704896540
transform 1 0 13616 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_150
timestamp 1704896540
transform 1 0 14352 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_157
timestamp 1704896540
transform 1 0 14996 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_163
timestamp 1704896540
transform 1 0 15548 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1704896540
transform 1 0 16100 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_181
timestamp 1704896540
transform 1 0 17204 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_189
timestamp 1704896540
transform 1 0 17940 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_204
timestamp 1704896540
transform 1 0 19320 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_216
timestamp 1704896540
transform 1 0 20424 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_225
timestamp 1704896540
transform 1 0 21252 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_258
timestamp 1704896540
transform 1 0 24288 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_277
timestamp 1704896540
transform 1 0 26036 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_3
timestamp 1704896540
transform 1 0 828 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_19
timestamp 1704896540
transform 1 0 2300 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_25
timestamp 1704896540
transform 1 0 2852 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_35
timestamp 1704896540
transform 1 0 3772 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_53
timestamp 1704896540
transform 1 0 5428 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_62
timestamp 1704896540
transform 1 0 6256 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_72
timestamp 1704896540
transform 1 0 7176 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_85
timestamp 1704896540
transform 1 0 8372 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_113
timestamp 1704896540
transform 1 0 10948 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1704896540
transform 1 0 13340 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_157
timestamp 1704896540
transform 1 0 14996 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_175
timestamp 1704896540
transform 1 0 16652 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_191
timestamp 1704896540
transform 1 0 18124 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_216
timestamp 1704896540
transform 1 0 20424 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_269
timestamp 1704896540
transform 1 0 25300 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_3
timestamp 1704896540
transform 1 0 828 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_7
timestamp 1704896540
transform 1 0 1196 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_16
timestamp 1704896540
transform 1 0 2024 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_35
timestamp 1704896540
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1704896540
transform 1 0 5612 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_57
timestamp 1704896540
transform 1 0 5796 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_110
timestamp 1704896540
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_116
timestamp 1704896540
transform 1 0 11224 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_128
timestamp 1704896540
transform 1 0 12328 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_140
timestamp 1704896540
transform 1 0 13432 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_153
timestamp 1704896540
transform 1 0 14628 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_169
timestamp 1704896540
transform 1 0 16100 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_188
timestamp 1704896540
transform 1 0 17848 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_202
timestamp 1704896540
transform 1 0 19136 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1704896540
transform 1 0 21068 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 1704896540
transform 1 0 26220 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1704896540
transform 1 0 3036 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_45
timestamp 1704896540
transform 1 0 4692 0 1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_52
timestamp 1704896540
transform 1 0 5336 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_64
timestamp 1704896540
transform 1 0 6440 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_68
timestamp 1704896540
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_93
timestamp 1704896540
transform 1 0 9108 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_120
timestamp 1704896540
transform 1 0 11592 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_141
timestamp 1704896540
transform 1 0 13524 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_165
timestamp 1704896540
transform 1 0 15732 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_169
timestamp 1704896540
transform 1 0 16100 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_184
timestamp 1704896540
transform 1 0 17480 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_210
timestamp 1704896540
transform 1 0 19872 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_222
timestamp 1704896540
transform 1 0 20976 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_267
timestamp 1704896540
transform 1 0 25116 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_287
timestamp 1704896540
transform 1 0 26956 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_3
timestamp 1704896540
transform 1 0 828 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_11
timestamp 1704896540
transform 1 0 1564 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_16
timestamp 1704896540
transform 1 0 2024 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_22
timestamp 1704896540
transform 1 0 2576 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_50
timestamp 1704896540
transform 1 0 5152 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_72
timestamp 1704896540
transform 1 0 7176 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_86
timestamp 1704896540
transform 1 0 8464 0 -1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_99
timestamp 1704896540
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1704896540
transform 1 0 10764 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_113
timestamp 1704896540
transform 1 0 10948 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_146
timestamp 1704896540
transform 1 0 13984 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_165
timestamp 1704896540
transform 1 0 15732 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_217
timestamp 1704896540
transform 1 0 20516 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_240
timestamp 1704896540
transform 1 0 22632 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_267
timestamp 1704896540
transform 1 0 25116 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_19
timestamp 1704896540
transform 1 0 2300 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1704896540
transform 1 0 3036 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_29
timestamp 1704896540
transform 1 0 3220 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_37
timestamp 1704896540
transform 1 0 3956 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_81
timestamp 1704896540
transform 1 0 8004 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_133
timestamp 1704896540
transform 1 0 12788 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_137
timestamp 1704896540
transform 1 0 13156 0 1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1704896540
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_153
timestamp 1704896540
transform 1 0 14628 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_157
timestamp 1704896540
transform 1 0 14996 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_162
timestamp 1704896540
transform 1 0 15456 0 1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 1704896540
transform 1 0 18676 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_209
timestamp 1704896540
transform 1 0 19780 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_221
timestamp 1704896540
transform 1 0 20884 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_233
timestamp 1704896540
transform 1 0 21988 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_253
timestamp 1704896540
transform 1 0 23828 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_270
timestamp 1704896540
transform 1 0 25392 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_3
timestamp 1704896540
transform 1 0 828 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_10
timestamp 1704896540
transform 1 0 1472 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_31
timestamp 1704896540
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_52
timestamp 1704896540
transform 1 0 5336 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_57
timestamp 1704896540
transform 1 0 5796 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_76
timestamp 1704896540
transform 1 0 7544 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_101
timestamp 1704896540
transform 1 0 9844 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_109
timestamp 1704896540
transform 1 0 10580 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_113
timestamp 1704896540
transform 1 0 10948 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_121
timestamp 1704896540
transform 1 0 11684 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_157
timestamp 1704896540
transform 1 0 14996 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_166
timestamp 1704896540
transform 1 0 15824 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_169
timestamp 1704896540
transform 1 0 16100 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_187
timestamp 1704896540
transform 1 0 17756 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_195
timestamp 1704896540
transform 1 0 18492 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_219
timestamp 1704896540
transform 1 0 20700 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1704896540
transform 1 0 21068 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_236
timestamp 1704896540
transform 1 0 22264 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_248
timestamp 1704896540
transform 1 0 23368 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_260
timestamp 1704896540
transform 1 0 24472 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_264
timestamp 1704896540
transform 1 0 24840 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_3
timestamp 1704896540
transform 1 0 828 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_22
timestamp 1704896540
transform 1 0 2576 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_37
timestamp 1704896540
transform 1 0 3956 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_54
timestamp 1704896540
transform 1 0 5520 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_62
timestamp 1704896540
transform 1 0 6256 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_73
timestamp 1704896540
transform 1 0 7268 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_81
timestamp 1704896540
transform 1 0 8004 0 1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1704896540
transform 1 0 8372 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_97
timestamp 1704896540
transform 1 0 9476 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_103
timestamp 1704896540
transform 1 0 10028 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1704896540
transform 1 0 13340 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_146
timestamp 1704896540
transform 1 0 13984 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_150
timestamp 1704896540
transform 1 0 14352 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_158
timestamp 1704896540
transform 1 0 15088 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_165
timestamp 1704896540
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_177
timestamp 1704896540
transform 1 0 16836 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_183
timestamp 1704896540
transform 1 0 17388 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_191
timestamp 1704896540
transform 1 0 18124 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1704896540
transform 1 0 18492 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_197
timestamp 1704896540
transform 1 0 18676 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_222
timestamp 1704896540
transform 1 0 20976 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_241
timestamp 1704896540
transform 1 0 22724 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_282
timestamp 1704896540
transform 1 0 26496 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_288
timestamp 1704896540
transform 1 0 27048 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1704896540
transform 1 0 828 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_15
timestamp 1704896540
transform 1 0 1932 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_39
timestamp 1704896540
transform 1 0 4140 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_54
timestamp 1704896540
transform 1 0 5520 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_57
timestamp 1704896540
transform 1 0 5796 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_76
timestamp 1704896540
transform 1 0 7544 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_83
timestamp 1704896540
transform 1 0 8188 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_107
timestamp 1704896540
transform 1 0 10396 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1704896540
transform 1 0 10764 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_113
timestamp 1704896540
transform 1 0 10948 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_123
timestamp 1704896540
transform 1 0 11868 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_131
timestamp 1704896540
transform 1 0 12604 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1704896540
transform 1 0 15916 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_206
timestamp 1704896540
transform 1 0 19504 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 1704896540
transform 1 0 21068 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_240
timestamp 1704896540
transform 1 0 22632 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_260
timestamp 1704896540
transform 1 0 24472 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_272
timestamp 1704896540
transform 1 0 25576 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_278
timestamp 1704896540
transform 1 0 26128 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_281
timestamp 1704896540
transform 1 0 26404 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_3
timestamp 1704896540
transform 1 0 828 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_7
timestamp 1704896540
transform 1 0 1196 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_15
timestamp 1704896540
transform 1 0 1932 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_45
timestamp 1704896540
transform 1 0 4692 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_59
timestamp 1704896540
transform 1 0 5980 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_85
timestamp 1704896540
transform 1 0 8372 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_108
timestamp 1704896540
transform 1 0 10488 0 1 16864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_117
timestamp 1704896540
transform 1 0 11316 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_129
timestamp 1704896540
transform 1 0 12420 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_137
timestamp 1704896540
transform 1 0 13156 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_141
timestamp 1704896540
transform 1 0 13524 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_167
timestamp 1704896540
transform 1 0 15916 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_187
timestamp 1704896540
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_197
timestamp 1704896540
transform 1 0 18676 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_223
timestamp 1704896540
transform 1 0 21068 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_231
timestamp 1704896540
transform 1 0 21804 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_239
timestamp 1704896540
transform 1 0 22540 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_247
timestamp 1704896540
transform 1 0 23276 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1704896540
transform 1 0 23644 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_256
timestamp 1704896540
transform 1 0 24104 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_265
timestamp 1704896540
transform 1 0 24932 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_271
timestamp 1704896540
transform 1 0 25484 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_26
timestamp 1704896540
transform 1 0 2944 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_54
timestamp 1704896540
transform 1 0 5520 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_63
timestamp 1704896540
transform 1 0 6348 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_90
timestamp 1704896540
transform 1 0 8832 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_97
timestamp 1704896540
transform 1 0 9476 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_107
timestamp 1704896540
transform 1 0 10396 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1704896540
transform 1 0 10764 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_116
timestamp 1704896540
transform 1 0 11224 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_122
timestamp 1704896540
transform 1 0 11776 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_142
timestamp 1704896540
transform 1 0 13616 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_169
timestamp 1704896540
transform 1 0 16100 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_182
timestamp 1704896540
transform 1 0 17296 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_186
timestamp 1704896540
transform 1 0 17664 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_190
timestamp 1704896540
transform 1 0 18032 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_194
timestamp 1704896540
transform 1 0 18400 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_203
timestamp 1704896540
transform 1 0 19228 0 -1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_212
timestamp 1704896540
transform 1 0 20056 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_238
timestamp 1704896540
transform 1 0 22448 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_265
timestamp 1704896540
transform 1 0 24932 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_284
timestamp 1704896540
transform 1 0 26680 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_288
timestamp 1704896540
transform 1 0 27048 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_3
timestamp 1704896540
transform 1 0 828 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_9
timestamp 1704896540
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_13
timestamp 1704896540
transform 1 0 1748 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_24
timestamp 1704896540
transform 1 0 2760 0 1 17952
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1704896540
transform 1 0 3220 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_41
timestamp 1704896540
transform 1 0 4324 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_52
timestamp 1704896540
transform 1 0 5336 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_67
timestamp 1704896540
transform 1 0 6716 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_79
timestamp 1704896540
transform 1 0 7820 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1704896540
transform 1 0 8188 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_85
timestamp 1704896540
transform 1 0 8372 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_93
timestamp 1704896540
transform 1 0 9108 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_130
timestamp 1704896540
transform 1 0 12512 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_136
timestamp 1704896540
transform 1 0 13064 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_141
timestamp 1704896540
transform 1 0 13524 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_147
timestamp 1704896540
transform 1 0 14076 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_176
timestamp 1704896540
transform 1 0 16744 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_197
timestamp 1704896540
transform 1 0 18676 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_216
timestamp 1704896540
transform 1 0 20424 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_230
timestamp 1704896540
transform 1 0 21712 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 1704896540
transform 1 0 23644 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_272
timestamp 1704896540
transform 1 0 25576 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1704896540
transform 1 0 828 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_15
timestamp 1704896540
transform 1 0 1932 0 -1 19040
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_37
timestamp 1704896540
transform 1 0 3956 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_49
timestamp 1704896540
transform 1 0 5060 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1704896540
transform 1 0 5612 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_63
timestamp 1704896540
transform 1 0 6348 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_113
timestamp 1704896540
transform 1 0 10948 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_122
timestamp 1704896540
transform 1 0 11776 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_126
timestamp 1704896540
transform 1 0 12144 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_133
timestamp 1704896540
transform 1 0 12788 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_165
timestamp 1704896540
transform 1 0 15732 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_201
timestamp 1704896540
transform 1 0 19044 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_223
timestamp 1704896540
transform 1 0 21068 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_247
timestamp 1704896540
transform 1 0 23276 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_259
timestamp 1704896540
transform 1 0 24380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_271
timestamp 1704896540
transform 1 0 25484 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_275
timestamp 1704896540
transform 1 0 25852 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_279
timestamp 1704896540
transform 1 0 26220 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_281
timestamp 1704896540
transform 1 0 26404 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_3
timestamp 1704896540
transform 1 0 828 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_8
timestamp 1704896540
transform 1 0 1288 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_12
timestamp 1704896540
transform 1 0 1656 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_32
timestamp 1704896540
transform 1 0 3496 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_36
timestamp 1704896540
transform 1 0 3864 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_43
timestamp 1704896540
transform 1 0 4508 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_59
timestamp 1704896540
transform 1 0 5980 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 1704896540
transform 1 0 8188 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_85
timestamp 1704896540
transform 1 0 8372 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_92
timestamp 1704896540
transform 1 0 9016 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_115
timestamp 1704896540
transform 1 0 11132 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_176
timestamp 1704896540
transform 1 0 16744 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_197
timestamp 1704896540
transform 1 0 18676 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_201
timestamp 1704896540
transform 1 0 19044 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_251
timestamp 1704896540
transform 1 0 23644 0 1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_253
timestamp 1704896540
transform 1 0 23828 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_265
timestamp 1704896540
transform 1 0 24932 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_271
timestamp 1704896540
transform 1 0 25484 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_288
timestamp 1704896540
transform 1 0 27048 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_27
timestamp 1704896540
transform 1 0 3036 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_40
timestamp 1704896540
transform 1 0 4232 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_50
timestamp 1704896540
transform 1 0 5152 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_57
timestamp 1704896540
transform 1 0 5796 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_74
timestamp 1704896540
transform 1 0 7360 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_86
timestamp 1704896540
transform 1 0 8464 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_93
timestamp 1704896540
transform 1 0 9108 0 -1 20128
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_100
timestamp 1704896540
transform 1 0 9752 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_127
timestamp 1704896540
transform 1 0 12236 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_154
timestamp 1704896540
transform 1 0 14720 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_162
timestamp 1704896540
transform 1 0 15456 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_169
timestamp 1704896540
transform 1 0 16100 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_178
timestamp 1704896540
transform 1 0 16928 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_198
timestamp 1704896540
transform 1 0 18768 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_218
timestamp 1704896540
transform 1 0 20608 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_232
timestamp 1704896540
transform 1 0 21896 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_273
timestamp 1704896540
transform 1 0 25668 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_279
timestamp 1704896540
transform 1 0 26220 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_281
timestamp 1704896540
transform 1 0 26404 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_3
timestamp 1704896540
transform 1 0 828 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_11
timestamp 1704896540
transform 1 0 1564 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_26
timestamp 1704896540
transform 1 0 2944 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_29
timestamp 1704896540
transform 1 0 3220 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_39
timestamp 1704896540
transform 1 0 4140 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_44
timestamp 1704896540
transform 1 0 4600 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_51
timestamp 1704896540
transform 1 0 5244 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_71
timestamp 1704896540
transform 1 0 7084 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_81
timestamp 1704896540
transform 1 0 8004 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_101
timestamp 1704896540
transform 1 0 9844 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_118
timestamp 1704896540
transform 1 0 11408 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_130
timestamp 1704896540
transform 1 0 12512 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_138
timestamp 1704896540
transform 1 0 13248 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_144
timestamp 1704896540
transform 1 0 13800 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_165
timestamp 1704896540
transform 1 0 15732 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_183
timestamp 1704896540
transform 1 0 17388 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_190
timestamp 1704896540
transform 1 0 18032 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_212
timestamp 1704896540
transform 1 0 20056 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_242
timestamp 1704896540
transform 1 0 22816 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_253
timestamp 1704896540
transform 1 0 23828 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_273
timestamp 1704896540
transform 1 0 25668 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_287
timestamp 1704896540
transform 1 0 26956 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_3
timestamp 1704896540
transform 1 0 828 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_26
timestamp 1704896540
transform 1 0 2944 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_30
timestamp 1704896540
transform 1 0 3312 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_54
timestamp 1704896540
transform 1 0 5520 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_57
timestamp 1704896540
transform 1 0 5796 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_91
timestamp 1704896540
transform 1 0 8924 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_100
timestamp 1704896540
transform 1 0 9752 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_113
timestamp 1704896540
transform 1 0 10948 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_131
timestamp 1704896540
transform 1 0 12604 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_155
timestamp 1704896540
transform 1 0 14812 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_163
timestamp 1704896540
transform 1 0 15548 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 1704896540
transform 1 0 15916 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_169
timestamp 1704896540
transform 1 0 16100 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_173
timestamp 1704896540
transform 1 0 16468 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_177
timestamp 1704896540
transform 1 0 16836 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_190
timestamp 1704896540
transform 1 0 18032 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 1704896540
transform 1 0 21068 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_240
timestamp 1704896540
transform 1 0 22632 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_246
timestamp 1704896540
transform 1 0 23184 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_252
timestamp 1704896540
transform 1 0 23736 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_260
timestamp 1704896540
transform 1 0 24472 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_269
timestamp 1704896540
transform 1 0 25300 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_273
timestamp 1704896540
transform 1 0 25668 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 1704896540
transform 1 0 26220 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_26
timestamp 1704896540
transform 1 0 2944 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_50
timestamp 1704896540
transform 1 0 5152 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_81
timestamp 1704896540
transform 1 0 8004 0 1 21216
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_90
timestamp 1704896540
transform 1 0 8832 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_102
timestamp 1704896540
transform 1 0 9936 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_120
timestamp 1704896540
transform 1 0 11592 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_150
timestamp 1704896540
transform 1 0 14352 0 1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_156
timestamp 1704896540
transform 1 0 14904 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_168
timestamp 1704896540
transform 1 0 16008 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_179
timestamp 1704896540
transform 1 0 17020 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_205
timestamp 1704896540
transform 1 0 19412 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_221
timestamp 1704896540
transform 1 0 20884 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_231
timestamp 1704896540
transform 1 0 21804 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_238
timestamp 1704896540
transform 1 0 22448 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_248
timestamp 1704896540
transform 1 0 23368 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_285
timestamp 1704896540
transform 1 0 26772 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_3
timestamp 1704896540
transform 1 0 828 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_16
timestamp 1704896540
transform 1 0 2024 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_24
timestamp 1704896540
transform 1 0 2760 0 -1 22304
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_30
timestamp 1704896540
transform 1 0 3312 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_42
timestamp 1704896540
transform 1 0 4416 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_46
timestamp 1704896540
transform 1 0 4784 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_71
timestamp 1704896540
transform 1 0 7084 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_91
timestamp 1704896540
transform 1 0 8924 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_98
timestamp 1704896540
transform 1 0 9568 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_110
timestamp 1704896540
transform 1 0 10672 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_116
timestamp 1704896540
transform 1 0 11224 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_120
timestamp 1704896540
transform 1 0 11592 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_137
timestamp 1704896540
transform 1 0 13156 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_173
timestamp 1704896540
transform 1 0 16468 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_179
timestamp 1704896540
transform 1 0 17020 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_184
timestamp 1704896540
transform 1 0 17480 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_189
timestamp 1704896540
transform 1 0 17940 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_197
timestamp 1704896540
transform 1 0 18676 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_222
timestamp 1704896540
transform 1 0 20976 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_225
timestamp 1704896540
transform 1 0 21252 0 -1 22304
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_263
timestamp 1704896540
transform 1 0 24748 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_275
timestamp 1704896540
transform 1 0 25852 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_279
timestamp 1704896540
transform 1 0 26220 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_281
timestamp 1704896540
transform 1 0 26404 0 -1 22304
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1704896540
transform 1 0 828 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_15
timestamp 1704896540
transform 1 0 1932 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_19
timestamp 1704896540
transform 1 0 2300 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1704896540
transform 1 0 3036 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_35
timestamp 1704896540
transform 1 0 3772 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 1704896540
transform 1 0 8188 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_85
timestamp 1704896540
transform 1 0 8372 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_102
timestamp 1704896540
transform 1 0 9936 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_121
timestamp 1704896540
transform 1 0 11684 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_131
timestamp 1704896540
transform 1 0 12604 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_151
timestamp 1704896540
transform 1 0 14444 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_190
timestamp 1704896540
transform 1 0 18032 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_197
timestamp 1704896540
transform 1 0 18676 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_205
timestamp 1704896540
transform 1 0 19412 0 1 22304
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_216
timestamp 1704896540
transform 1 0 20424 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_228
timestamp 1704896540
transform 1 0 21528 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_236
timestamp 1704896540
transform 1 0 22264 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_249
timestamp 1704896540
transform 1 0 23460 0 1 22304
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_256
timestamp 1704896540
transform 1 0 24104 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_268
timestamp 1704896540
transform 1 0 25208 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_287
timestamp 1704896540
transform 1 0 26956 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_19
timestamp 1704896540
transform 1 0 2300 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_34
timestamp 1704896540
transform 1 0 3680 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_47
timestamp 1704896540
transform 1 0 4876 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 1704896540
transform 1 0 5612 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_57
timestamp 1704896540
transform 1 0 5796 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_94
timestamp 1704896540
transform 1 0 9200 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_108
timestamp 1704896540
transform 1 0 10488 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_113
timestamp 1704896540
transform 1 0 10948 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_121
timestamp 1704896540
transform 1 0 11684 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_128
timestamp 1704896540
transform 1 0 12328 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_155
timestamp 1704896540
transform 1 0 14812 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_159
timestamp 1704896540
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_178
timestamp 1704896540
transform 1 0 16928 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_188
timestamp 1704896540
transform 1 0 17848 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_203
timestamp 1704896540
transform 1 0 19228 0 -1 23392
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_239
timestamp 1704896540
transform 1 0 22540 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_254
timestamp 1704896540
transform 1 0 23920 0 -1 23392
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_263
timestamp 1704896540
transform 1 0 24748 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_275
timestamp 1704896540
transform 1 0 25852 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_279
timestamp 1704896540
transform 1 0 26220 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_16
timestamp 1704896540
transform 1 0 2024 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1704896540
transform 1 0 3036 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_29
timestamp 1704896540
transform 1 0 3220 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_69
timestamp 1704896540
transform 1 0 6900 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_80
timestamp 1704896540
transform 1 0 7912 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_93
timestamp 1704896540
transform 1 0 9108 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_138
timestamp 1704896540
transform 1 0 13248 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_149
timestamp 1704896540
transform 1 0 14260 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_162
timestamp 1704896540
transform 1 0 15456 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_166
timestamp 1704896540
transform 1 0 15824 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_192
timestamp 1704896540
transform 1 0 18216 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_218
timestamp 1704896540
transform 1 0 20608 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_234
timestamp 1704896540
transform 1 0 22080 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_253
timestamp 1704896540
transform 1 0 23828 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_277
timestamp 1704896540
transform 1 0 26036 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_281
timestamp 1704896540
transform 1 0 26404 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_285
timestamp 1704896540
transform 1 0 26772 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_3
timestamp 1704896540
transform 1 0 828 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_11
timestamp 1704896540
transform 1 0 1564 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_21
timestamp 1704896540
transform 1 0 2484 0 -1 24480
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_26
timestamp 1704896540
transform 1 0 2944 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_38
timestamp 1704896540
transform 1 0 4048 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_47
timestamp 1704896540
transform 1 0 4876 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1704896540
transform 1 0 5612 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_57
timestamp 1704896540
transform 1 0 5796 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_91
timestamp 1704896540
transform 1 0 8924 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_101
timestamp 1704896540
transform 1 0 9844 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_109
timestamp 1704896540
transform 1 0 10580 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_125
timestamp 1704896540
transform 1 0 12052 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_137
timestamp 1704896540
transform 1 0 13156 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_145
timestamp 1704896540
transform 1 0 13892 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_164
timestamp 1704896540
transform 1 0 15640 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_178
timestamp 1704896540
transform 1 0 16928 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_184
timestamp 1704896540
transform 1 0 17480 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_190
timestamp 1704896540
transform 1 0 18032 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_198
timestamp 1704896540
transform 1 0 18768 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_204
timestamp 1704896540
transform 1 0 19320 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_220
timestamp 1704896540
transform 1 0 20792 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_225
timestamp 1704896540
transform 1 0 21252 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_235
timestamp 1704896540
transform 1 0 22172 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_239
timestamp 1704896540
transform 1 0 22540 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_265
timestamp 1704896540
transform 1 0 24932 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_281
timestamp 1704896540
transform 1 0 26404 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_287
timestamp 1704896540
transform 1 0 26956 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_3
timestamp 1704896540
transform 1 0 828 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_8
timestamp 1704896540
transform 1 0 1288 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_17
timestamp 1704896540
transform 1 0 2116 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_29
timestamp 1704896540
transform 1 0 3220 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_37
timestamp 1704896540
transform 1 0 3956 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_44
timestamp 1704896540
transform 1 0 4600 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_52
timestamp 1704896540
transform 1 0 5336 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_80
timestamp 1704896540
transform 1 0 7912 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_85
timestamp 1704896540
transform 1 0 8372 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_120
timestamp 1704896540
transform 1 0 11592 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_141
timestamp 1704896540
transform 1 0 13524 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_163
timestamp 1704896540
transform 1 0 15548 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_188
timestamp 1704896540
transform 1 0 17848 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_194
timestamp 1704896540
transform 1 0 18400 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_197
timestamp 1704896540
transform 1 0 18676 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_220
timestamp 1704896540
transform 1 0 20792 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_228
timestamp 1704896540
transform 1 0 21528 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_235
timestamp 1704896540
transform 1 0 22172 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_243
timestamp 1704896540
transform 1 0 22908 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_251
timestamp 1704896540
transform 1 0 23644 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_270
timestamp 1704896540
transform 1 0 25392 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_40
timestamp 1704896540
transform 1 0 4232 0 -1 25568
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 1704896540
transform 1 0 5796 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_74
timestamp 1704896540
transform 1 0 7360 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_83
timestamp 1704896540
transform 1 0 8188 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_94
timestamp 1704896540
transform 1 0 9200 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_110
timestamp 1704896540
transform 1 0 10672 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_113
timestamp 1704896540
transform 1 0 10948 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_136
timestamp 1704896540
transform 1 0 13064 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_144
timestamp 1704896540
transform 1 0 13800 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_148
timestamp 1704896540
transform 1 0 14168 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_159
timestamp 1704896540
transform 1 0 15180 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 1704896540
transform 1 0 15916 0 -1 25568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_169
timestamp 1704896540
transform 1 0 16100 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_181
timestamp 1704896540
transform 1 0 17204 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_203
timestamp 1704896540
transform 1 0 19228 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_211
timestamp 1704896540
transform 1 0 19964 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_216
timestamp 1704896540
transform 1 0 20424 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_225
timestamp 1704896540
transform 1 0 21252 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_246
timestamp 1704896540
transform 1 0 23184 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_256
timestamp 1704896540
transform 1 0 24104 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_260
timestamp 1704896540
transform 1 0 24472 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_265
timestamp 1704896540
transform 1 0 24932 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_281
timestamp 1704896540
transform 1 0 26404 0 -1 25568
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1704896540
transform 1 0 828 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_15
timestamp 1704896540
transform 1 0 1932 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_40
timestamp 1704896540
transform 1 0 4232 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_44
timestamp 1704896540
transform 1 0 4600 0 1 25568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_52
timestamp 1704896540
transform 1 0 5336 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_64
timestamp 1704896540
transform 1 0 6440 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_77
timestamp 1704896540
transform 1 0 7636 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_101
timestamp 1704896540
transform 1 0 9844 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_109
timestamp 1704896540
transform 1 0 10580 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_131
timestamp 1704896540
transform 1 0 12604 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_167
timestamp 1704896540
transform 1 0 15916 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_171
timestamp 1704896540
transform 1 0 16284 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_177
timestamp 1704896540
transform 1 0 16836 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_185
timestamp 1704896540
transform 1 0 17572 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_193
timestamp 1704896540
transform 1 0 18308 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_217
timestamp 1704896540
transform 1 0 20516 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_227
timestamp 1704896540
transform 1 0 21436 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_235
timestamp 1704896540
transform 1 0 22172 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_281
timestamp 1704896540
transform 1 0 26404 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_3
timestamp 1704896540
transform 1 0 828 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_9
timestamp 1704896540
transform 1 0 1380 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_17
timestamp 1704896540
transform 1 0 2116 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_32
timestamp 1704896540
transform 1 0 3496 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_36
timestamp 1704896540
transform 1 0 3864 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_43
timestamp 1704896540
transform 1 0 4508 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_49
timestamp 1704896540
transform 1 0 5060 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_64
timestamp 1704896540
transform 1 0 6440 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_82
timestamp 1704896540
transform 1 0 8096 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_96
timestamp 1704896540
transform 1 0 9384 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_106
timestamp 1704896540
transform 1 0 10304 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_113
timestamp 1704896540
transform 1 0 10948 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_129
timestamp 1704896540
transform 1 0 12420 0 -1 26656
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_138
timestamp 1704896540
transform 1 0 13248 0 -1 26656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_150
timestamp 1704896540
transform 1 0 14352 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_162
timestamp 1704896540
transform 1 0 15456 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_205
timestamp 1704896540
transform 1 0 19412 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_215
timestamp 1704896540
transform 1 0 20332 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_223
timestamp 1704896540
transform 1 0 21068 0 -1 26656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_232
timestamp 1704896540
transform 1 0 21896 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_244
timestamp 1704896540
transform 1 0 23000 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_248
timestamp 1704896540
transform 1 0 23368 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_252
timestamp 1704896540
transform 1 0 23736 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_258
timestamp 1704896540
transform 1 0 24288 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_267
timestamp 1704896540
transform 1 0 25116 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_271
timestamp 1704896540
transform 1 0 25484 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_275
timestamp 1704896540
transform 1 0 25852 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_279
timestamp 1704896540
transform 1 0 26220 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_281
timestamp 1704896540
transform 1 0 26404 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_26
timestamp 1704896540
transform 1 0 2944 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_29
timestamp 1704896540
transform 1 0 3220 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_40
timestamp 1704896540
transform 1 0 4232 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_50
timestamp 1704896540
transform 1 0 5152 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_54
timestamp 1704896540
transform 1 0 5520 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_85
timestamp 1704896540
transform 1 0 8372 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_113
timestamp 1704896540
transform 1 0 10948 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_123
timestamp 1704896540
transform 1 0 11868 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_131
timestamp 1704896540
transform 1 0 12604 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_139
timestamp 1704896540
transform 1 0 13340 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_148
timestamp 1704896540
transform 1 0 14168 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_160
timestamp 1704896540
transform 1 0 15272 0 1 26656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_168
timestamp 1704896540
transform 1 0 16008 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_180
timestamp 1704896540
transform 1 0 17112 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_188
timestamp 1704896540
transform 1 0 17848 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_205
timestamp 1704896540
transform 1 0 19412 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_217
timestamp 1704896540
transform 1 0 20516 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_230
timestamp 1704896540
transform 1 0 21712 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_236
timestamp 1704896540
transform 1 0 22264 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_244
timestamp 1704896540
transform 1 0 23000 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_248
timestamp 1704896540
transform 1 0 23368 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_270
timestamp 1704896540
transform 1 0 25392 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_288
timestamp 1704896540
transform 1 0 27048 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_3
timestamp 1704896540
transform 1 0 828 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_11
timestamp 1704896540
transform 1 0 1564 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_17
timestamp 1704896540
transform 1 0 2116 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_31
timestamp 1704896540
transform 1 0 3404 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_48
timestamp 1704896540
transform 1 0 4968 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_79
timestamp 1704896540
transform 1 0 7820 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_99
timestamp 1704896540
transform 1 0 9660 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_107
timestamp 1704896540
transform 1 0 10396 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_111
timestamp 1704896540
transform 1 0 10764 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_113
timestamp 1704896540
transform 1 0 10948 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_119
timestamp 1704896540
transform 1 0 11500 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_126
timestamp 1704896540
transform 1 0 12144 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_134
timestamp 1704896540
transform 1 0 12880 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_138
timestamp 1704896540
transform 1 0 13248 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_144
timestamp 1704896540
transform 1 0 13800 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_148
timestamp 1704896540
transform 1 0 14168 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_152
timestamp 1704896540
transform 1 0 14536 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_157
timestamp 1704896540
transform 1 0 14996 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_161
timestamp 1704896540
transform 1 0 15364 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_165
timestamp 1704896540
transform 1 0 15732 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_175
timestamp 1704896540
transform 1 0 16652 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_220
timestamp 1704896540
transform 1 0 20792 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_225
timestamp 1704896540
transform 1 0 21252 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_245
timestamp 1704896540
transform 1 0 23092 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_254
timestamp 1704896540
transform 1 0 23920 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_281
timestamp 1704896540
transform 1 0 26404 0 -1 27744
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1704896540
transform 1 0 828 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_15
timestamp 1704896540
transform 1 0 1932 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_21
timestamp 1704896540
transform 1 0 2484 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1704896540
transform 1 0 3036 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_32
timestamp 1704896540
transform 1 0 3496 0 1 27744
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_39
timestamp 1704896540
transform 1 0 4140 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_51
timestamp 1704896540
transform 1 0 5244 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_72
timestamp 1704896540
transform 1 0 7176 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_76
timestamp 1704896540
transform 1 0 7544 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_83
timestamp 1704896540
transform 1 0 8188 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_85
timestamp 1704896540
transform 1 0 8372 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_116
timestamp 1704896540
transform 1 0 11224 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_133
timestamp 1704896540
transform 1 0 12788 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_162
timestamp 1704896540
transform 1 0 15456 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_195
timestamp 1704896540
transform 1 0 18492 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_204
timestamp 1704896540
transform 1 0 19320 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_212
timestamp 1704896540
transform 1 0 20056 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_219
timestamp 1704896540
transform 1 0 20700 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_224
timestamp 1704896540
transform 1 0 21160 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_231
timestamp 1704896540
transform 1 0 21804 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_238
timestamp 1704896540
transform 1 0 22448 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_263
timestamp 1704896540
transform 1 0 24748 0 1 27744
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_270
timestamp 1704896540
transform 1 0 25392 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_282
timestamp 1704896540
transform 1 0 26496 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_288
timestamp 1704896540
transform 1 0 27048 0 1 27744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 1704896540
transform 1 0 828 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_15
timestamp 1704896540
transform 1 0 1932 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_37
timestamp 1704896540
transform 1 0 3956 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_41
timestamp 1704896540
transform 1 0 4324 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_47
timestamp 1704896540
transform 1 0 4876 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 1704896540
transform 1 0 5612 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_89
timestamp 1704896540
transform 1 0 8740 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_110
timestamp 1704896540
transform 1 0 10672 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_123
timestamp 1704896540
transform 1 0 11868 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_131
timestamp 1704896540
transform 1 0 12604 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_141
timestamp 1704896540
transform 1 0 13524 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_156
timestamp 1704896540
transform 1 0 14904 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_166
timestamp 1704896540
transform 1 0 15824 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_174
timestamp 1704896540
transform 1 0 16560 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_195
timestamp 1704896540
transform 1 0 18492 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_221
timestamp 1704896540
transform 1 0 20884 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_241
timestamp 1704896540
transform 1 0 22724 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_247
timestamp 1704896540
transform 1 0 23276 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_253
timestamp 1704896540
transform 1 0 23828 0 -1 28832
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_258
timestamp 1704896540
transform 1 0 24288 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_273
timestamp 1704896540
transform 1 0 25668 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_279
timestamp 1704896540
transform 1 0 26220 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_281
timestamp 1704896540
transform 1 0 26404 0 -1 28832
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_3
timestamp 1704896540
transform 1 0 828 0 1 28832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_15
timestamp 1704896540
transform 1 0 1932 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 1704896540
transform 1 0 3036 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_29
timestamp 1704896540
transform 1 0 3220 0 1 28832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_64
timestamp 1704896540
transform 1 0 6440 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_76
timestamp 1704896540
transform 1 0 7544 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_95
timestamp 1704896540
transform 1 0 9292 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_99
timestamp 1704896540
transform 1 0 9660 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_106
timestamp 1704896540
transform 1 0 10304 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_112
timestamp 1704896540
transform 1 0 10856 0 1 28832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_122
timestamp 1704896540
transform 1 0 11776 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_134
timestamp 1704896540
transform 1 0 12880 0 1 28832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_141
timestamp 1704896540
transform 1 0 13524 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_153
timestamp 1704896540
transform 1 0 14628 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_159
timestamp 1704896540
transform 1 0 15180 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_165
timestamp 1704896540
transform 1 0 15732 0 1 28832
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_180
timestamp 1704896540
transform 1 0 17112 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_192
timestamp 1704896540
transform 1 0 18216 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_204
timestamp 1704896540
transform 1 0 19320 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_218
timestamp 1704896540
transform 1 0 20608 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_224
timestamp 1704896540
transform 1 0 21160 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_230
timestamp 1704896540
transform 1 0 21712 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_236
timestamp 1704896540
transform 1 0 22264 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_251
timestamp 1704896540
transform 1 0 23644 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_253
timestamp 1704896540
transform 1 0 23828 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_287
timestamp 1704896540
transform 1 0 26956 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_20
timestamp 1704896540
transform 1 0 2392 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_24
timestamp 1704896540
transform 1 0 2760 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_32
timestamp 1704896540
transform 1 0 3496 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_38
timestamp 1704896540
transform 1 0 4048 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_53
timestamp 1704896540
transform 1 0 5428 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_74
timestamp 1704896540
transform 1 0 7360 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_80
timestamp 1704896540
transform 1 0 7912 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_97
timestamp 1704896540
transform 1 0 9476 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_103
timestamp 1704896540
transform 1 0 10028 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_113
timestamp 1704896540
transform 1 0 10948 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_118
timestamp 1704896540
transform 1 0 11408 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_129
timestamp 1704896540
transform 1 0 12420 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_148
timestamp 1704896540
transform 1 0 14168 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_167
timestamp 1704896540
transform 1 0 15916 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_222
timestamp 1704896540
transform 1 0 20976 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_257
timestamp 1704896540
transform 1 0 24196 0 -1 29920
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_268
timestamp 1704896540
transform 1 0 25208 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_3
timestamp 1704896540
transform 1 0 828 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_62
timestamp 1704896540
transform 1 0 6256 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_82
timestamp 1704896540
transform 1 0 8096 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_113
timestamp 1704896540
transform 1 0 10948 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_133
timestamp 1704896540
transform 1 0 12788 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_144
timestamp 1704896540
transform 1 0 13800 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_164
timestamp 1704896540
transform 1 0 15640 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_184
timestamp 1704896540
transform 1 0 17480 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_197
timestamp 1704896540
transform 1 0 18676 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_234
timestamp 1704896540
transform 1 0 22080 0 1 29920
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_272
timestamp 1704896540
transform 1 0 25576 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_284
timestamp 1704896540
transform 1 0 26680 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_288
timestamp 1704896540
transform 1 0 27048 0 1 29920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_3
timestamp 1704896540
transform 1 0 828 0 -1 31008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_15
timestamp 1704896540
transform 1 0 1932 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_27
timestamp 1704896540
transform 1 0 3036 0 -1 31008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_29
timestamp 1704896540
transform 1 0 3220 0 -1 31008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_41
timestamp 1704896540
transform 1 0 4324 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_53
timestamp 1704896540
transform 1 0 5428 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_73
timestamp 1704896540
transform 1 0 7268 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_83
timestamp 1704896540
transform 1 0 8188 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_88
timestamp 1704896540
transform 1 0 8648 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_93
timestamp 1704896540
transform 1 0 9108 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_101
timestamp 1704896540
transform 1 0 9844 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_110
timestamp 1704896540
transform 1 0 10672 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_113
timestamp 1704896540
transform 1 0 10948 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_121
timestamp 1704896540
transform 1 0 11684 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_129
timestamp 1704896540
transform 1 0 12420 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_138
timestamp 1704896540
transform 1 0 13248 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_150
timestamp 1704896540
transform 1 0 14352 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_158
timestamp 1704896540
transform 1 0 15088 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_166
timestamp 1704896540
transform 1 0 15824 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_179
timestamp 1704896540
transform 1 0 17020 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_183
timestamp 1704896540
transform 1 0 17388 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_195
timestamp 1704896540
transform 1 0 18492 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_204
timestamp 1704896540
transform 1 0 19320 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_222
timestamp 1704896540
transform 1 0 20976 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_225
timestamp 1704896540
transform 1 0 21252 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_233
timestamp 1704896540
transform 1 0 21988 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_238
timestamp 1704896540
transform 1 0 22448 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_244
timestamp 1704896540
transform 1 0 23000 0 -1 31008
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_263
timestamp 1704896540
transform 1 0 24748 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_275
timestamp 1704896540
transform 1 0 25852 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_279
timestamp 1704896540
transform 1 0 26220 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_281
timestamp 1704896540
transform 1 0 26404 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_285
timestamp 1704896540
transform 1 0 26772 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 17020 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1704896540
transform -1 0 15916 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1704896540
transform 1 0 20240 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1704896540
transform 1 0 19964 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1704896540
transform 1 0 24196 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1704896540
transform -1 0 23736 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1704896540
transform -1 0 20976 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1704896540
transform -1 0 19412 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1704896540
transform 1 0 6808 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1704896540
transform -1 0 20332 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1704896540
transform -1 0 13248 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1704896540
transform 1 0 17756 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1704896540
transform 1 0 15548 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1704896540
transform -1 0 7912 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1704896540
transform -1 0 7912 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1704896540
transform -1 0 18584 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1704896540
transform -1 0 16928 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1704896540
transform -1 0 21068 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1704896540
transform -1 0 7084 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1704896540
transform -1 0 19412 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1704896540
transform -1 0 21068 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1704896540
transform 1 0 7728 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1704896540
transform -1 0 7268 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1704896540
transform -1 0 8280 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1704896540
transform -1 0 20884 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1704896540
transform -1 0 20332 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1704896540
transform 1 0 23736 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1704896540
transform -1 0 23368 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1704896540
transform -1 0 19504 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1704896540
transform -1 0 19412 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1704896540
transform 1 0 21344 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1704896540
transform -1 0 20516 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1704896540
transform 1 0 20240 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1704896540
transform -1 0 9108 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1704896540
transform -1 0 5612 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1704896540
transform -1 0 3956 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1704896540
transform -1 0 20240 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1704896540
transform -1 0 20240 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1704896540
transform -1 0 24932 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1704896540
transform -1 0 25668 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1704896540
transform -1 0 27140 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1704896540
transform 1 0 24564 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1704896540
transform -1 0 24932 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1704896540
transform -1 0 27140 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1704896540
transform -1 0 19320 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1704896540
transform -1 0 24564 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1704896540
transform -1 0 22724 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1704896540
transform -1 0 8188 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1704896540
transform -1 0 19228 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1704896540
transform -1 0 9200 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1704896540
transform -1 0 27140 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1704896540
transform -1 0 19412 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1704896540
transform -1 0 27140 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1704896540
transform -1 0 27140 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1704896540
transform 1 0 24196 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1704896540
transform -1 0 26220 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1704896540
transform -1 0 25760 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1704896540
transform 1 0 23552 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1704896540
transform -1 0 27140 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1704896540
transform -1 0 21344 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1704896540
transform -1 0 27140 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1704896540
transform -1 0 25576 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1704896540
transform 1 0 24840 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1704896540
transform -1 0 24564 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1704896540
transform -1 0 27048 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1704896540
transform -1 0 8188 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1704896540
transform 1 0 6164 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1704896540
transform 1 0 17112 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1704896540
transform -1 0 3036 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1704896540
transform -1 0 2024 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1704896540
transform -1 0 23184 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1704896540
transform -1 0 5520 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1704896540
transform -1 0 23736 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1704896540
transform -1 0 4968 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1704896540
transform -1 0 26312 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1704896540
transform 1 0 5520 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1704896540
transform -1 0 2760 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1704896540
transform -1 0 2024 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1704896540
transform -1 0 8188 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1704896540
transform 1 0 9752 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1704896540
transform 1 0 16192 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1704896540
transform -1 0 17204 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1704896540
transform -1 0 20148 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 1704896540
transform -1 0 4048 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1704896540
transform 1 0 17940 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 1704896540
transform -1 0 8004 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1704896540
transform -1 0 6992 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 1704896540
transform 1 0 23460 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 1704896540
transform 1 0 11316 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1704896540
transform -1 0 12880 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 1704896540
transform -1 0 15364 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 1704896540
transform -1 0 13064 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 1704896540
transform -1 0 15824 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 1704896540
transform 1 0 10856 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 1704896540
transform -1 0 13432 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 1704896540
transform -1 0 10764 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 1704896540
transform -1 0 10304 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 1704896540
transform -1 0 27140 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 1704896540
transform 1 0 22080 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 1704896540
transform -1 0 15456 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 1704896540
transform -1 0 10856 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 1704896540
transform -1 0 9936 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 1704896540
transform -1 0 14720 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 1704896540
transform -1 0 13984 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 1704896540
transform -1 0 16836 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 1704896540
transform 1 0 9936 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 1704896540
transform 1 0 12696 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 1704896540
transform 1 0 18676 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 1704896540
transform 1 0 6532 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold110
timestamp 1704896540
transform 1 0 7728 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold111
timestamp 1704896540
transform -1 0 12604 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold112
timestamp 1704896540
transform 1 0 13800 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold113
timestamp 1704896540
transform -1 0 10672 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold114
timestamp 1704896540
transform -1 0 13984 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold115
timestamp 1704896540
transform 1 0 13616 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold116
timestamp 1704896540
transform -1 0 11684 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold117
timestamp 1704896540
transform -1 0 27140 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold118
timestamp 1704896540
transform -1 0 13708 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold119
timestamp 1704896540
transform -1 0 20424 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold120
timestamp 1704896540
transform -1 0 8096 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold121
timestamp 1704896540
transform 1 0 18032 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold122
timestamp 1704896540
transform 1 0 7268 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold123
timestamp 1704896540
transform -1 0 8832 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold124
timestamp 1704896540
transform 1 0 21804 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1704896540
transform -1 0 9108 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1704896540
transform -1 0 10672 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1704896540
transform 1 0 8372 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1704896540
transform 1 0 6348 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1704896540
transform -1 0 22448 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1704896540
transform -1 0 20976 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1704896540
transform -1 0 20608 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1704896540
transform -1 0 18492 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1704896540
transform -1 0 17020 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input10
timestamp 1704896540
transform 1 0 14720 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input11
timestamp 1704896540
transform 1 0 13064 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input12
timestamp 1704896540
transform 1 0 11776 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1704896540
transform 1 0 26496 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input14 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 23828 0 -1 31008
box -38 -48 958 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_56
timestamp 1704896540
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 27416 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_57
timestamp 1704896540
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 27416 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_58
timestamp 1704896540
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 27416 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_59
timestamp 1704896540
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 27416 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_60
timestamp 1704896540
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 27416 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_61
timestamp 1704896540
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 27416 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_62
timestamp 1704896540
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 27416 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_63
timestamp 1704896540
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 27416 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_64
timestamp 1704896540
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 27416 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_65
timestamp 1704896540
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 27416 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_66
timestamp 1704896540
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 27416 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_67
timestamp 1704896540
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 27416 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_68
timestamp 1704896540
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 27416 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_69
timestamp 1704896540
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1704896540
transform -1 0 27416 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_70
timestamp 1704896540
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1704896540
transform -1 0 27416 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_71
timestamp 1704896540
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1704896540
transform -1 0 27416 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_72
timestamp 1704896540
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1704896540
transform -1 0 27416 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_73
timestamp 1704896540
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1704896540
transform -1 0 27416 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_74
timestamp 1704896540
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1704896540
transform -1 0 27416 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_75
timestamp 1704896540
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1704896540
transform -1 0 27416 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_76
timestamp 1704896540
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1704896540
transform -1 0 27416 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_77
timestamp 1704896540
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1704896540
transform -1 0 27416 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_78
timestamp 1704896540
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1704896540
transform -1 0 27416 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_79
timestamp 1704896540
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1704896540
transform -1 0 27416 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_80
timestamp 1704896540
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1704896540
transform -1 0 27416 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_81
timestamp 1704896540
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1704896540
transform -1 0 27416 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_82
timestamp 1704896540
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1704896540
transform -1 0 27416 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_83
timestamp 1704896540
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1704896540
transform -1 0 27416 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_84
timestamp 1704896540
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1704896540
transform -1 0 27416 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_85
timestamp 1704896540
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1704896540
transform -1 0 27416 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_86
timestamp 1704896540
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1704896540
transform -1 0 27416 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_87
timestamp 1704896540
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1704896540
transform -1 0 27416 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_88
timestamp 1704896540
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1704896540
transform -1 0 27416 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_89
timestamp 1704896540
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1704896540
transform -1 0 27416 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_90
timestamp 1704896540
transform 1 0 552 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1704896540
transform -1 0 27416 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_91
timestamp 1704896540
transform 1 0 552 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1704896540
transform -1 0 27416 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_92
timestamp 1704896540
transform 1 0 552 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1704896540
transform -1 0 27416 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_93
timestamp 1704896540
transform 1 0 552 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1704896540
transform -1 0 27416 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_94
timestamp 1704896540
transform 1 0 552 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1704896540
transform -1 0 27416 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_95
timestamp 1704896540
transform 1 0 552 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1704896540
transform -1 0 27416 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_96
timestamp 1704896540
transform 1 0 552 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1704896540
transform -1 0 27416 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_97
timestamp 1704896540
transform 1 0 552 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 1704896540
transform -1 0 27416 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_98
timestamp 1704896540
transform 1 0 552 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 1704896540
transform -1 0 27416 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_99
timestamp 1704896540
transform 1 0 552 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 1704896540
transform -1 0 27416 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_100
timestamp 1704896540
transform 1 0 552 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 1704896540
transform -1 0 27416 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_101
timestamp 1704896540
transform 1 0 552 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 1704896540
transform -1 0 27416 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_102
timestamp 1704896540
transform 1 0 552 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 1704896540
transform -1 0 27416 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_103
timestamp 1704896540
transform 1 0 552 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 1704896540
transform -1 0 27416 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_104
timestamp 1704896540
transform 1 0 552 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 1704896540
transform -1 0 27416 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_105
timestamp 1704896540
transform 1 0 552 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 1704896540
transform -1 0 27416 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_106
timestamp 1704896540
transform 1 0 552 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp 1704896540
transform -1 0 27416 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_107
timestamp 1704896540
transform 1 0 552 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp 1704896540
transform -1 0 27416 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_108
timestamp 1704896540
transform 1 0 552 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp 1704896540
transform -1 0 27416 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_109
timestamp 1704896540
transform 1 0 552 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp 1704896540
transform -1 0 27416 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Left_110
timestamp 1704896540
transform 1 0 552 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Right_54
timestamp 1704896540
transform -1 0 27416 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Left_111
timestamp 1704896540
transform 1 0 552 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Right_55
timestamp 1704896540
transform -1 0 27416 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_112 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_113
timestamp 1704896540
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_114
timestamp 1704896540
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_115
timestamp 1704896540
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_116
timestamp 1704896540
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_117
timestamp 1704896540
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_118
timestamp 1704896540
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_119
timestamp 1704896540
transform 1 0 21160 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_120
timestamp 1704896540
transform 1 0 23736 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_121
timestamp 1704896540
transform 1 0 26312 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_122
timestamp 1704896540
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_123
timestamp 1704896540
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_124
timestamp 1704896540
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_125
timestamp 1704896540
transform 1 0 21160 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_126
timestamp 1704896540
transform 1 0 26312 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_127
timestamp 1704896540
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_128
timestamp 1704896540
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_129
timestamp 1704896540
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_130
timestamp 1704896540
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_131
timestamp 1704896540
transform 1 0 23736 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_132
timestamp 1704896540
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_133
timestamp 1704896540
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_134
timestamp 1704896540
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_135
timestamp 1704896540
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_136
timestamp 1704896540
transform 1 0 26312 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_137
timestamp 1704896540
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_138
timestamp 1704896540
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_139
timestamp 1704896540
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_140
timestamp 1704896540
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_141
timestamp 1704896540
transform 1 0 23736 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_142
timestamp 1704896540
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_143
timestamp 1704896540
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_144
timestamp 1704896540
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_145
timestamp 1704896540
transform 1 0 21160 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_146
timestamp 1704896540
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_147
timestamp 1704896540
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_148
timestamp 1704896540
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_149
timestamp 1704896540
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_150
timestamp 1704896540
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_151
timestamp 1704896540
transform 1 0 23736 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_152
timestamp 1704896540
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_153
timestamp 1704896540
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_154
timestamp 1704896540
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_155
timestamp 1704896540
transform 1 0 21160 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_156
timestamp 1704896540
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_157
timestamp 1704896540
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_158
timestamp 1704896540
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_159
timestamp 1704896540
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_160
timestamp 1704896540
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_161
timestamp 1704896540
transform 1 0 23736 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_162
timestamp 1704896540
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_163
timestamp 1704896540
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_164
timestamp 1704896540
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_165
timestamp 1704896540
transform 1 0 21160 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_166
timestamp 1704896540
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_167
timestamp 1704896540
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_168
timestamp 1704896540
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_169
timestamp 1704896540
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_170
timestamp 1704896540
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_171
timestamp 1704896540
transform 1 0 23736 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_172
timestamp 1704896540
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_173
timestamp 1704896540
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_174
timestamp 1704896540
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_175
timestamp 1704896540
transform 1 0 21160 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_176
timestamp 1704896540
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_177
timestamp 1704896540
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_178
timestamp 1704896540
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_179
timestamp 1704896540
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_180
timestamp 1704896540
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_181
timestamp 1704896540
transform 1 0 23736 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_182
timestamp 1704896540
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_183
timestamp 1704896540
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_184
timestamp 1704896540
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_185
timestamp 1704896540
transform 1 0 21160 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_186
timestamp 1704896540
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_187
timestamp 1704896540
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_188
timestamp 1704896540
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_189
timestamp 1704896540
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_190
timestamp 1704896540
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_191
timestamp 1704896540
transform 1 0 23736 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_192
timestamp 1704896540
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_193
timestamp 1704896540
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_194
timestamp 1704896540
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_195
timestamp 1704896540
transform 1 0 21160 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_196
timestamp 1704896540
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_197
timestamp 1704896540
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_198
timestamp 1704896540
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_199
timestamp 1704896540
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_200
timestamp 1704896540
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_201
timestamp 1704896540
transform 1 0 23736 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_202
timestamp 1704896540
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_203
timestamp 1704896540
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_204
timestamp 1704896540
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_205
timestamp 1704896540
transform 1 0 21160 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_206
timestamp 1704896540
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_207
timestamp 1704896540
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_208
timestamp 1704896540
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_209
timestamp 1704896540
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_210
timestamp 1704896540
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_211
timestamp 1704896540
transform 1 0 23736 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_212
timestamp 1704896540
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_213
timestamp 1704896540
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_214
timestamp 1704896540
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_215
timestamp 1704896540
transform 1 0 21160 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_216
timestamp 1704896540
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_217
timestamp 1704896540
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_218
timestamp 1704896540
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_219
timestamp 1704896540
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_220
timestamp 1704896540
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_221
timestamp 1704896540
transform 1 0 23736 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_222
timestamp 1704896540
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_223
timestamp 1704896540
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_224
timestamp 1704896540
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_225
timestamp 1704896540
transform 1 0 21160 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_226
timestamp 1704896540
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_227
timestamp 1704896540
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_228
timestamp 1704896540
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_229
timestamp 1704896540
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_230
timestamp 1704896540
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_231
timestamp 1704896540
transform 1 0 23736 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_232
timestamp 1704896540
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_233
timestamp 1704896540
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_234
timestamp 1704896540
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_235
timestamp 1704896540
transform 1 0 21160 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_236
timestamp 1704896540
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_237
timestamp 1704896540
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_238
timestamp 1704896540
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_239
timestamp 1704896540
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_240
timestamp 1704896540
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_241
timestamp 1704896540
transform 1 0 23736 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_242
timestamp 1704896540
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_243
timestamp 1704896540
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_244
timestamp 1704896540
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_245
timestamp 1704896540
transform 1 0 21160 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_246
timestamp 1704896540
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_247
timestamp 1704896540
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_248
timestamp 1704896540
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_249
timestamp 1704896540
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_250
timestamp 1704896540
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_251
timestamp 1704896540
transform 1 0 23736 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_252
timestamp 1704896540
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_253
timestamp 1704896540
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_254
timestamp 1704896540
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_255
timestamp 1704896540
transform 1 0 21160 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_256
timestamp 1704896540
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_257
timestamp 1704896540
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_258
timestamp 1704896540
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_259
timestamp 1704896540
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_260
timestamp 1704896540
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_261
timestamp 1704896540
transform 1 0 23736 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_262
timestamp 1704896540
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_263
timestamp 1704896540
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_264
timestamp 1704896540
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_265
timestamp 1704896540
transform 1 0 21160 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_266
timestamp 1704896540
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_267
timestamp 1704896540
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_268
timestamp 1704896540
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_269
timestamp 1704896540
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_270
timestamp 1704896540
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_271
timestamp 1704896540
transform 1 0 23736 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_272
timestamp 1704896540
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_273
timestamp 1704896540
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_274
timestamp 1704896540
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_275
timestamp 1704896540
transform 1 0 21160 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_276
timestamp 1704896540
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_277
timestamp 1704896540
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_278
timestamp 1704896540
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_279
timestamp 1704896540
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_280
timestamp 1704896540
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_281
timestamp 1704896540
transform 1 0 23736 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_282
timestamp 1704896540
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_283
timestamp 1704896540
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_284
timestamp 1704896540
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_285
timestamp 1704896540
transform 1 0 21160 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_286
timestamp 1704896540
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_287
timestamp 1704896540
transform 1 0 3128 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_288
timestamp 1704896540
transform 1 0 8280 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_289
timestamp 1704896540
transform 1 0 13432 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_290
timestamp 1704896540
transform 1 0 18584 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_291
timestamp 1704896540
transform 1 0 23736 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_292
timestamp 1704896540
transform 1 0 5704 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_293
timestamp 1704896540
transform 1 0 10856 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_294
timestamp 1704896540
transform 1 0 16008 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_295
timestamp 1704896540
transform 1 0 21160 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_296
timestamp 1704896540
transform 1 0 26312 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_297
timestamp 1704896540
transform 1 0 3128 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_298
timestamp 1704896540
transform 1 0 8280 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_299
timestamp 1704896540
transform 1 0 13432 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_300
timestamp 1704896540
transform 1 0 18584 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_301
timestamp 1704896540
transform 1 0 23736 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_302
timestamp 1704896540
transform 1 0 5704 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_303
timestamp 1704896540
transform 1 0 10856 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_304
timestamp 1704896540
transform 1 0 16008 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_305
timestamp 1704896540
transform 1 0 21160 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_306
timestamp 1704896540
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_307
timestamp 1704896540
transform 1 0 3128 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_308
timestamp 1704896540
transform 1 0 8280 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_309
timestamp 1704896540
transform 1 0 13432 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_310
timestamp 1704896540
transform 1 0 18584 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_311
timestamp 1704896540
transform 1 0 23736 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_312
timestamp 1704896540
transform 1 0 5704 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_313
timestamp 1704896540
transform 1 0 10856 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_314
timestamp 1704896540
transform 1 0 16008 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_315
timestamp 1704896540
transform 1 0 21160 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_316
timestamp 1704896540
transform 1 0 26312 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_317
timestamp 1704896540
transform 1 0 3128 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_318
timestamp 1704896540
transform 1 0 8280 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_319
timestamp 1704896540
transform 1 0 13432 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_320
timestamp 1704896540
transform 1 0 18584 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_321
timestamp 1704896540
transform 1 0 23736 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_322
timestamp 1704896540
transform 1 0 5704 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_323
timestamp 1704896540
transform 1 0 10856 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_324
timestamp 1704896540
transform 1 0 16008 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_325
timestamp 1704896540
transform 1 0 21160 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_326
timestamp 1704896540
transform 1 0 26312 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_327
timestamp 1704896540
transform 1 0 3128 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_328
timestamp 1704896540
transform 1 0 8280 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_329
timestamp 1704896540
transform 1 0 13432 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_330
timestamp 1704896540
transform 1 0 18584 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_331
timestamp 1704896540
transform 1 0 23736 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_332
timestamp 1704896540
transform 1 0 5704 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_333
timestamp 1704896540
transform 1 0 10856 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_334
timestamp 1704896540
transform 1 0 16008 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_335
timestamp 1704896540
transform 1 0 21160 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_336
timestamp 1704896540
transform 1 0 26312 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_337
timestamp 1704896540
transform 1 0 3128 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_338
timestamp 1704896540
transform 1 0 8280 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_339
timestamp 1704896540
transform 1 0 13432 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_340
timestamp 1704896540
transform 1 0 18584 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_341
timestamp 1704896540
transform 1 0 23736 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_342
timestamp 1704896540
transform 1 0 5704 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_343
timestamp 1704896540
transform 1 0 10856 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_344
timestamp 1704896540
transform 1 0 16008 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_345
timestamp 1704896540
transform 1 0 21160 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_346
timestamp 1704896540
transform 1 0 26312 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_347
timestamp 1704896540
transform 1 0 3128 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_348
timestamp 1704896540
transform 1 0 8280 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_349
timestamp 1704896540
transform 1 0 13432 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_350
timestamp 1704896540
transform 1 0 18584 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_351
timestamp 1704896540
transform 1 0 23736 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_352
timestamp 1704896540
transform 1 0 5704 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_353
timestamp 1704896540
transform 1 0 10856 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_354
timestamp 1704896540
transform 1 0 16008 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_355
timestamp 1704896540
transform 1 0 21160 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_356
timestamp 1704896540
transform 1 0 26312 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_357
timestamp 1704896540
transform 1 0 3128 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_358
timestamp 1704896540
transform 1 0 8280 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_359
timestamp 1704896540
transform 1 0 13432 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_360
timestamp 1704896540
transform 1 0 18584 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_361
timestamp 1704896540
transform 1 0 23736 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_362
timestamp 1704896540
transform 1 0 5704 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_363
timestamp 1704896540
transform 1 0 10856 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_364
timestamp 1704896540
transform 1 0 16008 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_365
timestamp 1704896540
transform 1 0 21160 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_366
timestamp 1704896540
transform 1 0 26312 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_367
timestamp 1704896540
transform 1 0 3128 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_368
timestamp 1704896540
transform 1 0 8280 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_369
timestamp 1704896540
transform 1 0 13432 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_370
timestamp 1704896540
transform 1 0 18584 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_371
timestamp 1704896540
transform 1 0 23736 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_372
timestamp 1704896540
transform 1 0 5704 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_373
timestamp 1704896540
transform 1 0 10856 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_374
timestamp 1704896540
transform 1 0 16008 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_375
timestamp 1704896540
transform 1 0 21160 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_376
timestamp 1704896540
transform 1 0 26312 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_377
timestamp 1704896540
transform 1 0 3128 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_378
timestamp 1704896540
transform 1 0 8280 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_379
timestamp 1704896540
transform 1 0 13432 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_380
timestamp 1704896540
transform 1 0 18584 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_381
timestamp 1704896540
transform 1 0 23736 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_382
timestamp 1704896540
transform 1 0 5704 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_383
timestamp 1704896540
transform 1 0 10856 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_384
timestamp 1704896540
transform 1 0 16008 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_385
timestamp 1704896540
transform 1 0 21160 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_386
timestamp 1704896540
transform 1 0 26312 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_387
timestamp 1704896540
transform 1 0 3128 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_388
timestamp 1704896540
transform 1 0 8280 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_389
timestamp 1704896540
transform 1 0 13432 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_390
timestamp 1704896540
transform 1 0 18584 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_391
timestamp 1704896540
transform 1 0 23736 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_392
timestamp 1704896540
transform 1 0 3128 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_393
timestamp 1704896540
transform 1 0 5704 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_394
timestamp 1704896540
transform 1 0 8280 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_395
timestamp 1704896540
transform 1 0 10856 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_396
timestamp 1704896540
transform 1 0 13432 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_397
timestamp 1704896540
transform 1 0 16008 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_398
timestamp 1704896540
transform 1 0 18584 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_399
timestamp 1704896540
transform 1 0 21160 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_400
timestamp 1704896540
transform 1 0 23736 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_401
timestamp 1704896540
transform 1 0 26312 0 -1 31008
box -38 -48 130 592
<< labels >>
rlabel metal2 s 14064 31008 14064 31008 4 VGND
rlabel metal1 s 13984 30464 13984 30464 4 VPWR
rlabel metal1 s 10672 17646 10672 17646 4 _0003_
rlabel metal1 s 19442 24650 19442 24650 4 _0004_
rlabel metal1 s 19810 23222 19810 23222 4 _0005_
rlabel metal1 s 18752 23562 18752 23562 4 _0006_
rlabel metal1 s 16866 23562 16866 23562 4 _0007_
rlabel metal1 s 8924 22202 8924 22202 4 _0008_
rlabel metal2 s 8689 25806 8689 25806 4 _0009_
rlabel metal2 s 9338 24514 9338 24514 4 _0010_
rlabel metal2 s 9982 23426 9982 23426 4 _0011_
rlabel metal1 s 10437 24718 10437 24718 4 _0012_
rlabel metal1 s 11679 25398 11679 25398 4 _0013_
rlabel metal2 s 11822 23392 11822 23392 4 _0014_
rlabel metal2 s 12650 24514 12650 24514 4 _0015_
rlabel metal2 s 13570 19006 13570 19006 4 _0016_
rlabel metal2 s 12282 19040 12282 19040 4 _0017_
rlabel metal1 s 12558 17306 12558 17306 4 _0018_
rlabel metal2 s 12466 15810 12466 15810 4 _0019_
rlabel metal1 s 13646 15606 13646 15606 4 _0020_
rlabel metal1 s 18844 17034 18844 17034 4 _0021_
rlabel metal1 s 17572 16218 17572 16218 4 _0022_
rlabel metal1 s 19350 15606 19350 15606 4 _0023_
rlabel metal2 s 19545 16014 19545 16014 4 _0024_
rlabel metal1 s 20741 5134 20741 5134 4 _0025_
rlabel metal2 s 25341 5134 25341 5134 4 _0026_
rlabel metal1 s 24778 7242 24778 7242 4 _0027_
rlabel metal1 s 21834 6154 21834 6154 4 _0028_
rlabel metal2 s 21569 7922 21569 7922 4 _0029_
rlabel metal2 s 20010 9282 20010 9282 4 _0030_
rlabel metal2 s 18436 6834 18436 6834 4 _0031_
rlabel metal1 s 17572 8602 17572 8602 4 _0032_
rlabel metal1 s 2576 29478 2576 29478 4 _0033_
rlabel metal1 s 13933 23222 13933 23222 4 _0034_
rlabel metal1 s 13708 20570 13708 20570 4 _0035_
rlabel metal2 s 11274 21454 11274 21454 4 _0036_
rlabel metal2 s 10253 20366 10253 20366 4 _0037_
rlabel metal1 s 11530 30090 11530 30090 4 _0038_
rlabel metal1 s 1932 15674 1932 15674 4 _0039_
rlabel metal1 s 1656 12954 1656 12954 4 _0040_
rlabel metal1 s 3956 13498 3956 13498 4 _0041_
rlabel metal2 s 1426 11492 1426 11492 4 _0042_
rlabel metal2 s 2617 12342 2617 12342 4 _0043_
rlabel metal1 s 4216 13430 4216 13430 4 _0044_
rlabel metal1 s 4043 11594 4043 11594 4 _0045_
rlabel metal1 s 10636 18802 10636 18802 4 _0046_
rlabel metal2 s 10994 17986 10994 17986 4 _0047_
rlabel metal2 s 9057 17102 9057 17102 4 _0048_
rlabel metal1 s 10610 15946 10610 15946 4 _0049_
rlabel metal1 s 5734 20298 5734 20298 4 _0050_
rlabel metal1 s 8050 20570 8050 20570 4 _0051_
rlabel metal2 s 9062 20162 9062 20162 4 _0052_
rlabel metal2 s 6762 19686 6762 19686 4 _0053_
rlabel metal2 s 7682 16898 7682 16898 4 _0054_
rlabel metal2 s 6389 16626 6389 16626 4 _0055_
rlabel metal2 s 7314 18598 7314 18598 4 _0056_
rlabel metal2 s 8602 18598 8602 18598 4 _0057_
rlabel metal1 s 13754 9146 13754 9146 4 _0058_
rlabel metal1 s 13570 10778 13570 10778 4 _0059_
rlabel metal1 s 14674 14042 14674 14042 4 _0060_
rlabel metal1 s 14025 12682 14025 12682 4 _0061_
rlabel metal2 s 15410 11458 15410 11458 4 _0062_
rlabel metal1 s 6844 26418 6844 26418 4 _0063_
rlabel metal2 s 7038 26758 7038 26758 4 _0064_
rlabel metal1 s 7666 24310 7666 24310 4 _0065_
rlabel metal2 s 6210 24514 6210 24514 4 _0066_
rlabel metal1 s 8836 23222 8836 23222 4 _0067_
rlabel metal2 s 6486 23426 6486 23426 4 _0068_
rlabel metal1 s 5883 22474 5883 22474 4 _0069_
rlabel metal2 s 8606 22066 8606 22066 4 _0070_
rlabel metal1 s 11311 9078 11311 9078 4 _0071_
rlabel metal1 s 11592 10234 11592 10234 4 _0072_
rlabel metal1 s 12144 14042 12144 14042 4 _0073_
rlabel metal1 s 11495 12682 11495 12682 4 _0074_
rlabel metal1 s 12466 11866 12466 11866 4 _0075_
rlabel metal2 s 20842 11254 20842 11254 4 _0076_
rlabel metal2 s 25622 28866 25622 28866 4 _0077_
rlabel metal2 s 22581 30158 22581 30158 4 _0078_
rlabel metal1 s 24660 30090 24660 30090 4 _0079_
rlabel metal1 s 24288 28730 24288 28730 4 _0080_
rlabel metal1 s 25672 27574 25672 27574 4 _0081_
rlabel metal1 s 25852 26554 25852 26554 4 _0082_
rlabel metal2 s 25254 25602 25254 25602 4 _0083_
rlabel metal2 s 23418 25806 23418 25806 4 _0084_
rlabel metal1 s 23322 24140 23322 24140 4 _0085_
rlabel metal1 s 24982 23562 24982 23562 4 _0086_
rlabel metal2 s 26082 24514 26082 24514 4 _0087_
rlabel metal2 s 25801 22542 25801 22542 4 _0088_
rlabel metal2 s 15497 12682 15497 12682 4 _0089_
rlabel metal2 s 6941 30158 6941 30158 4 _0090_
rlabel metal1 s 6854 28186 6854 28186 4 _0091_
rlabel metal1 s 8505 29682 8505 29682 4 _0092_
rlabel metal1 s 9598 30090 9598 30090 4 _0093_
rlabel metal1 s 9333 28662 9333 28662 4 _0094_
rlabel metal2 s 11638 27778 11638 27778 4 _0095_
rlabel metal1 s 13289 29750 13289 29750 4 _0096_
rlabel metal2 s 14490 27778 14490 27778 4 _0097_
rlabel metal1 s 15149 30090 15149 30090 4 _0098_
rlabel metal1 s 17070 30090 17070 30090 4 _0099_
rlabel metal2 s 17061 28594 17061 28594 4 _0100_
rlabel metal1 s 16054 27642 16054 27642 4 _0101_
rlabel metal2 s 18538 10268 18538 10268 4 _0102_
rlabel metal1 s 17771 10166 17771 10166 4 _0103_
rlabel metal1 s 16831 13430 16831 13430 4 _0104_
rlabel metal1 s 19131 12682 19131 12682 4 _0105_
rlabel metal2 s 16974 11458 16974 11458 4 _0106_
rlabel metal1 s 18124 14042 18124 14042 4 _0107_
rlabel metal1 s 20669 13430 20669 13430 4 _0108_
rlabel metal2 s 25622 21250 25622 21250 4 _0109_
rlabel metal1 s 24200 22066 24200 22066 4 _0110_
rlabel metal1 s 24936 21386 24936 21386 4 _0111_
rlabel metal1 s 24752 20298 24752 20298 4 _0112_
rlabel metal1 s 24752 19958 24752 19958 4 _0113_
rlabel metal2 s 23970 17714 23970 17714 4 _0114_
rlabel metal2 s 25806 19074 25806 19074 4 _0115_
rlabel metal2 s 26634 17986 26634 17986 4 _0116_
rlabel metal2 s 26082 16898 26082 16898 4 _0117_
rlabel metal1 s 25146 15946 25146 15946 4 _0118_
rlabel metal2 s 22581 14858 22581 14858 4 _0119_
rlabel metal2 s 23598 16558 23598 16558 4 _0120_
rlabel metal1 s 9931 10166 9931 10166 4 _0121_
rlabel metal2 s 10442 11458 10442 11458 4 _0122_
rlabel metal1 s 8827 13362 8827 13362 4 _0123_
rlabel metal1 s 10396 12954 10396 12954 4 _0124_
rlabel metal1 s 9399 12342 9399 12342 4 _0125_
rlabel metal1 s 5147 14858 5147 14858 4 _0126_
rlabel metal1 s 16702 20366 16702 20366 4 _0127_
rlabel metal1 s 14382 20298 14382 20298 4 _0128_
rlabel metal2 s 16698 18598 16698 18598 4 _0129_
rlabel metal1 s 17536 17102 17536 17102 4 _0130_
rlabel metal2 s 15778 17340 15778 17340 4 _0131_
rlabel metal2 s 16882 14722 16882 14722 4 _0132_
rlabel metal1 s 22325 10506 22325 10506 4 _0133_
rlabel metal1 s 25530 9962 25530 9962 4 _0134_
rlabel metal1 s 22949 11254 22949 11254 4 _0135_
rlabel metal2 s 22126 9690 22126 9690 4 _0136_
rlabel metal1 s 23552 10030 23552 10030 4 _0137_
rlabel metal1 s 24840 8942 24840 8942 4 _0138_
rlabel metal1 s 25668 8058 25668 8058 4 _0139_
rlabel metal1 s 25714 9146 25714 9146 4 _0140_
rlabel metal2 s 25530 10064 25530 10064 4 _0141_
rlabel metal1 s 25790 11594 25790 11594 4 _0142_
rlabel metal1 s 25024 12206 25024 12206 4 _0143_
rlabel metal1 s 26215 14858 26215 14858 4 _0144_
rlabel metal2 s 25801 13838 25801 13838 4 _0145_
rlabel metal1 s 23772 14450 23772 14450 4 _0146_
rlabel metal1 s 25530 13260 25530 13260 4 _0147_
rlabel metal1 s 22724 13294 22724 13294 4 _0148_
rlabel metal1 s 21615 12682 21615 12682 4 _0149_
rlabel metal1 s 20240 21658 20240 21658 4 _0150_
rlabel metal2 s 17434 21250 17434 21250 4 _0151_
rlabel metal1 s 19166 21046 19166 21046 4 _0152_
rlabel metal1 s 20235 19958 20235 19958 4 _0153_
rlabel metal1 s 17296 19482 17296 19482 4 _0154_
rlabel metal1 s 21206 18598 21206 18598 4 _0155_
rlabel metal1 s 17572 18394 17572 18394 4 _0156_
rlabel metal1 s 19361 18122 19361 18122 4 _0157_
rlabel metal1 s 8586 14858 8586 14858 4 _0158_
rlabel metal1 s 13800 25466 13800 25466 4 _0159_
rlabel metal1 s 14669 24242 14669 24242 4 _0160_
rlabel metal1 s 16038 24650 16038 24650 4 _0161_
rlabel metal2 s 15497 22542 15497 22542 4 _0162_
rlabel metal1 s 3716 29070 3716 29070 4 _0163_
rlabel metal2 s 4370 29954 4370 29954 4 _0164_
rlabel metal1 s 3859 27574 3859 27574 4 _0165_
rlabel metal1 s 3542 28186 3542 28186 4 _0166_
rlabel metal2 s 1150 26690 1150 26690 4 _0167_
rlabel metal2 s 3077 25330 3077 25330 4 _0168_
rlabel metal1 s 1104 24922 1104 24922 4 _0169_
rlabel metal2 s 1145 23154 1145 23154 4 _0170_
rlabel metal2 s 966 21250 966 21250 4 _0171_
rlabel metal1 s 2944 20842 2944 20842 4 _0172_
rlabel metal1 s 1104 19482 1104 19482 4 _0173_
rlabel metal1 s 3316 18870 3316 18870 4 _0174_
rlabel metal2 s 1145 17782 1145 17782 4 _0175_
rlabel metal1 s 1191 14858 1191 14858 4 _0176_
rlabel metal2 s 4374 17102 4374 17102 4 _0177_
rlabel metal1 s 2438 16626 2438 16626 4 _0178_
rlabel metal1 s 3864 15130 3864 15130 4 _0179_
rlabel metal2 s 6486 15844 6486 15844 4 _0180_
rlabel metal2 s 6757 13362 6757 13362 4 _0181_
rlabel metal1 s 5796 11866 5796 11866 4 _0182_
rlabel metal2 s 4922 9894 4922 9894 4 _0183_
rlabel metal2 s 6302 10268 6302 10268 4 _0184_
rlabel metal1 s 18768 28186 18768 28186 4 _0185_
rlabel metal1 s 18814 29274 18814 29274 4 _0186_
rlabel metal1 s 19223 30090 19223 30090 4 _0187_
rlabel metal2 s 17613 29682 17613 29682 4 _0188_
rlabel metal1 s 17894 27098 17894 27098 4 _0189_
rlabel metal1 s 18998 27098 18998 27098 4 _0190_
rlabel metal1 s 17878 25398 17878 25398 4 _0191_
rlabel metal1 s 18804 25806 18804 25806 4 _0192_
rlabel metal1 s 18262 14790 18262 14790 4 _0193_
rlabel metal1 s 8142 5338 8142 5338 4 _0194_
rlabel metal1 s 7114 7990 7114 7990 4 _0195_
rlabel metal2 s 5842 8058 5842 8058 4 _0196_
rlabel metal2 s 4278 8058 4278 8058 4 _0197_
rlabel metal1 s 2203 5134 2203 5134 4 _0198_
rlabel metal2 s 1145 7242 1145 7242 4 _0199_
rlabel metal2 s 1150 8806 1150 8806 4 _0200_
rlabel metal1 s 3312 9690 3312 9690 4 _0201_
rlabel metal2 s 3542 16429 3542 16429 4 _0202_
rlabel metal1 s 15548 5338 15548 5338 4 _0203_
rlabel metal1 s 16412 5134 16412 5134 4 _0204_
rlabel metal2 s 16417 7922 16417 7922 4 _0205_
rlabel metal1 s 14030 7514 14030 7514 4 _0206_
rlabel metal1 s 14310 6222 14310 6222 4 _0207_
rlabel metal1 s 11311 6902 11311 6902 4 _0208_
rlabel metal1 s 8970 5338 8970 5338 4 _0209_
rlabel metal1 s 9276 7990 9276 7990 4 _0210_
rlabel metal2 s 3082 21556 3082 21556 4 _0211_
rlabel metal1 s 8050 2618 8050 2618 4 _0212_
rlabel metal2 s 2990 1564 2990 1564 4 _0213_
rlabel metal1 s 2691 2482 2691 2482 4 _0214_
rlabel metal1 s 2507 782 2507 782 4 _0215_
rlabel metal2 s 1242 2108 1242 2108 4 _0216_
rlabel metal1 s 1242 1836 1242 1836 4 _0217_
rlabel metal2 s 8234 1836 8234 1836 4 _0218_
rlabel metal2 s 7038 1904 7038 1904 4 _0219_
rlabel metal1 s 5796 2278 5796 2278 4 _0220_
rlabel metal1 s 5474 3502 5474 3502 4 _0221_
rlabel metal2 s 5244 1870 5244 1870 4 _0222_
rlabel metal1 s 6854 2516 6854 2516 4 _0223_
rlabel metal2 s 4830 1564 4830 1564 4 _0224_
rlabel metal2 s 4554 1258 4554 1258 4 _0225_
rlabel metal2 s 3634 1564 3634 1564 4 _0226_
rlabel metal2 s 6302 5542 6302 5542 4 _0227_
rlabel metal2 s 7590 4454 7590 4454 4 _0228_
rlabel metal2 s 4922 5270 4922 5270 4 _0229_
rlabel metal2 s 5014 4964 5014 4964 4 _0230_
rlabel metal1 s 3496 4046 3496 4046 4 _0231_
rlabel metal2 s 1426 4828 1426 4828 4 _0232_
rlabel metal1 s 1886 4012 1886 4012 4 _0233_
rlabel metal1 s 4876 5338 4876 5338 4 _0234_
rlabel metal1 s 17342 1462 17342 1462 4 _0235_
rlabel metal1 s 11316 1394 11316 1394 4 _0236_
rlabel metal2 s 11270 1530 11270 1530 4 _0237_
rlabel metal2 s 9982 1836 9982 1836 4 _0238_
rlabel metal2 s 9706 1530 9706 1530 4 _0239_
rlabel metal1 s 9568 1870 9568 1870 4 _0240_
rlabel metal1 s 16560 782 16560 782 4 _0241_
rlabel metal2 s 16330 1836 16330 1836 4 _0242_
rlabel metal1 s 15594 2516 15594 2516 4 _0243_
rlabel metal2 s 14306 3332 14306 3332 4 _0244_
rlabel metal2 s 14260 1972 14260 1972 4 _0245_
rlabel metal1 s 13708 1394 13708 1394 4 _0246_
rlabel metal2 s 13018 1564 13018 1564 4 _0247_
rlabel metal1 s 12880 782 12880 782 4 _0248_
rlabel metal2 s 11914 2074 11914 2074 4 _0249_
rlabel metal2 s 12650 4964 12650 4964 4 _0250_
rlabel metal2 s 16514 3876 16514 3876 4 _0251_
rlabel metal1 s 16698 2924 16698 2924 4 _0252_
rlabel metal1 s 14398 4250 14398 4250 4 _0253_
rlabel metal1 s 13570 4794 13570 4794 4 _0254_
rlabel metal2 s 10810 4964 10810 4964 4 _0255_
rlabel metal1 s 12926 3570 12926 3570 4 _0256_
rlabel metal1 s 9706 4012 9706 4012 4 _0257_
rlabel metal1 s 24058 2924 24058 2924 4 _0258_
rlabel metal2 s 19826 2074 19826 2074 4 _0259_
rlabel metal1 s 20010 1428 20010 1428 4 _0260_
rlabel metal2 s 18998 1530 18998 1530 4 _0261_
rlabel metal1 s 18676 1394 18676 1394 4 _0262_
rlabel metal2 s 17710 1530 17710 1530 4 _0263_
rlabel metal1 s 25208 2822 25208 2822 4 _0264_
rlabel metal1 s 24058 2618 24058 2618 4 _0265_
rlabel metal1 s 23322 2346 23322 2346 4 _0266_
rlabel metal1 s 23460 1462 23460 1462 4 _0267_
rlabel metal1 s 22540 782 22540 782 4 _0268_
rlabel metal1 s 22172 2346 22172 2346 4 _0269_
rlabel metal1 s 21482 1836 21482 1836 4 _0270_
rlabel metal2 s 21574 1836 21574 1836 4 _0271_
rlabel metal2 s 20286 1530 20286 1530 4 _0272_
rlabel metal1 s 19504 3910 19504 3910 4 _0273_
rlabel metal1 s 24610 4012 24610 4012 4 _0274_
rlabel metal2 s 24794 3366 24794 3366 4 _0275_
rlabel metal1 s 22034 4760 22034 4760 4 _0276_
rlabel metal2 s 23230 4964 23230 4964 4 _0277_
rlabel metal2 s 19182 4964 19182 4964 4 _0278_
rlabel metal2 s 20746 4386 20746 4386 4 _0279_
rlabel metal2 s 18078 4828 18078 4828 4 _0280_
rlabel metal1 s 24410 27914 24410 27914 4 _0281_
rlabel metal2 s 24334 28390 24334 28390 4 _0282_
rlabel metal1 s 24058 27370 24058 27370 4 _0283_
rlabel metal2 s 24610 27676 24610 27676 4 _0284_
rlabel metal1 s 24978 27370 24978 27370 4 _0285_
rlabel metal1 s 24748 26894 24748 26894 4 _0286_
rlabel metal1 s 24702 27098 24702 27098 4 _0287_
rlabel metal2 s 25622 26588 25622 26588 4 _0288_
rlabel metal2 s 24334 26112 24334 26112 4 _0289_
rlabel metal2 s 24702 26112 24702 26112 4 _0290_
rlabel metal2 s 25070 25534 25070 25534 4 _0291_
rlabel metal1 s 23828 25126 23828 25126 4 _0292_
rlabel metal2 s 23414 25568 23414 25568 4 _0293_
rlabel metal1 s 23828 26010 23828 26010 4 _0294_
rlabel metal1 s 24242 24820 24242 24820 4 _0295_
rlabel metal2 s 23414 24446 23414 24446 4 _0296_
rlabel metal2 s 24518 23494 24518 23494 4 _0297_
rlabel metal2 s 25162 23732 25162 23732 4 _0298_
rlabel metal2 s 24702 24004 24702 24004 4 _0299_
rlabel metal2 s 25806 24310 25806 24310 4 _0300_
rlabel metal1 s 25676 24378 25676 24378 4 _0301_
rlabel metal1 s 26128 24242 26128 24242 4 _0302_
rlabel metal1 s 17066 27574 17066 27574 4 _0303_
rlabel metal1 s 16146 26010 16146 26010 4 _0304_
rlabel metal1 s 16376 26350 16376 26350 4 _0305_
rlabel metal1 s 16054 26486 16054 26486 4 _0306_
rlabel metal2 s 15686 27098 15686 27098 4 _0307_
rlabel metal2 s 14950 27098 14950 27098 4 _0308_
rlabel metal1 s 14536 26758 14536 26758 4 _0309_
rlabel metal2 s 12006 27098 12006 27098 4 _0310_
rlabel metal1 s 10672 28390 10672 28390 4 _0311_
rlabel metal2 s 11454 26656 11454 26656 4 _0312_
rlabel metal2 s 9430 26350 9430 26350 4 _0313_
rlabel metal1 s 9338 26792 9338 26792 4 _0314_
rlabel metal2 s 9154 26894 9154 26894 4 _0315_
rlabel metal1 s 9062 26928 9062 26928 4 _0316_
rlabel metal1 s 9798 26758 9798 26758 4 _0317_
rlabel metal1 s 10718 26894 10718 26894 4 _0318_
rlabel metal1 s 9890 26010 9890 26010 4 _0319_
rlabel metal1 s 10212 26894 10212 26894 4 _0320_
rlabel metal1 s 10810 26418 10810 26418 4 _0321_
rlabel metal2 s 13018 27098 13018 27098 4 _0322_
rlabel metal2 s 11638 26588 11638 26588 4 _0323_
rlabel metal1 s 12328 26486 12328 26486 4 _0324_
rlabel metal2 s 13846 27098 13846 27098 4 _0325_
rlabel metal2 s 12742 26588 12742 26588 4 _0326_
rlabel metal2 s 13018 26588 13018 26588 4 _0327_
rlabel metal1 s 13754 26554 13754 26554 4 _0328_
rlabel metal1 s 17296 26282 17296 26282 4 _0329_
rlabel metal1 s 14996 26826 14996 26826 4 _0330_
rlabel metal2 s 16330 26758 16330 26758 4 _0331_
rlabel metal1 s 16008 13362 16008 13362 4 _0332_
rlabel metal2 s 15686 12886 15686 12886 4 _0333_
rlabel metal1 s 15686 28594 15686 28594 4 _0334_
rlabel metal1 s 13754 28662 13754 28662 4 _0335_
rlabel metal1 s 6394 30736 6394 30736 4 _0336_
rlabel metal1 s 8372 28458 8372 28458 4 _0337_
rlabel metal2 s 8142 28424 8142 28424 4 _0338_
rlabel metal1 s 7314 27982 7314 27982 4 _0339_
rlabel metal1 s 10534 29648 10534 29648 4 _0340_
rlabel metal2 s 8602 29648 8602 29648 4 _0341_
rlabel metal1 s 8648 29206 8648 29206 4 _0342_
rlabel metal1 s 10488 29818 10488 29818 4 _0343_
rlabel metal2 s 10166 30328 10166 30328 4 _0344_
rlabel metal1 s 9338 30158 9338 30158 4 _0345_
rlabel metal1 s 10810 28458 10810 28458 4 _0346_
rlabel metal2 s 10166 28560 10166 28560 4 _0347_
rlabel metal2 s 9982 28628 9982 28628 4 _0348_
rlabel metal1 s 13486 27846 13486 27846 4 _0349_
rlabel metal1 s 11500 28390 11500 28390 4 _0350_
rlabel metal2 s 11822 27948 11822 27948 4 _0351_
rlabel metal1 s 13708 28594 13708 28594 4 _0352_
rlabel metal2 s 13294 28662 13294 28662 4 _0353_
rlabel metal1 s 13616 28730 13616 28730 4 _0354_
rlabel metal1 s 14536 29750 14536 29750 4 _0355_
rlabel metal1 s 14214 28424 14214 28424 4 _0356_
rlabel metal2 s 14306 27948 14306 27948 4 _0357_
rlabel metal1 s 15180 29546 15180 29546 4 _0358_
rlabel metal1 s 14996 29478 14996 29478 4 _0359_
rlabel metal2 s 15410 29988 15410 29988 4 _0360_
rlabel metal1 s 16146 28696 16146 28696 4 _0361_
rlabel metal2 s 15686 29376 15686 29376 4 _0362_
rlabel metal2 s 16146 29988 16146 29988 4 _0363_
rlabel metal2 s 16698 28254 16698 28254 4 _0364_
rlabel metal1 s 16422 28730 16422 28730 4 _0365_
rlabel metal1 s 16882 29036 16882 29036 4 _0366_
rlabel metal1 s 17526 13838 17526 13838 4 _0367_
rlabel metal1 s 18308 15334 18308 15334 4 _0368_
rlabel metal1 s 18492 10098 18492 10098 4 _0369_
rlabel metal1 s 18170 10540 18170 10540 4 _0370_
rlabel metal1 s 18400 13498 18400 13498 4 _0371_
rlabel metal2 s 18998 12070 18998 12070 4 _0372_
rlabel metal2 s 17158 11356 17158 11356 4 _0373_
rlabel metal1 s 18262 13872 18262 13872 4 _0374_
rlabel metal1 s 21482 15436 21482 15436 4 _0375_
rlabel metal2 s 22126 15657 22126 15657 4 _0376_
rlabel metal1 s 21666 15334 21666 15334 4 _0377_
rlabel metal1 s 21574 16048 21574 16048 4 _0378_
rlabel metal1 s 21390 15946 21390 15946 4 _0379_
rlabel metal1 s 22218 16150 22218 16150 4 _0380_
rlabel metal2 s 22402 16796 22402 16796 4 _0381_
rlabel metal1 s 21791 17714 21791 17714 4 _0382_
rlabel metal1 s 21022 18156 21022 18156 4 _0383_
rlabel metal1 s 21160 18054 21160 18054 4 _0384_
rlabel metal2 s 22494 18972 22494 18972 4 _0385_
rlabel metal1 s 21574 19856 21574 19856 4 _0386_
rlabel metal1 s 22770 19142 22770 19142 4 _0387_
rlabel metal1 s 21712 21386 21712 21386 4 _0388_
rlabel metal2 s 21022 21250 21022 21250 4 _0389_
rlabel metal1 s 21620 21114 21620 21114 4 _0390_
rlabel metal1 s 21206 21114 21206 21114 4 _0391_
rlabel metal2 s 22402 20842 22402 20842 4 _0392_
rlabel metal2 s 21666 20196 21666 20196 4 _0393_
rlabel metal1 s 22264 20366 22264 20366 4 _0394_
rlabel metal2 s 22586 20196 22586 20196 4 _0395_
rlabel metal2 s 22770 19754 22770 19754 4 _0396_
rlabel metal2 s 23046 19108 23046 19108 4 _0397_
rlabel metal1 s 21666 18292 21666 18292 4 _0398_
rlabel metal1 s 21620 16626 21620 16626 4 _0399_
rlabel metal2 s 21942 17238 21942 17238 4 _0400_
rlabel metal1 s 21344 17850 21344 17850 4 _0401_
rlabel metal2 s 21482 17714 21482 17714 4 _0402_
rlabel metal2 s 22034 16898 22034 16898 4 _0403_
rlabel metal1 s 22034 17680 22034 17680 4 _0404_
rlabel metal2 s 21482 13056 21482 13056 4 _0405_
rlabel metal2 s 20378 13396 20378 13396 4 _0406_
rlabel metal2 s 21298 13634 21298 13634 4 _0407_
rlabel metal2 s 21022 13668 21022 13668 4 _0408_
rlabel metal1 s 23184 19210 23184 19210 4 _0409_
rlabel metal1 s 23230 21318 23230 21318 4 _0410_
rlabel metal1 s 25346 20978 25346 20978 4 _0411_
rlabel metal1 s 22816 21930 22816 21930 4 _0412_
rlabel metal2 s 23054 22134 23054 22134 4 _0413_
rlabel metal2 s 23230 22372 23230 22372 4 _0414_
rlabel metal2 s 22770 21726 22770 21726 4 _0415_
rlabel metal1 s 22816 21658 22816 21658 4 _0416_
rlabel metal1 s 23414 21658 23414 21658 4 _0417_
rlabel metal2 s 23598 20026 23598 20026 4 _0418_
rlabel metal1 s 23460 20570 23460 20570 4 _0419_
rlabel metal1 s 23874 20366 23874 20366 4 _0420_
rlabel metal1 s 22034 18156 22034 18156 4 _0421_
rlabel metal1 s 23184 19686 23184 19686 4 _0422_
rlabel metal1 s 23966 19924 23966 19924 4 _0423_
rlabel metal1 s 23368 18326 23368 18326 4 _0424_
rlabel metal1 s 22632 18122 22632 18122 4 _0425_
rlabel metal1 s 23690 18190 23690 18190 4 _0426_
rlabel metal1 s 25208 18394 25208 18394 4 _0427_
rlabel metal1 s 24986 18054 24986 18054 4 _0428_
rlabel metal2 s 25530 18598 25530 18598 4 _0429_
rlabel metal1 s 25484 17578 25484 17578 4 _0430_
rlabel metal1 s 25806 17850 25806 17850 4 _0431_
rlabel metal2 s 26450 17612 26450 17612 4 _0432_
rlabel metal1 s 24978 16660 24978 16660 4 _0433_
rlabel metal2 s 25346 16864 25346 16864 4 _0434_
rlabel metal1 s 25714 16626 25714 16626 4 _0435_
rlabel metal1 s 24610 15674 24610 15674 4 _0436_
rlabel metal1 s 24426 15470 24426 15470 4 _0437_
rlabel metal1 s 23644 15674 23644 15674 4 _0438_
rlabel metal1 s 10442 12818 10442 12818 4 _0439_
rlabel metal1 s 10994 13872 10994 13872 4 _0440_
rlabel metal1 s 10672 10234 10672 10234 4 _0441_
rlabel metal2 s 10258 11628 10258 11628 4 _0442_
rlabel metal1 s 9384 12886 9384 12886 4 _0443_
rlabel metal1 s 10396 12750 10396 12750 4 _0444_
rlabel metal1 s 9706 11322 9706 11322 4 _0445_
rlabel metal1 s 10488 15470 10488 15470 4 _0446_
rlabel metal2 s 5106 15028 5106 15028 4 _0447_
rlabel metal2 s 15686 16932 15686 16932 4 _0448_
rlabel metal1 s 15548 16218 15548 16218 4 _0449_
rlabel metal2 s 15134 16388 15134 16388 4 _0450_
rlabel metal1 s 14950 16660 14950 16660 4 _0451_
rlabel metal1 s 14582 18224 14582 18224 4 _0452_
rlabel metal1 s 15042 17782 15042 17782 4 _0453_
rlabel metal1 s 14490 18870 14490 18870 4 _0454_
rlabel metal1 s 14674 19482 14674 19482 4 _0455_
rlabel metal1 s 14950 18190 14950 18190 4 _0456_
rlabel metal1 s 14398 17714 14398 17714 4 _0457_
rlabel metal2 s 14766 17068 14766 17068 4 _0458_
rlabel metal1 s 15594 16422 15594 16422 4 _0459_
rlabel metal2 s 15594 15028 15594 15028 4 _0460_
rlabel metal1 s 15226 20026 15226 20026 4 _0461_
rlabel metal2 s 16238 20230 16238 20230 4 _0462_
rlabel metal1 s 15916 19686 15916 19686 4 _0463_
rlabel metal2 s 15042 20298 15042 20298 4 _0464_
rlabel metal2 s 14858 20196 14858 20196 4 _0465_
rlabel metal1 s 15824 17714 15824 17714 4 _0466_
rlabel metal1 s 16100 18394 16100 18394 4 _0467_
rlabel metal1 s 16422 18190 16422 18190 4 _0468_
rlabel metal1 s 16330 17510 16330 17510 4 _0469_
rlabel metal1 s 16660 16762 16660 16762 4 _0470_
rlabel metal2 s 16974 17238 16974 17238 4 _0471_
rlabel metal1 s 18308 14926 18308 14926 4 _0472_
rlabel metal2 s 21758 14212 21758 14212 4 _0473_
rlabel metal1 s 21758 11560 21758 11560 4 _0474_
rlabel metal1 s 25990 8976 25990 8976 4 _0475_
rlabel metal2 s 24978 15198 24978 15198 4 _0476_
rlabel metal1 s 21988 11594 21988 11594 4 _0477_
rlabel metal2 s 23322 10404 23322 10404 4 _0478_
rlabel metal2 s 26266 8466 26266 8466 4 _0479_
rlabel metal2 s 24518 10812 24518 10812 4 _0480_
rlabel metal1 s 22448 12070 22448 12070 4 _0481_
rlabel metal1 s 22908 8602 22908 8602 4 _0482_
rlabel metal1 s 23184 8058 23184 8058 4 _0483_
rlabel metal1 s 24564 8058 24564 8058 4 _0484_
rlabel metal2 s 26818 7344 26818 7344 4 _0485_
rlabel metal2 s 26174 7922 26174 7922 4 _0486_
rlabel metal2 s 25070 10693 25070 10693 4 _0487_
rlabel metal1 s 25484 10166 25484 10166 4 _0488_
rlabel metal1 s 22954 13362 22954 13362 4 _0489_
rlabel metal1 s 26174 15402 26174 15402 4 _0490_
rlabel metal2 s 26910 14620 26910 14620 4 _0491_
rlabel metal1 s 23322 14382 23322 14382 4 _0492_
rlabel metal1 s 23552 13226 23552 13226 4 _0493_
rlabel metal1 s 23276 13362 23276 13362 4 _0494_
rlabel metal1 s 22034 12274 22034 12274 4 _0495_
rlabel metal1 s 21850 12104 21850 12104 4 _0496_
rlabel metal1 s 24334 9418 24334 9418 4 _0497_
rlabel metal1 s 22724 9350 22724 9350 4 _0498_
rlabel metal1 s 21942 12342 21942 12342 4 _0499_
rlabel metal1 s 22586 12410 22586 12410 4 _0500_
rlabel metal2 s 21850 12308 21850 12308 4 _0501_
rlabel metal1 s 21344 20366 21344 20366 4 _0502_
rlabel metal1 s 21482 20298 21482 20298 4 _0503_
rlabel metal1 s 7314 14450 7314 14450 4 _0504_
rlabel metal1 s 7176 14382 7176 14382 4 _0505_
rlabel metal2 s 7038 15674 7038 15674 4 _0506_
rlabel metal1 s 10258 16694 10258 16694 4 _0507_
rlabel metal1 s 9154 15606 9154 15606 4 _0508_
rlabel metal2 s 8786 14858 8786 14858 4 _0509_
rlabel metal2 s 9246 14892 9246 14892 4 _0510_
rlabel metal1 s 8602 15538 8602 15538 4 _0511_
rlabel metal1 s 14950 25466 14950 25466 4 _0512_
rlabel metal1 s 15226 23732 15226 23732 4 _0513_
rlabel metal1 s 14260 25330 14260 25330 4 _0514_
rlabel metal2 s 15134 24140 15134 24140 4 _0515_
rlabel metal2 s 14674 24276 14674 24276 4 _0516_
rlabel metal1 s 17020 24378 17020 24378 4 _0517_
rlabel metal1 s 15916 24378 15916 24378 4 _0518_
rlabel metal1 s 16284 23086 16284 23086 4 _0519_
rlabel metal1 s 15502 23086 15502 23086 4 _0520_
rlabel metal2 s 6302 17680 6302 17680 4 _0521_
rlabel metal2 s 5658 17306 5658 17306 4 _0522_
rlabel metal2 s 5474 16864 5474 16864 4 _0523_
rlabel metal1 s 4968 16762 4968 16762 4 _0524_
rlabel metal1 s 5198 18054 5198 18054 4 _0525_
rlabel metal1 s 6210 18122 6210 18122 4 _0526_
rlabel metal1 s 5474 17748 5474 17748 4 _0527_
rlabel metal1 s 5106 17306 5106 17306 4 _0528_
rlabel metal1 s 5152 18122 5152 18122 4 _0529_
rlabel metal2 s 6118 18598 6118 18598 4 _0530_
rlabel metal1 s 5474 18598 5474 18598 4 _0531_
rlabel metal1 s 5980 18938 5980 18938 4 _0532_
rlabel metal1 s 2346 19244 2346 19244 4 _0533_
rlabel metal1 s 3542 19890 3542 19890 4 _0534_
rlabel metal1 s 4324 20026 4324 20026 4 _0535_
rlabel metal2 s 4186 21148 4186 21148 4 _0536_
rlabel metal1 s 4324 20366 4324 20366 4 _0537_
rlabel metal1 s 2622 20332 2622 20332 4 _0538_
rlabel metal2 s 5474 21420 5474 21420 4 _0539_
rlabel metal2 s 4922 21080 4922 21080 4 _0540_
rlabel metal2 s 4738 20604 4738 20604 4 _0541_
rlabel metal1 s 4692 19822 4692 19822 4 _0542_
rlabel metal1 s 4508 17850 4508 17850 4 _0543_
rlabel metal1 s 5060 19890 5060 19890 4 _0544_
rlabel metal2 s 5658 19516 5658 19516 4 _0545_
rlabel metal2 s 5106 25126 5106 25126 4 _0546_
rlabel metal2 s 5658 27268 5658 27268 4 _0547_
rlabel metal1 s 6256 27506 6256 27506 4 _0548_
rlabel metal2 s 5934 27676 5934 27676 4 _0549_
rlabel metal2 s 5842 26860 5842 26860 4 _0550_
rlabel metal1 s 5336 24922 5336 24922 4 _0551_
rlabel metal2 s 4646 25670 4646 25670 4 _0552_
rlabel metal1 s 5428 26418 5428 26418 4 _0553_
rlabel metal2 s 5014 26044 5014 26044 4 _0554_
rlabel metal2 s 4462 25636 4462 25636 4 _0555_
rlabel metal2 s 4370 25024 4370 25024 4 _0556_
rlabel metal2 s 4048 23630 4048 23630 4 _0557_
rlabel metal1 s 4186 23120 4186 23120 4 _0558_
rlabel metal1 s 3864 23086 3864 23086 4 _0559_
rlabel metal1 s 4600 23290 4600 23290 4 _0560_
rlabel metal1 s 4554 23630 4554 23630 4 _0561_
rlabel metal1 s 4968 23834 4968 23834 4 _0562_
rlabel metal1 s 1334 23664 1334 23664 4 _0563_
rlabel metal1 s 2346 25874 2346 25874 4 _0564_
rlabel metal3 s 3818 23613 3818 23613 4 _0565_
rlabel metal1 s 5290 23834 5290 23834 4 _0566_
rlabel metal1 s 4462 22406 4462 22406 4 _0567_
rlabel metal2 s 4830 23324 4830 23324 4 _0568_
rlabel metal2 s 4554 22746 4554 22746 4 _0569_
rlabel metal1 s 4508 20570 4508 20570 4 _0570_
rlabel metal1 s 4554 20502 4554 20502 4 _0571_
rlabel metal2 s 4830 21556 4830 21556 4 _0572_
rlabel metal1 s 5060 22542 5060 22542 4 _0573_
rlabel metal2 s 5796 21114 5796 21114 4 _0574_
rlabel metal1 s 5244 19278 5244 19278 4 _0575_
rlabel metal1 s 5474 22508 5474 22508 4 _0576_
rlabel metal1 s 4784 19278 4784 19278 4 _0577_
rlabel metal1 s 4600 16014 4600 16014 4 _0578_
rlabel metal1 s 1978 19482 1978 19482 4 _0579_
rlabel metal1 s 2346 16694 2346 16694 4 _0580_
rlabel metal2 s 5842 29172 5842 29172 4 _0581_
rlabel metal1 s 5152 28390 5152 28390 4 _0582_
rlabel metal1 s 4822 28730 4822 28730 4 _0583_
rlabel metal1 s 4324 28730 4324 28730 4 _0584_
rlabel metal1 s 2622 26452 2622 26452 4 _0585_
rlabel metal1 s 4278 27030 4278 27030 4 _0586_
rlabel metal2 s 4186 27540 4186 27540 4 _0587_
rlabel metal1 s 3082 27302 3082 27302 4 _0588_
rlabel metal2 s 2714 27574 2714 27574 4 _0589_
rlabel metal1 s 3082 27642 3082 27642 4 _0590_
rlabel metal1 s 2392 26282 2392 26282 4 _0591_
rlabel metal2 s 2806 26826 2806 26826 4 _0592_
rlabel metal1 s 1840 26418 1840 26418 4 _0593_
rlabel metal1 s 2530 25772 2530 25772 4 _0594_
rlabel metal1 s 2684 24650 2684 24650 4 _0595_
rlabel metal1 s 2852 24922 2852 24922 4 _0596_
rlabel metal1 s 2392 24038 2392 24038 4 _0597_
rlabel metal2 s 1886 23800 1886 23800 4 _0598_
rlabel metal2 s 1878 24650 1878 24650 4 _0599_
rlabel metal1 s 1472 24718 1472 24718 4 _0600_
rlabel metal1 s 2116 22066 2116 22066 4 _0601_
rlabel metal1 s 1426 23834 1426 23834 4 _0602_
rlabel metal1 s 874 23698 874 23698 4 _0603_
rlabel metal2 s 2438 20570 2438 20570 4 _0604_
rlabel metal2 s 1418 21114 1418 21114 4 _0605_
rlabel metal1 s 1196 20978 1196 20978 4 _0606_
rlabel metal1 s 2392 22746 2392 22746 4 _0607_
rlabel metal1 s 2208 21590 2208 21590 4 _0608_
rlabel metal1 s 2622 20570 2622 20570 4 _0609_
rlabel metal2 s 2898 21148 2898 21148 4 _0610_
rlabel metal2 s 2346 20298 2346 20298 4 _0611_
rlabel metal1 s 2016 20230 2016 20230 4 _0612_
rlabel metal2 s 1242 19754 1242 19754 4 _0613_
rlabel metal1 s 2392 19414 2392 19414 4 _0614_
rlabel metal1 s 2208 19142 2208 19142 4 _0615_
rlabel metal2 s 2806 19686 2806 19686 4 _0616_
rlabel metal2 s 1886 17646 1886 17646 4 _0617_
rlabel metal1 s 1748 17034 1748 17034 4 _0618_
rlabel metal2 s 1334 17748 1334 17748 4 _0619_
rlabel metal1 s 1748 16218 1748 16218 4 _0620_
rlabel metal1 s 2246 15878 2246 15878 4 _0621_
rlabel metal1 s 1472 15538 1472 15538 4 _0622_
rlabel metal1 s 2484 17238 2484 17238 4 _0623_
rlabel metal2 s 2898 17272 2898 17272 4 _0624_
rlabel metal2 s 3082 17510 3082 17510 4 _0625_
rlabel metal2 s 7774 15130 7774 15130 4 _0626_
rlabel metal1 s 6670 15572 6670 15572 4 _0627_
rlabel metal2 s 6302 13804 6302 13804 4 _0628_
rlabel metal1 s 6808 12954 6808 12954 4 _0629_
rlabel metal1 s 6348 13498 6348 13498 4 _0630_
rlabel metal1 s 6256 11526 6256 11526 4 _0631_
rlabel metal2 s 6762 11492 6762 11492 4 _0632_
rlabel metal1 s 5796 10778 5796 10778 4 _0633_
rlabel metal2 s 6670 10404 6670 10404 4 _0634_
rlabel metal2 s 5106 9962 5106 9962 4 _0635_
rlabel metal1 s 5934 10642 5934 10642 4 _0636_
rlabel metal1 s 18032 24718 18032 24718 4 _0637_
rlabel metal1 s 17894 30872 17894 30872 4 _0638_
rlabel metal1 s 7636 6426 7636 6426 4 _0639_
rlabel metal2 s 7782 6086 7782 6086 4 _0640_
rlabel metal1 s 7912 5134 7912 5134 4 _0641_
rlabel metal1 s 7590 7276 7590 7276 4 _0642_
rlabel metal1 s 7820 7378 7820 7378 4 _0643_
rlabel metal1 s 6578 6868 6578 6868 4 _0644_
rlabel metal1 s 6992 7514 6992 7514 4 _0645_
rlabel metal1 s 6900 7786 6900 7786 4 _0646_
rlabel metal2 s 6486 7072 6486 7072 4 _0647_
rlabel metal1 s 6302 6800 6302 6800 4 _0648_
rlabel metal1 s 6210 6902 6210 6902 4 _0649_
rlabel metal1 s 5888 7378 5888 7378 4 _0650_
rlabel metal1 s 5980 6970 5980 6970 4 _0651_
rlabel metal1 s 6072 7514 6072 7514 4 _0652_
rlabel metal1 s 5106 6766 5106 6766 4 _0653_
rlabel metal2 s 4646 6596 4646 6596 4 _0654_
rlabel metal1 s 4968 7310 4968 7310 4 _0655_
rlabel metal1 s 4416 7446 4416 7446 4 _0656_
rlabel metal1 s 4416 6834 4416 6834 4 _0657_
rlabel metal2 s 4462 7718 4462 7718 4 _0658_
rlabel metal1 s 3496 6222 3496 6222 4 _0659_
rlabel metal1 s 2990 4692 2990 4692 4 _0660_
rlabel metal2 s 3174 5100 3174 5100 4 _0661_
rlabel metal1 s 3036 6222 3036 6222 4 _0662_
rlabel metal1 s 3450 6426 3450 6426 4 _0663_
rlabel metal2 s 3634 7072 3634 7072 4 _0664_
rlabel metal1 s 2622 5780 2622 5780 4 _0665_
rlabel metal1 s 2392 7514 2392 7514 4 _0666_
rlabel metal1 s 2576 7310 2576 7310 4 _0667_
rlabel metal1 s 3220 7378 3220 7378 4 _0668_
rlabel metal1 s 3266 6698 3266 6698 4 _0669_
rlabel metal1 s 2530 7888 2530 7888 4 _0670_
rlabel metal1 s 2668 6766 2668 6766 4 _0671_
rlabel metal2 s 2990 9146 2990 9146 4 _0672_
rlabel metal2 s 3175 9010 3175 9010 4 _0673_
rlabel metal2 s 3082 8602 3082 8602 4 _0674_
rlabel metal1 s 2392 8602 2392 8602 4 _0675_
rlabel metal2 s 2706 9078 2706 9078 4 _0676_
rlabel metal1 s 1334 8432 1334 8432 4 _0677_
rlabel metal1 s 3680 10438 3680 10438 4 _0678_
rlabel metal1 s 4232 9486 4232 9486 4 _0679_
rlabel metal1 s 2622 10030 2622 10030 4 _0680_
rlabel metal1 s 2668 9554 2668 9554 4 _0681_
rlabel metal1 s 3128 10574 3128 10574 4 _0682_
rlabel metal1 s 3266 9486 3266 9486 4 _0683_
rlabel metal1 s 15272 5338 15272 5338 4 _0684_
rlabel metal2 s 15594 5644 15594 5644 4 _0685_
rlabel metal1 s 15640 5134 15640 5134 4 _0686_
rlabel metal1 s 17848 5542 17848 5542 4 _0687_
rlabel metal1 s 17066 5814 17066 5814 4 _0688_
rlabel metal2 s 16606 5882 16606 5882 4 _0689_
rlabel metal2 s 16514 5984 16514 5984 4 _0690_
rlabel metal1 s 16146 5746 16146 5746 4 _0691_
rlabel metal2 s 16974 7072 16974 7072 4 _0692_
rlabel metal1 s 16790 6800 16790 6800 4 _0693_
rlabel metal1 s 17342 7412 17342 7412 4 _0694_
rlabel metal1 s 16284 7446 16284 7446 4 _0695_
rlabel metal1 s 16376 6970 16376 6970 4 _0696_
rlabel metal1 s 16468 7514 16468 7514 4 _0697_
rlabel metal2 s 15318 8160 15318 8160 4 _0698_
rlabel metal2 s 15134 8228 15134 8228 4 _0699_
rlabel metal2 s 15686 7718 15686 7718 4 _0700_
rlabel metal1 s 14536 7514 14536 7514 4 _0701_
rlabel metal1 s 13294 7956 13294 7956 4 _0702_
rlabel metal1 s 14352 7310 14352 7310 4 _0703_
rlabel metal2 s 14214 6358 14214 6358 4 _0704_
rlabel metal1 s 13570 6800 13570 6800 4 _0705_
rlabel metal2 s 13386 7412 13386 7412 4 _0706_
rlabel metal2 s 14030 7548 14030 7548 4 _0707_
rlabel metal1 s 12650 7412 12650 7412 4 _0708_
rlabel metal2 s 13110 7004 13110 7004 4 _0709_
rlabel metal2 s 12558 6630 12558 6630 4 _0710_
rlabel metal2 s 11546 6630 11546 6630 4 _0711_
rlabel metal2 s 12558 7140 12558 7140 4 _0712_
rlabel metal2 s 12098 7514 12098 7514 4 _0713_
rlabel metal1 s 11822 7344 11822 7344 4 _0714_
rlabel metal2 s 10074 6052 10074 6052 4 _0715_
rlabel metal1 s 10442 6222 10442 6222 4 _0716_
rlabel metal1 s 10626 6290 10626 6290 4 _0717_
rlabel metal1 s 9292 6426 9292 6426 4 _0718_
rlabel metal1 s 9676 6154 9676 6154 4 _0719_
rlabel metal2 s 9246 5746 9246 5746 4 _0720_
rlabel metal1 s 10304 8806 10304 8806 4 _0721_
rlabel metal1 s 11040 7310 11040 7310 4 _0722_
rlabel metal1 s 10166 7308 10166 7308 4 _0723_
rlabel metal1 s 9246 7514 9246 7514 4 _0724_
rlabel metal1 s 9660 8398 9660 8398 4 _0725_
rlabel metal1 s 8556 7922 8556 7922 4 _0726_
rlabel metal1 s 8556 14450 8556 14450 4 _0727_
rlabel metal1 s 12926 9452 12926 9452 4 _0728_
rlabel metal2 s 19642 11390 19642 11390 4 _0729_
rlabel metal1 s 13018 11016 13018 11016 4 _0730_
rlabel metal2 s 8970 10268 8970 10268 4 _0731_
rlabel metal1 s 6670 4760 6670 4760 4 _0732_
rlabel metal1 s 13570 9656 13570 9656 4 _0733_
rlabel metal2 s 9062 9452 9062 9452 4 _0734_
rlabel metal1 s 7130 5202 7130 5202 4 _0735_
rlabel metal1 s 6992 4658 6992 4658 4 _0736_
rlabel metal1 s 3542 2448 3542 2448 4 _0737_
rlabel metal1 s 12742 8908 12742 8908 4 _0738_
rlabel metal1 s 9062 9452 9062 9452 4 _0739_
rlabel metal1 s 6946 5100 6946 5100 4 _0740_
rlabel metal1 s 15594 10642 15594 10642 4 _0741_
rlabel metal2 s 9246 10846 9246 10846 4 _0742_
rlabel metal1 s 8832 10438 8832 10438 4 _0743_
rlabel metal1 s 7130 2482 7130 2482 4 _0744_
rlabel metal1 s 6302 5202 6302 5202 4 _0745_
rlabel metal1 s 6900 5202 6900 5202 4 _0746_
rlabel metal2 s 9016 4046 9016 4046 4 _0747_
rlabel metal1 s 7774 4080 7774 4080 4 _0748_
rlabel metal1 s 7820 3706 7820 3706 4 _0749_
rlabel metal1 s 7912 2482 7912 2482 4 _0750_
rlabel metal1 s 4554 2516 4554 2516 4 _0751_
rlabel metal1 s 8004 3910 8004 3910 4 _0752_
rlabel metal1 s 4370 1836 4370 1836 4 _0753_
rlabel metal1 s 3864 3638 3864 3638 4 _0754_
rlabel metal1 s 4876 2618 4876 2618 4 _0755_
rlabel metal1 s 5382 2482 5382 2482 4 _0756_
rlabel metal1 s 5658 2448 5658 2448 4 _0757_
rlabel metal1 s 4094 2992 4094 2992 4 _0758_
rlabel metal1 s 4600 3162 4600 3162 4 _0759_
rlabel metal1 s 4508 3570 4508 3570 4 _0760_
rlabel metal1 s 5106 3706 5106 3706 4 _0761_
rlabel metal1 s 6900 3502 6900 3502 4 _0762_
rlabel metal1 s 6486 3672 6486 3672 4 _0763_
rlabel metal1 s 1610 5100 1610 5100 4 _0764_
rlabel metal2 s 17894 10778 17894 10778 4 _0765_
rlabel metal1 s 13018 8976 13018 8976 4 _0766_
rlabel metal2 s 13294 9690 13294 9690 4 _0767_
rlabel metal1 s 12420 5066 12420 5066 4 _0768_
rlabel metal1 s 13156 12614 13156 12614 4 _0769_
rlabel metal1 s 11960 5134 11960 5134 4 _0770_
rlabel metal2 s 12742 4862 12742 4862 4 _0771_
rlabel metal1 s 12650 4080 12650 4080 4 _0772_
rlabel metal1 s 13018 8602 13018 8602 4 _0773_
rlabel metal2 s 12466 7089 12466 7089 4 _0774_
rlabel metal1 s 12518 10574 12518 10574 4 _0775_
rlabel metal1 s 12650 3468 12650 3468 4 _0776_
rlabel metal2 s 13570 3009 13570 3009 4 _0777_
rlabel metal1 s 11592 4522 11592 4522 4 _0778_
rlabel metal1 s 11592 4182 11592 4182 4 _0779_
rlabel metal1 s 11592 4590 11592 4590 4 _0780_
rlabel metal1 s 13294 1904 13294 1904 4 _0781_
rlabel metal1 s 15364 3162 15364 3162 4 _0782_
rlabel metal2 s 12834 3876 12834 3876 4 _0783_
rlabel metal1 s 14628 4182 14628 4182 4 _0784_
rlabel metal1 s 15778 4046 15778 4046 4 _0785_
rlabel metal2 s 16330 3740 16330 3740 4 _0786_
rlabel metal2 s 12834 3162 12834 3162 4 _0787_
rlabel metal1 s 13018 1836 13018 1836 4 _0788_
rlabel metal1 s 15686 2380 15686 2380 4 _0789_
rlabel metal1 s 16054 2822 16054 2822 4 _0790_
rlabel metal1 s 13938 2550 13938 2550 4 _0791_
rlabel metal1 s 13754 2924 13754 2924 4 _0792_
rlabel metal1 s 16054 2958 16054 2958 4 _0793_
rlabel metal1 s 13202 2924 13202 2924 4 _0794_
rlabel metal1 s 13156 3162 13156 3162 4 _0795_
rlabel metal1 s 14076 3706 14076 3706 4 _0796_
rlabel metal1 s 13570 4046 13570 4046 4 _0797_
rlabel metal1 s 13432 4250 13432 4250 4 _0798_
rlabel metal2 s 11086 4386 11086 4386 4 _0799_
rlabel metal1 s 16376 2482 16376 2482 4 _0800_
rlabel metal1 s 18262 12682 18262 12682 4 _0801_
rlabel metal1 s 16652 12614 16652 12614 4 _0802_
rlabel metal1 s 16146 9452 16146 9452 4 _0803_
rlabel metal1 s 23092 2618 23092 2618 4 _0804_
rlabel metal1 s 15548 10098 15548 10098 4 _0805_
rlabel metal1 s 16790 3978 16790 3978 4 _0806_
rlabel metal2 s 17894 3774 17894 3774 4 _0807_
rlabel metal1 s 18906 2448 18906 2448 4 _0808_
rlabel metal2 s 15962 9180 15962 9180 4 _0809_
rlabel metal1 s 17204 2958 17204 2958 4 _0810_
rlabel metal2 s 16238 10336 16238 10336 4 _0811_
rlabel metal1 s 17986 5168 17986 5168 4 _0812_
rlabel metal1 s 17710 2516 17710 2516 4 _0813_
rlabel metal1 s 18584 4182 18584 4182 4 _0814_
rlabel metal1 s 18354 3434 18354 3434 4 _0815_
rlabel metal1 s 19592 4114 19592 4114 4 _0816_
rlabel metal1 s 20516 2482 20516 2482 4 _0817_
rlabel metal1 s 23368 2958 23368 2958 4 _0818_
rlabel metal1 s 20838 4012 20838 4012 4 _0819_
rlabel metal1 s 23276 3910 23276 3910 4 _0820_
rlabel metal1 s 23782 2958 23782 2958 4 _0821_
rlabel metal1 s 24104 3162 24104 3162 4 _0822_
rlabel metal1 s 20332 3094 20332 3094 4 _0823_
rlabel metal1 s 20792 2482 20792 2482 4 _0824_
rlabel metal1 s 23138 3128 23138 3128 4 _0825_
rlabel metal1 s 23414 2482 23414 2482 4 _0826_
rlabel metal1 s 22264 2482 22264 2482 4 _0827_
rlabel metal1 s 22310 2992 22310 2992 4 _0828_
rlabel metal1 s 24840 2958 24840 2958 4 _0829_
rlabel metal1 s 19136 2618 19136 2618 4 _0830_
rlabel metal1 s 21114 3638 21114 3638 4 _0831_
rlabel metal2 s 21850 4182 21850 4182 4 _0832_
rlabel metal1 s 21988 4114 21988 4114 4 _0833_
rlabel metal1 s 23000 4250 23000 4250 4 _0834_
rlabel metal1 s 18768 4250 18768 4250 4 _0835_
rlabel metal2 s 25070 3162 25070 3162 4 _0836_
rlabel metal1 s 12420 22610 12420 22610 4 _0837_
rlabel metal1 s 12328 20978 12328 20978 4 _0838_
rlabel metal2 s 12466 20366 12466 20366 4 _0839_
rlabel metal1 s 16882 21862 16882 21862 4 _0840_
rlabel metal2 s 21850 17459 21850 17459 4 _0841_
rlabel metal1 s 16146 21318 16146 21318 4 _0842_
rlabel metal1 s 20194 24242 20194 24242 4 _0843_
rlabel metal2 s 12834 23018 12834 23018 4 _0844_
rlabel metal1 s 20148 22610 20148 22610 4 _0845_
rlabel metal1 s 19320 24378 19320 24378 4 _0846_
rlabel metal1 s 20148 22474 20148 22474 4 _0847_
rlabel metal2 s 19642 22950 19642 22950 4 _0848_
rlabel metal2 s 18906 23664 18906 23664 4 _0849_
rlabel metal1 s 18400 23290 18400 23290 4 _0850_
rlabel metal1 s 17572 23290 17572 23290 4 _0851_
rlabel metal1 s 16974 23290 16974 23290 4 _0852_
rlabel metal1 s 17664 21318 17664 21318 4 _0853_
rlabel metal1 s 14214 16728 14214 16728 4 _0854_
rlabel metal2 s 9522 22073 9522 22073 4 _0855_
rlabel metal1 s 12834 25160 12834 25160 4 _0856_
rlabel metal1 s 8058 25738 8058 25738 4 _0857_
rlabel metal1 s 9798 21964 9798 21964 4 _0858_
rlabel metal1 s 17480 18054 17480 18054 4 _0859_
rlabel metal1 s 8924 26418 8924 26418 4 _0860_
rlabel metal1 s 18538 18394 18538 18394 4 _0861_
rlabel metal1 s 9476 24242 9476 24242 4 _0862_
rlabel metal2 s 21298 20315 21298 20315 4 _0863_
rlabel metal2 s 10166 23596 10166 23596 4 _0864_
rlabel metal3 s 17250 19227 17250 19227 4 _0865_
rlabel metal2 s 9706 25772 9706 25772 4 _0866_
rlabel metal1 s 12374 25466 12374 25466 4 _0867_
rlabel metal1 s 12972 19686 12972 19686 4 _0868_
rlabel metal1 s 11960 23154 11960 23154 4 _0869_
rlabel metal1 s 12834 24276 12834 24276 4 _0870_
rlabel metal1 s 16836 20978 16836 20978 4 _0871_
rlabel metal1 s 12926 18802 12926 18802 4 _0872_
rlabel metal1 s 12780 19958 12780 19958 4 _0873_
rlabel metal2 s 13386 18972 13386 18972 4 _0874_
rlabel metal2 s 12466 19244 12466 19244 4 _0875_
rlabel metal1 s 12834 17136 12834 17136 4 _0876_
rlabel metal2 s 12650 15980 12650 15980 4 _0877_
rlabel metal1 s 13340 15538 13340 15538 4 _0878_
rlabel metal1 s 17802 17680 17802 17680 4 _0879_
rlabel metal1 s 2254 9996 2254 9996 4 _0880_
rlabel metal3 s 1702 15555 1702 15555 4 _0881_
rlabel metal1 s 18860 17782 18860 17782 4 _0882_
rlabel metal1 s 14996 14858 14996 14858 4 _0883_
rlabel metal1 s 13018 20944 13018 20944 4 _0884_
rlabel metal1 s 21804 5542 21804 5542 4 _0885_
rlabel metal2 s 21850 5610 21850 5610 4 _0886_
rlabel metal1 s 21206 5746 21206 5746 4 _0887_
rlabel metal2 s 24610 4964 24610 4964 4 _0888_
rlabel metal1 s 25162 5712 25162 5712 4 _0889_
rlabel metal1 s 24840 5542 24840 5542 4 _0890_
rlabel metal1 s 21068 14042 21068 14042 4 _0891_
rlabel metal2 s 24426 4896 24426 4896 4 _0892_
rlabel metal1 s 24932 4522 24932 4522 4 _0893_
rlabel metal2 s 25254 6358 25254 6358 4 _0894_
rlabel metal2 s 25438 6630 25438 6630 4 _0895_
rlabel metal1 s 25024 6834 25024 6834 4 _0896_
rlabel metal2 s 23598 7072 23598 7072 4 _0897_
rlabel metal1 s 25070 6154 25070 6154 4 _0898_
rlabel metal2 s 24610 6868 24610 6868 4 _0899_
rlabel metal2 s 23322 6630 23322 6630 4 _0900_
rlabel metal1 s 21758 7276 21758 7276 4 _0901_
rlabel metal2 s 23782 7038 23782 7038 4 _0902_
rlabel metal1 s 21574 6664 21574 6664 4 _0903_
rlabel metal2 s 22034 7106 22034 7106 4 _0904_
rlabel metal1 s 21574 6222 21574 6222 4 _0905_
rlabel metal1 s 23782 7956 23782 7956 4 _0906_
rlabel metal1 s 21482 8432 21482 8432 4 _0907_
rlabel metal2 s 21942 7548 21942 7548 4 _0908_
rlabel metal1 s 21620 8398 21620 8398 4 _0909_
rlabel metal1 s 17710 20332 17710 20332 4 _0910_
rlabel metal2 s 21758 7956 21758 7956 4 _0911_
rlabel metal1 s 20286 8432 20286 8432 4 _0912_
rlabel metal1 s 20470 8942 20470 8942 4 _0913_
rlabel metal1 s 21252 7922 21252 7922 4 _0914_
rlabel metal2 s 20838 8636 20838 8636 4 _0915_
rlabel metal1 s 20608 8398 20608 8398 4 _0916_
rlabel metal2 s 20470 8806 20470 8806 4 _0917_
rlabel metal1 s 19550 7446 19550 7446 4 _0918_
rlabel metal2 s 19734 7140 19734 7140 4 _0919_
rlabel metal1 s 19826 7888 19826 7888 4 _0920_
rlabel metal2 s 18906 7616 18906 7616 4 _0921_
rlabel metal1 s 19220 7174 19220 7174 4 _0922_
rlabel metal1 s 17940 6834 17940 6834 4 _0923_
rlabel metal1 s 19435 9010 19435 9010 4 _0924_
rlabel metal2 s 19550 9044 19550 9044 4 _0925_
rlabel metal2 s 18814 8602 18814 8602 4 _0926_
rlabel metal1 s 18492 8058 18492 8058 4 _0927_
rlabel metal1 s 18676 8534 18676 8534 4 _0928_
rlabel metal1 s 17802 8398 17802 8398 4 _0929_
rlabel metal1 s 12144 30770 12144 30770 4 _0930_
rlabel metal1 s 14306 30736 14306 30736 4 _0931_
rlabel metal1 s 14306 21522 14306 21522 4 _0932_
rlabel metal2 s 13202 22746 13202 22746 4 _0933_
rlabel metal1 s 13846 22746 13846 22746 4 _0934_
rlabel metal2 s 13110 21148 13110 21148 4 _0935_
rlabel metal2 s 13570 20570 13570 20570 4 _0936_
rlabel metal1 s 10672 22406 10672 22406 4 _0937_
rlabel metal1 s 10810 22066 10810 22066 4 _0938_
rlabel metal1 s 10350 20944 10350 20944 4 _0939_
rlabel metal1 s 10672 20978 10672 20978 4 _0940_
rlabel metal2 s 11730 29818 11730 29818 4 _0941_
rlabel metal2 s 1610 13498 1610 13498 4 _0942_
rlabel metal2 s 3442 11526 3442 11526 4 _0943_
rlabel metal1 s 2852 13430 2852 13430 4 _0944_
rlabel metal1 s 3542 13328 3542 13328 4 _0945_
rlabel metal1 s 1656 11186 1656 11186 4 _0946_
rlabel metal1 s 5152 13838 5152 13838 4 _0947_
rlabel metal1 s 2944 11322 2944 11322 4 _0948_
rlabel metal1 s 2622 11050 2622 11050 4 _0949_
rlabel metal2 s 3910 13532 3910 13532 4 _0950_
rlabel metal1 s 15870 12954 15870 12954 4 _0951_
rlabel metal1 s 6670 12614 6670 12614 4 _0952_
rlabel metal1 s 4232 12614 4232 12614 4 _0953_
rlabel metal2 s 11454 19346 11454 19346 4 _0954_
rlabel metal2 s 11730 19244 11730 19244 4 _0955_
rlabel metal1 s 11914 17850 11914 17850 4 _0956_
rlabel metal2 s 11178 17918 11178 17918 4 _0957_
rlabel metal2 s 10350 16150 10350 16150 4 _0958_
rlabel metal2 s 10258 17238 10258 17238 4 _0959_
rlabel metal1 s 9522 17714 9522 17714 4 _0960_
rlabel metal1 s 11546 15674 11546 15674 4 _0961_
rlabel metal1 s 10258 16014 10258 16014 4 _0962_
rlabel metal1 s 16054 22066 16054 22066 4 _0963_
rlabel metal1 s 9522 19856 9522 19856 4 _0964_
rlabel metal2 s 7498 20842 7498 20842 4 _0965_
rlabel metal1 s 8758 21012 8758 21012 4 _0966_
rlabel metal1 s 5566 21488 5566 21488 4 _0967_
rlabel metal1 s 8096 20366 8096 20366 4 _0968_
rlabel metal2 s 8878 20332 8878 20332 4 _0969_
rlabel metal1 s 6992 19278 6992 19278 4 _0970_
rlabel metal2 s 7866 17102 7866 17102 4 _0971_
rlabel metal2 s 6486 17306 6486 17306 4 _0972_
rlabel metal1 s 7590 18190 7590 18190 4 _0973_
rlabel metal1 s 8878 18190 8878 18190 4 _0974_
rlabel metal1 s 12558 14892 12558 14892 4 _0975_
rlabel metal1 s 15180 13838 15180 13838 4 _0976_
rlabel metal1 s 15134 13770 15134 13770 4 _0977_
rlabel metal1 s 14628 13498 14628 13498 4 _0978_
rlabel metal1 s 14122 9044 14122 9044 4 _0979_
rlabel metal1 s 13846 10540 13846 10540 4 _0980_
rlabel metal1 s 14950 13872 14950 13872 4 _0981_
rlabel metal1 s 14260 13158 14260 13158 4 _0982_
rlabel metal2 s 15594 11356 15594 11356 4 _0983_
rlabel metal1 s 17250 15538 17250 15538 4 _0984_
rlabel metal2 s 13018 22814 13018 22814 4 _0985_
rlabel metal1 s 6854 23120 6854 23120 4 _0986_
rlabel metal1 s 11914 9486 11914 9486 4 _0987_
rlabel metal1 s 12926 14824 12926 14824 4 _0988_
rlabel metal2 s 11730 9044 11730 9044 4 _0989_
rlabel metal1 s 11730 10064 11730 10064 4 _0990_
rlabel metal1 s 19458 13770 19458 13770 4 _0991_
rlabel metal1 s 12581 13974 12581 13974 4 _0992_
rlabel metal2 s 11730 12444 11730 12444 4 _0993_
rlabel metal1 s 12742 11560 12742 11560 4 _0994_
rlabel metal2 s 20930 26010 20930 26010 4 _0995_
rlabel metal1 s 20424 25806 20424 25806 4 _0996_
rlabel metal1 s 20884 26486 20884 26486 4 _0997_
rlabel metal1 s 21114 25942 21114 25942 4 _0998_
rlabel metal2 s 20930 26656 20930 26656 4 _0999_
rlabel metal1 s 21482 26860 21482 26860 4 _1000_
rlabel metal2 s 22770 27302 22770 27302 4 _1001_
rlabel metal2 s 22218 27676 22218 27676 4 _1002_
rlabel metal2 s 21390 29580 21390 29580 4 _1003_
rlabel metal2 s 22034 29750 22034 29750 4 _1004_
rlabel metal2 s 21482 29376 21482 29376 4 _1005_
rlabel metal2 s 20930 28526 20930 28526 4 _1006_
rlabel metal1 s 21919 27982 21919 27982 4 _1007_
rlabel metal1 s 21022 28050 21022 28050 4 _1008_
rlabel metal1 s 21068 27982 21068 27982 4 _1009_
rlabel metal2 s 21850 29954 21850 29954 4 _1010_
rlabel metal1 s 21114 27880 21114 27880 4 _1011_
rlabel metal2 s 21298 28628 21298 28628 4 _1012_
rlabel metal1 s 21390 27574 21390 27574 4 _1013_
rlabel metal2 s 23046 27132 23046 27132 4 _1014_
rlabel metal1 s 21666 27608 21666 27608 4 _1015_
rlabel metal1 s 21850 27438 21850 27438 4 _1016_
rlabel metal2 s 21574 26860 21574 26860 4 _1017_
rlabel metal1 s 21482 26282 21482 26282 4 _1018_
rlabel metal1 s 21574 23120 21574 23120 4 _1019_
rlabel metal1 s 21666 24276 21666 24276 4 _1020_
rlabel metal1 s 21206 23800 21206 23800 4 _1021_
rlabel metal1 s 21850 23188 21850 23188 4 _1022_
rlabel metal1 s 22034 23562 22034 23562 4 _1023_
rlabel metal1 s 21528 24650 21528 24650 4 _1024_
rlabel metal2 s 21022 23936 21022 23936 4 _1025_
rlabel metal1 s 22172 24378 22172 24378 4 _1026_
rlabel metal1 s 22264 24922 22264 24922 4 _1027_
rlabel metal2 s 22310 27846 22310 27846 4 _1028_
rlabel metal2 s 21206 27132 21206 27132 4 _1029_
rlabel metal2 s 22494 26180 22494 26180 4 _1030_
rlabel metal2 s 21298 24548 21298 24548 4 _1031_
rlabel metal2 s 6302 30124 6302 30124 4 _1032_
rlabel metal1 s 4738 14246 4738 14246 4 _1033_
rlabel metal1 s 5658 12614 5658 12614 4 _1034_
rlabel metal1 s 6532 29274 6532 29274 4 _1035_
rlabel metal2 s 21390 26554 21390 26554 4 _1036_
rlabel metal1 s 22126 25262 22126 25262 4 _1037_
rlabel metal1 s 20976 11798 20976 11798 4 _1038_
rlabel metal1 s 20930 11730 20930 11730 4 _1039_
rlabel metal1 s 24334 25398 24334 25398 4 _1040_
rlabel metal1 s 23552 29750 23552 29750 4 _1041_
rlabel metal1 s 15870 16592 15870 16592 4 _1042_
rlabel metal2 s 15502 20094 15502 20094 4 _1043_
rlabel metal2 s 25438 29070 25438 29070 4 _1044_
rlabel metal2 s 23414 29070 23414 29070 4 _1045_
rlabel metal2 s 23138 29376 23138 29376 4 _1046_
rlabel metal2 s 22954 30124 22954 30124 4 _1047_
rlabel metal1 s 23230 29682 23230 29682 4 _1048_
rlabel metal2 s 23782 29104 23782 29104 4 _1049_
rlabel metal2 s 24150 29988 24150 29988 4 _1050_
rlabel metal1 s 23414 27982 23414 27982 4 _1051_
rlabel metal2 s 12742 30532 12742 30532 4 active
rlabel metal1 s 7130 5610 7130 5610 4 amp_A.pwm_out\[0\]
rlabel metal2 s 8602 6018 8602 6018 4 amp_A.pwm_out\[1\]
rlabel metal1 s 5934 6256 5934 6256 4 amp_A.pwm_out\[2\]
rlabel metal1 s 4692 6222 4692 6222 4 amp_A.pwm_out\[3\]
rlabel metal1 s 3864 5066 3864 5066 4 amp_A.pwm_out\[4\]
rlabel metal1 s 2116 6834 2116 6834 4 amp_A.pwm_out\[5\]
rlabel metal1 s 2484 3910 2484 3910 4 amp_A.pwm_out\[6\]
rlabel metal1 s 4462 9384 4462 9384 4 amp_A.pwm_out\[7\]
rlabel metal2 s 15318 5695 15318 5695 4 amp_B.pwm_out\[0\]
rlabel metal1 s 17204 6222 17204 6222 4 amp_B.pwm_out\[1\]
rlabel metal1 s 17664 6834 17664 6834 4 amp_B.pwm_out\[2\]
rlabel metal1 s 15134 8364 15134 8364 4 amp_B.pwm_out\[3\]
rlabel metal1 s 14030 5848 14030 5848 4 amp_B.pwm_out\[4\]
rlabel metal2 s 11822 5780 11822 5780 4 amp_B.pwm_out\[5\]
rlabel metal1 s 10212 5746 10212 5746 4 amp_B.pwm_out\[6\]
rlabel metal1 s 11040 7922 11040 7922 4 amp_B.pwm_out\[7\]
rlabel metal1 s 21896 5814 21896 5814 4 amp_C.pwm_out\[0\]
rlabel metal1 s 25392 4726 25392 4726 4 amp_C.pwm_out\[1\]
rlabel metal1 s 25208 6222 25208 6222 4 amp_C.pwm_out\[2\]
rlabel metal2 s 22954 5270 22954 5270 4 amp_C.pwm_out\[3\]
rlabel metal2 s 24058 7871 24058 7871 4 amp_C.pwm_out\[4\]
rlabel metal1 s 19872 8398 19872 8398 4 amp_C.pwm_out\[5\]
rlabel metal2 s 20286 5814 20286 5814 4 amp_C.pwm_out\[6\]
rlabel metal2 s 18722 6596 18722 6596 4 amp_C.pwm_out\[7\]
rlabel metal1 s 10580 9894 10580 9894 4 amplitude_A\[0\]
rlabel metal2 s 9614 12036 9614 12036 4 amplitude_A\[1\]
rlabel metal1 s 9568 12818 9568 12818 4 amplitude_A\[2\]
rlabel metal2 s 9982 13532 9982 13532 4 amplitude_A\[3\]
rlabel metal1 s 12834 8398 12834 8398 4 amplitude_B\[0\]
rlabel metal2 s 12926 10812 12926 10812 4 amplitude_B\[1\]
rlabel metal1 s 13524 14382 13524 14382 4 amplitude_B\[2\]
rlabel metal2 s 13110 13022 13110 13022 4 amplitude_B\[3\]
rlabel metal2 s 15686 9826 15686 9826 4 amplitude_C\[0\]
rlabel metal2 s 15318 10642 15318 10642 4 amplitude_C\[1\]
rlabel metal1 s 16514 14382 16514 14382 4 amplitude_C\[2\]
rlabel metal1 s 15272 12614 15272 12614 4 amplitude_C\[3\]
rlabel metal1 s 8832 30770 8832 30770 4 bc1
rlabel metal1 s 10350 30770 10350 30770 4 bdir
rlabel metal2 s 9522 1418 9522 1418 4 channel_A_dac_ctrl[0]
rlabel metal1 s 2461 1394 2461 1394 4 channel_A_dac_ctrl[10]
rlabel metal2 s 3450 1418 3450 1418 4 channel_A_dac_ctrl[11]
rlabel metal2 s 2898 568 2898 568 4 channel_A_dac_ctrl[12]
rlabel metal2 s 2346 908 2346 908 4 channel_A_dac_ctrl[13]
rlabel metal2 s 1794 1112 1794 1112 4 channel_A_dac_ctrl[14]
rlabel metal2 s 8970 874 8970 874 4 channel_A_dac_ctrl[1]
rlabel metal2 s 8418 942 8418 942 4 channel_A_dac_ctrl[2]
rlabel metal2 s 7866 568 7866 568 4 channel_A_dac_ctrl[3]
rlabel metal2 s 7286 0 7342 400 4 channel_A_dac_ctrl[4]
port 14 nsew
rlabel metal2 s 6762 551 6762 551 4 channel_A_dac_ctrl[5]
rlabel metal2 s 6210 1418 6210 1418 4 channel_A_dac_ctrl[6]
rlabel metal2 s 5658 874 5658 874 4 channel_A_dac_ctrl[7]
rlabel metal2 s 5106 568 5106 568 4 channel_A_dac_ctrl[8]
rlabel metal2 s 4554 483 4554 483 4 channel_A_dac_ctrl[9]
rlabel metal1 s 4508 30294 4508 30294 4 channel_A_pwm_out
rlabel metal2 s 17802 942 17802 942 4 channel_B_dac_ctrl[0]
rlabel metal2 s 12282 551 12282 551 4 channel_B_dac_ctrl[10]
rlabel metal2 s 11730 568 11730 568 4 channel_B_dac_ctrl[11]
rlabel metal2 s 11178 942 11178 942 4 channel_B_dac_ctrl[12]
rlabel metal2 s 10626 568 10626 568 4 channel_B_dac_ctrl[13]
rlabel metal2 s 10074 1112 10074 1112 4 channel_B_dac_ctrl[14]
rlabel metal2 s 17250 568 17250 568 4 channel_B_dac_ctrl[1]
rlabel metal2 s 16698 874 16698 874 4 channel_B_dac_ctrl[2]
rlabel metal2 s 16146 1112 16146 1112 4 channel_B_dac_ctrl[3]
rlabel metal2 s 15594 874 15594 874 4 channel_B_dac_ctrl[4]
rlabel metal2 s 15042 568 15042 568 4 channel_B_dac_ctrl[5]
rlabel metal2 s 14490 874 14490 874 4 channel_B_dac_ctrl[6]
rlabel metal2 s 13910 0 13966 400 4 channel_B_dac_ctrl[7]
port 33 nsew
rlabel metal2 s 13386 568 13386 568 4 channel_B_dac_ctrl[8]
rlabel metal2 s 12834 1112 12834 1112 4 channel_B_dac_ctrl[9]
rlabel metal2 s 2990 30073 2990 30073 4 channel_B_pwm_out
rlabel metal2 s 26082 568 26082 568 4 channel_C_dac_ctrl[0]
rlabel metal2 s 20534 0 20590 400 4 channel_C_dac_ctrl[10]
port 38 nsew
rlabel metal2 s 20010 551 20010 551 4 channel_C_dac_ctrl[11]
rlabel metal2 s 19458 568 19458 568 4 channel_C_dac_ctrl[12]
rlabel metal2 s 18906 874 18906 874 4 channel_C_dac_ctrl[13]
rlabel metal2 s 18354 568 18354 568 4 channel_C_dac_ctrl[14]
rlabel metal2 s 25530 874 25530 874 4 channel_C_dac_ctrl[1]
rlabel metal2 s 24978 1112 24978 1112 4 channel_C_dac_ctrl[2]
rlabel metal2 s 24426 568 24426 568 4 channel_C_dac_ctrl[3]
rlabel metal2 s 23874 415 23874 415 4 channel_C_dac_ctrl[4]
rlabel metal2 s 23322 568 23322 568 4 channel_C_dac_ctrl[5]
rlabel metal2 s 22770 874 22770 874 4 channel_C_dac_ctrl[6]
rlabel metal2 s 22218 1112 22218 1112 4 channel_C_dac_ctrl[7]
rlabel metal2 s 21666 874 21666 874 4 channel_C_dac_ctrl[8]
rlabel metal2 s 21114 568 21114 568 4 channel_C_dac_ctrl[9]
rlabel metal1 s 1196 29818 1196 29818 4 channel_C_pwm_out
rlabel metal1 s 18906 18768 18906 18768 4 clk
rlabel metal1 s 2714 14552 2714 14552 4 clk_counter\[0\]
rlabel metal1 s 1978 14348 1978 14348 4 clk_counter\[1\]
rlabel metal1 s 3174 14484 3174 14484 4 clk_counter\[2\]
rlabel metal2 s 2254 11900 2254 11900 4 clk_counter\[3\]
rlabel metal1 s 3450 12818 3450 12818 4 clk_counter\[4\]
rlabel metal1 s 4692 12954 4692 12954 4 clk_counter\[5\]
rlabel metal1 s 4462 12716 4462 12716 4 clk_counter\[6\]
rlabel metal1 s 16836 18938 16836 18938 4 clknet_0_clk
rlabel metal4 s 12604 18020 12604 18020 4 clknet_1_0__leaf_clk
rlabel metal3 s 17618 19227 17618 19227 4 clknet_1_1__leaf_clk
rlabel metal2 s 8418 14178 8418 14178 4 clknet_leaf_0_clk
rlabel metal1 s 25346 21590 25346 21590 4 clknet_leaf_10_clk
rlabel metal2 s 27094 17986 27094 17986 4 clknet_leaf_11_clk
rlabel metal2 s 19274 15776 19274 15776 4 clknet_leaf_12_clk
rlabel metal2 s 20746 13056 20746 13056 4 clknet_leaf_13_clk
rlabel metal1 s 25392 16014 25392 16014 4 clknet_leaf_14_clk
rlabel metal2 s 21298 7072 21298 7072 4 clknet_leaf_15_clk
rlabel metal2 s 18170 6052 18170 6052 4 clknet_leaf_16_clk
rlabel metal2 s 16422 13056 16422 13056 4 clknet_leaf_17_clk
rlabel metal1 s 13616 9486 13616 9486 4 clknet_leaf_18_clk
rlabel metal1 s 874 9078 874 9078 4 clknet_leaf_19_clk
rlabel metal1 s 5842 19822 5842 19822 4 clknet_leaf_1_clk
rlabel metal1 s 874 12308 874 12308 4 clknet_leaf_20_clk
rlabel metal2 s 874 18768 874 18768 4 clknet_leaf_2_clk
rlabel metal1 s 966 25330 966 25330 4 clknet_leaf_3_clk
rlabel metal2 s 6486 27472 6486 27472 4 clknet_leaf_4_clk
rlabel metal1 s 7314 24718 7314 24718 4 clknet_leaf_5_clk
rlabel metal2 s 12650 27744 12650 27744 4 clknet_leaf_6_clk
rlabel metal1 s 14996 21998 14996 21998 4 clknet_leaf_7_clk
rlabel metal2 s 15962 24514 15962 24514 4 clknet_leaf_8_clk
rlabel metal1 s 19044 27506 19044 27506 4 clknet_leaf_9_clk
rlabel metal1 s 8096 30770 8096 30770 4 clock_select[0]
rlabel metal1 s 6578 30124 6578 30124 4 clock_select[1]
rlabel metal2 s 22034 31273 22034 31273 4 data[0]
rlabel metal1 s 20884 30838 20884 30838 4 data[1]
rlabel metal1 s 19918 30838 19918 30838 4 data[2]
rlabel metal1 s 18170 30838 18170 30838 4 data[3]
rlabel metal1 s 16790 30804 16790 30804 4 data[4]
rlabel metal1 s 14720 30770 14720 30770 4 data[5]
rlabel metal1 s 13156 30158 13156 30158 4 data[6]
rlabel metal1 s 11776 30770 11776 30770 4 data[7]
rlabel metal1 s 26588 30770 26588 30770 4 ena
rlabel metal1 s 9200 10982 9200 10982 4 envelope_A
rlabel metal1 s 13386 12750 13386 12750 4 envelope_B
rlabel metal1 s 15318 11866 15318 11866 4 envelope_C
rlabel metal2 s 11454 17884 11454 17884 4 envelope_generator.alternate
rlabel metal2 s 10166 16864 10166 16864 4 envelope_generator.attack
rlabel metal1 s 9522 16558 9522 16558 4 envelope_generator.continue_
rlabel metal1 s 6394 13396 6394 13396 4 envelope_generator.envelope_counter\[0\]
rlabel metal1 s 7544 12070 7544 12070 4 envelope_generator.envelope_counter\[1\]
rlabel metal1 s 7130 10064 7130 10064 4 envelope_generator.envelope_counter\[2\]
rlabel metal1 s 7682 9010 7682 9010 4 envelope_generator.envelope_counter\[3\]
rlabel metal1 s 8924 18598 8924 18598 4 envelope_generator.hold
rlabel metal2 s 9614 14620 9614 14620 4 envelope_generator.invert_output
rlabel metal2 s 6210 26860 6210 26860 4 envelope_generator.period\[0\]
rlabel metal1 s 8464 20570 8464 20570 4 envelope_generator.period\[10\]
rlabel metal1 s 7314 19788 7314 19788 4 envelope_generator.period\[11\]
rlabel metal1 s 7774 17306 7774 17306 4 envelope_generator.period\[12\]
rlabel metal2 s 7498 17204 7498 17204 4 envelope_generator.period\[13\]
rlabel metal2 s 6486 18904 6486 18904 4 envelope_generator.period\[14\]
rlabel metal1 s 8280 18938 8280 18938 4 envelope_generator.period\[15\]
rlabel metal1 s 6256 27642 6256 27642 4 envelope_generator.period\[1\]
rlabel metal1 s 8970 25262 8970 25262 4 envelope_generator.period\[2\]
rlabel metal1 s 6026 24582 6026 24582 4 envelope_generator.period\[3\]
rlabel metal1 s 7820 23018 7820 23018 4 envelope_generator.period\[4\]
rlabel metal1 s 6854 23528 6854 23528 4 envelope_generator.period\[5\]
rlabel metal2 s 6946 22236 6946 22236 4 envelope_generator.period\[6\]
rlabel metal2 s 7498 22372 7498 22372 4 envelope_generator.period\[7\]
rlabel metal1 s 6716 21454 6716 21454 4 envelope_generator.period\[8\]
rlabel metal1 s 5106 20876 5106 20876 4 envelope_generator.period\[9\]
rlabel metal1 s 6716 15130 6716 15130 4 envelope_generator.signal_edge.previous_signal_state_0
rlabel metal1 s 4922 15334 4922 15334 4 envelope_generator.signal_edge.signal
rlabel metal2 s 7774 14620 7774 14620 4 envelope_generator.stop
rlabel metal2 s 5382 27234 5382 27234 4 envelope_generator.tone.counter\[0\]
rlabel metal2 s 2254 20196 2254 20196 4 envelope_generator.tone.counter\[10\]
rlabel metal2 s 2530 19074 2530 19074 4 envelope_generator.tone.counter\[11\]
rlabel metal1 s 2392 18190 2392 18190 4 envelope_generator.tone.counter\[12\]
rlabel metal2 s 2530 15572 2530 15572 4 envelope_generator.tone.counter\[13\]
rlabel metal1 s 2438 17612 2438 17612 4 envelope_generator.tone.counter\[14\]
rlabel metal1 s 4094 17646 4094 17646 4 envelope_generator.tone.counter\[15\]
rlabel metal2 s 6118 29546 6118 29546 4 envelope_generator.tone.counter\[1\]
rlabel metal1 s 4830 25262 4830 25262 4 envelope_generator.tone.counter\[2\]
rlabel metal1 s 2645 26214 2645 26214 4 envelope_generator.tone.counter\[3\]
rlabel metal1 s 2714 26520 2714 26520 4 envelope_generator.tone.counter\[4\]
rlabel metal1 s 2300 24174 2300 24174 4 envelope_generator.tone.counter\[5\]
rlabel metal2 s 2254 24922 2254 24922 4 envelope_generator.tone.counter\[6\]
rlabel metal1 s 2944 23562 2944 23562 4 envelope_generator.tone.counter\[7\]
rlabel metal1 s 2438 21318 2438 21318 4 envelope_generator.tone.counter\[8\]
rlabel metal1 s 3312 20978 3312 20978 4 envelope_generator.tone.counter\[9\]
rlabel metal1 s 14720 21454 14720 21454 4 latched_register\[0\]
rlabel metal1 s 14582 21420 14582 21420 4 latched_register\[1\]
rlabel metal1 s 12489 21454 12489 21454 4 latched_register\[2\]
rlabel metal1 s 12650 22032 12650 22032 4 latched_register\[3\]
rlabel metal2 s 11270 30396 11270 30396 4 net1
rlabel metal2 s 19090 17884 19090 17884 4 net10
rlabel metal1 s 16054 13430 16054 13430 4 net100
rlabel metal2 s 20378 17238 20378 17238 4 net101
rlabel metal2 s 6486 21658 6486 21658 4 net102
rlabel metal2 s 18262 26044 18262 26044 4 net103
rlabel metal1 s 18032 17102 18032 17102 4 net104
rlabel metal1 s 8188 14518 8188 14518 4 net105
rlabel metal2 s 6573 14926 6573 14926 4 net106
rlabel metal1 s 6210 26928 6210 26928 4 net107
rlabel metal1 s 19504 27982 19504 27982 4 net108
rlabel metal1 s 18630 15504 18630 15504 4 net109
rlabel metal2 s 17710 18241 17710 18241 4 net11
rlabel metal2 s 24426 24548 24426 24548 4 net110
rlabel metal1 s 22627 23562 22627 23562 4 net111
rlabel metal1 s 18446 16014 18446 16014 4 net112
rlabel metal1 s 17250 26826 17250 26826 4 net113
rlabel metal2 s 21850 18972 21850 18972 4 net114
rlabel metal1 s 17986 26928 17986 26928 4 net115
rlabel metal1 s 21574 20400 21574 20400 4 net116
rlabel metal2 s 6854 24038 6854 24038 4 net117
rlabel metal1 s 4830 12274 4830 12274 4 net118
rlabel metal2 s 1886 15147 1886 15147 4 net119
rlabel metal1 s 14076 30702 14076 30702 4 net12
rlabel metal1 s 18446 21012 18446 21012 4 net120
rlabel metal1 s 18722 30736 18722 30736 4 net121
rlabel metal1 s 24288 13158 24288 13158 4 net122
rlabel metal2 s 24982 12750 24982 12750 4 net123
rlabel metal1 s 26312 11322 26312 11322 4 net124
rlabel metal1 s 25606 12682 25606 12682 4 net125
rlabel metal1 s 23782 14858 23782 14858 4 net126
rlabel metal1 s 25346 11696 25346 11696 4 net127
rlabel metal2 s 18906 8602 18906 8602 4 net128
rlabel metal1 s 23046 13396 23046 13396 4 net129
rlabel metal2 s 19458 31008 19458 31008 4 net13
rlabel metal2 s 22218 13634 22218 13634 4 net130
rlabel metal2 s 7130 22916 7130 22916 4 net131
rlabel metal1 s 18262 17850 18262 17850 4 net132
rlabel metal1 s 8326 25330 8326 25330 4 net133
rlabel metal1 s 26588 23290 26588 23290 4 net134
rlabel metal1 s 17802 19278 17802 19278 4 net135
rlabel metal1 s 26680 14450 26680 14450 4 net136
rlabel metal1 s 25852 9078 25852 9078 4 net137
rlabel metal1 s 24702 10132 24702 10132 4 net138
rlabel metal1 s 25361 11254 25361 11254 4 net139
rlabel metal1 s 16974 22066 16974 22066 4 net14
rlabel metal1 s 23552 10098 23552 10098 4 net140
rlabel metal2 s 23786 9010 23786 9010 4 net141
rlabel metal1 s 26588 15334 26588 15334 4 net142
rlabel metal1 s 20424 19482 20424 19482 4 net143
rlabel metal2 s 26450 8432 26450 8432 4 net144
rlabel metal1 s 24518 9044 24518 9044 4 net145
rlabel metal2 s 24982 8398 24982 8398 4 net146
rlabel metal1 s 23322 11662 23322 11662 4 net147
rlabel metal1 s 26128 7514 26128 7514 4 net148
rlabel metal1 s 7452 10098 7452 10098 4 net149
rlabel metal1 s 25162 782 25162 782 4 net15
rlabel metal1 s 6996 9418 6996 9418 4 net150
rlabel metal2 s 17526 14654 17526 14654 4 net151
rlabel metal2 s 1794 13260 1794 13260 4 net152
rlabel metal2 s 1334 13634 1334 13634 4 net153
rlabel metal1 s 22356 10098 22356 10098 4 net154
rlabel metal2 s 4646 15436 4646 15436 4 net155
rlabel metal1 s 23000 12750 23000 12750 4 net156
rlabel metal1 s 4232 10574 4232 10574 4 net157
rlabel metal1 s 24794 15504 24794 15504 4 net158
rlabel metal1 s 6854 12784 6854 12784 4 net159
rlabel metal2 s 24886 1666 24886 1666 4 net16
rlabel metal2 s 1886 11356 1886 11356 4 net160
rlabel metal1 s 1242 11866 1242 11866 4 net161
rlabel metal1 s 7268 30770 7268 30770 4 net162
rlabel metal1 s 10396 8330 10396 8330 4 net163
rlabel metal1 s 16698 19278 16698 19278 4 net164
rlabel metal1 s 16376 10778 16376 10778 4 net165
rlabel metal1 s 19136 9894 19136 9894 4 net166
rlabel metal2 s 3358 17068 3358 17068 4 net167
rlabel metal1 s 18906 13192 18906 13192 4 net168
rlabel metal2 s 7038 11662 7038 11662 4 net169
rlabel metal1 s 23644 986 23644 986 4 net17
rlabel metal1 s 5980 11662 5980 11662 4 net170
rlabel metal1 s 23736 15538 23736 15538 4 net171
rlabel metal2 s 11730 14620 11730 14620 4 net172
rlabel metal1 s 12052 8602 12052 8602 4 net173
rlabel metal1 s 14536 10778 14536 10778 4 net174
rlabel metal2 s 12282 10166 12282 10166 4 net175
rlabel metal2 s 15226 9792 15226 9792 4 net176
rlabel metal2 s 11178 10166 11178 10166 4 net177
rlabel metal2 s 12834 13056 12834 13056 4 net178
rlabel metal1 s 9798 12104 9798 12104 4 net179
rlabel metal1 s 23828 850 23828 850 4 net18
rlabel metal1 s 8418 26520 8418 26520 4 net180
rlabel metal1 s 24886 21012 24886 21012 4 net181
rlabel metal1 s 22954 10574 22954 10574 4 net182
rlabel metal1 s 14582 13158 14582 13158 4 net183
rlabel metal2 s 10166 22270 10166 22270 4 net184
rlabel metal1 s 9108 12954 9108 12954 4 net185
rlabel metal1 s 13340 19210 13340 19210 4 net186
rlabel metal1 s 13110 14042 13110 14042 4 net187
rlabel metal1 s 15824 14042 15824 14042 4 net188
rlabel metal1 s 10810 12954 10810 12954 4 net189
rlabel metal1 s 23552 1326 23552 1326 4 net19
rlabel metal2 s 13018 25534 13018 25534 4 net190
rlabel metal1 s 19504 14042 19504 14042 4 net191
rlabel metal1 s 7406 21658 7406 21658 4 net192
rlabel metal1 s 8280 19210 8280 19210 4 net193
rlabel metal1 s 11822 26010 11822 26010 4 net194
rlabel metal1 s 14398 17850 14398 17850 4 net195
rlabel metal2 s 7866 25602 7866 25602 4 net196
rlabel metal1 s 13248 16694 13248 16694 4 net197
rlabel metal1 s 14950 24650 14950 24650 4 net198
rlabel metal1 s 10764 24310 10764 24310 4 net199
rlabel metal2 s 11086 30362 11086 30362 4 net2
rlabel metal1 s 22310 782 22310 782 4 net20
rlabel metal1 s 25622 29682 25622 29682 4 net200
rlabel metal1 s 12972 19958 12972 19958 4 net201
rlabel metal2 s 19182 11968 19182 11968 4 net202
rlabel metal1 s 6808 17782 6808 17782 4 net203
rlabel metal2 s 18170 11968 18170 11968 4 net204
rlabel metal1 s 8372 21386 8372 21386 4 net205
rlabel metal2 s 6992 17782 6992 17782 4 net206
rlabel metal2 s 22494 11798 22494 11798 4 net207
rlabel metal2 s 22494 1632 22494 1632 4 net21
rlabel metal1 s 21482 986 21482 986 4 net22
rlabel metal2 s 21298 1156 21298 1156 4 net23
rlabel metal2 s 20010 1020 20010 1020 4 net24
rlabel metal1 s 19504 1870 19504 1870 4 net25
rlabel metal1 s 19504 1326 19504 1326 4 net26
rlabel metal2 s 18722 1360 18722 1360 4 net27
rlabel metal1 s 18262 1326 18262 1326 4 net28
rlabel metal1 s 17526 782 17526 782 4 net29
rlabel metal1 s 5842 30804 5842 30804 4 net3
rlabel metal1 s 19872 5270 19872 5270 4 net30
rlabel metal1 s 24288 4046 24288 4046 4 net31
rlabel metal1 s 24472 3502 24472 3502 4 net32
rlabel metal2 s 22126 4862 22126 4862 4 net33
rlabel metal2 s 22586 5372 22586 5372 4 net34
rlabel metal2 s 18906 5372 18906 5372 4 net35
rlabel metal1 s 19320 4658 19320 4658 4 net36
rlabel metal1 s 17894 4658 17894 4658 4 net37
rlabel metal2 s 17342 1632 17342 1632 4 net38
rlabel metal1 s 16330 782 16330 782 4 net39
rlabel metal2 s 6394 29614 6394 29614 4 net4
rlabel metal1 s 16054 1326 16054 1326 4 net40
rlabel metal2 s 15226 2108 15226 2108 4 net41
rlabel metal2 s 14582 1632 14582 1632 4 net42
rlabel metal1 s 14122 782 14122 782 4 net43
rlabel metal1 s 13524 986 13524 986 4 net44
rlabel metal1 s 13432 1394 13432 1394 4 net45
rlabel metal2 s 12282 1564 12282 1564 4 net46
rlabel metal1 s 11592 1870 11592 1870 4 net47
rlabel metal1 s 10994 1360 10994 1360 4 net48
rlabel metal1 s 10948 850 10948 850 4 net49
rlabel metal1 s 15870 21386 15870 21386 4 net5
rlabel metal1 s 9660 1326 9660 1326 4 net50
rlabel metal2 s 9430 1020 9430 1020 4 net51
rlabel metal2 s 9062 1428 9062 1428 4 net52
rlabel metal2 s 12558 5338 12558 5338 4 net53
rlabel metal2 s 16330 4284 16330 4284 4 net54
rlabel metal2 s 16422 3196 16422 3196 4 net55
rlabel metal1 s 14168 4590 14168 4590 4 net56
rlabel metal2 s 13478 4896 13478 4896 4 net57
rlabel metal1 s 10580 5134 10580 5134 4 net58
rlabel metal1 s 9246 3570 9246 3570 4 net59
rlabel metal1 s 17250 18224 17250 18224 4 net6
rlabel metal2 s 9430 4284 9430 4284 4 net60
rlabel metal1 s 8234 2482 8234 2482 4 net61
rlabel metal2 s 7958 1156 7958 1156 4 net62
rlabel metal1 s 6762 1360 6762 1360 4 net63
rlabel metal2 s 6762 1020 6762 1020 4 net64
rlabel metal2 s 6302 2108 6302 2108 4 net65
rlabel metal1 s 5796 1326 5796 1326 4 net66
rlabel metal1 s 6440 1258 6440 1258 4 net67
rlabel metal2 s 5474 1088 5474 1088 4 net68
rlabel metal2 s 4278 1360 4278 1360 4 net69
rlabel metal1 s 18492 23154 18492 23154 4 net7
rlabel metal1 s 3404 986 3404 986 4 net70
rlabel metal1 s 3496 918 3496 918 4 net71
rlabel metal1 s 2300 2414 2300 2414 4 net72
rlabel metal1 s 2070 782 2070 782 4 net73
rlabel metal1 s 1380 986 1380 986 4 net74
rlabel metal1 s 1012 986 1012 986 4 net75
rlabel metal1 s 6118 5746 6118 5746 4 net76
rlabel metal1 s 8510 4692 8510 4692 4 net77
rlabel metal1 s 4646 5780 4646 5780 4 net78
rlabel metal1 s 4140 5134 4140 5134 4 net79
rlabel metal1 s 13846 21454 13846 21454 4 net8
rlabel metal2 s 2990 4284 2990 4284 4 net80
rlabel metal2 s 1150 5100 1150 5100 4 net81
rlabel metal1 s 1564 4046 1564 4046 4 net82
rlabel metal2 s 4554 5984 4554 5984 4 net83
rlabel metal1 s 16146 17714 16146 17714 4 net84
rlabel metal1 s 14623 17034 14623 17034 4 net85
rlabel metal2 s 20838 21658 20838 21658 4 net86
rlabel metal1 s 20516 11526 20516 11526 4 net87
rlabel metal2 s 24426 16796 24426 16796 4 net88
rlabel metal2 s 23046 16422 23046 16422 4 net89
rlabel metal2 s 16790 30566 16790 30566 4 net9
rlabel metal1 s 19274 29104 19274 29104 4 net90
rlabel metal2 s 17986 21182 17986 21182 4 net91
rlabel metal1 s 7544 25806 7544 25806 4 net92
rlabel metal1 s 18078 26452 18078 26452 4 net93
rlabel metal1 s 12466 30770 12466 30770 4 net94
rlabel metal2 s 18446 28390 18446 28390 4 net95
rlabel metal1 s 16406 27914 16406 27914 4 net96
rlabel metal2 s 6762 24412 6762 24412 4 net97
rlabel metal2 s 7038 23324 7038 23324 4 net98
rlabel metal2 s 18078 30532 18078 30532 4 net99
rlabel metal1 s 20010 12206 20010 12206 4 noise_disable_A
rlabel metal2 s 17894 12036 17894 12036 4 noise_disable_B
rlabel metal2 s 18722 14042 18722 14042 4 noise_disable_C
rlabel metal1 s 17802 10540 17802 10540 4 noise_generator.lfsr\[0\]
rlabel metal2 s 27094 13124 27094 13124 4 noise_generator.lfsr\[10\]
rlabel metal1 s 26220 13158 26220 13158 4 noise_generator.lfsr\[11\]
rlabel metal1 s 26956 13362 26956 13362 4 noise_generator.lfsr\[12\]
rlabel metal2 s 25070 14790 25070 14790 4 noise_generator.lfsr\[13\]
rlabel metal2 s 24886 13124 24886 13124 4 noise_generator.lfsr\[14\]
rlabel metal1 s 24426 13940 24426 13940 4 noise_generator.lfsr\[15\]
rlabel metal1 s 23598 12852 23598 12852 4 noise_generator.lfsr\[16\]
rlabel metal1 s 23920 10574 23920 10574 4 noise_generator.lfsr\[1\]
rlabel metal1 s 23828 10982 23828 10982 4 noise_generator.lfsr\[2\]
rlabel metal2 s 22402 10370 22402 10370 4 noise_generator.lfsr\[3\]
rlabel metal1 s 23414 9554 23414 9554 4 noise_generator.lfsr\[4\]
rlabel metal1 s 25116 7922 25116 7922 4 noise_generator.lfsr\[5\]
rlabel metal1 s 24978 7990 24978 7990 4 noise_generator.lfsr\[6\]
rlabel metal2 s 27094 10302 27094 10302 4 noise_generator.lfsr\[7\]
rlabel metal1 s 26220 10778 26220 10778 4 noise_generator.lfsr\[8\]
rlabel metal1 s 26404 13362 26404 13362 4 noise_generator.lfsr\[9\]
rlabel metal2 s 14674 19618 14674 19618 4 noise_generator.period\[0\]
rlabel metal2 s 12926 19652 12926 19652 4 noise_generator.period\[1\]
rlabel metal1 s 13478 17850 13478 17850 4 noise_generator.period\[2\]
rlabel metal1 s 13708 16014 13708 16014 4 noise_generator.period\[3\]
rlabel metal1 s 14214 15946 14214 15946 4 noise_generator.period\[4\]
rlabel metal1 s 20608 14246 20608 14246 4 noise_generator.signal_edge.previous_signal_state_0
rlabel metal1 s 20884 14450 20884 14450 4 noise_generator.signal_edge.signal
rlabel metal1 s 15686 20570 15686 20570 4 noise_generator.tone.counter\[0\]
rlabel metal2 s 15318 19006 15318 19006 4 noise_generator.tone.counter\[1\]
rlabel metal1 s 15134 18224 15134 18224 4 noise_generator.tone.counter\[2\]
rlabel metal2 s 15318 17102 15318 17102 4 noise_generator.tone.counter\[3\]
rlabel metal1 s 15134 16626 15134 16626 4 noise_generator.tone.counter\[4\]
rlabel metal1 s 7314 5542 7314 5542 4 pwm_A.accumulator\[0\]
rlabel metal2 s 8234 7514 8234 7514 4 pwm_A.accumulator\[1\]
rlabel metal2 s 6624 6834 6624 6834 4 pwm_A.accumulator\[2\]
rlabel metal2 s 5106 7718 5106 7718 4 pwm_A.accumulator\[3\]
rlabel metal2 s 3082 5542 3082 5542 4 pwm_A.accumulator\[4\]
rlabel metal1 s 2300 6834 2300 6834 4 pwm_A.accumulator\[5\]
rlabel metal1 s 2162 8806 2162 8806 4 pwm_A.accumulator\[6\]
rlabel metal1 s 4508 10234 4508 10234 4 pwm_A.accumulator\[7\]
rlabel metal2 s 15502 6018 15502 6018 4 pwm_B.accumulator\[0\]
rlabel metal2 s 17894 6018 17894 6018 4 pwm_B.accumulator\[1\]
rlabel metal2 s 17802 7276 17802 7276 4 pwm_B.accumulator\[2\]
rlabel metal1 s 15272 7786 15272 7786 4 pwm_B.accumulator\[3\]
rlabel metal2 s 13570 5950 13570 5950 4 pwm_B.accumulator\[4\]
rlabel metal1 s 12558 6256 12558 6256 4 pwm_B.accumulator\[5\]
rlabel metal1 s 10212 5814 10212 5814 4 pwm_B.accumulator\[6\]
rlabel metal2 s 10626 8228 10626 8228 4 pwm_B.accumulator\[7\]
rlabel metal1 s 21712 5338 21712 5338 4 pwm_C.accumulator\[0\]
rlabel metal2 s 25714 5236 25714 5236 4 pwm_C.accumulator\[1\]
rlabel metal1 s 26128 6222 26128 6222 4 pwm_C.accumulator\[2\]
rlabel metal1 s 23230 6120 23230 6120 4 pwm_C.accumulator\[3\]
rlabel metal1 s 22770 7888 22770 7888 4 pwm_C.accumulator\[4\]
rlabel metal2 s 19642 8874 19642 8874 4 pwm_C.accumulator\[5\]
rlabel metal1 s 20010 6800 20010 6800 4 pwm_C.accumulator\[6\]
rlabel metal1 s 18814 8942 18814 8942 4 pwm_C.accumulator\[7\]
rlabel metal1 s 11362 15028 11362 15028 4 restart_envelope
rlabel metal1 s 23690 30770 23690 30770 4 rst_n
rlabel metal1 s 26956 29274 26956 29274 4 tone_A_generator.counter\[0\]
rlabel metal2 s 26910 24412 26910 24412 4 tone_A_generator.counter\[10\]
rlabel metal2 s 26910 22916 26910 22916 4 tone_A_generator.counter\[11\]
rlabel metal1 s 20286 27982 20286 27982 4 tone_A_generator.counter\[1\]
rlabel metal2 s 21482 29852 21482 29852 4 tone_A_generator.counter\[2\]
rlabel metal1 s 22011 30294 22011 30294 4 tone_A_generator.counter\[3\]
rlabel metal2 s 24242 27778 24242 27778 4 tone_A_generator.counter\[4\]
rlabel metal1 s 24426 26860 24426 26860 4 tone_A_generator.counter\[5\]
rlabel metal1 s 20746 26384 20746 26384 4 tone_A_generator.counter\[6\]
rlabel metal2 s 21022 26112 21022 26112 4 tone_A_generator.counter\[7\]
rlabel metal2 s 23782 24004 23782 24004 4 tone_A_generator.counter\[8\]
rlabel metal1 s 24610 24310 24610 24310 4 tone_A_generator.counter\[9\]
rlabel metal1 s 19872 11322 19872 11322 4 tone_A_generator.out
rlabel metal1 s 20746 28492 20746 28492 4 tone_A_generator.period\[0\]
rlabel metal1 s 19964 23766 19964 23766 4 tone_A_generator.period\[10\]
rlabel metal2 s 18170 24004 18170 24004 4 tone_A_generator.period\[11\]
rlabel metal1 s 20194 29580 20194 29580 4 tone_A_generator.period\[1\]
rlabel metal2 s 20470 29954 20470 29954 4 tone_A_generator.period\[2\]
rlabel metal1 s 21390 30294 21390 30294 4 tone_A_generator.period\[3\]
rlabel metal1 s 19780 26894 19780 26894 4 tone_A_generator.period\[4\]
rlabel metal1 s 20470 26826 20470 26826 4 tone_A_generator.period\[5\]
rlabel metal1 s 19274 25466 19274 25466 4 tone_A_generator.period\[6\]
rlabel metal1 s 20102 25704 20102 25704 4 tone_A_generator.period\[7\]
rlabel metal1 s 20838 24242 20838 24242 4 tone_A_generator.period\[8\]
rlabel metal1 s 21022 23018 21022 23018 4 tone_A_generator.period\[9\]
rlabel metal2 s 8050 30532 8050 30532 4 tone_B_generator.counter\[0\]
rlabel metal1 s 17572 26418 17572 26418 4 tone_B_generator.counter\[10\]
rlabel metal1 s 17756 28050 17756 28050 4 tone_B_generator.counter\[11\]
rlabel metal2 s 8510 27166 8510 27166 4 tone_B_generator.counter\[1\]
rlabel metal1 s 9292 29818 9292 29818 4 tone_B_generator.counter\[2\]
rlabel metal2 s 10626 29852 10626 29852 4 tone_B_generator.counter\[3\]
rlabel metal1 s 10994 28560 10994 28560 4 tone_B_generator.counter\[4\]
rlabel metal1 s 12098 27540 12098 27540 4 tone_B_generator.counter\[5\]
rlabel metal1 s 13294 29070 13294 29070 4 tone_B_generator.counter\[6\]
rlabel metal1 s 14352 28186 14352 28186 4 tone_B_generator.counter\[7\]
rlabel metal2 s 14582 29852 14582 29852 4 tone_B_generator.counter\[8\]
rlabel metal1 s 15778 29070 15778 29070 4 tone_B_generator.counter\[9\]
rlabel metal1 s 16698 12954 16698 12954 4 tone_B_generator.out
rlabel metal1 s 9844 22746 9844 22746 4 tone_B_generator.period\[0\]
rlabel metal1 s 17388 26350 17388 26350 4 tone_B_generator.period\[10\]
rlabel metal1 s 15686 23188 15686 23188 4 tone_B_generator.period\[11\]
rlabel metal2 s 9338 27234 9338 27234 4 tone_B_generator.period\[1\]
rlabel metal2 s 10166 26316 10166 26316 4 tone_B_generator.period\[2\]
rlabel metal1 s 10350 26010 10350 26010 4 tone_B_generator.period\[3\]
rlabel metal1 s 11316 26894 11316 26894 4 tone_B_generator.period\[4\]
rlabel metal2 s 12834 26384 12834 26384 4 tone_B_generator.period\[5\]
rlabel metal1 s 13202 23834 13202 23834 4 tone_B_generator.period\[6\]
rlabel metal1 s 13754 26860 13754 26860 4 tone_B_generator.period\[7\]
rlabel metal1 s 14674 26894 14674 26894 4 tone_B_generator.period\[8\]
rlabel metal2 s 15594 26962 15594 26962 4 tone_B_generator.period\[9\]
rlabel metal1 s 22494 20910 22494 20910 4 tone_C_generator.counter\[0\]
rlabel metal1 s 23644 15470 23644 15470 4 tone_C_generator.counter\[10\]
rlabel metal2 s 24150 16932 24150 16932 4 tone_C_generator.counter\[11\]
rlabel metal1 s 21160 20978 21160 20978 4 tone_C_generator.counter\[1\]
rlabel metal2 s 22218 21760 22218 21760 4 tone_C_generator.counter\[2\]
rlabel metal2 s 23230 20638 23230 20638 4 tone_C_generator.counter\[3\]
rlabel metal1 s 23414 19890 23414 19890 4 tone_C_generator.counter\[4\]
rlabel metal2 s 23230 18530 23230 18530 4 tone_C_generator.counter\[5\]
rlabel metal1 s 24840 18190 24840 18190 4 tone_C_generator.counter\[6\]
rlabel metal1 s 24794 17850 24794 17850 4 tone_C_generator.counter\[7\]
rlabel metal1 s 25392 17034 25392 17034 4 tone_C_generator.counter\[8\]
rlabel metal2 s 21666 16286 21666 16286 4 tone_C_generator.counter\[9\]
rlabel metal1 s 19366 13260 19366 13260 4 tone_C_generator.out
rlabel metal1 s 20930 21998 20930 21998 4 tone_C_generator.period\[0\]
rlabel metal1 s 20470 15674 20470 15674 4 tone_C_generator.period\[10\]
rlabel metal2 s 21114 15776 21114 15776 4 tone_C_generator.period\[11\]
rlabel metal1 s 19274 21556 19274 21556 4 tone_C_generator.period\[1\]
rlabel metal1 s 21827 21454 21827 21454 4 tone_C_generator.period\[2\]
rlabel metal1 s 21620 19958 21620 19958 4 tone_C_generator.period\[3\]
rlabel metal1 s 19688 20434 19688 20434 4 tone_C_generator.period\[4\]
rlabel metal1 s 21390 19210 21390 19210 4 tone_C_generator.period\[5\]
rlabel metal2 s 20930 18462 20930 18462 4 tone_C_generator.period\[6\]
rlabel metal1 s 21390 18394 21390 18394 4 tone_C_generator.period\[7\]
rlabel metal2 s 21022 16898 21022 16898 4 tone_C_generator.period\[8\]
rlabel metal1 s 19642 16626 19642 16626 4 tone_C_generator.period\[9\]
rlabel metal2 s 20102 10982 20102 10982 4 tone_disable_A
rlabel metal2 s 17066 10404 17066 10404 4 tone_disable_B
rlabel metal1 s 17802 13260 17802 13260 4 tone_disable_C
flabel metal4 s 27256 496 27576 31056 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 20540 496 20860 31056 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 13824 496 14144 31056 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 7108 496 7428 31056 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 23898 496 24218 31056 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 17182 496 17502 31056 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 10466 496 10786 31056 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 3750 496 4070 31056 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal2 s 8758 31600 8814 32000 0 FreeSans 280 90 0 0 bc1
port 3 nsew
flabel metal2 s 10230 31600 10286 32000 0 FreeSans 280 90 0 0 bdir
port 4 nsew
flabel metal2 s 9494 0 9550 400 0 FreeSans 280 90 0 0 channel_A_dac_ctrl[0]
port 5 nsew
flabel metal2 s 3974 0 4030 400 0 FreeSans 280 90 0 0 channel_A_dac_ctrl[10]
port 6 nsew
flabel metal2 s 3422 0 3478 400 0 FreeSans 280 90 0 0 channel_A_dac_ctrl[11]
port 7 nsew
flabel metal2 s 2870 0 2926 400 0 FreeSans 280 90 0 0 channel_A_dac_ctrl[12]
port 8 nsew
flabel metal2 s 2318 0 2374 400 0 FreeSans 280 90 0 0 channel_A_dac_ctrl[13]
port 9 nsew
flabel metal2 s 1766 0 1822 400 0 FreeSans 280 90 0 0 channel_A_dac_ctrl[14]
port 10 nsew
flabel metal2 s 8942 0 8998 400 0 FreeSans 280 90 0 0 channel_A_dac_ctrl[1]
port 11 nsew
flabel metal2 s 8390 0 8446 400 0 FreeSans 280 90 0 0 channel_A_dac_ctrl[2]
port 12 nsew
flabel metal2 s 7838 0 7894 400 0 FreeSans 280 90 0 0 channel_A_dac_ctrl[3]
port 13 nsew
flabel metal2 s 7314 200 7314 200 0 FreeSans 280 90 0 0 channel_A_dac_ctrl[4]
flabel metal2 s 6734 0 6790 400 0 FreeSans 280 90 0 0 channel_A_dac_ctrl[5]
port 15 nsew
flabel metal2 s 6182 0 6238 400 0 FreeSans 280 90 0 0 channel_A_dac_ctrl[6]
port 16 nsew
flabel metal2 s 5630 0 5686 400 0 FreeSans 280 90 0 0 channel_A_dac_ctrl[7]
port 17 nsew
flabel metal2 s 5078 0 5134 400 0 FreeSans 280 90 0 0 channel_A_dac_ctrl[8]
port 18 nsew
flabel metal2 s 4526 0 4582 400 0 FreeSans 280 90 0 0 channel_A_dac_ctrl[9]
port 19 nsew
flabel metal2 s 4342 31600 4398 32000 0 FreeSans 280 90 0 0 channel_A_pwm_out
port 20 nsew
flabel metal2 s 17774 0 17830 400 0 FreeSans 280 90 0 0 channel_B_dac_ctrl[0]
port 21 nsew
flabel metal2 s 12254 0 12310 400 0 FreeSans 280 90 0 0 channel_B_dac_ctrl[10]
port 22 nsew
flabel metal2 s 11702 0 11758 400 0 FreeSans 280 90 0 0 channel_B_dac_ctrl[11]
port 23 nsew
flabel metal2 s 11150 0 11206 400 0 FreeSans 280 90 0 0 channel_B_dac_ctrl[12]
port 24 nsew
flabel metal2 s 10598 0 10654 400 0 FreeSans 280 90 0 0 channel_B_dac_ctrl[13]
port 25 nsew
flabel metal2 s 10046 0 10102 400 0 FreeSans 280 90 0 0 channel_B_dac_ctrl[14]
port 26 nsew
flabel metal2 s 17222 0 17278 400 0 FreeSans 280 90 0 0 channel_B_dac_ctrl[1]
port 27 nsew
flabel metal2 s 16670 0 16726 400 0 FreeSans 280 90 0 0 channel_B_dac_ctrl[2]
port 28 nsew
flabel metal2 s 16118 0 16174 400 0 FreeSans 280 90 0 0 channel_B_dac_ctrl[3]
port 29 nsew
flabel metal2 s 15566 0 15622 400 0 FreeSans 280 90 0 0 channel_B_dac_ctrl[4]
port 30 nsew
flabel metal2 s 15014 0 15070 400 0 FreeSans 280 90 0 0 channel_B_dac_ctrl[5]
port 31 nsew
flabel metal2 s 14462 0 14518 400 0 FreeSans 280 90 0 0 channel_B_dac_ctrl[6]
port 32 nsew
flabel metal2 s 13938 200 13938 200 0 FreeSans 280 90 0 0 channel_B_dac_ctrl[7]
flabel metal2 s 13358 0 13414 400 0 FreeSans 280 90 0 0 channel_B_dac_ctrl[8]
port 34 nsew
flabel metal2 s 12806 0 12862 400 0 FreeSans 280 90 0 0 channel_B_dac_ctrl[9]
port 35 nsew
flabel metal2 s 2870 31600 2926 32000 0 FreeSans 280 90 0 0 channel_B_pwm_out
port 36 nsew
flabel metal2 s 26054 0 26110 400 0 FreeSans 280 90 0 0 channel_C_dac_ctrl[0]
port 37 nsew
flabel metal2 s 20562 200 20562 200 0 FreeSans 280 90 0 0 channel_C_dac_ctrl[10]
flabel metal2 s 19982 0 20038 400 0 FreeSans 280 90 0 0 channel_C_dac_ctrl[11]
port 39 nsew
flabel metal2 s 19430 0 19486 400 0 FreeSans 280 90 0 0 channel_C_dac_ctrl[12]
port 40 nsew
flabel metal2 s 18878 0 18934 400 0 FreeSans 280 90 0 0 channel_C_dac_ctrl[13]
port 41 nsew
flabel metal2 s 18326 0 18382 400 0 FreeSans 280 90 0 0 channel_C_dac_ctrl[14]
port 42 nsew
flabel metal2 s 25502 0 25558 400 0 FreeSans 280 90 0 0 channel_C_dac_ctrl[1]
port 43 nsew
flabel metal2 s 24950 0 25006 400 0 FreeSans 280 90 0 0 channel_C_dac_ctrl[2]
port 44 nsew
flabel metal2 s 24398 0 24454 400 0 FreeSans 280 90 0 0 channel_C_dac_ctrl[3]
port 45 nsew
flabel metal2 s 23846 0 23902 400 0 FreeSans 280 90 0 0 channel_C_dac_ctrl[4]
port 46 nsew
flabel metal2 s 23294 0 23350 400 0 FreeSans 280 90 0 0 channel_C_dac_ctrl[5]
port 47 nsew
flabel metal2 s 22742 0 22798 400 0 FreeSans 280 90 0 0 channel_C_dac_ctrl[6]
port 48 nsew
flabel metal2 s 22190 0 22246 400 0 FreeSans 280 90 0 0 channel_C_dac_ctrl[7]
port 49 nsew
flabel metal2 s 21638 0 21694 400 0 FreeSans 280 90 0 0 channel_C_dac_ctrl[8]
port 50 nsew
flabel metal2 s 21086 0 21142 400 0 FreeSans 280 90 0 0 channel_C_dac_ctrl[9]
port 51 nsew
flabel metal2 s 1398 31600 1454 32000 0 FreeSans 280 90 0 0 channel_C_pwm_out
port 52 nsew
flabel metal2 s 24950 31600 25006 32000 0 FreeSans 280 90 0 0 clk
port 53 nsew
flabel metal2 s 7286 31600 7342 32000 0 FreeSans 280 90 0 0 clock_select[0]
port 54 nsew
flabel metal2 s 5814 31600 5870 32000 0 FreeSans 280 90 0 0 clock_select[1]
port 55 nsew
flabel metal2 s 22006 31600 22062 32000 0 FreeSans 280 90 0 0 data[0]
port 56 nsew
flabel metal2 s 20534 31600 20590 32000 0 FreeSans 280 90 0 0 data[1]
port 57 nsew
flabel metal2 s 19062 31600 19118 32000 0 FreeSans 280 90 0 0 data[2]
port 58 nsew
flabel metal2 s 17590 31600 17646 32000 0 FreeSans 280 90 0 0 data[3]
port 59 nsew
flabel metal2 s 16118 31600 16174 32000 0 FreeSans 280 90 0 0 data[4]
port 60 nsew
flabel metal2 s 14646 31600 14702 32000 0 FreeSans 280 90 0 0 data[5]
port 61 nsew
flabel metal2 s 13174 31600 13230 32000 0 FreeSans 280 90 0 0 data[6]
port 62 nsew
flabel metal2 s 11702 31600 11758 32000 0 FreeSans 280 90 0 0 data[7]
port 63 nsew
flabel metal2 s 26422 31600 26478 32000 0 FreeSans 280 90 0 0 ena
port 64 nsew
flabel metal2 s 23478 31600 23534 32000 0 FreeSans 280 90 0 0 rst_n
port 65 nsew
<< properties >>
string FIXED_BBOX 0 0 28000 32000
string GDS_END 3701956
string GDS_FILE ../gds/ay8913.gds
string GDS_START 525914
<< end >>
