magic
tech sky130A
magscale 1 2
timestamp 1717253211
<< viali >>
rect 949 30889 983 30923
rect 9781 30821 9815 30855
rect 17877 30821 17911 30855
rect 19625 30821 19659 30855
rect 20269 30821 20303 30855
rect 23397 30821 23431 30855
rect 2073 30753 2107 30787
rect 3893 30753 3927 30787
rect 6101 30753 6135 30787
rect 7573 30753 7607 30787
rect 8585 30753 8619 30787
rect 8861 30753 8895 30787
rect 9505 30753 9539 30787
rect 9689 30753 9723 30787
rect 9873 30753 9907 30787
rect 10977 30753 11011 30787
rect 11989 30753 12023 30787
rect 12357 30753 12391 30787
rect 12541 30753 12575 30787
rect 14289 30753 14323 30787
rect 14749 30753 14783 30787
rect 15301 30753 15335 30787
rect 16221 30753 16255 30787
rect 16957 30753 16991 30787
rect 18061 30753 18095 30787
rect 19441 30753 19475 30787
rect 19533 30753 19567 30787
rect 19809 30753 19843 30787
rect 19993 30753 20027 30787
rect 21557 30753 21591 30787
rect 23305 30753 23339 30787
rect 23489 30753 23523 30787
rect 23673 30753 23707 30787
rect 23857 30753 23891 30787
rect 26709 30753 26743 30787
rect 2329 30685 2363 30719
rect 10149 30685 10183 30719
rect 10701 30685 10735 30719
rect 11253 30685 11287 30719
rect 11805 30685 11839 30719
rect 14105 30685 14139 30719
rect 20821 30685 20855 30719
rect 21741 30685 21775 30719
rect 22477 30685 22511 30719
rect 10057 30617 10091 30651
rect 11161 30617 11195 30651
rect 14473 30617 14507 30651
rect 17141 30617 17175 30651
rect 22293 30617 22327 30651
rect 3709 30549 3743 30583
rect 5917 30549 5951 30583
rect 7389 30549 7423 30583
rect 8493 30549 8527 30583
rect 9045 30549 9079 30583
rect 12173 30549 12207 30583
rect 12449 30549 12483 30583
rect 13553 30549 13587 30583
rect 14933 30549 14967 30583
rect 15117 30549 15151 30583
rect 16405 30549 16439 30583
rect 17785 30549 17819 30583
rect 18245 30549 18279 30583
rect 19257 30549 19291 30583
rect 20085 30549 20119 30583
rect 21373 30549 21407 30583
rect 23029 30549 23063 30583
rect 23121 30549 23155 30583
rect 24041 30549 24075 30583
rect 26525 30549 26559 30583
rect 5733 30345 5767 30379
rect 13185 30345 13219 30379
rect 15209 30345 15243 30379
rect 16221 30345 16255 30379
rect 20729 30345 20763 30379
rect 22661 30345 22695 30379
rect 2973 30277 3007 30311
rect 5181 30277 5215 30311
rect 6101 30277 6135 30311
rect 7757 30277 7791 30311
rect 13001 30277 13035 30311
rect 17049 30277 17083 30311
rect 4813 30209 4847 30243
rect 13829 30209 13863 30243
rect 16037 30209 16071 30243
rect 21281 30209 21315 30243
rect 24593 30209 24627 30243
rect 1593 30141 1627 30175
rect 3341 30141 3375 30175
rect 5825 30141 5859 30175
rect 5917 30141 5951 30175
rect 6193 30141 6227 30175
rect 9965 30141 9999 30175
rect 11529 30141 11563 30175
rect 11621 30141 11655 30175
rect 13093 30141 13127 30175
rect 13277 30141 13311 30175
rect 14096 30141 14130 30175
rect 15485 30141 15519 30175
rect 16313 30141 16347 30175
rect 16405 30141 16439 30175
rect 18162 30141 18196 30175
rect 18429 30141 18463 30175
rect 19349 30141 19383 30175
rect 19616 30141 19650 30175
rect 20821 30141 20855 30175
rect 22937 30141 22971 30175
rect 23305 30141 23339 30175
rect 23397 30141 23431 30175
rect 24041 30141 24075 30175
rect 24501 30141 24535 30175
rect 24685 30141 24719 30175
rect 24961 30141 24995 30175
rect 1860 30073 1894 30107
rect 3608 30073 3642 30107
rect 6438 30073 6472 30107
rect 8125 30073 8159 30107
rect 9698 30073 9732 30107
rect 11262 30073 11296 30107
rect 11888 30073 11922 30107
rect 15393 30073 15427 30107
rect 16681 30073 16715 30107
rect 21548 30073 21582 30107
rect 23029 30073 23063 30107
rect 23121 30073 23155 30107
rect 23489 30073 23523 30107
rect 24409 30073 24443 30107
rect 4721 30005 4755 30039
rect 5273 30005 5307 30039
rect 5365 30005 5399 30039
rect 7573 30005 7607 30039
rect 7665 30005 7699 30039
rect 8585 30005 8619 30039
rect 10149 30005 10183 30039
rect 15761 30005 15795 30039
rect 21005 30005 21039 30039
rect 22753 30005 22787 30039
rect 23857 30005 23891 30039
rect 24133 30005 24167 30039
rect 24225 30005 24259 30039
rect 24869 30005 24903 30039
rect 4077 29801 4111 29835
rect 6193 29801 6227 29835
rect 7021 29801 7055 29835
rect 7205 29801 7239 29835
rect 12357 29801 12391 29835
rect 12725 29801 12759 29835
rect 14381 29801 14415 29835
rect 15133 29801 15167 29835
rect 15301 29801 15335 29835
rect 16313 29801 16347 29835
rect 16773 29801 16807 29835
rect 22937 29801 22971 29835
rect 24317 29801 24351 29835
rect 24501 29801 24535 29835
rect 3893 29733 3927 29767
rect 4537 29733 4571 29767
rect 11222 29733 11256 29767
rect 12449 29733 12483 29767
rect 12909 29733 12943 29767
rect 14013 29733 14047 29767
rect 14491 29733 14525 29767
rect 14933 29733 14967 29767
rect 15623 29733 15657 29767
rect 15793 29733 15827 29767
rect 16497 29733 16531 29767
rect 16957 29733 16991 29767
rect 18622 29733 18656 29767
rect 1961 29665 1995 29699
rect 2217 29665 2251 29699
rect 3525 29665 3559 29699
rect 4261 29665 4295 29699
rect 4445 29665 4479 29699
rect 4721 29665 4755 29699
rect 5181 29665 5215 29699
rect 6009 29665 6043 29699
rect 6837 29665 6871 29699
rect 6929 29665 6963 29699
rect 7297 29665 7331 29699
rect 7748 29665 7782 29699
rect 8125 29665 8159 29699
rect 8309 29665 8343 29699
rect 8585 29665 8619 29699
rect 8677 29665 8711 29699
rect 8769 29665 8803 29699
rect 9689 29665 9723 29699
rect 10057 29665 10091 29699
rect 10241 29665 10275 29699
rect 10333 29665 10367 29699
rect 10425 29665 10459 29699
rect 13866 29665 13900 29699
rect 14197 29665 14231 29699
rect 14381 29665 14415 29699
rect 14657 29665 14691 29699
rect 16405 29665 16439 29699
rect 18889 29665 18923 29699
rect 19441 29665 19475 29699
rect 19708 29665 19742 29699
rect 22405 29665 22439 29699
rect 22934 29665 22968 29699
rect 23397 29665 23431 29699
rect 23489 29665 23523 29699
rect 23673 29665 23707 29699
rect 23857 29665 23891 29699
rect 24024 29665 24058 29699
rect 24442 29665 24476 29699
rect 24869 29665 24903 29699
rect 24961 29665 24995 29699
rect 25513 29665 25547 29699
rect 4353 29597 4387 29631
rect 5089 29597 5123 29631
rect 5825 29597 5859 29631
rect 7205 29597 7239 29631
rect 7573 29597 7607 29631
rect 9597 29597 9631 29631
rect 10977 29597 11011 29631
rect 12817 29597 12851 29631
rect 13645 29597 13679 29631
rect 22661 29597 22695 29631
rect 23765 29597 23799 29631
rect 5549 29529 5583 29563
rect 7389 29529 7423 29563
rect 10609 29529 10643 29563
rect 13369 29529 13403 29563
rect 16129 29529 16163 29563
rect 17325 29529 17359 29563
rect 22753 29529 22787 29563
rect 25053 29529 25087 29563
rect 3341 29461 3375 29495
rect 3893 29461 3927 29495
rect 4905 29461 4939 29495
rect 9413 29461 9447 29495
rect 13093 29461 13127 29495
rect 13737 29461 13771 29495
rect 14841 29461 14875 29495
rect 15117 29461 15151 29495
rect 15761 29461 15795 29495
rect 15945 29461 15979 29495
rect 16681 29461 16715 29495
rect 16957 29461 16991 29495
rect 17509 29461 17543 29495
rect 20821 29461 20855 29495
rect 21281 29461 21315 29495
rect 23305 29461 23339 29495
rect 24225 29461 24259 29495
rect 25237 29461 25271 29495
rect 3709 29257 3743 29291
rect 4537 29257 4571 29291
rect 4997 29257 5031 29291
rect 6469 29257 6503 29291
rect 6929 29257 6963 29291
rect 7481 29257 7515 29291
rect 8125 29257 8159 29291
rect 8677 29257 8711 29291
rect 13829 29257 13863 29291
rect 17141 29257 17175 29291
rect 17325 29257 17359 29291
rect 19533 29257 19567 29291
rect 24225 29257 24259 29291
rect 4261 29189 4295 29223
rect 5181 29189 5215 29223
rect 5457 29189 5491 29223
rect 16773 29189 16807 29223
rect 18521 29189 18555 29223
rect 23857 29189 23891 29223
rect 24593 29189 24627 29223
rect 25329 29189 25363 29223
rect 19993 29121 20027 29155
rect 20637 29121 20671 29155
rect 24961 29121 24995 29155
rect 3709 29053 3743 29087
rect 3893 29053 3927 29087
rect 4345 29055 4379 29089
rect 4445 29053 4479 29087
rect 4629 29053 4663 29087
rect 5273 29053 5307 29087
rect 6377 29053 6411 29087
rect 6653 29053 6687 29087
rect 6745 29053 6779 29087
rect 7205 29053 7239 29087
rect 7297 29053 7331 29087
rect 7573 29053 7607 29087
rect 7849 29053 7883 29087
rect 7941 29053 7975 29087
rect 8217 29053 8251 29087
rect 8861 29053 8895 29087
rect 9229 29053 9263 29087
rect 11897 29053 11931 29087
rect 12265 29053 12299 29087
rect 12357 29053 12391 29087
rect 13001 29053 13035 29087
rect 13553 29053 13587 29087
rect 13645 29053 13679 29087
rect 14013 29053 14047 29087
rect 14933 29053 14967 29087
rect 15117 29053 15151 29087
rect 15669 29053 15703 29087
rect 15761 29053 15795 29087
rect 17785 29053 17819 29087
rect 17969 29053 18003 29087
rect 18153 29053 18187 29087
rect 18337 29053 18371 29087
rect 18705 29053 18739 29087
rect 18981 29053 19015 29087
rect 19165 29053 19199 29087
rect 19257 29053 19291 29087
rect 19349 29053 19383 29087
rect 21281 29053 21315 29087
rect 21649 29053 21683 29087
rect 26709 29053 26743 29087
rect 4813 28985 4847 29019
rect 5018 28985 5052 29019
rect 7665 28985 7699 29019
rect 8953 28985 8987 29019
rect 9045 28985 9079 29019
rect 11069 28985 11103 29019
rect 11989 28985 12023 29019
rect 12081 28985 12115 29019
rect 15025 28985 15059 29019
rect 17141 28985 17175 29019
rect 17417 28985 17451 29019
rect 17601 28985 17635 29019
rect 18245 28985 18279 29019
rect 20729 28985 20763 29019
rect 24225 28985 24259 29019
rect 26442 28985 26476 29019
rect 7021 28917 7055 28951
rect 9597 28917 9631 28951
rect 11713 28917 11747 28951
rect 15577 28917 15611 28951
rect 15853 28917 15887 28951
rect 18889 28917 18923 28951
rect 21465 28917 21499 28951
rect 24409 28917 24443 28951
rect 24501 28917 24535 28951
rect 3249 28713 3283 28747
rect 7389 28713 7423 28747
rect 10057 28713 10091 28747
rect 16513 28713 16547 28747
rect 17417 28713 17451 28747
rect 24869 28713 24903 28747
rect 25697 28713 25731 28747
rect 4229 28645 4263 28679
rect 4445 28645 4479 28679
rect 11244 28645 11278 28679
rect 16313 28645 16347 28679
rect 17233 28645 17267 28679
rect 17877 28645 17911 28679
rect 19082 28645 19116 28679
rect 21548 28645 21582 28679
rect 25037 28645 25071 28679
rect 25237 28645 25271 28679
rect 2136 28577 2170 28611
rect 3525 28577 3559 28611
rect 3617 28577 3651 28611
rect 3801 28577 3835 28611
rect 5825 28577 5859 28611
rect 6081 28577 6115 28611
rect 7297 28577 7331 28611
rect 7481 28577 7515 28611
rect 7573 28577 7607 28611
rect 7757 28577 7791 28611
rect 8493 28577 8527 28611
rect 8585 28577 8619 28611
rect 8944 28577 8978 28611
rect 10701 28577 10735 28611
rect 13073 28577 13107 28611
rect 15485 28577 15519 28611
rect 15577 28577 15611 28611
rect 15761 28577 15795 28611
rect 17509 28577 17543 28611
rect 17693 28577 17727 28611
rect 19789 28577 19823 28611
rect 21281 28577 21315 28611
rect 23121 28577 23155 28611
rect 24593 28577 24627 28611
rect 25329 28577 25363 28611
rect 25504 28577 25538 28611
rect 25605 28577 25639 28611
rect 25881 28577 25915 28611
rect 1869 28509 1903 28543
rect 8677 28509 8711 28543
rect 10977 28509 11011 28543
rect 12817 28509 12851 28543
rect 14933 28509 14967 28543
rect 19349 28509 19383 28543
rect 19533 28509 19567 28543
rect 3985 28441 4019 28475
rect 7665 28441 7699 28475
rect 14197 28441 14231 28475
rect 16681 28441 16715 28475
rect 16865 28441 16899 28475
rect 17969 28441 18003 28475
rect 24777 28441 24811 28475
rect 4077 28373 4111 28407
rect 4261 28373 4295 28407
rect 7205 28373 7239 28407
rect 10149 28373 10183 28407
rect 12357 28373 12391 28407
rect 14289 28373 14323 28407
rect 15025 28373 15059 28407
rect 15393 28373 15427 28407
rect 15669 28373 15703 28407
rect 16497 28373 16531 28407
rect 17233 28373 17267 28407
rect 20913 28373 20947 28407
rect 22661 28373 22695 28407
rect 22937 28373 22971 28407
rect 25053 28373 25087 28407
rect 25421 28373 25455 28407
rect 26065 28373 26099 28407
rect 2237 28169 2271 28203
rect 4537 28169 4571 28203
rect 12725 28169 12759 28203
rect 16037 28169 16071 28203
rect 21649 28169 21683 28203
rect 21833 28169 21867 28203
rect 24961 28169 24995 28203
rect 25421 28169 25455 28203
rect 25605 28169 25639 28203
rect 3065 28101 3099 28135
rect 6837 28101 6871 28135
rect 10885 28101 10919 28135
rect 6929 28033 6963 28067
rect 9505 28033 9539 28067
rect 11529 28033 11563 28067
rect 16129 28033 16163 28067
rect 22293 28033 22327 28067
rect 2421 27965 2455 27999
rect 2697 27965 2731 27999
rect 3065 27965 3099 27999
rect 6653 27965 6687 27999
rect 6745 27965 6779 27999
rect 7941 27965 7975 27999
rect 8033 27965 8067 27999
rect 8677 27965 8711 27999
rect 9045 27965 9079 27999
rect 9137 27965 9171 27999
rect 9413 27965 9447 27999
rect 12541 27965 12575 27999
rect 12909 27965 12943 27999
rect 13001 27965 13035 27999
rect 13277 27965 13311 27999
rect 13553 27965 13587 27999
rect 13645 27965 13679 27999
rect 14657 27965 14691 27999
rect 14841 27965 14875 27999
rect 14933 27965 14967 27999
rect 15025 27965 15059 27999
rect 15209 27965 15243 27999
rect 15610 27965 15644 27999
rect 16405 27965 16439 27999
rect 16589 27965 16623 27999
rect 16681 27965 16715 27999
rect 16773 27965 16807 27999
rect 17141 27965 17175 27999
rect 22201 27965 22235 27999
rect 23857 27965 23891 27999
rect 24041 27965 24075 27999
rect 24133 27965 24167 27999
rect 24317 27965 24351 27999
rect 24409 27965 24443 27999
rect 25053 27965 25087 27999
rect 27077 27965 27111 27999
rect 2789 27897 2823 27931
rect 2973 27897 3007 27931
rect 3249 27897 3283 27931
rect 9229 27897 9263 27931
rect 9772 27897 9806 27931
rect 13093 27897 13127 27931
rect 17049 27897 17083 27931
rect 17386 27897 17420 27931
rect 19809 27897 19843 27931
rect 21557 27897 21591 27931
rect 22560 27897 22594 27931
rect 24593 27897 24627 27931
rect 24777 27897 24811 27931
rect 26810 27897 26844 27931
rect 2513 27829 2547 27863
rect 7757 27829 7791 27863
rect 8585 27829 8619 27863
rect 8861 27829 8895 27863
rect 10977 27829 11011 27863
rect 11989 27829 12023 27863
rect 15393 27829 15427 27863
rect 15485 27829 15519 27863
rect 15669 27829 15703 27863
rect 18521 27829 18555 27863
rect 21833 27829 21867 27863
rect 23673 27829 23707 27863
rect 25421 27829 25455 27863
rect 25697 27829 25731 27863
rect 3709 27625 3743 27659
rect 7205 27625 7239 27659
rect 8861 27625 8895 27659
rect 9597 27625 9631 27659
rect 9689 27625 9723 27659
rect 14933 27625 14967 27659
rect 22937 27625 22971 27659
rect 24961 27625 24995 27659
rect 25395 27625 25429 27659
rect 25697 27625 25731 27659
rect 2504 27557 2538 27591
rect 3877 27557 3911 27591
rect 4077 27557 4111 27591
rect 4537 27557 4571 27591
rect 15577 27557 15611 27591
rect 16589 27557 16623 27591
rect 16789 27557 16823 27591
rect 20085 27557 20119 27591
rect 22109 27557 22143 27591
rect 22753 27557 22787 27591
rect 24409 27557 24443 27591
rect 24777 27557 24811 27591
rect 25605 27557 25639 27591
rect 4353 27489 4387 27523
rect 4629 27489 4663 27523
rect 4813 27489 4847 27523
rect 5273 27489 5307 27523
rect 5825 27489 5859 27523
rect 6081 27489 6115 27523
rect 7665 27489 7699 27523
rect 7757 27489 7791 27523
rect 8033 27489 8067 27523
rect 8309 27489 8343 27523
rect 8493 27489 8527 27523
rect 8585 27489 8619 27523
rect 8677 27489 8711 27523
rect 9873 27489 9907 27523
rect 9965 27489 9999 27523
rect 10057 27489 10091 27523
rect 10241 27489 10275 27523
rect 10517 27489 10551 27523
rect 10977 27489 11011 27523
rect 11233 27489 11267 27523
rect 12817 27489 12851 27523
rect 13073 27489 13107 27523
rect 14473 27489 14507 27523
rect 14992 27489 15026 27523
rect 17049 27489 17083 27523
rect 17693 27489 17727 27523
rect 17969 27489 18003 27523
rect 19358 27489 19392 27523
rect 19625 27489 19659 27523
rect 19901 27489 19935 27523
rect 19993 27489 20027 27523
rect 20269 27489 20303 27523
rect 21281 27489 21315 27523
rect 22017 27489 22051 27523
rect 22192 27489 22226 27523
rect 23029 27489 23063 27523
rect 24501 27489 24535 27523
rect 24593 27489 24627 27523
rect 24869 27489 24903 27523
rect 25697 27489 25731 27523
rect 25881 27489 25915 27523
rect 2237 27421 2271 27455
rect 4721 27421 4755 27455
rect 8953 27421 8987 27455
rect 21833 27421 21867 27455
rect 23121 27421 23155 27455
rect 3617 27353 3651 27387
rect 5457 27353 5491 27387
rect 12357 27353 12391 27387
rect 14197 27353 14231 27387
rect 15117 27353 15151 27387
rect 15209 27353 15243 27387
rect 22385 27353 22419 27387
rect 3893 27285 3927 27319
rect 4169 27285 4203 27319
rect 7481 27285 7515 27319
rect 7941 27285 7975 27319
rect 10425 27285 10459 27319
rect 14565 27285 14599 27319
rect 15577 27285 15611 27319
rect 15761 27285 15795 27319
rect 16773 27285 16807 27319
rect 16957 27285 16991 27319
rect 17877 27285 17911 27319
rect 18245 27285 18279 27319
rect 19717 27285 19751 27319
rect 22753 27285 22787 27319
rect 25145 27285 25179 27319
rect 25237 27285 25271 27319
rect 25421 27285 25455 27319
rect 5089 27081 5123 27115
rect 5273 27081 5307 27115
rect 5365 27081 5399 27115
rect 5549 27081 5583 27115
rect 6745 27081 6779 27115
rect 7941 27081 7975 27115
rect 8401 27081 8435 27115
rect 8953 27081 8987 27115
rect 10977 27081 11011 27115
rect 12909 27081 12943 27115
rect 17693 27081 17727 27115
rect 17969 27081 18003 27115
rect 18337 27081 18371 27115
rect 19165 27081 19199 27115
rect 20913 27081 20947 27115
rect 21649 27081 21683 27115
rect 21925 27081 21959 27115
rect 22109 27081 22143 27115
rect 22753 27081 22787 27115
rect 23397 27081 23431 27115
rect 4721 27013 4755 27047
rect 6193 27013 6227 27047
rect 7021 27013 7055 27047
rect 7481 27013 7515 27047
rect 15853 27013 15887 27047
rect 17141 27013 17175 27047
rect 18153 27013 18187 27047
rect 21833 27013 21867 27047
rect 7205 26945 7239 26979
rect 7757 26945 7791 26979
rect 8769 26945 8803 26979
rect 14197 26945 14231 26979
rect 19533 26945 19567 26979
rect 2237 26877 2271 26911
rect 6009 26877 6043 26911
rect 6929 26877 6963 26911
rect 7113 26877 7147 26911
rect 7389 26877 7423 26911
rect 8033 26877 8067 26911
rect 8585 26877 8619 26911
rect 10333 26877 10367 26911
rect 11161 26877 11195 26911
rect 11529 26877 11563 26911
rect 11621 26877 11655 26911
rect 15393 26877 15427 26911
rect 15485 26877 15519 26911
rect 17049 26877 17083 26911
rect 17233 26877 17267 26911
rect 17509 26877 17543 26911
rect 18245 26877 18279 26911
rect 18705 26877 18739 26911
rect 18889 26877 18923 26911
rect 18981 26877 19015 26911
rect 19800 26877 19834 26911
rect 21189 26877 21223 26911
rect 21373 26877 21407 26911
rect 22385 26877 22419 26911
rect 23213 26877 23247 26911
rect 2421 26809 2455 26843
rect 5517 26809 5551 26843
rect 5733 26809 5767 26843
rect 5825 26809 5859 26843
rect 10066 26809 10100 26843
rect 11253 26809 11287 26843
rect 11345 26809 11379 26843
rect 15117 26809 15151 26843
rect 16221 26809 16255 26843
rect 17325 26809 17359 26843
rect 17785 26809 17819 26843
rect 21465 26809 21499 26843
rect 21681 26809 21715 26843
rect 22293 26809 22327 26843
rect 22558 26809 22592 26843
rect 25329 26809 25363 26843
rect 2605 26741 2639 26775
rect 5089 26741 5123 26775
rect 13553 26741 13587 26775
rect 15301 26741 15335 26775
rect 15669 26741 15703 26775
rect 15761 26741 15795 26775
rect 17985 26741 18019 26775
rect 18705 26741 18739 26775
rect 21281 26741 21315 26775
rect 22093 26741 22127 26775
rect 23673 26741 23707 26775
rect 26617 26741 26651 26775
rect 6561 26537 6595 26571
rect 12633 26537 12667 26571
rect 16773 26537 16807 26571
rect 17995 26537 18029 26571
rect 21833 26537 21867 26571
rect 22845 26537 22879 26571
rect 23305 26537 23339 26571
rect 24317 26537 24351 26571
rect 25513 26537 25547 26571
rect 2605 26469 2639 26503
rect 8953 26469 8987 26503
rect 11621 26469 11655 26503
rect 13001 26469 13035 26503
rect 17785 26469 17819 26503
rect 21449 26469 21483 26503
rect 21649 26469 21683 26503
rect 21925 26469 21959 26503
rect 23949 26469 23983 26503
rect 25329 26469 25363 26503
rect 25757 26469 25791 26503
rect 25973 26469 26007 26503
rect 949 26401 983 26435
rect 1216 26401 1250 26435
rect 3065 26401 3099 26435
rect 3249 26401 3283 26435
rect 3801 26401 3835 26435
rect 4997 26401 5031 26435
rect 5089 26401 5123 26435
rect 5273 26401 5307 26435
rect 5549 26401 5583 26435
rect 6285 26401 6319 26435
rect 7205 26401 7239 26435
rect 7297 26401 7331 26435
rect 7481 26401 7515 26435
rect 7573 26401 7607 26435
rect 8217 26401 8251 26435
rect 8309 26401 8343 26435
rect 8401 26401 8435 26435
rect 8585 26401 8619 26435
rect 8861 26401 8895 26435
rect 9045 26401 9079 26435
rect 9229 26401 9263 26435
rect 10057 26401 10091 26435
rect 10609 26401 10643 26435
rect 11437 26401 11471 26435
rect 11529 26401 11563 26435
rect 11805 26401 11839 26435
rect 11897 26401 11931 26435
rect 12817 26401 12851 26435
rect 12909 26401 12943 26435
rect 13185 26401 13219 26435
rect 13369 26401 13403 26435
rect 14381 26401 14415 26435
rect 15485 26401 15519 26435
rect 15577 26401 15611 26435
rect 15761 26401 15795 26435
rect 15853 26401 15887 26435
rect 16957 26401 16991 26435
rect 17601 26401 17635 26435
rect 19542 26401 19576 26435
rect 19809 26401 19843 26435
rect 20913 26401 20947 26435
rect 21741 26401 21775 26435
rect 22017 26401 22051 26435
rect 22385 26401 22419 26435
rect 23397 26401 23431 26435
rect 23489 26401 23523 26435
rect 23765 26401 23799 26435
rect 24041 26401 24075 26435
rect 24133 26401 24167 26435
rect 26249 26401 26283 26435
rect 6101 26333 6135 26367
rect 6929 26333 6963 26367
rect 7021 26333 7055 26367
rect 9321 26333 9355 26367
rect 9873 26333 9907 26367
rect 12541 26333 12575 26367
rect 16313 26333 16347 26367
rect 24961 26333 24995 26367
rect 2329 26265 2363 26299
rect 2973 26265 3007 26299
rect 6469 26265 6503 26299
rect 7757 26265 7791 26299
rect 13921 26265 13955 26299
rect 15301 26265 15335 26299
rect 16589 26265 16623 26299
rect 17141 26265 17175 26299
rect 17509 26265 17543 26299
rect 21281 26265 21315 26299
rect 23121 26265 23155 26299
rect 23673 26265 23707 26299
rect 2421 26197 2455 26231
rect 2605 26197 2639 26231
rect 3433 26197 3467 26231
rect 3617 26197 3651 26231
rect 5457 26197 5491 26231
rect 7297 26197 7331 26231
rect 8033 26197 8067 26231
rect 8677 26197 8711 26231
rect 11253 26197 11287 26231
rect 13645 26197 13679 26231
rect 13829 26197 13863 26231
rect 14289 26197 14323 26231
rect 17969 26197 18003 26231
rect 18153 26197 18187 26231
rect 18429 26197 18463 26231
rect 20729 26197 20763 26231
rect 21465 26197 21499 26231
rect 22477 26197 22511 26231
rect 25329 26197 25363 26231
rect 25605 26197 25639 26231
rect 25789 26197 25823 26231
rect 26065 26197 26099 26231
rect 1409 25993 1443 26027
rect 2881 25993 2915 26027
rect 7297 25993 7331 26027
rect 7941 25993 7975 26027
rect 11529 25993 11563 26027
rect 14933 25993 14967 26027
rect 18245 25993 18279 26027
rect 18429 25993 18463 26027
rect 18889 25993 18923 26027
rect 21741 25993 21775 26027
rect 22477 25993 22511 26027
rect 22845 25993 22879 26027
rect 23121 25993 23155 26027
rect 23489 25993 23523 26027
rect 23949 25993 23983 26027
rect 24593 25993 24627 26027
rect 25421 25993 25455 26027
rect 25697 25993 25731 26027
rect 2605 25925 2639 25959
rect 8493 25925 8527 25959
rect 13001 25925 13035 25959
rect 7757 25857 7791 25891
rect 13277 25857 13311 25891
rect 16589 25857 16623 25891
rect 20269 25857 20303 25891
rect 25053 25857 25087 25891
rect 1593 25789 1627 25823
rect 2329 25789 2363 25823
rect 2421 25789 2455 25823
rect 3249 25789 3283 25823
rect 4997 25789 5031 25823
rect 7021 25789 7055 25823
rect 7205 25789 7239 25823
rect 7481 25789 7515 25823
rect 7573 25789 7607 25823
rect 8033 25789 8067 25823
rect 8585 25789 8619 25823
rect 8677 25789 8711 25823
rect 10149 25789 10183 25823
rect 11621 25789 11655 25823
rect 13185 25789 13219 25823
rect 13369 25789 13403 25823
rect 14105 25789 14139 25823
rect 14381 25789 14415 25823
rect 14657 25789 14691 25823
rect 14749 25789 14783 25823
rect 17877 25789 17911 25823
rect 18061 25789 18095 25823
rect 18521 25789 18555 25823
rect 18705 25789 18739 25823
rect 21925 25789 21959 25823
rect 22109 25789 22143 25823
rect 22201 25789 22235 25823
rect 22385 25789 22419 25823
rect 23029 25789 23063 25823
rect 23857 25789 23891 25823
rect 24041 25789 24075 25823
rect 24501 25789 24535 25823
rect 24777 25789 24811 25823
rect 24961 25789 24995 25823
rect 27077 25789 27111 25823
rect 2697 25721 2731 25755
rect 3516 25721 3550 25755
rect 5264 25721 5298 25755
rect 8922 25721 8956 25755
rect 10416 25721 10450 25755
rect 11888 25721 11922 25755
rect 14565 25721 14599 25755
rect 16322 25721 16356 25755
rect 20536 25721 20570 25755
rect 26810 25721 26844 25755
rect 2897 25653 2931 25687
rect 3065 25653 3099 25687
rect 4629 25653 4663 25687
rect 6377 25653 6411 25687
rect 6469 25653 6503 25687
rect 10057 25653 10091 25687
rect 13553 25653 13587 25687
rect 15209 25653 15243 25687
rect 21649 25653 21683 25687
rect 24317 25653 24351 25687
rect 25421 25653 25455 25687
rect 25605 25653 25639 25687
rect 3801 25449 3835 25483
rect 5181 25449 5215 25483
rect 9321 25449 9355 25483
rect 11805 25449 11839 25483
rect 13645 25449 13679 25483
rect 13921 25449 13955 25483
rect 14013 25449 14047 25483
rect 24317 25449 24351 25483
rect 24869 25449 24903 25483
rect 26893 25449 26927 25483
rect 3617 25381 3651 25415
rect 8186 25381 8220 25415
rect 12081 25381 12115 25415
rect 13737 25381 13771 25415
rect 14933 25381 14967 25415
rect 15393 25381 15427 25415
rect 15593 25381 15627 25415
rect 18337 25381 18371 25415
rect 19165 25381 19199 25415
rect 20821 25381 20855 25415
rect 26433 25381 26467 25415
rect 1225 25313 1259 25347
rect 2237 25313 2271 25347
rect 2421 25313 2455 25347
rect 3249 25313 3283 25347
rect 4537 25313 4571 25347
rect 4721 25313 4755 25347
rect 4813 25313 4847 25347
rect 4905 25313 4939 25347
rect 7021 25313 7055 25347
rect 11989 25313 12023 25347
rect 12173 25313 12207 25347
rect 12357 25313 12391 25347
rect 13185 25313 13219 25347
rect 14105 25313 14139 25347
rect 16681 25313 16715 25347
rect 16865 25313 16899 25347
rect 18429 25313 18463 25347
rect 19257 25313 19291 25347
rect 19717 25313 19751 25347
rect 20269 25313 20303 25347
rect 20637 25313 20671 25347
rect 20729 25313 20763 25347
rect 21005 25313 21039 25347
rect 21281 25313 21315 25347
rect 25982 25313 26016 25347
rect 26249 25313 26283 25347
rect 26617 25313 26651 25347
rect 27077 25313 27111 25347
rect 7941 25245 7975 25279
rect 9965 25245 9999 25279
rect 14289 25245 14323 25279
rect 17969 25245 18003 25279
rect 21925 25245 21959 25279
rect 22569 25245 22603 25279
rect 23857 25245 23891 25279
rect 14565 25177 14599 25211
rect 22937 25177 22971 25211
rect 24225 25177 24259 25211
rect 1041 25109 1075 25143
rect 2605 25109 2639 25143
rect 3617 25109 3651 25143
rect 6929 25109 6963 25143
rect 9413 25109 9447 25143
rect 13461 25109 13495 25143
rect 14933 25109 14967 25143
rect 15117 25109 15151 25143
rect 15577 25109 15611 25143
rect 15761 25109 15795 25143
rect 16681 25109 16715 25143
rect 18153 25109 18187 25143
rect 20453 25109 20487 25143
rect 23029 25109 23063 25143
rect 26801 25109 26835 25143
rect 2237 24905 2271 24939
rect 2513 24905 2547 24939
rect 3433 24905 3467 24939
rect 6377 24905 6411 24939
rect 7297 24905 7331 24939
rect 8401 24905 8435 24939
rect 14013 24905 14047 24939
rect 14381 24905 14415 24939
rect 14933 24905 14967 24939
rect 15025 24905 15059 24939
rect 15209 24905 15243 24939
rect 16221 24905 16255 24939
rect 16405 24905 16439 24939
rect 24593 24905 24627 24939
rect 2329 24837 2363 24871
rect 2881 24837 2915 24871
rect 3249 24837 3283 24871
rect 4537 24837 4571 24871
rect 5733 24837 5767 24871
rect 15669 24837 15703 24871
rect 21557 24837 21591 24871
rect 22017 24837 22051 24871
rect 22753 24837 22787 24871
rect 23581 24837 23615 24871
rect 5181 24769 5215 24803
rect 6285 24769 6319 24803
rect 9781 24769 9815 24803
rect 11713 24769 11747 24803
rect 16589 24769 16623 24803
rect 16681 24769 16715 24803
rect 17049 24769 17083 24803
rect 20177 24769 20211 24803
rect 22109 24769 22143 24803
rect 23397 24769 23431 24803
rect 857 24701 891 24735
rect 4721 24701 4755 24735
rect 5825 24701 5859 24735
rect 6804 24701 6838 24735
rect 7021 24701 7055 24735
rect 7573 24701 7607 24735
rect 7757 24701 7791 24735
rect 10057 24701 10091 24735
rect 10149 24701 10183 24735
rect 10425 24701 10459 24735
rect 10517 24701 10551 24735
rect 13921 24701 13955 24735
rect 14749 24701 14783 24735
rect 15485 24701 15519 24735
rect 16037 24701 16071 24735
rect 16313 24701 16347 24735
rect 16773 24701 16807 24735
rect 17325 24701 17359 24735
rect 17417 24701 17451 24735
rect 18705 24701 18739 24735
rect 20444 24701 20478 24735
rect 22661 24701 22695 24735
rect 23029 24701 23063 24735
rect 23121 24701 23155 24735
rect 23489 24701 23523 24735
rect 24041 24701 24075 24735
rect 24225 24701 24259 24735
rect 24317 24701 24351 24735
rect 24869 24701 24903 24735
rect 25053 24701 25087 24735
rect 25145 24701 25179 24735
rect 25237 24701 25271 24735
rect 25605 24701 25639 24735
rect 3387 24667 3421 24701
rect 1124 24633 1158 24667
rect 3617 24633 3651 24667
rect 5089 24633 5123 24667
rect 5365 24633 5399 24667
rect 5549 24633 5583 24667
rect 7665 24633 7699 24667
rect 9514 24633 9548 24667
rect 10241 24633 10275 24667
rect 11980 24633 12014 24667
rect 14565 24633 14599 24667
rect 15393 24633 15427 24667
rect 16957 24633 16991 24667
rect 18950 24633 18984 24667
rect 21649 24633 21683 24667
rect 24561 24633 24595 24667
rect 24777 24633 24811 24667
rect 25850 24633 25884 24667
rect 2513 24565 2547 24599
rect 4813 24565 4847 24599
rect 4905 24565 4939 24599
rect 5457 24565 5491 24599
rect 5917 24565 5951 24599
rect 6745 24565 6779 24599
rect 6929 24565 6963 24599
rect 7481 24565 7515 24599
rect 9873 24565 9907 24599
rect 11161 24565 11195 24599
rect 13093 24565 13127 24599
rect 15193 24565 15227 24599
rect 15853 24565 15887 24599
rect 17601 24565 17635 24599
rect 20085 24565 20119 24599
rect 22937 24565 22971 24599
rect 23857 24565 23891 24599
rect 24409 24565 24443 24599
rect 25513 24565 25547 24599
rect 26985 24565 27019 24599
rect 4997 24361 5031 24395
rect 7665 24361 7699 24395
rect 8677 24361 8711 24395
rect 9413 24361 9447 24395
rect 10977 24361 11011 24395
rect 11713 24361 11747 24395
rect 14105 24361 14139 24395
rect 14657 24361 14691 24395
rect 15117 24361 15151 24395
rect 15485 24361 15519 24395
rect 16306 24361 16340 24395
rect 16589 24361 16623 24395
rect 17233 24361 17267 24395
rect 18061 24361 18095 24395
rect 18245 24361 18279 24395
rect 18889 24361 18923 24395
rect 23029 24361 23063 24395
rect 23942 24361 23976 24395
rect 25513 24361 25547 24395
rect 26433 24361 26467 24395
rect 2053 24293 2087 24327
rect 2513 24293 2547 24327
rect 2973 24293 3007 24327
rect 5641 24293 5675 24327
rect 10548 24293 10582 24327
rect 12909 24293 12943 24327
rect 13277 24293 13311 24327
rect 13737 24293 13771 24327
rect 13942 24293 13976 24327
rect 16405 24293 16439 24327
rect 19349 24293 19383 24327
rect 23857 24293 23891 24327
rect 24961 24293 24995 24327
rect 25161 24293 25195 24327
rect 1225 24225 1259 24259
rect 1869 24225 1903 24259
rect 2145 24225 2179 24259
rect 3138 24225 3172 24259
rect 3249 24225 3283 24259
rect 3516 24225 3550 24259
rect 4905 24225 4939 24259
rect 5273 24225 5307 24259
rect 6193 24225 6227 24259
rect 6285 24225 6319 24259
rect 6561 24225 6595 24259
rect 6837 24225 6871 24259
rect 7021 24225 7055 24259
rect 7113 24225 7147 24259
rect 7205 24225 7239 24259
rect 7389 24225 7423 24259
rect 7606 24225 7640 24259
rect 8033 24225 8067 24259
rect 8217 24225 8251 24259
rect 8401 24225 8435 24259
rect 8861 24225 8895 24259
rect 8953 24225 8987 24259
rect 9045 24225 9079 24259
rect 9229 24225 9263 24259
rect 10793 24225 10827 24259
rect 11897 24225 11931 24259
rect 11989 24225 12023 24259
rect 12081 24225 12115 24259
rect 12265 24225 12299 24259
rect 12725 24225 12759 24259
rect 12817 24225 12851 24259
rect 13001 24225 13035 24259
rect 14197 24225 14231 24259
rect 15025 24225 15059 24259
rect 15209 24225 15243 24259
rect 15577 24225 15611 24259
rect 16129 24225 16163 24259
rect 16221 24225 16255 24259
rect 16773 24225 16807 24259
rect 16865 24225 16899 24259
rect 16957 24225 16991 24259
rect 17141 24225 17175 24259
rect 17509 24225 17543 24259
rect 17601 24225 17635 24259
rect 17693 24225 17727 24259
rect 17877 24225 17911 24259
rect 18242 24225 18276 24259
rect 18613 24225 18647 24259
rect 19717 24225 19751 24259
rect 19984 24225 20018 24259
rect 22017 24225 22051 24259
rect 22569 24225 22603 24259
rect 23121 24225 23155 24259
rect 23213 24225 23247 24259
rect 23397 24225 23431 24259
rect 23765 24225 23799 24259
rect 24041 24225 24075 24259
rect 24685 24225 24719 24259
rect 25605 24225 25639 24259
rect 25973 24225 26007 24259
rect 26157 24225 26191 24259
rect 26985 24225 27019 24259
rect 1685 24157 1719 24191
rect 8125 24157 8159 24191
rect 11529 24157 11563 24191
rect 12633 24157 12667 24191
rect 14749 24157 14783 24191
rect 18705 24157 18739 24191
rect 21833 24157 21867 24191
rect 22477 24157 22511 24191
rect 23581 24157 23615 24191
rect 2697 24089 2731 24123
rect 4629 24089 4663 24123
rect 6009 24089 6043 24123
rect 8309 24089 8343 24123
rect 13645 24089 13679 24123
rect 14565 24089 14599 24123
rect 14841 24089 14875 24123
rect 15669 24089 15703 24123
rect 19073 24089 19107 24123
rect 21097 24089 21131 24123
rect 25329 24089 25363 24123
rect 1041 24021 1075 24055
rect 2513 24021 2547 24055
rect 2789 24021 2823 24055
rect 6469 24021 6503 24055
rect 6653 24021 6687 24055
rect 7481 24021 7515 24055
rect 13093 24021 13127 24055
rect 13277 24021 13311 24055
rect 13921 24021 13955 24055
rect 21281 24021 21315 24055
rect 22109 24021 22143 24055
rect 22845 24021 22879 24055
rect 24593 24021 24627 24055
rect 25145 24021 25179 24055
rect 26065 24021 26099 24055
rect 2237 23817 2271 23851
rect 3525 23817 3559 23851
rect 5181 23817 5215 23851
rect 8125 23817 8159 23851
rect 11345 23817 11379 23851
rect 12909 23817 12943 23851
rect 14473 23817 14507 23851
rect 14841 23817 14875 23851
rect 15761 23817 15795 23851
rect 18981 23817 19015 23851
rect 19993 23817 20027 23851
rect 24593 23817 24627 23851
rect 5089 23749 5123 23783
rect 7665 23749 7699 23783
rect 15209 23749 15243 23783
rect 9137 23681 9171 23715
rect 9689 23681 9723 23715
rect 23029 23681 23063 23715
rect 857 23613 891 23647
rect 1124 23613 1158 23647
rect 3341 23613 3375 23647
rect 4721 23613 4755 23647
rect 5554 23613 5588 23647
rect 7297 23613 7331 23647
rect 7389 23613 7423 23647
rect 7757 23613 7791 23647
rect 8217 23613 8251 23647
rect 8493 23613 8527 23647
rect 8677 23613 8711 23647
rect 8861 23613 8895 23647
rect 9965 23613 9999 23647
rect 11437 23613 11471 23647
rect 13093 23613 13127 23647
rect 14105 23613 14139 23647
rect 14289 23613 14323 23647
rect 14473 23613 14507 23647
rect 14749 23613 14783 23647
rect 15301 23613 15335 23647
rect 15577 23613 15611 23647
rect 18705 23613 18739 23647
rect 18797 23613 18831 23647
rect 18981 23613 19015 23647
rect 20177 23613 20211 23647
rect 20545 23613 20579 23647
rect 21833 23613 21867 23647
rect 22017 23613 22051 23647
rect 24777 23613 24811 23647
rect 24869 23613 24903 23647
rect 24961 23613 24995 23647
rect 25697 23613 25731 23647
rect 2697 23545 2731 23579
rect 2881 23545 2915 23579
rect 4813 23545 4847 23579
rect 5181 23545 5215 23579
rect 5365 23545 5399 23579
rect 5457 23545 5491 23579
rect 7481 23545 7515 23579
rect 8769 23545 8803 23579
rect 10210 23545 10244 23579
rect 11704 23545 11738 23579
rect 20269 23545 20303 23579
rect 20361 23545 20395 23579
rect 22477 23545 22511 23579
rect 25942 23545 25976 23579
rect 3065 23477 3099 23511
rect 4537 23477 4571 23511
rect 4905 23477 4939 23511
rect 7113 23477 7147 23511
rect 7849 23477 7883 23511
rect 9045 23477 9079 23511
rect 12817 23477 12851 23511
rect 13553 23477 13587 23511
rect 15393 23477 15427 23511
rect 21925 23477 21959 23511
rect 27077 23477 27111 23511
rect 2605 23273 2639 23307
rect 3065 23273 3099 23307
rect 3249 23273 3283 23307
rect 3509 23273 3543 23307
rect 5089 23273 5123 23307
rect 8125 23273 8159 23307
rect 14749 23273 14783 23307
rect 15301 23273 15335 23307
rect 16129 23273 16163 23307
rect 19349 23273 19383 23307
rect 21833 23273 21867 23307
rect 23305 23273 23339 23307
rect 23765 23273 23799 23307
rect 24501 23273 24535 23307
rect 25773 23273 25807 23307
rect 3709 23205 3743 23239
rect 4813 23205 4847 23239
rect 7113 23205 7147 23239
rect 7297 23205 7331 23239
rect 7481 23205 7515 23239
rect 9238 23205 9272 23239
rect 9689 23205 9723 23239
rect 11529 23205 11563 23239
rect 11621 23205 11655 23239
rect 12173 23205 12207 23239
rect 17242 23205 17276 23239
rect 22170 23205 22204 23239
rect 25513 23205 25547 23239
rect 25973 23205 26007 23239
rect 26617 23205 26651 23239
rect 2421 23137 2455 23171
rect 3985 23137 4019 23171
rect 4721 23137 4755 23171
rect 4905 23137 4939 23171
rect 5825 23137 5859 23171
rect 6837 23137 6871 23171
rect 7205 23137 7239 23171
rect 9873 23137 9907 23171
rect 9965 23137 9999 23171
rect 10149 23137 10183 23171
rect 10333 23137 10367 23171
rect 10425 23137 10459 23171
rect 10517 23137 10551 23171
rect 11437 23137 11471 23171
rect 11805 23137 11839 23171
rect 12081 23137 12115 23171
rect 12265 23137 12299 23171
rect 12449 23137 12483 23171
rect 14289 23137 14323 23171
rect 14841 23137 14875 23171
rect 18225 23137 18259 23171
rect 19993 23137 20027 23171
rect 20637 23137 20671 23171
rect 21465 23137 21499 23171
rect 23673 23137 23707 23171
rect 23857 23137 23891 23171
rect 23949 23137 23983 23171
rect 24133 23137 24167 23171
rect 24225 23137 24259 23171
rect 24317 23137 24351 23171
rect 25145 23137 25179 23171
rect 25421 23137 25455 23171
rect 26249 23137 26283 23171
rect 26433 23137 26467 23171
rect 26893 23137 26927 23171
rect 2237 23069 2271 23103
rect 7113 23069 7147 23103
rect 9505 23069 9539 23103
rect 12541 23069 12575 23103
rect 13093 23069 13127 23103
rect 17509 23069 17543 23103
rect 17969 23069 18003 23103
rect 20361 23069 20395 23103
rect 21373 23069 21407 23103
rect 21925 23069 21959 23103
rect 25053 23069 25087 23103
rect 2697 23001 2731 23035
rect 3341 23001 3375 23035
rect 4537 23001 4571 23035
rect 6929 23001 6963 23035
rect 15117 23001 15151 23035
rect 26801 23001 26835 23035
rect 3065 22933 3099 22967
rect 3525 22933 3559 22967
rect 3801 22933 3835 22967
rect 5917 22933 5951 22967
rect 6285 22933 6319 22967
rect 7481 22933 7515 22967
rect 10701 22933 10735 22967
rect 11253 22933 11287 22967
rect 11897 22933 11931 22967
rect 14381 22933 14415 22967
rect 19441 22933 19475 22967
rect 24869 22933 24903 22967
rect 25605 22933 25639 22967
rect 25789 22933 25823 22967
rect 26157 22933 26191 22967
rect 26985 22933 27019 22967
rect 2237 22729 2271 22763
rect 2513 22729 2547 22763
rect 6745 22729 6779 22763
rect 9137 22729 9171 22763
rect 13737 22729 13771 22763
rect 14013 22729 14047 22763
rect 17233 22729 17267 22763
rect 17877 22729 17911 22763
rect 18797 22729 18831 22763
rect 19533 22729 19567 22763
rect 23857 22729 23891 22763
rect 25237 22729 25271 22763
rect 25605 22729 25639 22763
rect 25697 22729 25731 22763
rect 2881 22661 2915 22695
rect 4813 22661 4847 22695
rect 6469 22661 6503 22695
rect 13921 22661 13955 22695
rect 23305 22661 23339 22695
rect 857 22593 891 22627
rect 5181 22593 5215 22627
rect 6193 22593 6227 22627
rect 9505 22593 9539 22627
rect 12633 22593 12667 22627
rect 16497 22593 16531 22627
rect 17141 22593 17175 22627
rect 21925 22593 21959 22627
rect 3433 22525 3467 22559
rect 5089 22525 5123 22559
rect 5273 22525 5307 22559
rect 5365 22525 5399 22559
rect 5825 22525 5859 22559
rect 6101 22525 6135 22559
rect 7021 22525 7055 22559
rect 7297 22525 7331 22559
rect 7481 22525 7515 22559
rect 7573 22525 7607 22559
rect 9321 22525 9355 22559
rect 9597 22525 9631 22559
rect 10241 22525 10275 22559
rect 12541 22525 12575 22559
rect 12725 22525 12759 22559
rect 12909 22525 12943 22559
rect 14013 22525 14047 22559
rect 14105 22525 14139 22559
rect 17417 22525 17451 22559
rect 17785 22525 17819 22559
rect 18061 22525 18095 22559
rect 18153 22525 18187 22559
rect 18429 22525 18463 22559
rect 18889 22525 18923 22559
rect 19073 22525 19107 22559
rect 19165 22525 19199 22559
rect 19349 22525 19383 22559
rect 19809 22525 19843 22559
rect 21281 22525 21315 22559
rect 21557 22525 21591 22559
rect 21649 22525 21683 22559
rect 24409 22525 24443 22559
rect 24593 22525 24627 22559
rect 24777 22525 24811 22559
rect 24869 22525 24903 22559
rect 24961 22525 24995 22559
rect 25421 22525 25455 22559
rect 27077 22525 27111 22559
rect 1124 22457 1158 22491
rect 3700 22457 3734 22491
rect 6310 22457 6344 22491
rect 7389 22457 7423 22491
rect 13553 22457 13587 22491
rect 14289 22457 14323 22491
rect 17509 22457 17543 22491
rect 17601 22457 17635 22491
rect 18245 22457 18279 22491
rect 20054 22457 20088 22491
rect 21465 22457 21499 22491
rect 22170 22457 22204 22491
rect 26810 22457 26844 22491
rect 2329 22389 2363 22423
rect 2513 22389 2547 22423
rect 4905 22389 4939 22423
rect 6561 22389 6595 22423
rect 7113 22389 7147 22423
rect 9689 22389 9723 22423
rect 11069 22389 11103 22423
rect 13753 22389 13787 22423
rect 21189 22389 21223 22423
rect 21833 22389 21867 22423
rect 1225 22185 1259 22219
rect 2421 22185 2455 22219
rect 3893 22185 3927 22219
rect 4077 22185 4111 22219
rect 5641 22185 5675 22219
rect 6285 22185 6319 22219
rect 6469 22185 6503 22219
rect 7573 22185 7607 22219
rect 10149 22185 10183 22219
rect 12817 22185 12851 22219
rect 14565 22185 14599 22219
rect 19625 22185 19659 22219
rect 19901 22185 19935 22219
rect 26893 22185 26927 22219
rect 2605 22117 2639 22151
rect 2789 22117 2823 22151
rect 11682 22117 11716 22151
rect 18061 22117 18095 22151
rect 26433 22117 26467 22151
rect 26649 22117 26683 22151
rect 1409 22049 1443 22083
rect 3525 22049 3559 22083
rect 5181 22049 5215 22083
rect 5825 22049 5859 22083
rect 6377 22049 6411 22083
rect 6653 22049 6687 22083
rect 7113 22049 7147 22083
rect 7481 22049 7515 22083
rect 7757 22049 7791 22083
rect 7941 22049 7975 22083
rect 8933 22049 8967 22083
rect 11437 22049 11471 22083
rect 14206 22049 14240 22083
rect 15689 22049 15723 22083
rect 15945 22049 15979 22083
rect 16405 22049 16439 22083
rect 16589 22049 16623 22083
rect 16681 22049 16715 22083
rect 16865 22049 16899 22083
rect 16957 22049 16991 22083
rect 17141 22049 17175 22083
rect 17877 22049 17911 22083
rect 17969 22049 18003 22083
rect 18245 22049 18279 22083
rect 18613 22049 18647 22083
rect 19441 22049 19475 22083
rect 19625 22049 19659 22083
rect 20061 22049 20095 22083
rect 20177 22049 20211 22083
rect 20269 22049 20303 22083
rect 20453 22049 20487 22083
rect 21281 22049 21315 22083
rect 21833 22049 21867 22083
rect 24869 22049 24903 22083
rect 24961 22049 24995 22083
rect 25697 22049 25731 22083
rect 26065 22049 26099 22083
rect 26157 22049 26191 22083
rect 27077 22049 27111 22083
rect 7297 21981 7331 22015
rect 8677 21981 8711 22015
rect 10701 21981 10735 22015
rect 14473 21981 14507 22015
rect 16129 21981 16163 22015
rect 17049 21981 17083 22015
rect 19257 21981 19291 22015
rect 22937 21981 22971 22015
rect 23581 21981 23615 22015
rect 25513 21981 25547 22015
rect 5457 21913 5491 21947
rect 6653 21913 6687 21947
rect 7113 21913 7147 21947
rect 10057 21913 10091 21947
rect 16773 21913 16807 21947
rect 23029 21913 23063 21947
rect 24777 21913 24811 21947
rect 26801 21913 26835 21947
rect 3893 21845 3927 21879
rect 6101 21845 6135 21879
rect 13093 21845 13127 21879
rect 16221 21845 16255 21879
rect 17693 21845 17727 21879
rect 22293 21845 22327 21879
rect 25881 21845 25915 21879
rect 26617 21845 26651 21879
rect 3893 21641 3927 21675
rect 4261 21641 4295 21675
rect 7849 21641 7883 21675
rect 8769 21641 8803 21675
rect 12081 21641 12115 21675
rect 13645 21641 13679 21675
rect 14197 21641 14231 21675
rect 16037 21641 16071 21675
rect 19901 21641 19935 21675
rect 24501 21641 24535 21675
rect 25053 21641 25087 21675
rect 26617 21641 26651 21675
rect 1317 21573 1351 21607
rect 6929 21573 6963 21607
rect 10057 21573 10091 21607
rect 19257 21573 19291 21607
rect 23213 21573 23247 21607
rect 24961 21573 24995 21607
rect 1501 21505 1535 21539
rect 1685 21505 1719 21539
rect 14841 21505 14875 21539
rect 15853 21505 15887 21539
rect 19165 21505 19199 21539
rect 23949 21505 23983 21539
rect 1041 21437 1075 21471
rect 1409 21437 1443 21471
rect 2329 21437 2363 21471
rect 2513 21437 2547 21471
rect 3525 21437 3559 21471
rect 3801 21437 3835 21471
rect 3893 21437 3927 21471
rect 3985 21437 4019 21471
rect 4905 21437 4939 21471
rect 4997 21437 5031 21471
rect 7113 21437 7147 21471
rect 7389 21437 7423 21471
rect 7941 21437 7975 21471
rect 8953 21437 8987 21471
rect 9137 21437 9171 21471
rect 9321 21437 9355 21471
rect 11170 21437 11204 21471
rect 11437 21437 11471 21471
rect 12265 21437 12299 21471
rect 12449 21437 12483 21471
rect 12541 21437 12575 21471
rect 13829 21437 13863 21471
rect 14013 21437 14047 21471
rect 14105 21437 14139 21471
rect 14381 21437 14415 21471
rect 15485 21437 15519 21471
rect 15761 21437 15795 21471
rect 18061 21437 18095 21471
rect 19441 21437 19475 21471
rect 19717 21437 19751 21471
rect 19901 21437 19935 21471
rect 21189 21437 21223 21471
rect 21373 21437 21407 21471
rect 21557 21437 21591 21471
rect 21833 21437 21867 21471
rect 23489 21437 23523 21471
rect 23581 21437 23615 21471
rect 23857 21437 23891 21471
rect 24376 21437 24410 21471
rect 25329 21437 25363 21471
rect 1317 21369 1351 21403
rect 1685 21369 1719 21403
rect 3709 21369 3743 21403
rect 5181 21369 5215 21403
rect 7297 21369 7331 21403
rect 9045 21369 9079 21403
rect 17816 21369 17850 21403
rect 19625 21369 19659 21403
rect 21465 21369 21499 21403
rect 22078 21369 22112 21403
rect 24593 21369 24627 21403
rect 1133 21301 1167 21335
rect 1777 21301 1811 21335
rect 2697 21301 2731 21335
rect 3341 21301 3375 21335
rect 4905 21301 4939 21335
rect 7481 21301 7515 21335
rect 16681 21301 16715 21335
rect 21741 21301 21775 21335
rect 24317 21301 24351 21335
rect 4997 21097 5031 21131
rect 5457 21097 5491 21131
rect 7113 21097 7147 21131
rect 7849 21097 7883 21131
rect 11161 21097 11195 21131
rect 14013 21097 14047 21131
rect 19349 21097 19383 21131
rect 23305 21097 23339 21131
rect 24041 21097 24075 21131
rect 24869 21097 24903 21131
rect 26433 21097 26467 21131
rect 26985 21097 27019 21131
rect 3525 21029 3559 21063
rect 7690 21029 7724 21063
rect 14197 21029 14231 21063
rect 14565 21029 14599 21063
rect 18214 21029 18248 21063
rect 22170 21029 22204 21063
rect 24225 21029 24259 21063
rect 25982 21029 26016 21063
rect 1777 20961 1811 20995
rect 3873 20961 3907 20995
rect 5319 20961 5353 20995
rect 5549 20961 5583 20995
rect 7205 20961 7239 20995
rect 7481 20961 7515 20995
rect 9065 20961 9099 20995
rect 10526 20961 10560 20995
rect 10977 20961 11011 20995
rect 12173 20961 12207 20995
rect 12265 20961 12299 20995
rect 12449 20961 12483 20995
rect 12725 20961 12759 20995
rect 13461 20961 13495 20995
rect 15117 20961 15151 20995
rect 15301 20961 15335 20995
rect 15393 20961 15427 20995
rect 17877 20961 17911 20995
rect 19625 20961 19659 20995
rect 20729 20961 20763 20995
rect 21281 20961 21315 20995
rect 21465 20961 21499 20995
rect 21557 20961 21591 20995
rect 21649 20961 21683 20995
rect 23949 20961 23983 20995
rect 26249 20961 26283 20995
rect 26617 20961 26651 20995
rect 26801 20961 26835 20995
rect 26893 20961 26927 20995
rect 27077 20961 27111 20995
rect 1593 20893 1627 20927
rect 3617 20893 3651 20927
rect 6653 20893 6687 20927
rect 7573 20893 7607 20927
rect 9321 20893 9355 20927
rect 10793 20893 10827 20927
rect 13737 20893 13771 20927
rect 14933 20893 14967 20927
rect 17969 20893 18003 20927
rect 21925 20893 21959 20927
rect 7021 20825 7055 20859
rect 15577 20825 15611 20859
rect 21833 20825 21867 20859
rect 24225 20825 24259 20859
rect 1041 20757 1075 20791
rect 5089 20757 5123 20791
rect 7941 20757 7975 20791
rect 9413 20757 9447 20791
rect 12541 20757 12575 20791
rect 13829 20757 13863 20791
rect 16405 20757 16439 20791
rect 19441 20757 19475 20791
rect 20913 20757 20947 20791
rect 2237 20553 2271 20587
rect 2881 20553 2915 20587
rect 3433 20553 3467 20587
rect 6929 20553 6963 20587
rect 7389 20553 7423 20587
rect 7757 20553 7791 20587
rect 14565 20553 14599 20587
rect 18153 20553 18187 20587
rect 3065 20485 3099 20519
rect 5089 20485 5123 20519
rect 3709 20417 3743 20451
rect 8401 20417 8435 20451
rect 9413 20417 9447 20451
rect 10333 20417 10367 20451
rect 11805 20417 11839 20451
rect 14289 20417 14323 20451
rect 16865 20417 16899 20451
rect 857 20349 891 20383
rect 1124 20349 1158 20383
rect 2513 20349 2547 20383
rect 5273 20349 5307 20383
rect 5457 20349 5491 20383
rect 5549 20349 5583 20383
rect 7849 20349 7883 20383
rect 12072 20349 12106 20383
rect 13645 20349 13679 20383
rect 13737 20349 13771 20383
rect 14105 20349 14139 20383
rect 16221 20349 16255 20383
rect 17509 20349 17543 20383
rect 17601 20349 17635 20383
rect 17785 20349 17819 20383
rect 17877 20349 17911 20383
rect 17969 20349 18003 20383
rect 18889 20349 18923 20383
rect 20545 20349 20579 20383
rect 20729 20349 20763 20383
rect 22026 20349 22060 20383
rect 22293 20349 22327 20383
rect 23673 20349 23707 20383
rect 25697 20349 25731 20383
rect 14611 20315 14645 20349
rect 3249 20281 3283 20315
rect 3449 20281 3483 20315
rect 3976 20281 4010 20315
rect 5365 20281 5399 20315
rect 5794 20281 5828 20315
rect 10600 20281 10634 20315
rect 14381 20281 14415 20315
rect 15954 20281 15988 20315
rect 19156 20281 19190 20315
rect 20361 20281 20395 20315
rect 25942 20281 25976 20315
rect 2881 20213 2915 20247
rect 3617 20213 3651 20247
rect 9045 20213 9079 20247
rect 10057 20213 10091 20247
rect 11713 20213 11747 20247
rect 13185 20213 13219 20247
rect 14749 20213 14783 20247
rect 14841 20213 14875 20247
rect 20269 20213 20303 20247
rect 20913 20213 20947 20247
rect 23489 20213 23523 20247
rect 27077 20213 27111 20247
rect 3893 20009 3927 20043
rect 4337 20009 4371 20043
rect 5365 20009 5399 20043
rect 7665 20009 7699 20043
rect 9229 20009 9263 20043
rect 9321 20009 9355 20043
rect 10425 20009 10459 20043
rect 11069 20009 11103 20043
rect 12633 20009 12667 20043
rect 13093 20009 13127 20043
rect 15209 20009 15243 20043
rect 15577 20009 15611 20043
rect 17141 20009 17175 20043
rect 19441 20009 19475 20043
rect 19809 20009 19843 20043
rect 21281 20009 21315 20043
rect 4537 19941 4571 19975
rect 9597 19941 9631 19975
rect 11345 19941 11379 19975
rect 15669 19941 15703 19975
rect 17478 19941 17512 19975
rect 22937 19941 22971 19975
rect 1409 19873 1443 19907
rect 4077 19873 4111 19907
rect 4997 19873 5031 19907
rect 6101 19873 6135 19907
rect 6929 19873 6963 19907
rect 8125 19873 8159 19907
rect 8677 19873 8711 19907
rect 8861 19873 8895 19907
rect 8953 19873 8987 19907
rect 9045 19873 9079 19907
rect 9505 19873 9539 19907
rect 9689 19873 9723 19907
rect 9873 19873 9907 19907
rect 10793 19873 10827 19907
rect 11253 19873 11287 19907
rect 11437 19873 11471 19907
rect 11621 19873 11655 19907
rect 11713 19873 11747 19907
rect 12357 19873 12391 19907
rect 13001 19873 13035 19907
rect 13737 19873 13771 19907
rect 14197 19873 14231 19907
rect 14876 19873 14910 19907
rect 16313 19873 16347 19907
rect 16957 19873 16991 19907
rect 19349 19873 19383 19907
rect 20085 19873 20119 19907
rect 20545 19873 20579 19907
rect 20821 19873 20855 19907
rect 20913 19873 20947 19907
rect 21097 19873 21131 19907
rect 21649 19873 21683 19907
rect 22201 19873 22235 19907
rect 27077 19873 27111 19907
rect 5089 19805 5123 19839
rect 6193 19805 6227 19839
rect 7573 19805 7607 19839
rect 9965 19805 9999 19839
rect 13185 19805 13219 19839
rect 15761 19805 15795 19839
rect 17233 19805 17267 19839
rect 19257 19805 19291 19839
rect 20269 19805 20303 19839
rect 21741 19805 21775 19839
rect 21833 19805 21867 19839
rect 4169 19737 4203 19771
rect 10333 19737 10367 19771
rect 10609 19737 10643 19771
rect 1225 19669 1259 19703
rect 4353 19669 4387 19703
rect 6377 19669 6411 19703
rect 7849 19669 7883 19703
rect 14657 19669 14691 19703
rect 16129 19669 16163 19703
rect 18613 19669 18647 19703
rect 19901 19669 19935 19703
rect 20361 19669 20395 19703
rect 22293 19669 22327 19703
rect 24409 19669 24443 19703
rect 26433 19669 26467 19703
rect 9229 19465 9263 19499
rect 12541 19465 12575 19499
rect 14105 19465 14139 19499
rect 14289 19465 14323 19499
rect 15761 19465 15795 19499
rect 17325 19465 17359 19499
rect 20085 19465 20119 19499
rect 23489 19465 23523 19499
rect 23673 19465 23707 19499
rect 25237 19465 25271 19499
rect 25053 19397 25087 19431
rect 14657 19329 14691 19363
rect 14933 19329 14967 19363
rect 15393 19329 15427 19363
rect 15853 19329 15887 19363
rect 17877 19329 17911 19363
rect 18521 19329 18555 19363
rect 21189 19329 21223 19363
rect 22109 19329 22143 19363
rect 24593 19329 24627 19363
rect 857 19261 891 19295
rect 1124 19261 1158 19295
rect 2605 19261 2639 19295
rect 2789 19261 2823 19295
rect 3525 19261 3559 19295
rect 4077 19261 4111 19295
rect 4353 19261 4387 19295
rect 4629 19261 4663 19295
rect 4721 19261 4755 19295
rect 5825 19261 5859 19295
rect 7665 19261 7699 19295
rect 8585 19261 8619 19295
rect 8677 19261 8711 19295
rect 8769 19261 8803 19295
rect 8861 19261 8895 19295
rect 9597 19261 9631 19295
rect 9781 19261 9815 19295
rect 9965 19261 9999 19295
rect 10425 19261 10459 19295
rect 10517 19261 10551 19295
rect 10885 19261 10919 19295
rect 11161 19261 11195 19295
rect 11805 19261 11839 19295
rect 11897 19261 11931 19295
rect 12265 19261 12299 19295
rect 12725 19261 12759 19295
rect 12909 19261 12943 19295
rect 12997 19261 13031 19295
rect 13645 19261 13679 19295
rect 13921 19261 13955 19295
rect 15209 19261 15243 19295
rect 15577 19261 15611 19295
rect 16120 19261 16154 19295
rect 17785 19261 17819 19295
rect 18337 19261 18371 19295
rect 21097 19261 21131 19295
rect 22293 19261 22327 19295
rect 22477 19261 22511 19295
rect 22569 19261 22603 19295
rect 22937 19261 22971 19295
rect 23213 19261 23247 19295
rect 24041 19261 24075 19295
rect 24317 19261 24351 19295
rect 24685 19261 24719 19295
rect 25145 19261 25179 19295
rect 25329 19261 25363 19295
rect 26801 19261 26835 19295
rect 4997 19193 5031 19227
rect 5089 19193 5123 19227
rect 5917 19193 5951 19227
rect 9045 19193 9079 19227
rect 9873 19193 9907 19227
rect 12081 19193 12115 19227
rect 12173 19193 12207 19227
rect 15025 19193 15059 19227
rect 17693 19193 17727 19227
rect 18797 19193 18831 19227
rect 23305 19193 23339 19227
rect 23521 19193 23555 19227
rect 23857 19193 23891 19227
rect 26534 19193 26568 19227
rect 2237 19125 2271 19159
rect 2697 19125 2731 19159
rect 3709 19125 3743 19159
rect 4445 19125 4479 19159
rect 5181 19125 5215 19159
rect 8401 19125 8435 19159
rect 9245 19125 9279 19159
rect 9413 19125 9447 19159
rect 10149 19125 10183 19159
rect 10241 19125 10275 19159
rect 12449 19125 12483 19159
rect 13645 19125 13679 19159
rect 14289 19125 14323 19159
rect 17233 19125 17267 19159
rect 18153 19125 18187 19159
rect 20637 19125 20671 19159
rect 21005 19125 21039 19159
rect 22845 19125 22879 19159
rect 23121 19125 23155 19159
rect 24225 19125 24259 19159
rect 25421 19125 25455 19159
rect 1501 18921 1535 18955
rect 1961 18921 1995 18955
rect 5457 18921 5491 18955
rect 7573 18921 7607 18955
rect 8125 18921 8159 18955
rect 8769 18921 8803 18955
rect 10333 18921 10367 18955
rect 11069 18921 11103 18955
rect 14657 18921 14691 18955
rect 16129 18921 16163 18955
rect 16589 18921 16623 18955
rect 20729 18921 20763 18955
rect 22569 18921 22603 18955
rect 24317 18921 24351 18955
rect 24593 18921 24627 18955
rect 24685 18921 24719 18955
rect 25605 18921 25639 18955
rect 25881 18921 25915 18955
rect 2688 18853 2722 18887
rect 8677 18853 8711 18887
rect 9996 18853 10030 18887
rect 14565 18853 14599 18887
rect 23204 18853 23238 18887
rect 25421 18853 25455 18887
rect 1041 18785 1075 18819
rect 2145 18785 2179 18819
rect 2421 18785 2455 18819
rect 3985 18785 4019 18819
rect 4252 18785 4286 18819
rect 5457 18785 5491 18819
rect 5641 18785 5675 18819
rect 6193 18785 6227 18819
rect 6460 18785 6494 18819
rect 8033 18785 8067 18819
rect 8217 18785 8251 18819
rect 8493 18785 8527 18819
rect 8769 18785 8803 18819
rect 10241 18785 10275 18819
rect 10517 18785 10551 18819
rect 12193 18785 12227 18819
rect 12449 18785 12483 18819
rect 12541 18785 12575 18819
rect 13737 18785 13771 18819
rect 13921 18785 13955 18819
rect 16497 18785 16531 18819
rect 17049 18785 17083 18819
rect 17325 18785 17359 18819
rect 17581 18785 17615 18819
rect 18981 18785 19015 18819
rect 19248 18785 19282 18819
rect 20637 18785 20671 18819
rect 20913 18785 20947 18819
rect 21925 18785 21959 18819
rect 22109 18785 22143 18819
rect 22201 18785 22235 18819
rect 22293 18785 22327 18819
rect 22937 18785 22971 18819
rect 24777 18785 24811 18819
rect 25697 18785 25731 18819
rect 2329 18717 2363 18751
rect 14749 18717 14783 18751
rect 16681 18717 16715 18751
rect 21097 18717 21131 18751
rect 24409 18717 24443 18751
rect 1409 18649 1443 18683
rect 8401 18649 8435 18683
rect 14197 18649 14231 18683
rect 17233 18649 17267 18683
rect 20361 18649 20395 18683
rect 24961 18649 24995 18683
rect 25053 18649 25087 18683
rect 3801 18581 3835 18615
rect 5365 18581 5399 18615
rect 7849 18581 7883 18615
rect 8861 18581 8895 18615
rect 12633 18581 12667 18615
rect 14105 18581 14139 18615
rect 18705 18581 18739 18615
rect 20453 18581 20487 18615
rect 25421 18581 25455 18615
rect 2789 18377 2823 18411
rect 6561 18377 6595 18411
rect 7297 18377 7331 18411
rect 10425 18377 10459 18411
rect 12449 18377 12483 18411
rect 15117 18377 15151 18411
rect 15853 18377 15887 18411
rect 17785 18377 17819 18411
rect 19809 18377 19843 18411
rect 21741 18377 21775 18411
rect 22569 18377 22603 18411
rect 23305 18377 23339 18411
rect 23673 18377 23707 18411
rect 24225 18377 24259 18411
rect 5181 18309 5215 18343
rect 7665 18309 7699 18343
rect 22661 18309 22695 18343
rect 23121 18309 23155 18343
rect 2686 18241 2720 18275
rect 2881 18241 2915 18275
rect 3985 18241 4019 18275
rect 6101 18241 6135 18275
rect 8769 18241 8803 18275
rect 11069 18241 11103 18275
rect 17509 18241 17543 18275
rect 18429 18241 18463 18275
rect 19257 18241 19291 18275
rect 20361 18241 20395 18275
rect 23397 18241 23431 18275
rect 1409 18173 1443 18207
rect 1869 18173 1903 18207
rect 2973 18173 3007 18207
rect 3433 18173 3467 18207
rect 4905 18173 4939 18207
rect 5825 18173 5859 18207
rect 6469 18173 6503 18207
rect 6653 18173 6687 18207
rect 8953 18173 8987 18207
rect 9045 18173 9079 18207
rect 9413 18173 9447 18207
rect 10057 18173 10091 18207
rect 11161 18173 11195 18207
rect 13737 18173 13771 18207
rect 15577 18173 15611 18207
rect 15669 18173 15703 18207
rect 16773 18173 16807 18207
rect 17233 18173 17267 18207
rect 18245 18173 18279 18207
rect 20617 18173 20651 18207
rect 22017 18173 22051 18207
rect 22293 18173 22327 18207
rect 22385 18173 22419 18207
rect 22845 18173 22879 18207
rect 22937 18173 22971 18207
rect 23213 18173 23247 18207
rect 23305 18173 23339 18207
rect 23949 18173 23983 18207
rect 24041 18173 24075 18207
rect 24133 18173 24167 18207
rect 24317 18173 24351 18207
rect 24593 18173 24627 18207
rect 25697 18173 25731 18207
rect 7297 18105 7331 18139
rect 14004 18105 14038 18139
rect 15209 18105 15243 18139
rect 15393 18105 15427 18139
rect 19349 18105 19383 18139
rect 19441 18105 19475 18139
rect 22201 18105 22235 18139
rect 24501 18105 24535 18139
rect 25964 18105 25998 18139
rect 1685 18037 1719 18071
rect 1777 18037 1811 18071
rect 7113 18037 7147 18071
rect 9505 18037 9539 18071
rect 18153 18037 18187 18071
rect 27077 18037 27111 18071
rect 2329 17833 2363 17867
rect 5457 17833 5491 17867
rect 7757 17833 7791 17867
rect 8493 17833 8527 17867
rect 8861 17833 8895 17867
rect 11897 17833 11931 17867
rect 15761 17833 15795 17867
rect 17601 17833 17635 17867
rect 18337 17833 18371 17867
rect 23121 17833 23155 17867
rect 25437 17833 25471 17867
rect 25605 17833 25639 17867
rect 25881 17833 25915 17867
rect 3893 17765 3927 17799
rect 11805 17765 11839 17799
rect 13645 17765 13679 17799
rect 16773 17765 16807 17799
rect 24225 17765 24259 17799
rect 24425 17765 24459 17799
rect 24777 17765 24811 17799
rect 24961 17765 24995 17799
rect 25237 17765 25271 17799
rect 857 17697 891 17731
rect 1124 17697 1158 17731
rect 2973 17697 3007 17731
rect 3617 17697 3651 17731
rect 4169 17697 4203 17731
rect 4629 17697 4663 17731
rect 4997 17697 5031 17731
rect 5181 17697 5215 17731
rect 5365 17697 5399 17731
rect 5641 17697 5675 17731
rect 6377 17697 6411 17731
rect 6644 17697 6678 17731
rect 8309 17697 8343 17731
rect 8401 17697 8435 17731
rect 8677 17697 8711 17731
rect 8953 17697 8987 17731
rect 9137 17697 9171 17731
rect 9229 17697 9263 17731
rect 9505 17697 9539 17731
rect 9689 17697 9723 17731
rect 9873 17697 9907 17731
rect 9965 17697 9999 17731
rect 10241 17697 10275 17731
rect 13010 17697 13044 17731
rect 13277 17697 13311 17731
rect 13369 17697 13403 17731
rect 13553 17697 13587 17731
rect 13737 17697 13771 17731
rect 14197 17697 14231 17731
rect 14381 17697 14415 17731
rect 14473 17697 14507 17731
rect 14657 17697 14691 17731
rect 15301 17697 15335 17731
rect 15393 17697 15427 17731
rect 16405 17697 16439 17731
rect 16865 17697 16899 17731
rect 17141 17697 17175 17731
rect 17785 17697 17819 17731
rect 18521 17697 18555 17731
rect 18705 17697 18739 17731
rect 19073 17697 19107 17731
rect 19809 17697 19843 17731
rect 21465 17697 21499 17731
rect 22385 17697 22419 17731
rect 22477 17697 22511 17731
rect 22753 17697 22787 17731
rect 23213 17697 23247 17731
rect 23949 17697 23983 17731
rect 24133 17697 24167 17731
rect 25145 17697 25179 17731
rect 25697 17697 25731 17731
rect 3341 17629 3375 17663
rect 3433 17629 3467 17663
rect 3525 17629 3559 17663
rect 3985 17629 4019 17663
rect 10057 17629 10091 17663
rect 11161 17629 11195 17663
rect 14013 17629 14047 17663
rect 19993 17629 20027 17663
rect 21281 17629 21315 17663
rect 2237 17561 2271 17595
rect 3801 17561 3835 17595
rect 4353 17561 4387 17595
rect 14565 17561 14599 17595
rect 3893 17493 3927 17527
rect 4445 17493 4479 17527
rect 8217 17493 8251 17527
rect 9413 17493 9447 17527
rect 10425 17493 10459 17527
rect 13921 17493 13955 17527
rect 14841 17493 14875 17527
rect 15209 17493 15243 17527
rect 15761 17493 15795 17527
rect 15945 17493 15979 17527
rect 17233 17493 17267 17527
rect 19257 17493 19291 17527
rect 19625 17493 19659 17527
rect 21649 17493 21683 17527
rect 22201 17493 22235 17527
rect 22661 17493 22695 17527
rect 24041 17493 24075 17527
rect 24409 17493 24443 17527
rect 24593 17493 24627 17527
rect 25421 17493 25455 17527
rect 1409 17289 1443 17323
rect 2789 17289 2823 17323
rect 4353 17289 4387 17323
rect 4537 17289 4571 17323
rect 6009 17289 6043 17323
rect 6193 17289 6227 17323
rect 6837 17289 6871 17323
rect 14013 17289 14047 17323
rect 17325 17289 17359 17323
rect 17509 17289 17543 17323
rect 20269 17289 20303 17323
rect 21833 17289 21867 17323
rect 25145 17289 25179 17323
rect 2605 17221 2639 17255
rect 3985 17221 4019 17255
rect 9781 17221 9815 17255
rect 10793 17221 10827 17255
rect 11989 17221 12023 17255
rect 23949 17221 23983 17255
rect 1869 17153 1903 17187
rect 6561 17153 6595 17187
rect 10241 17153 10275 17187
rect 10333 17153 10367 17187
rect 11253 17153 11287 17187
rect 18061 17153 18095 17187
rect 23489 17153 23523 17187
rect 25513 17153 25547 17187
rect 1593 17085 1627 17119
rect 1777 17085 1811 17119
rect 3801 17085 3835 17119
rect 4629 17085 4663 17119
rect 6101 17085 6135 17119
rect 7021 17085 7055 17119
rect 7757 17085 7791 17119
rect 8125 17085 8159 17119
rect 8217 17085 8251 17119
rect 8401 17085 8435 17119
rect 10057 17085 10091 17119
rect 10421 17085 10455 17119
rect 10609 17085 10643 17119
rect 10885 17085 10919 17119
rect 11161 17085 11195 17119
rect 13369 17085 13403 17119
rect 14197 17085 14231 17119
rect 16313 17085 16347 17119
rect 16589 17085 16623 17119
rect 16773 17085 16807 17119
rect 16865 17085 16899 17119
rect 17141 17085 17175 17119
rect 18889 17085 18923 17119
rect 20453 17085 20487 17119
rect 22523 17085 22557 17119
rect 22661 17085 22695 17119
rect 22753 17085 22787 17119
rect 22936 17085 22970 17119
rect 23029 17085 23063 17119
rect 23305 17085 23339 17119
rect 24041 17085 24075 17119
rect 24777 17085 24811 17119
rect 25237 17085 25271 17119
rect 25421 17085 25455 17119
rect 2973 17017 3007 17051
rect 4353 17017 4387 17051
rect 4896 17017 4930 17051
rect 8668 17017 8702 17051
rect 13124 17017 13158 17051
rect 13553 17017 13587 17051
rect 13737 17017 13771 17051
rect 13921 17017 13955 17051
rect 16129 17017 16163 17051
rect 17969 17017 18003 17051
rect 19156 17017 19190 17051
rect 20698 17017 20732 17051
rect 24685 17017 24719 17051
rect 24961 17017 24995 17051
rect 25780 17017 25814 17051
rect 2763 16949 2797 16983
rect 3249 16949 3283 16983
rect 8033 16949 8067 16983
rect 9873 16949 9907 16983
rect 11069 16949 11103 16983
rect 11897 16949 11931 16983
rect 14841 16949 14875 16983
rect 16313 16949 16347 16983
rect 16957 16949 16991 16983
rect 17877 16949 17911 16983
rect 22385 16949 22419 16983
rect 23121 16949 23155 16983
rect 24133 16949 24167 16983
rect 24317 16949 24351 16983
rect 24409 16949 24443 16983
rect 24501 16949 24535 16983
rect 25237 16949 25271 16983
rect 26893 16949 26927 16983
rect 2421 16745 2455 16779
rect 3249 16745 3283 16779
rect 7021 16745 7055 16779
rect 9045 16745 9079 16779
rect 10517 16745 10551 16779
rect 10977 16745 11011 16779
rect 13277 16745 13311 16779
rect 15209 16745 15243 16779
rect 16313 16745 16347 16779
rect 16589 16745 16623 16779
rect 18521 16745 18555 16779
rect 19073 16745 19107 16779
rect 19441 16745 19475 16779
rect 20545 16745 20579 16779
rect 21281 16745 21315 16779
rect 21649 16745 21683 16779
rect 21741 16745 21775 16779
rect 24225 16745 24259 16779
rect 24685 16745 24719 16779
rect 24869 16745 24903 16779
rect 25053 16745 25087 16779
rect 25513 16745 25547 16779
rect 25789 16745 25823 16779
rect 7941 16677 7975 16711
rect 9137 16677 9171 16711
rect 10149 16677 10183 16711
rect 19533 16677 19567 16711
rect 22937 16677 22971 16711
rect 9367 16643 9401 16677
rect 1041 16609 1075 16643
rect 1308 16609 1342 16643
rect 2697 16609 2731 16643
rect 2973 16609 3007 16643
rect 4373 16609 4407 16643
rect 6837 16609 6871 16643
rect 7021 16609 7055 16643
rect 7665 16609 7699 16643
rect 7849 16609 7883 16643
rect 8125 16609 8159 16643
rect 8309 16609 8343 16643
rect 8493 16609 8527 16643
rect 9965 16609 9999 16643
rect 10241 16609 10275 16643
rect 10333 16609 10367 16643
rect 12090 16609 12124 16643
rect 12357 16609 12391 16643
rect 13093 16609 13127 16643
rect 13829 16609 13863 16643
rect 14096 16609 14130 16643
rect 15485 16609 15519 16643
rect 15669 16609 15703 16643
rect 16129 16609 16163 16643
rect 16773 16609 16807 16643
rect 17049 16609 17083 16643
rect 17316 16609 17350 16643
rect 18705 16609 18739 16643
rect 20729 16609 20763 16643
rect 22477 16609 22511 16643
rect 22569 16609 22603 16643
rect 23029 16609 23063 16643
rect 23121 16609 23155 16643
rect 24041 16609 24075 16643
rect 24225 16609 24259 16643
rect 25145 16609 25179 16643
rect 25329 16609 25363 16643
rect 25605 16609 25639 16643
rect 2513 16541 2547 16575
rect 4629 16541 4663 16575
rect 7481 16541 7515 16575
rect 18889 16541 18923 16575
rect 19717 16541 19751 16575
rect 21833 16541 21867 16575
rect 24317 16541 24351 16575
rect 2881 16473 2915 16507
rect 18429 16473 18463 16507
rect 6653 16405 6687 16439
rect 7757 16405 7791 16439
rect 9321 16405 9355 16439
rect 9505 16405 9539 16439
rect 15301 16405 15335 16439
rect 22293 16405 22327 16439
rect 22845 16405 22879 16439
rect 23121 16405 23155 16439
rect 23397 16405 23431 16439
rect 24685 16405 24719 16439
rect 2697 16201 2731 16235
rect 5917 16201 5951 16235
rect 8861 16201 8895 16235
rect 11069 16201 11103 16235
rect 12173 16201 12207 16235
rect 14289 16201 14323 16235
rect 19993 16201 20027 16235
rect 25421 16201 25455 16235
rect 7389 16133 7423 16167
rect 20729 16133 20763 16167
rect 8033 16065 8067 16099
rect 15117 16065 15151 16099
rect 15209 16065 15243 16099
rect 15761 16065 15795 16099
rect 2053 15997 2087 16031
rect 2145 15997 2179 16031
rect 2237 15997 2271 16031
rect 2421 15997 2455 16031
rect 2513 15997 2547 16031
rect 2881 15997 2915 16031
rect 2973 15997 3007 16031
rect 3433 15997 3467 16031
rect 4537 15997 4571 16031
rect 6009 15997 6043 16031
rect 10149 15997 10183 16031
rect 10977 15997 11011 16031
rect 11253 15997 11287 16031
rect 11345 15997 11379 16031
rect 11621 15997 11655 16031
rect 14473 15997 14507 16031
rect 15025 15997 15059 16031
rect 15853 15997 15887 16031
rect 16129 15997 16163 16031
rect 16681 15997 16715 16031
rect 17509 15997 17543 16031
rect 18337 15997 18371 16031
rect 18429 15997 18463 16031
rect 20545 15997 20579 16031
rect 20913 15997 20947 16031
rect 21097 15997 21131 16031
rect 24133 15997 24167 16031
rect 26534 15997 26568 16031
rect 26801 15997 26835 16031
rect 3617 15929 3651 15963
rect 4804 15929 4838 15963
rect 6276 15929 6310 15963
rect 10701 15929 10735 15963
rect 11437 15929 11471 15963
rect 12081 15929 12115 15963
rect 18705 15929 18739 15963
rect 1777 15861 1811 15895
rect 3249 15861 3283 15895
rect 7481 15861 7515 15895
rect 14657 15861 14691 15895
rect 15485 15861 15519 15895
rect 17693 15861 17727 15895
rect 18153 15861 18187 15895
rect 20913 15861 20947 15895
rect 24225 15861 24259 15895
rect 2513 15657 2547 15691
rect 6745 15657 6779 15691
rect 9045 15657 9079 15691
rect 10517 15657 10551 15691
rect 15301 15657 15335 15691
rect 16129 15657 16163 15691
rect 18981 15657 19015 15691
rect 21005 15657 21039 15691
rect 22845 15657 22879 15691
rect 23213 15657 23247 15691
rect 7849 15589 7883 15623
rect 8049 15589 8083 15623
rect 10180 15589 10214 15623
rect 15853 15589 15887 15623
rect 17242 15589 17276 15623
rect 17846 15589 17880 15623
rect 22201 15589 22235 15623
rect 24041 15589 24075 15623
rect 24409 15589 24443 15623
rect 24593 15589 24627 15623
rect 1225 15521 1259 15555
rect 1317 15521 1351 15555
rect 1409 15521 1443 15555
rect 1593 15521 1627 15555
rect 1777 15521 1811 15555
rect 3516 15521 3550 15555
rect 5641 15521 5675 15555
rect 5917 15521 5951 15555
rect 6469 15521 6503 15555
rect 6561 15521 6595 15555
rect 6837 15521 6871 15555
rect 7297 15521 7331 15555
rect 10425 15521 10459 15555
rect 10701 15521 10735 15555
rect 11244 15521 11278 15555
rect 12449 15521 12483 15555
rect 12716 15521 12750 15555
rect 14289 15521 14323 15555
rect 15209 15521 15243 15555
rect 15761 15521 15795 15555
rect 15945 15521 15979 15555
rect 19349 15521 19383 15555
rect 19901 15521 19935 15555
rect 20729 15521 20763 15555
rect 22109 15521 22143 15555
rect 22293 15521 22327 15555
rect 22848 15521 22882 15555
rect 23213 15521 23247 15555
rect 23581 15521 23615 15555
rect 23673 15521 23707 15555
rect 23857 15521 23891 15555
rect 25421 15521 25455 15555
rect 3157 15453 3191 15487
rect 3249 15453 3283 15487
rect 5273 15453 5307 15487
rect 7481 15453 7515 15487
rect 8861 15453 8895 15487
rect 10977 15453 11011 15487
rect 14381 15453 14415 15487
rect 14473 15453 14507 15487
rect 15485 15453 15519 15487
rect 17509 15453 17543 15487
rect 17601 15453 17635 15487
rect 19441 15453 19475 15487
rect 20269 15453 20303 15487
rect 21281 15453 21315 15487
rect 22385 15453 22419 15487
rect 23305 15453 23339 15487
rect 4629 15385 4663 15419
rect 6193 15385 6227 15419
rect 8309 15385 8343 15419
rect 19349 15385 19383 15419
rect 22477 15385 22511 15419
rect 23489 15385 23523 15419
rect 949 15317 983 15351
rect 2421 15317 2455 15351
rect 4721 15317 4755 15351
rect 5549 15317 5583 15351
rect 8033 15317 8067 15351
rect 8217 15317 8251 15351
rect 12357 15317 12391 15351
rect 13829 15317 13863 15351
rect 13921 15317 13955 15351
rect 14841 15317 14875 15351
rect 21925 15317 21959 15351
rect 23029 15317 23063 15351
rect 24777 15317 24811 15351
rect 25605 15317 25639 15351
rect 949 15113 983 15147
rect 3893 15113 3927 15147
rect 5365 15113 5399 15147
rect 6561 15113 6595 15147
rect 6653 15113 6687 15147
rect 8217 15113 8251 15147
rect 13369 15113 13403 15147
rect 17601 15113 17635 15147
rect 19625 15113 19659 15147
rect 21373 15113 21407 15147
rect 23305 15113 23339 15147
rect 24869 15113 24903 15147
rect 25053 15113 25087 15147
rect 10425 15045 10459 15079
rect 12265 15045 12299 15079
rect 12725 15045 12759 15079
rect 15577 15045 15611 15079
rect 23949 15045 23983 15079
rect 1685 14977 1719 15011
rect 5917 14977 5951 15011
rect 6561 14977 6595 15011
rect 6837 14977 6871 15011
rect 11069 14977 11103 15011
rect 15209 14977 15243 15011
rect 15945 14977 15979 15011
rect 18153 14977 18187 15011
rect 21741 14977 21775 15011
rect 1593 14909 1627 14943
rect 1952 14909 1986 14943
rect 3249 14909 3283 14943
rect 3433 14909 3467 14943
rect 3525 14909 3559 14943
rect 3617 14909 3651 14943
rect 4077 14909 4111 14943
rect 6745 14909 6779 14943
rect 8493 14909 8527 14943
rect 8677 14909 8711 14943
rect 8953 14909 8987 14943
rect 9045 14909 9079 14943
rect 11805 14909 11839 14943
rect 12909 14909 12943 14943
rect 13093 14909 13127 14943
rect 13185 14909 13219 14943
rect 14289 14909 14323 14943
rect 14473 14909 14507 14943
rect 14657 14909 14691 14943
rect 14933 14909 14967 14943
rect 15577 14909 15611 14943
rect 17969 14909 18003 14943
rect 20749 14909 20783 14943
rect 21005 14909 21039 14943
rect 21649 14909 21683 14943
rect 22845 14909 22879 14943
rect 23489 14909 23523 14943
rect 24041 14909 24075 14943
rect 24133 14909 24167 14943
rect 24317 14909 24351 14943
rect 24409 14909 24443 14943
rect 24593 14909 24627 14943
rect 25329 14909 25363 14943
rect 26718 14909 26752 14943
rect 26985 14909 27019 14943
rect 6101 14841 6135 14875
rect 6285 14841 6319 14875
rect 6377 14841 6411 14875
rect 7104 14841 7138 14875
rect 9312 14841 9346 14875
rect 13645 14841 13679 14875
rect 14013 14841 14047 14875
rect 19441 14841 19475 14875
rect 24685 14841 24719 14875
rect 24901 14841 24935 14875
rect 25145 14841 25179 14875
rect 3065 14773 3099 14807
rect 8861 14773 8895 14807
rect 10517 14773 10551 14807
rect 11805 14773 11839 14807
rect 18061 14773 18095 14807
rect 19165 14773 19199 14807
rect 22293 14773 22327 14807
rect 23029 14773 23063 14807
rect 24133 14773 24167 14807
rect 24593 14773 24627 14807
rect 25513 14773 25547 14807
rect 25605 14773 25639 14807
rect 8125 14569 8159 14603
rect 9413 14569 9447 14603
rect 10133 14569 10167 14603
rect 13829 14569 13863 14603
rect 15301 14569 15335 14603
rect 24501 14569 24535 14603
rect 24593 14569 24627 14603
rect 25805 14569 25839 14603
rect 25973 14569 26007 14603
rect 1124 14501 1158 14535
rect 9013 14501 9047 14535
rect 9229 14501 9263 14535
rect 10333 14501 10367 14535
rect 12265 14501 12299 14535
rect 14166 14501 14200 14535
rect 20453 14501 20487 14535
rect 21557 14501 21591 14535
rect 22845 14501 22879 14535
rect 25329 14501 25363 14535
rect 25605 14501 25639 14535
rect 857 14433 891 14467
rect 2605 14433 2639 14467
rect 2789 14433 2823 14467
rect 2881 14433 2915 14467
rect 2973 14433 3007 14467
rect 4077 14433 4111 14467
rect 6745 14433 6779 14467
rect 7012 14433 7046 14467
rect 8309 14433 8343 14467
rect 8493 14433 8527 14467
rect 8677 14433 8711 14467
rect 8769 14433 8803 14467
rect 9597 14433 9631 14467
rect 9781 14433 9815 14467
rect 9873 14433 9907 14467
rect 10425 14433 10459 14467
rect 13645 14433 13679 14467
rect 16681 14433 16715 14467
rect 17693 14433 17727 14467
rect 18429 14433 18463 14467
rect 18889 14433 18923 14467
rect 19533 14433 19567 14467
rect 19993 14433 20027 14467
rect 20637 14433 20671 14467
rect 21465 14433 21499 14467
rect 21649 14433 21683 14467
rect 21833 14433 21867 14467
rect 22017 14433 22051 14467
rect 22661 14433 22695 14467
rect 22753 14433 22787 14467
rect 23029 14433 23063 14467
rect 23119 14423 23153 14457
rect 23237 14433 23271 14467
rect 24685 14433 24719 14467
rect 26065 14433 26099 14467
rect 26617 14433 26651 14467
rect 3249 14365 3283 14399
rect 3341 14365 3375 14399
rect 4629 14365 4663 14399
rect 4997 14365 5031 14399
rect 6561 14365 6595 14399
rect 10517 14365 10551 14399
rect 10977 14365 11011 14399
rect 12081 14365 12115 14399
rect 12173 14365 12207 14399
rect 13921 14365 13955 14399
rect 16865 14365 16899 14399
rect 17601 14365 17635 14399
rect 18153 14365 18187 14399
rect 19809 14365 19843 14399
rect 3985 14297 4019 14331
rect 5641 14297 5675 14331
rect 8861 14297 8895 14331
rect 9965 14297 9999 14331
rect 24869 14297 24903 14331
rect 24961 14297 24995 14331
rect 25513 14297 25547 14331
rect 26433 14297 26467 14331
rect 2237 14229 2271 14263
rect 5917 14229 5951 14263
rect 9045 14229 9079 14263
rect 10149 14229 10183 14263
rect 11621 14229 11655 14263
rect 12633 14229 12667 14263
rect 16497 14229 16531 14263
rect 19625 14229 19659 14263
rect 19717 14229 19751 14263
rect 20085 14229 20119 14263
rect 20821 14229 20855 14263
rect 21281 14229 21315 14263
rect 22293 14229 22327 14263
rect 22477 14229 22511 14263
rect 23305 14229 23339 14263
rect 24317 14229 24351 14263
rect 25329 14229 25363 14263
rect 25789 14229 25823 14263
rect 26249 14229 26283 14263
rect 1409 14025 1443 14059
rect 3249 14025 3283 14059
rect 6653 14025 6687 14059
rect 7021 14025 7055 14059
rect 7205 14025 7239 14059
rect 12725 14025 12759 14059
rect 17141 14025 17175 14059
rect 24961 14025 24995 14059
rect 25605 14025 25639 14059
rect 7297 13957 7331 13991
rect 17509 13957 17543 13991
rect 22845 13957 22879 13991
rect 23857 13957 23891 13991
rect 25329 13957 25363 13991
rect 4629 13889 4663 13923
rect 6193 13889 6227 13923
rect 7389 13889 7423 13923
rect 13093 13889 13127 13923
rect 14657 13889 14691 13923
rect 15761 13889 15795 13923
rect 18061 13889 18095 13923
rect 23489 13889 23523 13923
rect 24409 13889 24443 13923
rect 24869 13889 24903 13923
rect 1225 13821 1259 13855
rect 1501 13821 1535 13855
rect 2881 13821 2915 13855
rect 4362 13821 4396 13855
rect 5926 13821 5960 13855
rect 6745 13821 6779 13855
rect 6837 13821 6871 13855
rect 7021 13821 7055 13855
rect 7113 13821 7147 13855
rect 9045 13821 9079 13855
rect 11253 13821 11287 13855
rect 12909 13821 12943 13855
rect 13553 13821 13587 13855
rect 13737 13821 13771 13855
rect 14565 13821 14599 13855
rect 14841 13821 14875 13855
rect 15485 13821 15519 13855
rect 16017 13821 16051 13855
rect 17417 13821 17451 13855
rect 17969 13821 18003 13855
rect 19625 13821 19659 13855
rect 21465 13821 21499 13855
rect 24041 13821 24075 13855
rect 24133 13821 24167 13855
rect 25145 13821 25179 13855
rect 25237 13821 25271 13855
rect 26718 13821 26752 13855
rect 26985 13821 27019 13855
rect 1041 13753 1075 13787
rect 6285 13753 6319 13787
rect 6469 13753 6503 13787
rect 11520 13753 11554 13787
rect 21710 13753 21744 13787
rect 24501 13753 24535 13787
rect 2145 13685 2179 13719
rect 2237 13685 2271 13719
rect 4813 13685 4847 13719
rect 10333 13685 10367 13719
rect 12633 13685 12667 13719
rect 13921 13685 13955 13719
rect 14381 13685 14415 13719
rect 15025 13685 15059 13719
rect 15669 13685 15703 13719
rect 17233 13685 17267 13719
rect 17877 13685 17911 13719
rect 20913 13685 20947 13719
rect 22937 13685 22971 13719
rect 24593 13685 24627 13719
rect 2973 13481 3007 13515
rect 5365 13481 5399 13515
rect 9413 13481 9447 13515
rect 12265 13481 12299 13515
rect 15393 13481 15427 13515
rect 16129 13481 16163 13515
rect 16497 13481 16531 13515
rect 18429 13481 18463 13515
rect 18797 13481 18831 13515
rect 20453 13481 20487 13515
rect 22661 13481 22695 13515
rect 23397 13481 23431 13515
rect 24133 13481 24167 13515
rect 24869 13481 24903 13515
rect 1992 13413 2026 13447
rect 3249 13413 3283 13447
rect 3433 13413 3467 13447
rect 3985 13413 4019 13447
rect 4997 13413 5031 13447
rect 6184 13413 6218 13447
rect 10548 13413 10582 13447
rect 11713 13413 11747 13447
rect 16589 13413 16623 13447
rect 26004 13413 26038 13447
rect 2237 13345 2271 13379
rect 2329 13345 2363 13379
rect 2513 13345 2547 13379
rect 2605 13345 2639 13379
rect 2697 13345 2731 13379
rect 3617 13345 3651 13379
rect 3709 13345 3743 13379
rect 4169 13345 4203 13379
rect 4445 13345 4479 13379
rect 5917 13345 5951 13379
rect 8309 13345 8343 13379
rect 11897 13345 11931 13379
rect 12081 13345 12115 13379
rect 12173 13345 12207 13379
rect 12449 13345 12483 13379
rect 12541 13345 12575 13379
rect 12808 13345 12842 13379
rect 14013 13345 14047 13379
rect 14280 13345 14314 13379
rect 17049 13345 17083 13379
rect 17316 13345 17350 13379
rect 19910 13345 19944 13379
rect 20177 13345 20211 13379
rect 20637 13345 20671 13379
rect 20729 13345 20763 13379
rect 20821 13345 20855 13379
rect 21005 13345 21039 13379
rect 21281 13345 21315 13379
rect 21548 13345 21582 13379
rect 23029 13345 23063 13379
rect 23213 13345 23247 13379
rect 23581 13345 23615 13379
rect 23673 13345 23707 13379
rect 23857 13345 23891 13379
rect 23949 13345 23983 13379
rect 24041 13345 24075 13379
rect 24225 13345 24259 13379
rect 24501 13345 24535 13379
rect 26249 13345 26283 13379
rect 4813 13277 4847 13311
rect 4905 13277 4939 13311
rect 7941 13277 7975 13311
rect 8401 13277 8435 13311
rect 10793 13277 10827 13311
rect 11529 13277 11563 13311
rect 16681 13277 16715 13311
rect 22937 13277 22971 13311
rect 23121 13277 23155 13311
rect 24685 13277 24719 13311
rect 3893 13209 3927 13243
rect 4261 13209 4295 13243
rect 4353 13209 4387 13243
rect 7297 13209 7331 13243
rect 857 13141 891 13175
rect 3157 13141 3191 13175
rect 3709 13141 3743 13175
rect 7389 13141 7423 13175
rect 8585 13141 8619 13175
rect 10977 13141 11011 13175
rect 13921 13141 13955 13175
rect 22753 13141 22787 13175
rect 24317 13141 24351 13175
rect 1593 12937 1627 12971
rect 6285 12937 6319 12971
rect 7941 12937 7975 12971
rect 11713 12937 11747 12971
rect 11897 12937 11931 12971
rect 12817 12937 12851 12971
rect 14565 12937 14599 12971
rect 18153 12937 18187 12971
rect 19993 12937 20027 12971
rect 23213 12937 23247 12971
rect 24501 12937 24535 12971
rect 7113 12869 7147 12903
rect 13553 12869 13587 12903
rect 20545 12869 20579 12903
rect 24133 12869 24167 12903
rect 9689 12801 9723 12835
rect 9781 12801 9815 12835
rect 12725 12801 12759 12835
rect 14105 12801 14139 12835
rect 15209 12801 15243 12835
rect 16405 12801 16439 12835
rect 18521 12801 18555 12835
rect 19257 12801 19291 12835
rect 21833 12801 21867 12835
rect 23949 12801 23983 12835
rect 26893 12801 26927 12835
rect 1225 12733 1259 12767
rect 3065 12733 3099 12767
rect 3801 12733 3835 12767
rect 4261 12733 4295 12767
rect 4353 12733 4387 12767
rect 4445 12733 4479 12767
rect 4629 12733 4663 12767
rect 5273 12733 5307 12767
rect 5641 12733 5675 12767
rect 5825 12733 5859 12767
rect 5917 12733 5951 12767
rect 6009 12733 6043 12767
rect 6469 12733 6503 12767
rect 8033 12733 8067 12767
rect 10241 12733 10275 12767
rect 12173 12733 12207 12767
rect 12541 12733 12575 12767
rect 13001 12733 13035 12767
rect 14013 12733 14047 12767
rect 14933 12733 14967 12767
rect 16221 12733 16255 12767
rect 18337 12733 18371 12767
rect 18705 12733 18739 12767
rect 20177 12733 20211 12767
rect 20453 12733 20487 12767
rect 20729 12733 20763 12767
rect 20913 12733 20947 12767
rect 21281 12733 21315 12767
rect 22477 12733 22511 12767
rect 22753 12733 22787 12767
rect 22845 12733 22879 12767
rect 23121 12733 23155 12767
rect 23857 12733 23891 12767
rect 24041 12733 24075 12767
rect 25329 12733 25363 12767
rect 11759 12699 11793 12733
rect 1409 12665 1443 12699
rect 2798 12665 2832 12699
rect 4721 12665 4755 12699
rect 7021 12665 7055 12699
rect 7297 12665 7331 12699
rect 7481 12665 7515 12699
rect 9597 12665 9631 12699
rect 11529 12665 11563 12699
rect 13921 12665 13955 12699
rect 16313 12665 16347 12699
rect 18981 12665 19015 12699
rect 21097 12665 21131 12699
rect 21189 12665 21223 12699
rect 22937 12665 22971 12699
rect 23397 12665 23431 12699
rect 23581 12665 23615 12699
rect 26626 12665 26660 12699
rect 1685 12597 1719 12631
rect 3249 12597 3283 12631
rect 3985 12597 4019 12631
rect 7573 12597 7607 12631
rect 9229 12597 9263 12631
rect 10149 12597 10183 12631
rect 11989 12597 12023 12631
rect 12357 12597 12391 12631
rect 15025 12597 15059 12631
rect 15853 12597 15887 12631
rect 19901 12597 19935 12631
rect 20361 12597 20395 12631
rect 21465 12597 21499 12631
rect 22569 12597 22603 12631
rect 24501 12597 24535 12631
rect 24685 12597 24719 12631
rect 24777 12597 24811 12631
rect 25513 12597 25547 12631
rect 1409 12393 1443 12427
rect 2881 12393 2915 12427
rect 3433 12393 3467 12427
rect 7757 12393 7791 12427
rect 10149 12393 10183 12427
rect 15485 12393 15519 12427
rect 15945 12393 15979 12427
rect 19625 12393 19659 12427
rect 20729 12393 20763 12427
rect 22661 12393 22695 12427
rect 23397 12393 23431 12427
rect 23857 12393 23891 12427
rect 26249 12393 26283 12427
rect 26617 12393 26651 12427
rect 3792 12325 3826 12359
rect 5641 12325 5675 12359
rect 7306 12325 7340 12359
rect 8769 12325 8803 12359
rect 11336 12325 11370 12359
rect 12725 12325 12759 12359
rect 14473 12325 14507 12359
rect 17242 12325 17276 12359
rect 20269 12325 20303 12359
rect 21526 12325 21560 12359
rect 1041 12257 1075 12291
rect 1225 12257 1259 12291
rect 1501 12257 1535 12291
rect 1685 12257 1719 12291
rect 1777 12257 1811 12291
rect 1869 12257 1903 12291
rect 2973 12257 3007 12291
rect 3157 12257 3191 12291
rect 3249 12257 3283 12291
rect 4997 12257 5031 12291
rect 5181 12257 5215 12291
rect 5273 12257 5307 12291
rect 5365 12257 5399 12291
rect 7665 12257 7699 12291
rect 8309 12257 8343 12291
rect 8493 12257 8527 12291
rect 8861 12257 8895 12291
rect 9045 12257 9079 12291
rect 9321 12257 9355 12291
rect 10793 12257 10827 12291
rect 11069 12257 11103 12291
rect 14565 12257 14599 12291
rect 14749 12257 14783 12291
rect 15301 12257 15335 12291
rect 15761 12257 15795 12291
rect 17960 12257 17994 12291
rect 19533 12257 19567 12291
rect 20361 12257 20395 12291
rect 21281 12257 21315 12291
rect 23949 12257 23983 12291
rect 24869 12257 24903 12291
rect 25125 12257 25159 12291
rect 26433 12257 26467 12291
rect 2145 12189 2179 12223
rect 2237 12189 2271 12223
rect 3525 12189 3559 12223
rect 7573 12189 7607 12223
rect 9873 12189 9907 12223
rect 10057 12189 10091 12223
rect 15577 12189 15611 12223
rect 17509 12189 17543 12223
rect 17693 12189 17727 12223
rect 19717 12189 19751 12223
rect 20085 12189 20119 12223
rect 22845 12189 22879 12223
rect 23489 12189 23523 12223
rect 23673 12189 23707 12223
rect 24593 12189 24627 12223
rect 10517 12121 10551 12155
rect 16129 12121 16163 12155
rect 2973 12053 3007 12087
rect 4905 12053 4939 12087
rect 6193 12053 6227 12087
rect 9137 12053 9171 12087
rect 9597 12053 9631 12087
rect 10609 12053 10643 12087
rect 12449 12053 12483 12087
rect 14565 12053 14599 12087
rect 19073 12053 19107 12087
rect 19165 12053 19199 12087
rect 24041 12053 24075 12087
rect 9137 11849 9171 11883
rect 12449 11849 12483 11883
rect 17969 11849 18003 11883
rect 19073 11849 19107 11883
rect 23121 11849 23155 11883
rect 23305 11849 23339 11883
rect 23949 11849 23983 11883
rect 24777 11849 24811 11883
rect 24869 11849 24903 11883
rect 26801 11849 26835 11883
rect 4353 11781 4387 11815
rect 8217 11781 8251 11815
rect 15209 11781 15243 11815
rect 22477 11781 22511 11815
rect 2881 11713 2915 11747
rect 5365 11713 5399 11747
rect 9689 11713 9723 11747
rect 11897 11713 11931 11747
rect 11989 11713 12023 11747
rect 13185 11713 13219 11747
rect 15761 11713 15795 11747
rect 17601 11713 17635 11747
rect 20637 11713 20671 11747
rect 21097 11713 21131 11747
rect 1225 11645 1259 11679
rect 1409 11645 1443 11679
rect 1777 11645 1811 11679
rect 1869 11645 1903 11679
rect 1961 11645 1995 11679
rect 2145 11645 2179 11679
rect 4169 11645 4203 11679
rect 4537 11645 4571 11679
rect 4629 11645 4663 11679
rect 6837 11645 6871 11679
rect 8677 11645 8711 11679
rect 8769 11645 8803 11679
rect 8861 11645 8895 11679
rect 9045 11645 9079 11679
rect 9965 11645 9999 11679
rect 11437 11645 11471 11679
rect 12081 11645 12115 11679
rect 12909 11645 12943 11679
rect 13737 11645 13771 11679
rect 15669 11645 15703 11679
rect 17509 11645 17543 11679
rect 18153 11645 18187 11679
rect 18705 11645 18739 11679
rect 18889 11645 18923 11679
rect 20370 11645 20404 11679
rect 21364 11645 21398 11679
rect 22845 11645 22879 11679
rect 22937 11645 22971 11679
rect 23213 11645 23247 11679
rect 23489 11645 23523 11679
rect 23581 11645 23615 11679
rect 23857 11645 23891 11679
rect 24041 11645 24075 11679
rect 24133 11645 24167 11679
rect 24317 11645 24351 11679
rect 24409 11645 24443 11679
rect 24501 11645 24535 11679
rect 25237 11645 25271 11679
rect 1041 11577 1075 11611
rect 5273 11577 5307 11611
rect 5610 11577 5644 11611
rect 7104 11577 7138 11611
rect 10232 11577 10266 11611
rect 14004 11577 14038 11611
rect 15577 11577 15611 11611
rect 25053 11577 25087 11611
rect 25329 11577 25363 11611
rect 1501 11509 1535 11543
rect 2237 11509 2271 11543
rect 3525 11509 3559 11543
rect 6745 11509 6779 11543
rect 8401 11509 8435 11543
rect 11345 11509 11379 11543
rect 11621 11509 11655 11543
rect 12541 11509 12575 11543
rect 13001 11509 13035 11543
rect 15117 11509 15151 11543
rect 17049 11509 17083 11543
rect 17417 11509 17451 11543
rect 19257 11509 19291 11543
rect 22661 11509 22695 11543
rect 2237 11305 2271 11339
rect 4629 11305 4663 11339
rect 7113 11305 7147 11339
rect 7757 11305 7791 11339
rect 8953 11305 8987 11339
rect 9873 11305 9907 11339
rect 13461 11305 13495 11339
rect 14105 11305 14139 11339
rect 15025 11305 15059 11339
rect 16681 11305 16715 11339
rect 18245 11305 18279 11339
rect 19809 11305 19843 11339
rect 25973 11305 26007 11339
rect 4353 11237 4387 11271
rect 5917 11237 5951 11271
rect 7389 11237 7423 11271
rect 7573 11237 7607 11271
rect 9137 11237 9171 11271
rect 10241 11237 10275 11271
rect 12142 11237 12176 11271
rect 17018 11237 17052 11271
rect 22937 11237 22971 11271
rect 23918 11237 23952 11271
rect 1124 11169 1158 11203
rect 2605 11169 2639 11203
rect 2964 11169 2998 11203
rect 4169 11169 4203 11203
rect 4905 11169 4939 11203
rect 4997 11169 5031 11203
rect 5089 11169 5123 11203
rect 5273 11169 5307 11203
rect 6561 11169 6595 11203
rect 6653 11169 6687 11203
rect 6837 11169 6871 11203
rect 6929 11169 6963 11203
rect 8401 11169 8435 11203
rect 8493 11169 8527 11203
rect 9045 11169 9079 11203
rect 9505 11169 9539 11203
rect 9965 11169 9999 11203
rect 10057 11169 10091 11203
rect 11161 11169 11195 11203
rect 11904 11169 11938 11203
rect 13645 11169 13679 11203
rect 13829 11169 13863 11203
rect 14289 11169 14323 11203
rect 14381 11169 14415 11203
rect 14565 11169 14599 11203
rect 14841 11169 14875 11203
rect 16497 11169 16531 11203
rect 18429 11169 18463 11203
rect 19625 11169 19659 11203
rect 22661 11169 22695 11203
rect 22753 11169 22787 11203
rect 23581 11169 23615 11203
rect 25789 11169 25823 11203
rect 25881 11169 25915 11203
rect 857 11101 891 11135
rect 2697 11101 2731 11135
rect 4537 11101 4571 11135
rect 7205 11101 7239 11135
rect 9597 11101 9631 11135
rect 11345 11101 11379 11135
rect 14657 11101 14691 11135
rect 16773 11101 16807 11135
rect 18613 11101 18647 11135
rect 19441 11101 19475 11135
rect 23489 11101 23523 11135
rect 23673 11101 23707 11135
rect 25145 11101 25179 11135
rect 2421 11033 2455 11067
rect 4077 11033 4111 11067
rect 18153 11033 18187 11067
rect 22937 11033 22971 11067
rect 25053 11033 25087 11067
rect 6653 10965 6687 10999
rect 8585 10965 8619 10999
rect 10241 10965 10275 10999
rect 13277 10965 13311 10999
rect 14565 10965 14599 10999
rect 1501 10761 1535 10795
rect 7941 10761 7975 10795
rect 9597 10761 9631 10795
rect 24961 10761 24995 10795
rect 1409 10693 1443 10727
rect 6285 10693 6319 10727
rect 2053 10625 2087 10659
rect 4261 10625 4295 10659
rect 4905 10625 4939 10659
rect 5733 10625 5767 10659
rect 9229 10625 9263 10659
rect 10333 10625 10367 10659
rect 19533 10625 19567 10659
rect 21097 10625 21131 10659
rect 21649 10625 21683 10659
rect 22293 10625 22327 10659
rect 1041 10557 1075 10591
rect 1225 10557 1259 10591
rect 3065 10557 3099 10591
rect 3433 10557 3467 10591
rect 3617 10557 3651 10591
rect 3709 10557 3743 10591
rect 3801 10557 3835 10591
rect 5181 10557 5215 10591
rect 5273 10557 5307 10591
rect 5365 10557 5399 10591
rect 5549 10557 5583 10591
rect 6653 10557 6687 10591
rect 6745 10557 6779 10591
rect 6837 10557 6871 10591
rect 7021 10557 7055 10591
rect 7481 10557 7515 10591
rect 7573 10557 7607 10591
rect 7757 10557 7791 10591
rect 8217 10557 8251 10591
rect 9413 10557 9447 10591
rect 9505 10557 9539 10591
rect 10149 10557 10183 10591
rect 12173 10557 12207 10591
rect 12265 10557 12299 10591
rect 12449 10557 12483 10591
rect 12541 10557 12575 10591
rect 13185 10557 13219 10591
rect 13369 10557 13403 10591
rect 14933 10557 14967 10591
rect 15393 10557 15427 10591
rect 15577 10557 15611 10591
rect 16037 10557 16071 10591
rect 18705 10557 18739 10591
rect 18889 10557 18923 10591
rect 18981 10557 19015 10591
rect 19165 10557 19199 10591
rect 19717 10557 19751 10591
rect 20637 10557 20671 10591
rect 20729 10557 20763 10591
rect 20821 10557 20855 10591
rect 21005 10557 21039 10591
rect 21833 10557 21867 10591
rect 22109 10557 22143 10591
rect 24869 10557 24903 10591
rect 25053 10557 25087 10591
rect 7113 10489 7147 10523
rect 7297 10489 7331 10523
rect 9229 10489 9263 10523
rect 20361 10489 20395 10523
rect 2421 10421 2455 10455
rect 4077 10421 4111 10455
rect 4813 10421 4847 10455
rect 6377 10421 6411 10455
rect 8033 10421 8067 10455
rect 10977 10421 11011 10455
rect 11989 10421 12023 10455
rect 13277 10421 13311 10455
rect 14749 10421 14783 10455
rect 15209 10421 15243 10455
rect 16221 10421 16255 10455
rect 18797 10421 18831 10455
rect 19073 10421 19107 10455
rect 19901 10421 19935 10455
rect 21925 10421 21959 10455
rect 1869 10217 1903 10251
rect 4905 10217 4939 10251
rect 6285 10217 6319 10251
rect 9413 10217 9447 10251
rect 13461 10217 13495 10251
rect 13829 10217 13863 10251
rect 16129 10217 16163 10251
rect 17877 10217 17911 10251
rect 19349 10217 19383 10251
rect 19717 10217 19751 10251
rect 21281 10217 21315 10251
rect 3617 10149 3651 10183
rect 5825 10149 5859 10183
rect 9137 10149 9171 10183
rect 10548 10149 10582 10183
rect 14729 10149 14763 10183
rect 16497 10149 16531 10183
rect 1225 10081 1259 10115
rect 1409 10081 1443 10115
rect 1501 10081 1535 10115
rect 1593 10081 1627 10115
rect 2412 10081 2446 10115
rect 6101 10081 6135 10115
rect 7021 10081 7055 10115
rect 7205 10081 7239 10115
rect 7472 10081 7506 10115
rect 8953 10081 8987 10115
rect 10793 10081 10827 10115
rect 11069 10081 11103 10115
rect 11253 10081 11287 10115
rect 12081 10081 12115 10115
rect 12909 10081 12943 10115
rect 13001 10081 13035 10115
rect 13185 10081 13219 10115
rect 13277 10081 13311 10115
rect 13369 10081 13403 10115
rect 13553 10081 13587 10115
rect 14013 10081 14047 10115
rect 14105 10081 14139 10115
rect 14289 10081 14323 10115
rect 14381 10081 14415 10115
rect 17785 10081 17819 10115
rect 18521 10081 18555 10115
rect 18613 10081 18647 10115
rect 18797 10081 18831 10115
rect 18889 10081 18923 10115
rect 19257 10081 19291 10115
rect 20729 10081 20763 10115
rect 22394 10081 22428 10115
rect 22661 10081 22695 10115
rect 24685 10081 24719 10115
rect 2145 10013 2179 10047
rect 6009 10013 6043 10047
rect 14473 10013 14507 10047
rect 16589 10013 16623 10047
rect 16681 10013 16715 10047
rect 17969 10013 18003 10047
rect 19809 10013 19843 10047
rect 19993 10013 20027 10047
rect 20821 10013 20855 10047
rect 21097 10013 21131 10047
rect 8585 9945 8619 9979
rect 18337 9945 18371 9979
rect 3525 9877 3559 9911
rect 5825 9877 5859 9911
rect 6469 9877 6503 9911
rect 8769 9877 8803 9911
rect 12725 9877 12759 9911
rect 15853 9877 15887 9911
rect 17417 9877 17451 9911
rect 19073 9877 19107 9911
rect 24869 9877 24903 9911
rect 3801 9673 3835 9707
rect 5917 9673 5951 9707
rect 7389 9673 7423 9707
rect 8033 9673 8067 9707
rect 8217 9673 8251 9707
rect 10149 9673 10183 9707
rect 14933 9673 14967 9707
rect 17877 9673 17911 9707
rect 20361 9673 20395 9707
rect 3065 9605 3099 9639
rect 3709 9605 3743 9639
rect 9321 9605 9355 9639
rect 13185 9605 13219 9639
rect 20637 9605 20671 9639
rect 21741 9605 21775 9639
rect 24593 9605 24627 9639
rect 4537 9537 4571 9571
rect 6009 9537 6043 9571
rect 8861 9537 8895 9571
rect 9045 9537 9079 9571
rect 9873 9537 9907 9571
rect 11161 9537 11195 9571
rect 11897 9537 11931 9571
rect 15393 9537 15427 9571
rect 15577 9537 15611 9571
rect 18981 9537 19015 9571
rect 21281 9537 21315 9571
rect 22845 9537 22879 9571
rect 24133 9537 24167 9571
rect 25973 9537 26007 9571
rect 2237 9469 2271 9503
rect 2421 9469 2455 9503
rect 2605 9469 2639 9503
rect 2697 9469 2731 9503
rect 2789 9469 2823 9503
rect 3341 9469 3375 9503
rect 4445 9469 4479 9503
rect 4804 9469 4838 9503
rect 7665 9469 7699 9503
rect 8769 9469 8803 9503
rect 8953 9469 8987 9503
rect 9597 9469 9631 9503
rect 11069 9469 11103 9503
rect 12449 9469 12483 9503
rect 12633 9469 12667 9503
rect 13185 9469 13219 9503
rect 13369 9469 13403 9503
rect 14105 9469 14139 9503
rect 14197 9469 14231 9503
rect 14381 9469 14415 9503
rect 14473 9469 14507 9503
rect 15301 9469 15335 9503
rect 17233 9469 17267 9503
rect 17601 9469 17635 9503
rect 18061 9469 18095 9503
rect 18153 9469 18187 9503
rect 19237 9469 19271 9503
rect 20821 9469 20855 9503
rect 21097 9469 21131 9503
rect 21373 9469 21407 9503
rect 21557 9469 21591 9503
rect 22753 9469 22787 9503
rect 24041 9469 24075 9503
rect 25706 9469 25740 9503
rect 1970 9401 2004 9435
rect 3525 9401 3559 9435
rect 6276 9401 6310 9435
rect 8033 9401 8067 9435
rect 9689 9401 9723 9435
rect 10333 9401 10367 9435
rect 16966 9401 17000 9435
rect 857 9333 891 9367
rect 9229 9333 9263 9367
rect 9505 9333 9539 9367
rect 9965 9333 9999 9367
rect 10133 9333 10167 9367
rect 12541 9333 12575 9367
rect 13921 9333 13955 9367
rect 15853 9333 15887 9367
rect 17417 9333 17451 9367
rect 21005 9333 21039 9367
rect 23121 9333 23155 9367
rect 24409 9333 24443 9367
rect 1225 9129 1259 9163
rect 2789 9129 2823 9163
rect 3157 9129 3191 9163
rect 3433 9129 3467 9163
rect 5273 9129 5307 9163
rect 7849 9129 7883 9163
rect 9413 9129 9447 9163
rect 16589 9129 16623 9163
rect 18521 9129 18555 9163
rect 24777 9129 24811 9163
rect 3617 9061 3651 9095
rect 17397 9061 17431 9095
rect 19165 9061 19199 9095
rect 1777 8993 1811 9027
rect 1961 8993 1995 9027
rect 2145 8996 2179 9030
rect 2237 8993 2271 9027
rect 2329 8993 2363 9027
rect 2697 8993 2731 9027
rect 2973 8993 3007 9027
rect 3801 8993 3835 9027
rect 4160 8993 4194 9027
rect 7481 8993 7515 9027
rect 7946 8993 7980 9027
rect 8217 8993 8251 9027
rect 8493 8993 8527 9027
rect 8769 8993 8803 9027
rect 9045 8993 9079 9027
rect 11069 8993 11103 9027
rect 11437 8993 11471 9027
rect 13001 8993 13035 9027
rect 13093 8993 13127 9027
rect 13277 8993 13311 9027
rect 13369 8993 13403 9027
rect 14013 8993 14047 9027
rect 14105 8993 14139 9027
rect 14289 8993 14323 9027
rect 14381 8993 14415 9027
rect 14657 8993 14691 9027
rect 14841 8993 14875 9027
rect 14933 8993 14967 9027
rect 15117 8993 15151 9027
rect 16221 8993 16255 9027
rect 16405 8993 16439 9027
rect 18613 8993 18647 9027
rect 18705 8993 18739 9027
rect 18889 8993 18923 9027
rect 18981 8993 19015 9027
rect 19625 8993 19659 9027
rect 19717 8993 19751 9027
rect 19901 8993 19935 9027
rect 19993 8993 20027 9027
rect 20085 8993 20119 9027
rect 20269 8993 20303 9027
rect 22661 8993 22695 9027
rect 22845 8993 22879 9027
rect 22937 8993 22971 9027
rect 23397 8993 23431 9027
rect 23489 8993 23523 9027
rect 23581 8993 23615 9027
rect 23765 8993 23799 9027
rect 24593 8993 24627 9027
rect 2605 8925 2639 8959
rect 3893 8925 3927 8959
rect 7665 8925 7699 8959
rect 8953 8925 8987 8959
rect 12909 8925 12943 8959
rect 17141 8925 17175 8959
rect 20177 8925 20211 8959
rect 24409 8925 24443 8959
rect 8401 8857 8435 8891
rect 8585 8857 8619 8891
rect 22753 8857 22787 8891
rect 8033 8789 8067 8823
rect 9413 8789 9447 8823
rect 9597 8789 9631 8823
rect 13553 8789 13587 8823
rect 13829 8789 13863 8823
rect 14841 8789 14875 8823
rect 15117 8789 15151 8823
rect 19441 8789 19475 8823
rect 22477 8789 22511 8823
rect 23121 8789 23155 8823
rect 1409 8585 1443 8619
rect 2605 8585 2639 8619
rect 8125 8585 8159 8619
rect 10609 8585 10643 8619
rect 21741 8585 21775 8619
rect 22109 8585 22143 8619
rect 22937 8585 22971 8619
rect 23949 8585 23983 8619
rect 24041 8585 24075 8619
rect 1041 8517 1075 8551
rect 14105 8517 14139 8551
rect 16405 8517 16439 8551
rect 17601 8517 17635 8551
rect 23581 8517 23615 8551
rect 24317 8517 24351 8551
rect 25145 8517 25179 8551
rect 857 8449 891 8483
rect 1685 8449 1719 8483
rect 2053 8449 2087 8483
rect 2513 8449 2547 8483
rect 11069 8449 11103 8483
rect 12449 8449 12483 8483
rect 12633 8449 12667 8483
rect 20637 8449 20671 8483
rect 21925 8449 21959 8483
rect 24133 8449 24167 8483
rect 25421 8449 25455 8483
rect 1225 8381 1259 8415
rect 1317 8381 1351 8415
rect 1777 8381 1811 8415
rect 2237 8381 2271 8415
rect 2421 8381 2455 8415
rect 3249 8381 3283 8415
rect 5273 8381 5307 8415
rect 6745 8381 6779 8415
rect 9229 8381 9263 8415
rect 10977 8381 11011 8415
rect 12909 8381 12943 8415
rect 13277 8381 13311 8415
rect 14473 8381 14507 8415
rect 14933 8381 14967 8415
rect 15485 8381 15519 8415
rect 16221 8381 16255 8415
rect 17417 8381 17451 8415
rect 18337 8381 18371 8415
rect 18521 8381 18555 8415
rect 20453 8381 20487 8415
rect 21005 8381 21039 8415
rect 21097 8381 21131 8415
rect 21833 8381 21867 8415
rect 22201 8381 22235 8415
rect 23121 8381 23155 8415
rect 23213 8381 23247 8415
rect 23489 8381 23523 8415
rect 23673 8381 23707 8415
rect 23857 8381 23891 8415
rect 24225 8381 24259 8415
rect 24409 8381 24443 8415
rect 25605 8381 25639 8415
rect 2789 8313 2823 8347
rect 2973 8313 3007 8347
rect 3494 8313 3528 8347
rect 5540 8313 5574 8347
rect 7012 8313 7046 8347
rect 9496 8313 9530 8347
rect 12817 8313 12851 8347
rect 22937 8313 22971 8347
rect 24777 8313 24811 8347
rect 25789 8313 25823 8347
rect 4629 8245 4663 8279
rect 6653 8245 6687 8279
rect 11805 8245 11839 8279
rect 18429 8245 18463 8279
rect 19165 8245 19199 8279
rect 20913 8245 20947 8279
rect 21373 8245 21407 8279
rect 21925 8245 21959 8279
rect 25237 8245 25271 8279
rect 3249 8041 3283 8075
rect 4813 8041 4847 8075
rect 6377 8041 6411 8075
rect 9505 8041 9539 8075
rect 21925 8041 21959 8075
rect 22201 8041 22235 8075
rect 22753 8041 22787 8075
rect 23857 8041 23891 8075
rect 2513 7973 2547 8007
rect 2881 7973 2915 8007
rect 3065 7973 3099 8007
rect 3433 7973 3467 8007
rect 3617 7973 3651 8007
rect 3801 7973 3835 8007
rect 22569 7973 22603 8007
rect 22937 7973 22971 8007
rect 23489 7973 23523 8007
rect 24133 7973 24167 8007
rect 2789 7905 2823 7939
rect 3157 7905 3191 7939
rect 3985 7905 4019 7939
rect 4169 7905 4203 7939
rect 4445 7905 4479 7939
rect 4905 7905 4939 7939
rect 5089 7905 5123 7939
rect 5365 7905 5399 7939
rect 6561 7905 6595 7939
rect 6653 7905 6687 7939
rect 6837 7905 6871 7939
rect 9689 7905 9723 7939
rect 11897 7905 11931 7939
rect 11989 7905 12023 7939
rect 12265 7905 12299 7939
rect 12357 7905 12391 7939
rect 12541 7905 12575 7939
rect 12633 7905 12667 7939
rect 14197 7905 14231 7939
rect 14289 7905 14323 7939
rect 14473 7905 14507 7939
rect 14565 7905 14599 7939
rect 14841 7905 14875 7939
rect 15485 7905 15519 7939
rect 17242 7905 17276 7939
rect 17509 7905 17543 7939
rect 18714 7905 18748 7939
rect 19073 7905 19107 7939
rect 19165 7905 19199 7939
rect 19349 7905 19383 7939
rect 19441 7905 19475 7939
rect 19984 7905 20018 7939
rect 21281 7905 21315 7939
rect 21465 7905 21499 7939
rect 21649 7905 21683 7939
rect 21741 7905 21775 7939
rect 21833 7905 21867 7939
rect 22017 7905 22051 7939
rect 22109 7905 22143 7939
rect 22293 7905 22327 7939
rect 22845 7905 22879 7939
rect 23121 7905 23155 7939
rect 23213 7905 23247 7939
rect 23673 7905 23707 7939
rect 24041 7905 24075 7939
rect 24225 7905 24259 7939
rect 24501 7905 24535 7939
rect 25993 7905 26027 7939
rect 26249 7905 26283 7939
rect 26617 7905 26651 7939
rect 2513 7837 2547 7871
rect 4353 7837 4387 7871
rect 5549 7837 5583 7871
rect 7021 7837 7055 7871
rect 11529 7837 11563 7871
rect 14933 7837 14967 7871
rect 15393 7837 15427 7871
rect 18981 7837 19015 7871
rect 19717 7837 19751 7871
rect 22937 7837 22971 7871
rect 24777 7837 24811 7871
rect 2881 7769 2915 7803
rect 16129 7769 16163 7803
rect 21097 7769 21131 7803
rect 26433 7769 26467 7803
rect 2697 7701 2731 7735
rect 4997 7701 5031 7735
rect 5181 7701 5215 7735
rect 11713 7701 11747 7735
rect 12081 7701 12115 7735
rect 14013 7701 14047 7735
rect 15117 7701 15151 7735
rect 15761 7701 15795 7735
rect 17601 7701 17635 7735
rect 19625 7701 19659 7735
rect 22569 7701 22603 7735
rect 24317 7701 24351 7735
rect 24685 7701 24719 7735
rect 24869 7701 24903 7735
rect 2421 7497 2455 7531
rect 4261 7497 4295 7531
rect 4537 7497 4571 7531
rect 6653 7497 6687 7531
rect 12909 7497 12943 7531
rect 16313 7497 16347 7531
rect 17601 7497 17635 7531
rect 23673 7497 23707 7531
rect 25329 7497 25363 7531
rect 3525 7429 3559 7463
rect 3617 7429 3651 7463
rect 1409 7361 1443 7395
rect 4353 7361 4387 7395
rect 7021 7361 7055 7395
rect 8861 7361 8895 7395
rect 19809 7361 19843 7395
rect 25145 7361 25179 7395
rect 1869 7293 1903 7327
rect 2145 7293 2179 7327
rect 2329 7293 2363 7327
rect 3249 7293 3283 7327
rect 3433 7293 3467 7327
rect 3709 7293 3743 7327
rect 4077 7293 4111 7327
rect 4169 7293 4203 7327
rect 4445 7293 4479 7327
rect 4629 7293 4663 7327
rect 5273 7293 5307 7327
rect 6929 7293 6963 7327
rect 8677 7293 8711 7327
rect 10149 7293 10183 7327
rect 10241 7293 10275 7327
rect 10333 7293 10367 7327
rect 10517 7293 10551 7327
rect 12449 7293 12483 7327
rect 12725 7293 12759 7327
rect 13001 7293 13035 7327
rect 15945 7293 15979 7327
rect 16129 7293 16163 7327
rect 17233 7293 17267 7327
rect 17417 7293 17451 7327
rect 18981 7293 19015 7327
rect 19349 7293 19383 7327
rect 19533 7293 19567 7327
rect 21649 7293 21683 7327
rect 22293 7293 22327 7327
rect 25053 7293 25087 7327
rect 25513 7293 25547 7327
rect 25697 7293 25731 7327
rect 1777 7225 1811 7259
rect 2513 7225 2547 7259
rect 9873 7225 9907 7259
rect 12204 7225 12238 7259
rect 12541 7225 12575 7259
rect 22560 7225 22594 7259
rect 1685 7157 1719 7191
rect 5457 7157 5491 7191
rect 8493 7157 8527 7191
rect 11069 7157 11103 7191
rect 19717 7157 19751 7191
rect 25513 7157 25547 7191
rect 2329 6953 2363 6987
rect 6929 6953 6963 6987
rect 7481 6953 7515 6987
rect 10425 6953 10459 6987
rect 12449 6953 12483 6987
rect 12810 6953 12844 6987
rect 14473 6953 14507 6987
rect 15117 6953 15151 6987
rect 5374 6885 5408 6919
rect 12909 6885 12943 6919
rect 857 6817 891 6851
rect 1124 6817 1158 6851
rect 2789 6817 2823 6851
rect 3157 6817 3191 6851
rect 3249 6817 3283 6851
rect 3433 6817 3467 6851
rect 3801 6817 3835 6851
rect 3893 6817 3927 6851
rect 3985 6817 4019 6851
rect 4169 6817 4203 6851
rect 5641 6817 5675 6851
rect 6193 6817 6227 6851
rect 6377 6817 6411 6851
rect 7021 6817 7055 6851
rect 7297 6817 7331 6851
rect 7665 6817 7699 6851
rect 9054 6817 9088 6851
rect 9321 6817 9355 6851
rect 9965 6817 9999 6851
rect 10057 6817 10091 6851
rect 10241 6817 10275 6851
rect 11345 6817 11379 6851
rect 11529 6817 11563 6851
rect 11897 6817 11931 6851
rect 11989 6817 12023 6851
rect 12633 6817 12667 6851
rect 12725 6817 12759 6851
rect 13001 6817 13035 6851
rect 13257 6817 13291 6851
rect 14657 6817 14691 6851
rect 14933 6817 14967 6851
rect 15393 6817 15427 6851
rect 16589 6817 16623 6851
rect 16773 6817 16807 6851
rect 18889 6817 18923 6851
rect 19073 6817 19107 6851
rect 19257 6817 19291 6851
rect 19349 6817 19383 6851
rect 20637 6817 20671 6851
rect 20729 6817 20763 6851
rect 20913 6817 20947 6851
rect 21097 6817 21131 6851
rect 21281 6817 21315 6851
rect 21373 6817 21407 6851
rect 21465 6817 21499 6851
rect 21649 6817 21683 6851
rect 21925 6817 21959 6851
rect 23949 6817 23983 6851
rect 24133 6817 24167 6851
rect 24317 6817 24351 6851
rect 24409 6817 24443 6851
rect 25513 6817 25547 6851
rect 25697 6817 25731 6851
rect 25789 6817 25823 6851
rect 25973 6817 26007 6851
rect 3525 6749 3559 6783
rect 6285 6749 6319 6783
rect 6469 6749 6503 6783
rect 7113 6749 7147 6783
rect 11437 6749 11471 6783
rect 11621 6749 11655 6783
rect 15117 6749 15151 6783
rect 17969 6749 18003 6783
rect 3433 6681 3467 6715
rect 4261 6681 4295 6715
rect 6745 6681 6779 6715
rect 7849 6681 7883 6715
rect 14749 6681 14783 6715
rect 14841 6681 14875 6715
rect 18337 6681 18371 6715
rect 22661 6681 22695 6715
rect 2237 6613 2271 6647
rect 2513 6613 2547 6647
rect 7941 6613 7975 6647
rect 11713 6613 11747 6647
rect 11805 6613 11839 6647
rect 12081 6613 12115 6647
rect 14381 6613 14415 6647
rect 15301 6613 15335 6647
rect 16681 6613 16715 6647
rect 18429 6613 18463 6647
rect 19533 6613 19567 6647
rect 19993 6613 20027 6647
rect 24593 6613 24627 6647
rect 25697 6613 25731 6647
rect 25881 6613 25915 6647
rect 1409 6409 1443 6443
rect 1777 6409 1811 6443
rect 2145 6409 2179 6443
rect 2329 6409 2363 6443
rect 6653 6409 6687 6443
rect 7205 6409 7239 6443
rect 8861 6409 8895 6443
rect 11713 6409 11747 6443
rect 12357 6409 12391 6443
rect 13645 6409 13679 6443
rect 14197 6409 14231 6443
rect 14657 6409 14691 6443
rect 16037 6409 16071 6443
rect 17049 6409 17083 6443
rect 21373 6409 21407 6443
rect 22477 6409 22511 6443
rect 23581 6409 23615 6443
rect 25605 6409 25639 6443
rect 25973 6409 26007 6443
rect 8125 6341 8159 6375
rect 17325 6341 17359 6375
rect 18521 6341 18555 6375
rect 26617 6341 26651 6375
rect 1869 6273 1903 6307
rect 3709 6273 3743 6307
rect 7573 6273 7607 6307
rect 7757 6273 7791 6307
rect 8217 6273 8251 6307
rect 8493 6273 8527 6307
rect 13553 6273 13587 6307
rect 16865 6273 16899 6307
rect 17233 6273 17267 6307
rect 18245 6273 18279 6307
rect 20361 6273 20395 6307
rect 24225 6273 24259 6307
rect 26341 6273 26375 6307
rect 26525 6273 26559 6307
rect 1593 6205 1627 6239
rect 1961 6205 1995 6239
rect 2145 6205 2179 6239
rect 2237 6205 2271 6239
rect 2421 6205 2455 6239
rect 2697 6205 2731 6239
rect 3617 6205 3651 6239
rect 4813 6205 4847 6239
rect 5825 6205 5859 6239
rect 6561 6205 6595 6239
rect 6745 6205 6779 6239
rect 7389 6205 7423 6239
rect 7665 6205 7699 6239
rect 8585 6205 8619 6239
rect 11529 6205 11563 6239
rect 11621 6205 11655 6239
rect 11897 6205 11931 6239
rect 12173 6205 12207 6239
rect 12357 6205 12391 6239
rect 13737 6205 13771 6239
rect 13829 6205 13863 6239
rect 14105 6205 14139 6239
rect 14289 6205 14323 6239
rect 14381 6205 14415 6239
rect 15025 6205 15059 6239
rect 15117 6205 15151 6239
rect 15209 6205 15243 6239
rect 15393 6205 15427 6239
rect 15485 6205 15519 6239
rect 16221 6205 16255 6239
rect 16405 6205 16439 6239
rect 16497 6205 16531 6239
rect 16773 6205 16807 6239
rect 18153 6205 18187 6239
rect 20269 6205 20303 6239
rect 20637 6205 20671 6239
rect 21465 6205 21499 6239
rect 21741 6205 21775 6239
rect 22569 6205 22603 6239
rect 22845 6205 22879 6239
rect 23857 6205 23891 6239
rect 24492 6205 24526 6239
rect 26249 6205 26283 6239
rect 14657 6137 14691 6171
rect 14749 6137 14783 6171
rect 15669 6137 15703 6171
rect 17693 6137 17727 6171
rect 20002 6137 20036 6171
rect 26985 6137 27019 6171
rect 3985 6069 4019 6103
rect 10241 6069 10275 6103
rect 12081 6069 12115 6103
rect 14473 6069 14507 6103
rect 15853 6069 15887 6103
rect 18889 6069 18923 6103
rect 3709 5865 3743 5899
rect 4537 5865 4571 5899
rect 6837 5865 6871 5899
rect 7849 5865 7883 5899
rect 8125 5865 8159 5899
rect 9137 5865 9171 5899
rect 15025 5865 15059 5899
rect 17601 5865 17635 5899
rect 18429 5865 18463 5899
rect 22845 5865 22879 5899
rect 23397 5865 23431 5899
rect 24501 5865 24535 5899
rect 25421 5865 25455 5899
rect 10272 5797 10306 5831
rect 16681 5797 16715 5831
rect 2329 5729 2363 5763
rect 2697 5729 2731 5763
rect 2973 5729 3007 5763
rect 5273 5729 5307 5763
rect 5549 5729 5583 5763
rect 5825 5729 5859 5763
rect 6101 5729 6135 5763
rect 7757 5729 7791 5763
rect 7941 5729 7975 5763
rect 8033 5729 8067 5763
rect 8217 5729 8251 5763
rect 11161 5729 11195 5763
rect 12265 5729 12299 5763
rect 12357 5729 12391 5763
rect 12541 5729 12575 5763
rect 13277 5729 13311 5763
rect 14933 5729 14967 5763
rect 15117 5729 15151 5763
rect 16589 5729 16623 5763
rect 16773 5729 16807 5763
rect 17785 5729 17819 5763
rect 17969 5729 18003 5763
rect 18061 5729 18095 5763
rect 18153 5729 18187 5763
rect 18337 5729 18371 5763
rect 18429 5729 18463 5763
rect 18613 5729 18647 5763
rect 21005 5729 21039 5763
rect 22569 5729 22603 5763
rect 23029 5729 23063 5763
rect 23213 5729 23247 5763
rect 23765 5729 23799 5763
rect 25605 5729 25639 5763
rect 2605 5661 2639 5695
rect 10517 5661 10551 5695
rect 11069 5661 11103 5695
rect 13001 5661 13035 5695
rect 18245 5661 18279 5695
rect 23489 5661 23523 5695
rect 25881 5661 25915 5695
rect 14013 5593 14047 5627
rect 24593 5593 24627 5627
rect 25789 5593 25823 5627
rect 1317 5525 1351 5559
rect 2145 5525 2179 5559
rect 2513 5525 2547 5559
rect 6929 5525 6963 5559
rect 11529 5525 11563 5559
rect 11805 5525 11839 5559
rect 12725 5525 12759 5559
rect 14197 5525 14231 5559
rect 15669 5525 15703 5559
rect 2237 5321 2271 5355
rect 2697 5321 2731 5355
rect 5089 5321 5123 5355
rect 5917 5321 5951 5355
rect 7665 5321 7699 5355
rect 10241 5321 10275 5355
rect 12725 5321 12759 5355
rect 13001 5321 13035 5355
rect 15209 5321 15243 5355
rect 16589 5321 16623 5355
rect 21005 5321 21039 5355
rect 22753 5321 22787 5355
rect 23121 5321 23155 5355
rect 25881 5321 25915 5355
rect 26433 5321 26467 5355
rect 11253 5253 11287 5287
rect 21557 5253 21591 5287
rect 6653 5185 6687 5219
rect 8769 5185 8803 5219
rect 14197 5185 14231 5219
rect 21189 5185 21223 5219
rect 21649 5185 21683 5219
rect 26525 5185 26559 5219
rect 1133 5117 1167 5151
rect 1225 5117 1259 5151
rect 1501 5117 1535 5151
rect 2697 5117 2731 5151
rect 2881 5117 2915 5151
rect 4905 5117 4939 5151
rect 5733 5117 5767 5151
rect 6377 5117 6411 5151
rect 6929 5117 6963 5151
rect 8493 5117 8527 5151
rect 8585 5117 8619 5151
rect 10057 5117 10091 5151
rect 10517 5117 10551 5151
rect 10793 5117 10827 5151
rect 11989 5117 12023 5151
rect 12265 5117 12299 5151
rect 12541 5117 12575 5151
rect 12725 5117 12759 5151
rect 14473 5117 14507 5151
rect 15301 5117 15335 5151
rect 15577 5117 15611 5151
rect 15853 5117 15887 5151
rect 19625 5117 19659 5151
rect 19809 5117 19843 5151
rect 20545 5117 20579 5151
rect 20729 5117 20763 5151
rect 20821 5117 20855 5151
rect 21005 5117 21039 5151
rect 21741 5117 21775 5151
rect 21925 5117 21959 5151
rect 22201 5117 22235 5151
rect 22753 5117 22787 5151
rect 22937 5117 22971 5151
rect 24133 5117 24167 5151
rect 24593 5117 24627 5151
rect 26433 5117 26467 5151
rect 10425 5049 10459 5083
rect 19993 5049 20027 5083
rect 20269 5049 20303 5083
rect 20453 5049 20487 5083
rect 20637 5049 20671 5083
rect 6561 4981 6595 5015
rect 8769 4981 8803 5015
rect 15485 4981 15519 5015
rect 20085 4981 20119 5015
rect 22109 4981 22143 5015
rect 22293 4981 22327 5015
rect 26801 4981 26835 5015
rect 2237 4777 2271 4811
rect 5825 4777 5859 4811
rect 8217 4777 8251 4811
rect 9153 4777 9187 4811
rect 9781 4777 9815 4811
rect 14381 4777 14415 4811
rect 15117 4777 15151 4811
rect 18153 4777 18187 4811
rect 21481 4777 21515 4811
rect 23489 4777 23523 4811
rect 23949 4777 23983 4811
rect 25053 4777 25087 4811
rect 26157 4777 26191 4811
rect 26633 4777 26667 4811
rect 26801 4777 26835 4811
rect 3157 4709 3191 4743
rect 8953 4709 8987 4743
rect 11161 4709 11195 4743
rect 11529 4709 11563 4743
rect 12081 4709 12115 4743
rect 12725 4709 12759 4743
rect 21281 4709 21315 4743
rect 23029 4709 23063 4743
rect 25421 4709 25455 4743
rect 26433 4709 26467 4743
rect 1225 4641 1259 4675
rect 1501 4641 1535 4675
rect 2973 4641 3007 4675
rect 3249 4641 3283 4675
rect 3433 4641 3467 4675
rect 3525 4641 3559 4675
rect 3709 4641 3743 4675
rect 4905 4641 4939 4675
rect 5089 4641 5123 4675
rect 5181 4641 5215 4675
rect 6193 4641 6227 4675
rect 7481 4641 7515 4675
rect 7665 4641 7699 4675
rect 7941 4641 7975 4675
rect 8125 4641 8159 4675
rect 8401 4641 8435 4675
rect 8677 4641 8711 4675
rect 8861 4641 8895 4675
rect 9413 4641 9447 4675
rect 10517 4641 10551 4675
rect 10793 4641 10827 4675
rect 11345 4641 11379 4675
rect 11713 4641 11747 4675
rect 11897 4641 11931 4675
rect 11989 4641 12023 4675
rect 12173 4641 12207 4675
rect 12265 4641 12299 4675
rect 12449 4641 12483 4675
rect 13461 4641 13495 4675
rect 13645 4641 13679 4675
rect 13737 4641 13771 4675
rect 14197 4641 14231 4675
rect 14749 4641 14783 4675
rect 14933 4641 14967 4675
rect 16589 4641 16623 4675
rect 17509 4641 17543 4675
rect 17693 4641 17727 4675
rect 17969 4641 18003 4675
rect 19358 4641 19392 4675
rect 19901 4641 19935 4675
rect 22009 4641 22043 4675
rect 22293 4641 22327 4675
rect 23305 4641 23339 4675
rect 23765 4641 23799 4675
rect 24317 4641 24351 4675
rect 25145 4641 25179 4675
rect 25513 4641 25547 4675
rect 25697 4641 25731 4675
rect 25973 4641 26007 4675
rect 27077 4641 27111 4675
rect 2789 4573 2823 4607
rect 3617 4573 3651 4607
rect 4169 4573 4203 4607
rect 4629 4573 4663 4607
rect 4721 4573 4755 4607
rect 6101 4573 6135 4607
rect 7757 4573 7791 4607
rect 13185 4573 13219 4607
rect 13277 4573 13311 4607
rect 15945 4573 15979 4607
rect 16313 4573 16347 4607
rect 19625 4573 19659 4607
rect 23121 4573 23155 4607
rect 24041 4573 24075 4607
rect 25421 4573 25455 4607
rect 3433 4505 3467 4539
rect 4445 4505 4479 4539
rect 7665 4505 7699 4539
rect 9321 4505 9355 4539
rect 12265 4505 12299 4539
rect 13093 4505 13127 4539
rect 17325 4505 17359 4539
rect 19993 4505 20027 4539
rect 21649 4505 21683 4539
rect 25237 4505 25271 4539
rect 5365 4437 5399 4471
rect 6009 4437 6043 4471
rect 7113 4437 7147 4471
rect 9137 4437 9171 4471
rect 9597 4437 9631 4471
rect 10977 4437 11011 4471
rect 13921 4437 13955 4471
rect 14749 4437 14783 4471
rect 18245 4437 18279 4471
rect 21465 4437 21499 4471
rect 22201 4437 22235 4471
rect 22477 4437 22511 4471
rect 23121 4437 23155 4471
rect 26617 4437 26651 4471
rect 26893 4437 26927 4471
rect 4445 4233 4479 4267
rect 4629 4233 4663 4267
rect 6285 4233 6319 4267
rect 6561 4233 6595 4267
rect 8033 4233 8067 4267
rect 8585 4233 8619 4267
rect 8953 4233 8987 4267
rect 13093 4233 13127 4267
rect 17509 4233 17543 4267
rect 18061 4233 18095 4267
rect 18429 4233 18463 4267
rect 18889 4233 18923 4267
rect 19349 4233 19383 4267
rect 22937 4233 22971 4267
rect 23213 4233 23247 4267
rect 25421 4233 25455 4267
rect 3525 4165 3559 4199
rect 10701 4165 10735 4199
rect 20453 4165 20487 4199
rect 3249 4097 3283 4131
rect 3709 4097 3743 4131
rect 6193 4097 6227 4131
rect 17601 4097 17635 4131
rect 20545 4097 20579 4131
rect 21649 4097 21683 4131
rect 23121 4097 23155 4131
rect 23949 4097 23983 4131
rect 2053 4029 2087 4063
rect 2421 4029 2455 4063
rect 2605 4029 2639 4063
rect 3801 4029 3835 4063
rect 3985 4029 4019 4063
rect 4169 4029 4203 4063
rect 4813 4029 4847 4063
rect 5089 4029 5123 4063
rect 5365 4029 5399 4063
rect 5641 4029 5675 4063
rect 6377 4029 6411 4063
rect 6745 4029 6779 4063
rect 7021 4029 7055 4063
rect 7297 4029 7331 4063
rect 8585 4029 8619 4063
rect 8769 4029 8803 4063
rect 10250 4029 10284 4063
rect 10517 4029 10551 4063
rect 10609 4029 10643 4063
rect 11713 4029 11747 4063
rect 11897 4029 11931 4063
rect 13553 4029 13587 4063
rect 13921 4029 13955 4063
rect 15301 4029 15335 4063
rect 15577 4029 15611 4063
rect 16037 4029 16071 4063
rect 16129 4029 16163 4063
rect 16405 4029 16439 4063
rect 17325 4029 17359 4063
rect 17509 4029 17543 4063
rect 17785 4029 17819 4063
rect 18061 4029 18095 4063
rect 18153 4029 18187 4063
rect 19165 4029 19199 4063
rect 19717 4029 19751 4063
rect 19901 4029 19935 4063
rect 20085 4029 20119 4063
rect 20637 4029 20671 4063
rect 20821 4029 20855 4063
rect 20913 4029 20947 4063
rect 21311 4029 21345 4063
rect 21465 4029 21499 4063
rect 21557 4029 21591 4063
rect 21741 4029 21775 4063
rect 21833 4029 21867 4063
rect 22109 4029 22143 4063
rect 22477 4029 22511 4063
rect 22753 4029 22787 4063
rect 23305 4029 23339 4063
rect 24225 4029 24259 4063
rect 25053 4029 25087 4063
rect 25237 4029 25271 4063
rect 26810 4029 26844 4063
rect 27077 4029 27111 4063
rect 2789 3961 2823 3995
rect 4261 3961 4295 3995
rect 4461 3961 4495 3995
rect 6101 3961 6135 3995
rect 12909 3961 12943 3995
rect 13125 3961 13159 3995
rect 18705 3961 18739 3995
rect 22293 3961 22327 3995
rect 23029 3961 23063 3995
rect 2145 3893 2179 3927
rect 4905 3893 4939 3927
rect 5273 3893 5307 3927
rect 5457 3893 5491 3927
rect 5825 3893 5859 3927
rect 6929 3893 6963 3927
rect 9137 3893 9171 3927
rect 11805 3893 11839 3927
rect 13277 3893 13311 3927
rect 13645 3893 13679 3927
rect 14105 3893 14139 3927
rect 15485 3893 15519 3927
rect 15761 3893 15795 3927
rect 17141 3893 17175 3927
rect 17969 3893 18003 3927
rect 18905 3893 18939 3927
rect 19073 3893 19107 3927
rect 19809 3893 19843 3927
rect 21097 3893 21131 3927
rect 21925 3893 21959 3927
rect 22569 3893 22603 3927
rect 23489 3893 23523 3927
rect 24961 3893 24995 3927
rect 25697 3893 25731 3927
rect 3065 3689 3099 3723
rect 5089 3689 5123 3723
rect 6561 3689 6595 3723
rect 10701 3689 10735 3723
rect 13645 3689 13679 3723
rect 14933 3689 14967 3723
rect 15485 3689 15519 3723
rect 18061 3689 18095 3723
rect 23857 3689 23891 3723
rect 3709 3621 3743 3655
rect 5273 3621 5307 3655
rect 11713 3621 11747 3655
rect 13277 3621 13311 3655
rect 14013 3621 14047 3655
rect 15025 3621 15059 3655
rect 23029 3621 23063 3655
rect 2973 3553 3007 3587
rect 3157 3553 3191 3587
rect 3341 3553 3375 3587
rect 3434 3553 3468 3587
rect 4077 3553 4111 3587
rect 4261 3553 4295 3587
rect 4353 3553 4387 3587
rect 4537 3553 4571 3587
rect 4721 3553 4755 3587
rect 4905 3553 4939 3587
rect 5181 3553 5215 3587
rect 5457 3553 5491 3587
rect 5641 3553 5675 3587
rect 6101 3553 6135 3587
rect 6377 3553 6411 3587
rect 6653 3553 6687 3587
rect 7113 3553 7147 3587
rect 8677 3553 8711 3587
rect 8861 3553 8895 3587
rect 9137 3553 9171 3587
rect 9321 3553 9355 3587
rect 10609 3553 10643 3587
rect 10793 3553 10827 3587
rect 11528 3553 11562 3587
rect 11621 3553 11655 3587
rect 12449 3553 12483 3587
rect 12909 3553 12943 3587
rect 13093 3553 13127 3587
rect 13185 3553 13219 3587
rect 13369 3553 13403 3587
rect 13569 3575 13603 3609
rect 13829 3553 13863 3587
rect 14473 3553 14507 3587
rect 14565 3553 14599 3587
rect 14749 3553 14783 3587
rect 15301 3553 15335 3587
rect 15577 3553 15611 3587
rect 15761 3553 15795 3587
rect 16129 3553 16163 3587
rect 17785 3553 17819 3587
rect 17877 3553 17911 3587
rect 19533 3553 19567 3587
rect 19717 3553 19751 3587
rect 21373 3553 21407 3587
rect 21557 3553 21591 3587
rect 21649 3553 21683 3587
rect 21833 3553 21867 3587
rect 22109 3553 22143 3587
rect 22201 3553 22235 3587
rect 22661 3553 22695 3587
rect 22845 3553 22879 3587
rect 23121 3553 23155 3587
rect 23305 3553 23339 3587
rect 23673 3553 23707 3587
rect 23949 3553 23983 3587
rect 25421 3553 25455 3587
rect 25605 3553 25639 3587
rect 6193 3485 6227 3519
rect 6745 3485 6779 3519
rect 12173 3485 12207 3519
rect 12633 3485 12667 3519
rect 13001 3485 13035 3519
rect 15117 3485 15151 3519
rect 15945 3485 15979 3519
rect 16221 3485 16255 3519
rect 18061 3485 18095 3519
rect 25513 3485 25547 3519
rect 4537 3417 4571 3451
rect 7021 3417 7055 3451
rect 11989 3417 12023 3451
rect 23489 3417 23523 3451
rect 24133 3417 24167 3451
rect 4169 3349 4203 3383
rect 4905 3349 4939 3383
rect 6377 3349 6411 3383
rect 6653 3349 6687 3383
rect 7297 3349 7331 3383
rect 7481 3349 7515 3383
rect 9045 3349 9079 3383
rect 9229 3349 9263 3383
rect 11437 3349 11471 3383
rect 12265 3349 12299 3383
rect 15117 3349 15151 3383
rect 16129 3349 16163 3383
rect 16497 3349 16531 3383
rect 19625 3349 19659 3383
rect 21465 3349 21499 3383
rect 21741 3349 21775 3383
rect 22109 3349 22143 3383
rect 22477 3349 22511 3383
rect 23121 3349 23155 3383
rect 24225 3349 24259 3383
rect 6009 3145 6043 3179
rect 8217 3145 8251 3179
rect 8585 3145 8619 3179
rect 11897 3145 11931 3179
rect 13829 3145 13863 3179
rect 14197 3145 14231 3179
rect 14289 3145 14323 3179
rect 15485 3145 15519 3179
rect 15669 3145 15703 3179
rect 17877 3145 17911 3179
rect 18245 3145 18279 3179
rect 25513 3145 25547 3179
rect 26341 3145 26375 3179
rect 10701 3077 10735 3111
rect 17233 3077 17267 3111
rect 24961 3077 24995 3111
rect 3801 3009 3835 3043
rect 7205 3009 7239 3043
rect 9965 3009 9999 3043
rect 11161 3009 11195 3043
rect 15301 3009 15335 3043
rect 19441 3009 19475 3043
rect 20453 3009 20487 3043
rect 22109 3009 22143 3043
rect 23949 3009 23983 3043
rect 1685 2941 1719 2975
rect 1869 2941 1903 2975
rect 1961 2941 1995 2975
rect 2145 2941 2179 2975
rect 2237 2941 2271 2975
rect 2421 2941 2455 2975
rect 2697 2941 2731 2975
rect 2881 2941 2915 2975
rect 3433 2941 3467 2975
rect 6193 2941 6227 2975
rect 6377 2941 6411 2975
rect 6469 2941 6503 2975
rect 6653 2941 6687 2975
rect 6745 2941 6779 2975
rect 6929 2941 6963 2975
rect 7481 2941 7515 2975
rect 10241 2941 10275 2975
rect 10425 2941 10459 2975
rect 10517 2941 10551 2975
rect 10701 2941 10735 2975
rect 10793 2941 10827 2975
rect 10977 2941 11011 2975
rect 11069 2941 11103 2975
rect 11253 2941 11287 2975
rect 11713 2941 11747 2975
rect 12541 2941 12575 2975
rect 12725 2941 12759 2975
rect 12817 2941 12851 2975
rect 13001 2941 13035 2975
rect 13829 2941 13863 2975
rect 13921 2941 13955 2975
rect 14289 2941 14323 2975
rect 14473 2941 14507 2975
rect 14565 2941 14599 2975
rect 14749 2941 14783 2975
rect 15485 2941 15519 2975
rect 15945 2941 15979 2975
rect 16221 2941 16255 2975
rect 16497 2941 16531 2975
rect 18153 2941 18187 2975
rect 18337 2941 18371 2975
rect 19073 2941 19107 2975
rect 19257 2941 19291 2975
rect 19349 2941 19383 2975
rect 19533 2941 19567 2975
rect 19625 2941 19659 2975
rect 19809 2941 19843 2975
rect 19901 2941 19935 2975
rect 20085 2941 20119 2975
rect 20367 2941 20401 2975
rect 20545 2941 20579 2975
rect 21097 2941 21131 2975
rect 22017 2941 22051 2975
rect 22201 2941 22235 2975
rect 22293 2941 22327 2975
rect 22477 2941 22511 2975
rect 22569 2941 22603 2975
rect 22753 2941 22787 2975
rect 23397 2941 23431 2975
rect 24225 2941 24259 2975
rect 25237 2941 25271 2975
rect 25973 2941 26007 2975
rect 26249 2941 26283 2975
rect 26433 2941 26467 2975
rect 2329 2873 2363 2907
rect 3617 2873 3651 2907
rect 5641 2873 5675 2907
rect 5825 2873 5859 2907
rect 6837 2873 6871 2907
rect 9698 2873 9732 2907
rect 11529 2873 11563 2907
rect 15209 2873 15243 2907
rect 18061 2873 18095 2907
rect 20913 2873 20947 2907
rect 22385 2873 22419 2907
rect 25697 2873 25731 2907
rect 26157 2873 26191 2907
rect 1777 2805 1811 2839
rect 2053 2805 2087 2839
rect 2789 2805 2823 2839
rect 6285 2805 6319 2839
rect 6561 2805 6595 2839
rect 10333 2805 10367 2839
rect 10885 2805 10919 2839
rect 12725 2805 12759 2839
rect 12909 2805 12943 2839
rect 14657 2805 14691 2839
rect 16129 2805 16163 2839
rect 17693 2805 17727 2839
rect 17861 2805 17895 2839
rect 19165 2805 19199 2839
rect 19717 2805 19751 2839
rect 19993 2805 20027 2839
rect 20729 2805 20763 2839
rect 22661 2805 22695 2839
rect 25053 2805 25087 2839
rect 25329 2805 25363 2839
rect 25497 2805 25531 2839
rect 25789 2805 25823 2839
rect 5089 2601 5123 2635
rect 6193 2601 6227 2635
rect 6745 2601 6779 2635
rect 8887 2601 8921 2635
rect 9045 2601 9079 2635
rect 9321 2601 9355 2635
rect 13737 2601 13771 2635
rect 15301 2601 15335 2635
rect 18245 2601 18279 2635
rect 22201 2601 22235 2635
rect 22477 2601 22511 2635
rect 23213 2601 23247 2635
rect 25881 2601 25915 2635
rect 6009 2533 6043 2567
rect 8677 2533 8711 2567
rect 14657 2533 14691 2567
rect 15117 2533 15151 2567
rect 18337 2533 18371 2567
rect 18521 2533 18555 2567
rect 23029 2533 23063 2567
rect 24768 2533 24802 2567
rect 2513 2465 2547 2499
rect 2697 2465 2731 2499
rect 3433 2465 3467 2499
rect 3617 2465 3651 2499
rect 4353 2465 4387 2499
rect 4537 2465 4571 2499
rect 4629 2465 4663 2499
rect 4813 2465 4847 2499
rect 4997 2465 5031 2499
rect 5181 2465 5215 2499
rect 5365 2465 5399 2499
rect 5549 2465 5583 2499
rect 5825 2465 5859 2499
rect 6285 2465 6319 2499
rect 6469 2465 6503 2499
rect 6745 2465 6779 2499
rect 6929 2465 6963 2499
rect 9137 2465 9171 2499
rect 11713 2465 11747 2499
rect 11897 2465 11931 2499
rect 12173 2465 12207 2499
rect 12541 2465 12575 2499
rect 12725 2465 12759 2499
rect 12817 2465 12851 2499
rect 13001 2465 13035 2499
rect 13645 2465 13679 2499
rect 13829 2465 13863 2499
rect 14289 2465 14323 2499
rect 14473 2465 14507 2499
rect 14565 2465 14599 2499
rect 14749 2465 14783 2499
rect 14933 2465 14967 2499
rect 16221 2465 16255 2499
rect 16865 2465 16899 2499
rect 17121 2465 17155 2499
rect 20269 2465 20303 2499
rect 20545 2465 20579 2499
rect 20729 2465 20763 2499
rect 20821 2465 20855 2499
rect 21005 2465 21039 2499
rect 21281 2465 21315 2499
rect 21465 2465 21499 2499
rect 22109 2465 22143 2499
rect 22293 2465 22327 2499
rect 22385 2465 22419 2499
rect 22569 2465 22603 2499
rect 22845 2465 22879 2499
rect 23581 2465 23615 2499
rect 24409 2465 24443 2499
rect 24501 2465 24535 2499
rect 18705 2397 18739 2431
rect 23305 2397 23339 2431
rect 2697 2329 2731 2363
rect 6469 2329 6503 2363
rect 12817 2329 12851 2363
rect 20545 2329 20579 2363
rect 3617 2261 3651 2295
rect 4077 2261 4111 2295
rect 4537 2261 4571 2295
rect 4813 2261 4847 2295
rect 5549 2261 5583 2295
rect 7021 2261 7055 2295
rect 8861 2261 8895 2295
rect 10333 2261 10367 2295
rect 11897 2261 11931 2295
rect 11989 2261 12023 2295
rect 12725 2261 12759 2295
rect 14289 2261 14323 2295
rect 20453 2261 20487 2295
rect 21005 2261 21039 2295
rect 21281 2261 21315 2295
rect 17509 2057 17543 2091
rect 21373 2057 21407 2091
rect 4077 1921 4111 1955
rect 6745 1921 6779 1955
rect 10425 1921 10459 1955
rect 20177 1921 20211 1955
rect 949 1853 983 1887
rect 1317 1853 1351 1887
rect 1777 1853 1811 1887
rect 1869 1853 1903 1887
rect 2145 1853 2179 1887
rect 2973 1853 3007 1887
rect 3249 1853 3283 1887
rect 3709 1853 3743 1887
rect 3985 1853 4019 1887
rect 4353 1853 4387 1887
rect 5181 1853 5215 1887
rect 5273 1853 5307 1887
rect 5549 1853 5583 1887
rect 5825 1853 5859 1887
rect 6653 1853 6687 1887
rect 7021 1853 7055 1887
rect 7849 1853 7883 1887
rect 7941 1853 7975 1887
rect 9229 1853 9263 1887
rect 9321 1853 9355 1887
rect 10149 1853 10183 1887
rect 10517 1853 10551 1887
rect 10793 1853 10827 1887
rect 11621 1853 11655 1887
rect 11713 1853 11747 1887
rect 11989 1853 12023 1887
rect 12817 1853 12851 1887
rect 12909 1853 12943 1887
rect 13185 1853 13219 1887
rect 14197 1853 14231 1887
rect 14657 1853 14691 1887
rect 15117 1853 15151 1887
rect 15209 1853 15243 1887
rect 15485 1853 15519 1887
rect 16313 1853 16347 1887
rect 16405 1853 16439 1887
rect 16865 1853 16899 1887
rect 17693 1853 17727 1887
rect 18889 1853 18923 1887
rect 18981 1853 19015 1887
rect 19257 1853 19291 1887
rect 20085 1853 20119 1887
rect 20453 1853 20487 1887
rect 21281 1853 21315 1887
rect 21649 1853 21683 1887
rect 21925 1853 21959 1887
rect 22385 1853 22419 1887
rect 22661 1853 22695 1887
rect 23489 1853 23523 1887
rect 23857 1853 23891 1887
rect 24593 1853 24627 1887
rect 24869 1853 24903 1887
rect 25697 1853 25731 1887
rect 3525 1717 3559 1751
rect 949 1377 983 1411
rect 1225 1377 1259 1411
rect 2053 1377 2087 1411
rect 2421 1377 2455 1411
rect 3249 1377 3283 1411
rect 3617 1377 3651 1411
rect 4445 1377 4479 1411
rect 4537 1377 4571 1411
rect 4813 1377 4847 1411
rect 5641 1377 5675 1411
rect 5825 1377 5859 1411
rect 7113 1377 7147 1411
rect 7941 1377 7975 1411
rect 8309 1377 8343 1411
rect 9137 1377 9171 1411
rect 9873 1377 9907 1411
rect 10701 1377 10735 1411
rect 11345 1377 11379 1411
rect 12173 1377 12207 1411
rect 12541 1377 12575 1411
rect 13369 1377 13403 1411
rect 13737 1377 13771 1411
rect 14565 1377 14599 1411
rect 14657 1377 14691 1411
rect 14933 1377 14967 1411
rect 15761 1377 15795 1411
rect 16405 1377 16439 1411
rect 17233 1377 17267 1411
rect 17325 1377 17359 1411
rect 17601 1377 17635 1411
rect 18429 1377 18463 1411
rect 18521 1377 18555 1411
rect 19349 1377 19383 1411
rect 19993 1377 20027 1411
rect 20821 1377 20855 1411
rect 21281 1377 21315 1411
rect 21557 1377 21591 1411
rect 22385 1377 22419 1411
rect 22753 1377 22787 1411
rect 23581 1377 23615 1411
rect 23949 1377 23983 1411
rect 24777 1377 24811 1411
rect 25145 1377 25179 1411
rect 25973 1377 26007 1411
rect 2145 1309 2179 1343
rect 3341 1309 3375 1343
rect 6837 1309 6871 1343
rect 8033 1309 8067 1343
rect 9505 1309 9539 1343
rect 9597 1309 9631 1343
rect 11069 1309 11103 1343
rect 12265 1309 12299 1343
rect 13461 1309 13495 1343
rect 16129 1309 16163 1343
rect 19625 1309 19659 1343
rect 19717 1309 19751 1343
rect 22477 1309 22511 1343
rect 23673 1309 23707 1343
rect 24869 1309 24903 1343
rect 6285 1173 6319 1207
rect 6745 1173 6779 1207
rect 21097 1173 21131 1207
rect 2237 969 2271 1003
rect 8401 969 8435 1003
rect 10609 969 10643 1003
rect 11253 969 11287 1003
rect 11713 969 11747 1003
rect 13553 969 13587 1003
rect 15761 969 15795 1003
rect 17877 969 17911 1003
rect 18521 969 18555 1003
rect 22477 969 22511 1003
rect 22753 969 22787 1003
rect 23213 969 23247 1003
rect 25053 969 25087 1003
rect 25329 969 25363 1003
rect 949 833 983 867
rect 4445 833 4479 867
rect 5917 833 5951 867
rect 7113 833 7147 867
rect 9229 833 9263 867
rect 12265 833 12299 867
rect 14105 833 14139 867
rect 18245 833 18279 867
rect 18705 833 18739 867
rect 21005 833 21039 867
rect 21281 833 21315 867
rect 23857 833 23891 867
rect 1225 765 1259 799
rect 2053 765 2087 799
rect 3065 765 3099 799
rect 3249 765 3283 799
rect 3525 765 3559 799
rect 4353 765 4387 799
rect 4721 765 4755 799
rect 5549 765 5583 799
rect 6193 765 6227 799
rect 7021 765 7055 799
rect 7389 765 7423 799
rect 8217 765 8251 799
rect 9505 765 9539 799
rect 10333 765 10367 799
rect 12541 765 12575 799
rect 13369 765 13403 799
rect 14381 765 14415 799
rect 15209 765 15243 799
rect 16221 765 16255 799
rect 16497 765 16531 799
rect 17325 765 17359 799
rect 18981 765 19015 799
rect 19809 765 19843 799
rect 19901 765 19935 799
rect 20729 765 20763 799
rect 21557 765 21591 799
rect 22385 765 22419 799
rect 24133 765 24167 799
rect 24961 765 24995 799
<< metal1 >>
rect 13446 31152 13452 31204
rect 13504 31192 13510 31204
rect 21082 31192 21088 31204
rect 13504 31164 21088 31192
rect 13504 31152 13510 31164
rect 21082 31152 21088 31164
rect 21140 31152 21146 31204
rect 19426 31084 19432 31136
rect 19484 31124 19490 31136
rect 22738 31124 22744 31136
rect 19484 31096 22744 31124
rect 19484 31084 19490 31096
rect 22738 31084 22744 31096
rect 22796 31084 22802 31136
rect 552 31034 27576 31056
rect 552 30982 7114 31034
rect 7166 30982 7178 31034
rect 7230 30982 7242 31034
rect 7294 30982 7306 31034
rect 7358 30982 7370 31034
rect 7422 30982 13830 31034
rect 13882 30982 13894 31034
rect 13946 30982 13958 31034
rect 14010 30982 14022 31034
rect 14074 30982 14086 31034
rect 14138 30982 20546 31034
rect 20598 30982 20610 31034
rect 20662 30982 20674 31034
rect 20726 30982 20738 31034
rect 20790 30982 20802 31034
rect 20854 30982 27262 31034
rect 27314 30982 27326 31034
rect 27378 30982 27390 31034
rect 27442 30982 27454 31034
rect 27506 30982 27518 31034
rect 27570 30982 27576 31034
rect 552 30960 27576 30982
rect 937 30923 995 30929
rect 937 30889 949 30923
rect 983 30920 995 30923
rect 1394 30920 1400 30932
rect 983 30892 1400 30920
rect 983 30889 995 30892
rect 937 30883 995 30889
rect 1394 30880 1400 30892
rect 1452 30880 1458 30932
rect 5810 30880 5816 30932
rect 5868 30880 5874 30932
rect 7466 30880 7472 30932
rect 7524 30880 7530 30932
rect 8754 30880 8760 30932
rect 8812 30880 8818 30932
rect 11072 30892 13124 30920
rect 2038 30744 2044 30796
rect 2096 30793 2102 30796
rect 2096 30787 2119 30793
rect 2107 30753 2119 30787
rect 2096 30747 2119 30753
rect 2096 30744 2102 30747
rect 3510 30744 3516 30796
rect 3568 30784 3574 30796
rect 3881 30787 3939 30793
rect 3881 30784 3893 30787
rect 3568 30756 3893 30784
rect 3568 30744 3574 30756
rect 3881 30753 3893 30756
rect 3927 30753 3939 30787
rect 5828 30784 5856 30880
rect 6089 30787 6147 30793
rect 6089 30784 6101 30787
rect 5828 30756 6101 30784
rect 3881 30747 3939 30753
rect 6089 30753 6101 30756
rect 6135 30753 6147 30787
rect 7484 30784 7512 30880
rect 7561 30787 7619 30793
rect 7561 30784 7573 30787
rect 7484 30756 7573 30784
rect 6089 30747 6147 30753
rect 7561 30753 7573 30756
rect 7607 30753 7619 30787
rect 7561 30747 7619 30753
rect 8573 30787 8631 30793
rect 8573 30753 8585 30787
rect 8619 30753 8631 30787
rect 8772 30784 8800 30880
rect 9769 30855 9827 30861
rect 9769 30821 9781 30855
rect 9815 30852 9827 30855
rect 11072 30852 11100 30892
rect 9815 30824 11100 30852
rect 11164 30824 12572 30852
rect 9815 30821 9827 30824
rect 9769 30815 9827 30821
rect 8849 30787 8907 30793
rect 8849 30784 8861 30787
rect 8772 30756 8861 30784
rect 8573 30747 8631 30753
rect 8849 30753 8861 30756
rect 8895 30753 8907 30787
rect 8849 30747 8907 30753
rect 9493 30787 9551 30793
rect 9493 30753 9505 30787
rect 9539 30753 9551 30787
rect 9493 30747 9551 30753
rect 2314 30676 2320 30728
rect 2372 30676 2378 30728
rect 8588 30716 8616 30747
rect 9508 30716 9536 30747
rect 9674 30744 9680 30796
rect 9732 30744 9738 30796
rect 9858 30744 9864 30796
rect 9916 30744 9922 30796
rect 10318 30744 10324 30796
rect 10376 30784 10382 30796
rect 10965 30787 11023 30793
rect 10965 30784 10977 30787
rect 10376 30756 10977 30784
rect 10376 30744 10382 30756
rect 10965 30753 10977 30756
rect 11011 30753 11023 30787
rect 10965 30747 11023 30753
rect 10137 30719 10195 30725
rect 10137 30716 10149 30719
rect 8588 30688 8800 30716
rect 9508 30688 10149 30716
rect 8772 30592 8800 30688
rect 10137 30685 10149 30688
rect 10183 30685 10195 30719
rect 10137 30679 10195 30685
rect 10226 30676 10232 30728
rect 10284 30716 10290 30728
rect 10689 30719 10747 30725
rect 10689 30716 10701 30719
rect 10284 30688 10701 30716
rect 10284 30676 10290 30688
rect 10689 30685 10701 30688
rect 10735 30685 10747 30719
rect 10689 30679 10747 30685
rect 10045 30651 10103 30657
rect 10045 30617 10057 30651
rect 10091 30648 10103 30651
rect 11054 30648 11060 30660
rect 10091 30620 11060 30648
rect 10091 30617 10103 30620
rect 10045 30611 10103 30617
rect 11054 30608 11060 30620
rect 11112 30608 11118 30660
rect 11164 30657 11192 30824
rect 11698 30744 11704 30796
rect 11756 30784 11762 30796
rect 12544 30793 12572 30824
rect 11977 30787 12035 30793
rect 11977 30784 11989 30787
rect 11756 30756 11989 30784
rect 11756 30744 11762 30756
rect 11977 30753 11989 30756
rect 12023 30753 12035 30787
rect 11977 30747 12035 30753
rect 12345 30787 12403 30793
rect 12345 30753 12357 30787
rect 12391 30753 12403 30787
rect 12345 30747 12403 30753
rect 12529 30787 12587 30793
rect 12529 30753 12541 30787
rect 12575 30784 12587 30787
rect 12710 30784 12716 30796
rect 12575 30756 12716 30784
rect 12575 30753 12587 30756
rect 12529 30747 12587 30753
rect 11238 30676 11244 30728
rect 11296 30676 11302 30728
rect 11790 30676 11796 30728
rect 11848 30676 11854 30728
rect 12360 30716 12388 30747
rect 12710 30744 12716 30756
rect 12768 30744 12774 30796
rect 12434 30716 12440 30728
rect 12360 30688 12440 30716
rect 12406 30676 12440 30688
rect 12492 30676 12498 30728
rect 13096 30716 13124 30892
rect 16114 30880 16120 30932
rect 16172 30880 16178 30932
rect 19628 30892 20392 30920
rect 13170 30744 13176 30796
rect 13228 30784 13234 30796
rect 14277 30787 14335 30793
rect 14277 30784 14289 30787
rect 13228 30756 14289 30784
rect 13228 30744 13234 30756
rect 14277 30753 14289 30756
rect 14323 30753 14335 30787
rect 14277 30747 14335 30753
rect 14642 30744 14648 30796
rect 14700 30784 14706 30796
rect 14737 30787 14795 30793
rect 14737 30784 14749 30787
rect 14700 30756 14749 30784
rect 14700 30744 14706 30756
rect 14737 30753 14749 30756
rect 14783 30753 14795 30787
rect 14737 30747 14795 30753
rect 15286 30744 15292 30796
rect 15344 30744 15350 30796
rect 16132 30784 16160 30880
rect 19628 30864 19656 30892
rect 17586 30812 17592 30864
rect 17644 30852 17650 30864
rect 17865 30855 17923 30861
rect 17865 30852 17877 30855
rect 17644 30824 17877 30852
rect 17644 30812 17650 30824
rect 17865 30821 17877 30824
rect 17911 30821 17923 30855
rect 17865 30815 17923 30821
rect 17972 30824 19564 30852
rect 16209 30787 16267 30793
rect 16209 30784 16221 30787
rect 16132 30756 16221 30784
rect 16209 30753 16221 30756
rect 16255 30753 16267 30787
rect 16209 30747 16267 30753
rect 16758 30744 16764 30796
rect 16816 30784 16822 30796
rect 16945 30787 17003 30793
rect 16945 30784 16957 30787
rect 16816 30756 16957 30784
rect 16816 30744 16822 30756
rect 16945 30753 16957 30756
rect 16991 30753 17003 30787
rect 16945 30747 17003 30753
rect 13096 30688 13676 30716
rect 11149 30651 11207 30657
rect 11149 30617 11161 30651
rect 11195 30617 11207 30651
rect 12406 30648 12434 30676
rect 13648 30660 13676 30688
rect 14090 30676 14096 30728
rect 14148 30676 14154 30728
rect 17972 30716 18000 30824
rect 18046 30744 18052 30796
rect 18104 30744 18110 30796
rect 19426 30744 19432 30796
rect 19484 30744 19490 30796
rect 19536 30793 19564 30824
rect 19610 30812 19616 30864
rect 19668 30812 19674 30864
rect 19702 30812 19708 30864
rect 19760 30812 19766 30864
rect 20257 30855 20315 30861
rect 20257 30852 20269 30855
rect 19812 30824 20269 30852
rect 19521 30787 19579 30793
rect 19521 30753 19533 30787
rect 19567 30784 19579 30787
rect 19720 30784 19748 30812
rect 19812 30793 19840 30824
rect 20257 30821 20269 30824
rect 20303 30821 20315 30855
rect 20364 30852 20392 30892
rect 21082 30880 21088 30932
rect 21140 30920 21146 30932
rect 21140 30892 23428 30920
rect 21140 30880 21146 30892
rect 23400 30861 23428 30892
rect 23474 30880 23480 30932
rect 23532 30880 23538 30932
rect 26418 30880 26424 30932
rect 26476 30880 26482 30932
rect 23385 30855 23443 30861
rect 20364 30824 22692 30852
rect 20257 30815 20315 30821
rect 19567 30756 19748 30784
rect 19797 30787 19855 30793
rect 19567 30753 19579 30756
rect 19521 30747 19579 30753
rect 19797 30753 19809 30787
rect 19843 30753 19855 30787
rect 19797 30747 19855 30753
rect 19981 30787 20039 30793
rect 19981 30753 19993 30787
rect 20027 30753 20039 30787
rect 19981 30747 20039 30753
rect 21545 30787 21603 30793
rect 21545 30753 21557 30787
rect 21591 30784 21603 30787
rect 22002 30784 22008 30796
rect 21591 30756 22008 30784
rect 21591 30753 21603 30756
rect 21545 30747 21603 30753
rect 14476 30688 18000 30716
rect 11149 30611 11207 30617
rect 11256 30620 12434 30648
rect 3602 30540 3608 30592
rect 3660 30580 3666 30592
rect 3697 30583 3755 30589
rect 3697 30580 3709 30583
rect 3660 30552 3709 30580
rect 3660 30540 3666 30552
rect 3697 30549 3709 30552
rect 3743 30549 3755 30583
rect 3697 30543 3755 30549
rect 5902 30540 5908 30592
rect 5960 30540 5966 30592
rect 7374 30540 7380 30592
rect 7432 30540 7438 30592
rect 8478 30540 8484 30592
rect 8536 30540 8542 30592
rect 8754 30540 8760 30592
rect 8812 30540 8818 30592
rect 9033 30583 9091 30589
rect 9033 30549 9045 30583
rect 9079 30580 9091 30583
rect 11256 30580 11284 30620
rect 13630 30608 13636 30660
rect 13688 30648 13694 30660
rect 14476 30657 14504 30688
rect 19058 30676 19064 30728
rect 19116 30716 19122 30728
rect 19996 30716 20024 30747
rect 22002 30744 22008 30756
rect 22060 30744 22066 30796
rect 19116 30688 20024 30716
rect 19116 30676 19122 30688
rect 20806 30676 20812 30728
rect 20864 30676 20870 30728
rect 21726 30676 21732 30728
rect 21784 30676 21790 30728
rect 22462 30676 22468 30728
rect 22520 30676 22526 30728
rect 22664 30716 22692 30824
rect 23385 30821 23397 30855
rect 23431 30821 23443 30855
rect 23492 30852 23520 30880
rect 23492 30824 23888 30852
rect 23385 30815 23443 30821
rect 22738 30744 22744 30796
rect 22796 30784 22802 30796
rect 23860 30793 23888 30824
rect 23293 30787 23351 30793
rect 23293 30784 23305 30787
rect 22796 30756 23305 30784
rect 22796 30744 22802 30756
rect 23293 30753 23305 30756
rect 23339 30753 23351 30787
rect 23293 30747 23351 30753
rect 23477 30787 23535 30793
rect 23477 30753 23489 30787
rect 23523 30753 23535 30787
rect 23477 30747 23535 30753
rect 23661 30787 23719 30793
rect 23661 30753 23673 30787
rect 23707 30753 23719 30787
rect 23661 30747 23719 30753
rect 23845 30787 23903 30793
rect 23845 30753 23857 30787
rect 23891 30753 23903 30787
rect 26436 30784 26464 30880
rect 26697 30787 26755 30793
rect 26697 30784 26709 30787
rect 26436 30756 26709 30784
rect 23845 30747 23903 30753
rect 26697 30753 26709 30756
rect 26743 30753 26755 30787
rect 26697 30747 26755 30753
rect 23198 30716 23204 30728
rect 22664 30688 23204 30716
rect 23198 30676 23204 30688
rect 23256 30716 23262 30728
rect 23492 30716 23520 30747
rect 23256 30688 23520 30716
rect 23256 30676 23262 30688
rect 14461 30651 14519 30657
rect 14461 30648 14473 30651
rect 13688 30620 14473 30648
rect 13688 30608 13694 30620
rect 14461 30617 14473 30620
rect 14507 30617 14519 30651
rect 14461 30611 14519 30617
rect 14550 30608 14556 30660
rect 14608 30648 14614 30660
rect 17129 30651 17187 30657
rect 14608 30620 15148 30648
rect 14608 30608 14614 30620
rect 9079 30552 11284 30580
rect 9079 30549 9091 30552
rect 9033 30543 9091 30549
rect 12158 30540 12164 30592
rect 12216 30540 12222 30592
rect 12437 30583 12495 30589
rect 12437 30549 12449 30583
rect 12483 30580 12495 30583
rect 12618 30580 12624 30592
rect 12483 30552 12624 30580
rect 12483 30549 12495 30552
rect 12437 30543 12495 30549
rect 12618 30540 12624 30552
rect 12676 30540 12682 30592
rect 13538 30540 13544 30592
rect 13596 30540 13602 30592
rect 14642 30540 14648 30592
rect 14700 30580 14706 30592
rect 15120 30589 15148 30620
rect 17129 30617 17141 30651
rect 17175 30648 17187 30651
rect 18138 30648 18144 30660
rect 17175 30620 18144 30648
rect 17175 30617 17187 30620
rect 17129 30611 17187 30617
rect 18138 30608 18144 30620
rect 18196 30608 18202 30660
rect 22281 30651 22339 30657
rect 22281 30617 22293 30651
rect 22327 30648 22339 30651
rect 23676 30648 23704 30747
rect 22327 30620 23704 30648
rect 22327 30617 22339 30620
rect 22281 30611 22339 30617
rect 14921 30583 14979 30589
rect 14921 30580 14933 30583
rect 14700 30552 14933 30580
rect 14700 30540 14706 30552
rect 14921 30549 14933 30552
rect 14967 30549 14979 30583
rect 14921 30543 14979 30549
rect 15105 30583 15163 30589
rect 15105 30549 15117 30583
rect 15151 30549 15163 30583
rect 15105 30543 15163 30549
rect 16390 30540 16396 30592
rect 16448 30540 16454 30592
rect 17770 30540 17776 30592
rect 17828 30540 17834 30592
rect 18230 30540 18236 30592
rect 18288 30540 18294 30592
rect 19245 30583 19303 30589
rect 19245 30549 19257 30583
rect 19291 30580 19303 30583
rect 19518 30580 19524 30592
rect 19291 30552 19524 30580
rect 19291 30549 19303 30552
rect 19245 30543 19303 30549
rect 19518 30540 19524 30552
rect 19576 30540 19582 30592
rect 20070 30540 20076 30592
rect 20128 30540 20134 30592
rect 21358 30540 21364 30592
rect 21416 30540 21422 30592
rect 23014 30540 23020 30592
rect 23072 30540 23078 30592
rect 23106 30540 23112 30592
rect 23164 30540 23170 30592
rect 23566 30540 23572 30592
rect 23624 30580 23630 30592
rect 24029 30583 24087 30589
rect 24029 30580 24041 30583
rect 23624 30552 24041 30580
rect 23624 30540 23630 30552
rect 24029 30549 24041 30552
rect 24075 30549 24087 30583
rect 24029 30543 24087 30549
rect 26510 30540 26516 30592
rect 26568 30540 26574 30592
rect 552 30490 27416 30512
rect 552 30438 3756 30490
rect 3808 30438 3820 30490
rect 3872 30438 3884 30490
rect 3936 30438 3948 30490
rect 4000 30438 4012 30490
rect 4064 30438 10472 30490
rect 10524 30438 10536 30490
rect 10588 30438 10600 30490
rect 10652 30438 10664 30490
rect 10716 30438 10728 30490
rect 10780 30438 17188 30490
rect 17240 30438 17252 30490
rect 17304 30438 17316 30490
rect 17368 30438 17380 30490
rect 17432 30438 17444 30490
rect 17496 30438 23904 30490
rect 23956 30438 23968 30490
rect 24020 30438 24032 30490
rect 24084 30438 24096 30490
rect 24148 30438 24160 30490
rect 24212 30438 27416 30490
rect 552 30416 27416 30438
rect 5721 30379 5779 30385
rect 5721 30345 5733 30379
rect 5767 30376 5779 30379
rect 5902 30376 5908 30388
rect 5767 30348 5908 30376
rect 5767 30345 5779 30348
rect 5721 30339 5779 30345
rect 2866 30268 2872 30320
rect 2924 30308 2930 30320
rect 2961 30311 3019 30317
rect 2961 30308 2973 30311
rect 2924 30280 2973 30308
rect 2924 30268 2930 30280
rect 2961 30277 2973 30280
rect 3007 30277 3019 30311
rect 2961 30271 3019 30277
rect 5169 30311 5227 30317
rect 5169 30277 5181 30311
rect 5215 30308 5227 30311
rect 5736 30308 5764 30339
rect 5902 30336 5908 30348
rect 5960 30336 5966 30388
rect 13173 30379 13231 30385
rect 6012 30348 7420 30376
rect 5215 30280 5764 30308
rect 5215 30277 5227 30280
rect 5169 30271 5227 30277
rect 4801 30243 4859 30249
rect 4801 30209 4813 30243
rect 4847 30240 4859 30243
rect 6012 30240 6040 30348
rect 7392 30320 7420 30348
rect 13173 30345 13185 30379
rect 13219 30376 13231 30379
rect 13262 30376 13268 30388
rect 13219 30348 13268 30376
rect 13219 30345 13231 30348
rect 13173 30339 13231 30345
rect 13262 30336 13268 30348
rect 13320 30336 13326 30388
rect 14090 30376 14096 30388
rect 13832 30348 14096 30376
rect 6089 30311 6147 30317
rect 6089 30277 6101 30311
rect 6135 30277 6147 30311
rect 6089 30271 6147 30277
rect 4847 30212 6040 30240
rect 4847 30209 4859 30212
rect 4801 30203 4859 30209
rect 1581 30175 1639 30181
rect 1581 30141 1593 30175
rect 1627 30172 1639 30175
rect 2314 30172 2320 30184
rect 1627 30144 2320 30172
rect 1627 30141 1639 30144
rect 1581 30135 1639 30141
rect 1780 30048 1808 30144
rect 2314 30132 2320 30144
rect 2372 30172 2378 30184
rect 3329 30175 3387 30181
rect 3329 30172 3341 30175
rect 2372 30144 3341 30172
rect 2372 30132 2378 30144
rect 3329 30141 3341 30144
rect 3375 30172 3387 30175
rect 4522 30172 4528 30184
rect 3375 30144 4528 30172
rect 3375 30141 3387 30144
rect 3329 30135 3387 30141
rect 4522 30132 4528 30144
rect 4580 30132 4586 30184
rect 5828 30181 5856 30212
rect 5813 30175 5871 30181
rect 5813 30141 5825 30175
rect 5859 30141 5871 30175
rect 5813 30135 5871 30141
rect 5902 30132 5908 30184
rect 5960 30132 5966 30184
rect 6104 30172 6132 30271
rect 7374 30268 7380 30320
rect 7432 30268 7438 30320
rect 7745 30311 7803 30317
rect 7745 30308 7757 30311
rect 7576 30280 7757 30308
rect 6012 30144 6132 30172
rect 6181 30175 6239 30181
rect 1854 30113 1860 30116
rect 1848 30067 1860 30113
rect 1854 30064 1860 30067
rect 1912 30064 1918 30116
rect 3602 30113 3608 30116
rect 3596 30104 3608 30113
rect 3563 30076 3608 30104
rect 3596 30067 3608 30076
rect 3602 30064 3608 30067
rect 3660 30064 3666 30116
rect 5442 30104 5448 30116
rect 4724 30076 5448 30104
rect 1762 29996 1768 30048
rect 1820 29996 1826 30048
rect 4724 30045 4752 30076
rect 5442 30064 5448 30076
rect 5500 30064 5506 30116
rect 6012 30104 6040 30144
rect 6181 30141 6193 30175
rect 6227 30172 6239 30175
rect 6822 30172 6828 30184
rect 6227 30144 6828 30172
rect 6227 30141 6239 30144
rect 6181 30135 6239 30141
rect 6822 30132 6828 30144
rect 6880 30132 6886 30184
rect 6426 30107 6484 30113
rect 6426 30104 6438 30107
rect 6012 30076 6438 30104
rect 6426 30073 6438 30076
rect 6472 30073 6484 30107
rect 7466 30104 7472 30116
rect 6426 30067 6484 30073
rect 6656 30076 7472 30104
rect 4709 30039 4767 30045
rect 4709 30005 4721 30039
rect 4755 30005 4767 30039
rect 4709 29999 4767 30005
rect 5166 29996 5172 30048
rect 5224 30036 5230 30048
rect 5261 30039 5319 30045
rect 5261 30036 5273 30039
rect 5224 30008 5273 30036
rect 5224 29996 5230 30008
rect 5261 30005 5273 30008
rect 5307 30005 5319 30039
rect 5261 29999 5319 30005
rect 5353 30039 5411 30045
rect 5353 30005 5365 30039
rect 5399 30036 5411 30039
rect 5534 30036 5540 30048
rect 5399 30008 5540 30036
rect 5399 30005 5411 30008
rect 5353 29999 5411 30005
rect 5534 29996 5540 30008
rect 5592 29996 5598 30048
rect 5810 29996 5816 30048
rect 5868 30036 5874 30048
rect 6656 30036 6684 30076
rect 7466 30064 7472 30076
rect 7524 30064 7530 30116
rect 7576 30104 7604 30280
rect 7745 30277 7757 30280
rect 7791 30277 7803 30311
rect 7745 30271 7803 30277
rect 12986 30268 12992 30320
rect 13044 30308 13050 30320
rect 13832 30308 13860 30348
rect 14090 30336 14096 30348
rect 14148 30336 14154 30388
rect 15197 30379 15255 30385
rect 15197 30345 15209 30379
rect 15243 30376 15255 30379
rect 15654 30376 15660 30388
rect 15243 30348 15660 30376
rect 15243 30345 15255 30348
rect 15197 30339 15255 30345
rect 15654 30336 15660 30348
rect 15712 30336 15718 30388
rect 16209 30379 16267 30385
rect 16209 30345 16221 30379
rect 16255 30376 16267 30379
rect 16390 30376 16396 30388
rect 16255 30348 16396 30376
rect 16255 30345 16267 30348
rect 16209 30339 16267 30345
rect 16390 30336 16396 30348
rect 16448 30336 16454 30388
rect 20717 30379 20775 30385
rect 20717 30345 20729 30379
rect 20763 30376 20775 30379
rect 20806 30376 20812 30388
rect 20763 30348 20812 30376
rect 20763 30345 20775 30348
rect 20717 30339 20775 30345
rect 20806 30336 20812 30348
rect 20864 30336 20870 30388
rect 22462 30336 22468 30388
rect 22520 30376 22526 30388
rect 22646 30376 22652 30388
rect 22520 30348 22652 30376
rect 22520 30336 22526 30348
rect 22646 30336 22652 30348
rect 22704 30336 22710 30388
rect 26510 30336 26516 30388
rect 26568 30336 26574 30388
rect 13044 30280 13860 30308
rect 13044 30268 13050 30280
rect 17034 30268 17040 30320
rect 17092 30268 17098 30320
rect 26528 30308 26556 30336
rect 22572 30280 26556 30308
rect 12618 30200 12624 30252
rect 12676 30200 12682 30252
rect 12802 30200 12808 30252
rect 12860 30240 12866 30252
rect 13817 30243 13875 30249
rect 13817 30240 13829 30243
rect 12860 30212 13829 30240
rect 12860 30200 12866 30212
rect 13817 30209 13829 30212
rect 13863 30209 13875 30243
rect 16025 30243 16083 30249
rect 16025 30240 16037 30243
rect 13817 30203 13875 30209
rect 14844 30212 16037 30240
rect 9953 30175 10011 30181
rect 9953 30141 9965 30175
rect 9999 30172 10011 30175
rect 10962 30172 10968 30184
rect 9999 30144 10968 30172
rect 9999 30141 10011 30144
rect 9953 30135 10011 30141
rect 10962 30132 10968 30144
rect 11020 30172 11026 30184
rect 11517 30175 11575 30181
rect 11517 30172 11529 30175
rect 11020 30144 11529 30172
rect 11020 30132 11026 30144
rect 11517 30141 11529 30144
rect 11563 30172 11575 30175
rect 11609 30175 11667 30181
rect 11609 30172 11621 30175
rect 11563 30144 11621 30172
rect 11563 30141 11575 30144
rect 11517 30135 11575 30141
rect 11609 30141 11621 30144
rect 11655 30141 11667 30175
rect 12636 30172 12664 30200
rect 13078 30172 13084 30184
rect 12636 30144 13084 30172
rect 11609 30135 11667 30141
rect 13078 30132 13084 30144
rect 13136 30132 13142 30184
rect 13265 30175 13323 30181
rect 13265 30141 13277 30175
rect 13311 30172 13323 30175
rect 13538 30172 13544 30184
rect 13311 30144 13544 30172
rect 13311 30141 13323 30144
rect 13265 30135 13323 30141
rect 13538 30132 13544 30144
rect 13596 30132 13602 30184
rect 14084 30175 14142 30181
rect 14084 30141 14096 30175
rect 14130 30172 14142 30175
rect 14550 30172 14556 30184
rect 14130 30144 14556 30172
rect 14130 30141 14142 30144
rect 14084 30135 14142 30141
rect 14550 30132 14556 30144
rect 14608 30132 14614 30184
rect 14642 30132 14648 30184
rect 14700 30172 14706 30184
rect 14844 30172 14872 30212
rect 16025 30209 16037 30212
rect 16071 30240 16083 30243
rect 16942 30240 16948 30252
rect 16071 30212 16948 30240
rect 16071 30209 16083 30212
rect 16025 30203 16083 30209
rect 16942 30200 16948 30212
rect 17000 30240 17006 30252
rect 17310 30240 17316 30252
rect 17000 30212 17316 30240
rect 17000 30200 17006 30212
rect 17310 30200 17316 30212
rect 17368 30200 17374 30252
rect 21266 30200 21272 30252
rect 21324 30200 21330 30252
rect 14700 30144 14872 30172
rect 15473 30175 15531 30181
rect 14700 30132 14706 30144
rect 15473 30141 15485 30175
rect 15519 30141 15531 30175
rect 15473 30135 15531 30141
rect 16301 30175 16359 30181
rect 16301 30141 16313 30175
rect 16347 30141 16359 30175
rect 16301 30135 16359 30141
rect 8018 30104 8024 30116
rect 7576 30076 8024 30104
rect 5868 30008 6684 30036
rect 5868 29996 5874 30008
rect 6730 29996 6736 30048
rect 6788 30036 6794 30048
rect 7576 30045 7604 30076
rect 8018 30064 8024 30076
rect 8076 30064 8082 30116
rect 8113 30107 8171 30113
rect 8113 30073 8125 30107
rect 8159 30104 8171 30107
rect 8159 30076 8616 30104
rect 8159 30073 8171 30076
rect 8113 30067 8171 30073
rect 7561 30039 7619 30045
rect 7561 30036 7573 30039
rect 6788 30008 7573 30036
rect 6788 29996 6794 30008
rect 7561 30005 7573 30008
rect 7607 30005 7619 30039
rect 7561 29999 7619 30005
rect 7650 29996 7656 30048
rect 7708 29996 7714 30048
rect 8588 30045 8616 30076
rect 8662 30064 8668 30116
rect 8720 30104 8726 30116
rect 9686 30107 9744 30113
rect 9686 30104 9698 30107
rect 8720 30076 9698 30104
rect 8720 30064 8726 30076
rect 9686 30073 9698 30076
rect 9732 30073 9744 30107
rect 9686 30067 9744 30073
rect 11054 30064 11060 30116
rect 11112 30104 11118 30116
rect 11250 30107 11308 30113
rect 11250 30104 11262 30107
rect 11112 30076 11262 30104
rect 11112 30064 11118 30076
rect 11250 30073 11262 30076
rect 11296 30073 11308 30107
rect 11250 30067 11308 30073
rect 11876 30107 11934 30113
rect 11876 30073 11888 30107
rect 11922 30104 11934 30107
rect 13722 30104 13728 30116
rect 11922 30076 13728 30104
rect 11922 30073 11934 30076
rect 11876 30067 11934 30073
rect 13722 30064 13728 30076
rect 13780 30064 13786 30116
rect 14274 30064 14280 30116
rect 14332 30104 14338 30116
rect 14332 30076 14964 30104
rect 14332 30064 14338 30076
rect 8573 30039 8631 30045
rect 8573 30005 8585 30039
rect 8619 30036 8631 30039
rect 8754 30036 8760 30048
rect 8619 30008 8760 30036
rect 8619 30005 8631 30008
rect 8573 29999 8631 30005
rect 8754 29996 8760 30008
rect 8812 29996 8818 30048
rect 9582 29996 9588 30048
rect 9640 30036 9646 30048
rect 10137 30039 10195 30045
rect 10137 30036 10149 30039
rect 9640 30008 10149 30036
rect 9640 29996 9646 30008
rect 10137 30005 10149 30008
rect 10183 30036 10195 30039
rect 10226 30036 10232 30048
rect 10183 30008 10232 30036
rect 10183 30005 10195 30008
rect 10137 29999 10195 30005
rect 10226 29996 10232 30008
rect 10284 29996 10290 30048
rect 11146 29996 11152 30048
rect 11204 30036 11210 30048
rect 14642 30036 14648 30048
rect 11204 30008 14648 30036
rect 11204 29996 11210 30008
rect 14642 29996 14648 30008
rect 14700 29996 14706 30048
rect 14936 30036 14964 30076
rect 15102 30064 15108 30116
rect 15160 30104 15166 30116
rect 15381 30107 15439 30113
rect 15381 30104 15393 30107
rect 15160 30076 15393 30104
rect 15160 30064 15166 30076
rect 15381 30073 15393 30076
rect 15427 30073 15439 30107
rect 15488 30104 15516 30135
rect 15562 30104 15568 30116
rect 15488 30076 15568 30104
rect 15381 30067 15439 30073
rect 15562 30064 15568 30076
rect 15620 30104 15626 30116
rect 15620 30076 16160 30104
rect 15620 30064 15626 30076
rect 16132 30048 16160 30076
rect 15749 30039 15807 30045
rect 15749 30036 15761 30039
rect 14936 30008 15761 30036
rect 15749 30005 15761 30008
rect 15795 30005 15807 30039
rect 15749 29999 15807 30005
rect 16114 29996 16120 30048
rect 16172 29996 16178 30048
rect 16316 30036 16344 30135
rect 16390 30132 16396 30184
rect 16448 30132 16454 30184
rect 18138 30132 18144 30184
rect 18196 30181 18202 30184
rect 18196 30172 18208 30181
rect 18417 30175 18475 30181
rect 18196 30144 18241 30172
rect 18196 30135 18208 30144
rect 18417 30141 18429 30175
rect 18463 30172 18475 30175
rect 19337 30175 19395 30181
rect 19337 30172 19349 30175
rect 18463 30144 19349 30172
rect 18463 30141 18475 30144
rect 18417 30135 18475 30141
rect 19337 30141 19349 30144
rect 19383 30172 19395 30175
rect 19426 30172 19432 30184
rect 19383 30144 19432 30172
rect 19383 30141 19395 30144
rect 19337 30135 19395 30141
rect 18196 30132 18202 30135
rect 19426 30132 19432 30144
rect 19484 30132 19490 30184
rect 19604 30175 19662 30181
rect 19604 30141 19616 30175
rect 19650 30141 19662 30175
rect 19604 30135 19662 30141
rect 16574 30064 16580 30116
rect 16632 30104 16638 30116
rect 16669 30107 16727 30113
rect 16669 30104 16681 30107
rect 16632 30076 16681 30104
rect 16632 30064 16638 30076
rect 16669 30073 16681 30076
rect 16715 30073 16727 30107
rect 16669 30067 16727 30073
rect 17052 30076 19472 30104
rect 17052 30036 17080 30076
rect 16316 30008 17080 30036
rect 19444 30036 19472 30076
rect 19518 30064 19524 30116
rect 19576 30104 19582 30116
rect 19628 30104 19656 30135
rect 20438 30132 20444 30184
rect 20496 30172 20502 30184
rect 20809 30175 20867 30181
rect 20809 30172 20821 30175
rect 20496 30144 20821 30172
rect 20496 30132 20502 30144
rect 20809 30141 20821 30144
rect 20855 30141 20867 30175
rect 22572 30172 22600 30280
rect 22738 30200 22744 30252
rect 22796 30240 22802 30252
rect 22796 30212 22968 30240
rect 22796 30200 22802 30212
rect 20809 30135 20867 30141
rect 20916 30144 22600 30172
rect 20916 30104 20944 30144
rect 22646 30132 22652 30184
rect 22704 30172 22710 30184
rect 22940 30181 22968 30212
rect 23014 30200 23020 30252
rect 23072 30240 23078 30252
rect 24581 30243 24639 30249
rect 24581 30240 24593 30243
rect 23072 30212 23336 30240
rect 23072 30200 23078 30212
rect 23308 30181 23336 30212
rect 24044 30212 24593 30240
rect 24044 30181 24072 30212
rect 24581 30209 24593 30212
rect 24627 30209 24639 30243
rect 24581 30203 24639 30209
rect 22925 30175 22983 30181
rect 22704 30144 22876 30172
rect 22704 30132 22710 30144
rect 19576 30076 19656 30104
rect 20640 30076 20944 30104
rect 21536 30107 21594 30113
rect 19576 30064 19582 30076
rect 20640 30036 20668 30076
rect 21536 30073 21548 30107
rect 21582 30104 21594 30107
rect 21582 30076 22784 30104
rect 21582 30073 21594 30076
rect 21536 30067 21594 30073
rect 19444 30008 20668 30036
rect 20990 29996 20996 30048
rect 21048 29996 21054 30048
rect 22756 30045 22784 30076
rect 22741 30039 22799 30045
rect 22741 30005 22753 30039
rect 22787 30005 22799 30039
rect 22848 30036 22876 30144
rect 22925 30141 22937 30175
rect 22971 30141 22983 30175
rect 22925 30135 22983 30141
rect 23293 30175 23351 30181
rect 23293 30141 23305 30175
rect 23339 30141 23351 30175
rect 23293 30135 23351 30141
rect 23385 30175 23443 30181
rect 23385 30141 23397 30175
rect 23431 30141 23443 30175
rect 23385 30135 23443 30141
rect 24029 30175 24087 30181
rect 24029 30141 24041 30175
rect 24075 30141 24087 30175
rect 24489 30175 24547 30181
rect 24489 30172 24501 30175
rect 24029 30135 24087 30141
rect 24136 30144 24501 30172
rect 23014 30064 23020 30116
rect 23072 30064 23078 30116
rect 23109 30107 23167 30113
rect 23109 30073 23121 30107
rect 23155 30104 23167 30107
rect 23198 30104 23204 30116
rect 23155 30076 23204 30104
rect 23155 30073 23167 30076
rect 23109 30067 23167 30073
rect 23198 30064 23204 30076
rect 23256 30064 23262 30116
rect 23400 30036 23428 30135
rect 23474 30064 23480 30116
rect 23532 30104 23538 30116
rect 24136 30104 24164 30144
rect 24489 30141 24501 30144
rect 24535 30141 24547 30175
rect 24489 30135 24547 30141
rect 24673 30175 24731 30181
rect 24673 30141 24685 30175
rect 24719 30141 24731 30175
rect 24673 30135 24731 30141
rect 24949 30175 25007 30181
rect 24949 30141 24961 30175
rect 24995 30172 25007 30175
rect 24995 30144 25268 30172
rect 24995 30141 25007 30144
rect 24949 30135 25007 30141
rect 23532 30076 24164 30104
rect 23532 30064 23538 30076
rect 24394 30064 24400 30116
rect 24452 30064 24458 30116
rect 24688 30104 24716 30135
rect 24504 30076 24716 30104
rect 24504 30048 24532 30076
rect 25240 30048 25268 30144
rect 22848 30008 23428 30036
rect 22741 29999 22799 30005
rect 23658 29996 23664 30048
rect 23716 30036 23722 30048
rect 23845 30039 23903 30045
rect 23845 30036 23857 30039
rect 23716 30008 23857 30036
rect 23716 29996 23722 30008
rect 23845 30005 23857 30008
rect 23891 30005 23903 30039
rect 23845 29999 23903 30005
rect 23934 29996 23940 30048
rect 23992 30036 23998 30048
rect 24121 30039 24179 30045
rect 24121 30036 24133 30039
rect 23992 30008 24133 30036
rect 23992 29996 23998 30008
rect 24121 30005 24133 30008
rect 24167 30005 24179 30039
rect 24121 29999 24179 30005
rect 24210 29996 24216 30048
rect 24268 29996 24274 30048
rect 24486 29996 24492 30048
rect 24544 29996 24550 30048
rect 24854 29996 24860 30048
rect 24912 29996 24918 30048
rect 25222 29996 25228 30048
rect 25280 29996 25286 30048
rect 552 29946 27576 29968
rect 552 29894 7114 29946
rect 7166 29894 7178 29946
rect 7230 29894 7242 29946
rect 7294 29894 7306 29946
rect 7358 29894 7370 29946
rect 7422 29894 13830 29946
rect 13882 29894 13894 29946
rect 13946 29894 13958 29946
rect 14010 29894 14022 29946
rect 14074 29894 14086 29946
rect 14138 29894 20546 29946
rect 20598 29894 20610 29946
rect 20662 29894 20674 29946
rect 20726 29894 20738 29946
rect 20790 29894 20802 29946
rect 20854 29894 27262 29946
rect 27314 29894 27326 29946
rect 27378 29894 27390 29946
rect 27442 29894 27454 29946
rect 27506 29894 27518 29946
rect 27570 29894 27576 29946
rect 552 29872 27576 29894
rect 3510 29792 3516 29844
rect 3568 29832 3574 29844
rect 4065 29835 4123 29841
rect 4065 29832 4077 29835
rect 3568 29804 4077 29832
rect 3568 29792 3574 29804
rect 4065 29801 4077 29804
rect 4111 29801 4123 29835
rect 5810 29832 5816 29844
rect 4065 29795 4123 29801
rect 4724 29804 5816 29832
rect 3881 29767 3939 29773
rect 3881 29733 3893 29767
rect 3927 29764 3939 29767
rect 4154 29764 4160 29776
rect 3927 29736 4160 29764
rect 3927 29733 3939 29736
rect 3881 29727 3939 29733
rect 4154 29724 4160 29736
rect 4212 29724 4218 29776
rect 4525 29767 4583 29773
rect 4525 29764 4537 29767
rect 4264 29736 4537 29764
rect 1949 29699 2007 29705
rect 1949 29696 1961 29699
rect 1872 29668 1961 29696
rect 1872 29640 1900 29668
rect 1949 29665 1961 29668
rect 1995 29665 2007 29699
rect 1949 29659 2007 29665
rect 2038 29656 2044 29708
rect 2096 29696 2102 29708
rect 2205 29699 2263 29705
rect 2205 29696 2217 29699
rect 2096 29668 2217 29696
rect 2096 29656 2102 29668
rect 2205 29665 2217 29668
rect 2251 29665 2263 29699
rect 2205 29659 2263 29665
rect 3513 29699 3571 29705
rect 3513 29665 3525 29699
rect 3559 29696 3571 29699
rect 3602 29696 3608 29708
rect 3559 29668 3608 29696
rect 3559 29665 3571 29668
rect 3513 29659 3571 29665
rect 3602 29656 3608 29668
rect 3660 29696 3666 29708
rect 4264 29705 4292 29736
rect 4525 29733 4537 29736
rect 4571 29733 4583 29767
rect 4525 29727 4583 29733
rect 4724 29705 4752 29804
rect 5810 29792 5816 29804
rect 5868 29792 5874 29844
rect 5902 29792 5908 29844
rect 5960 29832 5966 29844
rect 6181 29835 6239 29841
rect 6181 29832 6193 29835
rect 5960 29804 6193 29832
rect 5960 29792 5966 29804
rect 6181 29801 6193 29804
rect 6227 29801 6239 29835
rect 6181 29795 6239 29801
rect 7009 29835 7067 29841
rect 7009 29801 7021 29835
rect 7055 29832 7067 29835
rect 7193 29835 7251 29841
rect 7055 29804 7144 29832
rect 7055 29801 7067 29804
rect 7009 29795 7067 29801
rect 6730 29764 6736 29776
rect 5184 29736 6736 29764
rect 5184 29705 5212 29736
rect 6730 29724 6736 29736
rect 6788 29724 6794 29776
rect 7116 29708 7144 29804
rect 7193 29801 7205 29835
rect 7239 29801 7251 29835
rect 7193 29795 7251 29801
rect 7208 29764 7236 29795
rect 7466 29792 7472 29844
rect 7524 29832 7530 29844
rect 7926 29832 7932 29844
rect 7524 29804 7932 29832
rect 7524 29792 7530 29804
rect 7926 29792 7932 29804
rect 7984 29832 7990 29844
rect 11790 29832 11796 29844
rect 7984 29804 8156 29832
rect 7984 29792 7990 29804
rect 7834 29764 7840 29776
rect 7208 29736 7840 29764
rect 7834 29724 7840 29736
rect 7892 29724 7898 29776
rect 4249 29699 4307 29705
rect 4249 29696 4261 29699
rect 3660 29668 4261 29696
rect 3660 29656 3666 29668
rect 4249 29665 4261 29668
rect 4295 29665 4307 29699
rect 4249 29659 4307 29665
rect 4433 29699 4491 29705
rect 4433 29665 4445 29699
rect 4479 29696 4491 29699
rect 4709 29699 4767 29705
rect 4709 29696 4721 29699
rect 4479 29668 4721 29696
rect 4479 29665 4491 29668
rect 4433 29659 4491 29665
rect 4709 29665 4721 29668
rect 4755 29665 4767 29699
rect 4709 29659 4767 29665
rect 5169 29699 5227 29705
rect 5169 29665 5181 29699
rect 5215 29665 5227 29699
rect 5997 29699 6055 29705
rect 5997 29696 6009 29699
rect 5169 29659 5227 29665
rect 5552 29668 6009 29696
rect 1854 29588 1860 29640
rect 1912 29588 1918 29640
rect 4341 29631 4399 29637
rect 4341 29597 4353 29631
rect 4387 29628 4399 29631
rect 5074 29628 5080 29640
rect 4387 29600 5080 29628
rect 4387 29597 4399 29600
rect 4341 29591 4399 29597
rect 5074 29588 5080 29600
rect 5132 29588 5138 29640
rect 5552 29569 5580 29668
rect 5997 29665 6009 29668
rect 6043 29665 6055 29699
rect 5997 29659 6055 29665
rect 6825 29699 6883 29705
rect 6825 29665 6837 29699
rect 6871 29665 6883 29699
rect 6825 29659 6883 29665
rect 5813 29631 5871 29637
rect 5813 29628 5825 29631
rect 5644 29600 5825 29628
rect 5537 29563 5595 29569
rect 3804 29532 4384 29560
rect 3329 29495 3387 29501
rect 3329 29461 3341 29495
rect 3375 29492 3387 29495
rect 3804 29492 3832 29532
rect 4356 29504 4384 29532
rect 4816 29532 5488 29560
rect 4816 29504 4844 29532
rect 3375 29464 3832 29492
rect 3881 29495 3939 29501
rect 3375 29461 3387 29464
rect 3329 29455 3387 29461
rect 3881 29461 3893 29495
rect 3927 29492 3939 29495
rect 4246 29492 4252 29504
rect 3927 29464 4252 29492
rect 3927 29461 3939 29464
rect 3881 29455 3939 29461
rect 4246 29452 4252 29464
rect 4304 29452 4310 29504
rect 4338 29452 4344 29504
rect 4396 29452 4402 29504
rect 4798 29452 4804 29504
rect 4856 29452 4862 29504
rect 4890 29452 4896 29504
rect 4948 29452 4954 29504
rect 5460 29492 5488 29532
rect 5537 29529 5549 29563
rect 5583 29529 5595 29563
rect 5537 29523 5595 29529
rect 5644 29492 5672 29600
rect 5813 29597 5825 29600
rect 5859 29597 5871 29631
rect 5813 29591 5871 29597
rect 6362 29588 6368 29640
rect 6420 29588 6426 29640
rect 6840 29628 6868 29659
rect 6914 29656 6920 29708
rect 6972 29656 6978 29708
rect 7098 29656 7104 29708
rect 7156 29656 7162 29708
rect 7742 29705 7748 29708
rect 7285 29699 7343 29705
rect 7285 29665 7297 29699
rect 7331 29696 7343 29699
rect 7331 29668 7696 29696
rect 7331 29665 7343 29668
rect 7285 29659 7343 29665
rect 7668 29640 7696 29668
rect 7736 29659 7748 29705
rect 7800 29696 7806 29708
rect 8128 29705 8156 29804
rect 9692 29804 11796 29832
rect 9582 29764 9588 29776
rect 8680 29736 9588 29764
rect 8113 29699 8171 29705
rect 7800 29668 7836 29696
rect 7742 29656 7748 29659
rect 7800 29656 7806 29668
rect 8113 29665 8125 29699
rect 8159 29665 8171 29699
rect 8113 29659 8171 29665
rect 8294 29656 8300 29708
rect 8352 29696 8358 29708
rect 8680 29705 8708 29736
rect 9582 29724 9588 29736
rect 9640 29724 9646 29776
rect 8573 29699 8631 29705
rect 8573 29696 8585 29699
rect 8352 29668 8585 29696
rect 8352 29656 8358 29668
rect 8573 29665 8585 29668
rect 8619 29665 8631 29699
rect 8573 29659 8631 29665
rect 8665 29699 8723 29705
rect 8665 29665 8677 29699
rect 8711 29665 8723 29699
rect 8665 29659 8723 29665
rect 8754 29656 8760 29708
rect 8812 29656 8818 29708
rect 9692 29705 9720 29804
rect 11790 29792 11796 29804
rect 11848 29832 11854 29844
rect 12345 29835 12403 29841
rect 12345 29832 12357 29835
rect 11848 29804 12357 29832
rect 11848 29792 11854 29804
rect 12345 29801 12357 29804
rect 12391 29801 12403 29835
rect 12345 29795 12403 29801
rect 12710 29792 12716 29844
rect 12768 29792 12774 29844
rect 12986 29832 12992 29844
rect 12912 29804 12992 29832
rect 9858 29764 9864 29776
rect 9784 29736 9864 29764
rect 9677 29699 9735 29705
rect 9677 29665 9689 29699
rect 9723 29665 9735 29699
rect 9677 29659 9735 29665
rect 7006 29628 7012 29640
rect 6840 29600 7012 29628
rect 7006 29588 7012 29600
rect 7064 29588 7070 29640
rect 7190 29588 7196 29640
rect 7248 29588 7254 29640
rect 7561 29631 7619 29637
rect 7561 29628 7573 29631
rect 7300 29600 7573 29628
rect 6380 29560 6408 29588
rect 7300 29560 7328 29600
rect 7561 29597 7573 29600
rect 7607 29597 7619 29631
rect 7561 29591 7619 29597
rect 7650 29588 7656 29640
rect 7708 29588 7714 29640
rect 9585 29631 9643 29637
rect 9585 29628 9597 29631
rect 7852 29600 9597 29628
rect 6380 29532 7328 29560
rect 7377 29563 7435 29569
rect 7377 29529 7389 29563
rect 7423 29529 7435 29563
rect 7377 29523 7435 29529
rect 5460 29464 5672 29492
rect 7098 29452 7104 29504
rect 7156 29492 7162 29504
rect 7392 29492 7420 29523
rect 7742 29520 7748 29572
rect 7800 29560 7806 29572
rect 7852 29560 7880 29600
rect 9585 29597 9597 29600
rect 9631 29597 9643 29631
rect 9585 29591 9643 29597
rect 9784 29560 9812 29736
rect 9858 29724 9864 29736
rect 9916 29764 9922 29776
rect 11210 29767 11268 29773
rect 11210 29764 11222 29767
rect 9916 29736 10456 29764
rect 9916 29724 9922 29736
rect 10045 29699 10103 29705
rect 10045 29665 10057 29699
rect 10091 29665 10103 29699
rect 10045 29659 10103 29665
rect 7800 29532 7880 29560
rect 8772 29532 9812 29560
rect 7800 29520 7806 29532
rect 8772 29504 8800 29532
rect 7558 29492 7564 29504
rect 7156 29464 7564 29492
rect 7156 29452 7162 29464
rect 7558 29452 7564 29464
rect 7616 29452 7622 29504
rect 8754 29452 8760 29504
rect 8812 29452 8818 29504
rect 9398 29452 9404 29504
rect 9456 29452 9462 29504
rect 10060 29492 10088 29659
rect 10226 29656 10232 29708
rect 10284 29656 10290 29708
rect 10318 29656 10324 29708
rect 10376 29656 10382 29708
rect 10428 29705 10456 29736
rect 10612 29736 11222 29764
rect 10413 29699 10471 29705
rect 10413 29665 10425 29699
rect 10459 29665 10471 29699
rect 10413 29659 10471 29665
rect 10612 29569 10640 29736
rect 11210 29733 11222 29736
rect 11256 29733 11268 29767
rect 11210 29727 11268 29733
rect 12434 29724 12440 29776
rect 12492 29724 12498 29776
rect 12912 29773 12940 29804
rect 12986 29792 12992 29804
rect 13044 29792 13050 29844
rect 14274 29832 14280 29844
rect 14016 29804 14280 29832
rect 14016 29773 14044 29804
rect 14274 29792 14280 29804
rect 14332 29792 14338 29844
rect 14369 29835 14427 29841
rect 14369 29801 14381 29835
rect 14415 29832 14427 29835
rect 15010 29832 15016 29844
rect 14415 29804 15016 29832
rect 14415 29801 14427 29804
rect 14369 29795 14427 29801
rect 15010 29792 15016 29804
rect 15068 29832 15074 29844
rect 15121 29835 15179 29841
rect 15121 29832 15133 29835
rect 15068 29804 15133 29832
rect 15068 29792 15074 29804
rect 15121 29801 15133 29804
rect 15167 29801 15179 29835
rect 15121 29795 15179 29801
rect 15286 29792 15292 29844
rect 15344 29792 15350 29844
rect 16114 29792 16120 29844
rect 16172 29832 16178 29844
rect 16301 29835 16359 29841
rect 16301 29832 16313 29835
rect 16172 29804 16313 29832
rect 16172 29792 16178 29804
rect 16301 29801 16313 29804
rect 16347 29832 16359 29835
rect 16347 29804 16620 29832
rect 16347 29801 16359 29804
rect 16301 29795 16359 29801
rect 12897 29767 12955 29773
rect 12897 29733 12909 29767
rect 12943 29733 12955 29767
rect 12897 29727 12955 29733
rect 14001 29767 14059 29773
rect 14001 29733 14013 29767
rect 14047 29733 14059 29767
rect 14001 29727 14059 29733
rect 14458 29724 14464 29776
rect 14516 29773 14522 29776
rect 14516 29767 14537 29773
rect 14525 29733 14537 29767
rect 14516 29727 14537 29733
rect 14921 29767 14979 29773
rect 14921 29733 14933 29767
rect 14967 29764 14979 29767
rect 15378 29764 15384 29776
rect 14967 29736 15384 29764
rect 14967 29733 14979 29736
rect 14921 29727 14979 29733
rect 14516 29724 14522 29727
rect 15378 29724 15384 29736
rect 15436 29724 15442 29776
rect 15562 29724 15568 29776
rect 15620 29773 15626 29776
rect 15620 29767 15669 29773
rect 15620 29733 15623 29767
rect 15657 29733 15669 29767
rect 15781 29767 15839 29773
rect 15781 29764 15793 29767
rect 15620 29727 15669 29733
rect 15764 29733 15793 29764
rect 15827 29764 15839 29767
rect 16206 29764 16212 29776
rect 15827 29736 16212 29764
rect 15827 29733 15839 29736
rect 15764 29727 15839 29733
rect 15620 29724 15626 29727
rect 13078 29656 13084 29708
rect 13136 29696 13142 29708
rect 13854 29699 13912 29705
rect 13854 29696 13866 29699
rect 13136 29668 13866 29696
rect 13136 29656 13142 29668
rect 13854 29665 13866 29668
rect 13900 29665 13912 29699
rect 13854 29659 13912 29665
rect 14185 29699 14243 29705
rect 14185 29665 14197 29699
rect 14231 29665 14243 29699
rect 14185 29659 14243 29665
rect 14369 29699 14427 29705
rect 14369 29665 14381 29699
rect 14415 29694 14427 29699
rect 14645 29699 14703 29705
rect 14645 29696 14657 29699
rect 14568 29694 14657 29696
rect 14415 29668 14657 29694
rect 14415 29666 14596 29668
rect 14415 29665 14427 29666
rect 14369 29659 14427 29665
rect 14645 29665 14657 29668
rect 14691 29665 14703 29699
rect 14645 29659 14703 29665
rect 10962 29588 10968 29640
rect 11020 29588 11026 29640
rect 12158 29588 12164 29640
rect 12216 29628 12222 29640
rect 12434 29628 12440 29640
rect 12216 29600 12440 29628
rect 12216 29588 12222 29600
rect 12434 29588 12440 29600
rect 12492 29588 12498 29640
rect 12805 29631 12863 29637
rect 12805 29597 12817 29631
rect 12851 29628 12863 29631
rect 13538 29628 13544 29640
rect 12851 29600 13544 29628
rect 12851 29597 12863 29600
rect 12805 29591 12863 29597
rect 13538 29588 13544 29600
rect 13596 29588 13602 29640
rect 13633 29631 13691 29637
rect 13633 29597 13645 29631
rect 13679 29597 13691 29631
rect 13633 29591 13691 29597
rect 10597 29563 10655 29569
rect 10597 29529 10609 29563
rect 10643 29529 10655 29563
rect 13354 29560 13360 29572
rect 10597 29523 10655 29529
rect 13004 29532 13360 29560
rect 13004 29504 13032 29532
rect 13354 29520 13360 29532
rect 13412 29520 13418 29572
rect 13446 29520 13452 29572
rect 13504 29560 13510 29572
rect 13648 29560 13676 29591
rect 13504 29532 13676 29560
rect 14200 29560 14228 29659
rect 14660 29628 14688 29659
rect 15562 29628 15568 29640
rect 14660 29600 15568 29628
rect 15562 29588 15568 29600
rect 15620 29588 15626 29640
rect 15764 29628 15792 29727
rect 16206 29724 16212 29736
rect 16264 29724 16270 29776
rect 16482 29724 16488 29776
rect 16540 29724 16546 29776
rect 16592 29764 16620 29804
rect 16758 29792 16764 29844
rect 16816 29792 16822 29844
rect 17034 29832 17040 29844
rect 16868 29804 17040 29832
rect 16868 29764 16896 29804
rect 17034 29792 17040 29804
rect 17092 29792 17098 29844
rect 20622 29792 20628 29844
rect 20680 29832 20686 29844
rect 22925 29835 22983 29841
rect 22925 29832 22937 29835
rect 20680 29804 22937 29832
rect 20680 29792 20686 29804
rect 22925 29801 22937 29804
rect 22971 29832 22983 29835
rect 22971 29804 23428 29832
rect 22971 29801 22983 29804
rect 22925 29795 22983 29801
rect 16592 29736 16896 29764
rect 16942 29724 16948 29776
rect 17000 29724 17006 29776
rect 18230 29724 18236 29776
rect 18288 29764 18294 29776
rect 18610 29767 18668 29773
rect 18610 29764 18622 29767
rect 18288 29736 18622 29764
rect 18288 29724 18294 29736
rect 18610 29733 18622 29736
rect 18656 29733 18668 29767
rect 18610 29727 18668 29733
rect 18966 29724 18972 29776
rect 19024 29764 19030 29776
rect 21542 29764 21548 29776
rect 19024 29736 21548 29764
rect 19024 29724 19030 29736
rect 21542 29724 21548 29736
rect 21600 29724 21606 29776
rect 23400 29764 23428 29804
rect 23842 29792 23848 29844
rect 23900 29832 23906 29844
rect 24305 29835 24363 29841
rect 23900 29804 24256 29832
rect 23900 29792 23906 29804
rect 23400 29736 23704 29764
rect 16393 29699 16451 29705
rect 16393 29696 16405 29699
rect 15672 29600 15792 29628
rect 15856 29668 16405 29696
rect 14458 29560 14464 29572
rect 14200 29532 14464 29560
rect 13504 29520 13510 29532
rect 14458 29520 14464 29532
rect 14516 29560 14522 29572
rect 14642 29560 14648 29572
rect 14516 29532 14648 29560
rect 14516 29520 14522 29532
rect 14642 29520 14648 29532
rect 14700 29560 14706 29572
rect 15672 29560 15700 29600
rect 14700 29532 15700 29560
rect 14700 29520 14706 29532
rect 11238 29492 11244 29504
rect 10060 29464 11244 29492
rect 11238 29452 11244 29464
rect 11296 29452 11302 29504
rect 12986 29452 12992 29504
rect 13044 29452 13050 29504
rect 13078 29452 13084 29504
rect 13136 29452 13142 29504
rect 13630 29452 13636 29504
rect 13688 29492 13694 29504
rect 13725 29495 13783 29501
rect 13725 29492 13737 29495
rect 13688 29464 13737 29492
rect 13688 29452 13694 29464
rect 13725 29461 13737 29464
rect 13771 29461 13783 29495
rect 13725 29455 13783 29461
rect 14829 29495 14887 29501
rect 14829 29461 14841 29495
rect 14875 29492 14887 29495
rect 15105 29495 15163 29501
rect 15105 29492 15117 29495
rect 14875 29464 15117 29492
rect 14875 29461 14887 29464
rect 14829 29455 14887 29461
rect 15105 29461 15117 29464
rect 15151 29461 15163 29495
rect 15105 29455 15163 29461
rect 15654 29452 15660 29504
rect 15712 29492 15718 29504
rect 15749 29495 15807 29501
rect 15749 29492 15761 29495
rect 15712 29464 15761 29492
rect 15712 29452 15718 29464
rect 15749 29461 15761 29464
rect 15795 29492 15807 29495
rect 15856 29492 15884 29668
rect 16393 29665 16405 29668
rect 16439 29665 16451 29699
rect 16393 29659 16451 29665
rect 17310 29656 17316 29708
rect 17368 29696 17374 29708
rect 18877 29699 18935 29705
rect 17368 29668 18828 29696
rect 17368 29656 17374 29668
rect 18800 29628 18828 29668
rect 18877 29665 18889 29699
rect 18923 29696 18935 29699
rect 19429 29699 19487 29705
rect 19429 29696 19441 29699
rect 18923 29668 19441 29696
rect 18923 29665 18935 29668
rect 18877 29659 18935 29665
rect 19429 29665 19441 29668
rect 19475 29696 19487 29699
rect 19518 29696 19524 29708
rect 19475 29668 19524 29696
rect 19475 29665 19487 29668
rect 19429 29659 19487 29665
rect 19518 29656 19524 29668
rect 19576 29656 19582 29708
rect 19702 29705 19708 29708
rect 19696 29659 19708 29705
rect 19702 29656 19708 29659
rect 19760 29656 19766 29708
rect 22393 29699 22451 29705
rect 22393 29665 22405 29699
rect 22439 29696 22451 29699
rect 22922 29696 22928 29708
rect 22439 29668 22784 29696
rect 22883 29668 22928 29696
rect 22439 29665 22451 29668
rect 22393 29659 22451 29665
rect 19242 29628 19248 29640
rect 16132 29600 17540 29628
rect 18800 29600 19248 29628
rect 16132 29572 16160 29600
rect 16114 29520 16120 29572
rect 16172 29520 16178 29572
rect 17034 29520 17040 29572
rect 17092 29560 17098 29572
rect 17313 29563 17371 29569
rect 17313 29560 17325 29563
rect 17092 29532 17325 29560
rect 17092 29520 17098 29532
rect 17313 29529 17325 29532
rect 17359 29529 17371 29563
rect 17313 29523 17371 29529
rect 15795 29464 15884 29492
rect 15795 29461 15807 29464
rect 15749 29455 15807 29461
rect 15930 29452 15936 29504
rect 15988 29452 15994 29504
rect 16666 29452 16672 29504
rect 16724 29452 16730 29504
rect 16758 29452 16764 29504
rect 16816 29492 16822 29504
rect 17512 29501 17540 29600
rect 19242 29588 19248 29600
rect 19300 29588 19306 29640
rect 22646 29588 22652 29640
rect 22704 29588 22710 29640
rect 22756 29628 22784 29668
rect 22922 29656 22928 29668
rect 22980 29656 22986 29708
rect 23382 29656 23388 29708
rect 23440 29656 23446 29708
rect 23676 29705 23704 29736
rect 23860 29705 23888 29792
rect 23477 29699 23535 29705
rect 23477 29665 23489 29699
rect 23523 29665 23535 29699
rect 23477 29659 23535 29665
rect 23661 29699 23719 29705
rect 23661 29665 23673 29699
rect 23707 29665 23719 29699
rect 23661 29659 23719 29665
rect 23845 29699 23903 29705
rect 23845 29665 23857 29699
rect 23891 29665 23903 29699
rect 23845 29659 23903 29665
rect 24012 29699 24070 29705
rect 24012 29665 24024 29699
rect 24058 29696 24070 29699
rect 24228 29696 24256 29804
rect 24305 29801 24317 29835
rect 24351 29832 24363 29835
rect 24394 29832 24400 29844
rect 24351 29804 24400 29832
rect 24351 29801 24363 29804
rect 24305 29795 24363 29801
rect 24394 29792 24400 29804
rect 24452 29792 24458 29844
rect 24489 29835 24547 29841
rect 24489 29801 24501 29835
rect 24535 29832 24547 29835
rect 24535 29804 24716 29832
rect 24535 29801 24547 29804
rect 24489 29795 24547 29801
rect 24688 29776 24716 29804
rect 24854 29792 24860 29844
rect 24912 29792 24918 29844
rect 24670 29724 24676 29776
rect 24728 29724 24734 29776
rect 24430 29699 24488 29705
rect 24430 29696 24442 29699
rect 24058 29694 24072 29696
rect 24058 29666 24164 29694
rect 24228 29668 24442 29696
rect 24058 29665 24070 29666
rect 24012 29659 24070 29665
rect 23106 29628 23112 29640
rect 22756 29600 23112 29628
rect 23106 29588 23112 29600
rect 23164 29588 23170 29640
rect 22741 29563 22799 29569
rect 22741 29529 22753 29563
rect 22787 29560 22799 29563
rect 23492 29560 23520 29659
rect 23750 29588 23756 29640
rect 23808 29588 23814 29640
rect 24136 29628 24164 29666
rect 24430 29665 24442 29668
rect 24476 29665 24488 29699
rect 24430 29659 24488 29665
rect 24688 29628 24716 29724
rect 24872 29705 24900 29792
rect 24857 29699 24915 29705
rect 24857 29665 24869 29699
rect 24903 29665 24915 29699
rect 24857 29659 24915 29665
rect 24949 29699 25007 29705
rect 24949 29665 24961 29699
rect 24995 29696 25007 29699
rect 25501 29699 25559 29705
rect 25501 29696 25513 29699
rect 24995 29668 25513 29696
rect 24995 29665 25007 29668
rect 24949 29659 25007 29665
rect 25501 29665 25513 29668
rect 25547 29696 25559 29699
rect 25958 29696 25964 29708
rect 25547 29668 25964 29696
rect 25547 29665 25559 29668
rect 25501 29659 25559 29665
rect 25958 29656 25964 29668
rect 26016 29656 26022 29708
rect 24136 29600 24716 29628
rect 24578 29560 24584 29572
rect 22787 29532 23428 29560
rect 23492 29532 24584 29560
rect 22787 29529 22799 29532
rect 22741 29523 22799 29529
rect 16945 29495 17003 29501
rect 16945 29492 16957 29495
rect 16816 29464 16957 29492
rect 16816 29452 16822 29464
rect 16945 29461 16957 29464
rect 16991 29461 17003 29495
rect 16945 29455 17003 29461
rect 17497 29495 17555 29501
rect 17497 29461 17509 29495
rect 17543 29492 17555 29495
rect 17586 29492 17592 29504
rect 17543 29464 17592 29492
rect 17543 29461 17555 29464
rect 17497 29455 17555 29461
rect 17586 29452 17592 29464
rect 17644 29452 17650 29504
rect 18138 29452 18144 29504
rect 18196 29492 18202 29504
rect 19150 29492 19156 29504
rect 18196 29464 19156 29492
rect 18196 29452 18202 29464
rect 19150 29452 19156 29464
rect 19208 29492 19214 29504
rect 19610 29492 19616 29504
rect 19208 29464 19616 29492
rect 19208 29452 19214 29464
rect 19610 29452 19616 29464
rect 19668 29492 19674 29504
rect 20070 29492 20076 29504
rect 19668 29464 20076 29492
rect 19668 29452 19674 29464
rect 20070 29452 20076 29464
rect 20128 29452 20134 29504
rect 20622 29452 20628 29504
rect 20680 29492 20686 29504
rect 20809 29495 20867 29501
rect 20809 29492 20821 29495
rect 20680 29464 20821 29492
rect 20680 29452 20686 29464
rect 20809 29461 20821 29464
rect 20855 29461 20867 29495
rect 20809 29455 20867 29461
rect 21269 29495 21327 29501
rect 21269 29461 21281 29495
rect 21315 29492 21327 29495
rect 21726 29492 21732 29504
rect 21315 29464 21732 29492
rect 21315 29461 21327 29464
rect 21269 29455 21327 29461
rect 21726 29452 21732 29464
rect 21784 29492 21790 29504
rect 22830 29492 22836 29504
rect 21784 29464 22836 29492
rect 21784 29452 21790 29464
rect 22830 29452 22836 29464
rect 22888 29452 22894 29504
rect 23290 29452 23296 29504
rect 23348 29452 23354 29504
rect 23400 29492 23428 29532
rect 24578 29520 24584 29532
rect 24636 29560 24642 29572
rect 25041 29563 25099 29569
rect 25041 29560 25053 29563
rect 24636 29532 25053 29560
rect 24636 29520 24642 29532
rect 25041 29529 25053 29532
rect 25087 29529 25099 29563
rect 25041 29523 25099 29529
rect 23750 29492 23756 29504
rect 23400 29464 23756 29492
rect 23750 29452 23756 29464
rect 23808 29452 23814 29504
rect 24210 29452 24216 29504
rect 24268 29452 24274 29504
rect 25222 29452 25228 29504
rect 25280 29452 25286 29504
rect 552 29402 27416 29424
rect 552 29350 3756 29402
rect 3808 29350 3820 29402
rect 3872 29350 3884 29402
rect 3936 29350 3948 29402
rect 4000 29350 4012 29402
rect 4064 29350 10472 29402
rect 10524 29350 10536 29402
rect 10588 29350 10600 29402
rect 10652 29350 10664 29402
rect 10716 29350 10728 29402
rect 10780 29350 17188 29402
rect 17240 29350 17252 29402
rect 17304 29350 17316 29402
rect 17368 29350 17380 29402
rect 17432 29350 17444 29402
rect 17496 29350 23904 29402
rect 23956 29350 23968 29402
rect 24020 29350 24032 29402
rect 24084 29350 24096 29402
rect 24148 29350 24160 29402
rect 24212 29350 27416 29402
rect 552 29328 27416 29350
rect 3602 29248 3608 29300
rect 3660 29288 3666 29300
rect 3697 29291 3755 29297
rect 3697 29288 3709 29291
rect 3660 29260 3709 29288
rect 3660 29248 3666 29260
rect 3697 29257 3709 29260
rect 3743 29257 3755 29291
rect 3697 29251 3755 29257
rect 4154 29248 4160 29300
rect 4212 29288 4218 29300
rect 4525 29291 4583 29297
rect 4525 29288 4537 29291
rect 4212 29260 4537 29288
rect 4212 29248 4218 29260
rect 4525 29257 4537 29260
rect 4571 29257 4583 29291
rect 4525 29251 4583 29257
rect 4890 29248 4896 29300
rect 4948 29288 4954 29300
rect 4985 29291 5043 29297
rect 4985 29288 4997 29291
rect 4948 29260 4997 29288
rect 4948 29248 4954 29260
rect 4985 29257 4997 29260
rect 5031 29257 5043 29291
rect 4985 29251 5043 29257
rect 5074 29248 5080 29300
rect 5132 29248 5138 29300
rect 6454 29248 6460 29300
rect 6512 29248 6518 29300
rect 6914 29248 6920 29300
rect 6972 29248 6978 29300
rect 7190 29248 7196 29300
rect 7248 29248 7254 29300
rect 7469 29291 7527 29297
rect 7469 29257 7481 29291
rect 7515 29288 7527 29291
rect 7650 29288 7656 29300
rect 7515 29260 7656 29288
rect 7515 29257 7527 29260
rect 7469 29251 7527 29257
rect 7650 29248 7656 29260
rect 7708 29248 7714 29300
rect 8113 29291 8171 29297
rect 8113 29257 8125 29291
rect 8159 29288 8171 29291
rect 8478 29288 8484 29300
rect 8159 29260 8484 29288
rect 8159 29257 8171 29260
rect 8113 29251 8171 29257
rect 8478 29248 8484 29260
rect 8536 29248 8542 29300
rect 8662 29248 8668 29300
rect 8720 29248 8726 29300
rect 9398 29248 9404 29300
rect 9456 29248 9462 29300
rect 9490 29248 9496 29300
rect 9548 29288 9554 29300
rect 9674 29288 9680 29300
rect 9548 29260 9680 29288
rect 9548 29248 9554 29260
rect 9674 29248 9680 29260
rect 9732 29288 9738 29300
rect 10226 29288 10232 29300
rect 9732 29260 10232 29288
rect 9732 29248 9738 29260
rect 10226 29248 10232 29260
rect 10284 29248 10290 29300
rect 10318 29248 10324 29300
rect 10376 29288 10382 29300
rect 11146 29288 11152 29300
rect 10376 29260 11152 29288
rect 10376 29248 10382 29260
rect 11146 29248 11152 29260
rect 11204 29248 11210 29300
rect 13262 29248 13268 29300
rect 13320 29248 13326 29300
rect 13538 29248 13544 29300
rect 13596 29248 13602 29300
rect 13722 29248 13728 29300
rect 13780 29288 13786 29300
rect 13817 29291 13875 29297
rect 13817 29288 13829 29291
rect 13780 29260 13829 29288
rect 13780 29248 13786 29260
rect 13817 29257 13829 29260
rect 13863 29257 13875 29291
rect 16574 29288 16580 29300
rect 13817 29251 13875 29257
rect 15580 29260 16580 29288
rect 4249 29223 4307 29229
rect 4249 29220 4261 29223
rect 3896 29192 4261 29220
rect 3050 29044 3056 29096
rect 3108 29084 3114 29096
rect 3896 29093 3924 29192
rect 4249 29189 4261 29192
rect 4295 29220 4307 29223
rect 4295 29192 4476 29220
rect 4295 29189 4307 29192
rect 4249 29183 4307 29189
rect 3697 29087 3755 29093
rect 3697 29084 3709 29087
rect 3108 29056 3709 29084
rect 3108 29044 3114 29056
rect 3697 29053 3709 29056
rect 3743 29053 3755 29087
rect 3697 29047 3755 29053
rect 3881 29087 3939 29093
rect 3881 29053 3893 29087
rect 3927 29053 3939 29087
rect 4333 29089 4391 29095
rect 4448 29093 4476 29192
rect 4333 29086 4345 29089
rect 3881 29047 3939 29053
rect 4232 29058 4345 29086
rect 3712 29016 3740 29047
rect 3970 29016 3976 29028
rect 3712 28988 3976 29016
rect 3970 28976 3976 28988
rect 4028 28976 4034 29028
rect 4232 29016 4260 29058
rect 4333 29055 4345 29058
rect 4379 29055 4391 29089
rect 4333 29049 4391 29055
rect 4433 29087 4491 29093
rect 4433 29053 4445 29087
rect 4479 29053 4491 29087
rect 4433 29047 4491 29053
rect 4614 29044 4620 29096
rect 4672 29044 4678 29096
rect 4232 28994 4292 29016
rect 4232 28988 4384 28994
rect 4264 28966 4384 28988
rect 4798 28976 4804 29028
rect 4856 28976 4862 29028
rect 5006 29019 5064 29025
rect 5006 28985 5018 29019
rect 5052 29016 5064 29019
rect 5092 29016 5120 29248
rect 5169 29223 5227 29229
rect 5169 29189 5181 29223
rect 5215 29189 5227 29223
rect 5169 29183 5227 29189
rect 5445 29223 5503 29229
rect 5445 29189 5457 29223
rect 5491 29220 5503 29223
rect 5902 29220 5908 29232
rect 5491 29192 5908 29220
rect 5491 29189 5503 29192
rect 5445 29183 5503 29189
rect 5184 29084 5212 29183
rect 5902 29180 5908 29192
rect 5960 29180 5966 29232
rect 6932 29152 6960 29248
rect 7208 29220 7236 29248
rect 7208 29192 7604 29220
rect 6932 29124 7328 29152
rect 5261 29087 5319 29093
rect 5261 29084 5273 29087
rect 5184 29056 5273 29084
rect 5261 29053 5273 29056
rect 5307 29053 5319 29087
rect 5261 29047 5319 29053
rect 5442 29044 5448 29096
rect 5500 29084 5506 29096
rect 6362 29084 6368 29096
rect 5500 29056 6368 29084
rect 5500 29044 5506 29056
rect 6362 29044 6368 29056
rect 6420 29044 6426 29096
rect 6638 29044 6644 29096
rect 6696 29044 6702 29096
rect 7300 29093 7328 29124
rect 7576 29093 7604 29192
rect 8294 29180 8300 29232
rect 8352 29180 8358 29232
rect 8312 29152 8340 29180
rect 7852 29124 8340 29152
rect 7852 29093 7880 29124
rect 6733 29087 6791 29093
rect 6733 29053 6745 29087
rect 6779 29053 6791 29087
rect 6733 29047 6791 29053
rect 7193 29087 7251 29093
rect 7193 29053 7205 29087
rect 7239 29053 7251 29087
rect 7193 29047 7251 29053
rect 7285 29087 7343 29093
rect 7285 29053 7297 29087
rect 7331 29053 7343 29087
rect 7285 29047 7343 29053
rect 7561 29087 7619 29093
rect 7561 29053 7573 29087
rect 7607 29053 7619 29087
rect 7561 29047 7619 29053
rect 7837 29087 7895 29093
rect 7837 29053 7849 29087
rect 7883 29053 7895 29087
rect 7837 29047 7895 29053
rect 5460 29016 5488 29044
rect 5052 28988 5120 29016
rect 5184 28988 5488 29016
rect 6748 29016 6776 29047
rect 7208 29016 7236 29047
rect 7466 29016 7472 29028
rect 6748 28988 7144 29016
rect 7208 28988 7472 29016
rect 5052 28985 5064 28988
rect 5006 28979 5064 28985
rect 4356 28948 4384 28966
rect 5184 28948 5212 28988
rect 4356 28920 5212 28948
rect 7006 28908 7012 28960
rect 7064 28908 7070 28960
rect 7116 28948 7144 28988
rect 7466 28976 7472 28988
rect 7524 28976 7530 29028
rect 7576 29016 7604 29047
rect 7926 29044 7932 29096
rect 7984 29044 7990 29096
rect 8018 29044 8024 29096
rect 8076 29084 8082 29096
rect 8205 29087 8263 29093
rect 8205 29084 8217 29087
rect 8076 29056 8217 29084
rect 8076 29044 8082 29056
rect 8205 29053 8217 29056
rect 8251 29053 8263 29087
rect 8205 29047 8263 29053
rect 8754 29044 8760 29096
rect 8812 29084 8818 29096
rect 8849 29087 8907 29093
rect 8849 29084 8861 29087
rect 8812 29056 8861 29084
rect 8812 29044 8818 29056
rect 8849 29053 8861 29056
rect 8895 29053 8907 29087
rect 9217 29087 9275 29093
rect 8849 29047 8907 29053
rect 8956 29056 9168 29084
rect 8956 29028 8984 29056
rect 7650 29016 7656 29028
rect 7576 28988 7656 29016
rect 7650 28976 7656 28988
rect 7708 28976 7714 29028
rect 8386 28976 8392 29028
rect 8444 28976 8450 29028
rect 8938 28976 8944 29028
rect 8996 28976 9002 29028
rect 9033 29019 9091 29025
rect 9033 28985 9045 29019
rect 9079 28985 9091 29019
rect 9140 29016 9168 29056
rect 9217 29053 9229 29087
rect 9263 29084 9275 29087
rect 9416 29084 9444 29248
rect 12434 29220 12440 29232
rect 9263 29056 9444 29084
rect 10152 29192 12440 29220
rect 9263 29053 9275 29056
rect 9217 29047 9275 29053
rect 10152 29016 10180 29192
rect 12434 29180 12440 29192
rect 12492 29220 12498 29232
rect 12492 29192 12940 29220
rect 12492 29180 12498 29192
rect 11885 29087 11943 29093
rect 11885 29053 11897 29087
rect 11931 29084 11943 29087
rect 12253 29087 12311 29093
rect 11931 29056 12204 29084
rect 11931 29053 11943 29056
rect 11885 29047 11943 29053
rect 9140 28988 10180 29016
rect 11057 29019 11115 29025
rect 9033 28979 9091 28985
rect 11057 28985 11069 29019
rect 11103 29016 11115 29019
rect 11606 29016 11612 29028
rect 11103 28988 11612 29016
rect 11103 28985 11115 28988
rect 11057 28979 11115 28985
rect 7742 28948 7748 28960
rect 7116 28920 7748 28948
rect 7742 28908 7748 28920
rect 7800 28908 7806 28960
rect 8404 28948 8432 28976
rect 9048 28948 9076 28979
rect 11606 28976 11612 28988
rect 11664 28976 11670 29028
rect 11974 28976 11980 29028
rect 12032 28976 12038 29028
rect 12066 28976 12072 29028
rect 12124 28976 12130 29028
rect 12176 29016 12204 29056
rect 12253 29053 12265 29087
rect 12299 29084 12311 29087
rect 12345 29087 12403 29093
rect 12345 29084 12357 29087
rect 12299 29056 12357 29084
rect 12299 29053 12311 29056
rect 12253 29047 12311 29053
rect 12345 29053 12357 29056
rect 12391 29053 12403 29087
rect 12345 29047 12403 29053
rect 12176 28988 12434 29016
rect 9490 28948 9496 28960
rect 8404 28920 9496 28948
rect 9490 28908 9496 28920
rect 9548 28908 9554 28960
rect 9585 28951 9643 28957
rect 9585 28917 9597 28951
rect 9631 28948 9643 28951
rect 9674 28948 9680 28960
rect 9631 28920 9680 28948
rect 9631 28917 9643 28920
rect 9585 28911 9643 28917
rect 9674 28908 9680 28920
rect 9732 28908 9738 28960
rect 11698 28908 11704 28960
rect 11756 28908 11762 28960
rect 12406 28948 12434 28988
rect 12618 28948 12624 28960
rect 12406 28920 12624 28948
rect 12618 28908 12624 28920
rect 12676 28908 12682 28960
rect 12912 28948 12940 29192
rect 12989 29087 13047 29093
rect 12989 29053 13001 29087
rect 13035 29053 13047 29087
rect 13280 29084 13308 29248
rect 13556 29220 13584 29248
rect 15580 29220 15608 29260
rect 16574 29248 16580 29260
rect 16632 29248 16638 29300
rect 16942 29248 16948 29300
rect 17000 29248 17006 29300
rect 17126 29248 17132 29300
rect 17184 29248 17190 29300
rect 17313 29291 17371 29297
rect 17313 29257 17325 29291
rect 17359 29288 17371 29291
rect 18046 29288 18052 29300
rect 17359 29260 18052 29288
rect 17359 29257 17371 29260
rect 17313 29251 17371 29257
rect 18046 29248 18052 29260
rect 18104 29248 18110 29300
rect 19334 29288 19340 29300
rect 18340 29260 19340 29288
rect 16114 29220 16120 29232
rect 13556 29192 15608 29220
rect 15672 29192 16120 29220
rect 13354 29112 13360 29164
rect 13412 29152 13418 29164
rect 15010 29152 15016 29164
rect 13412 29124 13676 29152
rect 13412 29112 13418 29124
rect 13648 29093 13676 29124
rect 14936 29124 15016 29152
rect 13541 29087 13599 29093
rect 13541 29084 13553 29087
rect 13280 29056 13553 29084
rect 12989 29047 13047 29053
rect 13541 29053 13553 29056
rect 13587 29053 13599 29087
rect 13541 29047 13599 29053
rect 13633 29087 13691 29093
rect 13633 29053 13645 29087
rect 13679 29053 13691 29087
rect 13633 29047 13691 29053
rect 14001 29087 14059 29093
rect 14001 29053 14013 29087
rect 14047 29084 14059 29087
rect 14458 29084 14464 29096
rect 14047 29056 14464 29084
rect 14047 29053 14059 29056
rect 14001 29047 14059 29053
rect 13004 29016 13032 29047
rect 14458 29044 14464 29056
rect 14516 29044 14522 29096
rect 14936 29093 14964 29124
rect 15010 29112 15016 29124
rect 15068 29112 15074 29164
rect 14921 29087 14979 29093
rect 14921 29053 14933 29087
rect 14967 29053 14979 29087
rect 14921 29047 14979 29053
rect 15102 29044 15108 29096
rect 15160 29044 15166 29096
rect 15672 29093 15700 29192
rect 16114 29180 16120 29192
rect 16172 29180 16178 29232
rect 16666 29180 16672 29232
rect 16724 29220 16730 29232
rect 16761 29223 16819 29229
rect 16761 29220 16773 29223
rect 16724 29192 16773 29220
rect 16724 29180 16730 29192
rect 16761 29189 16773 29192
rect 16807 29189 16819 29223
rect 16761 29183 16819 29189
rect 16960 29152 16988 29248
rect 15856 29124 16988 29152
rect 15657 29087 15715 29093
rect 15657 29053 15669 29087
rect 15703 29053 15715 29087
rect 15657 29047 15715 29053
rect 15746 29044 15752 29096
rect 15804 29044 15810 29096
rect 15013 29019 15071 29025
rect 13004 28988 13584 29016
rect 13556 28960 13584 28988
rect 15013 28985 15025 29019
rect 15059 29016 15071 29019
rect 15856 29016 15884 29124
rect 17034 29044 17040 29096
rect 17092 29044 17098 29096
rect 17773 29087 17831 29093
rect 17773 29084 17785 29087
rect 17144 29056 17785 29084
rect 15059 28988 15884 29016
rect 15059 28985 15071 28988
rect 15013 28979 15071 28985
rect 15930 28976 15936 29028
rect 15988 29016 15994 29028
rect 17052 29016 17080 29044
rect 17144 29025 17172 29056
rect 17773 29053 17785 29056
rect 17819 29053 17831 29087
rect 17773 29047 17831 29053
rect 17957 29087 18015 29093
rect 17957 29053 17969 29087
rect 18003 29053 18015 29087
rect 17957 29047 18015 29053
rect 15988 28988 17080 29016
rect 15988 28976 15994 28988
rect 13446 28948 13452 28960
rect 12912 28920 13452 28948
rect 13446 28908 13452 28920
rect 13504 28908 13510 28960
rect 13538 28908 13544 28960
rect 13596 28908 13602 28960
rect 15562 28908 15568 28960
rect 15620 28908 15626 28960
rect 15838 28908 15844 28960
rect 15896 28908 15902 28960
rect 16390 28908 16396 28960
rect 16448 28948 16454 28960
rect 16758 28948 16764 28960
rect 16448 28920 16764 28948
rect 16448 28908 16454 28920
rect 16758 28908 16764 28920
rect 16816 28908 16822 28960
rect 17052 28948 17080 28988
rect 17129 29019 17187 29025
rect 17129 28985 17141 29019
rect 17175 28985 17187 29019
rect 17405 29019 17463 29025
rect 17405 29016 17417 29019
rect 17129 28979 17187 28985
rect 17236 28988 17417 29016
rect 17236 28948 17264 28988
rect 17405 28985 17417 28988
rect 17451 28985 17463 29019
rect 17405 28979 17463 28985
rect 17586 28976 17592 29028
rect 17644 28976 17650 29028
rect 17972 29016 18000 29047
rect 18138 29044 18144 29096
rect 18196 29044 18202 29096
rect 18340 29093 18368 29260
rect 19334 29248 19340 29260
rect 19392 29248 19398 29300
rect 19521 29291 19579 29297
rect 19521 29257 19533 29291
rect 19567 29288 19579 29291
rect 19702 29288 19708 29300
rect 19567 29260 19708 29288
rect 19567 29257 19579 29260
rect 19521 29251 19579 29257
rect 19702 29248 19708 29260
rect 19760 29248 19766 29300
rect 23014 29288 23020 29300
rect 22066 29260 23020 29288
rect 18509 29223 18567 29229
rect 18509 29189 18521 29223
rect 18555 29220 18567 29223
rect 19610 29220 19616 29232
rect 18555 29192 19616 29220
rect 18555 29189 18567 29192
rect 18509 29183 18567 29189
rect 19610 29180 19616 29192
rect 19668 29180 19674 29232
rect 21542 29180 21548 29232
rect 21600 29220 21606 29232
rect 22066 29220 22094 29260
rect 23014 29248 23020 29260
rect 23072 29248 23078 29300
rect 23750 29248 23756 29300
rect 23808 29248 23814 29300
rect 24213 29291 24271 29297
rect 24213 29257 24225 29291
rect 24259 29288 24271 29291
rect 24302 29288 24308 29300
rect 24259 29260 24308 29288
rect 24259 29257 24271 29260
rect 24213 29251 24271 29257
rect 24302 29248 24308 29260
rect 24360 29248 24366 29300
rect 24394 29248 24400 29300
rect 24452 29248 24458 29300
rect 21600 29192 22094 29220
rect 23768 29220 23796 29248
rect 23845 29223 23903 29229
rect 23845 29220 23857 29223
rect 23768 29192 23857 29220
rect 21600 29180 21606 29192
rect 23845 29189 23857 29192
rect 23891 29189 23903 29223
rect 23845 29183 23903 29189
rect 19981 29155 20039 29161
rect 19981 29152 19993 29155
rect 18984 29124 19993 29152
rect 18325 29087 18383 29093
rect 18325 29053 18337 29087
rect 18371 29053 18383 29087
rect 18325 29047 18383 29053
rect 18690 29044 18696 29096
rect 18748 29044 18754 29096
rect 18984 29093 19012 29124
rect 19981 29121 19993 29124
rect 20027 29121 20039 29155
rect 19981 29115 20039 29121
rect 20622 29112 20628 29164
rect 20680 29112 20686 29164
rect 24302 29152 24308 29164
rect 24136 29124 24308 29152
rect 18969 29087 19027 29093
rect 18969 29053 18981 29087
rect 19015 29053 19027 29087
rect 18969 29047 19027 29053
rect 19150 29044 19156 29096
rect 19208 29044 19214 29096
rect 19242 29044 19248 29096
rect 19300 29044 19306 29096
rect 19334 29044 19340 29096
rect 19392 29084 19398 29096
rect 19794 29084 19800 29096
rect 19392 29056 19800 29084
rect 19392 29044 19398 29056
rect 19794 29044 19800 29056
rect 19852 29044 19858 29096
rect 21174 29044 21180 29096
rect 21232 29084 21238 29096
rect 21269 29087 21327 29093
rect 21269 29084 21281 29087
rect 21232 29056 21281 29084
rect 21232 29044 21238 29056
rect 21269 29053 21281 29056
rect 21315 29053 21327 29087
rect 21269 29047 21327 29053
rect 21634 29044 21640 29096
rect 21692 29044 21698 29096
rect 23290 29044 23296 29096
rect 23348 29084 23354 29096
rect 24136 29084 24164 29124
rect 24302 29112 24308 29124
rect 24360 29112 24366 29164
rect 24412 29152 24440 29248
rect 24578 29180 24584 29232
rect 24636 29180 24642 29232
rect 25317 29223 25375 29229
rect 25317 29189 25329 29223
rect 25363 29189 25375 29223
rect 25317 29183 25375 29189
rect 24949 29155 25007 29161
rect 24949 29152 24961 29155
rect 24412 29124 24961 29152
rect 23348 29056 24164 29084
rect 23348 29044 23354 29056
rect 17972 28988 18184 29016
rect 17052 28920 17264 28948
rect 18156 28948 18184 28988
rect 18230 28976 18236 29028
rect 18288 28976 18294 29028
rect 20717 29019 20775 29025
rect 20717 29016 20729 29019
rect 18340 28988 20729 29016
rect 18340 28948 18368 28988
rect 20717 28985 20729 28988
rect 20763 28985 20775 29019
rect 20717 28979 20775 28985
rect 24213 29019 24271 29025
rect 24213 28985 24225 29019
rect 24259 29016 24271 29019
rect 24412 29016 24440 29124
rect 24949 29121 24961 29124
rect 24995 29121 25007 29155
rect 24949 29115 25007 29121
rect 25332 29096 25360 29183
rect 24486 29044 24492 29096
rect 24544 29084 24550 29096
rect 24762 29084 24768 29096
rect 24544 29056 24768 29084
rect 24544 29044 24550 29056
rect 24762 29044 24768 29056
rect 24820 29084 24826 29096
rect 25314 29084 25320 29096
rect 24820 29056 25320 29084
rect 24820 29044 24826 29056
rect 25314 29044 25320 29056
rect 25372 29044 25378 29096
rect 26697 29087 26755 29093
rect 26697 29084 26709 29087
rect 26252 29056 26709 29084
rect 24259 28988 24440 29016
rect 24259 28985 24271 28988
rect 24213 28979 24271 28985
rect 26252 28960 26280 29056
rect 26697 29053 26709 29056
rect 26743 29053 26755 29087
rect 26697 29047 26755 29053
rect 26418 28976 26424 29028
rect 26476 29025 26482 29028
rect 26476 28979 26488 29025
rect 26476 28976 26482 28979
rect 18156 28920 18368 28948
rect 18874 28908 18880 28960
rect 18932 28908 18938 28960
rect 21453 28951 21511 28957
rect 21453 28917 21465 28951
rect 21499 28948 21511 28951
rect 21726 28948 21732 28960
rect 21499 28920 21732 28948
rect 21499 28917 21511 28920
rect 21453 28911 21511 28917
rect 21726 28908 21732 28920
rect 21784 28908 21790 28960
rect 24394 28908 24400 28960
rect 24452 28908 24458 28960
rect 24486 28908 24492 28960
rect 24544 28908 24550 28960
rect 26234 28908 26240 28960
rect 26292 28908 26298 28960
rect 552 28858 27576 28880
rect 552 28806 7114 28858
rect 7166 28806 7178 28858
rect 7230 28806 7242 28858
rect 7294 28806 7306 28858
rect 7358 28806 7370 28858
rect 7422 28806 13830 28858
rect 13882 28806 13894 28858
rect 13946 28806 13958 28858
rect 14010 28806 14022 28858
rect 14074 28806 14086 28858
rect 14138 28806 20546 28858
rect 20598 28806 20610 28858
rect 20662 28806 20674 28858
rect 20726 28806 20738 28858
rect 20790 28806 20802 28858
rect 20854 28806 27262 28858
rect 27314 28806 27326 28858
rect 27378 28806 27390 28858
rect 27442 28806 27454 28858
rect 27506 28806 27518 28858
rect 27570 28806 27576 28858
rect 552 28784 27576 28806
rect 3234 28704 3240 28756
rect 3292 28744 3298 28756
rect 6638 28744 6644 28756
rect 3292 28716 3832 28744
rect 3292 28704 3298 28716
rect 2130 28617 2136 28620
rect 2124 28571 2136 28617
rect 2130 28568 2136 28571
rect 2188 28568 2194 28620
rect 3513 28611 3571 28617
rect 3513 28577 3525 28611
rect 3559 28577 3571 28611
rect 3513 28571 3571 28577
rect 1854 28500 1860 28552
rect 1912 28500 1918 28552
rect 3528 28540 3556 28571
rect 3602 28568 3608 28620
rect 3660 28568 3666 28620
rect 3804 28617 3832 28716
rect 4908 28716 6644 28744
rect 4246 28685 4252 28688
rect 4217 28679 4252 28685
rect 4217 28645 4229 28679
rect 4217 28639 4252 28645
rect 4246 28636 4252 28639
rect 4304 28636 4310 28688
rect 4430 28636 4436 28688
rect 4488 28676 4494 28688
rect 4798 28676 4804 28688
rect 4488 28648 4804 28676
rect 4488 28636 4494 28648
rect 4798 28636 4804 28648
rect 4856 28636 4862 28688
rect 3789 28611 3847 28617
rect 3789 28577 3801 28611
rect 3835 28608 3847 28611
rect 4908 28608 4936 28716
rect 6638 28704 6644 28716
rect 6696 28744 6702 28756
rect 7282 28744 7288 28756
rect 6696 28716 7288 28744
rect 6696 28704 6702 28716
rect 7282 28704 7288 28716
rect 7340 28704 7346 28756
rect 7377 28747 7435 28753
rect 7377 28713 7389 28747
rect 7423 28744 7435 28747
rect 7466 28744 7472 28756
rect 7423 28716 7472 28744
rect 7423 28713 7435 28716
rect 7377 28707 7435 28713
rect 7466 28704 7472 28716
rect 7524 28704 7530 28756
rect 7558 28704 7564 28756
rect 7616 28704 7622 28756
rect 10045 28747 10103 28753
rect 10045 28744 10057 28747
rect 8588 28716 10057 28744
rect 7576 28676 7604 28704
rect 5828 28648 6868 28676
rect 5828 28617 5856 28648
rect 3835 28580 4936 28608
rect 5813 28611 5871 28617
rect 3835 28577 3847 28580
rect 3789 28571 3847 28577
rect 5813 28577 5825 28611
rect 5859 28577 5871 28611
rect 5813 28571 5871 28577
rect 5902 28568 5908 28620
rect 5960 28608 5966 28620
rect 6069 28611 6127 28617
rect 6069 28608 6081 28611
rect 5960 28580 6081 28608
rect 5960 28568 5966 28580
rect 6069 28577 6081 28580
rect 6115 28577 6127 28611
rect 6069 28571 6127 28577
rect 6840 28552 6868 28648
rect 7484 28648 7604 28676
rect 7190 28568 7196 28620
rect 7248 28606 7254 28620
rect 7484 28617 7512 28648
rect 7285 28611 7343 28617
rect 7285 28606 7297 28611
rect 7248 28578 7297 28606
rect 7248 28568 7254 28578
rect 7285 28577 7297 28578
rect 7331 28577 7343 28611
rect 7285 28571 7343 28577
rect 7469 28611 7527 28617
rect 7469 28577 7481 28611
rect 7515 28577 7527 28611
rect 7469 28571 7527 28577
rect 7558 28568 7564 28620
rect 7616 28568 7622 28620
rect 7742 28568 7748 28620
rect 7800 28608 7806 28620
rect 8588 28617 8616 28716
rect 10045 28713 10057 28716
rect 10091 28713 10103 28747
rect 10045 28707 10103 28713
rect 8938 28617 8944 28620
rect 8481 28611 8539 28617
rect 8481 28608 8493 28611
rect 7800 28580 8493 28608
rect 7800 28568 7806 28580
rect 8481 28577 8493 28580
rect 8527 28577 8539 28611
rect 8481 28571 8539 28577
rect 8573 28611 8631 28617
rect 8573 28577 8585 28611
rect 8619 28577 8631 28611
rect 8573 28571 8631 28577
rect 8932 28571 8944 28617
rect 8938 28568 8944 28571
rect 8996 28568 9002 28620
rect 10060 28608 10088 28707
rect 15378 28704 15384 28756
rect 15436 28744 15442 28756
rect 15436 28716 15700 28744
rect 15436 28704 15442 28716
rect 11232 28679 11290 28685
rect 11232 28645 11244 28679
rect 11278 28676 11290 28679
rect 11698 28676 11704 28688
rect 11278 28648 11704 28676
rect 11278 28645 11290 28648
rect 11232 28639 11290 28645
rect 11698 28636 11704 28648
rect 11756 28636 11762 28688
rect 14550 28636 14556 28688
rect 14608 28676 14614 28688
rect 15672 28676 15700 28716
rect 15930 28704 15936 28756
rect 15988 28744 15994 28756
rect 16501 28747 16559 28753
rect 16501 28744 16513 28747
rect 15988 28716 16513 28744
rect 15988 28704 15994 28716
rect 16501 28713 16513 28716
rect 16547 28713 16559 28747
rect 16501 28707 16559 28713
rect 17405 28747 17463 28753
rect 17405 28713 17417 28747
rect 17451 28744 17463 28747
rect 18690 28744 18696 28756
rect 17451 28716 18696 28744
rect 17451 28713 17463 28716
rect 17405 28707 17463 28713
rect 18690 28704 18696 28716
rect 18748 28704 18754 28756
rect 24857 28747 24915 28753
rect 24857 28713 24869 28747
rect 24903 28713 24915 28747
rect 24857 28707 24915 28713
rect 16301 28679 16359 28685
rect 14608 28648 15608 28676
rect 15672 28648 16068 28676
rect 14608 28636 14614 28648
rect 10689 28611 10747 28617
rect 10689 28608 10701 28611
rect 10060 28580 10701 28608
rect 10689 28577 10701 28580
rect 10735 28577 10747 28611
rect 10689 28571 10747 28577
rect 12710 28568 12716 28620
rect 12768 28608 12774 28620
rect 15580 28617 15608 28648
rect 13061 28611 13119 28617
rect 13061 28608 13073 28611
rect 12768 28580 13073 28608
rect 12768 28568 12774 28580
rect 13061 28577 13073 28580
rect 13107 28577 13119 28611
rect 13061 28571 13119 28577
rect 15473 28611 15531 28617
rect 15473 28577 15485 28611
rect 15519 28577 15531 28611
rect 15473 28571 15531 28577
rect 15565 28611 15623 28617
rect 15565 28577 15577 28611
rect 15611 28577 15623 28611
rect 15565 28571 15623 28577
rect 4246 28540 4252 28552
rect 3528 28512 4252 28540
rect 1872 28404 1900 28500
rect 3528 28472 3556 28512
rect 4246 28500 4252 28512
rect 4304 28500 4310 28552
rect 6822 28500 6828 28552
rect 6880 28540 6886 28552
rect 8665 28543 8723 28549
rect 8665 28540 8677 28543
rect 6880 28512 8677 28540
rect 6880 28500 6886 28512
rect 8665 28509 8677 28512
rect 8711 28509 8723 28543
rect 8665 28503 8723 28509
rect 2792 28444 3556 28472
rect 3973 28475 4031 28481
rect 2792 28416 2820 28444
rect 3973 28441 3985 28475
rect 4019 28472 4031 28475
rect 4019 28444 4292 28472
rect 4019 28441 4031 28444
rect 3973 28435 4031 28441
rect 2222 28404 2228 28416
rect 1872 28376 2228 28404
rect 2222 28364 2228 28376
rect 2280 28364 2286 28416
rect 2774 28364 2780 28416
rect 2832 28364 2838 28416
rect 3418 28364 3424 28416
rect 3476 28404 3482 28416
rect 4264 28413 4292 28444
rect 6914 28432 6920 28484
rect 6972 28472 6978 28484
rect 7653 28475 7711 28481
rect 7653 28472 7665 28475
rect 6972 28444 7665 28472
rect 6972 28432 6978 28444
rect 7653 28441 7665 28444
rect 7699 28441 7711 28475
rect 7653 28435 7711 28441
rect 7926 28432 7932 28484
rect 7984 28432 7990 28484
rect 4065 28407 4123 28413
rect 4065 28404 4077 28407
rect 3476 28376 4077 28404
rect 3476 28364 3482 28376
rect 4065 28373 4077 28376
rect 4111 28373 4123 28407
rect 4065 28367 4123 28373
rect 4249 28407 4307 28413
rect 4249 28373 4261 28407
rect 4295 28373 4307 28407
rect 4249 28367 4307 28373
rect 7193 28407 7251 28413
rect 7193 28373 7205 28407
rect 7239 28404 7251 28407
rect 7944 28404 7972 28432
rect 7239 28376 7972 28404
rect 8680 28404 8708 28503
rect 10962 28500 10968 28552
rect 11020 28500 11026 28552
rect 12802 28500 12808 28552
rect 12860 28500 12866 28552
rect 14921 28543 14979 28549
rect 14921 28509 14933 28543
rect 14967 28509 14979 28543
rect 15488 28540 15516 28571
rect 15654 28568 15660 28620
rect 15712 28608 15718 28620
rect 15749 28611 15807 28617
rect 15749 28608 15761 28611
rect 15712 28580 15761 28608
rect 15712 28568 15718 28580
rect 15749 28577 15761 28580
rect 15795 28608 15807 28611
rect 15930 28608 15936 28620
rect 15795 28580 15936 28608
rect 15795 28577 15807 28580
rect 15749 28571 15807 28577
rect 15930 28568 15936 28580
rect 15988 28568 15994 28620
rect 16040 28608 16068 28648
rect 16301 28645 16313 28679
rect 16347 28676 16359 28679
rect 16347 28648 16620 28676
rect 16347 28645 16359 28648
rect 16301 28639 16359 28645
rect 16390 28608 16396 28620
rect 16040 28580 16396 28608
rect 16390 28568 16396 28580
rect 16448 28568 16454 28620
rect 16592 28552 16620 28648
rect 16666 28636 16672 28688
rect 16724 28636 16730 28688
rect 17221 28679 17279 28685
rect 17221 28645 17233 28679
rect 17267 28676 17279 28679
rect 17865 28679 17923 28685
rect 17865 28676 17877 28679
rect 17267 28648 17877 28676
rect 17267 28645 17279 28648
rect 17221 28639 17279 28645
rect 17865 28645 17877 28648
rect 17911 28645 17923 28679
rect 17865 28639 17923 28645
rect 18874 28636 18880 28688
rect 18932 28676 18938 28688
rect 19070 28679 19128 28685
rect 19070 28676 19082 28679
rect 18932 28648 19082 28676
rect 18932 28636 18938 28648
rect 19070 28645 19082 28648
rect 19116 28645 19128 28679
rect 21536 28679 21594 28685
rect 19070 28639 19128 28645
rect 19536 28648 21312 28676
rect 16684 28608 16712 28636
rect 17497 28611 17555 28617
rect 17497 28608 17509 28611
rect 16684 28580 17509 28608
rect 17497 28577 17509 28580
rect 17543 28608 17555 28611
rect 17586 28608 17592 28620
rect 17543 28580 17592 28608
rect 17543 28577 17555 28580
rect 17497 28571 17555 28577
rect 17586 28568 17592 28580
rect 17644 28568 17650 28620
rect 17681 28611 17739 28617
rect 17681 28577 17693 28611
rect 17727 28608 17739 28611
rect 17727 28580 18000 28608
rect 17727 28577 17739 28580
rect 17681 28571 17739 28577
rect 16574 28540 16580 28552
rect 15488 28512 16580 28540
rect 14921 28503 14979 28509
rect 10980 28472 11008 28500
rect 9692 28444 11008 28472
rect 14185 28475 14243 28481
rect 9692 28416 9720 28444
rect 14185 28441 14197 28475
rect 14231 28472 14243 28475
rect 14936 28472 14964 28503
rect 16574 28500 16580 28512
rect 16632 28540 16638 28552
rect 17696 28540 17724 28571
rect 16632 28512 17724 28540
rect 16632 28500 16638 28512
rect 14231 28444 15792 28472
rect 14231 28441 14243 28444
rect 14185 28435 14243 28441
rect 9674 28404 9680 28416
rect 8680 28376 9680 28404
rect 7239 28373 7251 28376
rect 7193 28367 7251 28373
rect 9674 28364 9680 28376
rect 9732 28364 9738 28416
rect 10134 28364 10140 28416
rect 10192 28364 10198 28416
rect 12345 28407 12403 28413
rect 12345 28373 12357 28407
rect 12391 28404 12403 28407
rect 13538 28404 13544 28416
rect 12391 28376 13544 28404
rect 12391 28373 12403 28376
rect 12345 28367 12403 28373
rect 13538 28364 13544 28376
rect 13596 28364 13602 28416
rect 14274 28364 14280 28416
rect 14332 28364 14338 28416
rect 15013 28407 15071 28413
rect 15013 28373 15025 28407
rect 15059 28404 15071 28407
rect 15286 28404 15292 28416
rect 15059 28376 15292 28404
rect 15059 28373 15071 28376
rect 15013 28367 15071 28373
rect 15286 28364 15292 28376
rect 15344 28364 15350 28416
rect 15396 28413 15424 28444
rect 15764 28416 15792 28444
rect 16666 28432 16672 28484
rect 16724 28472 16730 28484
rect 17972 28481 18000 28580
rect 19536 28552 19564 28648
rect 21284 28620 21312 28648
rect 21536 28645 21548 28679
rect 21582 28676 21594 28679
rect 21726 28676 21732 28688
rect 21582 28648 21732 28676
rect 21582 28645 21594 28648
rect 21536 28639 21594 28645
rect 21726 28636 21732 28648
rect 21784 28636 21790 28688
rect 19610 28568 19616 28620
rect 19668 28608 19674 28620
rect 19777 28611 19835 28617
rect 19777 28608 19789 28611
rect 19668 28580 19789 28608
rect 19668 28568 19674 28580
rect 19777 28577 19789 28580
rect 19823 28577 19835 28611
rect 19777 28571 19835 28577
rect 21266 28568 21272 28620
rect 21324 28568 21330 28620
rect 23106 28568 23112 28620
rect 23164 28568 23170 28620
rect 24581 28611 24639 28617
rect 24581 28577 24593 28611
rect 24627 28608 24639 28611
rect 24872 28608 24900 28707
rect 25314 28704 25320 28756
rect 25372 28704 25378 28756
rect 25682 28704 25688 28756
rect 25740 28704 25746 28756
rect 25038 28685 25044 28688
rect 25025 28679 25044 28685
rect 25025 28645 25037 28679
rect 25025 28639 25044 28645
rect 25038 28636 25044 28639
rect 25096 28636 25102 28688
rect 25222 28636 25228 28688
rect 25280 28636 25286 28688
rect 25332 28676 25360 28704
rect 25332 28648 25452 28676
rect 24627 28580 24900 28608
rect 25317 28611 25375 28617
rect 24627 28577 24639 28580
rect 24581 28571 24639 28577
rect 25317 28577 25329 28611
rect 25363 28577 25375 28611
rect 25424 28608 25452 28648
rect 25492 28611 25550 28617
rect 25492 28608 25504 28611
rect 25424 28580 25504 28608
rect 25317 28571 25375 28577
rect 25492 28577 25504 28580
rect 25538 28577 25550 28611
rect 25492 28571 25550 28577
rect 19337 28543 19395 28549
rect 19337 28509 19349 28543
rect 19383 28540 19395 28543
rect 19518 28540 19524 28552
rect 19383 28512 19524 28540
rect 19383 28509 19395 28512
rect 19337 28503 19395 28509
rect 19518 28500 19524 28512
rect 19576 28500 19582 28552
rect 25332 28540 25360 28571
rect 25590 28568 25596 28620
rect 25648 28568 25654 28620
rect 25866 28568 25872 28620
rect 25924 28568 25930 28620
rect 26418 28568 26424 28620
rect 26476 28568 26482 28620
rect 24596 28512 25360 28540
rect 16853 28475 16911 28481
rect 16853 28472 16865 28475
rect 16724 28444 16865 28472
rect 16724 28432 16730 28444
rect 16853 28441 16865 28444
rect 16899 28441 16911 28475
rect 16853 28435 16911 28441
rect 17957 28475 18015 28481
rect 17957 28441 17969 28475
rect 18003 28441 18015 28475
rect 17957 28435 18015 28441
rect 24596 28416 24624 28512
rect 24765 28475 24823 28481
rect 24765 28441 24777 28475
rect 24811 28472 24823 28475
rect 26436 28472 26464 28568
rect 24811 28444 26464 28472
rect 24811 28441 24823 28444
rect 24765 28435 24823 28441
rect 15381 28407 15439 28413
rect 15381 28373 15393 28407
rect 15427 28373 15439 28407
rect 15381 28367 15439 28373
rect 15654 28364 15660 28416
rect 15712 28364 15718 28416
rect 15746 28364 15752 28416
rect 15804 28364 15810 28416
rect 16114 28364 16120 28416
rect 16172 28404 16178 28416
rect 16485 28407 16543 28413
rect 16485 28404 16497 28407
rect 16172 28376 16497 28404
rect 16172 28364 16178 28376
rect 16485 28373 16497 28376
rect 16531 28373 16543 28407
rect 16485 28367 16543 28373
rect 16758 28364 16764 28416
rect 16816 28404 16822 28416
rect 17126 28404 17132 28416
rect 16816 28376 17132 28404
rect 16816 28364 16822 28376
rect 17126 28364 17132 28376
rect 17184 28404 17190 28416
rect 17221 28407 17279 28413
rect 17221 28404 17233 28407
rect 17184 28376 17233 28404
rect 17184 28364 17190 28376
rect 17221 28373 17233 28376
rect 17267 28373 17279 28407
rect 17221 28367 17279 28373
rect 20901 28407 20959 28413
rect 20901 28373 20913 28407
rect 20947 28404 20959 28407
rect 21174 28404 21180 28416
rect 20947 28376 21180 28404
rect 20947 28373 20959 28376
rect 20901 28367 20959 28373
rect 21174 28364 21180 28376
rect 21232 28404 21238 28416
rect 22002 28404 22008 28416
rect 21232 28376 22008 28404
rect 21232 28364 21238 28376
rect 22002 28364 22008 28376
rect 22060 28364 22066 28416
rect 22649 28407 22707 28413
rect 22649 28373 22661 28407
rect 22695 28404 22707 28407
rect 22830 28404 22836 28416
rect 22695 28376 22836 28404
rect 22695 28373 22707 28376
rect 22649 28367 22707 28373
rect 22830 28364 22836 28376
rect 22888 28364 22894 28416
rect 22922 28364 22928 28416
rect 22980 28364 22986 28416
rect 24578 28364 24584 28416
rect 24636 28364 24642 28416
rect 25038 28364 25044 28416
rect 25096 28364 25102 28416
rect 25130 28364 25136 28416
rect 25188 28404 25194 28416
rect 25409 28407 25467 28413
rect 25409 28404 25421 28407
rect 25188 28376 25421 28404
rect 25188 28364 25194 28376
rect 25409 28373 25421 28376
rect 25455 28404 25467 28407
rect 25774 28404 25780 28416
rect 25455 28376 25780 28404
rect 25455 28373 25467 28376
rect 25409 28367 25467 28373
rect 25774 28364 25780 28376
rect 25832 28364 25838 28416
rect 26050 28364 26056 28416
rect 26108 28364 26114 28416
rect 552 28314 27416 28336
rect 552 28262 3756 28314
rect 3808 28262 3820 28314
rect 3872 28262 3884 28314
rect 3936 28262 3948 28314
rect 4000 28262 4012 28314
rect 4064 28262 10472 28314
rect 10524 28262 10536 28314
rect 10588 28262 10600 28314
rect 10652 28262 10664 28314
rect 10716 28262 10728 28314
rect 10780 28262 17188 28314
rect 17240 28262 17252 28314
rect 17304 28262 17316 28314
rect 17368 28262 17380 28314
rect 17432 28262 17444 28314
rect 17496 28262 23904 28314
rect 23956 28262 23968 28314
rect 24020 28262 24032 28314
rect 24084 28262 24096 28314
rect 24148 28262 24160 28314
rect 24212 28262 27416 28314
rect 552 28240 27416 28262
rect 2130 28160 2136 28212
rect 2188 28200 2194 28212
rect 2225 28203 2283 28209
rect 2225 28200 2237 28203
rect 2188 28172 2237 28200
rect 2188 28160 2194 28172
rect 2225 28169 2237 28172
rect 2271 28169 2283 28203
rect 3418 28200 3424 28212
rect 2225 28163 2283 28169
rect 2746 28172 3424 28200
rect 2746 28064 2774 28172
rect 3418 28160 3424 28172
rect 3476 28160 3482 28212
rect 4522 28160 4528 28212
rect 4580 28160 4586 28212
rect 7006 28160 7012 28212
rect 7064 28160 7070 28212
rect 9674 28200 9680 28212
rect 9508 28172 9680 28200
rect 3050 28092 3056 28144
rect 3108 28092 3114 28144
rect 3234 28092 3240 28144
rect 3292 28092 3298 28144
rect 6546 28092 6552 28144
rect 6604 28132 6610 28144
rect 6825 28135 6883 28141
rect 6825 28132 6837 28135
rect 6604 28104 6837 28132
rect 6604 28092 6610 28104
rect 6825 28101 6837 28104
rect 6871 28101 6883 28135
rect 6825 28095 6883 28101
rect 2424 28036 2774 28064
rect 2424 28005 2452 28036
rect 2409 27999 2467 28005
rect 2409 27965 2421 27999
rect 2455 27965 2467 27999
rect 2409 27959 2467 27965
rect 2685 27999 2743 28005
rect 2685 27965 2697 27999
rect 2731 27996 2743 27999
rect 2866 27996 2872 28008
rect 2731 27968 2872 27996
rect 2731 27965 2743 27968
rect 2685 27959 2743 27965
rect 2866 27956 2872 27968
rect 2924 27956 2930 28008
rect 3053 27999 3111 28005
rect 3053 27965 3065 27999
rect 3099 27996 3111 27999
rect 3252 27996 3280 28092
rect 6917 28067 6975 28073
rect 6917 28033 6929 28067
rect 6963 28064 6975 28067
rect 7024 28064 7052 28160
rect 6963 28036 7052 28064
rect 6963 28033 6975 28036
rect 6917 28027 6975 28033
rect 8754 28024 8760 28076
rect 8812 28064 8818 28076
rect 9214 28064 9220 28076
rect 8812 28036 9076 28064
rect 8812 28024 8818 28036
rect 3099 27968 3280 27996
rect 6641 27999 6699 28005
rect 3099 27965 3111 27968
rect 3053 27959 3111 27965
rect 6641 27965 6653 27999
rect 6687 27965 6699 27999
rect 6641 27959 6699 27965
rect 2774 27888 2780 27940
rect 2832 27888 2838 27940
rect 2961 27931 3019 27937
rect 2961 27897 2973 27931
rect 3007 27897 3019 27931
rect 2961 27891 3019 27897
rect 2498 27820 2504 27872
rect 2556 27820 2562 27872
rect 2976 27860 3004 27891
rect 3234 27888 3240 27940
rect 3292 27888 3298 27940
rect 3602 27888 3608 27940
rect 3660 27888 3666 27940
rect 6656 27928 6684 27959
rect 6730 27956 6736 28008
rect 6788 27956 6794 28008
rect 7929 27999 7987 28005
rect 7929 27965 7941 27999
rect 7975 27965 7987 27999
rect 7929 27959 7987 27965
rect 7558 27928 7564 27940
rect 6656 27900 7564 27928
rect 7558 27888 7564 27900
rect 7616 27928 7622 27940
rect 7834 27928 7840 27940
rect 7616 27900 7840 27928
rect 7616 27888 7622 27900
rect 7834 27888 7840 27900
rect 7892 27888 7898 27940
rect 3620 27860 3648 27888
rect 7944 27872 7972 27959
rect 8018 27956 8024 28008
rect 8076 27956 8082 28008
rect 8665 27999 8723 28005
rect 8665 27965 8677 27999
rect 8711 27996 8723 27999
rect 8846 27996 8852 28008
rect 8711 27968 8852 27996
rect 8711 27965 8723 27968
rect 8665 27959 8723 27965
rect 8846 27956 8852 27968
rect 8904 27956 8910 28008
rect 9048 28005 9076 28036
rect 9140 28036 9220 28064
rect 9140 28005 9168 28036
rect 9214 28024 9220 28036
rect 9272 28024 9278 28076
rect 9508 28073 9536 28172
rect 9674 28160 9680 28172
rect 9732 28160 9738 28212
rect 12710 28160 12716 28212
rect 12768 28160 12774 28212
rect 13446 28160 13452 28212
rect 13504 28160 13510 28212
rect 14274 28160 14280 28212
rect 14332 28160 14338 28212
rect 15838 28160 15844 28212
rect 15896 28200 15902 28212
rect 16025 28203 16083 28209
rect 16025 28200 16037 28203
rect 15896 28172 16037 28200
rect 15896 28160 15902 28172
rect 16025 28169 16037 28172
rect 16071 28169 16083 28203
rect 16025 28163 16083 28169
rect 16574 28160 16580 28212
rect 16632 28160 16638 28212
rect 16666 28160 16672 28212
rect 16724 28160 16730 28212
rect 21634 28160 21640 28212
rect 21692 28160 21698 28212
rect 21821 28203 21879 28209
rect 21821 28169 21833 28203
rect 21867 28200 21879 28203
rect 22186 28200 22192 28212
rect 21867 28172 22192 28200
rect 21867 28169 21879 28172
rect 21821 28163 21879 28169
rect 22186 28160 22192 28172
rect 22244 28160 22250 28212
rect 22646 28200 22652 28212
rect 22296 28172 22652 28200
rect 10870 28092 10876 28144
rect 10928 28132 10934 28144
rect 13464 28132 13492 28160
rect 10928 28104 11560 28132
rect 10928 28092 10934 28104
rect 11532 28073 11560 28104
rect 13004 28104 13492 28132
rect 9493 28067 9551 28073
rect 9493 28033 9505 28067
rect 9539 28033 9551 28067
rect 9493 28027 9551 28033
rect 11517 28067 11575 28073
rect 11517 28033 11529 28067
rect 11563 28033 11575 28067
rect 11517 28027 11575 28033
rect 9033 27999 9091 28005
rect 9033 27965 9045 27999
rect 9079 27965 9091 27999
rect 9033 27959 9091 27965
rect 9125 27999 9183 28005
rect 9125 27965 9137 27999
rect 9171 27996 9183 27999
rect 9171 27968 9352 27996
rect 9171 27965 9183 27968
rect 9125 27959 9183 27965
rect 8386 27888 8392 27940
rect 8444 27928 8450 27940
rect 9217 27931 9275 27937
rect 9217 27928 9229 27931
rect 8444 27900 9229 27928
rect 8444 27888 8450 27900
rect 9217 27897 9229 27900
rect 9263 27897 9275 27931
rect 9324 27928 9352 27968
rect 9398 27956 9404 28008
rect 9456 27956 9462 28008
rect 11698 27996 11704 28008
rect 9692 27968 11704 27996
rect 9692 27928 9720 27968
rect 11698 27956 11704 27968
rect 11756 27956 11762 28008
rect 12526 27956 12532 28008
rect 12584 27956 12590 28008
rect 12618 27956 12624 28008
rect 12676 27996 12682 28008
rect 13004 28005 13032 28104
rect 14292 28064 14320 28160
rect 15286 28132 15292 28144
rect 13280 28036 14320 28064
rect 14660 28104 15292 28132
rect 13280 28005 13308 28036
rect 12897 27999 12955 28005
rect 12897 27996 12909 27999
rect 12676 27968 12909 27996
rect 12676 27956 12682 27968
rect 12897 27965 12909 27968
rect 12943 27965 12955 27999
rect 12897 27959 12955 27965
rect 12989 27999 13047 28005
rect 12989 27965 13001 27999
rect 13035 27965 13047 27999
rect 12989 27959 13047 27965
rect 13265 27999 13323 28005
rect 13265 27965 13277 27999
rect 13311 27965 13323 27999
rect 13265 27959 13323 27965
rect 13538 27956 13544 28008
rect 13596 27956 13602 28008
rect 13633 27999 13691 28005
rect 13633 27965 13645 27999
rect 13679 27996 13691 27999
rect 14550 27996 14556 28008
rect 13679 27968 14556 27996
rect 13679 27965 13691 27968
rect 13633 27959 13691 27965
rect 14550 27956 14556 27968
rect 14608 27956 14614 28008
rect 14660 28005 14688 28104
rect 15286 28092 15292 28104
rect 15344 28092 15350 28144
rect 16117 28067 16175 28073
rect 15128 28036 15641 28064
rect 14645 27999 14703 28005
rect 14645 27965 14657 27999
rect 14691 27965 14703 27999
rect 14645 27959 14703 27965
rect 14829 27999 14887 28005
rect 14829 27965 14841 27999
rect 14875 27965 14887 27999
rect 14829 27959 14887 27965
rect 14921 27999 14979 28005
rect 14921 27965 14933 27999
rect 14967 27965 14979 27999
rect 14921 27959 14979 27965
rect 9766 27937 9772 27940
rect 9324 27900 9720 27928
rect 9217 27891 9275 27897
rect 9760 27891 9772 27937
rect 9766 27888 9772 27891
rect 9824 27888 9830 27940
rect 2976 27832 3648 27860
rect 7742 27820 7748 27872
rect 7800 27820 7806 27872
rect 7926 27820 7932 27872
rect 7984 27820 7990 27872
rect 8570 27820 8576 27872
rect 8628 27820 8634 27872
rect 8849 27863 8907 27869
rect 8849 27829 8861 27863
rect 8895 27860 8907 27863
rect 9858 27860 9864 27872
rect 8895 27832 9864 27860
rect 8895 27829 8907 27832
rect 8849 27823 8907 27829
rect 9858 27820 9864 27832
rect 9916 27820 9922 27872
rect 10962 27820 10968 27872
rect 11020 27820 11026 27872
rect 11514 27820 11520 27872
rect 11572 27860 11578 27872
rect 11977 27863 12035 27869
rect 11977 27860 11989 27863
rect 11572 27832 11989 27860
rect 11572 27820 11578 27832
rect 11977 27829 11989 27832
rect 12023 27829 12035 27863
rect 12544 27860 12572 27956
rect 13078 27888 13084 27940
rect 13136 27888 13142 27940
rect 14844 27872 14872 27959
rect 14936 27928 14964 27959
rect 15010 27956 15016 28008
rect 15068 27996 15074 28008
rect 15128 27996 15156 28036
rect 15613 28005 15641 28036
rect 16117 28033 16129 28067
rect 16163 28064 16175 28067
rect 16592 28064 16620 28160
rect 16163 28036 16620 28064
rect 16163 28033 16175 28036
rect 16117 28027 16175 28033
rect 16684 28005 16712 28160
rect 16942 28064 16948 28076
rect 16776 28036 16948 28064
rect 16776 28005 16804 28036
rect 16942 28024 16948 28036
rect 17000 28024 17006 28076
rect 21266 28024 21272 28076
rect 21324 28064 21330 28076
rect 22296 28073 22324 28172
rect 22646 28160 22652 28172
rect 22704 28160 22710 28212
rect 23290 28160 23296 28212
rect 23348 28160 23354 28212
rect 24949 28203 25007 28209
rect 24949 28169 24961 28203
rect 24995 28200 25007 28203
rect 25038 28200 25044 28212
rect 24995 28172 25044 28200
rect 24995 28169 25007 28172
rect 24949 28163 25007 28169
rect 25038 28160 25044 28172
rect 25096 28160 25102 28212
rect 25409 28203 25467 28209
rect 25409 28169 25421 28203
rect 25455 28169 25467 28203
rect 25409 28163 25467 28169
rect 25593 28203 25651 28209
rect 25593 28169 25605 28203
rect 25639 28200 25651 28203
rect 25866 28200 25872 28212
rect 25639 28172 25872 28200
rect 25639 28169 25651 28172
rect 25593 28163 25651 28169
rect 23308 28132 23336 28160
rect 25222 28132 25228 28144
rect 23308 28104 25228 28132
rect 25222 28092 25228 28104
rect 25280 28132 25286 28144
rect 25424 28132 25452 28163
rect 25866 28160 25872 28172
rect 25924 28160 25930 28212
rect 26050 28160 26056 28212
rect 26108 28160 26114 28212
rect 25280 28104 25452 28132
rect 25280 28092 25286 28104
rect 22281 28067 22339 28073
rect 22281 28064 22293 28067
rect 21324 28036 22293 28064
rect 21324 28024 21330 28036
rect 22281 28033 22293 28036
rect 22327 28033 22339 28067
rect 22281 28027 22339 28033
rect 23308 28036 25360 28064
rect 15068 27968 15156 27996
rect 15197 27999 15255 28005
rect 15068 27956 15074 27968
rect 15197 27965 15209 27999
rect 15243 27965 15255 27999
rect 15197 27959 15255 27965
rect 15598 27999 15656 28005
rect 15598 27965 15610 27999
rect 15644 27965 15656 27999
rect 15598 27959 15656 27965
rect 16393 27999 16451 28005
rect 16393 27965 16405 27999
rect 16439 27965 16451 27999
rect 16393 27959 16451 27965
rect 16577 27999 16635 28005
rect 16577 27965 16589 27999
rect 16623 27965 16635 27999
rect 16577 27959 16635 27965
rect 16669 27999 16727 28005
rect 16669 27965 16681 27999
rect 16715 27965 16727 27999
rect 16669 27959 16727 27965
rect 16761 27999 16819 28005
rect 16761 27965 16773 27999
rect 16807 27965 16819 27999
rect 16761 27959 16819 27965
rect 15102 27928 15108 27940
rect 14936 27900 15108 27928
rect 15102 27888 15108 27900
rect 15160 27888 15166 27940
rect 15212 27928 15240 27959
rect 15212 27900 15608 27928
rect 15580 27872 15608 27900
rect 16408 27872 16436 27959
rect 14826 27860 14832 27872
rect 12544 27832 14832 27860
rect 11977 27823 12035 27829
rect 14826 27820 14832 27832
rect 14884 27820 14890 27872
rect 15378 27820 15384 27872
rect 15436 27820 15442 27872
rect 15470 27820 15476 27872
rect 15528 27820 15534 27872
rect 15562 27820 15568 27872
rect 15620 27860 15626 27872
rect 15657 27863 15715 27869
rect 15657 27860 15669 27863
rect 15620 27832 15669 27860
rect 15620 27820 15626 27832
rect 15657 27829 15669 27832
rect 15703 27829 15715 27863
rect 15657 27823 15715 27829
rect 16390 27820 16396 27872
rect 16448 27820 16454 27872
rect 16592 27860 16620 27959
rect 17126 27956 17132 28008
rect 17184 27996 17190 28008
rect 17770 27996 17776 28008
rect 17184 27968 17776 27996
rect 17184 27956 17190 27968
rect 17770 27956 17776 27968
rect 17828 27956 17834 28008
rect 22189 27999 22247 28005
rect 22189 27965 22201 27999
rect 22235 27996 22247 27999
rect 22370 27996 22376 28008
rect 22235 27968 22376 27996
rect 22235 27965 22247 27968
rect 22189 27959 22247 27965
rect 22370 27956 22376 27968
rect 22428 27956 22434 28008
rect 23308 27996 23336 28036
rect 22480 27968 23336 27996
rect 17037 27931 17095 27937
rect 17037 27897 17049 27931
rect 17083 27928 17095 27931
rect 17374 27931 17432 27937
rect 17374 27928 17386 27931
rect 17083 27900 17386 27928
rect 17083 27897 17095 27900
rect 17037 27891 17095 27897
rect 17374 27897 17386 27900
rect 17420 27897 17432 27931
rect 17374 27891 17432 27897
rect 19797 27931 19855 27937
rect 19797 27897 19809 27931
rect 19843 27897 19855 27931
rect 19797 27891 19855 27897
rect 21545 27931 21603 27937
rect 21545 27897 21557 27931
rect 21591 27928 21603 27931
rect 22480 27928 22508 27968
rect 23658 27956 23664 28008
rect 23716 27996 23722 28008
rect 23845 27999 23903 28005
rect 23845 27996 23857 27999
rect 23716 27968 23857 27996
rect 23716 27956 23722 27968
rect 23845 27965 23857 27968
rect 23891 27965 23903 27999
rect 23845 27959 23903 27965
rect 24029 27999 24087 28005
rect 24029 27965 24041 27999
rect 24075 27965 24087 27999
rect 24029 27959 24087 27965
rect 24121 27999 24179 28005
rect 24121 27965 24133 27999
rect 24167 27996 24179 27999
rect 24210 27996 24216 28008
rect 24167 27968 24216 27996
rect 24167 27965 24179 27968
rect 24121 27959 24179 27965
rect 21591 27900 22508 27928
rect 22548 27931 22606 27937
rect 21591 27897 21603 27900
rect 21545 27891 21603 27897
rect 22548 27897 22560 27931
rect 22594 27928 22606 27931
rect 22922 27928 22928 27940
rect 22594 27900 22928 27928
rect 22594 27897 22606 27900
rect 22548 27891 22606 27897
rect 16666 27860 16672 27872
rect 16592 27832 16672 27860
rect 16666 27820 16672 27832
rect 16724 27820 16730 27872
rect 17218 27820 17224 27872
rect 17276 27860 17282 27872
rect 18322 27860 18328 27872
rect 17276 27832 18328 27860
rect 17276 27820 17282 27832
rect 18322 27820 18328 27832
rect 18380 27820 18386 27872
rect 18506 27820 18512 27872
rect 18564 27820 18570 27872
rect 19518 27820 19524 27872
rect 19576 27860 19582 27872
rect 19812 27860 19840 27891
rect 22922 27888 22928 27900
rect 22980 27888 22986 27940
rect 23566 27888 23572 27940
rect 23624 27928 23630 27940
rect 24044 27928 24072 27959
rect 24210 27956 24216 27968
rect 24268 27956 24274 28008
rect 24305 27999 24363 28005
rect 24305 27965 24317 27999
rect 24351 27965 24363 27999
rect 24305 27959 24363 27965
rect 23624 27900 24072 27928
rect 24320 27928 24348 27959
rect 24394 27956 24400 28008
rect 24452 27956 24458 28008
rect 24486 27956 24492 28008
rect 24544 27956 24550 28008
rect 25041 27999 25099 28005
rect 25041 27965 25053 27999
rect 25087 27996 25099 27999
rect 25222 27996 25228 28008
rect 25087 27968 25228 27996
rect 25087 27965 25099 27968
rect 25041 27959 25099 27965
rect 25222 27956 25228 27968
rect 25280 27956 25286 28008
rect 24504 27928 24532 27956
rect 25332 27940 25360 28036
rect 24320 27900 24532 27928
rect 23624 27888 23630 27900
rect 19576 27832 19840 27860
rect 19576 27820 19582 27832
rect 21818 27820 21824 27872
rect 21876 27820 21882 27872
rect 22186 27820 22192 27872
rect 22244 27860 22250 27872
rect 22646 27860 22652 27872
rect 22244 27832 22652 27860
rect 22244 27820 22250 27832
rect 22646 27820 22652 27832
rect 22704 27860 22710 27872
rect 23290 27860 23296 27872
rect 22704 27832 23296 27860
rect 22704 27820 22710 27832
rect 23290 27820 23296 27832
rect 23348 27820 23354 27872
rect 23382 27820 23388 27872
rect 23440 27860 23446 27872
rect 23661 27863 23719 27869
rect 23661 27860 23673 27863
rect 23440 27832 23673 27860
rect 23440 27820 23446 27832
rect 23661 27829 23673 27832
rect 23707 27829 23719 27863
rect 24044 27860 24072 27900
rect 24578 27888 24584 27940
rect 24636 27888 24642 27940
rect 24762 27888 24768 27940
rect 24820 27888 24826 27940
rect 25314 27888 25320 27940
rect 25372 27888 25378 27940
rect 26068 27928 26096 28160
rect 26234 27956 26240 28008
rect 26292 27996 26298 28008
rect 27065 27999 27123 28005
rect 27065 27996 27077 27999
rect 26292 27968 27077 27996
rect 26292 27956 26298 27968
rect 27065 27965 27077 27968
rect 27111 27965 27123 27999
rect 27065 27959 27123 27965
rect 26798 27931 26856 27937
rect 26798 27928 26810 27931
rect 26068 27900 26810 27928
rect 26798 27897 26810 27900
rect 26844 27897 26856 27931
rect 26798 27891 26856 27897
rect 24486 27860 24492 27872
rect 24044 27832 24492 27860
rect 23661 27823 23719 27829
rect 24486 27820 24492 27832
rect 24544 27820 24550 27872
rect 25409 27863 25467 27869
rect 25409 27829 25421 27863
rect 25455 27860 25467 27863
rect 25498 27860 25504 27872
rect 25455 27832 25504 27860
rect 25455 27829 25467 27832
rect 25409 27823 25467 27829
rect 25498 27820 25504 27832
rect 25556 27820 25562 27872
rect 25590 27820 25596 27872
rect 25648 27860 25654 27872
rect 25685 27863 25743 27869
rect 25685 27860 25697 27863
rect 25648 27832 25697 27860
rect 25648 27820 25654 27832
rect 25685 27829 25697 27832
rect 25731 27829 25743 27863
rect 25685 27823 25743 27829
rect 552 27770 27576 27792
rect 552 27718 7114 27770
rect 7166 27718 7178 27770
rect 7230 27718 7242 27770
rect 7294 27718 7306 27770
rect 7358 27718 7370 27770
rect 7422 27718 13830 27770
rect 13882 27718 13894 27770
rect 13946 27718 13958 27770
rect 14010 27718 14022 27770
rect 14074 27718 14086 27770
rect 14138 27718 20546 27770
rect 20598 27718 20610 27770
rect 20662 27718 20674 27770
rect 20726 27718 20738 27770
rect 20790 27718 20802 27770
rect 20854 27718 27262 27770
rect 27314 27718 27326 27770
rect 27378 27718 27390 27770
rect 27442 27718 27454 27770
rect 27506 27718 27518 27770
rect 27570 27718 27576 27770
rect 552 27696 27576 27718
rect 2866 27616 2872 27668
rect 2924 27656 2930 27668
rect 3697 27659 3755 27665
rect 3697 27656 3709 27659
rect 2924 27628 3709 27656
rect 2924 27616 2930 27628
rect 3697 27625 3709 27628
rect 3743 27625 3755 27659
rect 4430 27656 4436 27668
rect 3697 27619 3755 27625
rect 4080 27628 4436 27656
rect 2498 27597 2504 27600
rect 2492 27588 2504 27597
rect 2459 27560 2504 27588
rect 2492 27551 2504 27560
rect 2498 27548 2504 27551
rect 2556 27548 2562 27600
rect 4080 27597 4108 27628
rect 4430 27616 4436 27628
rect 4488 27616 4494 27668
rect 7193 27659 7251 27665
rect 7193 27625 7205 27659
rect 7239 27625 7251 27659
rect 7193 27619 7251 27625
rect 8849 27659 8907 27665
rect 8849 27625 8861 27659
rect 8895 27656 8907 27659
rect 8938 27656 8944 27668
rect 8895 27628 8944 27656
rect 8895 27625 8907 27628
rect 8849 27619 8907 27625
rect 3865 27591 3923 27597
rect 3865 27557 3877 27591
rect 3911 27588 3923 27591
rect 4065 27591 4123 27597
rect 3911 27560 4016 27588
rect 3911 27557 3923 27560
rect 3865 27551 3923 27557
rect 2222 27412 2228 27464
rect 2280 27412 2286 27464
rect 3988 27452 4016 27560
rect 4065 27557 4077 27591
rect 4111 27557 4123 27591
rect 4065 27551 4123 27557
rect 4246 27548 4252 27600
rect 4304 27588 4310 27600
rect 4525 27591 4583 27597
rect 4525 27588 4537 27591
rect 4304 27560 4537 27588
rect 4304 27548 4310 27560
rect 4525 27557 4537 27560
rect 4571 27588 4583 27591
rect 7208 27588 7236 27619
rect 8938 27616 8944 27628
rect 8996 27616 9002 27668
rect 9398 27616 9404 27668
rect 9456 27656 9462 27668
rect 9585 27659 9643 27665
rect 9585 27656 9597 27659
rect 9456 27628 9597 27656
rect 9456 27616 9462 27628
rect 9585 27625 9597 27628
rect 9631 27625 9643 27659
rect 9585 27619 9643 27625
rect 9677 27659 9735 27665
rect 9677 27625 9689 27659
rect 9723 27656 9735 27659
rect 9766 27656 9772 27668
rect 9723 27628 9772 27656
rect 9723 27625 9735 27628
rect 9677 27619 9735 27625
rect 9766 27616 9772 27628
rect 9824 27616 9830 27668
rect 10962 27656 10968 27668
rect 10244 27628 10968 27656
rect 4571 27560 4936 27588
rect 4571 27557 4583 27560
rect 4525 27551 4583 27557
rect 4341 27523 4399 27529
rect 4341 27489 4353 27523
rect 4387 27520 4399 27523
rect 4614 27520 4620 27532
rect 4387 27492 4620 27520
rect 4387 27489 4399 27492
rect 4341 27483 4399 27489
rect 4614 27480 4620 27492
rect 4672 27480 4678 27532
rect 4801 27523 4859 27529
rect 4801 27489 4813 27523
rect 4847 27520 4859 27523
rect 4908 27520 4936 27560
rect 5828 27560 6868 27588
rect 7208 27560 7788 27588
rect 4847 27492 4936 27520
rect 4847 27489 4859 27492
rect 4801 27483 4859 27489
rect 5258 27480 5264 27532
rect 5316 27480 5322 27532
rect 5828 27529 5856 27560
rect 6840 27532 6868 27560
rect 5813 27523 5871 27529
rect 5813 27489 5825 27523
rect 5859 27489 5871 27523
rect 6069 27523 6127 27529
rect 6069 27520 6081 27523
rect 5813 27483 5871 27489
rect 5920 27492 6081 27520
rect 4709 27455 4767 27461
rect 4709 27452 4721 27455
rect 3988 27424 4721 27452
rect 4709 27421 4721 27424
rect 4755 27421 4767 27455
rect 5920 27452 5948 27492
rect 6069 27489 6081 27492
rect 6115 27489 6127 27523
rect 6069 27483 6127 27489
rect 6822 27480 6828 27532
rect 6880 27480 6886 27532
rect 7760 27529 7788 27560
rect 8312 27560 10180 27588
rect 7653 27523 7711 27529
rect 7653 27489 7665 27523
rect 7699 27489 7711 27523
rect 7653 27483 7711 27489
rect 7745 27523 7803 27529
rect 7745 27489 7757 27523
rect 7791 27520 7803 27523
rect 7834 27520 7840 27532
rect 7791 27492 7840 27520
rect 7791 27489 7803 27492
rect 7745 27483 7803 27489
rect 4709 27415 4767 27421
rect 5460 27424 5948 27452
rect 7668 27452 7696 27483
rect 7834 27480 7840 27492
rect 7892 27480 7898 27532
rect 8018 27480 8024 27532
rect 8076 27480 8082 27532
rect 8312 27529 8340 27560
rect 10152 27532 10180 27560
rect 8297 27523 8355 27529
rect 8297 27489 8309 27523
rect 8343 27489 8355 27523
rect 8297 27483 8355 27489
rect 8386 27480 8392 27532
rect 8444 27520 8450 27532
rect 8481 27523 8539 27529
rect 8481 27520 8493 27523
rect 8444 27492 8493 27520
rect 8444 27480 8450 27492
rect 8481 27489 8493 27492
rect 8527 27489 8539 27523
rect 8481 27483 8539 27489
rect 8573 27523 8631 27529
rect 8573 27489 8585 27523
rect 8619 27489 8631 27523
rect 8573 27483 8631 27489
rect 8665 27524 8723 27529
rect 8754 27524 8760 27532
rect 8665 27523 8760 27524
rect 8665 27489 8677 27523
rect 8711 27496 8760 27523
rect 8711 27489 8723 27496
rect 8665 27483 8723 27489
rect 8588 27452 8616 27483
rect 8754 27480 8760 27496
rect 8812 27520 8818 27532
rect 9582 27520 9588 27532
rect 8812 27492 9588 27520
rect 8812 27480 8818 27492
rect 9582 27480 9588 27492
rect 9640 27520 9646 27532
rect 9861 27524 9919 27529
rect 9692 27523 9919 27524
rect 9692 27520 9873 27523
rect 9640 27496 9873 27520
rect 9640 27492 9720 27496
rect 9640 27480 9646 27492
rect 9861 27489 9873 27496
rect 9907 27489 9919 27523
rect 9861 27483 9919 27489
rect 9950 27480 9956 27532
rect 10008 27480 10014 27532
rect 10045 27523 10103 27529
rect 10045 27489 10057 27523
rect 10091 27489 10103 27523
rect 10045 27483 10103 27489
rect 7668 27424 8156 27452
rect 8588 27424 8708 27452
rect 3602 27344 3608 27396
rect 3660 27384 3666 27396
rect 5460 27393 5488 27424
rect 5445 27387 5503 27393
rect 3660 27356 4660 27384
rect 3660 27344 3666 27356
rect 4632 27328 4660 27356
rect 5445 27353 5457 27387
rect 5491 27353 5503 27387
rect 8018 27384 8024 27396
rect 5445 27347 5503 27353
rect 6748 27356 8024 27384
rect 3881 27319 3939 27325
rect 3881 27285 3893 27319
rect 3927 27316 3939 27319
rect 4157 27319 4215 27325
rect 4157 27316 4169 27319
rect 3927 27288 4169 27316
rect 3927 27285 3939 27288
rect 3881 27279 3939 27285
rect 4157 27285 4169 27288
rect 4203 27285 4215 27319
rect 4157 27279 4215 27285
rect 4614 27276 4620 27328
rect 4672 27316 4678 27328
rect 6748 27316 6776 27356
rect 8018 27344 8024 27356
rect 8076 27344 8082 27396
rect 8128 27384 8156 27424
rect 8570 27384 8576 27396
rect 8128 27356 8576 27384
rect 8570 27344 8576 27356
rect 8628 27344 8634 27396
rect 8680 27384 8708 27424
rect 8846 27412 8852 27464
rect 8904 27452 8910 27464
rect 8941 27455 8999 27461
rect 8941 27452 8953 27455
rect 8904 27424 8953 27452
rect 8904 27412 8910 27424
rect 8941 27421 8953 27424
rect 8987 27421 8999 27455
rect 8941 27415 8999 27421
rect 10060 27396 10088 27483
rect 10134 27480 10140 27532
rect 10192 27480 10198 27532
rect 10244 27529 10272 27628
rect 10962 27616 10968 27628
rect 11020 27616 11026 27668
rect 14826 27616 14832 27668
rect 14884 27656 14890 27668
rect 14921 27659 14979 27665
rect 14921 27656 14933 27659
rect 14884 27628 14933 27656
rect 14884 27616 14890 27628
rect 14921 27625 14933 27628
rect 14967 27625 14979 27659
rect 14921 27619 14979 27625
rect 16390 27616 16396 27668
rect 16448 27656 16454 27668
rect 16666 27656 16672 27668
rect 16448 27628 16672 27656
rect 16448 27616 16454 27628
rect 16666 27616 16672 27628
rect 16724 27616 16730 27668
rect 17218 27656 17224 27668
rect 16792 27628 17224 27656
rect 16792 27614 16820 27628
rect 17218 27616 17224 27628
rect 17276 27616 17282 27668
rect 17770 27616 17776 27668
rect 17828 27656 17834 27668
rect 17828 27628 19656 27656
rect 17828 27616 17834 27628
rect 10870 27588 10876 27600
rect 10520 27560 10876 27588
rect 10520 27529 10548 27560
rect 10870 27548 10876 27560
rect 10928 27548 10934 27600
rect 10980 27560 12434 27588
rect 10980 27532 11008 27560
rect 10229 27523 10287 27529
rect 10229 27489 10241 27523
rect 10275 27489 10287 27523
rect 10229 27483 10287 27489
rect 10505 27523 10563 27529
rect 10505 27489 10517 27523
rect 10551 27489 10563 27523
rect 10505 27483 10563 27489
rect 10962 27480 10968 27532
rect 11020 27480 11026 27532
rect 11054 27480 11060 27532
rect 11112 27520 11118 27532
rect 11221 27523 11279 27529
rect 11221 27520 11233 27523
rect 11112 27492 11233 27520
rect 11112 27480 11118 27492
rect 11221 27489 11233 27492
rect 11267 27489 11279 27523
rect 12406 27520 12434 27560
rect 15562 27548 15568 27600
rect 15620 27548 15626 27600
rect 16776 27597 16820 27614
rect 16577 27591 16635 27597
rect 16577 27557 16589 27591
rect 16623 27588 16635 27591
rect 16776 27591 16835 27597
rect 16623 27560 16712 27588
rect 16776 27560 16789 27591
rect 16623 27557 16635 27560
rect 16577 27551 16635 27557
rect 12802 27520 12808 27532
rect 12406 27492 12808 27520
rect 11221 27483 11279 27489
rect 12802 27480 12808 27492
rect 12860 27480 12866 27532
rect 12894 27480 12900 27532
rect 12952 27520 12958 27532
rect 13061 27523 13119 27529
rect 13061 27520 13073 27523
rect 12952 27492 13073 27520
rect 12952 27480 12958 27492
rect 13061 27489 13073 27492
rect 13107 27489 13119 27523
rect 13061 27483 13119 27489
rect 14461 27523 14519 27529
rect 14461 27489 14473 27523
rect 14507 27520 14519 27523
rect 14550 27520 14556 27532
rect 14507 27492 14556 27520
rect 14507 27489 14519 27492
rect 14461 27483 14519 27489
rect 14550 27480 14556 27492
rect 14608 27480 14614 27532
rect 14980 27523 15038 27529
rect 14980 27489 14992 27523
rect 15026 27520 15038 27523
rect 15102 27520 15108 27532
rect 15026 27492 15108 27520
rect 15026 27489 15038 27492
rect 14980 27483 15038 27489
rect 15102 27480 15108 27492
rect 15160 27480 15166 27532
rect 16684 27452 16712 27560
rect 16777 27557 16789 27560
rect 16823 27557 16835 27591
rect 16777 27551 16835 27557
rect 18506 27548 18512 27600
rect 18564 27548 18570 27600
rect 16942 27480 16948 27532
rect 17000 27520 17006 27532
rect 17037 27523 17095 27529
rect 17037 27520 17049 27523
rect 17000 27492 17049 27520
rect 17000 27480 17006 27492
rect 17037 27489 17049 27492
rect 17083 27489 17095 27523
rect 17037 27483 17095 27489
rect 17681 27523 17739 27529
rect 17681 27489 17693 27523
rect 17727 27520 17739 27523
rect 17957 27523 18015 27529
rect 17957 27520 17969 27523
rect 17727 27492 17969 27520
rect 17727 27489 17739 27492
rect 17681 27483 17739 27489
rect 17957 27489 17969 27492
rect 18003 27520 18015 27523
rect 18524 27520 18552 27548
rect 18003 27492 18552 27520
rect 18003 27489 18015 27492
rect 17957 27483 18015 27489
rect 17696 27452 17724 27483
rect 19334 27480 19340 27532
rect 19392 27529 19398 27532
rect 19392 27483 19404 27529
rect 19392 27480 19398 27483
rect 19518 27480 19524 27532
rect 19576 27520 19582 27532
rect 19628 27529 19656 27628
rect 21542 27616 21548 27668
rect 21600 27656 21606 27668
rect 22925 27659 22983 27665
rect 21600 27628 22232 27656
rect 21600 27616 21606 27628
rect 20070 27548 20076 27600
rect 20128 27548 20134 27600
rect 21818 27548 21824 27600
rect 21876 27588 21882 27600
rect 22097 27591 22155 27597
rect 22097 27588 22109 27591
rect 21876 27560 22109 27588
rect 21876 27548 21882 27560
rect 22097 27557 22109 27560
rect 22143 27557 22155 27591
rect 22097 27551 22155 27557
rect 19613 27523 19671 27529
rect 19613 27520 19625 27523
rect 19576 27492 19625 27520
rect 19576 27480 19582 27492
rect 19613 27489 19625 27492
rect 19659 27489 19671 27523
rect 19613 27483 19671 27489
rect 19794 27480 19800 27532
rect 19852 27520 19858 27532
rect 19889 27523 19947 27529
rect 19889 27520 19901 27523
rect 19852 27492 19901 27520
rect 19852 27480 19858 27492
rect 19889 27489 19901 27492
rect 19935 27489 19947 27523
rect 19889 27483 19947 27489
rect 19978 27480 19984 27532
rect 20036 27480 20042 27532
rect 20257 27523 20315 27529
rect 20257 27489 20269 27523
rect 20303 27520 20315 27523
rect 21269 27523 21327 27529
rect 21269 27520 21281 27523
rect 20303 27492 21281 27520
rect 20303 27489 20315 27492
rect 20257 27483 20315 27489
rect 21269 27489 21281 27492
rect 21315 27489 21327 27523
rect 21269 27483 21327 27489
rect 21726 27480 21732 27532
rect 21784 27520 21790 27532
rect 22204 27529 22232 27628
rect 22925 27625 22937 27659
rect 22971 27656 22983 27659
rect 23106 27656 23112 27668
rect 22971 27628 23112 27656
rect 22971 27625 22983 27628
rect 22925 27619 22983 27625
rect 23106 27616 23112 27628
rect 23164 27616 23170 27668
rect 24578 27656 24584 27668
rect 24044 27628 24584 27656
rect 22738 27548 22744 27600
rect 22796 27548 22802 27600
rect 22830 27548 22836 27600
rect 22888 27588 22894 27600
rect 22888 27560 23060 27588
rect 22888 27548 22894 27560
rect 22005 27523 22063 27529
rect 22180 27526 22238 27529
rect 22005 27520 22017 27523
rect 21784 27492 22017 27520
rect 21784 27480 21790 27492
rect 22005 27489 22017 27492
rect 22051 27489 22063 27523
rect 22005 27483 22063 27489
rect 22173 27523 22238 27526
rect 22173 27489 22192 27523
rect 22226 27489 22238 27523
rect 22173 27483 22238 27489
rect 16684 27424 17724 27452
rect 21821 27455 21879 27461
rect 21821 27421 21833 27455
rect 21867 27452 21879 27455
rect 22173 27452 22201 27483
rect 22278 27480 22284 27532
rect 22336 27520 22342 27532
rect 22922 27520 22928 27532
rect 22336 27492 22928 27520
rect 22336 27480 22342 27492
rect 22922 27480 22928 27492
rect 22980 27480 22986 27532
rect 23032 27529 23060 27560
rect 23017 27523 23075 27529
rect 23017 27489 23029 27523
rect 23063 27489 23075 27523
rect 23017 27483 23075 27489
rect 23109 27455 23167 27461
rect 23109 27452 23121 27455
rect 21867 27424 21901 27452
rect 22173 27424 23121 27452
rect 21867 27421 21879 27424
rect 21821 27415 21879 27421
rect 23109 27421 23121 27424
rect 23155 27421 23167 27455
rect 23109 27415 23167 27421
rect 9306 27384 9312 27396
rect 8680 27356 9312 27384
rect 9306 27344 9312 27356
rect 9364 27344 9370 27396
rect 10042 27344 10048 27396
rect 10100 27344 10106 27396
rect 12345 27387 12403 27393
rect 12345 27353 12357 27387
rect 12391 27384 12403 27387
rect 12526 27384 12532 27396
rect 12391 27356 12532 27384
rect 12391 27353 12403 27356
rect 12345 27347 12403 27353
rect 12526 27344 12532 27356
rect 12584 27344 12590 27396
rect 14182 27344 14188 27396
rect 14240 27384 14246 27396
rect 15010 27384 15016 27396
rect 14240 27356 15016 27384
rect 14240 27344 14246 27356
rect 15010 27344 15016 27356
rect 15068 27344 15074 27396
rect 15105 27387 15163 27393
rect 15105 27353 15117 27387
rect 15151 27384 15163 27387
rect 15194 27384 15200 27396
rect 15151 27356 15200 27384
rect 15151 27353 15163 27356
rect 15105 27347 15163 27353
rect 15194 27344 15200 27356
rect 15252 27344 15258 27396
rect 15930 27384 15936 27396
rect 15304 27356 15936 27384
rect 4672 27288 6776 27316
rect 4672 27276 4678 27288
rect 7282 27276 7288 27328
rect 7340 27316 7346 27328
rect 7469 27319 7527 27325
rect 7469 27316 7481 27319
rect 7340 27288 7481 27316
rect 7340 27276 7346 27288
rect 7469 27285 7481 27288
rect 7515 27285 7527 27319
rect 7469 27279 7527 27285
rect 7926 27276 7932 27328
rect 7984 27316 7990 27328
rect 10413 27319 10471 27325
rect 10413 27316 10425 27319
rect 7984 27288 10425 27316
rect 7984 27276 7990 27288
rect 10413 27285 10425 27288
rect 10459 27285 10471 27319
rect 10413 27279 10471 27285
rect 14553 27319 14611 27325
rect 14553 27285 14565 27319
rect 14599 27316 14611 27319
rect 15304 27316 15332 27356
rect 15930 27344 15936 27356
rect 15988 27344 15994 27396
rect 18414 27384 18420 27396
rect 16500 27356 18420 27384
rect 16500 27328 16528 27356
rect 18414 27344 18420 27356
rect 18472 27344 18478 27396
rect 21836 27384 21864 27415
rect 22278 27384 22284 27396
rect 21744 27356 22284 27384
rect 14599 27288 15332 27316
rect 14599 27285 14611 27288
rect 14553 27279 14611 27285
rect 15378 27276 15384 27328
rect 15436 27316 15442 27328
rect 15565 27319 15623 27325
rect 15565 27316 15577 27319
rect 15436 27288 15577 27316
rect 15436 27276 15442 27288
rect 15565 27285 15577 27288
rect 15611 27285 15623 27319
rect 15565 27279 15623 27285
rect 15749 27319 15807 27325
rect 15749 27285 15761 27319
rect 15795 27316 15807 27319
rect 15838 27316 15844 27328
rect 15795 27288 15844 27316
rect 15795 27285 15807 27288
rect 15749 27279 15807 27285
rect 15838 27276 15844 27288
rect 15896 27276 15902 27328
rect 16482 27276 16488 27328
rect 16540 27276 16546 27328
rect 16574 27276 16580 27328
rect 16632 27316 16638 27328
rect 16761 27319 16819 27325
rect 16761 27316 16773 27319
rect 16632 27288 16773 27316
rect 16632 27276 16638 27288
rect 16761 27285 16773 27288
rect 16807 27285 16819 27319
rect 16761 27279 16819 27285
rect 16942 27276 16948 27328
rect 17000 27276 17006 27328
rect 17770 27276 17776 27328
rect 17828 27316 17834 27328
rect 17865 27319 17923 27325
rect 17865 27316 17877 27319
rect 17828 27288 17877 27316
rect 17828 27276 17834 27288
rect 17865 27285 17877 27288
rect 17911 27285 17923 27319
rect 17865 27279 17923 27285
rect 18046 27276 18052 27328
rect 18104 27316 18110 27328
rect 18233 27319 18291 27325
rect 18233 27316 18245 27319
rect 18104 27288 18245 27316
rect 18104 27276 18110 27288
rect 18233 27285 18245 27288
rect 18279 27285 18291 27319
rect 18233 27279 18291 27285
rect 19705 27319 19763 27325
rect 19705 27285 19717 27319
rect 19751 27316 19763 27319
rect 19794 27316 19800 27328
rect 19751 27288 19800 27316
rect 19751 27285 19763 27288
rect 19705 27279 19763 27285
rect 19794 27276 19800 27288
rect 19852 27276 19858 27328
rect 20898 27276 20904 27328
rect 20956 27316 20962 27328
rect 21744 27316 21772 27356
rect 22278 27344 22284 27356
rect 22336 27344 22342 27396
rect 22373 27387 22431 27393
rect 22373 27353 22385 27387
rect 22419 27384 22431 27387
rect 24044 27384 24072 27628
rect 24578 27616 24584 27628
rect 24636 27656 24642 27668
rect 24949 27659 25007 27665
rect 24949 27656 24961 27659
rect 24636 27628 24961 27656
rect 24636 27616 24642 27628
rect 24949 27625 24961 27628
rect 24995 27656 25007 27659
rect 25383 27659 25441 27665
rect 25383 27656 25395 27659
rect 24995 27628 25395 27656
rect 24995 27625 25007 27628
rect 24949 27619 25007 27625
rect 25383 27625 25395 27628
rect 25429 27625 25441 27659
rect 25383 27619 25441 27625
rect 25498 27616 25504 27668
rect 25556 27656 25562 27668
rect 25685 27659 25743 27665
rect 25685 27656 25697 27659
rect 25556 27628 25697 27656
rect 25556 27616 25562 27628
rect 25685 27625 25697 27628
rect 25731 27625 25743 27659
rect 25685 27619 25743 27625
rect 24397 27591 24455 27597
rect 24397 27557 24409 27591
rect 24443 27588 24455 27591
rect 24670 27588 24676 27600
rect 24443 27560 24676 27588
rect 24443 27557 24455 27560
rect 24397 27551 24455 27557
rect 24670 27548 24676 27560
rect 24728 27548 24734 27600
rect 24765 27591 24823 27597
rect 24765 27557 24777 27591
rect 24811 27588 24823 27591
rect 25590 27588 25596 27600
rect 24811 27560 25596 27588
rect 24811 27557 24823 27560
rect 24765 27551 24823 27557
rect 25590 27548 25596 27560
rect 25648 27548 25654 27600
rect 24489 27523 24547 27529
rect 24489 27489 24501 27523
rect 24535 27520 24547 27523
rect 24578 27520 24584 27532
rect 24535 27492 24584 27520
rect 24535 27489 24547 27492
rect 24489 27483 24547 27489
rect 24578 27480 24584 27492
rect 24636 27480 24642 27532
rect 24854 27480 24860 27532
rect 24912 27480 24918 27532
rect 25682 27480 25688 27532
rect 25740 27480 25746 27532
rect 25774 27480 25780 27532
rect 25832 27520 25838 27532
rect 25869 27523 25927 27529
rect 25869 27520 25881 27523
rect 25832 27492 25881 27520
rect 25832 27480 25838 27492
rect 25869 27489 25881 27492
rect 25915 27489 25927 27523
rect 25869 27483 25927 27489
rect 24872 27452 24900 27480
rect 24872 27424 25452 27452
rect 22419 27356 24072 27384
rect 22419 27353 22431 27356
rect 22373 27347 22431 27353
rect 20956 27288 21772 27316
rect 20956 27276 20962 27288
rect 22186 27276 22192 27328
rect 22244 27316 22250 27328
rect 22388 27316 22416 27347
rect 22244 27288 22416 27316
rect 22244 27276 22250 27288
rect 22646 27276 22652 27328
rect 22704 27316 22710 27328
rect 22741 27319 22799 27325
rect 22741 27316 22753 27319
rect 22704 27288 22753 27316
rect 22704 27276 22710 27288
rect 22741 27285 22753 27288
rect 22787 27285 22799 27319
rect 22741 27279 22799 27285
rect 25130 27276 25136 27328
rect 25188 27276 25194 27328
rect 25222 27276 25228 27328
rect 25280 27276 25286 27328
rect 25424 27325 25452 27424
rect 25409 27319 25467 27325
rect 25409 27285 25421 27319
rect 25455 27285 25467 27319
rect 25409 27279 25467 27285
rect 552 27226 27416 27248
rect 552 27174 3756 27226
rect 3808 27174 3820 27226
rect 3872 27174 3884 27226
rect 3936 27174 3948 27226
rect 4000 27174 4012 27226
rect 4064 27174 10472 27226
rect 10524 27174 10536 27226
rect 10588 27174 10600 27226
rect 10652 27174 10664 27226
rect 10716 27174 10728 27226
rect 10780 27174 17188 27226
rect 17240 27174 17252 27226
rect 17304 27174 17316 27226
rect 17368 27174 17380 27226
rect 17432 27174 17444 27226
rect 17496 27174 23904 27226
rect 23956 27174 23968 27226
rect 24020 27174 24032 27226
rect 24084 27174 24096 27226
rect 24148 27174 24160 27226
rect 24212 27174 27416 27226
rect 552 27152 27416 27174
rect 4246 27072 4252 27124
rect 4304 27072 4310 27124
rect 5077 27115 5135 27121
rect 5077 27081 5089 27115
rect 5123 27081 5135 27115
rect 5077 27075 5135 27081
rect 4264 27044 4292 27072
rect 4709 27047 4767 27053
rect 4709 27044 4721 27047
rect 4264 27016 4721 27044
rect 4709 27013 4721 27016
rect 4755 27013 4767 27047
rect 5092 27044 5120 27075
rect 5258 27072 5264 27124
rect 5316 27072 5322 27124
rect 5350 27072 5356 27124
rect 5408 27072 5414 27124
rect 5537 27115 5595 27121
rect 5537 27081 5549 27115
rect 5583 27112 5595 27115
rect 6086 27112 6092 27124
rect 5583 27084 6092 27112
rect 5583 27081 5595 27084
rect 5537 27075 5595 27081
rect 6086 27072 6092 27084
rect 6144 27072 6150 27124
rect 6730 27072 6736 27124
rect 6788 27072 6794 27124
rect 7929 27115 7987 27121
rect 6840 27084 7880 27112
rect 6181 27047 6239 27053
rect 6181 27044 6193 27047
rect 5092 27016 5396 27044
rect 4709 27007 4767 27013
rect 4724 26976 4752 27007
rect 5258 26976 5264 26988
rect 4724 26948 5264 26976
rect 5258 26936 5264 26948
rect 5316 26936 5322 26988
rect 2225 26911 2283 26917
rect 2225 26877 2237 26911
rect 2271 26908 2283 26911
rect 2498 26908 2504 26920
rect 2271 26880 2504 26908
rect 2271 26877 2283 26880
rect 2225 26871 2283 26877
rect 2498 26868 2504 26880
rect 2556 26868 2562 26920
rect 5074 26868 5080 26920
rect 5132 26868 5138 26920
rect 5368 26908 5396 27016
rect 5644 27016 6193 27044
rect 5644 26908 5672 27016
rect 6181 27013 6193 27016
rect 6227 27013 6239 27047
rect 6181 27007 6239 27013
rect 5997 26911 6055 26917
rect 5997 26908 6009 26911
rect 5368 26880 5672 26908
rect 5736 26880 6009 26908
rect 2314 26800 2320 26852
rect 2372 26840 2378 26852
rect 2409 26843 2467 26849
rect 2409 26840 2421 26843
rect 2372 26812 2421 26840
rect 2372 26800 2378 26812
rect 2409 26809 2421 26812
rect 2455 26809 2467 26843
rect 5092 26840 5120 26868
rect 5736 26849 5764 26880
rect 5997 26877 6009 26880
rect 6043 26908 6055 26911
rect 6840 26908 6868 27084
rect 7009 27047 7067 27053
rect 7009 27013 7021 27047
rect 7055 27044 7067 27047
rect 7466 27044 7472 27056
rect 7055 27016 7472 27044
rect 7055 27013 7067 27016
rect 7009 27007 7067 27013
rect 7466 27004 7472 27016
rect 7524 27004 7530 27056
rect 7852 26988 7880 27084
rect 7929 27081 7941 27115
rect 7975 27112 7987 27115
rect 8389 27115 8447 27121
rect 8389 27112 8401 27115
rect 7975 27084 8401 27112
rect 7975 27081 7987 27084
rect 7929 27075 7987 27081
rect 8389 27081 8401 27084
rect 8435 27081 8447 27115
rect 8389 27075 8447 27081
rect 8846 27072 8852 27124
rect 8904 27112 8910 27124
rect 8941 27115 8999 27121
rect 8941 27112 8953 27115
rect 8904 27084 8953 27112
rect 8904 27072 8910 27084
rect 8941 27081 8953 27084
rect 8987 27081 8999 27115
rect 8941 27075 8999 27081
rect 9030 27072 9036 27124
rect 9088 27112 9094 27124
rect 10042 27112 10048 27124
rect 9088 27084 10048 27112
rect 9088 27072 9094 27084
rect 10042 27072 10048 27084
rect 10100 27072 10106 27124
rect 10965 27115 11023 27121
rect 10965 27081 10977 27115
rect 11011 27112 11023 27115
rect 11054 27112 11060 27124
rect 11011 27084 11060 27112
rect 11011 27081 11023 27084
rect 10965 27075 11023 27081
rect 11054 27072 11060 27084
rect 11112 27072 11118 27124
rect 12802 27072 12808 27124
rect 12860 27112 12866 27124
rect 12897 27115 12955 27121
rect 12897 27112 12909 27115
rect 12860 27084 12909 27112
rect 12860 27072 12866 27084
rect 12897 27081 12909 27084
rect 12943 27081 12955 27115
rect 12897 27075 12955 27081
rect 15194 27072 15200 27124
rect 15252 27072 15258 27124
rect 16942 27072 16948 27124
rect 17000 27072 17006 27124
rect 17681 27115 17739 27121
rect 17681 27081 17693 27115
rect 17727 27112 17739 27115
rect 17957 27115 18015 27121
rect 17957 27112 17969 27115
rect 17727 27084 17969 27112
rect 17727 27081 17739 27084
rect 17681 27075 17739 27081
rect 17957 27081 17969 27084
rect 18003 27081 18015 27115
rect 17957 27075 18015 27081
rect 18046 27072 18052 27124
rect 18104 27072 18110 27124
rect 18322 27072 18328 27124
rect 18380 27072 18386 27124
rect 18414 27072 18420 27124
rect 18472 27072 18478 27124
rect 19153 27115 19211 27121
rect 19153 27081 19165 27115
rect 19199 27112 19211 27115
rect 19334 27112 19340 27124
rect 19199 27084 19340 27112
rect 19199 27081 19211 27084
rect 19153 27075 19211 27081
rect 19334 27072 19340 27084
rect 19392 27072 19398 27124
rect 19545 27084 20475 27112
rect 7193 26979 7251 26985
rect 7193 26945 7205 26979
rect 7239 26976 7251 26979
rect 7282 26976 7288 26988
rect 7239 26948 7288 26976
rect 7239 26945 7251 26948
rect 7193 26939 7251 26945
rect 7282 26936 7288 26948
rect 7340 26936 7346 26988
rect 7742 26936 7748 26988
rect 7800 26936 7806 26988
rect 7834 26936 7840 26988
rect 7892 26976 7898 26988
rect 8757 26979 8815 26985
rect 8757 26976 8769 26979
rect 7892 26948 8769 26976
rect 7892 26936 7898 26948
rect 8757 26945 8769 26948
rect 8803 26945 8815 26979
rect 8757 26939 8815 26945
rect 14182 26936 14188 26988
rect 14240 26936 14246 26988
rect 6043 26880 6868 26908
rect 6917 26911 6975 26917
rect 6043 26877 6055 26880
rect 5997 26871 6055 26877
rect 6917 26877 6929 26911
rect 6963 26877 6975 26911
rect 6917 26871 6975 26877
rect 7101 26911 7159 26917
rect 7101 26877 7113 26911
rect 7147 26877 7159 26911
rect 7101 26871 7159 26877
rect 5505 26843 5563 26849
rect 5505 26840 5517 26843
rect 5092 26812 5517 26840
rect 2409 26803 2467 26809
rect 5505 26809 5517 26812
rect 5551 26809 5563 26843
rect 5505 26803 5563 26809
rect 5721 26843 5779 26849
rect 5721 26809 5733 26843
rect 5767 26809 5779 26843
rect 5721 26803 5779 26809
rect 5810 26800 5816 26852
rect 5868 26800 5874 26852
rect 6932 26784 6960 26871
rect 2590 26732 2596 26784
rect 2648 26732 2654 26784
rect 2682 26732 2688 26784
rect 2740 26772 2746 26784
rect 5077 26775 5135 26781
rect 5077 26772 5089 26775
rect 2740 26744 5089 26772
rect 2740 26732 2746 26744
rect 5077 26741 5089 26744
rect 5123 26741 5135 26775
rect 5077 26735 5135 26741
rect 6914 26732 6920 26784
rect 6972 26732 6978 26784
rect 7006 26732 7012 26784
rect 7064 26772 7070 26784
rect 7116 26772 7144 26871
rect 7300 26840 7328 26936
rect 7377 26911 7435 26917
rect 7377 26877 7389 26911
rect 7423 26908 7435 26911
rect 7760 26908 7788 26936
rect 7423 26880 7788 26908
rect 8021 26911 8079 26917
rect 7423 26877 7435 26880
rect 7377 26871 7435 26877
rect 8021 26877 8033 26911
rect 8067 26877 8079 26911
rect 8021 26871 8079 26877
rect 8036 26840 8064 26871
rect 8570 26868 8576 26920
rect 8628 26868 8634 26920
rect 9674 26868 9680 26920
rect 9732 26908 9738 26920
rect 10321 26911 10379 26917
rect 10321 26908 10333 26911
rect 9732 26880 10333 26908
rect 9732 26868 9738 26880
rect 10321 26877 10333 26880
rect 10367 26877 10379 26911
rect 10321 26871 10379 26877
rect 11149 26911 11207 26917
rect 11149 26877 11161 26911
rect 11195 26908 11207 26911
rect 11422 26908 11428 26920
rect 11195 26880 11428 26908
rect 11195 26877 11207 26880
rect 11149 26871 11207 26877
rect 11422 26868 11428 26880
rect 11480 26868 11486 26920
rect 11514 26868 11520 26920
rect 11572 26868 11578 26920
rect 11606 26868 11612 26920
rect 11664 26868 11670 26920
rect 12802 26868 12808 26920
rect 12860 26908 12866 26920
rect 13630 26908 13636 26920
rect 12860 26880 13636 26908
rect 12860 26868 12866 26880
rect 13630 26868 13636 26880
rect 13688 26868 13694 26920
rect 15212 26908 15240 27072
rect 15286 27004 15292 27056
rect 15344 27044 15350 27056
rect 15841 27047 15899 27053
rect 15841 27044 15853 27047
rect 15344 27016 15853 27044
rect 15344 27004 15350 27016
rect 15841 27013 15853 27016
rect 15887 27013 15899 27047
rect 15841 27007 15899 27013
rect 15381 26911 15439 26917
rect 15381 26908 15393 26911
rect 15212 26880 15393 26908
rect 15381 26877 15393 26880
rect 15427 26877 15439 26911
rect 15381 26871 15439 26877
rect 15473 26911 15531 26917
rect 15473 26877 15485 26911
rect 15519 26908 15531 26911
rect 15654 26908 15660 26920
rect 15519 26880 15660 26908
rect 15519 26877 15531 26880
rect 15473 26871 15531 26877
rect 15654 26868 15660 26880
rect 15712 26868 15718 26920
rect 16960 26908 16988 27072
rect 17129 27047 17187 27053
rect 17129 27013 17141 27047
rect 17175 27044 17187 27047
rect 17862 27044 17868 27056
rect 17175 27016 17868 27044
rect 17175 27013 17187 27016
rect 17129 27007 17187 27013
rect 17862 27004 17868 27016
rect 17920 27004 17926 27056
rect 18064 26976 18092 27072
rect 18141 27047 18199 27053
rect 18141 27013 18153 27047
rect 18187 27013 18199 27047
rect 18432 27044 18460 27072
rect 19545 27044 19573 27084
rect 18432 27016 19573 27044
rect 20447 27044 20475 27084
rect 20898 27072 20904 27124
rect 20956 27072 20962 27124
rect 21450 27072 21456 27124
rect 21508 27112 21514 27124
rect 21637 27115 21695 27121
rect 21637 27112 21649 27115
rect 21508 27084 21649 27112
rect 21508 27072 21514 27084
rect 21637 27081 21649 27084
rect 21683 27081 21695 27115
rect 21637 27075 21695 27081
rect 21910 27072 21916 27124
rect 21968 27072 21974 27124
rect 22097 27115 22155 27121
rect 22097 27081 22109 27115
rect 22143 27112 22155 27115
rect 22462 27112 22468 27124
rect 22143 27084 22468 27112
rect 22143 27081 22155 27084
rect 22097 27075 22155 27081
rect 22462 27072 22468 27084
rect 22520 27112 22526 27124
rect 22520 27084 22600 27112
rect 22520 27072 22526 27084
rect 21266 27044 21272 27056
rect 20447 27016 21272 27044
rect 18141 27007 18199 27013
rect 17236 26948 18092 26976
rect 18156 26976 18184 27007
rect 21266 27004 21272 27016
rect 21324 27004 21330 27056
rect 21821 27047 21879 27053
rect 21821 27013 21833 27047
rect 21867 27044 21879 27047
rect 22572 27044 22600 27084
rect 22738 27072 22744 27124
rect 22796 27072 22802 27124
rect 22830 27072 22836 27124
rect 22888 27072 22894 27124
rect 23382 27072 23388 27124
rect 23440 27072 23446 27124
rect 22848 27044 22876 27072
rect 21867 27016 21956 27044
rect 22572 27016 22876 27044
rect 21867 27013 21879 27016
rect 21821 27007 21879 27013
rect 18156 26948 19012 26976
rect 17236 26917 17264 26948
rect 17037 26911 17095 26917
rect 17037 26908 17049 26911
rect 16960 26880 17049 26908
rect 17037 26877 17049 26880
rect 17083 26877 17095 26911
rect 17037 26871 17095 26877
rect 17221 26911 17279 26917
rect 17221 26877 17233 26911
rect 17267 26908 17279 26911
rect 17494 26910 17500 26920
rect 17420 26908 17500 26910
rect 17267 26882 17500 26908
rect 17267 26880 17448 26882
rect 17267 26877 17279 26880
rect 17221 26871 17279 26877
rect 7300 26812 8064 26840
rect 9858 26800 9864 26852
rect 9916 26840 9922 26852
rect 10054 26843 10112 26849
rect 10054 26840 10066 26843
rect 9916 26812 10066 26840
rect 9916 26800 9922 26812
rect 10054 26809 10066 26812
rect 10100 26809 10112 26843
rect 10054 26803 10112 26809
rect 11054 26800 11060 26852
rect 11112 26840 11118 26852
rect 11241 26843 11299 26849
rect 11241 26840 11253 26843
rect 11112 26812 11253 26840
rect 11112 26800 11118 26812
rect 11241 26809 11253 26812
rect 11287 26809 11299 26843
rect 11241 26803 11299 26809
rect 11330 26800 11336 26852
rect 11388 26800 11394 26852
rect 15105 26843 15163 26849
rect 15105 26809 15117 26843
rect 15151 26840 15163 26843
rect 15562 26840 15568 26852
rect 15151 26812 15568 26840
rect 15151 26809 15163 26812
rect 15105 26803 15163 26809
rect 15562 26800 15568 26812
rect 15620 26840 15626 26852
rect 16209 26843 16267 26849
rect 16209 26840 16221 26843
rect 15620 26812 16221 26840
rect 15620 26800 15626 26812
rect 16209 26809 16221 26812
rect 16255 26809 16267 26843
rect 17052 26840 17080 26871
rect 17494 26868 17500 26882
rect 17552 26868 17558 26920
rect 18233 26911 18291 26917
rect 18233 26908 18245 26911
rect 17880 26880 18245 26908
rect 17313 26843 17371 26849
rect 17313 26840 17325 26843
rect 17052 26812 17325 26840
rect 16209 26803 16267 26809
rect 17313 26809 17325 26812
rect 17359 26809 17371 26843
rect 17313 26803 17371 26809
rect 7650 26772 7656 26784
rect 7064 26744 7656 26772
rect 7064 26732 7070 26744
rect 7650 26732 7656 26744
rect 7708 26732 7714 26784
rect 13538 26732 13544 26784
rect 13596 26732 13602 26784
rect 15289 26775 15347 26781
rect 15289 26741 15301 26775
rect 15335 26772 15347 26775
rect 15378 26772 15384 26784
rect 15335 26744 15384 26772
rect 15335 26741 15347 26744
rect 15289 26735 15347 26741
rect 15378 26732 15384 26744
rect 15436 26732 15442 26784
rect 15654 26732 15660 26784
rect 15712 26732 15718 26784
rect 15746 26732 15752 26784
rect 15804 26732 15810 26784
rect 17328 26772 17356 26803
rect 17402 26800 17408 26852
rect 17460 26840 17466 26852
rect 17773 26843 17831 26849
rect 17773 26840 17785 26843
rect 17460 26812 17785 26840
rect 17460 26800 17466 26812
rect 17773 26809 17785 26812
rect 17819 26809 17831 26843
rect 17773 26803 17831 26809
rect 17880 26772 17908 26880
rect 18233 26877 18245 26880
rect 18279 26877 18291 26911
rect 18233 26871 18291 26877
rect 18506 26868 18512 26920
rect 18564 26908 18570 26920
rect 18984 26917 19012 26948
rect 19518 26936 19524 26988
rect 19576 26936 19582 26988
rect 21542 26976 21548 26988
rect 21192 26948 21548 26976
rect 19794 26917 19800 26920
rect 18693 26911 18751 26917
rect 18693 26908 18705 26911
rect 18564 26880 18705 26908
rect 18564 26868 18570 26880
rect 18693 26877 18705 26880
rect 18739 26877 18751 26911
rect 18693 26871 18751 26877
rect 18877 26911 18935 26917
rect 18877 26877 18889 26911
rect 18923 26877 18935 26911
rect 18877 26871 18935 26877
rect 18969 26911 19027 26917
rect 18969 26877 18981 26911
rect 19015 26877 19027 26911
rect 19788 26908 19800 26917
rect 19755 26880 19800 26908
rect 18969 26871 19027 26877
rect 19788 26871 19800 26880
rect 18892 26840 18920 26871
rect 19794 26868 19800 26871
rect 19852 26868 19858 26920
rect 21192 26917 21220 26948
rect 21542 26936 21548 26948
rect 21600 26936 21606 26988
rect 21928 26976 21956 27016
rect 22186 26976 22192 26988
rect 21928 26948 22192 26976
rect 22186 26936 22192 26948
rect 22244 26936 22250 26988
rect 21177 26911 21235 26917
rect 21177 26877 21189 26911
rect 21223 26877 21235 26911
rect 21177 26871 21235 26877
rect 21266 26868 21272 26920
rect 21324 26908 21330 26920
rect 21361 26911 21419 26917
rect 21361 26908 21373 26911
rect 21324 26880 21373 26908
rect 21324 26868 21330 26880
rect 21361 26877 21373 26880
rect 21407 26877 21419 26911
rect 22370 26908 22376 26920
rect 21361 26871 21419 26877
rect 22029 26880 22376 26908
rect 18248 26812 18920 26840
rect 21453 26843 21511 26849
rect 17328 26744 17908 26772
rect 17954 26732 17960 26784
rect 18012 26781 18018 26784
rect 18012 26775 18031 26781
rect 18019 26772 18031 26775
rect 18248 26772 18276 26812
rect 21453 26809 21465 26843
rect 21499 26840 21511 26843
rect 21542 26840 21548 26852
rect 21499 26812 21548 26840
rect 21499 26809 21511 26812
rect 21453 26803 21511 26809
rect 21542 26800 21548 26812
rect 21600 26800 21606 26852
rect 21669 26843 21727 26849
rect 21669 26809 21681 26843
rect 21715 26840 21727 26843
rect 21818 26840 21824 26852
rect 21715 26812 21824 26840
rect 21715 26809 21727 26812
rect 21669 26803 21727 26809
rect 21818 26800 21824 26812
rect 21876 26800 21882 26852
rect 22029 26840 22057 26880
rect 22370 26868 22376 26880
rect 22428 26868 22434 26920
rect 22922 26868 22928 26920
rect 22980 26908 22986 26920
rect 23201 26911 23259 26917
rect 23201 26908 23213 26911
rect 22980 26880 23213 26908
rect 22980 26868 22986 26880
rect 23201 26877 23213 26880
rect 23247 26877 23259 26911
rect 23201 26871 23259 26877
rect 23474 26868 23480 26920
rect 23532 26908 23538 26920
rect 24670 26908 24676 26920
rect 23532 26880 24676 26908
rect 23532 26868 23538 26880
rect 24670 26868 24676 26880
rect 24728 26868 24734 26920
rect 21928 26812 22057 26840
rect 22281 26843 22339 26849
rect 18019 26744 18276 26772
rect 18019 26741 18031 26744
rect 18012 26735 18031 26741
rect 18012 26732 18018 26735
rect 18690 26732 18696 26784
rect 18748 26732 18754 26784
rect 21269 26775 21327 26781
rect 21269 26741 21281 26775
rect 21315 26772 21327 26775
rect 21928 26772 21956 26812
rect 22281 26809 22293 26843
rect 22327 26840 22339 26843
rect 22546 26843 22604 26849
rect 22546 26840 22558 26843
rect 22327 26812 22558 26840
rect 22327 26809 22339 26812
rect 22281 26803 22339 26809
rect 22546 26809 22558 26812
rect 22592 26809 22604 26843
rect 22546 26803 22604 26809
rect 22094 26781 22100 26784
rect 21315 26744 21956 26772
rect 22081 26775 22100 26781
rect 21315 26741 21327 26744
rect 21269 26735 21327 26741
rect 22081 26741 22093 26775
rect 22081 26735 22100 26741
rect 22094 26732 22100 26735
rect 22152 26732 22158 26784
rect 22296 26772 22324 26803
rect 25314 26800 25320 26852
rect 25372 26800 25378 26852
rect 23014 26772 23020 26784
rect 22296 26744 23020 26772
rect 23014 26732 23020 26744
rect 23072 26772 23078 26784
rect 23382 26772 23388 26784
rect 23072 26744 23388 26772
rect 23072 26732 23078 26744
rect 23382 26732 23388 26744
rect 23440 26732 23446 26784
rect 23474 26732 23480 26784
rect 23532 26772 23538 26784
rect 23661 26775 23719 26781
rect 23661 26772 23673 26775
rect 23532 26744 23673 26772
rect 23532 26732 23538 26744
rect 23661 26741 23673 26744
rect 23707 26741 23719 26775
rect 23661 26735 23719 26741
rect 26234 26732 26240 26784
rect 26292 26772 26298 26784
rect 26605 26775 26663 26781
rect 26605 26772 26617 26775
rect 26292 26744 26617 26772
rect 26292 26732 26298 26744
rect 26605 26741 26617 26744
rect 26651 26741 26663 26775
rect 26605 26735 26663 26741
rect 552 26682 27576 26704
rect 552 26630 7114 26682
rect 7166 26630 7178 26682
rect 7230 26630 7242 26682
rect 7294 26630 7306 26682
rect 7358 26630 7370 26682
rect 7422 26630 13830 26682
rect 13882 26630 13894 26682
rect 13946 26630 13958 26682
rect 14010 26630 14022 26682
rect 14074 26630 14086 26682
rect 14138 26630 20546 26682
rect 20598 26630 20610 26682
rect 20662 26630 20674 26682
rect 20726 26630 20738 26682
rect 20790 26630 20802 26682
rect 20854 26630 27262 26682
rect 27314 26630 27326 26682
rect 27378 26630 27390 26682
rect 27442 26630 27454 26682
rect 27506 26630 27518 26682
rect 27570 26630 27576 26682
rect 552 26608 27576 26630
rect 2222 26568 2228 26580
rect 952 26540 2228 26568
rect 952 26441 980 26540
rect 2222 26528 2228 26540
rect 2280 26568 2286 26580
rect 2280 26540 2728 26568
rect 2280 26528 2286 26540
rect 2593 26503 2651 26509
rect 2593 26469 2605 26503
rect 2639 26469 2651 26503
rect 2700 26500 2728 26540
rect 5810 26528 5816 26580
rect 5868 26528 5874 26580
rect 6549 26571 6607 26577
rect 6549 26537 6561 26571
rect 6595 26568 6607 26571
rect 7006 26568 7012 26580
rect 6595 26540 7012 26568
rect 6595 26537 6607 26540
rect 6549 26531 6607 26537
rect 7006 26528 7012 26540
rect 7064 26528 7070 26580
rect 7466 26528 7472 26580
rect 7524 26528 7530 26580
rect 9582 26568 9588 26580
rect 8864 26540 9588 26568
rect 2700 26472 2820 26500
rect 2593 26463 2651 26469
rect 1210 26441 1216 26444
rect 937 26435 995 26441
rect 937 26401 949 26435
rect 983 26401 995 26435
rect 937 26395 995 26401
rect 1204 26395 1216 26441
rect 1210 26392 1216 26395
rect 1268 26392 1274 26444
rect 2608 26432 2636 26463
rect 2682 26432 2688 26444
rect 2608 26404 2688 26432
rect 2682 26392 2688 26404
rect 2740 26392 2746 26444
rect 2314 26256 2320 26308
rect 2372 26256 2378 26308
rect 2406 26188 2412 26240
rect 2464 26188 2470 26240
rect 2590 26188 2596 26240
rect 2648 26188 2654 26240
rect 2792 26228 2820 26472
rect 3053 26435 3111 26441
rect 3053 26432 3065 26435
rect 2976 26404 3065 26432
rect 2976 26308 3004 26404
rect 3053 26401 3065 26404
rect 3099 26401 3111 26435
rect 3053 26395 3111 26401
rect 3237 26435 3295 26441
rect 3237 26401 3249 26435
rect 3283 26432 3295 26435
rect 3326 26432 3332 26444
rect 3283 26404 3332 26432
rect 3283 26401 3295 26404
rect 3237 26395 3295 26401
rect 3326 26392 3332 26404
rect 3384 26392 3390 26444
rect 3510 26392 3516 26444
rect 3568 26432 3574 26444
rect 3789 26435 3847 26441
rect 3789 26432 3801 26435
rect 3568 26404 3801 26432
rect 3568 26392 3574 26404
rect 3789 26401 3801 26404
rect 3835 26401 3847 26435
rect 3789 26395 3847 26401
rect 4982 26392 4988 26444
rect 5040 26392 5046 26444
rect 5077 26435 5135 26441
rect 5077 26401 5089 26435
rect 5123 26401 5135 26435
rect 5077 26395 5135 26401
rect 5261 26435 5319 26441
rect 5261 26401 5273 26435
rect 5307 26432 5319 26435
rect 5537 26435 5595 26441
rect 5537 26432 5549 26435
rect 5307 26404 5549 26432
rect 5307 26401 5319 26404
rect 5261 26395 5319 26401
rect 5537 26401 5549 26404
rect 5583 26432 5595 26435
rect 5828 26432 5856 26528
rect 5583 26404 5856 26432
rect 6273 26435 6331 26441
rect 5583 26401 5595 26404
rect 5537 26395 5595 26401
rect 6273 26401 6285 26435
rect 6319 26432 6331 26435
rect 7098 26432 7104 26444
rect 6319 26404 7104 26432
rect 6319 26401 6331 26404
rect 6273 26395 6331 26401
rect 5092 26308 5120 26395
rect 7098 26392 7104 26404
rect 7156 26392 7162 26444
rect 7484 26441 7512 26528
rect 8864 26500 8892 26540
rect 9582 26528 9588 26540
rect 9640 26568 9646 26580
rect 9674 26568 9680 26580
rect 9640 26540 9680 26568
rect 9640 26528 9646 26540
rect 9674 26528 9680 26540
rect 9732 26528 9738 26580
rect 12066 26528 12072 26580
rect 12124 26528 12130 26580
rect 12621 26571 12679 26577
rect 12621 26537 12633 26571
rect 12667 26568 12679 26571
rect 12894 26568 12900 26580
rect 12667 26540 12900 26568
rect 12667 26537 12679 26540
rect 12621 26531 12679 26537
rect 12894 26528 12900 26540
rect 12952 26528 12958 26580
rect 13538 26528 13544 26580
rect 13596 26528 13602 26580
rect 15746 26528 15752 26580
rect 15804 26528 15810 26580
rect 15838 26528 15844 26580
rect 15896 26528 15902 26580
rect 16761 26571 16819 26577
rect 16761 26537 16773 26571
rect 16807 26537 16819 26571
rect 16761 26531 16819 26537
rect 8220 26472 8892 26500
rect 7193 26435 7251 26441
rect 7193 26401 7205 26435
rect 7239 26432 7251 26435
rect 7285 26435 7343 26441
rect 7285 26432 7297 26435
rect 7239 26404 7297 26432
rect 7239 26401 7251 26404
rect 7193 26395 7251 26401
rect 7285 26401 7297 26404
rect 7331 26401 7343 26435
rect 7285 26395 7343 26401
rect 7469 26435 7527 26441
rect 7469 26401 7481 26435
rect 7515 26401 7527 26435
rect 7469 26395 7527 26401
rect 7558 26392 7564 26444
rect 7616 26392 7622 26444
rect 8220 26441 8248 26472
rect 8205 26435 8263 26441
rect 8205 26401 8217 26435
rect 8251 26401 8263 26435
rect 8205 26395 8263 26401
rect 8297 26435 8355 26441
rect 8297 26401 8309 26435
rect 8343 26401 8355 26435
rect 8297 26395 8355 26401
rect 6089 26367 6147 26373
rect 6089 26333 6101 26367
rect 6135 26364 6147 26367
rect 6178 26364 6184 26376
rect 6135 26336 6184 26364
rect 6135 26333 6147 26336
rect 6089 26327 6147 26333
rect 6178 26324 6184 26336
rect 6236 26324 6242 26376
rect 6917 26367 6975 26373
rect 6917 26364 6929 26367
rect 6380 26336 6929 26364
rect 2958 26256 2964 26308
rect 3016 26256 3022 26308
rect 5074 26256 5080 26308
rect 5132 26256 5138 26308
rect 3142 26228 3148 26240
rect 2792 26200 3148 26228
rect 3142 26188 3148 26200
rect 3200 26188 3206 26240
rect 3418 26188 3424 26240
rect 3476 26188 3482 26240
rect 3602 26188 3608 26240
rect 3660 26188 3666 26240
rect 5442 26188 5448 26240
rect 5500 26188 5506 26240
rect 5626 26188 5632 26240
rect 5684 26228 5690 26240
rect 6380 26228 6408 26336
rect 6917 26333 6929 26336
rect 6963 26333 6975 26367
rect 6917 26327 6975 26333
rect 7006 26324 7012 26376
rect 7064 26324 7070 26376
rect 8312 26364 8340 26395
rect 8386 26392 8392 26444
rect 8444 26392 8450 26444
rect 8864 26441 8892 26472
rect 8941 26503 8999 26509
rect 8941 26469 8953 26503
rect 8987 26500 8999 26503
rect 11146 26500 11152 26512
rect 8987 26472 11152 26500
rect 8987 26469 8999 26472
rect 8941 26463 8999 26469
rect 11146 26460 11152 26472
rect 11204 26460 11210 26512
rect 11330 26460 11336 26512
rect 11388 26500 11394 26512
rect 11609 26503 11667 26509
rect 11609 26500 11621 26503
rect 11388 26472 11621 26500
rect 11388 26460 11394 26472
rect 11609 26469 11621 26472
rect 11655 26500 11667 26503
rect 12084 26500 12112 26528
rect 12250 26500 12256 26512
rect 11655 26472 12256 26500
rect 11655 26469 11667 26472
rect 11609 26463 11667 26469
rect 12250 26460 12256 26472
rect 12308 26500 12314 26512
rect 12989 26503 13047 26509
rect 12989 26500 13001 26503
rect 12308 26472 13001 26500
rect 12308 26460 12314 26472
rect 12989 26469 13001 26472
rect 13035 26500 13047 26503
rect 13078 26500 13084 26512
rect 13035 26472 13084 26500
rect 13035 26469 13047 26472
rect 12989 26463 13047 26469
rect 13078 26460 13084 26472
rect 13136 26460 13142 26512
rect 13556 26500 13584 26528
rect 15654 26500 15660 26512
rect 13188 26472 13584 26500
rect 15488 26472 15660 26500
rect 8573 26435 8631 26441
rect 8573 26401 8585 26435
rect 8619 26401 8631 26435
rect 8573 26395 8631 26401
rect 8849 26435 8907 26441
rect 8849 26401 8861 26435
rect 8895 26401 8907 26435
rect 8849 26395 8907 26401
rect 8478 26364 8484 26376
rect 8312 26336 8484 26364
rect 8478 26324 8484 26336
rect 8536 26324 8542 26376
rect 8588 26364 8616 26395
rect 9030 26392 9036 26444
rect 9088 26392 9094 26444
rect 9217 26435 9275 26441
rect 9217 26401 9229 26435
rect 9263 26432 9275 26435
rect 10045 26435 10103 26441
rect 10045 26432 10057 26435
rect 9263 26404 10057 26432
rect 9263 26401 9275 26404
rect 9217 26395 9275 26401
rect 10045 26401 10057 26404
rect 10091 26401 10103 26435
rect 10045 26395 10103 26401
rect 10134 26392 10140 26444
rect 10192 26432 10198 26444
rect 10597 26435 10655 26441
rect 10597 26432 10609 26435
rect 10192 26404 10609 26432
rect 10192 26392 10198 26404
rect 10597 26401 10609 26404
rect 10643 26401 10655 26435
rect 10597 26395 10655 26401
rect 11422 26392 11428 26444
rect 11480 26392 11486 26444
rect 11517 26435 11575 26441
rect 11517 26401 11529 26435
rect 11563 26432 11575 26435
rect 11698 26432 11704 26444
rect 11563 26404 11704 26432
rect 11563 26401 11575 26404
rect 11517 26395 11575 26401
rect 11698 26392 11704 26404
rect 11756 26392 11762 26444
rect 11793 26435 11851 26441
rect 11793 26401 11805 26435
rect 11839 26432 11851 26435
rect 11885 26435 11943 26441
rect 11885 26432 11897 26435
rect 11839 26404 11897 26432
rect 11839 26401 11851 26404
rect 11793 26395 11851 26401
rect 11885 26401 11897 26404
rect 11931 26401 11943 26435
rect 11885 26395 11943 26401
rect 12066 26392 12072 26444
rect 12124 26432 12130 26444
rect 12618 26432 12624 26444
rect 12124 26404 12624 26432
rect 12124 26392 12130 26404
rect 12618 26392 12624 26404
rect 12676 26432 12682 26444
rect 12805 26435 12863 26441
rect 12805 26432 12817 26435
rect 12676 26404 12817 26432
rect 12676 26392 12682 26404
rect 12805 26401 12817 26404
rect 12851 26401 12863 26435
rect 12805 26395 12863 26401
rect 12894 26392 12900 26444
rect 12952 26392 12958 26444
rect 13188 26441 13216 26472
rect 13173 26435 13231 26441
rect 13173 26401 13185 26435
rect 13219 26401 13231 26435
rect 13173 26395 13231 26401
rect 13357 26435 13415 26441
rect 13357 26401 13369 26435
rect 13403 26432 13415 26435
rect 13446 26432 13452 26444
rect 13403 26404 13452 26432
rect 13403 26401 13415 26404
rect 13357 26395 13415 26401
rect 13446 26392 13452 26404
rect 13504 26392 13510 26444
rect 14274 26392 14280 26444
rect 14332 26432 14338 26444
rect 15488 26441 15516 26472
rect 15654 26460 15660 26472
rect 15712 26460 15718 26512
rect 14369 26435 14427 26441
rect 14369 26432 14381 26435
rect 14332 26404 14381 26432
rect 14332 26392 14338 26404
rect 14369 26401 14381 26404
rect 14415 26401 14427 26435
rect 14369 26395 14427 26401
rect 15473 26435 15531 26441
rect 15473 26401 15485 26435
rect 15519 26401 15531 26435
rect 15473 26395 15531 26401
rect 15562 26392 15568 26444
rect 15620 26392 15626 26444
rect 15764 26441 15792 26528
rect 15856 26441 15884 26528
rect 16776 26444 16804 26531
rect 17494 26528 17500 26580
rect 17552 26528 17558 26580
rect 17983 26571 18041 26577
rect 17983 26537 17995 26571
rect 18029 26568 18041 26571
rect 18690 26568 18696 26580
rect 18029 26540 18696 26568
rect 18029 26537 18041 26540
rect 17983 26531 18041 26537
rect 18690 26528 18696 26540
rect 18748 26528 18754 26580
rect 19518 26528 19524 26580
rect 19576 26528 19582 26580
rect 21266 26528 21272 26580
rect 21324 26568 21330 26580
rect 21726 26568 21732 26580
rect 21324 26540 21732 26568
rect 21324 26528 21330 26540
rect 15749 26435 15807 26441
rect 15749 26401 15761 26435
rect 15795 26401 15807 26435
rect 15749 26395 15807 26401
rect 15841 26435 15899 26441
rect 15841 26401 15853 26435
rect 15887 26401 15899 26435
rect 15841 26395 15899 26401
rect 16758 26392 16764 26444
rect 16816 26432 16822 26444
rect 16945 26435 17003 26441
rect 16945 26432 16957 26435
rect 16816 26404 16957 26432
rect 16816 26392 16822 26404
rect 16945 26401 16957 26404
rect 16991 26401 17003 26435
rect 17512 26432 17540 26528
rect 17773 26503 17831 26509
rect 17773 26469 17785 26503
rect 17819 26469 17831 26503
rect 19536 26500 19564 26528
rect 19536 26472 19840 26500
rect 17773 26463 17831 26469
rect 17589 26435 17647 26441
rect 17589 26432 17601 26435
rect 17512 26404 17601 26432
rect 16945 26395 17003 26401
rect 17589 26401 17601 26404
rect 17635 26401 17647 26435
rect 17589 26395 17647 26401
rect 9309 26367 9367 26373
rect 9309 26364 9321 26367
rect 8588 26336 9321 26364
rect 9309 26333 9321 26336
rect 9355 26333 9367 26367
rect 9309 26327 9367 26333
rect 9858 26324 9864 26376
rect 9916 26324 9922 26376
rect 11440 26364 11468 26392
rect 12084 26364 12112 26392
rect 11440 26336 12112 26364
rect 12526 26324 12532 26376
rect 12584 26364 12590 26376
rect 14292 26364 14320 26392
rect 12584 26336 14320 26364
rect 12584 26324 12590 26336
rect 15930 26324 15936 26376
rect 15988 26364 15994 26376
rect 16301 26367 16359 26373
rect 16301 26364 16313 26367
rect 15988 26336 16313 26364
rect 15988 26324 15994 26336
rect 16301 26333 16313 26336
rect 16347 26333 16359 26367
rect 17402 26364 17408 26376
rect 16301 26327 16359 26333
rect 17144 26336 17408 26364
rect 6457 26299 6515 26305
rect 6457 26265 6469 26299
rect 6503 26296 6515 26299
rect 6503 26268 7328 26296
rect 6503 26265 6515 26268
rect 6457 26259 6515 26265
rect 6932 26240 6960 26268
rect 5684 26200 6408 26228
rect 5684 26188 5690 26200
rect 6914 26188 6920 26240
rect 6972 26188 6978 26240
rect 7300 26237 7328 26268
rect 7742 26256 7748 26308
rect 7800 26256 7806 26308
rect 8386 26256 8392 26308
rect 8444 26296 8450 26308
rect 9030 26296 9036 26308
rect 8444 26268 9036 26296
rect 8444 26256 8450 26268
rect 9030 26256 9036 26268
rect 9088 26256 9094 26308
rect 13909 26299 13967 26305
rect 13909 26265 13921 26299
rect 13955 26296 13967 26299
rect 14182 26296 14188 26308
rect 13955 26268 14188 26296
rect 13955 26265 13967 26268
rect 13909 26259 13967 26265
rect 14182 26256 14188 26268
rect 14240 26256 14246 26308
rect 15286 26256 15292 26308
rect 15344 26256 15350 26308
rect 16574 26256 16580 26308
rect 16632 26256 16638 26308
rect 16666 26256 16672 26308
rect 16724 26296 16730 26308
rect 17144 26305 17172 26336
rect 17402 26324 17408 26336
rect 17460 26364 17466 26376
rect 17788 26364 17816 26463
rect 19812 26444 19840 26472
rect 19518 26392 19524 26444
rect 19576 26441 19582 26444
rect 19576 26395 19588 26441
rect 19576 26392 19582 26395
rect 19794 26392 19800 26444
rect 19852 26392 19858 26444
rect 20901 26435 20959 26441
rect 20901 26401 20913 26435
rect 20947 26432 20959 26435
rect 20947 26404 21312 26432
rect 20947 26401 20959 26404
rect 20901 26395 20959 26401
rect 17460 26336 17816 26364
rect 17460 26324 17466 26336
rect 17129 26299 17187 26305
rect 17129 26296 17141 26299
rect 16724 26268 17141 26296
rect 16724 26256 16730 26268
rect 16868 26240 16896 26268
rect 17129 26265 17141 26268
rect 17175 26265 17187 26299
rect 17129 26259 17187 26265
rect 17497 26299 17555 26305
rect 17497 26265 17509 26299
rect 17543 26296 17555 26299
rect 17586 26296 17592 26308
rect 17543 26268 17592 26296
rect 17543 26265 17555 26268
rect 17497 26259 17555 26265
rect 17586 26256 17592 26268
rect 17644 26256 17650 26308
rect 21284 26305 21312 26404
rect 21269 26299 21327 26305
rect 21269 26265 21281 26299
rect 21315 26265 21327 26299
rect 21269 26259 21327 26265
rect 7285 26231 7343 26237
rect 7285 26197 7297 26231
rect 7331 26197 7343 26231
rect 7285 26191 7343 26197
rect 8018 26188 8024 26240
rect 8076 26188 8082 26240
rect 8665 26231 8723 26237
rect 8665 26197 8677 26231
rect 8711 26228 8723 26231
rect 8754 26228 8760 26240
rect 8711 26200 8760 26228
rect 8711 26197 8723 26200
rect 8665 26191 8723 26197
rect 8754 26188 8760 26200
rect 8812 26188 8818 26240
rect 11238 26188 11244 26240
rect 11296 26188 11302 26240
rect 13633 26231 13691 26237
rect 13633 26197 13645 26231
rect 13679 26228 13691 26231
rect 13722 26228 13728 26240
rect 13679 26200 13728 26228
rect 13679 26197 13691 26200
rect 13633 26191 13691 26197
rect 13722 26188 13728 26200
rect 13780 26188 13786 26240
rect 13814 26188 13820 26240
rect 13872 26188 13878 26240
rect 14277 26231 14335 26237
rect 14277 26197 14289 26231
rect 14323 26228 14335 26231
rect 14550 26228 14556 26240
rect 14323 26200 14556 26228
rect 14323 26197 14335 26200
rect 14277 26191 14335 26197
rect 14550 26188 14556 26200
rect 14608 26188 14614 26240
rect 16850 26188 16856 26240
rect 16908 26188 16914 26240
rect 17954 26188 17960 26240
rect 18012 26188 18018 26240
rect 18138 26188 18144 26240
rect 18196 26188 18202 26240
rect 18414 26188 18420 26240
rect 18472 26188 18478 26240
rect 20714 26188 20720 26240
rect 20772 26188 20778 26240
rect 21376 26228 21404 26540
rect 21726 26528 21732 26540
rect 21784 26568 21790 26580
rect 21821 26571 21879 26577
rect 21821 26568 21833 26571
rect 21784 26540 21833 26568
rect 21784 26528 21790 26540
rect 21821 26537 21833 26540
rect 21867 26537 21879 26571
rect 21821 26531 21879 26537
rect 22462 26528 22468 26580
rect 22520 26528 22526 26580
rect 22833 26571 22891 26577
rect 22833 26537 22845 26571
rect 22879 26568 22891 26571
rect 23293 26571 23351 26577
rect 23293 26568 23305 26571
rect 22879 26540 23305 26568
rect 22879 26537 22891 26540
rect 22833 26531 22891 26537
rect 23293 26537 23305 26540
rect 23339 26537 23351 26571
rect 23293 26531 23351 26537
rect 24302 26528 24308 26580
rect 24360 26528 24366 26580
rect 25501 26571 25559 26577
rect 25501 26537 25513 26571
rect 25547 26568 25559 26571
rect 25547 26540 26280 26568
rect 25547 26537 25559 26540
rect 25501 26531 25559 26537
rect 21437 26503 21495 26509
rect 21437 26469 21449 26503
rect 21483 26500 21495 26503
rect 21542 26500 21548 26512
rect 21483 26472 21548 26500
rect 21483 26469 21495 26472
rect 21437 26463 21495 26469
rect 21542 26460 21548 26472
rect 21600 26460 21606 26512
rect 21637 26503 21695 26509
rect 21637 26469 21649 26503
rect 21683 26500 21695 26503
rect 21683 26472 21864 26500
rect 21683 26469 21695 26472
rect 21637 26463 21695 26469
rect 21729 26435 21787 26441
rect 21729 26432 21741 26435
rect 21468 26404 21741 26432
rect 21468 26376 21496 26404
rect 21729 26401 21741 26404
rect 21775 26401 21787 26435
rect 21836 26432 21864 26472
rect 21910 26460 21916 26512
rect 21968 26460 21974 26512
rect 21836 26404 21956 26432
rect 21729 26395 21787 26401
rect 21450 26324 21456 26376
rect 21508 26324 21514 26376
rect 21928 26364 21956 26404
rect 22002 26392 22008 26444
rect 22060 26392 22066 26444
rect 22373 26435 22431 26441
rect 22373 26401 22385 26435
rect 22419 26432 22431 26435
rect 22480 26432 22508 26528
rect 23937 26503 23995 26509
rect 23937 26469 23949 26503
rect 23983 26500 23995 26503
rect 24394 26500 24400 26512
rect 23983 26472 24400 26500
rect 23983 26469 23995 26472
rect 23937 26463 23995 26469
rect 24394 26460 24400 26472
rect 24452 26460 24458 26512
rect 24946 26460 24952 26512
rect 25004 26500 25010 26512
rect 25317 26503 25375 26509
rect 25317 26500 25329 26503
rect 25004 26472 25329 26500
rect 25004 26460 25010 26472
rect 25317 26469 25329 26472
rect 25363 26469 25375 26503
rect 25745 26503 25803 26509
rect 25745 26500 25757 26503
rect 25317 26463 25375 26469
rect 25424 26472 25757 26500
rect 22419 26404 22508 26432
rect 22419 26401 22431 26404
rect 22373 26395 22431 26401
rect 22830 26392 22836 26444
rect 22888 26432 22894 26444
rect 23385 26435 23443 26441
rect 23385 26432 23397 26435
rect 22888 26404 23397 26432
rect 22888 26392 22894 26404
rect 23385 26401 23397 26404
rect 23431 26401 23443 26435
rect 23385 26395 23443 26401
rect 23474 26392 23480 26444
rect 23532 26392 23538 26444
rect 23753 26435 23811 26441
rect 23753 26432 23765 26435
rect 23584 26404 23765 26432
rect 22646 26364 22652 26376
rect 21928 26336 22652 26364
rect 21928 26240 21956 26336
rect 22646 26324 22652 26336
rect 22704 26324 22710 26376
rect 23584 26364 23612 26404
rect 23753 26401 23765 26404
rect 23799 26401 23811 26435
rect 23753 26395 23811 26401
rect 24029 26435 24087 26441
rect 24029 26401 24041 26435
rect 24075 26401 24087 26435
rect 24029 26395 24087 26401
rect 24121 26435 24179 26441
rect 24121 26401 24133 26435
rect 24167 26432 24179 26435
rect 24302 26432 24308 26444
rect 24167 26404 24308 26432
rect 24167 26401 24179 26404
rect 24121 26395 24179 26401
rect 24044 26364 24072 26395
rect 24302 26392 24308 26404
rect 24360 26392 24366 26444
rect 25130 26392 25136 26444
rect 25188 26392 25194 26444
rect 25222 26392 25228 26444
rect 25280 26432 25286 26444
rect 25424 26432 25452 26472
rect 25745 26469 25757 26472
rect 25791 26469 25803 26503
rect 25745 26463 25803 26469
rect 25958 26460 25964 26512
rect 26016 26460 26022 26512
rect 26252 26441 26280 26540
rect 25280 26404 25452 26432
rect 26237 26435 26295 26441
rect 25280 26392 25286 26404
rect 26237 26401 26249 26435
rect 26283 26401 26295 26435
rect 26237 26395 26295 26401
rect 23124 26336 23612 26364
rect 23676 26336 24072 26364
rect 23124 26308 23152 26336
rect 23106 26256 23112 26308
rect 23164 26256 23170 26308
rect 23566 26256 23572 26308
rect 23624 26296 23630 26308
rect 23676 26305 23704 26336
rect 24854 26324 24860 26376
rect 24912 26364 24918 26376
rect 24949 26367 25007 26373
rect 24949 26364 24961 26367
rect 24912 26336 24961 26364
rect 24912 26324 24918 26336
rect 24949 26333 24961 26336
rect 24995 26364 25007 26367
rect 25148 26364 25176 26392
rect 26142 26364 26148 26376
rect 24995 26336 26148 26364
rect 24995 26333 25007 26336
rect 24949 26327 25007 26333
rect 26142 26324 26148 26336
rect 26200 26324 26206 26376
rect 23661 26299 23719 26305
rect 23661 26296 23673 26299
rect 23624 26268 23673 26296
rect 23624 26256 23630 26268
rect 23661 26265 23673 26268
rect 23707 26265 23719 26299
rect 23661 26259 23719 26265
rect 25240 26268 25728 26296
rect 21453 26231 21511 26237
rect 21453 26228 21465 26231
rect 21376 26200 21465 26228
rect 21453 26197 21465 26200
rect 21499 26197 21511 26231
rect 21453 26191 21511 26197
rect 21910 26188 21916 26240
rect 21968 26188 21974 26240
rect 22278 26188 22284 26240
rect 22336 26228 22342 26240
rect 22465 26231 22523 26237
rect 22465 26228 22477 26231
rect 22336 26200 22477 26228
rect 22336 26188 22342 26200
rect 22465 26197 22477 26200
rect 22511 26197 22523 26231
rect 22465 26191 22523 26197
rect 24578 26188 24584 26240
rect 24636 26228 24642 26240
rect 25240 26228 25268 26268
rect 24636 26200 25268 26228
rect 25317 26231 25375 26237
rect 24636 26188 24642 26200
rect 25317 26197 25329 26231
rect 25363 26228 25375 26231
rect 25406 26228 25412 26240
rect 25363 26200 25412 26228
rect 25363 26197 25375 26200
rect 25317 26191 25375 26197
rect 25406 26188 25412 26200
rect 25464 26188 25470 26240
rect 25498 26188 25504 26240
rect 25556 26228 25562 26240
rect 25593 26231 25651 26237
rect 25593 26228 25605 26231
rect 25556 26200 25605 26228
rect 25556 26188 25562 26200
rect 25593 26197 25605 26200
rect 25639 26197 25651 26231
rect 25700 26228 25728 26268
rect 25777 26231 25835 26237
rect 25777 26228 25789 26231
rect 25700 26200 25789 26228
rect 25593 26191 25651 26197
rect 25777 26197 25789 26200
rect 25823 26197 25835 26231
rect 25777 26191 25835 26197
rect 26050 26188 26056 26240
rect 26108 26188 26114 26240
rect 552 26138 27416 26160
rect 552 26086 3756 26138
rect 3808 26086 3820 26138
rect 3872 26086 3884 26138
rect 3936 26086 3948 26138
rect 4000 26086 4012 26138
rect 4064 26086 10472 26138
rect 10524 26086 10536 26138
rect 10588 26086 10600 26138
rect 10652 26086 10664 26138
rect 10716 26086 10728 26138
rect 10780 26086 17188 26138
rect 17240 26086 17252 26138
rect 17304 26086 17316 26138
rect 17368 26086 17380 26138
rect 17432 26086 17444 26138
rect 17496 26086 23904 26138
rect 23956 26086 23968 26138
rect 24020 26086 24032 26138
rect 24084 26086 24096 26138
rect 24148 26086 24160 26138
rect 24212 26086 27416 26138
rect 552 26064 27416 26086
rect 1210 25984 1216 26036
rect 1268 26024 1274 26036
rect 1397 26027 1455 26033
rect 1397 26024 1409 26027
rect 1268 25996 1409 26024
rect 1268 25984 1274 25996
rect 1397 25993 1409 25996
rect 1443 25993 1455 26027
rect 1397 25987 1455 25993
rect 2406 25984 2412 26036
rect 2464 25984 2470 26036
rect 2869 26027 2927 26033
rect 2869 26024 2881 26027
rect 2516 25996 2881 26024
rect 2424 25888 2452 25984
rect 1596 25860 2452 25888
rect 1596 25829 1624 25860
rect 1581 25823 1639 25829
rect 1581 25789 1593 25823
rect 1627 25789 1639 25823
rect 1581 25783 1639 25789
rect 2314 25780 2320 25832
rect 2372 25780 2378 25832
rect 2406 25780 2412 25832
rect 2464 25780 2470 25832
rect 2332 25752 2360 25780
rect 2516 25752 2544 25996
rect 2869 25993 2881 25996
rect 2915 26024 2927 26027
rect 4522 26024 4528 26036
rect 2915 25996 4528 26024
rect 2915 25993 2927 25996
rect 2869 25987 2927 25993
rect 4522 25984 4528 25996
rect 4580 25984 4586 26036
rect 7098 25984 7104 26036
rect 7156 26024 7162 26036
rect 7285 26027 7343 26033
rect 7285 26024 7297 26027
rect 7156 25996 7297 26024
rect 7156 25984 7162 25996
rect 7285 25993 7297 25996
rect 7331 26024 7343 26027
rect 7929 26027 7987 26033
rect 7929 26024 7941 26027
rect 7331 25996 7941 26024
rect 7331 25993 7343 25996
rect 7285 25987 7343 25993
rect 7929 25993 7941 25996
rect 7975 25993 7987 26027
rect 9858 26024 9864 26036
rect 7929 25987 7987 25993
rect 8588 25996 9864 26024
rect 2593 25959 2651 25965
rect 2593 25925 2605 25959
rect 2639 25956 2651 25959
rect 2958 25956 2964 25968
rect 2639 25928 2964 25956
rect 2639 25925 2651 25928
rect 2593 25919 2651 25925
rect 2958 25916 2964 25928
rect 3016 25916 3022 25968
rect 7006 25916 7012 25968
rect 7064 25956 7070 25968
rect 8481 25959 8539 25965
rect 8481 25956 8493 25959
rect 7064 25928 8493 25956
rect 7064 25916 7070 25928
rect 6288 25860 7512 25888
rect 3142 25780 3148 25832
rect 3200 25820 3206 25832
rect 3237 25823 3295 25829
rect 3237 25820 3249 25823
rect 3200 25792 3249 25820
rect 3200 25780 3206 25792
rect 3237 25789 3249 25792
rect 3283 25820 3295 25823
rect 4985 25823 5043 25829
rect 4985 25820 4997 25823
rect 3283 25792 4997 25820
rect 3283 25789 3295 25792
rect 3237 25783 3295 25789
rect 4985 25789 4997 25792
rect 5031 25789 5043 25823
rect 6288 25820 6316 25860
rect 7484 25829 7512 25860
rect 7576 25829 7604 25928
rect 8481 25925 8493 25928
rect 8527 25925 8539 25959
rect 8481 25919 8539 25925
rect 7650 25848 7656 25900
rect 7708 25888 7714 25900
rect 7745 25891 7803 25897
rect 7745 25888 7757 25891
rect 7708 25860 7757 25888
rect 7708 25848 7714 25860
rect 7745 25857 7757 25860
rect 7791 25857 7803 25891
rect 7745 25851 7803 25857
rect 8588 25829 8616 25996
rect 9858 25984 9864 25996
rect 9916 25984 9922 26036
rect 11517 26027 11575 26033
rect 11517 25993 11529 26027
rect 11563 26024 11575 26027
rect 12526 26024 12532 26036
rect 11563 25996 12532 26024
rect 11563 25993 11575 25996
rect 11517 25987 11575 25993
rect 12526 25984 12532 25996
rect 12584 25984 12590 26036
rect 14921 26027 14979 26033
rect 14921 25993 14933 26027
rect 14967 26024 14979 26027
rect 15562 26024 15568 26036
rect 14967 25996 15568 26024
rect 14967 25993 14979 25996
rect 14921 25987 14979 25993
rect 15562 25984 15568 25996
rect 15620 25984 15626 26036
rect 17954 25984 17960 26036
rect 18012 26024 18018 26036
rect 18233 26027 18291 26033
rect 18233 26024 18245 26027
rect 18012 25996 18245 26024
rect 18012 25984 18018 25996
rect 18233 25993 18245 25996
rect 18279 25993 18291 26027
rect 18233 25987 18291 25993
rect 18417 26027 18475 26033
rect 18417 25993 18429 26027
rect 18463 26024 18475 26027
rect 18506 26024 18512 26036
rect 18463 25996 18512 26024
rect 18463 25993 18475 25996
rect 18417 25987 18475 25993
rect 12989 25959 13047 25965
rect 12989 25925 13001 25959
rect 13035 25956 13047 25959
rect 13170 25956 13176 25968
rect 13035 25928 13176 25956
rect 13035 25925 13047 25928
rect 12989 25919 13047 25925
rect 13170 25916 13176 25928
rect 13228 25956 13234 25968
rect 13722 25956 13728 25968
rect 13228 25928 13728 25956
rect 13228 25916 13234 25928
rect 13722 25916 13728 25928
rect 13780 25916 13786 25968
rect 18432 25956 18460 25987
rect 18506 25984 18512 25996
rect 18564 25984 18570 26036
rect 18877 26027 18935 26033
rect 18877 25993 18889 26027
rect 18923 26024 18935 26027
rect 19518 26024 19524 26036
rect 18923 25996 19524 26024
rect 18923 25993 18935 25996
rect 18877 25987 18935 25993
rect 19518 25984 19524 25996
rect 19576 25984 19582 26036
rect 21542 25984 21548 26036
rect 21600 26024 21606 26036
rect 21729 26027 21787 26033
rect 21729 26024 21741 26027
rect 21600 25996 21741 26024
rect 21600 25984 21606 25996
rect 21729 25993 21741 25996
rect 21775 25993 21787 26027
rect 21729 25987 21787 25993
rect 22278 25984 22284 26036
rect 22336 25984 22342 26036
rect 22462 25984 22468 26036
rect 22520 25984 22526 26036
rect 22830 25984 22836 26036
rect 22888 25984 22894 26036
rect 22922 25984 22928 26036
rect 22980 26024 22986 26036
rect 23109 26027 23167 26033
rect 23109 26024 23121 26027
rect 22980 25996 23121 26024
rect 22980 25984 22986 25996
rect 23109 25993 23121 25996
rect 23155 25993 23167 26027
rect 23109 25987 23167 25993
rect 23477 26027 23535 26033
rect 23477 25993 23489 26027
rect 23523 26024 23535 26027
rect 23566 26024 23572 26036
rect 23523 25996 23572 26024
rect 23523 25993 23535 25996
rect 23477 25987 23535 25993
rect 23566 25984 23572 25996
rect 23624 25984 23630 26036
rect 23937 26027 23995 26033
rect 23937 25993 23949 26027
rect 23983 26024 23995 26027
rect 24302 26024 24308 26036
rect 23983 25996 24308 26024
rect 23983 25993 23995 25996
rect 23937 25987 23995 25993
rect 24302 25984 24308 25996
rect 24360 25984 24366 26036
rect 24581 26027 24639 26033
rect 24581 25993 24593 26027
rect 24627 26024 24639 26027
rect 24946 26024 24952 26036
rect 24627 25996 24952 26024
rect 24627 25993 24639 25996
rect 24581 25987 24639 25993
rect 24946 25984 24952 25996
rect 25004 25984 25010 26036
rect 25406 26024 25412 26036
rect 25056 25996 25412 26024
rect 18064 25928 18460 25956
rect 13265 25891 13323 25897
rect 13265 25857 13277 25891
rect 13311 25888 13323 25891
rect 16577 25891 16635 25897
rect 13311 25860 14780 25888
rect 13311 25857 13323 25860
rect 13265 25851 13323 25857
rect 7009 25823 7067 25829
rect 7009 25820 7021 25823
rect 4985 25783 5043 25789
rect 5644 25792 6316 25820
rect 6380 25792 7021 25820
rect 2332 25724 2544 25752
rect 2685 25755 2743 25761
rect 2685 25721 2697 25755
rect 2731 25752 2743 25755
rect 3326 25752 3332 25764
rect 2731 25724 3332 25752
rect 2731 25721 2743 25724
rect 2685 25715 2743 25721
rect 3326 25712 3332 25724
rect 3384 25712 3390 25764
rect 3504 25755 3562 25761
rect 3504 25721 3516 25755
rect 3550 25752 3562 25755
rect 3602 25752 3608 25764
rect 3550 25724 3608 25752
rect 3550 25721 3562 25724
rect 3504 25715 3562 25721
rect 3602 25712 3608 25724
rect 3660 25712 3666 25764
rect 5258 25761 5264 25764
rect 5252 25715 5264 25761
rect 5258 25712 5264 25715
rect 5316 25712 5322 25764
rect 2498 25644 2504 25696
rect 2556 25684 2562 25696
rect 2866 25684 2872 25696
rect 2924 25693 2930 25696
rect 2924 25687 2943 25693
rect 2556 25656 2872 25684
rect 2556 25644 2562 25656
rect 2866 25644 2872 25656
rect 2931 25684 2943 25687
rect 2931 25656 3017 25684
rect 2931 25653 2943 25656
rect 2924 25647 2943 25653
rect 2924 25644 2930 25647
rect 3050 25644 3056 25696
rect 3108 25644 3114 25696
rect 3344 25684 3372 25712
rect 5644 25696 5672 25792
rect 4617 25687 4675 25693
rect 4617 25684 4629 25687
rect 3344 25656 4629 25684
rect 4617 25653 4629 25656
rect 4663 25684 4675 25687
rect 5626 25684 5632 25696
rect 4663 25656 5632 25684
rect 4663 25653 4675 25656
rect 4617 25647 4675 25653
rect 5626 25644 5632 25656
rect 5684 25644 5690 25696
rect 5718 25644 5724 25696
rect 5776 25684 5782 25696
rect 6178 25684 6184 25696
rect 5776 25656 6184 25684
rect 5776 25644 5782 25656
rect 6178 25644 6184 25656
rect 6236 25684 6242 25696
rect 6380 25693 6408 25792
rect 7009 25789 7021 25792
rect 7055 25820 7067 25823
rect 7193 25823 7251 25829
rect 7193 25820 7205 25823
rect 7055 25792 7205 25820
rect 7055 25789 7067 25792
rect 7009 25783 7067 25789
rect 7193 25789 7205 25792
rect 7239 25789 7251 25823
rect 7193 25783 7251 25789
rect 7469 25823 7527 25829
rect 7469 25789 7481 25823
rect 7515 25789 7527 25823
rect 7469 25783 7527 25789
rect 7561 25823 7619 25829
rect 7561 25789 7573 25823
rect 7607 25789 7619 25823
rect 7561 25783 7619 25789
rect 8021 25823 8079 25829
rect 8021 25789 8033 25823
rect 8067 25789 8079 25823
rect 8021 25783 8079 25789
rect 8573 25823 8631 25829
rect 8573 25789 8585 25823
rect 8619 25789 8631 25823
rect 8573 25783 8631 25789
rect 8665 25823 8723 25829
rect 8665 25789 8677 25823
rect 8711 25820 8723 25823
rect 10137 25823 10195 25829
rect 10137 25820 10149 25823
rect 8711 25792 10149 25820
rect 8711 25789 8723 25792
rect 8665 25783 8723 25789
rect 10137 25789 10149 25792
rect 10183 25820 10195 25823
rect 10962 25820 10968 25832
rect 10183 25792 10968 25820
rect 10183 25789 10195 25792
rect 10137 25783 10195 25789
rect 8036 25752 8064 25783
rect 10962 25780 10968 25792
rect 11020 25820 11026 25832
rect 11609 25823 11667 25829
rect 11609 25820 11621 25823
rect 11020 25792 11621 25820
rect 11020 25780 11026 25792
rect 11609 25789 11621 25792
rect 11655 25789 11667 25823
rect 11609 25783 11667 25789
rect 13173 25823 13231 25829
rect 13173 25789 13185 25823
rect 13219 25789 13231 25823
rect 13173 25783 13231 25789
rect 13357 25823 13415 25829
rect 13357 25789 13369 25823
rect 13403 25820 13415 25823
rect 13630 25820 13636 25832
rect 13403 25792 13636 25820
rect 13403 25789 13415 25792
rect 13357 25783 13415 25789
rect 8036 25724 8708 25752
rect 6365 25687 6423 25693
rect 6365 25684 6377 25687
rect 6236 25656 6377 25684
rect 6236 25644 6242 25656
rect 6365 25653 6377 25656
rect 6411 25653 6423 25687
rect 6365 25647 6423 25653
rect 6454 25644 6460 25696
rect 6512 25644 6518 25696
rect 8680 25684 8708 25724
rect 8754 25712 8760 25764
rect 8812 25752 8818 25764
rect 8910 25755 8968 25761
rect 8910 25752 8922 25755
rect 8812 25724 8922 25752
rect 8812 25712 8818 25724
rect 8910 25721 8922 25724
rect 8956 25721 8968 25755
rect 8910 25715 8968 25721
rect 10404 25755 10462 25761
rect 10404 25721 10416 25755
rect 10450 25752 10462 25755
rect 11238 25752 11244 25764
rect 10450 25724 11244 25752
rect 10450 25721 10462 25724
rect 10404 25715 10462 25721
rect 11238 25712 11244 25724
rect 11296 25712 11302 25764
rect 11882 25761 11888 25764
rect 11876 25715 11888 25761
rect 11882 25712 11888 25715
rect 11940 25712 11946 25764
rect 13188 25752 13216 25783
rect 13630 25780 13636 25792
rect 13688 25780 13694 25832
rect 13722 25780 13728 25832
rect 13780 25820 13786 25832
rect 14093 25823 14151 25829
rect 14093 25820 14105 25823
rect 13780 25792 14105 25820
rect 13780 25780 13786 25792
rect 14093 25789 14105 25792
rect 14139 25789 14151 25823
rect 14093 25783 14151 25789
rect 14182 25780 14188 25832
rect 14240 25780 14246 25832
rect 14366 25780 14372 25832
rect 14424 25780 14430 25832
rect 14752 25829 14780 25860
rect 16577 25857 16589 25891
rect 16623 25888 16635 25891
rect 17034 25888 17040 25900
rect 16623 25860 17040 25888
rect 16623 25857 16635 25860
rect 16577 25851 16635 25857
rect 17034 25848 17040 25860
rect 17092 25848 17098 25900
rect 14645 25823 14703 25829
rect 14645 25820 14657 25823
rect 14476 25792 14657 25820
rect 14200 25752 14228 25780
rect 13188 25724 14228 25752
rect 10045 25687 10103 25693
rect 10045 25684 10057 25687
rect 8680 25656 10057 25684
rect 10045 25653 10057 25656
rect 10091 25684 10103 25687
rect 10134 25684 10140 25696
rect 10091 25656 10140 25684
rect 10091 25653 10103 25656
rect 10045 25647 10103 25653
rect 10134 25644 10140 25656
rect 10192 25644 10198 25696
rect 13538 25644 13544 25696
rect 13596 25644 13602 25696
rect 13814 25644 13820 25696
rect 13872 25684 13878 25696
rect 14476 25684 14504 25792
rect 14645 25789 14657 25792
rect 14691 25789 14703 25823
rect 14645 25783 14703 25789
rect 14737 25823 14795 25829
rect 14737 25789 14749 25823
rect 14783 25789 14795 25823
rect 14737 25783 14795 25789
rect 17862 25780 17868 25832
rect 17920 25780 17926 25832
rect 18064 25829 18092 25928
rect 18414 25848 18420 25900
rect 18472 25888 18478 25900
rect 18472 25860 18552 25888
rect 18472 25848 18478 25860
rect 18049 25823 18107 25829
rect 18049 25789 18061 25823
rect 18095 25789 18107 25823
rect 18049 25783 18107 25789
rect 18138 25780 18144 25832
rect 18196 25780 18202 25832
rect 18524 25829 18552 25860
rect 19794 25848 19800 25900
rect 19852 25888 19858 25900
rect 20257 25891 20315 25897
rect 20257 25888 20269 25891
rect 19852 25860 20269 25888
rect 19852 25848 19858 25860
rect 20257 25857 20269 25860
rect 20303 25857 20315 25891
rect 22296 25888 22324 25984
rect 22848 25888 22876 25984
rect 24486 25916 24492 25968
rect 24544 25956 24550 25968
rect 24762 25956 24768 25968
rect 24544 25928 24768 25956
rect 24544 25916 24550 25928
rect 24762 25916 24768 25928
rect 24820 25916 24826 25968
rect 25056 25956 25084 25996
rect 25406 25984 25412 25996
rect 25464 25984 25470 26036
rect 25685 26027 25743 26033
rect 25685 25993 25697 26027
rect 25731 26024 25743 26027
rect 25958 26024 25964 26036
rect 25731 25996 25964 26024
rect 25731 25993 25743 25996
rect 25685 25987 25743 25993
rect 25958 25984 25964 25996
rect 26016 25984 26022 26036
rect 24964 25928 25084 25956
rect 20257 25851 20315 25857
rect 21836 25860 22140 25888
rect 22296 25860 22416 25888
rect 22848 25860 23428 25888
rect 21836 25832 21864 25860
rect 18509 25823 18567 25829
rect 18509 25789 18521 25823
rect 18555 25789 18567 25823
rect 18509 25783 18567 25789
rect 18693 25823 18751 25829
rect 18693 25789 18705 25823
rect 18739 25789 18751 25823
rect 18693 25783 18751 25789
rect 14553 25755 14611 25761
rect 14553 25721 14565 25755
rect 14599 25752 14611 25755
rect 15838 25752 15844 25764
rect 14599 25724 15844 25752
rect 14599 25721 14611 25724
rect 14553 25715 14611 25721
rect 15838 25712 15844 25724
rect 15896 25712 15902 25764
rect 16298 25712 16304 25764
rect 16356 25761 16362 25764
rect 16356 25715 16368 25761
rect 18156 25752 18184 25780
rect 18708 25752 18736 25783
rect 21818 25780 21824 25832
rect 21876 25780 21882 25832
rect 21913 25823 21971 25829
rect 21913 25789 21925 25823
rect 21959 25820 21971 25823
rect 22002 25820 22008 25832
rect 21959 25792 22008 25820
rect 21959 25789 21971 25792
rect 21913 25783 21971 25789
rect 18156 25724 18736 25752
rect 20524 25755 20582 25761
rect 20524 25721 20536 25755
rect 20570 25752 20582 25755
rect 20714 25752 20720 25764
rect 20570 25724 20720 25752
rect 20570 25721 20582 25724
rect 20524 25715 20582 25721
rect 16356 25712 16362 25715
rect 20714 25712 20720 25724
rect 20772 25712 20778 25764
rect 21928 25752 21956 25783
rect 22002 25780 22008 25792
rect 22060 25780 22066 25832
rect 22112 25829 22140 25860
rect 22097 25823 22155 25829
rect 22097 25789 22109 25823
rect 22143 25789 22155 25823
rect 22097 25783 22155 25789
rect 22189 25823 22247 25829
rect 22189 25789 22201 25823
rect 22235 25820 22247 25823
rect 22278 25820 22284 25832
rect 22235 25792 22284 25820
rect 22235 25789 22247 25792
rect 22189 25783 22247 25789
rect 22278 25780 22284 25792
rect 22336 25780 22342 25832
rect 22388 25829 22416 25860
rect 22373 25823 22431 25829
rect 22373 25789 22385 25823
rect 22419 25789 22431 25823
rect 22373 25783 22431 25789
rect 23014 25780 23020 25832
rect 23072 25780 23078 25832
rect 23400 25820 23428 25860
rect 23474 25848 23480 25900
rect 23532 25888 23538 25900
rect 24964 25888 24992 25928
rect 23532 25860 24072 25888
rect 23532 25848 23538 25860
rect 24044 25829 24072 25860
rect 24504 25860 24992 25888
rect 25041 25891 25099 25897
rect 24504 25829 24532 25860
rect 25041 25857 25053 25891
rect 25087 25888 25099 25891
rect 25087 25860 25452 25888
rect 25087 25857 25099 25860
rect 25041 25851 25099 25857
rect 25424 25832 25452 25860
rect 23845 25823 23903 25829
rect 23845 25820 23857 25823
rect 23400 25792 23857 25820
rect 23845 25789 23857 25792
rect 23891 25789 23903 25823
rect 23845 25783 23903 25789
rect 24029 25823 24087 25829
rect 24029 25789 24041 25823
rect 24075 25789 24087 25823
rect 24029 25783 24087 25789
rect 24489 25823 24547 25829
rect 24489 25789 24501 25823
rect 24535 25789 24547 25823
rect 24489 25783 24547 25789
rect 21652 25724 21956 25752
rect 21652 25696 21680 25724
rect 24504 25696 24532 25783
rect 24578 25780 24584 25832
rect 24636 25820 24642 25832
rect 24765 25823 24823 25829
rect 24765 25820 24777 25823
rect 24636 25792 24777 25820
rect 24636 25780 24642 25792
rect 24765 25789 24777 25792
rect 24811 25789 24823 25823
rect 24765 25783 24823 25789
rect 24949 25823 25007 25829
rect 24949 25789 24961 25823
rect 24995 25820 25007 25823
rect 25222 25820 25228 25832
rect 24995 25792 25228 25820
rect 24995 25789 25007 25792
rect 24949 25783 25007 25789
rect 25222 25780 25228 25792
rect 25280 25780 25286 25832
rect 25406 25780 25412 25832
rect 25464 25780 25470 25832
rect 26234 25780 26240 25832
rect 26292 25820 26298 25832
rect 27065 25823 27123 25829
rect 27065 25820 27077 25823
rect 26292 25792 27077 25820
rect 26292 25780 26298 25792
rect 27065 25789 27077 25792
rect 27111 25789 27123 25823
rect 27065 25783 27123 25789
rect 26786 25712 26792 25764
rect 26844 25761 26850 25764
rect 26844 25715 26856 25761
rect 26844 25712 26850 25715
rect 13872 25656 14504 25684
rect 13872 25644 13878 25656
rect 15194 25644 15200 25696
rect 15252 25644 15258 25696
rect 21634 25644 21640 25696
rect 21692 25644 21698 25696
rect 24302 25644 24308 25696
rect 24360 25644 24366 25696
rect 24486 25644 24492 25696
rect 24544 25644 24550 25696
rect 25409 25687 25467 25693
rect 25409 25653 25421 25687
rect 25455 25684 25467 25687
rect 25498 25684 25504 25696
rect 25455 25656 25504 25684
rect 25455 25653 25467 25656
rect 25409 25647 25467 25653
rect 25498 25644 25504 25656
rect 25556 25644 25562 25696
rect 25590 25644 25596 25696
rect 25648 25644 25654 25696
rect 552 25594 27576 25616
rect 552 25542 7114 25594
rect 7166 25542 7178 25594
rect 7230 25542 7242 25594
rect 7294 25542 7306 25594
rect 7358 25542 7370 25594
rect 7422 25542 13830 25594
rect 13882 25542 13894 25594
rect 13946 25542 13958 25594
rect 14010 25542 14022 25594
rect 14074 25542 14086 25594
rect 14138 25542 20546 25594
rect 20598 25542 20610 25594
rect 20662 25542 20674 25594
rect 20726 25542 20738 25594
rect 20790 25542 20802 25594
rect 20854 25542 27262 25594
rect 27314 25542 27326 25594
rect 27378 25542 27390 25594
rect 27442 25542 27454 25594
rect 27506 25542 27518 25594
rect 27570 25542 27576 25594
rect 552 25520 27576 25542
rect 3050 25440 3056 25492
rect 3108 25440 3114 25492
rect 3418 25440 3424 25492
rect 3476 25440 3482 25492
rect 3510 25440 3516 25492
rect 3568 25480 3574 25492
rect 3789 25483 3847 25489
rect 3789 25480 3801 25483
rect 3568 25452 3801 25480
rect 3568 25440 3574 25452
rect 3789 25449 3801 25452
rect 3835 25449 3847 25483
rect 3789 25443 3847 25449
rect 5169 25483 5227 25489
rect 5169 25449 5181 25483
rect 5215 25480 5227 25483
rect 5258 25480 5264 25492
rect 5215 25452 5264 25480
rect 5215 25449 5227 25452
rect 5169 25443 5227 25449
rect 5258 25440 5264 25452
rect 5316 25440 5322 25492
rect 5442 25440 5448 25492
rect 5500 25440 5506 25492
rect 6454 25440 6460 25492
rect 6512 25440 6518 25492
rect 9309 25483 9367 25489
rect 9309 25449 9321 25483
rect 9355 25480 9367 25483
rect 9858 25480 9864 25492
rect 9355 25452 9864 25480
rect 9355 25449 9367 25452
rect 9309 25443 9367 25449
rect 9858 25440 9864 25452
rect 9916 25440 9922 25492
rect 11793 25483 11851 25489
rect 11793 25449 11805 25483
rect 11839 25480 11851 25483
rect 11882 25480 11888 25492
rect 11839 25452 11888 25480
rect 11839 25449 11851 25452
rect 11793 25443 11851 25449
rect 11882 25440 11888 25452
rect 11940 25440 11946 25492
rect 13538 25480 13544 25492
rect 12360 25452 13544 25480
rect 1210 25304 1216 25356
rect 1268 25304 1274 25356
rect 2222 25304 2228 25356
rect 2280 25304 2286 25356
rect 2406 25304 2412 25356
rect 2464 25304 2470 25356
rect 3068 25344 3096 25440
rect 3436 25412 3464 25440
rect 3605 25415 3663 25421
rect 3605 25412 3617 25415
rect 3436 25384 3617 25412
rect 3605 25381 3617 25384
rect 3651 25381 3663 25415
rect 5460 25412 5488 25440
rect 3605 25375 3663 25381
rect 4724 25384 5488 25412
rect 3237 25347 3295 25353
rect 3237 25344 3249 25347
rect 3068 25316 3249 25344
rect 3237 25313 3249 25316
rect 3283 25313 3295 25347
rect 3237 25307 3295 25313
rect 3252 25276 3280 25307
rect 4430 25304 4436 25356
rect 4488 25344 4494 25356
rect 4724 25353 4752 25384
rect 4525 25347 4583 25353
rect 4525 25344 4537 25347
rect 4488 25316 4537 25344
rect 4488 25304 4494 25316
rect 4525 25313 4537 25316
rect 4571 25313 4583 25347
rect 4525 25307 4583 25313
rect 4709 25347 4767 25353
rect 4709 25313 4721 25347
rect 4755 25313 4767 25347
rect 4709 25307 4767 25313
rect 4801 25347 4859 25353
rect 4801 25313 4813 25347
rect 4847 25313 4859 25347
rect 4801 25307 4859 25313
rect 4893 25347 4951 25353
rect 4893 25313 4905 25347
rect 4939 25344 4951 25347
rect 6472 25344 6500 25440
rect 8018 25372 8024 25424
rect 8076 25412 8082 25424
rect 8174 25415 8232 25421
rect 8174 25412 8186 25415
rect 8076 25384 8186 25412
rect 8076 25372 8082 25384
rect 8174 25381 8186 25384
rect 8220 25381 8232 25415
rect 8174 25375 8232 25381
rect 9950 25372 9956 25424
rect 10008 25412 10014 25424
rect 12069 25415 12127 25421
rect 12069 25412 12081 25415
rect 10008 25384 12081 25412
rect 10008 25372 10014 25384
rect 12069 25381 12081 25384
rect 12115 25381 12127 25415
rect 12069 25375 12127 25381
rect 4939 25316 6500 25344
rect 7009 25347 7067 25353
rect 4939 25313 4951 25316
rect 4893 25307 4951 25313
rect 7009 25313 7021 25347
rect 7055 25344 7067 25347
rect 11977 25347 12035 25353
rect 7055 25316 9076 25344
rect 7055 25313 7067 25316
rect 7009 25307 7067 25313
rect 4816 25276 4844 25307
rect 9048 25288 9076 25316
rect 11977 25313 11989 25347
rect 12023 25313 12035 25347
rect 11977 25307 12035 25313
rect 12161 25347 12219 25353
rect 12161 25313 12173 25347
rect 12207 25344 12219 25347
rect 12250 25344 12256 25356
rect 12207 25316 12256 25344
rect 12207 25313 12219 25316
rect 12161 25307 12219 25313
rect 3252 25248 4844 25276
rect 6822 25236 6828 25288
rect 6880 25276 6886 25288
rect 7929 25279 7987 25285
rect 7929 25276 7941 25279
rect 6880 25248 7941 25276
rect 6880 25236 6886 25248
rect 7929 25245 7941 25248
rect 7975 25245 7987 25279
rect 7929 25239 7987 25245
rect 9030 25236 9036 25288
rect 9088 25276 9094 25288
rect 9953 25279 10011 25285
rect 9953 25276 9965 25279
rect 9088 25248 9965 25276
rect 9088 25236 9094 25248
rect 9953 25245 9965 25248
rect 9999 25245 10011 25279
rect 11992 25276 12020 25307
rect 12250 25304 12256 25316
rect 12308 25304 12314 25356
rect 12360 25353 12388 25452
rect 13538 25440 13544 25452
rect 13596 25440 13602 25492
rect 13630 25440 13636 25492
rect 13688 25480 13694 25492
rect 13909 25483 13967 25489
rect 13909 25480 13921 25483
rect 13688 25452 13921 25480
rect 13688 25440 13694 25452
rect 13909 25449 13921 25452
rect 13955 25449 13967 25483
rect 13909 25443 13967 25449
rect 14001 25483 14059 25489
rect 14001 25449 14013 25483
rect 14047 25480 14059 25483
rect 14182 25480 14188 25492
rect 14047 25452 14188 25480
rect 14047 25449 14059 25452
rect 14001 25443 14059 25449
rect 14182 25440 14188 25452
rect 14240 25440 14246 25492
rect 14826 25440 14832 25492
rect 14884 25480 14890 25492
rect 16850 25480 16856 25492
rect 14884 25452 16856 25480
rect 14884 25440 14890 25452
rect 16850 25440 16856 25452
rect 16908 25440 16914 25492
rect 17954 25440 17960 25492
rect 18012 25440 18018 25492
rect 19702 25440 19708 25492
rect 19760 25440 19766 25492
rect 20070 25440 20076 25492
rect 20128 25480 20134 25492
rect 20530 25480 20536 25492
rect 20128 25452 20536 25480
rect 20128 25440 20134 25452
rect 20530 25440 20536 25452
rect 20588 25480 20594 25492
rect 24305 25483 24363 25489
rect 20588 25452 20852 25480
rect 20588 25440 20594 25452
rect 13722 25372 13728 25424
rect 13780 25372 13786 25424
rect 14918 25372 14924 25424
rect 14976 25372 14982 25424
rect 15381 25415 15439 25421
rect 15381 25381 15393 25415
rect 15427 25381 15439 25415
rect 15381 25375 15439 25381
rect 12345 25347 12403 25353
rect 12345 25313 12357 25347
rect 12391 25313 12403 25347
rect 12345 25307 12403 25313
rect 13170 25304 13176 25356
rect 13228 25304 13234 25356
rect 14090 25304 14096 25356
rect 14148 25304 14154 25356
rect 15396 25344 15424 25375
rect 15470 25372 15476 25424
rect 15528 25412 15534 25424
rect 15581 25415 15639 25421
rect 15581 25412 15593 25415
rect 15528 25384 15593 25412
rect 15528 25372 15534 25384
rect 15581 25381 15593 25384
rect 15627 25381 15639 25415
rect 16868 25412 16896 25440
rect 16868 25384 17908 25412
rect 15581 25375 15639 25381
rect 16390 25344 16396 25356
rect 15396 25316 16396 25344
rect 16390 25304 16396 25316
rect 16448 25304 16454 25356
rect 16669 25347 16727 25353
rect 16669 25313 16681 25347
rect 16715 25313 16727 25347
rect 16669 25307 16727 25313
rect 16853 25347 16911 25353
rect 16853 25313 16865 25347
rect 16899 25344 16911 25347
rect 17034 25344 17040 25356
rect 16899 25316 17040 25344
rect 16899 25313 16911 25316
rect 16853 25307 16911 25313
rect 14277 25279 14335 25285
rect 11992 25248 12112 25276
rect 9953 25239 10011 25245
rect 12084 25152 12112 25248
rect 14277 25245 14289 25279
rect 14323 25276 14335 25279
rect 14366 25276 14372 25288
rect 14323 25248 14372 25276
rect 14323 25245 14335 25248
rect 14277 25239 14335 25245
rect 14366 25236 14372 25248
rect 14424 25276 14430 25288
rect 16684 25276 16712 25307
rect 17034 25304 17040 25316
rect 17092 25344 17098 25356
rect 17770 25344 17776 25356
rect 17092 25316 17776 25344
rect 17092 25304 17098 25316
rect 17770 25304 17776 25316
rect 17828 25304 17834 25356
rect 16942 25276 16948 25288
rect 14424 25248 15424 25276
rect 16684 25248 16948 25276
rect 14424 25236 14430 25248
rect 13814 25168 13820 25220
rect 13872 25208 13878 25220
rect 14553 25211 14611 25217
rect 13872 25180 14504 25208
rect 13872 25168 13878 25180
rect 1029 25143 1087 25149
rect 1029 25109 1041 25143
rect 1075 25140 1087 25143
rect 1118 25140 1124 25152
rect 1075 25112 1124 25140
rect 1075 25109 1087 25112
rect 1029 25103 1087 25109
rect 1118 25100 1124 25112
rect 1176 25100 1182 25152
rect 2590 25100 2596 25152
rect 2648 25100 2654 25152
rect 3605 25143 3663 25149
rect 3605 25109 3617 25143
rect 3651 25140 3663 25143
rect 4430 25140 4436 25152
rect 3651 25112 4436 25140
rect 3651 25109 3663 25112
rect 3605 25103 3663 25109
rect 4430 25100 4436 25112
rect 4488 25100 4494 25152
rect 6914 25100 6920 25152
rect 6972 25100 6978 25152
rect 9398 25100 9404 25152
rect 9456 25100 9462 25152
rect 10134 25100 10140 25152
rect 10192 25140 10198 25152
rect 11054 25140 11060 25152
rect 10192 25112 11060 25140
rect 10192 25100 10198 25112
rect 11054 25100 11060 25112
rect 11112 25100 11118 25152
rect 12066 25100 12072 25152
rect 12124 25100 12130 25152
rect 13446 25100 13452 25152
rect 13504 25140 13510 25152
rect 13722 25140 13728 25152
rect 13504 25112 13728 25140
rect 13504 25100 13510 25112
rect 13722 25100 13728 25112
rect 13780 25140 13786 25152
rect 13998 25140 14004 25152
rect 13780 25112 14004 25140
rect 13780 25100 13786 25112
rect 13998 25100 14004 25112
rect 14056 25100 14062 25152
rect 14476 25140 14504 25180
rect 14553 25177 14565 25211
rect 14599 25208 14611 25211
rect 14642 25208 14648 25220
rect 14599 25180 14648 25208
rect 14599 25177 14611 25180
rect 14553 25171 14611 25177
rect 14642 25168 14648 25180
rect 14700 25208 14706 25220
rect 15010 25208 15016 25220
rect 14700 25180 15016 25208
rect 14700 25168 14706 25180
rect 15010 25168 15016 25180
rect 15068 25168 15074 25220
rect 15396 25152 15424 25248
rect 16942 25236 16948 25248
rect 17000 25236 17006 25288
rect 17880 25276 17908 25384
rect 17972 25344 18000 25440
rect 18322 25372 18328 25424
rect 18380 25412 18386 25424
rect 19153 25415 19211 25421
rect 19153 25412 19165 25415
rect 18380 25384 19165 25412
rect 18380 25372 18386 25384
rect 19153 25381 19165 25384
rect 19199 25381 19211 25415
rect 19720 25412 19748 25440
rect 20346 25412 20352 25424
rect 19720 25384 20352 25412
rect 19153 25375 19211 25381
rect 20346 25372 20352 25384
rect 20404 25412 20410 25424
rect 20824 25421 20852 25452
rect 24305 25449 24317 25483
rect 24351 25480 24363 25483
rect 24486 25480 24492 25492
rect 24351 25452 24492 25480
rect 24351 25449 24363 25452
rect 24305 25443 24363 25449
rect 24486 25440 24492 25452
rect 24544 25440 24550 25492
rect 24578 25440 24584 25492
rect 24636 25480 24642 25492
rect 24857 25483 24915 25489
rect 24857 25480 24869 25483
rect 24636 25452 24869 25480
rect 24636 25440 24642 25452
rect 24857 25449 24869 25452
rect 24903 25449 24915 25483
rect 24857 25443 24915 25449
rect 25590 25440 25596 25492
rect 25648 25480 25654 25492
rect 25648 25452 26740 25480
rect 25648 25440 25654 25452
rect 20809 25415 20867 25421
rect 20404 25384 20668 25412
rect 20404 25372 20410 25384
rect 18417 25347 18475 25353
rect 18417 25344 18429 25347
rect 17972 25316 18429 25344
rect 18417 25313 18429 25316
rect 18463 25313 18475 25347
rect 18417 25307 18475 25313
rect 19245 25347 19303 25353
rect 19245 25313 19257 25347
rect 19291 25344 19303 25347
rect 19705 25347 19763 25353
rect 19705 25344 19717 25347
rect 19291 25316 19717 25344
rect 19291 25313 19303 25316
rect 19245 25307 19303 25313
rect 19705 25313 19717 25316
rect 19751 25313 19763 25347
rect 19705 25307 19763 25313
rect 20070 25304 20076 25356
rect 20128 25344 20134 25356
rect 20640 25353 20668 25384
rect 20809 25381 20821 25415
rect 20855 25381 20867 25415
rect 26050 25412 26056 25424
rect 20809 25375 20867 25381
rect 25976 25384 26056 25412
rect 20257 25347 20315 25353
rect 20257 25344 20269 25347
rect 20128 25316 20269 25344
rect 20128 25304 20134 25316
rect 20257 25313 20269 25316
rect 20303 25313 20315 25347
rect 20257 25307 20315 25313
rect 20625 25347 20683 25353
rect 20625 25313 20637 25347
rect 20671 25313 20683 25347
rect 20625 25307 20683 25313
rect 20717 25347 20775 25353
rect 20717 25313 20729 25347
rect 20763 25344 20775 25347
rect 20898 25344 20904 25356
rect 20763 25316 20904 25344
rect 20763 25313 20775 25316
rect 20717 25307 20775 25313
rect 20898 25304 20904 25316
rect 20956 25304 20962 25356
rect 25976 25353 26004 25384
rect 26050 25372 26056 25384
rect 26108 25372 26114 25424
rect 26142 25372 26148 25424
rect 26200 25412 26206 25424
rect 26421 25415 26479 25421
rect 26421 25412 26433 25415
rect 26200 25384 26433 25412
rect 26200 25372 26206 25384
rect 26421 25381 26433 25384
rect 26467 25381 26479 25415
rect 26421 25375 26479 25381
rect 20993 25347 21051 25353
rect 20993 25313 21005 25347
rect 21039 25344 21051 25347
rect 21269 25347 21327 25353
rect 21269 25344 21281 25347
rect 21039 25316 21281 25344
rect 21039 25313 21051 25316
rect 20993 25307 21051 25313
rect 21269 25313 21281 25316
rect 21315 25313 21327 25347
rect 21269 25307 21327 25313
rect 25970 25347 26028 25353
rect 25970 25313 25982 25347
rect 26016 25313 26028 25347
rect 25970 25307 26028 25313
rect 26234 25304 26240 25356
rect 26292 25304 26298 25356
rect 26326 25304 26332 25356
rect 26384 25344 26390 25356
rect 26605 25347 26663 25353
rect 26605 25344 26617 25347
rect 26384 25316 26617 25344
rect 26384 25304 26390 25316
rect 26605 25313 26617 25316
rect 26651 25313 26663 25347
rect 26712 25344 26740 25452
rect 26786 25440 26792 25492
rect 26844 25480 26850 25492
rect 26881 25483 26939 25489
rect 26881 25480 26893 25483
rect 26844 25452 26893 25480
rect 26844 25440 26850 25452
rect 26881 25449 26893 25452
rect 26927 25449 26939 25483
rect 26881 25443 26939 25449
rect 27065 25347 27123 25353
rect 27065 25344 27077 25347
rect 26712 25316 27077 25344
rect 26605 25307 26663 25313
rect 27065 25313 27077 25316
rect 27111 25313 27123 25347
rect 27065 25307 27123 25313
rect 17957 25279 18015 25285
rect 17957 25276 17969 25279
rect 17880 25248 17969 25276
rect 17957 25245 17969 25248
rect 18003 25245 18015 25279
rect 17957 25239 18015 25245
rect 21913 25279 21971 25285
rect 21913 25245 21925 25279
rect 21959 25276 21971 25279
rect 22002 25276 22008 25288
rect 21959 25248 22008 25276
rect 21959 25245 21971 25248
rect 21913 25239 21971 25245
rect 22002 25236 22008 25248
rect 22060 25236 22066 25288
rect 22554 25236 22560 25288
rect 22612 25236 22618 25288
rect 23750 25236 23756 25288
rect 23808 25276 23814 25288
rect 23845 25279 23903 25285
rect 23845 25276 23857 25279
rect 23808 25248 23857 25276
rect 23808 25236 23814 25248
rect 23845 25245 23857 25248
rect 23891 25245 23903 25279
rect 23845 25239 23903 25245
rect 22922 25168 22928 25220
rect 22980 25168 22986 25220
rect 24213 25211 24271 25217
rect 24213 25177 24225 25211
rect 24259 25208 24271 25211
rect 24670 25208 24676 25220
rect 24259 25180 24676 25208
rect 24259 25177 24271 25180
rect 24213 25171 24271 25177
rect 24670 25168 24676 25180
rect 24728 25168 24734 25220
rect 14826 25140 14832 25152
rect 14476 25112 14832 25140
rect 14826 25100 14832 25112
rect 14884 25140 14890 25152
rect 14921 25143 14979 25149
rect 14921 25140 14933 25143
rect 14884 25112 14933 25140
rect 14884 25100 14890 25112
rect 14921 25109 14933 25112
rect 14967 25109 14979 25143
rect 14921 25103 14979 25109
rect 15105 25143 15163 25149
rect 15105 25109 15117 25143
rect 15151 25140 15163 25143
rect 15194 25140 15200 25152
rect 15151 25112 15200 25140
rect 15151 25109 15163 25112
rect 15105 25103 15163 25109
rect 15194 25100 15200 25112
rect 15252 25100 15258 25152
rect 15378 25100 15384 25152
rect 15436 25100 15442 25152
rect 15565 25143 15623 25149
rect 15565 25109 15577 25143
rect 15611 25140 15623 25143
rect 15654 25140 15660 25152
rect 15611 25112 15660 25140
rect 15611 25109 15623 25112
rect 15565 25103 15623 25109
rect 15654 25100 15660 25112
rect 15712 25100 15718 25152
rect 15746 25100 15752 25152
rect 15804 25100 15810 25152
rect 16666 25100 16672 25152
rect 16724 25100 16730 25152
rect 18138 25100 18144 25152
rect 18196 25100 18202 25152
rect 20438 25100 20444 25152
rect 20496 25100 20502 25152
rect 23014 25100 23020 25152
rect 23072 25100 23078 25152
rect 25498 25100 25504 25152
rect 25556 25140 25562 25152
rect 26789 25143 26847 25149
rect 26789 25140 26801 25143
rect 25556 25112 26801 25140
rect 25556 25100 25562 25112
rect 26789 25109 26801 25112
rect 26835 25109 26847 25143
rect 26789 25103 26847 25109
rect 552 25050 27416 25072
rect 552 24998 3756 25050
rect 3808 24998 3820 25050
rect 3872 24998 3884 25050
rect 3936 24998 3948 25050
rect 4000 24998 4012 25050
rect 4064 24998 10472 25050
rect 10524 24998 10536 25050
rect 10588 24998 10600 25050
rect 10652 24998 10664 25050
rect 10716 24998 10728 25050
rect 10780 24998 17188 25050
rect 17240 24998 17252 25050
rect 17304 24998 17316 25050
rect 17368 24998 17380 25050
rect 17432 24998 17444 25050
rect 17496 24998 23904 25050
rect 23956 24998 23968 25050
rect 24020 24998 24032 25050
rect 24084 24998 24096 25050
rect 24148 24998 24160 25050
rect 24212 24998 27416 25050
rect 552 24976 27416 24998
rect 2225 24939 2283 24945
rect 2225 24905 2237 24939
rect 2271 24936 2283 24939
rect 2406 24936 2412 24948
rect 2271 24908 2412 24936
rect 2271 24905 2283 24908
rect 2225 24899 2283 24905
rect 2406 24896 2412 24908
rect 2464 24896 2470 24948
rect 2501 24939 2559 24945
rect 2501 24905 2513 24939
rect 2547 24936 2559 24939
rect 2590 24936 2596 24948
rect 2547 24908 2596 24936
rect 2547 24905 2559 24908
rect 2501 24899 2559 24905
rect 2590 24896 2596 24908
rect 2648 24896 2654 24948
rect 3050 24896 3056 24948
rect 3108 24936 3114 24948
rect 3421 24939 3479 24945
rect 3421 24936 3433 24939
rect 3108 24908 3433 24936
rect 3108 24896 3114 24908
rect 3421 24905 3433 24908
rect 3467 24936 3479 24939
rect 4798 24936 4804 24948
rect 3467 24908 4804 24936
rect 3467 24905 3479 24908
rect 3421 24899 3479 24905
rect 4798 24896 4804 24908
rect 4856 24896 4862 24948
rect 6365 24939 6423 24945
rect 6365 24905 6377 24939
rect 6411 24936 6423 24939
rect 6914 24936 6920 24948
rect 6411 24908 6920 24936
rect 6411 24905 6423 24908
rect 6365 24899 6423 24905
rect 6914 24896 6920 24908
rect 6972 24896 6978 24948
rect 7285 24939 7343 24945
rect 7285 24905 7297 24939
rect 7331 24936 7343 24939
rect 8389 24939 8447 24945
rect 8389 24936 8401 24939
rect 7331 24908 8401 24936
rect 7331 24905 7343 24908
rect 7285 24899 7343 24905
rect 8389 24905 8401 24908
rect 8435 24936 8447 24939
rect 9030 24936 9036 24948
rect 8435 24908 9036 24936
rect 8435 24905 8447 24908
rect 8389 24899 8447 24905
rect 9030 24896 9036 24908
rect 9088 24896 9094 24948
rect 10962 24896 10968 24948
rect 11020 24896 11026 24948
rect 14001 24939 14059 24945
rect 14001 24905 14013 24939
rect 14047 24905 14059 24939
rect 14001 24899 14059 24905
rect 2317 24871 2375 24877
rect 2317 24837 2329 24871
rect 2363 24837 2375 24871
rect 2317 24831 2375 24837
rect 2332 24800 2360 24831
rect 1872 24772 2360 24800
rect 2424 24800 2452 24896
rect 2866 24828 2872 24880
rect 2924 24868 2930 24880
rect 3237 24871 3295 24877
rect 3237 24868 3249 24871
rect 2924 24840 3249 24868
rect 2924 24828 2930 24840
rect 3237 24837 3249 24840
rect 3283 24837 3295 24871
rect 3237 24831 3295 24837
rect 4522 24828 4528 24880
rect 4580 24868 4586 24880
rect 4580 24840 5304 24868
rect 4580 24828 4586 24840
rect 2424 24772 3648 24800
rect 845 24735 903 24741
rect 845 24701 857 24735
rect 891 24701 903 24735
rect 1872 24732 1900 24772
rect 3418 24732 3424 24744
rect 845 24695 903 24701
rect 1228 24704 1900 24732
rect 2332 24704 3424 24732
rect 860 24596 888 24695
rect 1228 24676 1256 24704
rect 1118 24673 1124 24676
rect 1112 24664 1124 24673
rect 1079 24636 1124 24664
rect 1112 24627 1124 24636
rect 1118 24624 1124 24627
rect 1176 24624 1182 24676
rect 1210 24624 1216 24676
rect 1268 24624 1274 24676
rect 1854 24624 1860 24676
rect 1912 24664 1918 24676
rect 2332 24664 2360 24704
rect 3375 24701 3424 24704
rect 3142 24664 3148 24676
rect 1912 24636 2360 24664
rect 2424 24636 3148 24664
rect 1912 24624 1918 24636
rect 2424 24596 2452 24636
rect 3142 24624 3148 24636
rect 3200 24624 3206 24676
rect 3375 24667 3387 24701
rect 3421 24692 3424 24701
rect 3476 24692 3482 24744
rect 3620 24732 3648 24772
rect 5074 24760 5080 24812
rect 5132 24800 5138 24812
rect 5169 24803 5227 24809
rect 5169 24800 5181 24803
rect 5132 24772 5181 24800
rect 5132 24760 5138 24772
rect 5169 24769 5181 24772
rect 5215 24769 5227 24803
rect 5276 24800 5304 24840
rect 5718 24828 5724 24880
rect 5776 24828 5782 24880
rect 6454 24828 6460 24880
rect 6512 24868 6518 24880
rect 10980 24868 11008 24896
rect 14016 24868 14044 24899
rect 14090 24896 14096 24948
rect 14148 24936 14154 24948
rect 14369 24939 14427 24945
rect 14369 24936 14381 24939
rect 14148 24908 14381 24936
rect 14148 24896 14154 24908
rect 14369 24905 14381 24908
rect 14415 24905 14427 24939
rect 14369 24899 14427 24905
rect 14918 24896 14924 24948
rect 14976 24896 14982 24948
rect 15010 24896 15016 24948
rect 15068 24896 15074 24948
rect 15197 24939 15255 24945
rect 15197 24905 15209 24939
rect 15243 24936 15255 24939
rect 15562 24936 15568 24948
rect 15243 24908 15568 24936
rect 15243 24905 15255 24908
rect 15197 24899 15255 24905
rect 15562 24896 15568 24908
rect 15620 24896 15626 24948
rect 15746 24896 15752 24948
rect 15804 24936 15810 24948
rect 16209 24939 16267 24945
rect 16209 24936 16221 24939
rect 15804 24908 16221 24936
rect 15804 24896 15810 24908
rect 16209 24905 16221 24908
rect 16255 24905 16267 24939
rect 16209 24899 16267 24905
rect 16298 24896 16304 24948
rect 16356 24896 16362 24948
rect 16390 24896 16396 24948
rect 16448 24896 16454 24948
rect 21450 24936 21456 24948
rect 16500 24908 21456 24936
rect 14274 24868 14280 24880
rect 6512 24840 7144 24868
rect 10980 24840 11744 24868
rect 14016 24840 14280 24868
rect 6512 24828 6518 24840
rect 6273 24803 6331 24809
rect 6273 24800 6285 24803
rect 5276 24772 6285 24800
rect 5169 24763 5227 24769
rect 6273 24769 6285 24772
rect 6319 24800 6331 24803
rect 6319 24772 7052 24800
rect 6319 24769 6331 24772
rect 6273 24763 6331 24769
rect 4709 24735 4767 24741
rect 4709 24732 4721 24735
rect 3620 24704 4721 24732
rect 3421 24670 3438 24692
rect 3620 24673 3648 24704
rect 4709 24701 4721 24704
rect 4755 24732 4767 24735
rect 5813 24735 5871 24741
rect 5813 24732 5825 24735
rect 4755 24704 5825 24732
rect 4755 24701 4767 24704
rect 4709 24695 4767 24701
rect 5813 24701 5825 24704
rect 5859 24701 5871 24735
rect 5813 24695 5871 24701
rect 6792 24735 6850 24741
rect 6792 24701 6804 24735
rect 6838 24732 6850 24735
rect 6914 24732 6920 24744
rect 6838 24704 6920 24732
rect 6838 24701 6850 24704
rect 6792 24695 6850 24701
rect 6914 24692 6920 24704
rect 6972 24692 6978 24744
rect 7024 24741 7052 24772
rect 7009 24735 7067 24741
rect 7009 24701 7021 24735
rect 7055 24701 7067 24735
rect 7009 24695 7067 24701
rect 7116 24732 7144 24840
rect 11716 24809 11744 24840
rect 14274 24828 14280 24840
rect 14332 24828 14338 24880
rect 14458 24828 14464 24880
rect 14516 24868 14522 24880
rect 14826 24868 14832 24880
rect 14516 24840 14832 24868
rect 14516 24828 14522 24840
rect 14826 24828 14832 24840
rect 14884 24828 14890 24880
rect 9769 24803 9827 24809
rect 9769 24769 9781 24803
rect 9815 24800 9827 24803
rect 11701 24803 11759 24809
rect 9815 24772 11100 24800
rect 9815 24769 9827 24772
rect 9769 24763 9827 24769
rect 11072 24744 11100 24772
rect 11701 24769 11713 24803
rect 11747 24769 11759 24803
rect 11701 24763 11759 24769
rect 13446 24760 13452 24812
rect 13504 24800 13510 24812
rect 13814 24800 13820 24812
rect 13504 24772 13820 24800
rect 13504 24760 13510 24772
rect 13814 24760 13820 24772
rect 13872 24760 13878 24812
rect 14182 24800 14188 24812
rect 13924 24772 14188 24800
rect 7558 24732 7564 24744
rect 7116 24704 7564 24732
rect 3421 24667 3433 24670
rect 3375 24661 3433 24667
rect 3605 24667 3663 24673
rect 3605 24633 3617 24667
rect 3651 24633 3663 24667
rect 3605 24627 3663 24633
rect 5077 24667 5135 24673
rect 5077 24633 5089 24667
rect 5123 24664 5135 24667
rect 5353 24667 5411 24673
rect 5353 24664 5365 24667
rect 5123 24636 5365 24664
rect 5123 24633 5135 24636
rect 5077 24627 5135 24633
rect 5353 24633 5365 24636
rect 5399 24633 5411 24667
rect 5353 24627 5411 24633
rect 5537 24667 5595 24673
rect 5537 24633 5549 24667
rect 5583 24664 5595 24667
rect 5626 24664 5632 24676
rect 5583 24636 5632 24664
rect 5583 24633 5595 24636
rect 5537 24627 5595 24633
rect 5626 24624 5632 24636
rect 5684 24624 5690 24676
rect 860 24568 2452 24596
rect 2501 24599 2559 24605
rect 2501 24565 2513 24599
rect 2547 24596 2559 24599
rect 2682 24596 2688 24608
rect 2547 24568 2688 24596
rect 2547 24565 2559 24568
rect 2501 24559 2559 24565
rect 2682 24556 2688 24568
rect 2740 24556 2746 24608
rect 4798 24556 4804 24608
rect 4856 24556 4862 24608
rect 4890 24556 4896 24608
rect 4948 24556 4954 24608
rect 5442 24556 5448 24608
rect 5500 24556 5506 24608
rect 5905 24599 5963 24605
rect 5905 24565 5917 24599
rect 5951 24596 5963 24599
rect 6733 24599 6791 24605
rect 6733 24596 6745 24599
rect 5951 24568 6745 24596
rect 5951 24565 5963 24568
rect 5905 24559 5963 24565
rect 6733 24565 6745 24568
rect 6779 24596 6791 24599
rect 6822 24596 6828 24608
rect 6779 24568 6828 24596
rect 6779 24565 6791 24568
rect 6733 24559 6791 24565
rect 6822 24556 6828 24568
rect 6880 24556 6886 24608
rect 6917 24599 6975 24605
rect 6917 24565 6929 24599
rect 6963 24596 6975 24599
rect 7116 24596 7144 24704
rect 7558 24692 7564 24704
rect 7616 24692 7622 24744
rect 7745 24735 7803 24741
rect 7745 24701 7757 24735
rect 7791 24732 7803 24735
rect 7834 24732 7840 24744
rect 7791 24704 7840 24732
rect 7791 24701 7803 24704
rect 7745 24695 7803 24701
rect 7834 24692 7840 24704
rect 7892 24692 7898 24744
rect 10042 24732 10048 24744
rect 9784 24704 10048 24732
rect 7650 24624 7656 24676
rect 7708 24624 7714 24676
rect 8662 24624 8668 24676
rect 8720 24664 8726 24676
rect 9502 24667 9560 24673
rect 9502 24664 9514 24667
rect 8720 24636 9514 24664
rect 8720 24624 8726 24636
rect 9502 24633 9514 24636
rect 9548 24633 9560 24667
rect 9502 24627 9560 24633
rect 6963 24568 7144 24596
rect 6963 24565 6975 24568
rect 6917 24559 6975 24565
rect 7466 24556 7472 24608
rect 7524 24556 7530 24608
rect 8846 24556 8852 24608
rect 8904 24596 8910 24608
rect 9784 24596 9812 24704
rect 10042 24692 10048 24704
rect 10100 24692 10106 24744
rect 10134 24692 10140 24744
rect 10192 24692 10198 24744
rect 10410 24692 10416 24744
rect 10468 24692 10474 24744
rect 10505 24735 10563 24741
rect 10505 24701 10517 24735
rect 10551 24701 10563 24735
rect 10505 24695 10563 24701
rect 10226 24624 10232 24676
rect 10284 24624 10290 24676
rect 10318 24624 10324 24676
rect 10376 24664 10382 24676
rect 10520 24664 10548 24695
rect 11054 24692 11060 24744
rect 11112 24692 11118 24744
rect 13924 24741 13952 24772
rect 14182 24760 14188 24772
rect 14240 24800 14246 24812
rect 14550 24800 14556 24812
rect 14240 24772 14556 24800
rect 14240 24760 14246 24772
rect 14550 24760 14556 24772
rect 14608 24760 14614 24812
rect 15102 24800 15108 24812
rect 14752 24772 15108 24800
rect 13909 24735 13967 24741
rect 13909 24701 13921 24735
rect 13955 24701 13967 24735
rect 13909 24695 13967 24701
rect 10376 24636 10548 24664
rect 11968 24667 12026 24673
rect 10376 24624 10382 24636
rect 11968 24633 11980 24667
rect 12014 24664 12026 24667
rect 12894 24664 12900 24676
rect 12014 24636 12900 24664
rect 12014 24633 12026 24636
rect 11968 24627 12026 24633
rect 12894 24624 12900 24636
rect 12952 24624 12958 24676
rect 8904 24568 9812 24596
rect 8904 24556 8910 24568
rect 9858 24556 9864 24608
rect 9916 24556 9922 24608
rect 11149 24599 11207 24605
rect 11149 24565 11161 24599
rect 11195 24596 11207 24599
rect 11790 24596 11796 24608
rect 11195 24568 11796 24596
rect 11195 24565 11207 24568
rect 11149 24559 11207 24565
rect 11790 24556 11796 24568
rect 11848 24556 11854 24608
rect 13078 24556 13084 24608
rect 13136 24596 13142 24608
rect 13924 24596 13952 24695
rect 13998 24692 14004 24744
rect 14056 24732 14062 24744
rect 14752 24741 14780 24772
rect 15102 24760 15108 24772
rect 15160 24760 15166 24812
rect 15194 24760 15200 24812
rect 15252 24760 15258 24812
rect 14737 24735 14795 24741
rect 14737 24732 14749 24735
rect 14056 24704 14749 24732
rect 14056 24692 14062 24704
rect 14737 24701 14749 24704
rect 14783 24701 14795 24735
rect 15212 24732 15240 24760
rect 15473 24735 15531 24741
rect 15473 24732 15485 24735
rect 15212 24704 15485 24732
rect 14737 24695 14795 24701
rect 15473 24701 15485 24704
rect 15519 24701 15531 24735
rect 15580 24732 15608 24896
rect 15657 24871 15715 24877
rect 15657 24837 15669 24871
rect 15703 24868 15715 24871
rect 16316 24868 16344 24896
rect 15703 24840 16344 24868
rect 15703 24837 15715 24840
rect 15657 24831 15715 24837
rect 16500 24800 16528 24908
rect 21450 24896 21456 24908
rect 21508 24936 21514 24948
rect 24118 24936 24124 24948
rect 21508 24908 24124 24936
rect 21508 24896 21514 24908
rect 24118 24896 24124 24908
rect 24176 24896 24182 24948
rect 24581 24939 24639 24945
rect 24581 24905 24593 24939
rect 24627 24936 24639 24939
rect 24762 24936 24768 24948
rect 24627 24908 24768 24936
rect 24627 24905 24639 24908
rect 24581 24899 24639 24905
rect 24762 24896 24768 24908
rect 24820 24896 24826 24948
rect 25866 24936 25872 24948
rect 24872 24908 25872 24936
rect 21545 24871 21603 24877
rect 16592 24840 16804 24868
rect 16592 24812 16620 24840
rect 16040 24772 16528 24800
rect 16040 24741 16068 24772
rect 16574 24760 16580 24812
rect 16632 24760 16638 24812
rect 16666 24760 16672 24812
rect 16724 24760 16730 24812
rect 16776 24800 16804 24840
rect 21545 24837 21557 24871
rect 21591 24868 21603 24871
rect 22002 24868 22008 24880
rect 21591 24840 22008 24868
rect 21591 24837 21603 24840
rect 21545 24831 21603 24837
rect 22002 24828 22008 24840
rect 22060 24828 22066 24880
rect 22741 24871 22799 24877
rect 22741 24837 22753 24871
rect 22787 24868 22799 24871
rect 23569 24871 23627 24877
rect 23569 24868 23581 24871
rect 22787 24840 23581 24868
rect 22787 24837 22799 24840
rect 22741 24831 22799 24837
rect 23569 24837 23581 24840
rect 23615 24837 23627 24871
rect 23569 24831 23627 24837
rect 24302 24828 24308 24880
rect 24360 24868 24366 24880
rect 24872 24868 24900 24908
rect 25866 24896 25872 24908
rect 25924 24896 25930 24948
rect 25406 24868 25412 24880
rect 24360 24840 24900 24868
rect 24360 24828 24366 24840
rect 17037 24803 17095 24809
rect 17037 24800 17049 24803
rect 16776 24772 17049 24800
rect 17037 24769 17049 24772
rect 17083 24769 17095 24803
rect 17037 24763 17095 24769
rect 19794 24760 19800 24812
rect 19852 24800 19858 24812
rect 20165 24803 20223 24809
rect 20165 24800 20177 24803
rect 19852 24772 20177 24800
rect 19852 24760 19858 24772
rect 20165 24769 20177 24772
rect 20211 24769 20223 24803
rect 20165 24763 20223 24769
rect 21818 24760 21824 24812
rect 21876 24760 21882 24812
rect 22097 24803 22155 24809
rect 22097 24769 22109 24803
rect 22143 24800 22155 24803
rect 22554 24800 22560 24812
rect 22143 24772 22560 24800
rect 22143 24769 22155 24772
rect 22097 24763 22155 24769
rect 22554 24760 22560 24772
rect 22612 24800 22618 24812
rect 23290 24800 23296 24812
rect 22612 24772 23296 24800
rect 22612 24760 22618 24772
rect 23290 24760 23296 24772
rect 23348 24760 23354 24812
rect 23385 24803 23443 24809
rect 23385 24769 23397 24803
rect 23431 24800 23443 24803
rect 23431 24772 24440 24800
rect 23431 24769 23443 24772
rect 23385 24763 23443 24769
rect 16025 24735 16083 24741
rect 16025 24732 16037 24735
rect 15580 24704 16037 24732
rect 15473 24695 15531 24701
rect 16025 24701 16037 24704
rect 16071 24701 16083 24735
rect 16025 24695 16083 24701
rect 16298 24692 16304 24744
rect 16356 24692 16362 24744
rect 16761 24735 16819 24741
rect 16761 24701 16773 24735
rect 16807 24701 16819 24735
rect 16761 24695 16819 24701
rect 17313 24735 17371 24741
rect 17313 24701 17325 24735
rect 17359 24701 17371 24735
rect 17313 24695 17371 24701
rect 14458 24624 14464 24676
rect 14516 24664 14522 24676
rect 14553 24667 14611 24673
rect 14553 24664 14565 24667
rect 14516 24636 14565 24664
rect 14516 24624 14522 24636
rect 14553 24633 14565 24636
rect 14599 24633 14611 24667
rect 15381 24667 15439 24673
rect 15381 24664 15393 24667
rect 14553 24627 14611 24633
rect 14752 24636 15393 24664
rect 14752 24608 14780 24636
rect 15381 24633 15393 24636
rect 15427 24633 15439 24667
rect 16776 24664 16804 24695
rect 16945 24667 17003 24673
rect 16945 24664 16957 24667
rect 16776 24636 16957 24664
rect 15381 24627 15439 24633
rect 16945 24633 16957 24636
rect 16991 24633 17003 24667
rect 17328 24664 17356 24695
rect 17402 24692 17408 24744
rect 17460 24692 17466 24744
rect 18138 24692 18144 24744
rect 18196 24692 18202 24744
rect 18693 24735 18751 24741
rect 18693 24701 18705 24735
rect 18739 24732 18751 24735
rect 19812 24732 19840 24760
rect 20438 24741 20444 24744
rect 20432 24732 20444 24741
rect 18739 24704 19840 24732
rect 20399 24704 20444 24732
rect 18739 24701 18751 24704
rect 18693 24695 18751 24701
rect 20432 24695 20444 24704
rect 20438 24692 20444 24695
rect 20496 24692 20502 24744
rect 21836 24732 21864 24760
rect 22646 24732 22652 24744
rect 21836 24704 22652 24732
rect 22646 24692 22652 24704
rect 22704 24692 22710 24744
rect 23014 24692 23020 24744
rect 23072 24692 23078 24744
rect 23106 24692 23112 24744
rect 23164 24692 23170 24744
rect 23474 24692 23480 24744
rect 23532 24692 23538 24744
rect 24029 24735 24087 24741
rect 24029 24701 24041 24735
rect 24075 24732 24087 24735
rect 24118 24732 24124 24744
rect 24075 24704 24124 24732
rect 24075 24701 24087 24704
rect 24029 24695 24087 24701
rect 24118 24692 24124 24704
rect 24176 24692 24182 24744
rect 24213 24735 24271 24741
rect 24213 24701 24225 24735
rect 24259 24701 24271 24735
rect 24213 24695 24271 24701
rect 18156 24664 18184 24692
rect 18938 24667 18996 24673
rect 18938 24664 18950 24667
rect 17328 24636 18092 24664
rect 18156 24636 18950 24664
rect 16945 24627 17003 24633
rect 13136 24568 13952 24596
rect 13136 24556 13142 24568
rect 14734 24556 14740 24608
rect 14792 24556 14798 24608
rect 15194 24605 15200 24608
rect 15181 24599 15200 24605
rect 15181 24565 15193 24599
rect 15181 24559 15200 24565
rect 15194 24556 15200 24559
rect 15252 24556 15258 24608
rect 15654 24556 15660 24608
rect 15712 24596 15718 24608
rect 15841 24599 15899 24605
rect 15841 24596 15853 24599
rect 15712 24568 15853 24596
rect 15712 24556 15718 24568
rect 15841 24565 15853 24568
rect 15887 24596 15899 24599
rect 15930 24596 15936 24608
rect 15887 24568 15936 24596
rect 15887 24565 15899 24568
rect 15841 24559 15899 24565
rect 15930 24556 15936 24568
rect 15988 24556 15994 24608
rect 16960 24596 16988 24627
rect 17218 24596 17224 24608
rect 16960 24568 17224 24596
rect 17218 24556 17224 24568
rect 17276 24556 17282 24608
rect 17310 24556 17316 24608
rect 17368 24596 17374 24608
rect 17589 24599 17647 24605
rect 17589 24596 17601 24599
rect 17368 24568 17601 24596
rect 17368 24556 17374 24568
rect 17589 24565 17601 24568
rect 17635 24565 17647 24599
rect 18064 24596 18092 24636
rect 18938 24633 18950 24636
rect 18984 24633 18996 24667
rect 18938 24627 18996 24633
rect 21634 24624 21640 24676
rect 21692 24624 21698 24676
rect 18506 24596 18512 24608
rect 18064 24568 18512 24596
rect 17589 24559 17647 24565
rect 18506 24556 18512 24568
rect 18564 24556 18570 24608
rect 19702 24556 19708 24608
rect 19760 24596 19766 24608
rect 20070 24596 20076 24608
rect 19760 24568 20076 24596
rect 19760 24556 19766 24568
rect 20070 24556 20076 24568
rect 20128 24556 20134 24608
rect 22830 24556 22836 24608
rect 22888 24596 22894 24608
rect 22925 24599 22983 24605
rect 22925 24596 22937 24599
rect 22888 24568 22937 24596
rect 22888 24556 22894 24568
rect 22925 24565 22937 24568
rect 22971 24565 22983 24599
rect 22925 24559 22983 24565
rect 23750 24556 23756 24608
rect 23808 24596 23814 24608
rect 23845 24599 23903 24605
rect 23845 24596 23857 24599
rect 23808 24568 23857 24596
rect 23808 24556 23814 24568
rect 23845 24565 23857 24568
rect 23891 24565 23903 24599
rect 24228 24596 24256 24695
rect 24302 24692 24308 24744
rect 24360 24692 24366 24744
rect 24412 24664 24440 24772
rect 24872 24741 24900 24840
rect 25148 24840 25412 24868
rect 25148 24741 25176 24840
rect 25406 24828 25412 24840
rect 25464 24828 25470 24880
rect 25240 24772 25728 24800
rect 25240 24741 25268 24772
rect 24857 24735 24915 24741
rect 24857 24701 24869 24735
rect 24903 24701 24915 24735
rect 24857 24695 24915 24701
rect 25041 24735 25099 24741
rect 25041 24701 25053 24735
rect 25087 24701 25099 24735
rect 25041 24695 25099 24701
rect 25133 24735 25191 24741
rect 25133 24701 25145 24735
rect 25179 24701 25191 24735
rect 25133 24695 25191 24701
rect 25225 24735 25283 24741
rect 25225 24701 25237 24735
rect 25271 24701 25283 24735
rect 25225 24695 25283 24701
rect 24549 24667 24607 24673
rect 24549 24664 24561 24667
rect 24412 24636 24561 24664
rect 24549 24633 24561 24636
rect 24595 24633 24607 24667
rect 24549 24627 24607 24633
rect 24762 24624 24768 24676
rect 24820 24624 24826 24676
rect 25056 24664 25084 24695
rect 25498 24692 25504 24744
rect 25556 24732 25562 24744
rect 25593 24735 25651 24741
rect 25593 24732 25605 24735
rect 25556 24704 25605 24732
rect 25556 24692 25562 24704
rect 25593 24701 25605 24704
rect 25639 24701 25651 24735
rect 25700 24732 25728 24772
rect 25700 24704 26464 24732
rect 25593 24695 25651 24701
rect 25406 24664 25412 24676
rect 25056 24636 25412 24664
rect 25406 24624 25412 24636
rect 25464 24624 25470 24676
rect 25838 24667 25896 24673
rect 25838 24664 25850 24667
rect 25516 24636 25850 24664
rect 25516 24605 25544 24636
rect 25838 24633 25850 24636
rect 25884 24633 25896 24667
rect 25838 24627 25896 24633
rect 26436 24608 26464 24704
rect 24397 24599 24455 24605
rect 24397 24596 24409 24599
rect 24228 24568 24409 24596
rect 23845 24559 23903 24565
rect 24397 24565 24409 24568
rect 24443 24565 24455 24599
rect 24397 24559 24455 24565
rect 25501 24599 25559 24605
rect 25501 24565 25513 24599
rect 25547 24565 25559 24599
rect 25501 24559 25559 24565
rect 26418 24556 26424 24608
rect 26476 24556 26482 24608
rect 26970 24556 26976 24608
rect 27028 24556 27034 24608
rect 552 24506 27576 24528
rect 552 24454 7114 24506
rect 7166 24454 7178 24506
rect 7230 24454 7242 24506
rect 7294 24454 7306 24506
rect 7358 24454 7370 24506
rect 7422 24454 13830 24506
rect 13882 24454 13894 24506
rect 13946 24454 13958 24506
rect 14010 24454 14022 24506
rect 14074 24454 14086 24506
rect 14138 24454 20546 24506
rect 20598 24454 20610 24506
rect 20662 24454 20674 24506
rect 20726 24454 20738 24506
rect 20790 24454 20802 24506
rect 20854 24454 27262 24506
rect 27314 24454 27326 24506
rect 27378 24454 27390 24506
rect 27442 24454 27454 24506
rect 27506 24454 27518 24506
rect 27570 24454 27576 24506
rect 552 24432 27576 24454
rect 3050 24392 3056 24404
rect 2976 24364 3056 24392
rect 2041 24327 2099 24333
rect 2041 24293 2053 24327
rect 2087 24324 2099 24327
rect 2222 24324 2228 24336
rect 2087 24296 2228 24324
rect 2087 24293 2099 24296
rect 2041 24287 2099 24293
rect 1213 24259 1271 24265
rect 1213 24225 1225 24259
rect 1259 24225 1271 24259
rect 1213 24219 1271 24225
rect 1228 24120 1256 24219
rect 1854 24216 1860 24268
rect 1912 24216 1918 24268
rect 2056 24256 2084 24287
rect 2222 24284 2228 24296
rect 2280 24284 2286 24336
rect 2501 24327 2559 24333
rect 2501 24293 2513 24327
rect 2547 24324 2559 24327
rect 2774 24324 2780 24336
rect 2547 24296 2780 24324
rect 2547 24293 2559 24296
rect 2501 24287 2559 24293
rect 2774 24284 2780 24296
rect 2832 24284 2838 24336
rect 2976 24333 3004 24364
rect 3050 24352 3056 24364
rect 3108 24352 3114 24404
rect 3142 24352 3148 24404
rect 3200 24352 3206 24404
rect 4985 24395 5043 24401
rect 4985 24361 4997 24395
rect 5031 24392 5043 24395
rect 5031 24364 6960 24392
rect 5031 24361 5043 24364
rect 4985 24355 5043 24361
rect 2961 24327 3019 24333
rect 2961 24293 2973 24327
rect 3007 24293 3019 24327
rect 3160 24324 3188 24352
rect 3160 24296 3280 24324
rect 2961 24287 3019 24293
rect 2133 24259 2191 24265
rect 2133 24256 2145 24259
rect 2056 24228 2145 24256
rect 2133 24225 2145 24228
rect 2179 24225 2191 24259
rect 2133 24219 2191 24225
rect 1673 24191 1731 24197
rect 1673 24157 1685 24191
rect 1719 24188 1731 24191
rect 2976 24188 3004 24287
rect 3252 24265 3280 24296
rect 4798 24284 4804 24336
rect 4856 24324 4862 24336
rect 5629 24327 5687 24333
rect 4856 24296 4936 24324
rect 4856 24284 4862 24296
rect 3510 24265 3516 24268
rect 3126 24259 3184 24265
rect 3126 24256 3138 24259
rect 1719 24160 3004 24188
rect 3068 24228 3138 24256
rect 1719 24157 1731 24160
rect 1673 24151 1731 24157
rect 2685 24123 2743 24129
rect 2685 24120 2697 24123
rect 1228 24092 2697 24120
rect 2685 24089 2697 24092
rect 2731 24089 2743 24123
rect 2685 24083 2743 24089
rect 1029 24055 1087 24061
rect 1029 24021 1041 24055
rect 1075 24052 1087 24055
rect 1118 24052 1124 24064
rect 1075 24024 1124 24052
rect 1075 24021 1087 24024
rect 1029 24015 1087 24021
rect 1118 24012 1124 24024
rect 1176 24012 1182 24064
rect 2501 24055 2559 24061
rect 2501 24021 2513 24055
rect 2547 24052 2559 24055
rect 2777 24055 2835 24061
rect 2777 24052 2789 24055
rect 2547 24024 2789 24052
rect 2547 24021 2559 24024
rect 2501 24015 2559 24021
rect 2777 24021 2789 24024
rect 2823 24021 2835 24055
rect 3068 24052 3096 24228
rect 3126 24225 3138 24228
rect 3172 24225 3184 24259
rect 3126 24219 3184 24225
rect 3237 24259 3295 24265
rect 3237 24225 3249 24259
rect 3283 24225 3295 24259
rect 3237 24219 3295 24225
rect 3504 24219 3516 24265
rect 3510 24216 3516 24219
rect 3568 24216 3574 24268
rect 4908 24265 4936 24296
rect 5629 24293 5641 24327
rect 5675 24324 5687 24327
rect 6086 24324 6092 24336
rect 5675 24296 6092 24324
rect 5675 24293 5687 24296
rect 5629 24287 5687 24293
rect 6086 24284 6092 24296
rect 6144 24284 6150 24336
rect 6932 24324 6960 24364
rect 7006 24352 7012 24404
rect 7064 24392 7070 24404
rect 7064 24364 7604 24392
rect 7064 24352 7070 24364
rect 7576 24324 7604 24364
rect 7650 24352 7656 24404
rect 7708 24352 7714 24404
rect 7760 24364 8432 24392
rect 7760 24324 7788 24364
rect 6932 24296 7512 24324
rect 7576 24296 7788 24324
rect 8404 24324 8432 24364
rect 8662 24352 8668 24404
rect 8720 24352 8726 24404
rect 9401 24395 9459 24401
rect 9401 24361 9413 24395
rect 9447 24392 9459 24395
rect 10318 24392 10324 24404
rect 9447 24364 10324 24392
rect 9447 24361 9459 24364
rect 9401 24355 9459 24361
rect 9416 24324 9444 24355
rect 10318 24352 10324 24364
rect 10376 24352 10382 24404
rect 10410 24352 10416 24404
rect 10468 24392 10474 24404
rect 10965 24395 11023 24401
rect 10965 24392 10977 24395
rect 10468 24364 10977 24392
rect 10468 24352 10474 24364
rect 10965 24361 10977 24364
rect 11011 24361 11023 24395
rect 10965 24355 11023 24361
rect 11701 24395 11759 24401
rect 11701 24361 11713 24395
rect 11747 24361 11759 24395
rect 11701 24355 11759 24361
rect 10226 24324 10232 24336
rect 8404 24296 9444 24324
rect 9646 24296 10232 24324
rect 4893 24259 4951 24265
rect 4893 24225 4905 24259
rect 4939 24225 4951 24259
rect 4893 24219 4951 24225
rect 5258 24216 5264 24268
rect 5316 24216 5322 24268
rect 6178 24216 6184 24268
rect 6236 24216 6242 24268
rect 6273 24259 6331 24265
rect 6273 24225 6285 24259
rect 6319 24225 6331 24259
rect 6273 24219 6331 24225
rect 6288 24188 6316 24219
rect 6454 24216 6460 24268
rect 6512 24256 6518 24268
rect 6549 24259 6607 24265
rect 6549 24256 6561 24259
rect 6512 24228 6561 24256
rect 6512 24216 6518 24228
rect 6549 24225 6561 24228
rect 6595 24225 6607 24259
rect 6549 24219 6607 24225
rect 6822 24216 6828 24268
rect 6880 24216 6886 24268
rect 7006 24216 7012 24268
rect 7064 24216 7070 24268
rect 7116 24265 7144 24296
rect 7484 24266 7512 24296
rect 7484 24265 7604 24266
rect 7101 24259 7159 24265
rect 7101 24225 7113 24259
rect 7147 24225 7159 24259
rect 7101 24219 7159 24225
rect 7193 24259 7251 24265
rect 7193 24225 7205 24259
rect 7239 24256 7251 24259
rect 7377 24259 7435 24265
rect 7239 24228 7328 24256
rect 7239 24225 7251 24228
rect 7193 24219 7251 24225
rect 6288 24160 7232 24188
rect 4617 24123 4675 24129
rect 4617 24089 4629 24123
rect 4663 24120 4675 24123
rect 4890 24120 4896 24132
rect 4663 24092 4896 24120
rect 4663 24089 4675 24092
rect 4617 24083 4675 24089
rect 3418 24052 3424 24064
rect 3068 24024 3424 24052
rect 2777 24015 2835 24021
rect 3418 24012 3424 24024
rect 3476 24012 3482 24064
rect 3602 24012 3608 24064
rect 3660 24052 3666 24064
rect 4632 24052 4660 24083
rect 4890 24080 4896 24092
rect 4948 24120 4954 24132
rect 5997 24123 6055 24129
rect 4948 24092 5488 24120
rect 4948 24080 4954 24092
rect 3660 24024 4660 24052
rect 5460 24052 5488 24092
rect 5997 24089 6009 24123
rect 6043 24120 6055 24123
rect 6546 24120 6552 24132
rect 6043 24092 6552 24120
rect 6043 24089 6055 24092
rect 5997 24083 6055 24089
rect 6546 24080 6552 24092
rect 6604 24080 6610 24132
rect 6656 24092 6960 24120
rect 6362 24052 6368 24064
rect 5460 24024 6368 24052
rect 3660 24012 3666 24024
rect 6362 24012 6368 24024
rect 6420 24012 6426 24064
rect 6454 24012 6460 24064
rect 6512 24012 6518 24064
rect 6656 24061 6684 24092
rect 6932 24064 6960 24092
rect 6641 24055 6699 24061
rect 6641 24021 6653 24055
rect 6687 24021 6699 24055
rect 6641 24015 6699 24021
rect 6914 24012 6920 24064
rect 6972 24012 6978 24064
rect 7204 24052 7232 24160
rect 7300 24120 7328 24228
rect 7377 24225 7389 24259
rect 7423 24225 7435 24259
rect 7484 24259 7652 24265
rect 7484 24238 7606 24259
rect 7576 24228 7606 24238
rect 7377 24219 7435 24225
rect 7594 24225 7606 24228
rect 7640 24225 7652 24259
rect 7594 24219 7652 24225
rect 7392 24188 7420 24219
rect 7926 24216 7932 24268
rect 7984 24256 7990 24268
rect 8021 24259 8079 24265
rect 8021 24256 8033 24259
rect 7984 24228 8033 24256
rect 7984 24216 7990 24228
rect 8021 24225 8033 24228
rect 8067 24256 8079 24259
rect 8205 24259 8263 24265
rect 8205 24256 8217 24259
rect 8067 24228 8217 24256
rect 8067 24225 8079 24228
rect 8021 24219 8079 24225
rect 8205 24225 8217 24228
rect 8251 24225 8263 24259
rect 8205 24219 8263 24225
rect 8389 24259 8447 24265
rect 8389 24225 8401 24259
rect 8435 24225 8447 24259
rect 8389 24219 8447 24225
rect 7466 24188 7472 24200
rect 7392 24160 7472 24188
rect 7466 24148 7472 24160
rect 7524 24148 7530 24200
rect 8110 24148 8116 24200
rect 8168 24188 8174 24200
rect 8404 24188 8432 24219
rect 8846 24216 8852 24268
rect 8904 24216 8910 24268
rect 8938 24216 8944 24268
rect 8996 24216 9002 24268
rect 9033 24259 9091 24265
rect 9033 24225 9045 24259
rect 9079 24225 9091 24259
rect 9033 24219 9091 24225
rect 9217 24259 9275 24265
rect 9217 24225 9229 24259
rect 9263 24256 9275 24259
rect 9398 24256 9404 24268
rect 9263 24228 9404 24256
rect 9263 24225 9275 24228
rect 9217 24219 9275 24225
rect 8168 24160 8432 24188
rect 8168 24148 8174 24160
rect 8570 24148 8576 24200
rect 8628 24188 8634 24200
rect 9048 24188 9076 24219
rect 9398 24216 9404 24228
rect 9456 24216 9462 24268
rect 9646 24256 9674 24296
rect 10226 24284 10232 24296
rect 10284 24284 10290 24336
rect 10536 24327 10594 24333
rect 10536 24293 10548 24327
rect 10582 24324 10594 24327
rect 11716 24324 11744 24355
rect 11790 24352 11796 24404
rect 11848 24392 11854 24404
rect 13078 24392 13084 24404
rect 11848 24364 12296 24392
rect 11848 24352 11854 24364
rect 10582 24296 11744 24324
rect 10582 24293 10594 24296
rect 10536 24287 10594 24293
rect 9508 24228 9674 24256
rect 9508 24188 9536 24228
rect 10042 24216 10048 24268
rect 10100 24256 10106 24268
rect 10781 24259 10839 24265
rect 10100 24228 10732 24256
rect 10100 24216 10106 24228
rect 8628 24160 9536 24188
rect 10704 24188 10732 24228
rect 10781 24225 10793 24259
rect 10827 24256 10839 24259
rect 10962 24256 10968 24268
rect 10827 24228 10968 24256
rect 10827 24225 10839 24228
rect 10781 24219 10839 24225
rect 10962 24216 10968 24228
rect 11020 24216 11026 24268
rect 11885 24259 11943 24265
rect 11885 24256 11897 24259
rect 11072 24228 11897 24256
rect 11072 24188 11100 24228
rect 11885 24225 11897 24228
rect 11931 24225 11943 24259
rect 11885 24219 11943 24225
rect 11977 24259 12035 24265
rect 11977 24225 11989 24259
rect 12023 24225 12035 24259
rect 11977 24219 12035 24225
rect 12069 24259 12127 24265
rect 12069 24225 12081 24259
rect 12115 24256 12127 24259
rect 12158 24256 12164 24268
rect 12115 24228 12164 24256
rect 12115 24225 12127 24228
rect 12069 24219 12127 24225
rect 11517 24191 11575 24197
rect 11517 24188 11529 24191
rect 10704 24160 11100 24188
rect 11348 24160 11529 24188
rect 8628 24148 8634 24160
rect 7300 24092 7696 24120
rect 7668 24064 7696 24092
rect 7926 24080 7932 24132
rect 7984 24120 7990 24132
rect 8297 24123 8355 24129
rect 8297 24120 8309 24123
rect 7984 24092 8309 24120
rect 7984 24080 7990 24092
rect 8297 24089 8309 24092
rect 8343 24089 8355 24123
rect 8297 24083 8355 24089
rect 11348 24064 11376 24160
rect 11517 24157 11529 24160
rect 11563 24157 11575 24191
rect 11517 24151 11575 24157
rect 11992 24120 12020 24219
rect 12158 24216 12164 24228
rect 12216 24216 12222 24268
rect 12268 24265 12296 24364
rect 12728 24364 13084 24392
rect 12728 24265 12756 24364
rect 13078 24352 13084 24364
rect 13136 24352 13142 24404
rect 14093 24395 14151 24401
rect 14093 24361 14105 24395
rect 14139 24361 14151 24395
rect 14093 24355 14151 24361
rect 14645 24395 14703 24401
rect 14645 24361 14657 24395
rect 14691 24392 14703 24395
rect 15105 24395 15163 24401
rect 15105 24392 15117 24395
rect 14691 24364 15117 24392
rect 14691 24361 14703 24364
rect 14645 24355 14703 24361
rect 15105 24361 15117 24364
rect 15151 24361 15163 24395
rect 15105 24355 15163 24361
rect 12897 24327 12955 24333
rect 12897 24293 12909 24327
rect 12943 24324 12955 24327
rect 13265 24327 13323 24333
rect 13265 24324 13277 24327
rect 12943 24296 13277 24324
rect 12943 24293 12955 24296
rect 12897 24287 12955 24293
rect 13265 24293 13277 24296
rect 13311 24293 13323 24327
rect 13265 24287 13323 24293
rect 13722 24284 13728 24336
rect 13780 24284 13786 24336
rect 13930 24327 13988 24333
rect 13930 24293 13942 24327
rect 13976 24324 13988 24327
rect 14108 24324 14136 24355
rect 15194 24352 15200 24404
rect 15252 24352 15258 24404
rect 15286 24352 15292 24404
rect 15344 24352 15350 24404
rect 15470 24352 15476 24404
rect 15528 24352 15534 24404
rect 16298 24401 16304 24404
rect 16294 24392 16304 24401
rect 16259 24364 16304 24392
rect 16294 24355 16304 24364
rect 16298 24352 16304 24355
rect 16356 24352 16362 24404
rect 16574 24352 16580 24404
rect 16632 24352 16638 24404
rect 17218 24352 17224 24404
rect 17276 24352 17282 24404
rect 17310 24352 17316 24404
rect 17368 24352 17374 24404
rect 17402 24352 17408 24404
rect 17460 24352 17466 24404
rect 18049 24395 18107 24401
rect 18049 24392 18061 24395
rect 17696 24364 18061 24392
rect 15212 24324 15240 24352
rect 13976 24296 14044 24324
rect 14108 24296 15240 24324
rect 15304 24324 15332 24352
rect 16393 24327 16451 24333
rect 15304 24296 16160 24324
rect 13976 24293 13988 24296
rect 13930 24287 13988 24293
rect 12253 24259 12311 24265
rect 12253 24225 12265 24259
rect 12299 24225 12311 24259
rect 12253 24219 12311 24225
rect 12713 24259 12771 24265
rect 12713 24225 12725 24259
rect 12759 24225 12771 24259
rect 12713 24219 12771 24225
rect 12805 24259 12863 24265
rect 12805 24225 12817 24259
rect 12851 24225 12863 24259
rect 12805 24219 12863 24225
rect 12989 24259 13047 24265
rect 12989 24225 13001 24259
rect 13035 24256 13047 24259
rect 13814 24256 13820 24268
rect 13035 24228 13820 24256
rect 13035 24225 13047 24228
rect 12989 24219 13047 24225
rect 12621 24191 12679 24197
rect 12621 24157 12633 24191
rect 12667 24188 12679 24191
rect 12820 24188 12848 24219
rect 13814 24216 13820 24228
rect 13872 24216 13878 24268
rect 14016 24188 14044 24296
rect 14185 24259 14243 24265
rect 14185 24225 14197 24259
rect 14231 24256 14243 24259
rect 14231 24228 14964 24256
rect 14231 24225 14243 24228
rect 14185 24219 14243 24225
rect 14274 24188 14280 24200
rect 12667 24160 13216 24188
rect 14016 24160 14280 24188
rect 12667 24157 12679 24160
rect 12621 24151 12679 24157
rect 12802 24120 12808 24132
rect 11992 24092 12808 24120
rect 12802 24080 12808 24092
rect 12860 24080 12866 24132
rect 13188 24064 13216 24160
rect 14274 24148 14280 24160
rect 14332 24148 14338 24200
rect 14734 24148 14740 24200
rect 14792 24148 14798 24200
rect 14936 24188 14964 24228
rect 15010 24216 15016 24268
rect 15068 24216 15074 24268
rect 15197 24259 15255 24265
rect 15197 24225 15209 24259
rect 15243 24256 15255 24259
rect 15378 24256 15384 24268
rect 15243 24228 15384 24256
rect 15243 24225 15255 24228
rect 15197 24219 15255 24225
rect 15378 24216 15384 24228
rect 15436 24216 15442 24268
rect 15562 24216 15568 24268
rect 15620 24216 15626 24268
rect 16132 24265 16160 24296
rect 16393 24293 16405 24327
rect 16439 24324 16451 24327
rect 17328 24324 17356 24352
rect 16439 24296 17356 24324
rect 17420 24324 17448 24352
rect 17696 24324 17724 24364
rect 18049 24361 18061 24364
rect 18095 24361 18107 24395
rect 18049 24355 18107 24361
rect 18233 24395 18291 24401
rect 18233 24361 18245 24395
rect 18279 24361 18291 24395
rect 18233 24355 18291 24361
rect 17420 24296 17724 24324
rect 18248 24324 18276 24355
rect 18506 24352 18512 24404
rect 18564 24392 18570 24404
rect 18877 24395 18935 24401
rect 18877 24392 18889 24395
rect 18564 24364 18889 24392
rect 18564 24352 18570 24364
rect 18877 24361 18889 24364
rect 18923 24361 18935 24395
rect 18877 24355 18935 24361
rect 22646 24352 22652 24404
rect 22704 24352 22710 24404
rect 22922 24352 22928 24404
rect 22980 24392 22986 24404
rect 23017 24395 23075 24401
rect 23017 24392 23029 24395
rect 22980 24364 23029 24392
rect 22980 24352 22986 24364
rect 23017 24361 23029 24364
rect 23063 24361 23075 24395
rect 23017 24355 23075 24361
rect 19334 24324 19340 24336
rect 18248 24296 19340 24324
rect 16439 24293 16451 24296
rect 16393 24287 16451 24293
rect 16117 24259 16175 24265
rect 16117 24225 16129 24259
rect 16163 24225 16175 24259
rect 16117 24219 16175 24225
rect 16209 24259 16267 24265
rect 16209 24225 16221 24259
rect 16255 24256 16267 24259
rect 16255 24228 16436 24256
rect 16255 24225 16267 24228
rect 16209 24219 16267 24225
rect 16408 24200 16436 24228
rect 16758 24216 16764 24268
rect 16816 24216 16822 24268
rect 16853 24259 16911 24265
rect 16853 24225 16865 24259
rect 16899 24225 16911 24259
rect 16853 24219 16911 24225
rect 15470 24188 15476 24200
rect 14936 24160 15476 24188
rect 15470 24148 15476 24160
rect 15528 24148 15534 24200
rect 16390 24148 16396 24200
rect 16448 24148 16454 24200
rect 13633 24123 13691 24129
rect 13633 24089 13645 24123
rect 13679 24120 13691 24123
rect 14458 24120 14464 24132
rect 13679 24092 14464 24120
rect 13679 24089 13691 24092
rect 13633 24083 13691 24089
rect 14458 24080 14464 24092
rect 14516 24080 14522 24132
rect 14553 24123 14611 24129
rect 14553 24089 14565 24123
rect 14599 24089 14611 24123
rect 14553 24083 14611 24089
rect 14829 24123 14887 24129
rect 14829 24089 14841 24123
rect 14875 24120 14887 24123
rect 15657 24123 15715 24129
rect 15657 24120 15669 24123
rect 14875 24092 15669 24120
rect 14875 24089 14887 24092
rect 14829 24083 14887 24089
rect 15657 24089 15669 24092
rect 15703 24089 15715 24123
rect 16776 24120 16804 24216
rect 16868 24188 16896 24219
rect 16942 24216 16948 24268
rect 17000 24216 17006 24268
rect 17034 24216 17040 24268
rect 17092 24256 17098 24268
rect 17129 24259 17187 24265
rect 17129 24256 17141 24259
rect 17092 24228 17141 24256
rect 17092 24216 17098 24228
rect 17129 24225 17141 24228
rect 17175 24225 17187 24259
rect 17129 24219 17187 24225
rect 17494 24216 17500 24268
rect 17552 24216 17558 24268
rect 17696 24265 17724 24296
rect 19334 24284 19340 24296
rect 19392 24284 19398 24336
rect 17589 24259 17647 24265
rect 17589 24225 17601 24259
rect 17635 24225 17647 24259
rect 17589 24219 17647 24225
rect 17681 24259 17739 24265
rect 17681 24225 17693 24259
rect 17727 24225 17739 24259
rect 17681 24219 17739 24225
rect 17865 24259 17923 24265
rect 17865 24225 17877 24259
rect 17911 24225 17923 24259
rect 17865 24219 17923 24225
rect 18230 24259 18288 24265
rect 18230 24225 18242 24259
rect 18276 24256 18288 24259
rect 18322 24256 18328 24268
rect 18276 24228 18328 24256
rect 18276 24225 18288 24228
rect 18230 24219 18288 24225
rect 17512 24188 17540 24216
rect 16868 24160 17540 24188
rect 17604 24120 17632 24219
rect 17880 24188 17908 24219
rect 18322 24216 18328 24228
rect 18380 24216 18386 24268
rect 18414 24216 18420 24268
rect 18472 24256 18478 24268
rect 18601 24259 18659 24265
rect 18601 24256 18613 24259
rect 18472 24228 18613 24256
rect 18472 24216 18478 24228
rect 18601 24225 18613 24228
rect 18647 24256 18659 24259
rect 18782 24256 18788 24268
rect 18647 24228 18788 24256
rect 18647 24225 18659 24228
rect 18601 24219 18659 24225
rect 18782 24216 18788 24228
rect 18840 24216 18846 24268
rect 19705 24259 19763 24265
rect 19705 24225 19717 24259
rect 19751 24256 19763 24259
rect 19794 24256 19800 24268
rect 19751 24228 19800 24256
rect 19751 24225 19763 24228
rect 19705 24219 19763 24225
rect 19794 24216 19800 24228
rect 19852 24216 19858 24268
rect 19978 24265 19984 24268
rect 19972 24219 19984 24265
rect 19978 24216 19984 24219
rect 20036 24216 20042 24268
rect 21634 24216 21640 24268
rect 21692 24256 21698 24268
rect 22005 24259 22063 24265
rect 22005 24256 22017 24259
rect 21692 24228 22017 24256
rect 21692 24216 21698 24228
rect 22005 24225 22017 24228
rect 22051 24225 22063 24259
rect 22005 24219 22063 24225
rect 22557 24259 22615 24265
rect 22557 24225 22569 24259
rect 22603 24256 22615 24259
rect 22664 24256 22692 24352
rect 22603 24228 22692 24256
rect 23032 24256 23060 24355
rect 23474 24352 23480 24404
rect 23532 24352 23538 24404
rect 23658 24352 23664 24404
rect 23716 24352 23722 24404
rect 23930 24395 23988 24401
rect 23930 24361 23942 24395
rect 23976 24392 23988 24395
rect 24302 24392 24308 24404
rect 23976 24364 24308 24392
rect 23976 24361 23988 24364
rect 23930 24355 23988 24361
rect 24302 24352 24308 24364
rect 24360 24352 24366 24404
rect 24854 24352 24860 24404
rect 24912 24392 24918 24404
rect 24912 24364 25084 24392
rect 24912 24352 24918 24364
rect 23109 24259 23167 24265
rect 23109 24256 23121 24259
rect 23032 24228 23121 24256
rect 22603 24225 22615 24228
rect 22557 24219 22615 24225
rect 23109 24225 23121 24228
rect 23155 24225 23167 24259
rect 23109 24219 23167 24225
rect 23201 24259 23259 24265
rect 23201 24225 23213 24259
rect 23247 24225 23259 24259
rect 23201 24219 23259 24225
rect 17880 24160 18460 24188
rect 16776 24092 17632 24120
rect 15657 24083 15715 24089
rect 7374 24052 7380 24064
rect 7204 24024 7380 24052
rect 7374 24012 7380 24024
rect 7432 24052 7438 24064
rect 7469 24055 7527 24061
rect 7469 24052 7481 24055
rect 7432 24024 7481 24052
rect 7432 24012 7438 24024
rect 7469 24021 7481 24024
rect 7515 24021 7527 24055
rect 7469 24015 7527 24021
rect 7650 24012 7656 24064
rect 7708 24052 7714 24064
rect 11330 24052 11336 24064
rect 7708 24024 11336 24052
rect 7708 24012 7714 24024
rect 11330 24012 11336 24024
rect 11388 24012 11394 24064
rect 13078 24012 13084 24064
rect 13136 24012 13142 24064
rect 13170 24012 13176 24064
rect 13228 24012 13234 24064
rect 13265 24055 13323 24061
rect 13265 24021 13277 24055
rect 13311 24052 13323 24055
rect 13446 24052 13452 24064
rect 13311 24024 13452 24052
rect 13311 24021 13323 24024
rect 13265 24015 13323 24021
rect 13446 24012 13452 24024
rect 13504 24012 13510 24064
rect 13909 24055 13967 24061
rect 13909 24021 13921 24055
rect 13955 24052 13967 24055
rect 14182 24052 14188 24064
rect 13955 24024 14188 24052
rect 13955 24021 13967 24024
rect 13909 24015 13967 24021
rect 14182 24012 14188 24024
rect 14240 24012 14246 24064
rect 14568 24052 14596 24083
rect 18432 24064 18460 24160
rect 18690 24148 18696 24200
rect 18748 24148 18754 24200
rect 21821 24191 21879 24197
rect 21821 24157 21833 24191
rect 21867 24188 21879 24191
rect 22465 24191 22523 24197
rect 21867 24160 21901 24188
rect 21867 24157 21879 24160
rect 21821 24151 21879 24157
rect 22465 24157 22477 24191
rect 22511 24188 22523 24191
rect 22830 24188 22836 24200
rect 22511 24160 22836 24188
rect 22511 24157 22523 24160
rect 22465 24151 22523 24157
rect 19061 24123 19119 24129
rect 19061 24089 19073 24123
rect 19107 24120 19119 24123
rect 19702 24120 19708 24132
rect 19107 24092 19708 24120
rect 19107 24089 19119 24092
rect 19061 24083 19119 24089
rect 19702 24080 19708 24092
rect 19760 24080 19766 24132
rect 21085 24123 21143 24129
rect 21085 24089 21097 24123
rect 21131 24120 21143 24123
rect 21836 24120 21864 24151
rect 22830 24148 22836 24160
rect 22888 24188 22894 24200
rect 23216 24188 23244 24219
rect 23290 24216 23296 24268
rect 23348 24256 23354 24268
rect 23385 24259 23443 24265
rect 23385 24256 23397 24259
rect 23348 24228 23397 24256
rect 23348 24216 23354 24228
rect 23385 24225 23397 24228
rect 23431 24225 23443 24259
rect 23385 24219 23443 24225
rect 22888 24160 23244 24188
rect 22888 24148 22894 24160
rect 21131 24092 22876 24120
rect 21131 24089 21143 24092
rect 21085 24083 21143 24089
rect 15194 24052 15200 24064
rect 14568 24024 15200 24052
rect 15194 24012 15200 24024
rect 15252 24012 15258 24064
rect 18414 24012 18420 24064
rect 18472 24012 18478 24064
rect 21266 24012 21272 24064
rect 21324 24012 21330 24064
rect 22002 24012 22008 24064
rect 22060 24052 22066 24064
rect 22848 24061 22876 24092
rect 22097 24055 22155 24061
rect 22097 24052 22109 24055
rect 22060 24024 22109 24052
rect 22060 24012 22066 24024
rect 22097 24021 22109 24024
rect 22143 24021 22155 24055
rect 22097 24015 22155 24021
rect 22833 24055 22891 24061
rect 22833 24021 22845 24055
rect 22879 24052 22891 24055
rect 23492 24052 23520 24352
rect 23676 24256 23704 24352
rect 23845 24327 23903 24333
rect 23845 24293 23857 24327
rect 23891 24324 23903 24327
rect 24762 24324 24768 24336
rect 23891 24296 24768 24324
rect 23891 24293 23903 24296
rect 23845 24287 23903 24293
rect 24762 24284 24768 24296
rect 24820 24284 24826 24336
rect 24949 24327 25007 24333
rect 24949 24293 24961 24327
rect 24995 24293 25007 24327
rect 25056 24324 25084 24364
rect 25406 24352 25412 24404
rect 25464 24392 25470 24404
rect 25501 24395 25559 24401
rect 25501 24392 25513 24395
rect 25464 24364 25513 24392
rect 25464 24352 25470 24364
rect 25501 24361 25513 24364
rect 25547 24361 25559 24395
rect 25501 24355 25559 24361
rect 26418 24352 26424 24404
rect 26476 24352 26482 24404
rect 26970 24352 26976 24404
rect 27028 24352 27034 24404
rect 25149 24327 25207 24333
rect 25149 24324 25161 24327
rect 25056 24296 25161 24324
rect 24949 24287 25007 24293
rect 25149 24293 25161 24296
rect 25195 24293 25207 24327
rect 26988 24324 27016 24352
rect 25149 24287 25207 24293
rect 25240 24296 27016 24324
rect 23753 24259 23811 24265
rect 23753 24256 23765 24259
rect 23676 24228 23765 24256
rect 23753 24225 23765 24228
rect 23799 24225 23811 24259
rect 23753 24219 23811 24225
rect 24029 24259 24087 24265
rect 24029 24225 24041 24259
rect 24075 24256 24087 24259
rect 24673 24259 24731 24265
rect 24075 24228 24624 24256
rect 24075 24225 24087 24228
rect 24029 24219 24087 24225
rect 23569 24191 23627 24197
rect 23569 24157 23581 24191
rect 23615 24188 23627 24191
rect 24394 24188 24400 24200
rect 23615 24160 24400 24188
rect 23615 24157 23627 24160
rect 23569 24151 23627 24157
rect 24394 24148 24400 24160
rect 24452 24148 24458 24200
rect 24596 24188 24624 24228
rect 24673 24225 24685 24259
rect 24719 24256 24731 24259
rect 24964 24256 24992 24287
rect 25240 24256 25268 24296
rect 24719 24228 25268 24256
rect 25593 24259 25651 24265
rect 24719 24225 24731 24228
rect 24673 24219 24731 24225
rect 25593 24225 25605 24259
rect 25639 24256 25651 24259
rect 25961 24259 26019 24265
rect 25961 24256 25973 24259
rect 25639 24228 25973 24256
rect 25639 24225 25651 24228
rect 25593 24219 25651 24225
rect 25961 24225 25973 24228
rect 26007 24225 26019 24259
rect 25961 24219 26019 24225
rect 26145 24259 26203 24265
rect 26145 24225 26157 24259
rect 26191 24256 26203 24259
rect 26234 24256 26240 24268
rect 26191 24228 26240 24256
rect 26191 24225 26203 24228
rect 26145 24219 26203 24225
rect 25038 24188 25044 24200
rect 24596 24160 25044 24188
rect 25038 24148 25044 24160
rect 25096 24148 25102 24200
rect 25317 24123 25375 24129
rect 25317 24089 25329 24123
rect 25363 24120 25375 24123
rect 25608 24120 25636 24219
rect 25976 24188 26004 24219
rect 26234 24216 26240 24228
rect 26292 24216 26298 24268
rect 26988 24265 27016 24296
rect 26973 24259 27031 24265
rect 26973 24225 26985 24259
rect 27019 24225 27031 24259
rect 26973 24219 27031 24225
rect 25976 24160 26464 24188
rect 25363 24092 25636 24120
rect 25363 24089 25375 24092
rect 25317 24083 25375 24089
rect 26436 24064 26464 24160
rect 22879 24024 23520 24052
rect 22879 24021 22891 24024
rect 22833 24015 22891 24021
rect 24578 24012 24584 24064
rect 24636 24012 24642 24064
rect 25133 24055 25191 24061
rect 25133 24021 25145 24055
rect 25179 24052 25191 24055
rect 25958 24052 25964 24064
rect 25179 24024 25964 24052
rect 25179 24021 25191 24024
rect 25133 24015 25191 24021
rect 25958 24012 25964 24024
rect 26016 24012 26022 24064
rect 26050 24012 26056 24064
rect 26108 24012 26114 24064
rect 26418 24012 26424 24064
rect 26476 24012 26482 24064
rect 552 23962 27416 23984
rect 552 23910 3756 23962
rect 3808 23910 3820 23962
rect 3872 23910 3884 23962
rect 3936 23910 3948 23962
rect 4000 23910 4012 23962
rect 4064 23910 10472 23962
rect 10524 23910 10536 23962
rect 10588 23910 10600 23962
rect 10652 23910 10664 23962
rect 10716 23910 10728 23962
rect 10780 23910 17188 23962
rect 17240 23910 17252 23962
rect 17304 23910 17316 23962
rect 17368 23910 17380 23962
rect 17432 23910 17444 23962
rect 17496 23910 23904 23962
rect 23956 23910 23968 23962
rect 24020 23910 24032 23962
rect 24084 23910 24096 23962
rect 24148 23910 24160 23962
rect 24212 23910 27416 23962
rect 552 23888 27416 23910
rect 2225 23851 2283 23857
rect 2225 23817 2237 23851
rect 2271 23848 2283 23851
rect 3050 23848 3056 23860
rect 2271 23820 3056 23848
rect 2271 23817 2283 23820
rect 2225 23811 2283 23817
rect 3050 23808 3056 23820
rect 3108 23808 3114 23860
rect 3510 23808 3516 23860
rect 3568 23808 3574 23860
rect 5169 23851 5227 23857
rect 5169 23817 5181 23851
rect 5215 23848 5227 23851
rect 5258 23848 5264 23860
rect 5215 23820 5264 23848
rect 5215 23817 5227 23820
rect 5169 23811 5227 23817
rect 4706 23740 4712 23792
rect 4764 23780 4770 23792
rect 5077 23783 5135 23789
rect 5077 23780 5089 23783
rect 4764 23752 5089 23780
rect 4764 23740 4770 23752
rect 5077 23749 5089 23752
rect 5123 23749 5135 23783
rect 5077 23743 5135 23749
rect 842 23604 848 23656
rect 900 23604 906 23656
rect 1118 23653 1124 23656
rect 1112 23644 1124 23653
rect 1079 23616 1124 23644
rect 1112 23607 1124 23616
rect 1118 23604 1124 23607
rect 1176 23604 1182 23656
rect 3326 23604 3332 23656
rect 3384 23604 3390 23656
rect 3602 23604 3608 23656
rect 3660 23604 3666 23656
rect 4709 23647 4767 23653
rect 4709 23613 4721 23647
rect 4755 23644 4767 23647
rect 5184 23644 5212 23811
rect 5258 23808 5264 23820
rect 5316 23808 5322 23860
rect 6454 23808 6460 23860
rect 6512 23808 6518 23860
rect 6546 23808 6552 23860
rect 6604 23848 6610 23860
rect 6914 23848 6920 23860
rect 6604 23820 6920 23848
rect 6604 23808 6610 23820
rect 6914 23808 6920 23820
rect 6972 23808 6978 23860
rect 8110 23808 8116 23860
rect 8168 23808 8174 23860
rect 9858 23808 9864 23860
rect 9916 23808 9922 23860
rect 10226 23808 10232 23860
rect 10284 23848 10290 23860
rect 10284 23820 11284 23848
rect 10284 23808 10290 23820
rect 4755 23616 5212 23644
rect 4755 23613 4767 23616
rect 4709 23607 4767 23613
rect 5534 23604 5540 23656
rect 5592 23653 5598 23656
rect 5592 23644 5600 23653
rect 5592 23616 5637 23644
rect 5592 23607 5600 23616
rect 5592 23604 5598 23607
rect 2682 23536 2688 23588
rect 2740 23536 2746 23588
rect 2869 23579 2927 23585
rect 2869 23545 2881 23579
rect 2915 23576 2927 23579
rect 3620 23576 3648 23604
rect 2915 23548 3648 23576
rect 4801 23579 4859 23585
rect 2915 23545 2927 23548
rect 2869 23539 2927 23545
rect 4801 23545 4813 23579
rect 4847 23576 4859 23579
rect 4847 23548 5028 23576
rect 4847 23545 4859 23548
rect 4801 23539 4859 23545
rect 5000 23520 5028 23548
rect 5166 23536 5172 23588
rect 5224 23536 5230 23588
rect 5350 23536 5356 23588
rect 5408 23536 5414 23588
rect 5445 23579 5503 23585
rect 5445 23545 5457 23579
rect 5491 23545 5503 23579
rect 6472 23576 6500 23808
rect 7558 23740 7564 23792
rect 7616 23780 7622 23792
rect 7653 23783 7711 23789
rect 7653 23780 7665 23783
rect 7616 23752 7665 23780
rect 7616 23740 7622 23752
rect 7653 23749 7665 23752
rect 7699 23749 7711 23783
rect 7653 23743 7711 23749
rect 8220 23752 9720 23780
rect 7300 23684 7972 23712
rect 7300 23653 7328 23684
rect 7944 23656 7972 23684
rect 8220 23656 8248 23752
rect 9692 23721 9720 23752
rect 9125 23715 9183 23721
rect 9125 23712 9137 23715
rect 8496 23684 9137 23712
rect 7285 23647 7343 23653
rect 7285 23613 7297 23647
rect 7331 23613 7343 23647
rect 7285 23607 7343 23613
rect 7374 23604 7380 23656
rect 7432 23604 7438 23656
rect 7558 23604 7564 23656
rect 7616 23644 7622 23656
rect 7745 23647 7803 23653
rect 7745 23644 7757 23647
rect 7616 23616 7757 23644
rect 7616 23604 7622 23616
rect 7745 23613 7757 23616
rect 7791 23613 7803 23647
rect 7745 23607 7803 23613
rect 7834 23604 7840 23656
rect 7892 23604 7898 23656
rect 7926 23604 7932 23656
rect 7984 23604 7990 23656
rect 8202 23604 8208 23656
rect 8260 23604 8266 23656
rect 8496 23653 8524 23684
rect 9125 23681 9137 23684
rect 9171 23681 9183 23715
rect 9125 23675 9183 23681
rect 9677 23715 9735 23721
rect 9677 23681 9689 23715
rect 9723 23681 9735 23715
rect 9677 23675 9735 23681
rect 8481 23647 8539 23653
rect 8481 23613 8493 23647
rect 8527 23613 8539 23647
rect 8481 23607 8539 23613
rect 8570 23604 8576 23656
rect 8628 23644 8634 23656
rect 8665 23647 8723 23653
rect 8665 23644 8677 23647
rect 8628 23616 8677 23644
rect 8628 23604 8634 23616
rect 8665 23613 8677 23616
rect 8711 23613 8723 23647
rect 8665 23607 8723 23613
rect 8846 23604 8852 23656
rect 8904 23604 8910 23656
rect 7469 23579 7527 23585
rect 6472 23548 7236 23576
rect 5445 23539 5503 23545
rect 3050 23468 3056 23520
rect 3108 23468 3114 23520
rect 3510 23468 3516 23520
rect 3568 23508 3574 23520
rect 4525 23511 4583 23517
rect 4525 23508 4537 23511
rect 3568 23480 4537 23508
rect 3568 23468 3574 23480
rect 4525 23477 4537 23480
rect 4571 23477 4583 23511
rect 4525 23471 4583 23477
rect 4890 23468 4896 23520
rect 4948 23468 4954 23520
rect 4982 23468 4988 23520
rect 5040 23468 5046 23520
rect 5258 23468 5264 23520
rect 5316 23508 5322 23520
rect 5460 23508 5488 23539
rect 5316 23480 5488 23508
rect 5316 23468 5322 23480
rect 7006 23468 7012 23520
rect 7064 23508 7070 23520
rect 7101 23511 7159 23517
rect 7101 23508 7113 23511
rect 7064 23480 7113 23508
rect 7064 23468 7070 23480
rect 7101 23477 7113 23480
rect 7147 23477 7159 23511
rect 7208 23508 7236 23548
rect 7469 23545 7481 23579
rect 7515 23576 7527 23579
rect 7852 23576 7880 23604
rect 7515 23548 7880 23576
rect 8757 23579 8815 23585
rect 7515 23545 7527 23548
rect 7469 23539 7527 23545
rect 8757 23545 8769 23579
rect 8803 23576 8815 23579
rect 9306 23576 9312 23588
rect 8803 23548 9312 23576
rect 8803 23545 8815 23548
rect 8757 23539 8815 23545
rect 9306 23536 9312 23548
rect 9364 23536 9370 23588
rect 9876 23576 9904 23808
rect 11256 23780 11284 23820
rect 11330 23808 11336 23860
rect 11388 23808 11394 23860
rect 12158 23848 12164 23860
rect 11440 23820 12164 23848
rect 11440 23780 11468 23820
rect 12158 23808 12164 23820
rect 12216 23808 12222 23860
rect 12894 23808 12900 23860
rect 12952 23808 12958 23860
rect 13078 23808 13084 23860
rect 13136 23808 13142 23860
rect 14458 23808 14464 23860
rect 14516 23808 14522 23860
rect 14829 23851 14887 23857
rect 14829 23817 14841 23851
rect 14875 23848 14887 23851
rect 15562 23848 15568 23860
rect 14875 23820 15568 23848
rect 14875 23817 14887 23820
rect 14829 23811 14887 23817
rect 11256 23752 11468 23780
rect 9953 23647 10011 23653
rect 9953 23613 9965 23647
rect 9999 23644 10011 23647
rect 11054 23644 11060 23656
rect 9999 23616 11060 23644
rect 9999 23613 10011 23616
rect 9953 23607 10011 23613
rect 11054 23604 11060 23616
rect 11112 23644 11118 23656
rect 13096 23653 13124 23808
rect 13814 23740 13820 23792
rect 13872 23780 13878 23792
rect 13872 23752 14504 23780
rect 13872 23740 13878 23752
rect 13170 23672 13176 23724
rect 13228 23712 13234 23724
rect 13228 23684 14320 23712
rect 13228 23672 13234 23684
rect 14292 23653 14320 23684
rect 14476 23653 14504 23752
rect 14734 23740 14740 23792
rect 14792 23740 14798 23792
rect 14752 23653 14780 23740
rect 11425 23647 11483 23653
rect 11425 23644 11437 23647
rect 11112 23616 11437 23644
rect 11112 23604 11118 23616
rect 11425 23613 11437 23616
rect 11471 23613 11483 23647
rect 11425 23607 11483 23613
rect 13081 23647 13139 23653
rect 13081 23613 13093 23647
rect 13127 23613 13139 23647
rect 13081 23607 13139 23613
rect 14093 23647 14151 23653
rect 14093 23613 14105 23647
rect 14139 23613 14151 23647
rect 14093 23607 14151 23613
rect 14277 23647 14335 23653
rect 14277 23613 14289 23647
rect 14323 23613 14335 23647
rect 14277 23607 14335 23613
rect 14461 23647 14519 23653
rect 14461 23613 14473 23647
rect 14507 23613 14519 23647
rect 14461 23607 14519 23613
rect 14737 23647 14795 23653
rect 14737 23613 14749 23647
rect 14783 23613 14795 23647
rect 14737 23607 14795 23613
rect 10198 23579 10256 23585
rect 10198 23576 10210 23579
rect 9876 23548 10210 23576
rect 10198 23545 10210 23548
rect 10244 23545 10256 23579
rect 10198 23539 10256 23545
rect 11692 23579 11750 23585
rect 11692 23545 11704 23579
rect 11738 23576 11750 23579
rect 11882 23576 11888 23588
rect 11738 23548 11888 23576
rect 11738 23545 11750 23548
rect 11692 23539 11750 23545
rect 11882 23536 11888 23548
rect 11940 23536 11946 23588
rect 14108 23576 14136 23607
rect 14844 23576 14872 23811
rect 15562 23808 15568 23820
rect 15620 23808 15626 23860
rect 15749 23851 15807 23857
rect 15749 23817 15761 23851
rect 15795 23848 15807 23851
rect 15838 23848 15844 23860
rect 15795 23820 15844 23848
rect 15795 23817 15807 23820
rect 15749 23811 15807 23817
rect 15838 23808 15844 23820
rect 15896 23808 15902 23860
rect 18414 23808 18420 23860
rect 18472 23848 18478 23860
rect 18969 23851 19027 23857
rect 18969 23848 18981 23851
rect 18472 23820 18981 23848
rect 18472 23808 18478 23820
rect 18969 23817 18981 23820
rect 19015 23817 19027 23851
rect 18969 23811 19027 23817
rect 19978 23808 19984 23860
rect 20036 23808 20042 23860
rect 20346 23808 20352 23860
rect 20404 23808 20410 23860
rect 21266 23808 21272 23860
rect 21324 23808 21330 23860
rect 24581 23851 24639 23857
rect 24581 23817 24593 23851
rect 24627 23848 24639 23851
rect 24762 23848 24768 23860
rect 24627 23820 24768 23848
rect 24627 23817 24639 23820
rect 24581 23811 24639 23817
rect 24762 23808 24768 23820
rect 24820 23808 24826 23860
rect 15194 23740 15200 23792
rect 15252 23740 15258 23792
rect 18506 23740 18512 23792
rect 18564 23740 18570 23792
rect 15212 23644 15240 23740
rect 18524 23712 18552 23740
rect 18524 23684 19012 23712
rect 15289 23647 15347 23653
rect 15289 23644 15301 23647
rect 15212 23616 15301 23644
rect 15289 23613 15301 23616
rect 15335 23613 15347 23647
rect 15289 23607 15347 23613
rect 15470 23604 15476 23656
rect 15528 23644 15534 23656
rect 15565 23647 15623 23653
rect 15565 23644 15577 23647
rect 15528 23616 15577 23644
rect 15528 23604 15534 23616
rect 15565 23613 15577 23616
rect 15611 23613 15623 23647
rect 15565 23607 15623 23613
rect 18693 23647 18751 23653
rect 18693 23613 18705 23647
rect 18739 23613 18751 23647
rect 18693 23607 18751 23613
rect 12820 23548 14872 23576
rect 7837 23511 7895 23517
rect 7837 23508 7849 23511
rect 7208 23480 7849 23508
rect 7101 23471 7159 23477
rect 7837 23477 7849 23480
rect 7883 23477 7895 23511
rect 7837 23471 7895 23477
rect 9030 23468 9036 23520
rect 9088 23468 9094 23520
rect 12820 23517 12848 23548
rect 18708 23520 18736 23607
rect 18782 23604 18788 23656
rect 18840 23604 18846 23656
rect 18984 23653 19012 23684
rect 18969 23647 19027 23653
rect 18969 23613 18981 23647
rect 19015 23613 19027 23647
rect 18969 23607 19027 23613
rect 19610 23604 19616 23656
rect 19668 23644 19674 23656
rect 20165 23647 20223 23653
rect 20165 23644 20177 23647
rect 19668 23616 20177 23644
rect 19668 23604 19674 23616
rect 20165 23613 20177 23616
rect 20211 23644 20223 23647
rect 20364 23644 20392 23808
rect 20211 23616 20392 23644
rect 20211 23613 20223 23616
rect 20165 23607 20223 23613
rect 20438 23604 20444 23656
rect 20496 23604 20502 23656
rect 20533 23647 20591 23653
rect 20533 23613 20545 23647
rect 20579 23644 20591 23647
rect 21284 23644 21312 23808
rect 22646 23672 22652 23724
rect 22704 23712 22710 23724
rect 23017 23715 23075 23721
rect 23017 23712 23029 23715
rect 22704 23684 23029 23712
rect 22704 23672 22710 23684
rect 23017 23681 23029 23684
rect 23063 23681 23075 23715
rect 23017 23675 23075 23681
rect 24228 23684 25820 23712
rect 20579 23616 21312 23644
rect 20579 23613 20591 23616
rect 20533 23607 20591 23613
rect 21818 23604 21824 23656
rect 21876 23604 21882 23656
rect 21910 23604 21916 23656
rect 21968 23644 21974 23656
rect 22005 23647 22063 23653
rect 22005 23644 22017 23647
rect 21968 23616 22017 23644
rect 21968 23604 21974 23616
rect 22005 23613 22017 23616
rect 22051 23644 22063 23647
rect 24228 23644 24256 23684
rect 25792 23656 25820 23684
rect 22051 23616 24256 23644
rect 22051 23613 22063 23616
rect 22005 23607 22063 23613
rect 24486 23604 24492 23656
rect 24544 23644 24550 23656
rect 24765 23647 24823 23653
rect 24765 23644 24777 23647
rect 24544 23616 24777 23644
rect 24544 23604 24550 23616
rect 24765 23613 24777 23616
rect 24811 23613 24823 23647
rect 24765 23607 24823 23613
rect 24857 23647 24915 23653
rect 24857 23613 24869 23647
rect 24903 23613 24915 23647
rect 24857 23607 24915 23613
rect 19426 23536 19432 23588
rect 19484 23576 19490 23588
rect 20257 23579 20315 23585
rect 20257 23576 20269 23579
rect 19484 23548 20269 23576
rect 19484 23536 19490 23548
rect 20257 23545 20269 23548
rect 20303 23545 20315 23579
rect 20257 23539 20315 23545
rect 20349 23579 20407 23585
rect 20349 23545 20361 23579
rect 20395 23576 20407 23579
rect 20456 23576 20484 23604
rect 20395 23548 20484 23576
rect 20395 23545 20407 23548
rect 20349 23539 20407 23545
rect 22094 23536 22100 23588
rect 22152 23576 22158 23588
rect 22465 23579 22523 23585
rect 22465 23576 22477 23579
rect 22152 23548 22477 23576
rect 22152 23536 22158 23548
rect 22465 23545 22477 23548
rect 22511 23545 22523 23579
rect 22465 23539 22523 23545
rect 24394 23536 24400 23588
rect 24452 23576 24458 23588
rect 24872 23576 24900 23607
rect 24946 23604 24952 23656
rect 25004 23604 25010 23656
rect 25498 23644 25504 23656
rect 25240 23616 25504 23644
rect 24452 23548 24900 23576
rect 24452 23536 24458 23548
rect 12805 23511 12863 23517
rect 12805 23477 12817 23511
rect 12851 23477 12863 23511
rect 12805 23471 12863 23477
rect 13538 23468 13544 23520
rect 13596 23468 13602 23520
rect 14734 23468 14740 23520
rect 14792 23508 14798 23520
rect 15010 23508 15016 23520
rect 14792 23480 15016 23508
rect 14792 23468 14798 23480
rect 15010 23468 15016 23480
rect 15068 23508 15074 23520
rect 15381 23511 15439 23517
rect 15381 23508 15393 23511
rect 15068 23480 15393 23508
rect 15068 23468 15074 23480
rect 15381 23477 15393 23480
rect 15427 23477 15439 23511
rect 15381 23471 15439 23477
rect 18690 23468 18696 23520
rect 18748 23468 18754 23520
rect 19518 23468 19524 23520
rect 19576 23508 19582 23520
rect 19794 23508 19800 23520
rect 19576 23480 19800 23508
rect 19576 23468 19582 23480
rect 19794 23468 19800 23480
rect 19852 23468 19858 23520
rect 21913 23511 21971 23517
rect 21913 23477 21925 23511
rect 21959 23508 21971 23511
rect 22186 23508 22192 23520
rect 21959 23480 22192 23508
rect 21959 23477 21971 23480
rect 21913 23471 21971 23477
rect 22186 23468 22192 23480
rect 22244 23468 22250 23520
rect 23474 23468 23480 23520
rect 23532 23508 23538 23520
rect 25240 23508 25268 23616
rect 25498 23604 25504 23616
rect 25556 23644 25562 23656
rect 25685 23647 25743 23653
rect 25685 23644 25697 23647
rect 25556 23616 25697 23644
rect 25556 23604 25562 23616
rect 25685 23613 25697 23616
rect 25731 23613 25743 23647
rect 25685 23607 25743 23613
rect 25774 23604 25780 23656
rect 25832 23604 25838 23656
rect 25590 23536 25596 23588
rect 25648 23576 25654 23588
rect 25930 23579 25988 23585
rect 25930 23576 25942 23579
rect 25648 23548 25942 23576
rect 25648 23536 25654 23548
rect 25930 23545 25942 23548
rect 25976 23545 25988 23579
rect 25930 23539 25988 23545
rect 23532 23480 25268 23508
rect 23532 23468 23538 23480
rect 26234 23468 26240 23520
rect 26292 23508 26298 23520
rect 27065 23511 27123 23517
rect 27065 23508 27077 23511
rect 26292 23480 27077 23508
rect 26292 23468 26298 23480
rect 27065 23477 27077 23480
rect 27111 23477 27123 23511
rect 27065 23471 27123 23477
rect 552 23418 27576 23440
rect 552 23366 7114 23418
rect 7166 23366 7178 23418
rect 7230 23366 7242 23418
rect 7294 23366 7306 23418
rect 7358 23366 7370 23418
rect 7422 23366 13830 23418
rect 13882 23366 13894 23418
rect 13946 23366 13958 23418
rect 14010 23366 14022 23418
rect 14074 23366 14086 23418
rect 14138 23366 20546 23418
rect 20598 23366 20610 23418
rect 20662 23366 20674 23418
rect 20726 23366 20738 23418
rect 20790 23366 20802 23418
rect 20854 23366 27262 23418
rect 27314 23366 27326 23418
rect 27378 23366 27390 23418
rect 27442 23366 27454 23418
rect 27506 23366 27518 23418
rect 27570 23366 27576 23418
rect 552 23344 27576 23366
rect 2593 23307 2651 23313
rect 2593 23273 2605 23307
rect 2639 23304 2651 23307
rect 2682 23304 2688 23316
rect 2639 23276 2688 23304
rect 2639 23273 2651 23276
rect 2593 23267 2651 23273
rect 2682 23264 2688 23276
rect 2740 23264 2746 23316
rect 2774 23264 2780 23316
rect 2832 23304 2838 23316
rect 3053 23307 3111 23313
rect 3053 23304 3065 23307
rect 2832 23276 3065 23304
rect 2832 23264 2838 23276
rect 3053 23273 3065 23276
rect 3099 23273 3111 23307
rect 3053 23267 3111 23273
rect 3237 23307 3295 23313
rect 3237 23273 3249 23307
rect 3283 23304 3295 23307
rect 3326 23304 3332 23316
rect 3283 23276 3332 23304
rect 3283 23273 3295 23276
rect 3237 23267 3295 23273
rect 3326 23264 3332 23276
rect 3384 23264 3390 23316
rect 3510 23313 3516 23316
rect 3497 23307 3516 23313
rect 3497 23304 3509 23307
rect 3436 23276 3509 23304
rect 2409 23171 2467 23177
rect 2409 23137 2421 23171
rect 2455 23168 2467 23171
rect 2866 23168 2872 23180
rect 2455 23140 2872 23168
rect 2455 23137 2467 23140
rect 2409 23131 2467 23137
rect 2866 23128 2872 23140
rect 2924 23168 2930 23180
rect 3436 23168 3464 23276
rect 3497 23273 3509 23276
rect 3497 23267 3516 23273
rect 3510 23264 3516 23267
rect 3568 23264 3574 23316
rect 4890 23264 4896 23316
rect 4948 23264 4954 23316
rect 5077 23307 5135 23313
rect 5077 23273 5089 23307
rect 5123 23304 5135 23307
rect 5442 23304 5448 23316
rect 5123 23276 5448 23304
rect 5123 23273 5135 23276
rect 5077 23267 5135 23273
rect 5442 23264 5448 23276
rect 5500 23264 5506 23316
rect 6914 23264 6920 23316
rect 6972 23304 6978 23316
rect 8113 23307 8171 23313
rect 6972 23276 7420 23304
rect 6972 23264 6978 23276
rect 3602 23196 3608 23248
rect 3660 23236 3666 23248
rect 3697 23239 3755 23245
rect 3697 23236 3709 23239
rect 3660 23208 3709 23236
rect 3660 23196 3666 23208
rect 3697 23205 3709 23208
rect 3743 23205 3755 23239
rect 3697 23199 3755 23205
rect 4801 23239 4859 23245
rect 4801 23205 4813 23239
rect 4847 23236 4859 23239
rect 4908 23236 4936 23264
rect 7101 23239 7159 23245
rect 4847 23208 5212 23236
rect 4847 23205 4859 23208
rect 4801 23199 4859 23205
rect 5184 23180 5212 23208
rect 7101 23205 7113 23239
rect 7147 23236 7159 23239
rect 7285 23239 7343 23245
rect 7285 23236 7297 23239
rect 7147 23208 7297 23236
rect 7147 23205 7159 23208
rect 7101 23199 7159 23205
rect 7285 23205 7297 23208
rect 7331 23205 7343 23239
rect 7285 23199 7343 23205
rect 2924 23140 3464 23168
rect 3973 23171 4031 23177
rect 2924 23128 2930 23140
rect 3973 23137 3985 23171
rect 4019 23168 4031 23171
rect 4062 23168 4068 23180
rect 4019 23140 4068 23168
rect 4019 23137 4031 23140
rect 3973 23131 4031 23137
rect 4062 23128 4068 23140
rect 4120 23128 4126 23180
rect 4706 23128 4712 23180
rect 4764 23128 4770 23180
rect 4893 23171 4951 23177
rect 4893 23137 4905 23171
rect 4939 23168 4951 23171
rect 4982 23168 4988 23180
rect 4939 23140 4988 23168
rect 4939 23137 4951 23140
rect 4893 23131 4951 23137
rect 4982 23128 4988 23140
rect 5040 23128 5046 23180
rect 5166 23128 5172 23180
rect 5224 23128 5230 23180
rect 5813 23171 5871 23177
rect 5813 23137 5825 23171
rect 5859 23168 5871 23171
rect 6086 23168 6092 23180
rect 5859 23140 6092 23168
rect 5859 23137 5871 23140
rect 5813 23131 5871 23137
rect 6086 23128 6092 23140
rect 6144 23128 6150 23180
rect 6822 23128 6828 23180
rect 6880 23128 6886 23180
rect 7006 23128 7012 23180
rect 7064 23168 7070 23180
rect 7193 23171 7251 23177
rect 7064 23140 7144 23168
rect 7064 23128 7070 23140
rect 2222 23060 2228 23112
rect 2280 23060 2286 23112
rect 3418 23060 3424 23112
rect 3476 23060 3482 23112
rect 7116 23109 7144 23140
rect 7193 23137 7205 23171
rect 7239 23168 7251 23171
rect 7392 23168 7420 23276
rect 8113 23273 8125 23307
rect 8159 23304 8171 23307
rect 8202 23304 8208 23316
rect 8159 23276 8208 23304
rect 8159 23273 8171 23276
rect 8113 23267 8171 23273
rect 8202 23264 8208 23276
rect 8260 23264 8266 23316
rect 9950 23264 9956 23316
rect 10008 23304 10014 23316
rect 10410 23304 10416 23316
rect 10008 23276 10416 23304
rect 10008 23264 10014 23276
rect 10410 23264 10416 23276
rect 10468 23264 10474 23316
rect 11900 23276 12296 23304
rect 7469 23239 7527 23245
rect 7469 23205 7481 23239
rect 7515 23236 7527 23239
rect 7742 23236 7748 23248
rect 7515 23208 7748 23236
rect 7515 23205 7527 23208
rect 7469 23199 7527 23205
rect 7742 23196 7748 23208
rect 7800 23196 7806 23248
rect 9030 23196 9036 23248
rect 9088 23236 9094 23248
rect 9226 23239 9284 23245
rect 9226 23236 9238 23239
rect 9088 23208 9238 23236
rect 9088 23196 9094 23208
rect 9226 23205 9238 23208
rect 9272 23205 9284 23239
rect 9226 23199 9284 23205
rect 9674 23196 9680 23248
rect 9732 23196 9738 23248
rect 10060 23208 10548 23236
rect 10060 23180 10088 23208
rect 7239 23140 7420 23168
rect 7239 23137 7251 23140
rect 7193 23131 7251 23137
rect 9858 23128 9864 23180
rect 9916 23128 9922 23180
rect 9950 23128 9956 23180
rect 10008 23128 10014 23180
rect 10042 23128 10048 23180
rect 10100 23128 10106 23180
rect 10134 23128 10140 23180
rect 10192 23128 10198 23180
rect 10226 23128 10232 23180
rect 10284 23168 10290 23180
rect 10321 23171 10379 23177
rect 10321 23168 10333 23171
rect 10284 23140 10333 23168
rect 10284 23128 10290 23140
rect 10321 23137 10333 23140
rect 10367 23137 10379 23171
rect 10321 23131 10379 23137
rect 10410 23128 10416 23180
rect 10468 23128 10474 23180
rect 10520 23177 10548 23208
rect 11146 23196 11152 23248
rect 11204 23236 11210 23248
rect 11514 23236 11520 23248
rect 11204 23208 11520 23236
rect 11204 23196 11210 23208
rect 11514 23196 11520 23208
rect 11572 23196 11578 23248
rect 11609 23239 11667 23245
rect 11609 23205 11621 23239
rect 11655 23236 11667 23239
rect 11900 23236 11928 23276
rect 12161 23239 12219 23245
rect 12161 23236 12173 23239
rect 11655 23208 11928 23236
rect 11992 23208 12173 23236
rect 11655 23205 11667 23208
rect 11609 23199 11667 23205
rect 11992 23180 12020 23208
rect 12161 23205 12173 23208
rect 12207 23205 12219 23239
rect 12161 23199 12219 23205
rect 12268 23180 12296 23276
rect 14734 23264 14740 23316
rect 14792 23264 14798 23316
rect 15289 23307 15347 23313
rect 15289 23273 15301 23307
rect 15335 23304 15347 23307
rect 15470 23304 15476 23316
rect 15335 23276 15476 23304
rect 15335 23273 15347 23276
rect 15289 23267 15347 23273
rect 15470 23264 15476 23276
rect 15528 23264 15534 23316
rect 16117 23307 16175 23313
rect 16117 23273 16129 23307
rect 16163 23304 16175 23307
rect 16574 23304 16580 23316
rect 16163 23276 16580 23304
rect 16163 23273 16175 23276
rect 16117 23267 16175 23273
rect 16574 23264 16580 23276
rect 16632 23304 16638 23316
rect 16942 23304 16948 23316
rect 16632 23276 16948 23304
rect 16632 23264 16638 23276
rect 16942 23264 16948 23276
rect 17000 23264 17006 23316
rect 19334 23264 19340 23316
rect 19392 23264 19398 23316
rect 21818 23264 21824 23316
rect 21876 23264 21882 23316
rect 22278 23304 22284 23316
rect 21928 23276 22284 23304
rect 17034 23196 17040 23248
rect 17092 23236 17098 23248
rect 17230 23239 17288 23245
rect 17230 23236 17242 23239
rect 17092 23208 17242 23236
rect 17092 23196 17098 23208
rect 17230 23205 17242 23208
rect 17276 23205 17288 23239
rect 17230 23199 17288 23205
rect 10505 23171 10563 23177
rect 10505 23137 10517 23171
rect 10551 23137 10563 23171
rect 10505 23131 10563 23137
rect 11054 23128 11060 23180
rect 11112 23128 11118 23180
rect 11425 23171 11483 23177
rect 11425 23137 11437 23171
rect 11471 23137 11483 23171
rect 11425 23131 11483 23137
rect 11793 23171 11851 23177
rect 11793 23137 11805 23171
rect 11839 23137 11851 23171
rect 11793 23131 11851 23137
rect 7101 23103 7159 23109
rect 7101 23069 7113 23103
rect 7147 23069 7159 23103
rect 7101 23063 7159 23069
rect 9493 23103 9551 23109
rect 9493 23069 9505 23103
rect 9539 23100 9551 23103
rect 11072 23100 11100 23128
rect 9539 23072 11100 23100
rect 11440 23100 11468 23131
rect 11808 23100 11836 23131
rect 11974 23128 11980 23180
rect 12032 23128 12038 23180
rect 12066 23128 12072 23180
rect 12124 23128 12130 23180
rect 12250 23128 12256 23180
rect 12308 23128 12314 23180
rect 12437 23171 12495 23177
rect 12437 23137 12449 23171
rect 12483 23168 12495 23171
rect 13538 23168 13544 23180
rect 12483 23140 13544 23168
rect 12483 23137 12495 23140
rect 12437 23131 12495 23137
rect 13538 23128 13544 23140
rect 13596 23128 13602 23180
rect 14274 23168 14280 23180
rect 13832 23140 14280 23168
rect 12529 23103 12587 23109
rect 12529 23100 12541 23103
rect 11440 23072 11560 23100
rect 11808 23072 12541 23100
rect 9539 23069 9551 23072
rect 9493 23063 9551 23069
rect 2685 23035 2743 23041
rect 2685 23001 2697 23035
rect 2731 23032 2743 23035
rect 3329 23035 3387 23041
rect 3329 23032 3341 23035
rect 2731 23004 3341 23032
rect 2731 23001 2743 23004
rect 2685 22995 2743 23001
rect 3329 23001 3341 23004
rect 3375 23032 3387 23035
rect 3436 23032 3464 23060
rect 4522 23032 4528 23044
rect 3375 23004 3464 23032
rect 3528 23004 4528 23032
rect 3375 23001 3387 23004
rect 3329 22995 3387 23001
rect 3050 22924 3056 22976
rect 3108 22924 3114 22976
rect 3528 22973 3556 23004
rect 4522 22992 4528 23004
rect 4580 22992 4586 23044
rect 6917 23035 6975 23041
rect 6917 23001 6929 23035
rect 6963 23032 6975 23035
rect 7650 23032 7656 23044
rect 6963 23004 7656 23032
rect 6963 23001 6975 23004
rect 6917 22995 6975 23001
rect 7650 22992 7656 23004
rect 7708 22992 7714 23044
rect 11532 23032 11560 23072
rect 12529 23069 12541 23072
rect 12575 23069 12587 23103
rect 12529 23063 12587 23069
rect 12802 23060 12808 23112
rect 12860 23100 12866 23112
rect 13081 23103 13139 23109
rect 13081 23100 13093 23103
rect 12860 23072 13093 23100
rect 12860 23060 12866 23072
rect 13081 23069 13093 23072
rect 13127 23069 13139 23103
rect 13081 23063 13139 23069
rect 12066 23032 12072 23044
rect 11532 23004 12072 23032
rect 12066 22992 12072 23004
rect 12124 22992 12130 23044
rect 3513 22967 3571 22973
rect 3513 22933 3525 22967
rect 3559 22933 3571 22967
rect 3513 22927 3571 22933
rect 3602 22924 3608 22976
rect 3660 22964 3666 22976
rect 3789 22967 3847 22973
rect 3789 22964 3801 22967
rect 3660 22936 3801 22964
rect 3660 22924 3666 22936
rect 3789 22933 3801 22936
rect 3835 22933 3847 22967
rect 3789 22927 3847 22933
rect 5534 22924 5540 22976
rect 5592 22964 5598 22976
rect 5905 22967 5963 22973
rect 5905 22964 5917 22967
rect 5592 22936 5917 22964
rect 5592 22924 5598 22936
rect 5905 22933 5917 22936
rect 5951 22933 5963 22967
rect 5905 22927 5963 22933
rect 6270 22924 6276 22976
rect 6328 22924 6334 22976
rect 7466 22924 7472 22976
rect 7524 22924 7530 22976
rect 10689 22967 10747 22973
rect 10689 22933 10701 22967
rect 10735 22964 10747 22967
rect 11146 22964 11152 22976
rect 10735 22936 11152 22964
rect 10735 22933 10747 22936
rect 10689 22927 10747 22933
rect 11146 22924 11152 22936
rect 11204 22924 11210 22976
rect 11238 22924 11244 22976
rect 11296 22924 11302 22976
rect 11882 22924 11888 22976
rect 11940 22924 11946 22976
rect 13096 22964 13124 23063
rect 13832 23044 13860 23140
rect 14274 23128 14280 23140
rect 14332 23168 14338 23180
rect 14829 23171 14887 23177
rect 14829 23168 14841 23171
rect 14332 23140 14841 23168
rect 14332 23128 14338 23140
rect 14829 23137 14841 23140
rect 14875 23137 14887 23171
rect 14829 23131 14887 23137
rect 17862 23128 17868 23180
rect 17920 23168 17926 23180
rect 18213 23171 18271 23177
rect 18213 23168 18225 23171
rect 17920 23140 18225 23168
rect 17920 23128 17926 23140
rect 18213 23137 18225 23140
rect 18259 23137 18271 23171
rect 19352 23168 19380 23264
rect 21928 23236 21956 23276
rect 22278 23264 22284 23276
rect 22336 23264 22342 23316
rect 22646 23264 22652 23316
rect 22704 23304 22710 23316
rect 23293 23307 23351 23313
rect 23293 23304 23305 23307
rect 22704 23276 23305 23304
rect 22704 23264 22710 23276
rect 23293 23273 23305 23276
rect 23339 23273 23351 23307
rect 23293 23267 23351 23273
rect 23753 23307 23811 23313
rect 23753 23273 23765 23307
rect 23799 23304 23811 23307
rect 24394 23304 24400 23316
rect 23799 23276 24400 23304
rect 23799 23273 23811 23276
rect 23753 23267 23811 23273
rect 24394 23264 24400 23276
rect 24452 23264 24458 23316
rect 24486 23264 24492 23316
rect 24544 23304 24550 23316
rect 25761 23307 25819 23313
rect 24544 23276 25636 23304
rect 24544 23264 24550 23276
rect 22186 23245 22192 23248
rect 20640 23208 21956 23236
rect 22158 23239 22192 23245
rect 20640 23177 20668 23208
rect 22158 23205 22170 23239
rect 22158 23199 22192 23205
rect 22186 23196 22192 23199
rect 22244 23196 22250 23248
rect 24578 23236 24584 23248
rect 23952 23208 24584 23236
rect 19981 23171 20039 23177
rect 19981 23168 19993 23171
rect 19352 23140 19993 23168
rect 18213 23131 18271 23137
rect 19981 23137 19993 23140
rect 20027 23137 20039 23171
rect 20625 23171 20683 23177
rect 20625 23168 20637 23171
rect 19981 23131 20039 23137
rect 20088 23140 20637 23168
rect 17497 23103 17555 23109
rect 17497 23069 17509 23103
rect 17543 23100 17555 23103
rect 17954 23100 17960 23112
rect 17543 23072 17960 23100
rect 17543 23069 17555 23072
rect 17497 23063 17555 23069
rect 17954 23060 17960 23072
rect 18012 23060 18018 23112
rect 13814 22992 13820 23044
rect 13872 22992 13878 23044
rect 15105 23035 15163 23041
rect 15105 23032 15117 23035
rect 14384 23004 15117 23032
rect 14384 22973 14412 23004
rect 15105 23001 15117 23004
rect 15151 23001 15163 23035
rect 20088 23032 20116 23140
rect 20625 23137 20637 23140
rect 20671 23137 20683 23171
rect 20625 23131 20683 23137
rect 21453 23171 21511 23177
rect 21453 23137 21465 23171
rect 21499 23168 21511 23171
rect 22002 23168 22008 23180
rect 21499 23140 22008 23168
rect 21499 23137 21511 23140
rect 21453 23131 21511 23137
rect 22002 23128 22008 23140
rect 22060 23128 22066 23180
rect 23952 23177 23980 23208
rect 24578 23196 24584 23208
rect 24636 23196 24642 23248
rect 24946 23196 24952 23248
rect 25004 23236 25010 23248
rect 25501 23239 25559 23245
rect 25501 23236 25513 23239
rect 25004 23208 25513 23236
rect 25004 23196 25010 23208
rect 25501 23205 25513 23208
rect 25547 23205 25559 23239
rect 25501 23199 25559 23205
rect 23661 23171 23719 23177
rect 23661 23168 23673 23171
rect 23584 23140 23673 23168
rect 20346 23060 20352 23112
rect 20404 23100 20410 23112
rect 21361 23103 21419 23109
rect 21361 23100 21373 23103
rect 20404 23072 21373 23100
rect 20404 23060 20410 23072
rect 21361 23069 21373 23072
rect 21407 23069 21419 23103
rect 21361 23063 21419 23069
rect 21910 23060 21916 23112
rect 21968 23060 21974 23112
rect 23584 23100 23612 23140
rect 23661 23137 23673 23140
rect 23707 23137 23719 23171
rect 23661 23131 23719 23137
rect 23845 23171 23903 23177
rect 23845 23137 23857 23171
rect 23891 23168 23903 23171
rect 23937 23171 23995 23177
rect 23937 23168 23949 23171
rect 23891 23140 23949 23168
rect 23891 23137 23903 23140
rect 23845 23131 23903 23137
rect 23937 23137 23949 23140
rect 23983 23137 23995 23171
rect 23937 23131 23995 23137
rect 24121 23171 24179 23177
rect 24121 23137 24133 23171
rect 24167 23137 24179 23171
rect 24121 23131 24179 23137
rect 24213 23171 24271 23177
rect 24213 23137 24225 23171
rect 24259 23137 24271 23171
rect 24213 23131 24271 23137
rect 24305 23171 24363 23177
rect 24305 23137 24317 23171
rect 24351 23168 24363 23171
rect 24394 23168 24400 23180
rect 24351 23140 24400 23168
rect 24351 23137 24363 23140
rect 24305 23131 24363 23137
rect 24136 23100 24164 23131
rect 23584 23072 24164 23100
rect 24228 23100 24256 23131
rect 24394 23128 24400 23140
rect 24452 23128 24458 23180
rect 25130 23128 25136 23180
rect 25188 23128 25194 23180
rect 25409 23171 25467 23177
rect 25409 23137 25421 23171
rect 25455 23168 25467 23171
rect 25608 23168 25636 23276
rect 25761 23273 25773 23307
rect 25807 23304 25819 23307
rect 26050 23304 26056 23316
rect 25807 23276 26056 23304
rect 25807 23273 25819 23276
rect 25761 23267 25819 23273
rect 26050 23264 26056 23276
rect 26108 23264 26114 23316
rect 26234 23264 26240 23316
rect 26292 23264 26298 23316
rect 25866 23196 25872 23248
rect 25924 23236 25930 23248
rect 25961 23239 26019 23245
rect 25961 23236 25973 23239
rect 25924 23208 25973 23236
rect 25924 23196 25930 23208
rect 25961 23205 25973 23208
rect 26007 23205 26019 23239
rect 25961 23199 26019 23205
rect 26252 23236 26280 23264
rect 26605 23239 26663 23245
rect 26605 23236 26617 23239
rect 26252 23208 26617 23236
rect 26252 23177 26280 23208
rect 26605 23205 26617 23208
rect 26651 23205 26663 23239
rect 26605 23199 26663 23205
rect 25455 23140 25636 23168
rect 26237 23171 26295 23177
rect 25455 23137 25467 23140
rect 25409 23131 25467 23137
rect 26237 23137 26249 23171
rect 26283 23137 26295 23171
rect 26237 23131 26295 23137
rect 26418 23128 26424 23180
rect 26476 23128 26482 23180
rect 26881 23171 26939 23177
rect 26881 23137 26893 23171
rect 26927 23137 26939 23171
rect 26881 23131 26939 23137
rect 24486 23100 24492 23112
rect 24228 23072 24492 23100
rect 15105 22995 15163 23001
rect 18892 23004 20116 23032
rect 14369 22967 14427 22973
rect 14369 22964 14381 22967
rect 13096 22936 14381 22964
rect 14369 22933 14381 22936
rect 14415 22933 14427 22967
rect 14369 22927 14427 22933
rect 15010 22924 15016 22976
rect 15068 22964 15074 22976
rect 18892 22964 18920 23004
rect 15068 22936 18920 22964
rect 15068 22924 15074 22936
rect 18966 22924 18972 22976
rect 19024 22964 19030 22976
rect 19429 22967 19487 22973
rect 19429 22964 19441 22967
rect 19024 22936 19441 22964
rect 19024 22924 19030 22936
rect 19429 22933 19441 22936
rect 19475 22933 19487 22967
rect 21928 22964 21956 23060
rect 23584 22976 23612 23072
rect 24486 23060 24492 23072
rect 24544 23060 24550 23112
rect 24670 23060 24676 23112
rect 24728 23100 24734 23112
rect 25041 23103 25099 23109
rect 25041 23100 25053 23103
rect 24728 23072 25053 23100
rect 24728 23060 24734 23072
rect 25041 23069 25053 23072
rect 25087 23069 25099 23103
rect 25041 23063 25099 23069
rect 25682 23060 25688 23112
rect 25740 23100 25746 23112
rect 26896 23100 26924 23131
rect 25740 23072 26924 23100
rect 25740 23060 25746 23072
rect 26789 23035 26847 23041
rect 26789 23032 26801 23035
rect 25792 23004 26801 23032
rect 23474 22964 23480 22976
rect 21928 22936 23480 22964
rect 19429 22927 19487 22933
rect 23474 22924 23480 22936
rect 23532 22924 23538 22976
rect 23566 22924 23572 22976
rect 23624 22924 23630 22976
rect 24857 22967 24915 22973
rect 24857 22933 24869 22967
rect 24903 22964 24915 22967
rect 25038 22964 25044 22976
rect 24903 22936 25044 22964
rect 24903 22933 24915 22936
rect 24857 22927 24915 22933
rect 25038 22924 25044 22936
rect 25096 22924 25102 22976
rect 25406 22924 25412 22976
rect 25464 22964 25470 22976
rect 25792 22973 25820 23004
rect 26789 23001 26801 23004
rect 26835 23001 26847 23035
rect 26789 22995 26847 23001
rect 25593 22967 25651 22973
rect 25593 22964 25605 22967
rect 25464 22936 25605 22964
rect 25464 22924 25470 22936
rect 25593 22933 25605 22936
rect 25639 22933 25651 22967
rect 25593 22927 25651 22933
rect 25777 22967 25835 22973
rect 25777 22933 25789 22967
rect 25823 22933 25835 22967
rect 25777 22927 25835 22933
rect 26142 22924 26148 22976
rect 26200 22924 26206 22976
rect 26970 22924 26976 22976
rect 27028 22924 27034 22976
rect 552 22874 27416 22896
rect 552 22822 3756 22874
rect 3808 22822 3820 22874
rect 3872 22822 3884 22874
rect 3936 22822 3948 22874
rect 4000 22822 4012 22874
rect 4064 22822 10472 22874
rect 10524 22822 10536 22874
rect 10588 22822 10600 22874
rect 10652 22822 10664 22874
rect 10716 22822 10728 22874
rect 10780 22822 17188 22874
rect 17240 22822 17252 22874
rect 17304 22822 17316 22874
rect 17368 22822 17380 22874
rect 17432 22822 17444 22874
rect 17496 22822 23904 22874
rect 23956 22822 23968 22874
rect 24020 22822 24032 22874
rect 24084 22822 24096 22874
rect 24148 22822 24160 22874
rect 24212 22822 27416 22874
rect 552 22800 27416 22822
rect 2222 22720 2228 22772
rect 2280 22720 2286 22772
rect 2498 22720 2504 22772
rect 2556 22720 2562 22772
rect 2958 22760 2964 22772
rect 2608 22732 2964 22760
rect 2240 22692 2268 22720
rect 2608 22692 2636 22732
rect 2958 22720 2964 22732
rect 3016 22760 3022 22772
rect 4522 22760 4528 22772
rect 3016 22732 4528 22760
rect 3016 22720 3022 22732
rect 4522 22720 4528 22732
rect 4580 22760 4586 22772
rect 5442 22760 5448 22772
rect 4580 22732 5448 22760
rect 4580 22720 4586 22732
rect 5442 22720 5448 22732
rect 5500 22760 5506 22772
rect 6733 22763 6791 22769
rect 6733 22760 6745 22763
rect 5500 22732 6745 22760
rect 5500 22720 5506 22732
rect 6733 22729 6745 22732
rect 6779 22729 6791 22763
rect 6733 22723 6791 22729
rect 8386 22720 8392 22772
rect 8444 22760 8450 22772
rect 9125 22763 9183 22769
rect 9125 22760 9137 22763
rect 8444 22732 9137 22760
rect 8444 22720 8450 22732
rect 9125 22729 9137 22732
rect 9171 22729 9183 22763
rect 9125 22723 9183 22729
rect 11974 22720 11980 22772
rect 12032 22760 12038 22772
rect 12032 22732 13676 22760
rect 12032 22720 12038 22732
rect 2240 22664 2636 22692
rect 2682 22652 2688 22704
rect 2740 22692 2746 22704
rect 2869 22695 2927 22701
rect 2869 22692 2881 22695
rect 2740 22664 2881 22692
rect 2740 22652 2746 22664
rect 2869 22661 2881 22664
rect 2915 22661 2927 22695
rect 2869 22655 2927 22661
rect 4706 22652 4712 22704
rect 4764 22692 4770 22704
rect 4801 22695 4859 22701
rect 4801 22692 4813 22695
rect 4764 22664 4813 22692
rect 4764 22652 4770 22664
rect 4801 22661 4813 22664
rect 4847 22692 4859 22695
rect 6457 22695 6515 22701
rect 4847 22664 5396 22692
rect 4847 22661 4859 22664
rect 4801 22655 4859 22661
rect 842 22584 848 22636
rect 900 22584 906 22636
rect 5169 22627 5227 22633
rect 5169 22624 5181 22627
rect 5000 22596 5181 22624
rect 5000 22568 5028 22596
rect 5169 22593 5181 22596
rect 5215 22593 5227 22627
rect 5169 22587 5227 22593
rect 3418 22516 3424 22568
rect 3476 22516 3482 22568
rect 4982 22516 4988 22568
rect 5040 22516 5046 22568
rect 5074 22516 5080 22568
rect 5132 22516 5138 22568
rect 5368 22565 5396 22664
rect 6457 22661 6469 22695
rect 6503 22661 6515 22695
rect 6457 22655 6515 22661
rect 6181 22627 6239 22633
rect 6181 22593 6193 22627
rect 6227 22624 6239 22627
rect 6270 22624 6276 22636
rect 6227 22596 6276 22624
rect 6227 22593 6239 22596
rect 6181 22587 6239 22593
rect 6270 22584 6276 22596
rect 6328 22584 6334 22636
rect 6472 22624 6500 22655
rect 6638 22652 6644 22704
rect 6696 22692 6702 22704
rect 6696 22664 9352 22692
rect 6696 22652 6702 22664
rect 7926 22624 7932 22636
rect 6472 22596 6960 22624
rect 5261 22559 5319 22565
rect 5261 22556 5273 22559
rect 5184 22528 5273 22556
rect 1112 22491 1170 22497
rect 1112 22457 1124 22491
rect 1158 22488 1170 22491
rect 1210 22488 1216 22500
rect 1158 22460 1216 22488
rect 1158 22457 1170 22460
rect 1112 22451 1170 22457
rect 1210 22448 1216 22460
rect 1268 22448 1274 22500
rect 3688 22491 3746 22497
rect 3688 22457 3700 22491
rect 3734 22457 3746 22491
rect 3688 22451 3746 22457
rect 2314 22380 2320 22432
rect 2372 22380 2378 22432
rect 2501 22423 2559 22429
rect 2501 22389 2513 22423
rect 2547 22420 2559 22423
rect 2774 22420 2780 22432
rect 2547 22392 2780 22420
rect 2547 22389 2559 22392
rect 2501 22383 2559 22389
rect 2774 22380 2780 22392
rect 2832 22420 2838 22432
rect 3142 22420 3148 22432
rect 2832 22392 3148 22420
rect 2832 22380 2838 22392
rect 3142 22380 3148 22392
rect 3200 22380 3206 22432
rect 3602 22380 3608 22432
rect 3660 22420 3666 22432
rect 3712 22420 3740 22451
rect 3660 22392 3740 22420
rect 3660 22380 3666 22392
rect 4890 22380 4896 22432
rect 4948 22380 4954 22432
rect 5092 22420 5120 22516
rect 5184 22500 5212 22528
rect 5261 22525 5273 22528
rect 5307 22525 5319 22559
rect 5261 22519 5319 22525
rect 5353 22559 5411 22565
rect 5353 22525 5365 22559
rect 5399 22556 5411 22559
rect 5534 22556 5540 22568
rect 5399 22528 5540 22556
rect 5399 22525 5411 22528
rect 5353 22519 5411 22525
rect 5534 22516 5540 22528
rect 5592 22516 5598 22568
rect 5810 22516 5816 22568
rect 5868 22516 5874 22568
rect 6089 22559 6147 22565
rect 6089 22525 6101 22559
rect 6135 22556 6147 22559
rect 6135 22528 6592 22556
rect 6135 22525 6147 22528
rect 6089 22519 6147 22525
rect 5166 22448 5172 22500
rect 5224 22448 5230 22500
rect 6270 22448 6276 22500
rect 6328 22497 6334 22500
rect 6328 22491 6356 22497
rect 6344 22457 6356 22491
rect 6328 22451 6356 22457
rect 6328 22448 6334 22451
rect 6564 22432 6592 22528
rect 6932 22488 6960 22596
rect 7392 22596 7932 22624
rect 7006 22516 7012 22568
rect 7064 22516 7070 22568
rect 7098 22516 7104 22568
rect 7156 22556 7162 22568
rect 7285 22559 7343 22565
rect 7285 22556 7297 22559
rect 7156 22528 7297 22556
rect 7156 22516 7162 22528
rect 7285 22525 7297 22528
rect 7331 22525 7343 22559
rect 7285 22519 7343 22525
rect 7392 22497 7420 22596
rect 7926 22584 7932 22596
rect 7984 22584 7990 22636
rect 7469 22559 7527 22565
rect 7469 22525 7481 22559
rect 7515 22525 7527 22559
rect 7469 22519 7527 22525
rect 7561 22559 7619 22565
rect 7561 22525 7573 22559
rect 7607 22556 7619 22559
rect 7742 22556 7748 22568
rect 7607 22528 7748 22556
rect 7607 22525 7619 22528
rect 7561 22519 7619 22525
rect 7377 22491 7435 22497
rect 7377 22488 7389 22491
rect 6932 22460 7389 22488
rect 7377 22457 7389 22460
rect 7423 22457 7435 22491
rect 7484 22488 7512 22519
rect 7742 22516 7748 22528
rect 7800 22516 7806 22568
rect 9324 22565 9352 22664
rect 12066 22652 12072 22704
rect 12124 22692 12130 22704
rect 12124 22664 12664 22692
rect 12124 22652 12130 22664
rect 9493 22627 9551 22633
rect 9493 22593 9505 22627
rect 9539 22624 9551 22627
rect 9858 22624 9864 22636
rect 9539 22596 9864 22624
rect 9539 22593 9551 22596
rect 9493 22587 9551 22593
rect 9858 22584 9864 22596
rect 9916 22624 9922 22636
rect 12434 22624 12440 22636
rect 9916 22596 12440 22624
rect 9916 22584 9922 22596
rect 12434 22584 12440 22596
rect 12492 22584 12498 22636
rect 12636 22633 12664 22664
rect 12621 22627 12679 22633
rect 12621 22593 12633 22627
rect 12667 22593 12679 22627
rect 13648 22624 13676 22732
rect 13722 22720 13728 22772
rect 13780 22760 13786 22772
rect 14001 22763 14059 22769
rect 14001 22760 14013 22763
rect 13780 22732 14013 22760
rect 13780 22720 13786 22732
rect 14001 22729 14013 22732
rect 14047 22729 14059 22763
rect 14001 22723 14059 22729
rect 17034 22720 17040 22772
rect 17092 22760 17098 22772
rect 17221 22763 17279 22769
rect 17221 22760 17233 22763
rect 17092 22732 17233 22760
rect 17092 22720 17098 22732
rect 17221 22729 17233 22732
rect 17267 22729 17279 22763
rect 17221 22723 17279 22729
rect 17862 22720 17868 22772
rect 17920 22720 17926 22772
rect 18690 22720 18696 22772
rect 18748 22760 18754 22772
rect 18785 22763 18843 22769
rect 18785 22760 18797 22763
rect 18748 22732 18797 22760
rect 18748 22720 18754 22732
rect 18785 22729 18797 22732
rect 18831 22729 18843 22763
rect 18785 22723 18843 22729
rect 19521 22763 19579 22769
rect 19521 22729 19533 22763
rect 19567 22760 19579 22763
rect 20438 22760 20444 22772
rect 19567 22732 20444 22760
rect 19567 22729 19579 22732
rect 19521 22723 19579 22729
rect 20438 22720 20444 22732
rect 20496 22720 20502 22772
rect 23845 22763 23903 22769
rect 23845 22760 23857 22763
rect 21284 22732 23857 22760
rect 13909 22695 13967 22701
rect 13909 22661 13921 22695
rect 13955 22692 13967 22695
rect 14274 22692 14280 22704
rect 13955 22664 14280 22692
rect 13955 22661 13967 22664
rect 13909 22655 13967 22661
rect 14274 22652 14280 22664
rect 14332 22652 14338 22704
rect 19334 22692 19340 22704
rect 17052 22664 19340 22692
rect 16485 22627 16543 22633
rect 13648 22596 16436 22624
rect 12621 22587 12679 22593
rect 9309 22559 9367 22565
rect 9309 22525 9321 22559
rect 9355 22525 9367 22559
rect 9309 22519 9367 22525
rect 9585 22559 9643 22565
rect 9585 22525 9597 22559
rect 9631 22525 9643 22559
rect 9585 22519 9643 22525
rect 7834 22488 7840 22500
rect 7484 22460 7840 22488
rect 7377 22451 7435 22457
rect 7834 22448 7840 22460
rect 7892 22448 7898 22500
rect 9600 22488 9628 22519
rect 10042 22516 10048 22568
rect 10100 22556 10106 22568
rect 10229 22559 10287 22565
rect 10229 22556 10241 22559
rect 10100 22528 10241 22556
rect 10100 22516 10106 22528
rect 10229 22525 10241 22528
rect 10275 22525 10287 22559
rect 10229 22519 10287 22525
rect 10870 22516 10876 22568
rect 10928 22516 10934 22568
rect 11606 22516 11612 22568
rect 11664 22556 11670 22568
rect 12529 22559 12587 22565
rect 12529 22556 12541 22559
rect 11664 22528 12541 22556
rect 11664 22516 11670 22528
rect 12529 22525 12541 22528
rect 12575 22525 12587 22559
rect 12529 22519 12587 22525
rect 12713 22559 12771 22565
rect 12713 22525 12725 22559
rect 12759 22525 12771 22559
rect 12713 22519 12771 22525
rect 9950 22488 9956 22500
rect 9600 22460 9956 22488
rect 9950 22448 9956 22460
rect 10008 22488 10014 22500
rect 10888 22488 10916 22516
rect 10008 22460 10916 22488
rect 10980 22460 11284 22488
rect 10008 22448 10014 22460
rect 5626 22420 5632 22432
rect 5092 22392 5632 22420
rect 5626 22380 5632 22392
rect 5684 22380 5690 22432
rect 6546 22380 6552 22432
rect 6604 22380 6610 22432
rect 7101 22423 7159 22429
rect 7101 22389 7113 22423
rect 7147 22420 7159 22423
rect 7466 22420 7472 22432
rect 7147 22392 7472 22420
rect 7147 22389 7159 22392
rect 7101 22383 7159 22389
rect 7466 22380 7472 22392
rect 7524 22380 7530 22432
rect 9674 22380 9680 22432
rect 9732 22380 9738 22432
rect 10318 22380 10324 22432
rect 10376 22420 10382 22432
rect 10980 22420 11008 22460
rect 10376 22392 11008 22420
rect 10376 22380 10382 22392
rect 11054 22380 11060 22432
rect 11112 22380 11118 22432
rect 11256 22420 11284 22460
rect 12434 22448 12440 22500
rect 12492 22488 12498 22500
rect 12728 22488 12756 22519
rect 12894 22516 12900 22568
rect 12952 22516 12958 22568
rect 13814 22516 13820 22568
rect 13872 22556 13878 22568
rect 14001 22559 14059 22565
rect 14001 22556 14013 22559
rect 13872 22528 14013 22556
rect 13872 22516 13878 22528
rect 14001 22525 14013 22528
rect 14047 22525 14059 22559
rect 14001 22519 14059 22525
rect 14093 22559 14151 22565
rect 14093 22525 14105 22559
rect 14139 22556 14151 22559
rect 14642 22556 14648 22568
rect 14139 22528 14648 22556
rect 14139 22525 14151 22528
rect 14093 22519 14151 22525
rect 14642 22516 14648 22528
rect 14700 22516 14706 22568
rect 15010 22516 15016 22568
rect 15068 22516 15074 22568
rect 12492 22460 12756 22488
rect 12492 22448 12498 22460
rect 13446 22448 13452 22500
rect 13504 22488 13510 22500
rect 13541 22491 13599 22497
rect 13541 22488 13553 22491
rect 13504 22460 13553 22488
rect 13504 22448 13510 22460
rect 13541 22457 13553 22460
rect 13587 22457 13599 22491
rect 13541 22451 13599 22457
rect 14277 22491 14335 22497
rect 14277 22457 14289 22491
rect 14323 22488 14335 22491
rect 14550 22488 14556 22500
rect 14323 22460 14556 22488
rect 14323 22457 14335 22460
rect 14277 22451 14335 22457
rect 14550 22448 14556 22460
rect 14608 22488 14614 22500
rect 15028 22488 15056 22516
rect 14608 22460 15056 22488
rect 16408 22488 16436 22596
rect 16485 22593 16497 22627
rect 16531 22624 16543 22627
rect 16574 22624 16580 22636
rect 16531 22596 16580 22624
rect 16531 22593 16543 22596
rect 16485 22587 16543 22593
rect 16574 22584 16580 22596
rect 16632 22584 16638 22636
rect 17052 22488 17080 22664
rect 19334 22652 19340 22664
rect 19392 22692 19398 22704
rect 19392 22664 19840 22692
rect 19392 22652 19398 22664
rect 17129 22627 17187 22633
rect 17129 22593 17141 22627
rect 17175 22624 17187 22627
rect 18230 22624 18236 22636
rect 17175 22596 17816 22624
rect 17175 22593 17187 22596
rect 17129 22587 17187 22593
rect 17402 22516 17408 22568
rect 17460 22556 17466 22568
rect 17788 22565 17816 22596
rect 18156 22596 18236 22624
rect 17773 22559 17831 22565
rect 17460 22528 17724 22556
rect 17460 22516 17466 22528
rect 17497 22491 17555 22497
rect 17497 22488 17509 22491
rect 16408 22460 17509 22488
rect 14608 22448 14614 22460
rect 17497 22457 17509 22460
rect 17543 22457 17555 22491
rect 17497 22451 17555 22457
rect 17589 22491 17647 22497
rect 17589 22457 17601 22491
rect 17635 22457 17647 22491
rect 17696 22488 17724 22528
rect 17773 22525 17785 22559
rect 17819 22525 17831 22559
rect 17773 22519 17831 22525
rect 17862 22516 17868 22568
rect 17920 22556 17926 22568
rect 18156 22565 18184 22596
rect 18230 22584 18236 22596
rect 18288 22584 18294 22636
rect 18966 22624 18972 22636
rect 18432 22596 18972 22624
rect 18432 22565 18460 22596
rect 18966 22584 18972 22596
rect 19024 22584 19030 22636
rect 19812 22624 19840 22664
rect 19812 22596 19932 22624
rect 18049 22559 18107 22565
rect 18049 22556 18061 22559
rect 17920 22528 18061 22556
rect 17920 22516 17926 22528
rect 18049 22525 18061 22528
rect 18095 22525 18107 22559
rect 18049 22519 18107 22525
rect 18141 22559 18199 22565
rect 18141 22525 18153 22559
rect 18187 22525 18199 22559
rect 18141 22519 18199 22525
rect 18417 22559 18475 22565
rect 18417 22525 18429 22559
rect 18463 22525 18475 22559
rect 18417 22519 18475 22525
rect 18877 22559 18935 22565
rect 18877 22525 18889 22559
rect 18923 22525 18935 22559
rect 18877 22519 18935 22525
rect 17880 22488 17908 22516
rect 17696 22460 17908 22488
rect 18233 22491 18291 22497
rect 17589 22451 17647 22457
rect 18233 22457 18245 22491
rect 18279 22457 18291 22491
rect 18892 22488 18920 22519
rect 19058 22516 19064 22568
rect 19116 22516 19122 22568
rect 19150 22516 19156 22568
rect 19208 22516 19214 22568
rect 19334 22516 19340 22568
rect 19392 22516 19398 22568
rect 19426 22516 19432 22568
rect 19484 22556 19490 22568
rect 19797 22559 19855 22565
rect 19797 22556 19809 22559
rect 19484 22528 19809 22556
rect 19484 22516 19490 22528
rect 19797 22525 19809 22528
rect 19843 22525 19855 22559
rect 19904 22556 19932 22596
rect 21284 22565 21312 22732
rect 23845 22729 23857 22732
rect 23891 22729 23903 22763
rect 23845 22723 23903 22729
rect 24946 22720 24952 22772
rect 25004 22760 25010 22772
rect 25225 22763 25283 22769
rect 25225 22760 25237 22763
rect 25004 22732 25237 22760
rect 25004 22720 25010 22732
rect 25225 22729 25237 22732
rect 25271 22729 25283 22763
rect 25225 22723 25283 22729
rect 25590 22720 25596 22772
rect 25648 22720 25654 22772
rect 25682 22720 25688 22772
rect 25740 22720 25746 22772
rect 23293 22695 23351 22701
rect 23293 22661 23305 22695
rect 23339 22692 23351 22695
rect 23566 22692 23572 22704
rect 23339 22664 23572 22692
rect 23339 22661 23351 22664
rect 23293 22655 23351 22661
rect 23566 22652 23572 22664
rect 23624 22652 23630 22704
rect 24394 22652 24400 22704
rect 24452 22692 24458 22704
rect 24854 22692 24860 22704
rect 24452 22664 24860 22692
rect 24452 22652 24458 22664
rect 24854 22652 24860 22664
rect 24912 22652 24918 22704
rect 21910 22584 21916 22636
rect 21968 22584 21974 22636
rect 25498 22584 25504 22636
rect 25556 22584 25562 22636
rect 21269 22559 21327 22565
rect 19904 22528 20208 22556
rect 19797 22519 19855 22525
rect 19242 22488 19248 22500
rect 18892 22460 19248 22488
rect 18233 22451 18291 22457
rect 13170 22420 13176 22432
rect 11256 22392 13176 22420
rect 13170 22380 13176 22392
rect 13228 22380 13234 22432
rect 13630 22380 13636 22432
rect 13688 22420 13694 22432
rect 13741 22423 13799 22429
rect 13741 22420 13753 22423
rect 13688 22392 13753 22420
rect 13688 22380 13694 22392
rect 13741 22389 13753 22392
rect 13787 22389 13799 22423
rect 13741 22383 13799 22389
rect 16666 22380 16672 22432
rect 16724 22420 16730 22432
rect 17034 22420 17040 22432
rect 16724 22392 17040 22420
rect 16724 22380 16730 22392
rect 17034 22380 17040 22392
rect 17092 22380 17098 22432
rect 17604 22420 17632 22451
rect 17678 22420 17684 22432
rect 17604 22392 17684 22420
rect 17678 22380 17684 22392
rect 17736 22420 17742 22432
rect 18248 22420 18276 22451
rect 19242 22448 19248 22460
rect 19300 22448 19306 22500
rect 19886 22448 19892 22500
rect 19944 22488 19950 22500
rect 20042 22491 20100 22497
rect 20042 22488 20054 22491
rect 19944 22460 20054 22488
rect 19944 22448 19950 22460
rect 20042 22457 20054 22460
rect 20088 22457 20100 22491
rect 20180 22488 20208 22528
rect 21269 22525 21281 22559
rect 21315 22525 21327 22559
rect 21545 22559 21603 22565
rect 21545 22556 21557 22559
rect 21269 22519 21327 22525
rect 21376 22528 21557 22556
rect 21376 22500 21404 22528
rect 21545 22525 21557 22528
rect 21591 22525 21603 22559
rect 21545 22519 21603 22525
rect 21634 22516 21640 22568
rect 21692 22516 21698 22568
rect 24397 22559 24455 22565
rect 24397 22525 24409 22559
rect 24443 22525 24455 22559
rect 24397 22519 24455 22525
rect 21358 22488 21364 22500
rect 20180 22460 21364 22488
rect 20042 22451 20100 22457
rect 21358 22448 21364 22460
rect 21416 22448 21422 22500
rect 21450 22448 21456 22500
rect 21508 22448 21514 22500
rect 22158 22491 22216 22497
rect 22158 22488 22170 22491
rect 22066 22460 22170 22488
rect 17736 22392 18276 22420
rect 21177 22423 21235 22429
rect 17736 22380 17742 22392
rect 21177 22389 21189 22423
rect 21223 22420 21235 22423
rect 21726 22420 21732 22432
rect 21223 22392 21732 22420
rect 21223 22389 21235 22392
rect 21177 22383 21235 22389
rect 21726 22380 21732 22392
rect 21784 22380 21790 22432
rect 21821 22423 21879 22429
rect 21821 22389 21833 22423
rect 21867 22420 21879 22423
rect 22066 22420 22094 22460
rect 22158 22457 22170 22460
rect 22204 22457 22216 22491
rect 22158 22451 22216 22457
rect 23566 22448 23572 22500
rect 23624 22488 23630 22500
rect 24412 22488 24440 22519
rect 24578 22516 24584 22568
rect 24636 22516 24642 22568
rect 24765 22559 24823 22565
rect 24765 22556 24777 22559
rect 24688 22528 24777 22556
rect 24688 22500 24716 22528
rect 24765 22525 24777 22528
rect 24811 22525 24823 22559
rect 24765 22519 24823 22525
rect 24854 22516 24860 22568
rect 24912 22516 24918 22568
rect 24949 22559 25007 22565
rect 24949 22525 24961 22559
rect 24995 22525 25007 22559
rect 24949 22519 25007 22525
rect 23624 22460 24440 22488
rect 23624 22448 23630 22460
rect 24670 22448 24676 22500
rect 24728 22448 24734 22500
rect 24964 22488 24992 22519
rect 25406 22516 25412 22568
rect 25464 22516 25470 22568
rect 25516 22556 25544 22584
rect 26510 22556 26516 22568
rect 25516 22528 26516 22556
rect 26510 22516 26516 22528
rect 26568 22556 26574 22568
rect 27065 22559 27123 22565
rect 27065 22556 27077 22559
rect 26568 22528 27077 22556
rect 26568 22516 26574 22528
rect 27065 22525 27077 22528
rect 27111 22525 27123 22559
rect 27065 22519 27123 22525
rect 26142 22488 26148 22500
rect 24964 22460 26148 22488
rect 21867 22392 22094 22420
rect 21867 22389 21879 22392
rect 21821 22383 21879 22389
rect 24486 22380 24492 22432
rect 24544 22420 24550 22432
rect 24964 22420 24992 22460
rect 26142 22448 26148 22460
rect 26200 22448 26206 22500
rect 26786 22448 26792 22500
rect 26844 22497 26850 22500
rect 26844 22451 26856 22497
rect 26844 22448 26850 22451
rect 24544 22392 24992 22420
rect 24544 22380 24550 22392
rect 552 22330 27576 22352
rect 552 22278 7114 22330
rect 7166 22278 7178 22330
rect 7230 22278 7242 22330
rect 7294 22278 7306 22330
rect 7358 22278 7370 22330
rect 7422 22278 13830 22330
rect 13882 22278 13894 22330
rect 13946 22278 13958 22330
rect 14010 22278 14022 22330
rect 14074 22278 14086 22330
rect 14138 22278 20546 22330
rect 20598 22278 20610 22330
rect 20662 22278 20674 22330
rect 20726 22278 20738 22330
rect 20790 22278 20802 22330
rect 20854 22278 27262 22330
rect 27314 22278 27326 22330
rect 27378 22278 27390 22330
rect 27442 22278 27454 22330
rect 27506 22278 27518 22330
rect 27570 22278 27576 22330
rect 552 22256 27576 22278
rect 1210 22176 1216 22228
rect 1268 22176 1274 22228
rect 2314 22216 2320 22228
rect 1780 22188 2320 22216
rect 1397 22083 1455 22089
rect 1397 22049 1409 22083
rect 1443 22080 1455 22083
rect 1780 22080 1808 22188
rect 2314 22176 2320 22188
rect 2372 22176 2378 22228
rect 2409 22219 2467 22225
rect 2409 22185 2421 22219
rect 2455 22216 2467 22219
rect 2498 22216 2504 22228
rect 2455 22188 2504 22216
rect 2455 22185 2467 22188
rect 2409 22179 2467 22185
rect 2498 22176 2504 22188
rect 2556 22176 2562 22228
rect 2958 22216 2964 22228
rect 2608 22188 2964 22216
rect 2608 22157 2636 22188
rect 2958 22176 2964 22188
rect 3016 22176 3022 22228
rect 3142 22176 3148 22228
rect 3200 22216 3206 22228
rect 3881 22219 3939 22225
rect 3881 22216 3893 22219
rect 3200 22188 3893 22216
rect 3200 22176 3206 22188
rect 3881 22185 3893 22188
rect 3927 22185 3939 22219
rect 3881 22179 3939 22185
rect 4062 22176 4068 22228
rect 4120 22176 4126 22228
rect 5629 22219 5687 22225
rect 5629 22185 5641 22219
rect 5675 22216 5687 22219
rect 5810 22216 5816 22228
rect 5675 22188 5816 22216
rect 5675 22185 5687 22188
rect 5629 22179 5687 22185
rect 5810 22176 5816 22188
rect 5868 22216 5874 22228
rect 5868 22188 6132 22216
rect 5868 22176 5874 22188
rect 2593 22151 2651 22157
rect 2593 22117 2605 22151
rect 2639 22117 2651 22151
rect 2593 22111 2651 22117
rect 2777 22151 2835 22157
rect 2777 22117 2789 22151
rect 2823 22148 2835 22151
rect 2866 22148 2872 22160
rect 2823 22120 2872 22148
rect 2823 22117 2835 22120
rect 2777 22111 2835 22117
rect 2866 22108 2872 22120
rect 2924 22148 2930 22160
rect 2924 22120 3556 22148
rect 2924 22108 2930 22120
rect 3528 22089 3556 22120
rect 1443 22052 1808 22080
rect 3513 22083 3571 22089
rect 1443 22049 1455 22052
rect 1397 22043 1455 22049
rect 3513 22049 3525 22083
rect 3559 22080 3571 22083
rect 5169 22083 5227 22089
rect 3559 22052 3593 22080
rect 3559 22049 3571 22052
rect 3513 22043 3571 22049
rect 5169 22049 5181 22083
rect 5215 22049 5227 22083
rect 5169 22043 5227 22049
rect 5184 22012 5212 22043
rect 5534 22040 5540 22092
rect 5592 22080 5598 22092
rect 5813 22083 5871 22089
rect 5813 22080 5825 22083
rect 5592 22052 5825 22080
rect 5592 22040 5598 22052
rect 5813 22049 5825 22052
rect 5859 22049 5871 22083
rect 5813 22043 5871 22049
rect 5994 22012 6000 22024
rect 5184 21984 6000 22012
rect 5994 21972 6000 21984
rect 6052 21972 6058 22024
rect 6104 22012 6132 22188
rect 6270 22176 6276 22228
rect 6328 22176 6334 22228
rect 6362 22176 6368 22228
rect 6420 22176 6426 22228
rect 6457 22219 6515 22225
rect 6457 22185 6469 22219
rect 6503 22216 6515 22219
rect 6546 22216 6552 22228
rect 6503 22188 6552 22216
rect 6503 22185 6515 22188
rect 6457 22179 6515 22185
rect 6546 22176 6552 22188
rect 6604 22176 6610 22228
rect 7466 22176 7472 22228
rect 7524 22176 7530 22228
rect 7561 22219 7619 22225
rect 7561 22185 7573 22219
rect 7607 22216 7619 22219
rect 7650 22216 7656 22228
rect 7607 22188 7656 22216
rect 7607 22185 7619 22188
rect 7561 22179 7619 22185
rect 7650 22176 7656 22188
rect 7708 22176 7714 22228
rect 10134 22176 10140 22228
rect 10192 22176 10198 22228
rect 12802 22176 12808 22228
rect 12860 22176 12866 22228
rect 14553 22219 14611 22225
rect 14553 22185 14565 22219
rect 14599 22216 14611 22219
rect 14642 22216 14648 22228
rect 14599 22188 14648 22216
rect 14599 22185 14611 22188
rect 14553 22179 14611 22185
rect 14642 22176 14648 22188
rect 14700 22176 14706 22228
rect 16574 22176 16580 22228
rect 16632 22216 16638 22228
rect 17678 22216 17684 22228
rect 16632 22188 17684 22216
rect 16632 22176 16638 22188
rect 17678 22176 17684 22188
rect 17736 22216 17742 22228
rect 17736 22188 18092 22216
rect 17736 22176 17742 22188
rect 6380 22089 6408 22176
rect 6365 22083 6423 22089
rect 6365 22049 6377 22083
rect 6411 22049 6423 22083
rect 6365 22043 6423 22049
rect 6641 22083 6699 22089
rect 6641 22049 6653 22083
rect 6687 22049 6699 22083
rect 6641 22043 6699 22049
rect 6656 22012 6684 22043
rect 6730 22040 6736 22092
rect 6788 22080 6794 22092
rect 7484 22089 7512 22176
rect 11238 22108 11244 22160
rect 11296 22148 11302 22160
rect 18064 22157 18092 22188
rect 19150 22176 19156 22228
rect 19208 22216 19214 22228
rect 19208 22188 19472 22216
rect 19208 22176 19214 22188
rect 11670 22151 11728 22157
rect 11670 22148 11682 22151
rect 11296 22120 11682 22148
rect 11296 22108 11302 22120
rect 11670 22117 11682 22120
rect 11716 22117 11728 22151
rect 18049 22151 18107 22157
rect 11670 22111 11728 22117
rect 15580 22120 15976 22148
rect 7101 22083 7159 22089
rect 7101 22080 7113 22083
rect 6788 22052 7113 22080
rect 6788 22040 6794 22052
rect 7101 22049 7113 22052
rect 7147 22049 7159 22083
rect 7101 22043 7159 22049
rect 7469 22083 7527 22089
rect 7469 22049 7481 22083
rect 7515 22049 7527 22083
rect 7469 22043 7527 22049
rect 7558 22040 7564 22092
rect 7616 22040 7622 22092
rect 7742 22040 7748 22092
rect 7800 22040 7806 22092
rect 7926 22040 7932 22092
rect 7984 22040 7990 22092
rect 8754 22040 8760 22092
rect 8812 22080 8818 22092
rect 8921 22083 8979 22089
rect 8921 22080 8933 22083
rect 8812 22052 8933 22080
rect 8812 22040 8818 22052
rect 8921 22049 8933 22052
rect 8967 22049 8979 22083
rect 8921 22043 8979 22049
rect 11054 22040 11060 22092
rect 11112 22080 11118 22092
rect 11422 22080 11428 22092
rect 11112 22052 11428 22080
rect 11112 22040 11118 22052
rect 11422 22040 11428 22052
rect 11480 22040 11486 22092
rect 14182 22040 14188 22092
rect 14240 22089 14246 22092
rect 14240 22043 14252 22089
rect 15580 22080 15608 22120
rect 15948 22089 15976 22120
rect 16132 22120 17172 22148
rect 14936 22052 15608 22080
rect 15677 22083 15735 22089
rect 14240 22040 14246 22043
rect 6104 21984 6684 22012
rect 7006 21972 7012 22024
rect 7064 22012 7070 22024
rect 7285 22015 7343 22021
rect 7064 21984 7236 22012
rect 7064 21972 7070 21984
rect 5442 21904 5448 21956
rect 5500 21904 5506 21956
rect 6638 21904 6644 21956
rect 6696 21904 6702 21956
rect 6914 21904 6920 21956
rect 6972 21944 6978 21956
rect 7101 21947 7159 21953
rect 7101 21944 7113 21947
rect 6972 21916 7113 21944
rect 6972 21904 6978 21916
rect 7101 21913 7113 21916
rect 7147 21913 7159 21947
rect 7208 21944 7236 21984
rect 7285 21981 7297 22015
rect 7331 22012 7343 22015
rect 7576 22012 7604 22040
rect 7331 21984 7604 22012
rect 7331 21981 7343 21984
rect 7285 21975 7343 21981
rect 8018 21972 8024 22024
rect 8076 22012 8082 22024
rect 8665 22015 8723 22021
rect 8665 22012 8677 22015
rect 8076 21984 8677 22012
rect 8076 21972 8082 21984
rect 8665 21981 8677 21984
rect 8711 21981 8723 22015
rect 10689 22015 10747 22021
rect 10689 22012 10701 22015
rect 8665 21975 8723 21981
rect 10152 21984 10701 22012
rect 8202 21944 8208 21956
rect 7208 21916 8208 21944
rect 7101 21907 7159 21913
rect 8202 21904 8208 21916
rect 8260 21904 8266 21956
rect 10042 21904 10048 21956
rect 10100 21904 10106 21956
rect 3881 21879 3939 21885
rect 3881 21845 3893 21879
rect 3927 21876 3939 21879
rect 4890 21876 4896 21888
rect 3927 21848 4896 21876
rect 3927 21845 3939 21848
rect 3881 21839 3939 21845
rect 4890 21836 4896 21848
rect 4948 21836 4954 21888
rect 6086 21836 6092 21888
rect 6144 21876 6150 21888
rect 10060 21876 10088 21904
rect 10152 21888 10180 21984
rect 10689 21981 10701 21984
rect 10735 21981 10747 22015
rect 10689 21975 10747 21981
rect 14461 22015 14519 22021
rect 14461 21981 14473 22015
rect 14507 21981 14519 22015
rect 14461 21975 14519 21981
rect 6144 21848 10088 21876
rect 6144 21836 6150 21848
rect 10134 21836 10140 21888
rect 10192 21836 10198 21888
rect 13081 21879 13139 21885
rect 13081 21845 13093 21879
rect 13127 21876 13139 21879
rect 13814 21876 13820 21888
rect 13127 21848 13820 21876
rect 13127 21845 13139 21848
rect 13081 21839 13139 21845
rect 13814 21836 13820 21848
rect 13872 21836 13878 21888
rect 14476 21876 14504 21975
rect 14936 21876 14964 22052
rect 15677 22049 15689 22083
rect 15723 22080 15735 22083
rect 15933 22083 15991 22089
rect 15723 22052 15884 22080
rect 15723 22049 15735 22052
rect 15677 22043 15735 22049
rect 15856 22012 15884 22052
rect 15933 22049 15945 22083
rect 15979 22080 15991 22083
rect 15979 22052 16013 22080
rect 15979 22049 15991 22052
rect 15933 22043 15991 22049
rect 16132 22024 16160 22120
rect 16393 22083 16451 22089
rect 16393 22049 16405 22083
rect 16439 22049 16451 22083
rect 16393 22043 16451 22049
rect 15856 21984 16068 22012
rect 16040 21944 16068 21984
rect 16114 21972 16120 22024
rect 16172 21972 16178 22024
rect 16298 21972 16304 22024
rect 16356 22012 16362 22024
rect 16408 22012 16436 22043
rect 16574 22040 16580 22092
rect 16632 22040 16638 22092
rect 16666 22040 16672 22092
rect 16724 22040 16730 22092
rect 16850 22040 16856 22092
rect 16908 22040 16914 22092
rect 17144 22089 17172 22120
rect 18049 22117 18061 22151
rect 18095 22117 18107 22151
rect 19168 22148 19196 22176
rect 18049 22111 18107 22117
rect 18708 22120 19196 22148
rect 16945 22083 17003 22089
rect 16945 22049 16957 22083
rect 16991 22049 17003 22083
rect 16945 22043 17003 22049
rect 17129 22083 17187 22089
rect 17129 22049 17141 22083
rect 17175 22080 17187 22083
rect 17175 22052 17632 22080
rect 17175 22049 17187 22052
rect 17129 22043 17187 22049
rect 16356 21984 16436 22012
rect 16356 21972 16362 21984
rect 16761 21947 16819 21953
rect 16761 21944 16773 21947
rect 16040 21916 16773 21944
rect 16761 21913 16773 21916
rect 16807 21913 16819 21947
rect 16761 21907 16819 21913
rect 15746 21876 15752 21888
rect 14476 21848 15752 21876
rect 15746 21836 15752 21848
rect 15804 21836 15810 21888
rect 16206 21836 16212 21888
rect 16264 21876 16270 21888
rect 16960 21876 16988 22043
rect 17037 22015 17095 22021
rect 17037 21981 17049 22015
rect 17083 21981 17095 22015
rect 17037 21975 17095 21981
rect 17052 21944 17080 21975
rect 17402 21944 17408 21956
rect 17052 21916 17408 21944
rect 17402 21904 17408 21916
rect 17460 21904 17466 21956
rect 17604 21944 17632 22052
rect 17770 22040 17776 22092
rect 17828 22080 17834 22092
rect 17865 22083 17923 22089
rect 17865 22080 17877 22083
rect 17828 22052 17877 22080
rect 17828 22040 17834 22052
rect 17865 22049 17877 22052
rect 17911 22049 17923 22083
rect 17865 22043 17923 22049
rect 17957 22083 18015 22089
rect 17957 22049 17969 22083
rect 18003 22049 18015 22083
rect 17957 22043 18015 22049
rect 18233 22083 18291 22089
rect 18233 22049 18245 22083
rect 18279 22080 18291 22083
rect 18601 22083 18659 22089
rect 18601 22080 18613 22083
rect 18279 22052 18613 22080
rect 18279 22049 18291 22052
rect 18233 22043 18291 22049
rect 18601 22049 18613 22052
rect 18647 22049 18659 22083
rect 18601 22043 18659 22049
rect 17972 22012 18000 22043
rect 18708 22024 18736 22120
rect 19058 22040 19064 22092
rect 19116 22080 19122 22092
rect 19444 22089 19472 22188
rect 19610 22176 19616 22228
rect 19668 22176 19674 22228
rect 19886 22176 19892 22228
rect 19944 22176 19950 22228
rect 20346 22176 20352 22228
rect 20404 22216 20410 22228
rect 24486 22216 24492 22228
rect 20404 22188 24492 22216
rect 20404 22176 20410 22188
rect 24486 22176 24492 22188
rect 24544 22176 24550 22228
rect 26786 22176 26792 22228
rect 26844 22216 26850 22228
rect 26881 22219 26939 22225
rect 26881 22216 26893 22219
rect 26844 22188 26893 22216
rect 26844 22176 26850 22188
rect 26881 22185 26893 22188
rect 26927 22185 26939 22219
rect 26881 22179 26939 22185
rect 25866 22148 25872 22160
rect 20057 22120 21680 22148
rect 19429 22083 19487 22089
rect 19116 22052 19380 22080
rect 19116 22040 19122 22052
rect 18046 22012 18052 22024
rect 17972 21984 18052 22012
rect 18046 21972 18052 21984
rect 18104 22012 18110 22024
rect 18506 22012 18512 22024
rect 18104 21984 18512 22012
rect 18104 21972 18110 21984
rect 18506 21972 18512 21984
rect 18564 21972 18570 22024
rect 18690 21972 18696 22024
rect 18748 21972 18754 22024
rect 19242 21972 19248 22024
rect 19300 21972 19306 22024
rect 19352 22012 19380 22052
rect 19429 22049 19441 22083
rect 19475 22080 19487 22083
rect 19613 22083 19671 22089
rect 19475 22052 19509 22080
rect 19475 22049 19487 22052
rect 19429 22043 19487 22049
rect 19613 22049 19625 22083
rect 19659 22049 19671 22083
rect 19613 22043 19671 22049
rect 19628 22012 19656 22043
rect 19886 22040 19892 22092
rect 19944 22080 19950 22092
rect 20057 22089 20085 22120
rect 21652 22092 21680 22120
rect 25700 22120 25872 22148
rect 20049 22083 20107 22089
rect 20049 22080 20061 22083
rect 19944 22052 20061 22080
rect 19944 22040 19950 22052
rect 20049 22049 20061 22052
rect 20095 22049 20107 22083
rect 20049 22043 20107 22049
rect 20165 22083 20223 22089
rect 20165 22049 20177 22083
rect 20211 22049 20223 22083
rect 20165 22043 20223 22049
rect 20257 22083 20315 22089
rect 20257 22049 20269 22083
rect 20303 22049 20315 22083
rect 20257 22043 20315 22049
rect 20441 22083 20499 22089
rect 20441 22049 20453 22083
rect 20487 22080 20499 22083
rect 21269 22083 21327 22089
rect 21269 22080 21281 22083
rect 20487 22052 21281 22080
rect 20487 22049 20499 22052
rect 20441 22043 20499 22049
rect 21269 22049 21281 22052
rect 21315 22049 21327 22083
rect 21269 22043 21327 22049
rect 19352 21984 19656 22012
rect 19150 21944 19156 21956
rect 17604 21916 19156 21944
rect 19150 21904 19156 21916
rect 19208 21904 19214 21956
rect 19978 21904 19984 21956
rect 20036 21944 20042 21956
rect 20184 21944 20212 22043
rect 20272 22012 20300 22043
rect 21358 22040 21364 22092
rect 21416 22040 21422 22092
rect 21450 22040 21456 22092
rect 21508 22040 21514 22092
rect 21634 22040 21640 22092
rect 21692 22040 21698 22092
rect 21726 22040 21732 22092
rect 21784 22080 21790 22092
rect 21821 22083 21879 22089
rect 21821 22080 21833 22083
rect 21784 22052 21833 22080
rect 21784 22040 21790 22052
rect 21821 22049 21833 22052
rect 21867 22080 21879 22083
rect 24394 22080 24400 22092
rect 21867 22052 24400 22080
rect 21867 22049 21879 22052
rect 21821 22043 21879 22049
rect 24394 22040 24400 22052
rect 24452 22040 24458 22092
rect 25700 22089 25728 22120
rect 25866 22108 25872 22120
rect 25924 22148 25930 22160
rect 26421 22151 26479 22157
rect 26421 22148 26433 22151
rect 25924 22120 26433 22148
rect 25924 22108 25930 22120
rect 26421 22117 26433 22120
rect 26467 22117 26479 22151
rect 26421 22111 26479 22117
rect 26637 22151 26695 22157
rect 26637 22117 26649 22151
rect 26683 22148 26695 22151
rect 26970 22148 26976 22160
rect 26683 22120 26976 22148
rect 26683 22117 26695 22120
rect 26637 22111 26695 22117
rect 26970 22108 26976 22120
rect 27028 22108 27034 22160
rect 24857 22083 24915 22089
rect 24857 22049 24869 22083
rect 24903 22080 24915 22083
rect 24949 22083 25007 22089
rect 24949 22080 24961 22083
rect 24903 22052 24961 22080
rect 24903 22049 24915 22052
rect 24857 22043 24915 22049
rect 24949 22049 24961 22052
rect 24995 22049 25007 22083
rect 24949 22043 25007 22049
rect 25685 22083 25743 22089
rect 25685 22049 25697 22083
rect 25731 22049 25743 22083
rect 25685 22043 25743 22049
rect 26053 22083 26111 22089
rect 26053 22049 26065 22083
rect 26099 22049 26111 22083
rect 26053 22043 26111 22049
rect 26145 22083 26203 22089
rect 26145 22049 26157 22083
rect 26191 22080 26203 22083
rect 27065 22083 27123 22089
rect 26191 22052 26464 22080
rect 26191 22049 26203 22052
rect 26145 22043 26203 22049
rect 21376 22012 21404 22040
rect 20272 21984 21404 22012
rect 20898 21944 20904 21956
rect 20036 21916 20904 21944
rect 20036 21904 20042 21916
rect 20898 21904 20904 21916
rect 20956 21904 20962 21956
rect 16264 21848 16988 21876
rect 17681 21879 17739 21885
rect 16264 21836 16270 21848
rect 17681 21845 17693 21879
rect 17727 21876 17739 21879
rect 17862 21876 17868 21888
rect 17727 21848 17868 21876
rect 17727 21845 17739 21848
rect 17681 21839 17739 21845
rect 17862 21836 17868 21848
rect 17920 21836 17926 21888
rect 21082 21836 21088 21888
rect 21140 21876 21146 21888
rect 21468 21876 21496 22040
rect 22922 21972 22928 22024
rect 22980 21972 22986 22024
rect 23566 21972 23572 22024
rect 23624 21972 23630 22024
rect 25498 21972 25504 22024
rect 25556 21972 25562 22024
rect 21818 21904 21824 21956
rect 21876 21944 21882 21956
rect 23017 21947 23075 21953
rect 23017 21944 23029 21947
rect 21876 21916 23029 21944
rect 21876 21904 21882 21916
rect 23017 21913 23029 21916
rect 23063 21913 23075 21947
rect 23017 21907 23075 21913
rect 24394 21904 24400 21956
rect 24452 21944 24458 21956
rect 24765 21947 24823 21953
rect 24765 21944 24777 21947
rect 24452 21916 24777 21944
rect 24452 21904 24458 21916
rect 24765 21913 24777 21916
rect 24811 21944 24823 21947
rect 26068 21944 26096 22043
rect 24811 21916 26096 21944
rect 24811 21913 24823 21916
rect 24765 21907 24823 21913
rect 26436 21888 26464 22052
rect 27065 22049 27077 22083
rect 27111 22049 27123 22083
rect 27065 22043 27123 22049
rect 26789 21947 26847 21953
rect 26789 21913 26801 21947
rect 26835 21944 26847 21947
rect 27080 21944 27108 22043
rect 26835 21916 27108 21944
rect 26835 21913 26847 21916
rect 26789 21907 26847 21913
rect 21140 21848 21496 21876
rect 21140 21836 21146 21848
rect 21542 21836 21548 21888
rect 21600 21876 21606 21888
rect 22281 21879 22339 21885
rect 22281 21876 22293 21879
rect 21600 21848 22293 21876
rect 21600 21836 21606 21848
rect 22281 21845 22293 21848
rect 22327 21845 22339 21879
rect 22281 21839 22339 21845
rect 25866 21836 25872 21888
rect 25924 21836 25930 21888
rect 26418 21836 26424 21888
rect 26476 21876 26482 21888
rect 26605 21879 26663 21885
rect 26605 21876 26617 21879
rect 26476 21848 26617 21876
rect 26476 21836 26482 21848
rect 26605 21845 26617 21848
rect 26651 21845 26663 21879
rect 26605 21839 26663 21845
rect 552 21786 27416 21808
rect 552 21734 3756 21786
rect 3808 21734 3820 21786
rect 3872 21734 3884 21786
rect 3936 21734 3948 21786
rect 4000 21734 4012 21786
rect 4064 21734 10472 21786
rect 10524 21734 10536 21786
rect 10588 21734 10600 21786
rect 10652 21734 10664 21786
rect 10716 21734 10728 21786
rect 10780 21734 17188 21786
rect 17240 21734 17252 21786
rect 17304 21734 17316 21786
rect 17368 21734 17380 21786
rect 17432 21734 17444 21786
rect 17496 21734 23904 21786
rect 23956 21734 23968 21786
rect 24020 21734 24032 21786
rect 24084 21734 24096 21786
rect 24148 21734 24160 21786
rect 24212 21734 27416 21786
rect 552 21712 27416 21734
rect 3786 21672 3792 21684
rect 3528 21644 3792 21672
rect 3528 21616 3556 21644
rect 3786 21632 3792 21644
rect 3844 21672 3850 21684
rect 3881 21675 3939 21681
rect 3881 21672 3893 21675
rect 3844 21644 3893 21672
rect 3844 21632 3850 21644
rect 3881 21641 3893 21644
rect 3927 21641 3939 21675
rect 3881 21635 3939 21641
rect 4249 21675 4307 21681
rect 4249 21641 4261 21675
rect 4295 21672 4307 21675
rect 5258 21672 5264 21684
rect 4295 21644 5264 21672
rect 4295 21641 4307 21644
rect 4249 21635 4307 21641
rect 5258 21632 5264 21644
rect 5316 21632 5322 21684
rect 5994 21632 6000 21684
rect 6052 21672 6058 21684
rect 7006 21672 7012 21684
rect 6052 21644 7012 21672
rect 6052 21632 6058 21644
rect 7006 21632 7012 21644
rect 7064 21632 7070 21684
rect 7742 21632 7748 21684
rect 7800 21632 7806 21684
rect 7837 21675 7895 21681
rect 7837 21641 7849 21675
rect 7883 21641 7895 21675
rect 7837 21635 7895 21641
rect 1305 21607 1363 21613
rect 1305 21573 1317 21607
rect 1351 21604 1363 21607
rect 1351 21576 1624 21604
rect 1351 21573 1363 21576
rect 1305 21567 1363 21573
rect 1489 21539 1547 21545
rect 1489 21536 1501 21539
rect 1044 21508 1501 21536
rect 1044 21477 1072 21508
rect 1489 21505 1501 21508
rect 1535 21505 1547 21539
rect 1489 21499 1547 21505
rect 1596 21480 1624 21576
rect 3510 21564 3516 21616
rect 3568 21564 3574 21616
rect 6917 21607 6975 21613
rect 6917 21573 6929 21607
rect 6963 21604 6975 21607
rect 7760 21604 7788 21632
rect 6963 21576 7788 21604
rect 6963 21573 6975 21576
rect 6917 21567 6975 21573
rect 1673 21539 1731 21545
rect 1673 21505 1685 21539
rect 1719 21536 1731 21539
rect 5166 21536 5172 21548
rect 1719 21508 2452 21536
rect 1719 21505 1731 21508
rect 1673 21499 1731 21505
rect 2424 21480 2452 21508
rect 3528 21508 3924 21536
rect 1029 21471 1087 21477
rect 1029 21437 1041 21471
rect 1075 21437 1087 21471
rect 1397 21471 1455 21477
rect 1397 21468 1409 21471
rect 1029 21431 1087 21437
rect 1228 21440 1409 21468
rect 1044 21344 1072 21431
rect 1026 21292 1032 21344
rect 1084 21292 1090 21344
rect 1121 21335 1179 21341
rect 1121 21301 1133 21335
rect 1167 21332 1179 21335
rect 1228 21332 1256 21440
rect 1397 21437 1409 21440
rect 1443 21437 1455 21471
rect 1397 21431 1455 21437
rect 1578 21428 1584 21480
rect 1636 21428 1642 21480
rect 2222 21428 2228 21480
rect 2280 21468 2286 21480
rect 2317 21471 2375 21477
rect 2317 21468 2329 21471
rect 2280 21440 2329 21468
rect 2280 21428 2286 21440
rect 2317 21437 2329 21440
rect 2363 21437 2375 21471
rect 2317 21431 2375 21437
rect 1305 21403 1363 21409
rect 1305 21369 1317 21403
rect 1351 21400 1363 21403
rect 1673 21403 1731 21409
rect 1673 21400 1685 21403
rect 1351 21372 1685 21400
rect 1351 21369 1363 21372
rect 1305 21363 1363 21369
rect 1673 21369 1685 21372
rect 1719 21369 1731 21403
rect 2332 21400 2360 21431
rect 2406 21428 2412 21480
rect 2464 21428 2470 21480
rect 2501 21471 2559 21477
rect 2501 21437 2513 21471
rect 2547 21468 2559 21471
rect 2774 21468 2780 21480
rect 2547 21440 2780 21468
rect 2547 21437 2559 21440
rect 2501 21431 2559 21437
rect 2774 21428 2780 21440
rect 2832 21428 2838 21480
rect 3418 21428 3424 21480
rect 3476 21468 3482 21480
rect 3528 21477 3556 21508
rect 3513 21471 3571 21477
rect 3513 21468 3525 21471
rect 3476 21440 3525 21468
rect 3476 21428 3482 21440
rect 3513 21437 3525 21440
rect 3559 21437 3571 21471
rect 3513 21431 3571 21437
rect 3786 21428 3792 21480
rect 3844 21428 3850 21480
rect 3896 21477 3924 21508
rect 4908 21508 5172 21536
rect 4908 21477 4936 21508
rect 5166 21496 5172 21508
rect 5224 21536 5230 21548
rect 5534 21536 5540 21548
rect 5224 21508 5540 21536
rect 5224 21496 5230 21508
rect 5534 21496 5540 21508
rect 5592 21496 5598 21548
rect 7742 21496 7748 21548
rect 7800 21536 7806 21548
rect 7852 21536 7880 21635
rect 8202 21632 8208 21684
rect 8260 21632 8266 21684
rect 8754 21632 8760 21684
rect 8812 21632 8818 21684
rect 12069 21675 12127 21681
rect 12069 21641 12081 21675
rect 12115 21672 12127 21675
rect 12250 21672 12256 21684
rect 12115 21644 12256 21672
rect 12115 21641 12127 21644
rect 12069 21635 12127 21641
rect 12250 21632 12256 21644
rect 12308 21632 12314 21684
rect 13630 21632 13636 21684
rect 13688 21632 13694 21684
rect 14182 21632 14188 21684
rect 14240 21632 14246 21684
rect 16025 21675 16083 21681
rect 16025 21641 16037 21675
rect 16071 21672 16083 21675
rect 16666 21672 16672 21684
rect 16071 21644 16672 21672
rect 16071 21641 16083 21644
rect 16025 21635 16083 21641
rect 16666 21632 16672 21644
rect 16724 21632 16730 21684
rect 19334 21672 19340 21684
rect 17144 21644 19340 21672
rect 8220 21604 8248 21632
rect 10045 21607 10103 21613
rect 10045 21604 10057 21607
rect 8220 21576 10057 21604
rect 10045 21573 10057 21576
rect 10091 21604 10103 21607
rect 10134 21604 10140 21616
rect 10091 21576 10140 21604
rect 10091 21573 10103 21576
rect 10045 21567 10103 21573
rect 10134 21564 10140 21576
rect 10192 21564 10198 21616
rect 16206 21604 16212 21616
rect 12912 21576 16212 21604
rect 12912 21548 12940 21576
rect 16206 21564 16212 21576
rect 16264 21564 16270 21616
rect 16298 21564 16304 21616
rect 16356 21604 16362 21616
rect 17144 21604 17172 21644
rect 19334 21632 19340 21644
rect 19392 21632 19398 21684
rect 19886 21632 19892 21684
rect 19944 21632 19950 21684
rect 21542 21632 21548 21684
rect 21600 21632 21606 21684
rect 23566 21632 23572 21684
rect 23624 21632 23630 21684
rect 24489 21675 24547 21681
rect 24489 21641 24501 21675
rect 24535 21672 24547 21675
rect 24670 21672 24676 21684
rect 24535 21644 24676 21672
rect 24535 21641 24547 21644
rect 24489 21635 24547 21641
rect 24670 21632 24676 21644
rect 24728 21632 24734 21684
rect 25041 21675 25099 21681
rect 25041 21641 25053 21675
rect 25087 21672 25099 21675
rect 25130 21672 25136 21684
rect 25087 21644 25136 21672
rect 25087 21641 25099 21644
rect 25041 21635 25099 21641
rect 25130 21632 25136 21644
rect 25188 21632 25194 21684
rect 25498 21632 25504 21684
rect 25556 21632 25562 21684
rect 25682 21632 25688 21684
rect 25740 21632 25746 21684
rect 26510 21632 26516 21684
rect 26568 21672 26574 21684
rect 26605 21675 26663 21681
rect 26605 21672 26617 21675
rect 26568 21644 26617 21672
rect 26568 21632 26574 21644
rect 26605 21641 26617 21644
rect 26651 21641 26663 21675
rect 26605 21635 26663 21641
rect 16356 21576 17172 21604
rect 16356 21564 16362 21576
rect 18322 21564 18328 21616
rect 18380 21604 18386 21616
rect 19058 21604 19064 21616
rect 18380 21576 19064 21604
rect 18380 21564 18386 21576
rect 19058 21564 19064 21576
rect 19116 21604 19122 21616
rect 19245 21607 19303 21613
rect 19245 21604 19257 21607
rect 19116 21576 19257 21604
rect 19116 21564 19122 21576
rect 19245 21573 19257 21576
rect 19291 21604 19303 21607
rect 19291 21576 19932 21604
rect 19291 21573 19303 21576
rect 19245 21567 19303 21573
rect 9582 21536 9588 21548
rect 7800 21508 7880 21536
rect 9140 21508 9588 21536
rect 7800 21496 7806 21508
rect 3881 21471 3939 21477
rect 3881 21437 3893 21471
rect 3927 21437 3939 21471
rect 3881 21431 3939 21437
rect 3973 21471 4031 21477
rect 3973 21437 3985 21471
rect 4019 21437 4031 21471
rect 3973 21431 4031 21437
rect 4893 21471 4951 21477
rect 4893 21437 4905 21471
rect 4939 21437 4951 21471
rect 4893 21431 4951 21437
rect 3697 21403 3755 21409
rect 3697 21400 3709 21403
rect 2332 21372 3709 21400
rect 1673 21363 1731 21369
rect 3697 21369 3709 21372
rect 3743 21400 3755 21403
rect 3988 21400 4016 21431
rect 4982 21428 4988 21480
rect 5040 21428 5046 21480
rect 7006 21428 7012 21480
rect 7064 21468 7070 21480
rect 7101 21471 7159 21477
rect 7101 21468 7113 21471
rect 7064 21440 7113 21468
rect 7064 21428 7070 21440
rect 7101 21437 7113 21440
rect 7147 21437 7159 21471
rect 7101 21431 7159 21437
rect 7377 21471 7435 21477
rect 7377 21437 7389 21471
rect 7423 21468 7435 21471
rect 7929 21471 7987 21477
rect 7423 21440 7696 21468
rect 7423 21437 7435 21440
rect 7377 21431 7435 21437
rect 3743 21372 4016 21400
rect 5169 21403 5227 21409
rect 3743 21369 3755 21372
rect 3697 21363 3755 21369
rect 5169 21369 5181 21403
rect 5215 21400 5227 21403
rect 5442 21400 5448 21412
rect 5215 21372 5448 21400
rect 5215 21369 5227 21372
rect 5169 21363 5227 21369
rect 5442 21360 5448 21372
rect 5500 21360 5506 21412
rect 7285 21403 7343 21409
rect 7285 21369 7297 21403
rect 7331 21400 7343 21403
rect 7558 21400 7564 21412
rect 7331 21372 7564 21400
rect 7331 21369 7343 21372
rect 7285 21363 7343 21369
rect 7558 21360 7564 21372
rect 7616 21360 7622 21412
rect 7668 21344 7696 21440
rect 7929 21437 7941 21471
rect 7975 21437 7987 21471
rect 7929 21431 7987 21437
rect 7944 21344 7972 21431
rect 8846 21428 8852 21480
rect 8904 21468 8910 21480
rect 9140 21477 9168 21508
rect 9582 21496 9588 21508
rect 9640 21536 9646 21548
rect 10226 21536 10232 21548
rect 9640 21508 10232 21536
rect 9640 21496 9646 21508
rect 10226 21496 10232 21508
rect 10284 21536 10290 21548
rect 10410 21536 10416 21548
rect 10284 21508 10416 21536
rect 10284 21496 10290 21508
rect 10410 21496 10416 21508
rect 10468 21496 10474 21548
rect 12894 21496 12900 21548
rect 12952 21496 12958 21548
rect 14642 21536 14648 21548
rect 14016 21508 14648 21536
rect 8941 21471 8999 21477
rect 8941 21468 8953 21471
rect 8904 21440 8953 21468
rect 8904 21428 8910 21440
rect 8941 21437 8953 21440
rect 8987 21437 8999 21471
rect 8941 21431 8999 21437
rect 9125 21471 9183 21477
rect 9125 21437 9137 21471
rect 9171 21437 9183 21471
rect 9125 21431 9183 21437
rect 9309 21471 9367 21477
rect 9309 21437 9321 21471
rect 9355 21468 9367 21471
rect 9674 21468 9680 21480
rect 9355 21440 9680 21468
rect 9355 21437 9367 21440
rect 9309 21431 9367 21437
rect 9674 21428 9680 21440
rect 9732 21428 9738 21480
rect 11146 21428 11152 21480
rect 11204 21477 11210 21480
rect 11204 21431 11216 21477
rect 11204 21428 11210 21431
rect 11422 21428 11428 21480
rect 11480 21468 11486 21480
rect 11790 21468 11796 21480
rect 11480 21440 11796 21468
rect 11480 21428 11486 21440
rect 11790 21428 11796 21440
rect 11848 21428 11854 21480
rect 12253 21471 12311 21477
rect 12253 21437 12265 21471
rect 12299 21437 12311 21471
rect 12253 21431 12311 21437
rect 9033 21403 9091 21409
rect 9033 21369 9045 21403
rect 9079 21400 9091 21403
rect 9214 21400 9220 21412
rect 9079 21372 9220 21400
rect 9079 21369 9091 21372
rect 9033 21363 9091 21369
rect 9214 21360 9220 21372
rect 9272 21400 9278 21412
rect 9858 21400 9864 21412
rect 9272 21372 9864 21400
rect 9272 21360 9278 21372
rect 9858 21360 9864 21372
rect 9916 21400 9922 21412
rect 10962 21400 10968 21412
rect 9916 21372 10968 21400
rect 9916 21360 9922 21372
rect 10962 21360 10968 21372
rect 11020 21360 11026 21412
rect 12268 21400 12296 21431
rect 12434 21428 12440 21480
rect 12492 21428 12498 21480
rect 12529 21471 12587 21477
rect 12529 21437 12541 21471
rect 12575 21468 12587 21471
rect 12912 21468 12940 21496
rect 12575 21440 12940 21468
rect 12575 21437 12587 21440
rect 12529 21431 12587 21437
rect 13814 21428 13820 21480
rect 13872 21428 13878 21480
rect 14016 21477 14044 21508
rect 14642 21496 14648 21508
rect 14700 21536 14706 21548
rect 14829 21539 14887 21545
rect 14829 21536 14841 21539
rect 14700 21508 14841 21536
rect 14700 21496 14706 21508
rect 14829 21505 14841 21508
rect 14875 21505 14887 21539
rect 14829 21499 14887 21505
rect 15841 21539 15899 21545
rect 15841 21505 15853 21539
rect 15887 21536 15899 21539
rect 15887 21508 16988 21536
rect 15887 21505 15899 21508
rect 15841 21499 15899 21505
rect 14001 21471 14059 21477
rect 14001 21437 14013 21471
rect 14047 21437 14059 21471
rect 14001 21431 14059 21437
rect 14093 21471 14151 21477
rect 14093 21437 14105 21471
rect 14139 21437 14151 21471
rect 14093 21431 14151 21437
rect 12802 21400 12808 21412
rect 12268 21372 12808 21400
rect 12802 21360 12808 21372
rect 12860 21360 12866 21412
rect 14108 21400 14136 21431
rect 14366 21428 14372 21480
rect 14424 21428 14430 21480
rect 15473 21471 15531 21477
rect 15473 21437 15485 21471
rect 15519 21468 15531 21471
rect 15749 21471 15807 21477
rect 15749 21468 15761 21471
rect 15519 21440 15761 21468
rect 15519 21437 15531 21440
rect 15473 21431 15531 21437
rect 15749 21437 15761 21440
rect 15795 21437 15807 21471
rect 15749 21431 15807 21437
rect 14182 21400 14188 21412
rect 14108 21372 14188 21400
rect 14182 21360 14188 21372
rect 14240 21400 14246 21412
rect 15856 21400 15884 21499
rect 14240 21372 15884 21400
rect 14240 21360 14246 21372
rect 1765 21335 1823 21341
rect 1765 21332 1777 21335
rect 1167 21304 1777 21332
rect 1167 21301 1179 21304
rect 1121 21295 1179 21301
rect 1765 21301 1777 21304
rect 1811 21301 1823 21335
rect 1765 21295 1823 21301
rect 2682 21292 2688 21344
rect 2740 21292 2746 21344
rect 3326 21292 3332 21344
rect 3384 21292 3390 21344
rect 4890 21292 4896 21344
rect 4948 21292 4954 21344
rect 7466 21292 7472 21344
rect 7524 21292 7530 21344
rect 7650 21292 7656 21344
rect 7708 21292 7714 21344
rect 7926 21292 7932 21344
rect 7984 21292 7990 21344
rect 12820 21332 12848 21360
rect 14274 21332 14280 21344
rect 12820 21304 14280 21332
rect 14274 21292 14280 21304
rect 14332 21292 14338 21344
rect 14366 21292 14372 21344
rect 14424 21332 14430 21344
rect 16114 21332 16120 21344
rect 14424 21304 16120 21332
rect 14424 21292 14430 21304
rect 16114 21292 16120 21304
rect 16172 21292 16178 21344
rect 16669 21335 16727 21341
rect 16669 21301 16681 21335
rect 16715 21332 16727 21335
rect 16850 21332 16856 21344
rect 16715 21304 16856 21332
rect 16715 21301 16727 21304
rect 16669 21295 16727 21301
rect 16850 21292 16856 21304
rect 16908 21292 16914 21344
rect 16960 21332 16988 21508
rect 19150 21496 19156 21548
rect 19208 21536 19214 21548
rect 19208 21508 19748 21536
rect 19208 21496 19214 21508
rect 17954 21428 17960 21480
rect 18012 21468 18018 21480
rect 18049 21471 18107 21477
rect 18049 21468 18061 21471
rect 18012 21440 18061 21468
rect 18012 21428 18018 21440
rect 18049 21437 18061 21440
rect 18095 21437 18107 21471
rect 18049 21431 18107 21437
rect 19334 21428 19340 21480
rect 19392 21468 19398 21480
rect 19720 21477 19748 21508
rect 19904 21477 19932 21576
rect 21560 21536 21588 21632
rect 23201 21607 23259 21613
rect 23201 21573 23213 21607
rect 23247 21604 23259 21607
rect 23584 21604 23612 21632
rect 23247 21576 23612 21604
rect 23247 21573 23259 21576
rect 23201 21567 23259 21573
rect 23584 21536 23612 21576
rect 24949 21607 25007 21613
rect 24949 21573 24961 21607
rect 24995 21604 25007 21607
rect 25516 21604 25544 21632
rect 24995 21576 25544 21604
rect 24995 21573 25007 21576
rect 24949 21567 25007 21573
rect 21192 21508 21588 21536
rect 23492 21508 23612 21536
rect 23937 21539 23995 21545
rect 21192 21477 21220 21508
rect 19429 21471 19487 21477
rect 19429 21468 19441 21471
rect 19392 21440 19441 21468
rect 19392 21428 19398 21440
rect 19429 21437 19441 21440
rect 19475 21437 19487 21471
rect 19429 21431 19487 21437
rect 19705 21471 19763 21477
rect 19705 21437 19717 21471
rect 19751 21437 19763 21471
rect 19705 21431 19763 21437
rect 19889 21471 19947 21477
rect 19889 21437 19901 21471
rect 19935 21437 19947 21471
rect 19889 21431 19947 21437
rect 21177 21471 21235 21477
rect 21177 21437 21189 21471
rect 21223 21437 21235 21471
rect 21177 21431 21235 21437
rect 21358 21428 21364 21480
rect 21416 21428 21422 21480
rect 21545 21471 21603 21477
rect 21545 21437 21557 21471
rect 21591 21468 21603 21471
rect 21634 21468 21640 21480
rect 21591 21440 21640 21468
rect 21591 21437 21603 21440
rect 21545 21431 21603 21437
rect 21634 21428 21640 21440
rect 21692 21428 21698 21480
rect 23492 21477 23520 21508
rect 23937 21505 23949 21539
rect 23983 21536 23995 21539
rect 24026 21536 24032 21548
rect 23983 21508 24032 21536
rect 23983 21505 23995 21508
rect 23937 21499 23995 21505
rect 24026 21496 24032 21508
rect 24084 21536 24090 21548
rect 25700 21536 25728 21632
rect 24084 21508 25728 21536
rect 24084 21496 24090 21508
rect 21821 21471 21879 21477
rect 21821 21437 21833 21471
rect 21867 21437 21879 21471
rect 21821 21431 21879 21437
rect 23477 21471 23535 21477
rect 23477 21437 23489 21471
rect 23523 21437 23535 21471
rect 23477 21431 23535 21437
rect 23569 21471 23627 21477
rect 23569 21437 23581 21471
rect 23615 21468 23627 21471
rect 23842 21468 23848 21480
rect 23615 21440 23848 21468
rect 23615 21437 23627 21440
rect 23569 21431 23627 21437
rect 17804 21403 17862 21409
rect 17804 21369 17816 21403
rect 17850 21400 17862 21403
rect 18138 21400 18144 21412
rect 17850 21372 18144 21400
rect 17850 21369 17862 21372
rect 17804 21363 17862 21369
rect 18138 21360 18144 21372
rect 18196 21360 18202 21412
rect 19613 21403 19671 21409
rect 19613 21369 19625 21403
rect 19659 21400 19671 21403
rect 21376 21400 21404 21428
rect 19659 21372 21404 21400
rect 21453 21403 21511 21409
rect 19659 21369 19671 21372
rect 19613 21363 19671 21369
rect 21453 21369 21465 21403
rect 21499 21369 21511 21403
rect 21453 21363 21511 21369
rect 20346 21332 20352 21344
rect 16960 21304 20352 21332
rect 20346 21292 20352 21304
rect 20404 21292 20410 21344
rect 20438 21292 20444 21344
rect 20496 21332 20502 21344
rect 21468 21332 21496 21363
rect 20496 21304 21496 21332
rect 20496 21292 20502 21304
rect 21726 21292 21732 21344
rect 21784 21292 21790 21344
rect 21836 21332 21864 21431
rect 23842 21428 23848 21440
rect 23900 21428 23906 21480
rect 24394 21477 24400 21480
rect 24364 21471 24400 21477
rect 24364 21437 24376 21471
rect 24364 21431 24400 21437
rect 24394 21428 24400 21431
rect 24452 21428 24458 21480
rect 25314 21428 25320 21480
rect 25372 21428 25378 21480
rect 21910 21360 21916 21412
rect 21968 21400 21974 21412
rect 22066 21403 22124 21409
rect 22066 21400 22078 21403
rect 21968 21372 22078 21400
rect 21968 21360 21974 21372
rect 22066 21369 22078 21372
rect 22112 21369 22124 21403
rect 22066 21363 22124 21369
rect 22922 21360 22928 21412
rect 22980 21360 22986 21412
rect 24581 21403 24639 21409
rect 24581 21369 24593 21403
rect 24627 21369 24639 21403
rect 24581 21363 24639 21369
rect 22278 21332 22284 21344
rect 21836 21304 22284 21332
rect 22278 21292 22284 21304
rect 22336 21292 22342 21344
rect 22940 21332 22968 21360
rect 24305 21335 24363 21341
rect 24305 21332 24317 21335
rect 22940 21304 24317 21332
rect 24305 21301 24317 21304
rect 24351 21332 24363 21335
rect 24596 21332 24624 21363
rect 24351 21304 24624 21332
rect 24351 21301 24363 21304
rect 24305 21295 24363 21301
rect 552 21242 27576 21264
rect 552 21190 7114 21242
rect 7166 21190 7178 21242
rect 7230 21190 7242 21242
rect 7294 21190 7306 21242
rect 7358 21190 7370 21242
rect 7422 21190 13830 21242
rect 13882 21190 13894 21242
rect 13946 21190 13958 21242
rect 14010 21190 14022 21242
rect 14074 21190 14086 21242
rect 14138 21190 20546 21242
rect 20598 21190 20610 21242
rect 20662 21190 20674 21242
rect 20726 21190 20738 21242
rect 20790 21190 20802 21242
rect 20854 21190 27262 21242
rect 27314 21190 27326 21242
rect 27378 21190 27390 21242
rect 27442 21190 27454 21242
rect 27506 21190 27518 21242
rect 27570 21190 27576 21242
rect 552 21168 27576 21190
rect 2682 21088 2688 21140
rect 2740 21088 2746 21140
rect 3418 21088 3424 21140
rect 3476 21128 3482 21140
rect 4985 21131 5043 21137
rect 4985 21128 4997 21131
rect 3476 21100 4997 21128
rect 3476 21088 3482 21100
rect 4985 21097 4997 21100
rect 5031 21097 5043 21131
rect 4985 21091 5043 21097
rect 5074 21088 5080 21140
rect 5132 21128 5138 21140
rect 5445 21131 5503 21137
rect 5445 21128 5457 21131
rect 5132 21100 5457 21128
rect 5132 21088 5138 21100
rect 5445 21097 5457 21100
rect 5491 21097 5503 21131
rect 5445 21091 5503 21097
rect 7006 21088 7012 21140
rect 7064 21128 7070 21140
rect 7101 21131 7159 21137
rect 7101 21128 7113 21131
rect 7064 21100 7113 21128
rect 7064 21088 7070 21100
rect 7101 21097 7113 21100
rect 7147 21097 7159 21131
rect 7101 21091 7159 21097
rect 842 20952 848 21004
rect 900 20992 906 21004
rect 1765 20995 1823 21001
rect 1765 20992 1777 20995
rect 900 20964 1777 20992
rect 900 20952 906 20964
rect 1765 20961 1777 20964
rect 1811 20961 1823 20995
rect 2700 20992 2728 21088
rect 3234 21020 3240 21072
rect 3292 21060 3298 21072
rect 3513 21063 3571 21069
rect 3513 21060 3525 21063
rect 3292 21032 3525 21060
rect 3292 21020 3298 21032
rect 3513 21029 3525 21032
rect 3559 21060 3571 21063
rect 3559 21032 5948 21060
rect 3559 21029 3571 21032
rect 3513 21023 3571 21029
rect 5920 21004 5948 21032
rect 3861 20995 3919 21001
rect 3861 20992 3873 20995
rect 2700 20964 3873 20992
rect 1765 20955 1823 20961
rect 3861 20961 3873 20964
rect 3907 20961 3919 20995
rect 3861 20955 3919 20961
rect 5307 20995 5365 21001
rect 5307 20961 5319 20995
rect 5353 20992 5365 20995
rect 5537 20995 5595 21001
rect 5353 20964 5488 20992
rect 5353 20961 5365 20964
rect 5307 20955 5365 20961
rect 1578 20884 1584 20936
rect 1636 20884 1642 20936
rect 1780 20924 1808 20955
rect 3602 20924 3608 20936
rect 1780 20896 3608 20924
rect 3602 20884 3608 20896
rect 3660 20884 3666 20936
rect 5460 20924 5488 20964
rect 5537 20961 5549 20995
rect 5583 20992 5595 20995
rect 5810 20992 5816 21004
rect 5583 20964 5816 20992
rect 5583 20961 5595 20964
rect 5537 20955 5595 20961
rect 5810 20952 5816 20964
rect 5868 20952 5874 21004
rect 5902 20952 5908 21004
rect 5960 20952 5966 21004
rect 7116 20992 7144 21091
rect 7466 21088 7472 21140
rect 7524 21088 7530 21140
rect 7834 21088 7840 21140
rect 7892 21088 7898 21140
rect 10410 21088 10416 21140
rect 10468 21128 10474 21140
rect 11149 21131 11207 21137
rect 11149 21128 11161 21131
rect 10468 21100 11161 21128
rect 10468 21088 10474 21100
rect 11149 21097 11161 21100
rect 11195 21097 11207 21131
rect 11149 21091 11207 21097
rect 12434 21088 12440 21140
rect 12492 21128 12498 21140
rect 14001 21131 14059 21137
rect 12492 21100 13952 21128
rect 12492 21088 12498 21100
rect 7484 21060 7512 21088
rect 7678 21063 7736 21069
rect 7678 21060 7690 21063
rect 7484 21032 7690 21060
rect 7678 21029 7690 21032
rect 7724 21029 7736 21063
rect 7678 21023 7736 21029
rect 13262 21020 13268 21072
rect 13320 21020 13326 21072
rect 7193 20995 7251 21001
rect 7193 20992 7205 20995
rect 7116 20964 7205 20992
rect 7193 20961 7205 20964
rect 7239 20961 7251 20995
rect 7193 20955 7251 20961
rect 7466 20952 7472 21004
rect 7524 20952 7530 21004
rect 9053 20995 9111 21001
rect 9053 20961 9065 20995
rect 9099 20992 9111 20995
rect 9214 20992 9220 21004
rect 9099 20964 9220 20992
rect 9099 20961 9111 20964
rect 9053 20955 9111 20961
rect 9214 20952 9220 20964
rect 9272 20952 9278 21004
rect 9950 20952 9956 21004
rect 10008 20992 10014 21004
rect 10514 20995 10572 21001
rect 10514 20992 10526 20995
rect 10008 20964 10526 20992
rect 10008 20952 10014 20964
rect 10514 20961 10526 20964
rect 10560 20961 10572 20995
rect 10514 20955 10572 20961
rect 10962 20952 10968 21004
rect 11020 20952 11026 21004
rect 11790 20952 11796 21004
rect 11848 20952 11854 21004
rect 12161 20995 12219 21001
rect 12161 20961 12173 20995
rect 12207 20961 12219 20995
rect 12161 20955 12219 20961
rect 12253 20995 12311 21001
rect 12253 20961 12265 20995
rect 12299 20961 12311 20995
rect 12253 20955 12311 20961
rect 12437 20995 12495 21001
rect 12437 20961 12449 20995
rect 12483 20992 12495 20995
rect 12713 20995 12771 21001
rect 12713 20992 12725 20995
rect 12483 20964 12725 20992
rect 12483 20961 12495 20964
rect 12437 20955 12495 20961
rect 12713 20961 12725 20964
rect 12759 20961 12771 20995
rect 13280 20992 13308 21020
rect 13449 20995 13507 21001
rect 13449 20992 13461 20995
rect 13280 20964 13461 20992
rect 12713 20955 12771 20961
rect 13449 20961 13461 20964
rect 13495 20961 13507 20995
rect 13924 20992 13952 21100
rect 14001 21097 14013 21131
rect 14047 21097 14059 21131
rect 14001 21091 14059 21097
rect 14016 21060 14044 21091
rect 14274 21088 14280 21140
rect 14332 21128 14338 21140
rect 16298 21128 16304 21140
rect 14332 21100 16304 21128
rect 14332 21088 14338 21100
rect 16298 21088 16304 21100
rect 16356 21088 16362 21140
rect 17862 21088 17868 21140
rect 17920 21088 17926 21140
rect 19242 21088 19248 21140
rect 19300 21128 19306 21140
rect 19337 21131 19395 21137
rect 19337 21128 19349 21131
rect 19300 21100 19349 21128
rect 19300 21088 19306 21100
rect 19337 21097 19349 21100
rect 19383 21097 19395 21131
rect 19337 21091 19395 21097
rect 21726 21088 21732 21140
rect 21784 21128 21790 21140
rect 21784 21100 22094 21128
rect 21784 21088 21790 21100
rect 14185 21063 14243 21069
rect 14185 21060 14197 21063
rect 14016 21032 14197 21060
rect 14185 21029 14197 21032
rect 14231 21029 14243 21063
rect 14185 21023 14243 21029
rect 14553 21063 14611 21069
rect 14553 21029 14565 21063
rect 14599 21060 14611 21063
rect 17880 21060 17908 21088
rect 18202 21063 18260 21069
rect 18202 21060 18214 21063
rect 14599 21032 16712 21060
rect 17880 21032 18214 21060
rect 14599 21029 14611 21032
rect 14553 21023 14611 21029
rect 14568 20992 14596 21023
rect 16684 21004 16712 21032
rect 18202 21029 18214 21032
rect 18248 21029 18260 21063
rect 18202 21023 18260 21029
rect 18414 21020 18420 21072
rect 18472 21060 18478 21072
rect 20438 21060 20444 21072
rect 18472 21032 20444 21060
rect 18472 21020 18478 21032
rect 20438 21020 20444 21032
rect 20496 21020 20502 21072
rect 21910 21060 21916 21072
rect 21284 21032 21772 21060
rect 13924 20964 14596 20992
rect 15105 20995 15163 21001
rect 13449 20955 13507 20961
rect 15105 20961 15117 20995
rect 15151 20992 15163 20995
rect 15194 20992 15200 21004
rect 15151 20964 15200 20992
rect 15151 20961 15163 20964
rect 15105 20955 15163 20961
rect 6641 20927 6699 20933
rect 5460 20896 5580 20924
rect 5552 20800 5580 20896
rect 6641 20893 6653 20927
rect 6687 20893 6699 20927
rect 6641 20887 6699 20893
rect 7561 20927 7619 20933
rect 7561 20893 7573 20927
rect 7607 20924 7619 20927
rect 7650 20924 7656 20936
rect 7607 20896 7656 20924
rect 7607 20893 7619 20896
rect 7561 20887 7619 20893
rect 1029 20791 1087 20797
rect 1029 20757 1041 20791
rect 1075 20788 1087 20791
rect 1118 20788 1124 20800
rect 1075 20760 1124 20788
rect 1075 20757 1087 20760
rect 1029 20751 1087 20757
rect 1118 20748 1124 20760
rect 1176 20748 1182 20800
rect 5074 20748 5080 20800
rect 5132 20748 5138 20800
rect 5534 20748 5540 20800
rect 5592 20788 5598 20800
rect 6656 20788 6684 20887
rect 7650 20884 7656 20896
rect 7708 20884 7714 20936
rect 9309 20927 9367 20933
rect 9309 20893 9321 20927
rect 9355 20924 9367 20927
rect 9766 20924 9772 20936
rect 9355 20896 9772 20924
rect 9355 20893 9367 20896
rect 9309 20887 9367 20893
rect 9766 20884 9772 20896
rect 9824 20884 9830 20936
rect 10781 20927 10839 20933
rect 10781 20893 10793 20927
rect 10827 20924 10839 20927
rect 11808 20924 11836 20952
rect 10827 20896 11836 20924
rect 10827 20893 10839 20896
rect 10781 20887 10839 20893
rect 7006 20816 7012 20868
rect 7064 20856 7070 20868
rect 12176 20856 12204 20955
rect 12268 20924 12296 20955
rect 15194 20952 15200 20964
rect 15252 20952 15258 21004
rect 15289 20995 15347 21001
rect 15289 20961 15301 20995
rect 15335 20992 15347 20995
rect 15381 20995 15439 21001
rect 15381 20992 15393 20995
rect 15335 20964 15393 20992
rect 15335 20961 15347 20964
rect 15289 20955 15347 20961
rect 15381 20961 15393 20964
rect 15427 20961 15439 20995
rect 15381 20955 15439 20961
rect 16666 20952 16672 21004
rect 16724 20952 16730 21004
rect 17865 20995 17923 21001
rect 17865 20961 17877 20995
rect 17911 20992 17923 20995
rect 18046 20992 18052 21004
rect 17911 20964 18052 20992
rect 17911 20961 17923 20964
rect 17865 20955 17923 20961
rect 18046 20952 18052 20964
rect 18104 20952 18110 21004
rect 18506 20952 18512 21004
rect 18564 20992 18570 21004
rect 19150 20992 19156 21004
rect 18564 20964 19156 20992
rect 18564 20952 18570 20964
rect 19150 20952 19156 20964
rect 19208 20952 19214 21004
rect 19610 20952 19616 21004
rect 19668 20952 19674 21004
rect 20717 20995 20775 21001
rect 20717 20961 20729 20995
rect 20763 20992 20775 20995
rect 20990 20992 20996 21004
rect 20763 20964 20996 20992
rect 20763 20961 20775 20964
rect 20717 20955 20775 20961
rect 20990 20952 20996 20964
rect 21048 20952 21054 21004
rect 21284 21001 21312 21032
rect 21744 21004 21772 21032
rect 21836 21032 21916 21060
rect 21269 20995 21327 21001
rect 21269 20961 21281 20995
rect 21315 20961 21327 20995
rect 21269 20955 21327 20961
rect 21358 20952 21364 21004
rect 21416 20992 21422 21004
rect 21453 20995 21511 21001
rect 21453 20992 21465 20995
rect 21416 20964 21465 20992
rect 21416 20952 21422 20964
rect 21453 20961 21465 20964
rect 21499 20961 21511 20995
rect 21453 20955 21511 20961
rect 21545 20995 21603 21001
rect 21545 20961 21557 20995
rect 21591 20961 21603 20995
rect 21545 20955 21603 20961
rect 12618 20924 12624 20936
rect 12268 20896 12624 20924
rect 12618 20884 12624 20896
rect 12676 20884 12682 20936
rect 13630 20884 13636 20936
rect 13688 20924 13694 20936
rect 13725 20927 13783 20933
rect 13725 20924 13737 20927
rect 13688 20896 13737 20924
rect 13688 20884 13694 20896
rect 13725 20893 13737 20896
rect 13771 20893 13783 20927
rect 13725 20887 13783 20893
rect 14921 20927 14979 20933
rect 14921 20893 14933 20927
rect 14967 20924 14979 20927
rect 17954 20924 17960 20936
rect 14967 20896 15148 20924
rect 14967 20893 14979 20896
rect 14921 20887 14979 20893
rect 15120 20856 15148 20896
rect 16408 20896 17960 20924
rect 7064 20828 8432 20856
rect 12176 20828 15148 20856
rect 7064 20816 7070 20828
rect 7834 20788 7840 20800
rect 5592 20760 7840 20788
rect 5592 20748 5598 20760
rect 7834 20748 7840 20760
rect 7892 20748 7898 20800
rect 7926 20748 7932 20800
rect 7984 20748 7990 20800
rect 8404 20788 8432 20828
rect 15120 20800 15148 20828
rect 15565 20859 15623 20865
rect 15565 20825 15577 20859
rect 15611 20856 15623 20859
rect 15930 20856 15936 20868
rect 15611 20828 15936 20856
rect 15611 20825 15623 20828
rect 15565 20819 15623 20825
rect 15930 20816 15936 20828
rect 15988 20816 15994 20868
rect 9398 20788 9404 20800
rect 8404 20760 9404 20788
rect 9398 20748 9404 20760
rect 9456 20748 9462 20800
rect 12342 20748 12348 20800
rect 12400 20788 12406 20800
rect 12529 20791 12587 20797
rect 12529 20788 12541 20791
rect 12400 20760 12541 20788
rect 12400 20748 12406 20760
rect 12529 20757 12541 20760
rect 12575 20757 12587 20791
rect 12529 20751 12587 20757
rect 13817 20791 13875 20797
rect 13817 20757 13829 20791
rect 13863 20788 13875 20791
rect 14090 20788 14096 20800
rect 13863 20760 14096 20788
rect 13863 20757 13875 20760
rect 13817 20751 13875 20757
rect 14090 20748 14096 20760
rect 14148 20748 14154 20800
rect 15102 20748 15108 20800
rect 15160 20748 15166 20800
rect 15838 20748 15844 20800
rect 15896 20788 15902 20800
rect 16408 20797 16436 20896
rect 17954 20884 17960 20896
rect 18012 20884 18018 20936
rect 19168 20924 19196 20952
rect 20254 20924 20260 20936
rect 19168 20896 20260 20924
rect 20254 20884 20260 20896
rect 20312 20924 20318 20936
rect 21560 20924 21588 20955
rect 21634 20952 21640 21004
rect 21692 20952 21698 21004
rect 21726 20952 21732 21004
rect 21784 20952 21790 21004
rect 20312 20896 21588 20924
rect 20312 20884 20318 20896
rect 16666 20816 16672 20868
rect 16724 20816 16730 20868
rect 21836 20865 21864 21032
rect 21910 21020 21916 21032
rect 21968 21020 21974 21072
rect 22066 21060 22094 21100
rect 22922 21088 22928 21140
rect 22980 21128 22986 21140
rect 23293 21131 23351 21137
rect 23293 21128 23305 21131
rect 22980 21100 23305 21128
rect 22980 21088 22986 21100
rect 23293 21097 23305 21100
rect 23339 21097 23351 21131
rect 23293 21091 23351 21097
rect 23842 21088 23848 21140
rect 23900 21088 23906 21140
rect 24026 21088 24032 21140
rect 24084 21088 24090 21140
rect 24857 21131 24915 21137
rect 24857 21097 24869 21131
rect 24903 21128 24915 21131
rect 25498 21128 25504 21140
rect 24903 21100 25504 21128
rect 24903 21097 24915 21100
rect 24857 21091 24915 21097
rect 25498 21088 25504 21100
rect 25556 21088 25562 21140
rect 25866 21088 25872 21140
rect 25924 21088 25930 21140
rect 26418 21088 26424 21140
rect 26476 21088 26482 21140
rect 26970 21088 26976 21140
rect 27028 21088 27034 21140
rect 22158 21063 22216 21069
rect 22158 21060 22170 21063
rect 22066 21032 22170 21060
rect 22158 21029 22170 21032
rect 22204 21029 22216 21063
rect 22158 21023 22216 21029
rect 23860 20992 23888 21088
rect 24213 21063 24271 21069
rect 24213 21029 24225 21063
rect 24259 21060 24271 21063
rect 25130 21060 25136 21072
rect 24259 21032 25136 21060
rect 24259 21029 24271 21032
rect 24213 21023 24271 21029
rect 25130 21020 25136 21032
rect 25188 21020 25194 21072
rect 25884 21060 25912 21088
rect 25970 21063 26028 21069
rect 25970 21060 25982 21063
rect 25884 21032 25982 21060
rect 25970 21029 25982 21032
rect 26016 21029 26028 21063
rect 25970 21023 26028 21029
rect 26142 21020 26148 21072
rect 26200 21020 26206 21072
rect 23937 20995 23995 21001
rect 23937 20992 23949 20995
rect 23860 20964 23949 20992
rect 23937 20961 23949 20964
rect 23983 20961 23995 20995
rect 23937 20955 23995 20961
rect 21913 20927 21971 20933
rect 21913 20893 21925 20927
rect 21959 20893 21971 20927
rect 26160 20924 26188 21020
rect 26237 20995 26295 21001
rect 26237 20961 26249 20995
rect 26283 20992 26295 20995
rect 26510 20992 26516 21004
rect 26283 20964 26516 20992
rect 26283 20961 26295 20964
rect 26237 20955 26295 20961
rect 26510 20952 26516 20964
rect 26568 20952 26574 21004
rect 26605 20995 26663 21001
rect 26605 20961 26617 20995
rect 26651 20992 26663 20995
rect 26694 20992 26700 21004
rect 26651 20964 26700 20992
rect 26651 20961 26663 20964
rect 26605 20955 26663 20961
rect 26694 20952 26700 20964
rect 26752 20952 26758 21004
rect 26789 20995 26847 21001
rect 26789 20961 26801 20995
rect 26835 20992 26847 20995
rect 26881 20995 26939 21001
rect 26881 20992 26893 20995
rect 26835 20964 26893 20992
rect 26835 20961 26847 20964
rect 26789 20955 26847 20961
rect 26881 20961 26893 20964
rect 26927 20961 26939 20995
rect 26881 20955 26939 20961
rect 26804 20924 26832 20955
rect 26970 20952 26976 21004
rect 27028 20992 27034 21004
rect 27065 20995 27123 21001
rect 27065 20992 27077 20995
rect 27028 20964 27077 20992
rect 27028 20952 27034 20964
rect 27065 20961 27077 20964
rect 27111 20961 27123 20995
rect 27065 20955 27123 20961
rect 26160 20896 26832 20924
rect 21913 20887 21971 20893
rect 21821 20859 21879 20865
rect 21821 20825 21833 20859
rect 21867 20825 21879 20859
rect 21821 20819 21879 20825
rect 16393 20791 16451 20797
rect 16393 20788 16405 20791
rect 15896 20760 16405 20788
rect 15896 20748 15902 20760
rect 16393 20757 16405 20760
rect 16439 20757 16451 20791
rect 16684 20788 16712 20816
rect 18690 20788 18696 20800
rect 16684 20760 18696 20788
rect 16393 20751 16451 20757
rect 18690 20748 18696 20760
rect 18748 20748 18754 20800
rect 19334 20748 19340 20800
rect 19392 20788 19398 20800
rect 19429 20791 19487 20797
rect 19429 20788 19441 20791
rect 19392 20760 19441 20788
rect 19392 20748 19398 20760
rect 19429 20757 19441 20760
rect 19475 20757 19487 20791
rect 19429 20751 19487 20757
rect 20898 20748 20904 20800
rect 20956 20748 20962 20800
rect 21928 20788 21956 20887
rect 24213 20859 24271 20865
rect 24213 20825 24225 20859
rect 24259 20856 24271 20859
rect 24578 20856 24584 20868
rect 24259 20828 24584 20856
rect 24259 20825 24271 20828
rect 24213 20819 24271 20825
rect 24578 20816 24584 20828
rect 24636 20816 24642 20868
rect 22278 20788 22284 20800
rect 21928 20760 22284 20788
rect 22278 20748 22284 20760
rect 22336 20748 22342 20800
rect 552 20698 27416 20720
rect 552 20646 3756 20698
rect 3808 20646 3820 20698
rect 3872 20646 3884 20698
rect 3936 20646 3948 20698
rect 4000 20646 4012 20698
rect 4064 20646 10472 20698
rect 10524 20646 10536 20698
rect 10588 20646 10600 20698
rect 10652 20646 10664 20698
rect 10716 20646 10728 20698
rect 10780 20646 17188 20698
rect 17240 20646 17252 20698
rect 17304 20646 17316 20698
rect 17368 20646 17380 20698
rect 17432 20646 17444 20698
rect 17496 20646 23904 20698
rect 23956 20646 23968 20698
rect 24020 20646 24032 20698
rect 24084 20646 24096 20698
rect 24148 20646 24160 20698
rect 24212 20646 27416 20698
rect 552 20624 27416 20646
rect 2222 20544 2228 20596
rect 2280 20544 2286 20596
rect 2774 20544 2780 20596
rect 2832 20544 2838 20596
rect 2869 20587 2927 20593
rect 2869 20553 2881 20587
rect 2915 20584 2927 20587
rect 3326 20584 3332 20596
rect 2915 20556 3332 20584
rect 2915 20553 2927 20556
rect 2869 20547 2927 20553
rect 3326 20544 3332 20556
rect 3384 20544 3390 20596
rect 3421 20587 3479 20593
rect 3421 20553 3433 20587
rect 3467 20584 3479 20587
rect 3510 20584 3516 20596
rect 3467 20556 3516 20584
rect 3467 20553 3479 20556
rect 3421 20547 3479 20553
rect 842 20340 848 20392
rect 900 20340 906 20392
rect 1118 20389 1124 20392
rect 1112 20380 1124 20389
rect 1079 20352 1124 20380
rect 1112 20343 1124 20352
rect 1118 20340 1124 20343
rect 1176 20340 1182 20392
rect 2240 20312 2268 20544
rect 2792 20516 2820 20544
rect 3053 20519 3111 20525
rect 3053 20516 3065 20519
rect 2792 20488 3065 20516
rect 3053 20485 3065 20488
rect 3099 20485 3111 20519
rect 3436 20516 3464 20547
rect 3510 20544 3516 20556
rect 3568 20544 3574 20596
rect 3602 20544 3608 20596
rect 3660 20544 3666 20596
rect 4982 20544 4988 20596
rect 5040 20584 5046 20596
rect 6917 20587 6975 20593
rect 6917 20584 6929 20587
rect 5040 20556 6929 20584
rect 5040 20544 5046 20556
rect 6917 20553 6929 20556
rect 6963 20553 6975 20587
rect 6917 20547 6975 20553
rect 7377 20587 7435 20593
rect 7377 20553 7389 20587
rect 7423 20584 7435 20587
rect 7466 20584 7472 20596
rect 7423 20556 7472 20584
rect 7423 20553 7435 20556
rect 7377 20547 7435 20553
rect 3053 20479 3111 20485
rect 3344 20488 3464 20516
rect 3344 20460 3372 20488
rect 3326 20408 3332 20460
rect 3384 20408 3390 20460
rect 3620 20448 3648 20544
rect 5077 20519 5135 20525
rect 5077 20485 5089 20519
rect 5123 20516 5135 20519
rect 5534 20516 5540 20528
rect 5123 20488 5540 20516
rect 5123 20485 5135 20488
rect 5077 20479 5135 20485
rect 5534 20476 5540 20488
rect 5592 20476 5598 20528
rect 3697 20451 3755 20457
rect 3697 20448 3709 20451
rect 3620 20420 3709 20448
rect 3697 20417 3709 20420
rect 3743 20417 3755 20451
rect 3697 20411 3755 20417
rect 5184 20420 5488 20448
rect 2314 20340 2320 20392
rect 2372 20380 2378 20392
rect 2501 20383 2559 20389
rect 2501 20380 2513 20383
rect 2372 20352 2513 20380
rect 2372 20340 2378 20352
rect 2501 20349 2513 20352
rect 2547 20380 2559 20383
rect 2547 20352 3648 20380
rect 2547 20349 2559 20352
rect 2501 20343 2559 20349
rect 3237 20315 3295 20321
rect 3237 20312 3249 20315
rect 2240 20284 3249 20312
rect 3237 20281 3249 20284
rect 3283 20281 3295 20315
rect 3237 20275 3295 20281
rect 3418 20272 3424 20324
rect 3476 20321 3482 20324
rect 3476 20315 3495 20321
rect 3483 20281 3495 20315
rect 3476 20275 3495 20281
rect 3476 20272 3482 20275
rect 2866 20204 2872 20256
rect 2924 20204 2930 20256
rect 3620 20253 3648 20352
rect 4430 20340 4436 20392
rect 4488 20380 4494 20392
rect 5184 20380 5212 20420
rect 5460 20389 5488 20420
rect 4488 20352 5212 20380
rect 5261 20383 5319 20389
rect 4488 20340 4494 20352
rect 5261 20349 5273 20383
rect 5307 20349 5319 20383
rect 5261 20343 5319 20349
rect 5445 20383 5503 20389
rect 5445 20349 5457 20383
rect 5491 20349 5503 20383
rect 5445 20343 5503 20349
rect 5537 20383 5595 20389
rect 5537 20349 5549 20383
rect 5583 20380 5595 20383
rect 6270 20380 6276 20392
rect 5583 20352 6276 20380
rect 5583 20349 5595 20352
rect 5537 20343 5595 20349
rect 3970 20321 3976 20324
rect 3964 20275 3976 20321
rect 3970 20272 3976 20275
rect 4028 20272 4034 20324
rect 5276 20256 5304 20343
rect 6270 20340 6276 20352
rect 6328 20340 6334 20392
rect 6932 20380 6960 20547
rect 7466 20544 7472 20556
rect 7524 20544 7530 20596
rect 7745 20587 7803 20593
rect 7745 20553 7757 20587
rect 7791 20584 7803 20587
rect 7926 20584 7932 20596
rect 7791 20556 7932 20584
rect 7791 20553 7803 20556
rect 7745 20547 7803 20553
rect 7926 20544 7932 20556
rect 7984 20584 7990 20596
rect 7984 20556 8432 20584
rect 7984 20544 7990 20556
rect 8404 20457 8432 20556
rect 8570 20544 8576 20596
rect 8628 20584 8634 20596
rect 14182 20584 14188 20596
rect 8628 20556 14188 20584
rect 8628 20544 8634 20556
rect 14182 20544 14188 20556
rect 14240 20544 14246 20596
rect 14553 20587 14611 20593
rect 14553 20553 14565 20587
rect 14599 20584 14611 20587
rect 14826 20584 14832 20596
rect 14599 20556 14832 20584
rect 14599 20553 14611 20556
rect 14553 20547 14611 20553
rect 14826 20544 14832 20556
rect 14884 20544 14890 20596
rect 14936 20556 17908 20584
rect 14458 20516 14464 20528
rect 13096 20488 14464 20516
rect 8389 20451 8447 20457
rect 8389 20417 8401 20451
rect 8435 20417 8447 20451
rect 8389 20411 8447 20417
rect 9398 20408 9404 20460
rect 9456 20408 9462 20460
rect 9766 20408 9772 20460
rect 9824 20448 9830 20460
rect 10226 20448 10232 20460
rect 9824 20420 10232 20448
rect 9824 20408 9830 20420
rect 10226 20408 10232 20420
rect 10284 20448 10290 20460
rect 10321 20451 10379 20457
rect 10321 20448 10333 20451
rect 10284 20420 10333 20448
rect 10284 20408 10290 20420
rect 10321 20417 10333 20420
rect 10367 20417 10379 20451
rect 10321 20411 10379 20417
rect 11790 20408 11796 20460
rect 11848 20408 11854 20460
rect 7742 20380 7748 20392
rect 6932 20352 7748 20380
rect 7742 20340 7748 20352
rect 7800 20380 7806 20392
rect 7837 20383 7895 20389
rect 7837 20380 7849 20383
rect 7800 20352 7849 20380
rect 7800 20340 7806 20352
rect 7837 20349 7849 20352
rect 7883 20349 7895 20383
rect 7837 20343 7895 20349
rect 12060 20383 12118 20389
rect 12060 20349 12072 20383
rect 12106 20380 12118 20383
rect 12342 20380 12348 20392
rect 12106 20352 12348 20380
rect 12106 20349 12118 20352
rect 12060 20343 12118 20349
rect 12342 20340 12348 20352
rect 12400 20340 12406 20392
rect 5353 20315 5411 20321
rect 5353 20281 5365 20315
rect 5399 20312 5411 20315
rect 5782 20315 5840 20321
rect 5782 20312 5794 20315
rect 5399 20284 5794 20312
rect 5399 20281 5411 20284
rect 5353 20275 5411 20281
rect 5782 20281 5794 20284
rect 5828 20281 5840 20315
rect 5782 20275 5840 20281
rect 9398 20272 9404 20324
rect 9456 20312 9462 20324
rect 10588 20315 10646 20321
rect 9456 20284 10180 20312
rect 9456 20272 9462 20284
rect 3605 20247 3663 20253
rect 3605 20213 3617 20247
rect 3651 20213 3663 20247
rect 3605 20207 3663 20213
rect 5258 20204 5264 20256
rect 5316 20204 5322 20256
rect 9030 20204 9036 20256
rect 9088 20204 9094 20256
rect 10042 20204 10048 20256
rect 10100 20204 10106 20256
rect 10152 20244 10180 20284
rect 10588 20281 10600 20315
rect 10634 20312 10646 20315
rect 11054 20312 11060 20324
rect 10634 20284 11060 20312
rect 10634 20281 10646 20284
rect 10588 20275 10646 20281
rect 11054 20272 11060 20284
rect 11112 20272 11118 20324
rect 11330 20272 11336 20324
rect 11388 20312 11394 20324
rect 13096 20312 13124 20488
rect 14458 20476 14464 20488
rect 14516 20516 14522 20528
rect 14936 20516 14964 20556
rect 14516 20488 14964 20516
rect 14516 20476 14522 20488
rect 13262 20408 13268 20460
rect 13320 20448 13326 20460
rect 14182 20448 14188 20460
rect 13320 20420 14188 20448
rect 13320 20408 13326 20420
rect 13630 20380 13636 20392
rect 11388 20284 13124 20312
rect 13188 20352 13636 20380
rect 11388 20272 11394 20284
rect 11146 20244 11152 20256
rect 10152 20216 11152 20244
rect 11146 20204 11152 20216
rect 11204 20204 11210 20256
rect 11701 20247 11759 20253
rect 11701 20213 11713 20247
rect 11747 20244 11759 20247
rect 12526 20244 12532 20256
rect 11747 20216 12532 20244
rect 11747 20213 11759 20216
rect 11701 20207 11759 20213
rect 12526 20204 12532 20216
rect 12584 20204 12590 20256
rect 13078 20204 13084 20256
rect 13136 20244 13142 20256
rect 13188 20253 13216 20352
rect 13630 20340 13636 20352
rect 13688 20340 13694 20392
rect 13740 20389 13768 20420
rect 14182 20408 14188 20420
rect 14240 20408 14246 20460
rect 14277 20451 14335 20457
rect 14277 20417 14289 20451
rect 14323 20448 14335 20451
rect 14366 20448 14372 20460
rect 14323 20420 14372 20448
rect 14323 20417 14335 20420
rect 14277 20411 14335 20417
rect 14366 20408 14372 20420
rect 14424 20408 14430 20460
rect 14476 20420 14872 20448
rect 13725 20383 13783 20389
rect 13725 20349 13737 20383
rect 13771 20349 13783 20383
rect 13725 20343 13783 20349
rect 14090 20340 14096 20392
rect 14148 20380 14154 20392
rect 14476 20380 14504 20420
rect 14148 20352 14504 20380
rect 14148 20340 14154 20352
rect 14599 20349 14657 20355
rect 14599 20346 14611 20349
rect 13173 20247 13231 20253
rect 13173 20244 13185 20247
rect 13136 20216 13185 20244
rect 13136 20204 13142 20216
rect 13173 20213 13185 20216
rect 13219 20213 13231 20247
rect 13648 20244 13676 20340
rect 14369 20315 14427 20321
rect 14369 20312 14381 20315
rect 14292 20284 14381 20312
rect 14292 20244 14320 20284
rect 14369 20281 14381 20284
rect 14415 20281 14427 20315
rect 14584 20315 14611 20346
rect 14645 20315 14657 20349
rect 14584 20312 14657 20315
rect 14584 20284 14688 20312
rect 14369 20275 14427 20281
rect 14660 20256 14688 20284
rect 14844 20256 14872 20420
rect 16850 20408 16856 20460
rect 16908 20408 16914 20460
rect 17880 20448 17908 20556
rect 18138 20544 18144 20596
rect 18196 20544 18202 20596
rect 19978 20584 19984 20596
rect 18248 20556 19984 20584
rect 18248 20448 18276 20556
rect 19978 20544 19984 20556
rect 20036 20544 20042 20596
rect 20806 20516 20812 20528
rect 17880 20420 18276 20448
rect 19904 20488 20812 20516
rect 16209 20383 16267 20389
rect 16209 20380 16221 20383
rect 15856 20352 16221 20380
rect 15856 20324 15884 20352
rect 16209 20349 16221 20352
rect 16255 20349 16267 20383
rect 16209 20343 16267 20349
rect 17497 20383 17555 20389
rect 17497 20349 17509 20383
rect 17543 20380 17555 20383
rect 17589 20383 17647 20389
rect 17589 20380 17601 20383
rect 17543 20352 17601 20380
rect 17543 20349 17555 20352
rect 17497 20343 17555 20349
rect 17589 20349 17601 20352
rect 17635 20349 17647 20383
rect 17589 20343 17647 20349
rect 17678 20340 17684 20392
rect 17736 20380 17742 20392
rect 17880 20389 17908 20420
rect 17773 20383 17831 20389
rect 17773 20380 17785 20383
rect 17736 20352 17785 20380
rect 17736 20340 17742 20352
rect 17773 20349 17785 20352
rect 17819 20349 17831 20383
rect 17773 20343 17831 20349
rect 17865 20383 17923 20389
rect 17865 20349 17877 20383
rect 17911 20349 17923 20383
rect 17865 20343 17923 20349
rect 17954 20340 17960 20392
rect 18012 20340 18018 20392
rect 18506 20340 18512 20392
rect 18564 20340 18570 20392
rect 18877 20383 18935 20389
rect 18877 20349 18889 20383
rect 18923 20380 18935 20383
rect 18966 20380 18972 20392
rect 18923 20352 18972 20380
rect 18923 20349 18935 20352
rect 18877 20343 18935 20349
rect 18966 20340 18972 20352
rect 19024 20340 19030 20392
rect 19904 20380 19932 20488
rect 20806 20476 20812 20488
rect 20864 20476 20870 20528
rect 20548 20420 20852 20448
rect 20548 20389 20576 20420
rect 20824 20392 20852 20420
rect 19076 20352 19932 20380
rect 20533 20383 20591 20389
rect 15838 20272 15844 20324
rect 15896 20272 15902 20324
rect 15930 20272 15936 20324
rect 15988 20321 15994 20324
rect 15988 20312 16000 20321
rect 18524 20312 18552 20340
rect 19076 20312 19104 20352
rect 20533 20349 20545 20383
rect 20579 20349 20591 20383
rect 20533 20343 20591 20349
rect 20717 20383 20775 20389
rect 20717 20349 20729 20383
rect 20763 20349 20775 20383
rect 20717 20343 20775 20349
rect 15988 20284 16033 20312
rect 18524 20284 19104 20312
rect 19144 20315 19202 20321
rect 15988 20275 16000 20284
rect 19144 20281 19156 20315
rect 19190 20312 19202 20315
rect 19334 20312 19340 20324
rect 19190 20284 19340 20312
rect 19190 20281 19202 20284
rect 19144 20275 19202 20281
rect 15988 20272 15994 20275
rect 19334 20272 19340 20284
rect 19392 20272 19398 20324
rect 20349 20315 20407 20321
rect 20349 20312 20361 20315
rect 19628 20284 20361 20312
rect 13648 20216 14320 20244
rect 13173 20207 13231 20213
rect 14642 20204 14648 20256
rect 14700 20204 14706 20256
rect 14734 20204 14740 20256
rect 14792 20204 14798 20256
rect 14826 20204 14832 20256
rect 14884 20244 14890 20256
rect 15286 20244 15292 20256
rect 14884 20216 15292 20244
rect 14884 20204 14890 20216
rect 15286 20204 15292 20216
rect 15344 20204 15350 20256
rect 19518 20204 19524 20256
rect 19576 20244 19582 20256
rect 19628 20244 19656 20284
rect 20349 20281 20361 20284
rect 20395 20281 20407 20315
rect 20349 20275 20407 20281
rect 20732 20312 20760 20343
rect 20806 20340 20812 20392
rect 20864 20340 20870 20392
rect 20898 20340 20904 20392
rect 20956 20380 20962 20392
rect 22014 20383 22072 20389
rect 22014 20380 22026 20383
rect 20956 20352 22026 20380
rect 20956 20340 20962 20352
rect 22014 20349 22026 20352
rect 22060 20349 22072 20383
rect 22014 20343 22072 20349
rect 22278 20340 22284 20392
rect 22336 20380 22342 20392
rect 23014 20380 23020 20392
rect 22336 20352 23020 20380
rect 22336 20340 22342 20352
rect 23014 20340 23020 20352
rect 23072 20340 23078 20392
rect 23658 20340 23664 20392
rect 23716 20340 23722 20392
rect 25685 20383 25743 20389
rect 25685 20349 25697 20383
rect 25731 20380 25743 20383
rect 26234 20380 26240 20392
rect 25731 20352 26240 20380
rect 25731 20349 25743 20352
rect 25685 20343 25743 20349
rect 26234 20340 26240 20352
rect 26292 20380 26298 20392
rect 26510 20380 26516 20392
rect 26292 20352 26516 20380
rect 26292 20340 26298 20352
rect 26510 20340 26516 20352
rect 26568 20340 26574 20392
rect 20732 20284 22232 20312
rect 19576 20216 19656 20244
rect 20257 20247 20315 20253
rect 19576 20204 19582 20216
rect 20257 20213 20269 20247
rect 20303 20244 20315 20247
rect 20732 20244 20760 20284
rect 22204 20256 22232 20284
rect 25590 20272 25596 20324
rect 25648 20312 25654 20324
rect 25930 20315 25988 20321
rect 25930 20312 25942 20315
rect 25648 20284 25942 20312
rect 25648 20272 25654 20284
rect 25930 20281 25942 20284
rect 25976 20281 25988 20315
rect 25930 20275 25988 20281
rect 20303 20216 20760 20244
rect 20901 20247 20959 20253
rect 20303 20213 20315 20216
rect 20257 20207 20315 20213
rect 20901 20213 20913 20247
rect 20947 20244 20959 20247
rect 22094 20244 22100 20256
rect 20947 20216 22100 20244
rect 20947 20213 20959 20216
rect 20901 20207 20959 20213
rect 22094 20204 22100 20216
rect 22152 20204 22158 20256
rect 22186 20204 22192 20256
rect 22244 20204 22250 20256
rect 23474 20204 23480 20256
rect 23532 20204 23538 20256
rect 27062 20204 27068 20256
rect 27120 20204 27126 20256
rect 552 20154 27576 20176
rect 552 20102 7114 20154
rect 7166 20102 7178 20154
rect 7230 20102 7242 20154
rect 7294 20102 7306 20154
rect 7358 20102 7370 20154
rect 7422 20102 13830 20154
rect 13882 20102 13894 20154
rect 13946 20102 13958 20154
rect 14010 20102 14022 20154
rect 14074 20102 14086 20154
rect 14138 20102 20546 20154
rect 20598 20102 20610 20154
rect 20662 20102 20674 20154
rect 20726 20102 20738 20154
rect 20790 20102 20802 20154
rect 20854 20102 27262 20154
rect 27314 20102 27326 20154
rect 27378 20102 27390 20154
rect 27442 20102 27454 20154
rect 27506 20102 27518 20154
rect 27570 20102 27576 20154
rect 552 20080 27576 20102
rect 3881 20043 3939 20049
rect 3881 20009 3893 20043
rect 3927 20040 3939 20043
rect 3970 20040 3976 20052
rect 3927 20012 3976 20040
rect 3927 20009 3939 20012
rect 3881 20003 3939 20009
rect 3970 20000 3976 20012
rect 4028 20000 4034 20052
rect 4325 20043 4383 20049
rect 4325 20009 4337 20043
rect 4371 20040 4383 20043
rect 5074 20040 5080 20052
rect 4371 20012 5080 20040
rect 4371 20009 4383 20012
rect 4325 20003 4383 20009
rect 5074 20000 5080 20012
rect 5132 20000 5138 20052
rect 5258 20000 5264 20052
rect 5316 20040 5322 20052
rect 5353 20043 5411 20049
rect 5353 20040 5365 20043
rect 5316 20012 5365 20040
rect 5316 20000 5322 20012
rect 5353 20009 5365 20012
rect 5399 20009 5411 20043
rect 5353 20003 5411 20009
rect 7650 20000 7656 20052
rect 7708 20000 7714 20052
rect 8478 20000 8484 20052
rect 8536 20040 8542 20052
rect 8938 20040 8944 20052
rect 8536 20012 8944 20040
rect 8536 20000 8542 20012
rect 8938 20000 8944 20012
rect 8996 20000 9002 20052
rect 9030 20000 9036 20052
rect 9088 20000 9094 20052
rect 9214 20000 9220 20052
rect 9272 20000 9278 20052
rect 9309 20043 9367 20049
rect 9309 20009 9321 20043
rect 9355 20040 9367 20043
rect 9950 20040 9956 20052
rect 9355 20012 9956 20040
rect 9355 20009 9367 20012
rect 9309 20003 9367 20009
rect 9950 20000 9956 20012
rect 10008 20000 10014 20052
rect 10413 20043 10471 20049
rect 10413 20009 10425 20043
rect 10459 20040 10471 20043
rect 10962 20040 10968 20052
rect 10459 20012 10968 20040
rect 10459 20009 10471 20012
rect 10413 20003 10471 20009
rect 10962 20000 10968 20012
rect 11020 20000 11026 20052
rect 11054 20000 11060 20052
rect 11112 20000 11118 20052
rect 12618 20000 12624 20052
rect 12676 20000 12682 20052
rect 12986 20000 12992 20052
rect 13044 20000 13050 20052
rect 13078 20000 13084 20052
rect 13136 20000 13142 20052
rect 14182 20000 14188 20052
rect 14240 20040 14246 20052
rect 14642 20040 14648 20052
rect 14240 20012 14648 20040
rect 14240 20000 14246 20012
rect 14642 20000 14648 20012
rect 14700 20000 14706 20052
rect 15194 20000 15200 20052
rect 15252 20000 15258 20052
rect 15562 20000 15568 20052
rect 15620 20040 15626 20052
rect 17129 20043 17187 20049
rect 15620 20012 17080 20040
rect 15620 20000 15626 20012
rect 2866 19932 2872 19984
rect 2924 19972 2930 19984
rect 2924 19944 4292 19972
rect 2924 19932 2930 19944
rect 1394 19864 1400 19916
rect 1452 19864 1458 19916
rect 4065 19907 4123 19913
rect 4065 19873 4077 19907
rect 4111 19904 4123 19907
rect 4264 19904 4292 19944
rect 4430 19932 4436 19984
rect 4488 19972 4494 19984
rect 4525 19975 4583 19981
rect 4525 19972 4537 19975
rect 4488 19944 4537 19972
rect 4488 19932 4494 19944
rect 4525 19941 4537 19944
rect 4571 19941 4583 19975
rect 6546 19972 6552 19984
rect 4525 19935 4583 19941
rect 4908 19944 6552 19972
rect 4908 19904 4936 19944
rect 6546 19932 6552 19944
rect 6604 19932 6610 19984
rect 9048 19972 9076 20000
rect 8680 19944 9076 19972
rect 9585 19975 9643 19981
rect 4111 19876 4200 19904
rect 4264 19876 4936 19904
rect 4111 19873 4123 19876
rect 4065 19867 4123 19873
rect 4172 19777 4200 19876
rect 4982 19864 4988 19916
rect 5040 19864 5046 19916
rect 6089 19907 6147 19913
rect 6089 19873 6101 19907
rect 6135 19904 6147 19907
rect 6917 19907 6975 19913
rect 6917 19904 6929 19907
rect 6135 19876 6929 19904
rect 6135 19873 6147 19876
rect 6089 19867 6147 19873
rect 6917 19873 6929 19876
rect 6963 19873 6975 19907
rect 6917 19867 6975 19873
rect 7834 19864 7840 19916
rect 7892 19904 7898 19916
rect 8680 19913 8708 19944
rect 9585 19941 9597 19975
rect 9631 19972 9643 19975
rect 11330 19972 11336 19984
rect 9631 19944 11336 19972
rect 9631 19941 9643 19944
rect 9585 19935 9643 19941
rect 11330 19932 11336 19944
rect 11388 19932 11394 19984
rect 13004 19972 13032 20000
rect 12912 19944 13032 19972
rect 8113 19907 8171 19913
rect 8113 19904 8125 19907
rect 7892 19876 8125 19904
rect 7892 19864 7898 19876
rect 8113 19873 8125 19876
rect 8159 19873 8171 19907
rect 8113 19867 8171 19873
rect 8665 19907 8723 19913
rect 8665 19873 8677 19907
rect 8711 19873 8723 19907
rect 8849 19907 8907 19913
rect 8849 19904 8861 19907
rect 8665 19867 8723 19873
rect 8772 19876 8861 19904
rect 5077 19839 5135 19845
rect 5077 19805 5089 19839
rect 5123 19836 5135 19839
rect 5442 19836 5448 19848
rect 5123 19808 5448 19836
rect 5123 19805 5135 19808
rect 5077 19799 5135 19805
rect 5442 19796 5448 19808
rect 5500 19836 5506 19848
rect 6181 19839 6239 19845
rect 6181 19836 6193 19839
rect 5500 19808 6193 19836
rect 5500 19796 5506 19808
rect 6181 19805 6193 19808
rect 6227 19805 6239 19839
rect 6181 19799 6239 19805
rect 4157 19771 4215 19777
rect 4157 19737 4169 19771
rect 4203 19737 4215 19771
rect 6196 19768 6224 19799
rect 7558 19796 7564 19848
rect 7616 19796 7622 19848
rect 8570 19796 8576 19848
rect 8628 19796 8634 19848
rect 8588 19768 8616 19796
rect 6196 19740 8616 19768
rect 4157 19731 4215 19737
rect 1118 19660 1124 19712
rect 1176 19700 1182 19712
rect 1213 19703 1271 19709
rect 1213 19700 1225 19703
rect 1176 19672 1225 19700
rect 1176 19660 1182 19672
rect 1213 19669 1225 19672
rect 1259 19669 1271 19703
rect 1213 19663 1271 19669
rect 4341 19703 4399 19709
rect 4341 19669 4353 19703
rect 4387 19700 4399 19703
rect 4890 19700 4896 19712
rect 4387 19672 4896 19700
rect 4387 19669 4399 19672
rect 4341 19663 4399 19669
rect 4890 19660 4896 19672
rect 4948 19660 4954 19712
rect 6362 19660 6368 19712
rect 6420 19660 6426 19712
rect 7006 19660 7012 19712
rect 7064 19700 7070 19712
rect 7837 19703 7895 19709
rect 7837 19700 7849 19703
rect 7064 19672 7849 19700
rect 7064 19660 7070 19672
rect 7837 19669 7849 19672
rect 7883 19669 7895 19703
rect 8772 19700 8800 19876
rect 8849 19873 8861 19876
rect 8895 19873 8907 19907
rect 8849 19867 8907 19873
rect 8938 19864 8944 19916
rect 8996 19864 9002 19916
rect 9033 19907 9091 19913
rect 9033 19873 9045 19907
rect 9079 19904 9091 19907
rect 9493 19907 9551 19913
rect 9493 19904 9505 19907
rect 9079 19876 9505 19904
rect 9079 19873 9091 19876
rect 9033 19867 9091 19873
rect 9493 19873 9505 19876
rect 9539 19873 9551 19907
rect 9493 19867 9551 19873
rect 9048 19836 9076 19867
rect 8864 19808 9076 19836
rect 9508 19836 9536 19867
rect 9674 19864 9680 19916
rect 9732 19864 9738 19916
rect 9861 19907 9919 19913
rect 9861 19873 9873 19907
rect 9907 19904 9919 19907
rect 10042 19904 10048 19916
rect 9907 19876 10048 19904
rect 9907 19873 9919 19876
rect 9861 19867 9919 19873
rect 10042 19864 10048 19876
rect 10100 19864 10106 19916
rect 10781 19907 10839 19913
rect 10781 19873 10793 19907
rect 10827 19873 10839 19907
rect 10781 19867 10839 19873
rect 9953 19839 10011 19845
rect 9953 19836 9965 19839
rect 9508 19808 9965 19836
rect 8864 19780 8892 19808
rect 9953 19805 9965 19808
rect 9999 19836 10011 19839
rect 9999 19808 10640 19836
rect 9999 19805 10011 19808
rect 9953 19799 10011 19805
rect 8846 19728 8852 19780
rect 8904 19728 8910 19780
rect 9582 19728 9588 19780
rect 9640 19728 9646 19780
rect 10612 19777 10640 19808
rect 10321 19771 10379 19777
rect 10321 19737 10333 19771
rect 10367 19737 10379 19771
rect 10321 19731 10379 19737
rect 10597 19771 10655 19777
rect 10597 19737 10609 19771
rect 10643 19737 10655 19771
rect 10796 19768 10824 19867
rect 11238 19864 11244 19916
rect 11296 19864 11302 19916
rect 11422 19864 11428 19916
rect 11480 19864 11486 19916
rect 11609 19907 11667 19913
rect 11609 19873 11621 19907
rect 11655 19904 11667 19907
rect 11701 19907 11759 19913
rect 11701 19904 11713 19907
rect 11655 19876 11713 19904
rect 11655 19873 11667 19876
rect 11609 19867 11667 19873
rect 11701 19873 11713 19876
rect 11747 19873 11759 19907
rect 11701 19867 11759 19873
rect 12345 19907 12403 19913
rect 12345 19873 12357 19907
rect 12391 19904 12403 19907
rect 12526 19904 12532 19916
rect 12391 19876 12532 19904
rect 12391 19873 12403 19876
rect 12345 19867 12403 19873
rect 12526 19864 12532 19876
rect 12584 19864 12590 19916
rect 12912 19836 12940 19944
rect 15286 19932 15292 19984
rect 15344 19972 15350 19984
rect 15657 19975 15715 19981
rect 15657 19972 15669 19975
rect 15344 19944 15669 19972
rect 15344 19932 15350 19944
rect 15657 19941 15669 19944
rect 15703 19941 15715 19975
rect 15657 19935 15715 19941
rect 12986 19864 12992 19916
rect 13044 19864 13050 19916
rect 13630 19864 13636 19916
rect 13688 19904 13694 19916
rect 13725 19907 13783 19913
rect 13725 19904 13737 19907
rect 13688 19876 13737 19904
rect 13688 19864 13694 19876
rect 13725 19873 13737 19876
rect 13771 19873 13783 19907
rect 13725 19867 13783 19873
rect 14182 19864 14188 19916
rect 14240 19864 14246 19916
rect 14864 19907 14922 19913
rect 14864 19873 14876 19907
rect 14910 19904 14922 19907
rect 15304 19904 15332 19932
rect 14910 19876 15332 19904
rect 14910 19873 14922 19876
rect 14864 19867 14922 19873
rect 16022 19864 16028 19916
rect 16080 19904 16086 19916
rect 16301 19907 16359 19913
rect 16301 19904 16313 19907
rect 16080 19876 16313 19904
rect 16080 19864 16086 19876
rect 16301 19873 16313 19876
rect 16347 19873 16359 19907
rect 16301 19867 16359 19873
rect 16942 19864 16948 19916
rect 17000 19864 17006 19916
rect 17052 19904 17080 20012
rect 17129 20009 17141 20043
rect 17175 20009 17187 20043
rect 17129 20003 17187 20009
rect 17144 19972 17172 20003
rect 18966 20000 18972 20052
rect 19024 20040 19030 20052
rect 19334 20040 19340 20052
rect 19024 20012 19340 20040
rect 19024 20000 19030 20012
rect 19334 20000 19340 20012
rect 19392 20000 19398 20052
rect 19429 20043 19487 20049
rect 19429 20009 19441 20043
rect 19475 20040 19487 20043
rect 19518 20040 19524 20052
rect 19475 20012 19524 20040
rect 19475 20009 19487 20012
rect 19429 20003 19487 20009
rect 19518 20000 19524 20012
rect 19576 20000 19582 20052
rect 19610 20000 19616 20052
rect 19668 20040 19674 20052
rect 19797 20043 19855 20049
rect 19797 20040 19809 20043
rect 19668 20012 19809 20040
rect 19668 20000 19674 20012
rect 19797 20009 19809 20012
rect 19843 20009 19855 20043
rect 19797 20003 19855 20009
rect 20990 20000 20996 20052
rect 21048 20040 21054 20052
rect 21269 20043 21327 20049
rect 21269 20040 21281 20043
rect 21048 20012 21281 20040
rect 21048 20000 21054 20012
rect 21269 20009 21281 20012
rect 21315 20009 21327 20043
rect 21269 20003 21327 20009
rect 17466 19975 17524 19981
rect 17466 19972 17478 19975
rect 17144 19944 17478 19972
rect 17466 19941 17478 19944
rect 17512 19941 17524 19975
rect 17466 19935 17524 19941
rect 18046 19932 18052 19984
rect 18104 19972 18110 19984
rect 22925 19975 22983 19981
rect 22925 19972 22937 19975
rect 18104 19944 22937 19972
rect 18104 19932 18110 19944
rect 22925 19941 22937 19944
rect 22971 19972 22983 19975
rect 25314 19972 25320 19984
rect 22971 19944 25320 19972
rect 22971 19941 22983 19944
rect 22925 19935 22983 19941
rect 25314 19932 25320 19944
rect 25372 19932 25378 19984
rect 19337 19907 19395 19913
rect 17052 19876 18276 19904
rect 13173 19839 13231 19845
rect 13173 19836 13185 19839
rect 12912 19808 13185 19836
rect 13173 19805 13185 19808
rect 13219 19836 13231 19839
rect 14642 19836 14648 19848
rect 13219 19808 14648 19836
rect 13219 19805 13231 19808
rect 13173 19799 13231 19805
rect 14642 19796 14648 19808
rect 14700 19836 14706 19848
rect 15749 19839 15807 19845
rect 15749 19836 15761 19839
rect 14700 19808 15761 19836
rect 14700 19796 14706 19808
rect 15749 19805 15761 19808
rect 15795 19805 15807 19839
rect 15749 19799 15807 19805
rect 17221 19839 17279 19845
rect 17221 19805 17233 19839
rect 17267 19805 17279 19839
rect 17221 19799 17279 19805
rect 14090 19768 14096 19780
rect 10796 19740 14096 19768
rect 10597 19731 10655 19737
rect 9600 19700 9628 19728
rect 8772 19672 9628 19700
rect 10336 19700 10364 19731
rect 14090 19728 14096 19740
rect 14148 19728 14154 19780
rect 10962 19700 10968 19712
rect 10336 19672 10968 19700
rect 7837 19663 7895 19669
rect 10962 19660 10968 19672
rect 11020 19660 11026 19712
rect 11146 19660 11152 19712
rect 11204 19700 11210 19712
rect 14550 19700 14556 19712
rect 11204 19672 14556 19700
rect 11204 19660 11210 19672
rect 14550 19660 14556 19672
rect 14608 19660 14614 19712
rect 14645 19703 14703 19709
rect 14645 19669 14657 19703
rect 14691 19700 14703 19703
rect 15010 19700 15016 19712
rect 14691 19672 15016 19700
rect 14691 19669 14703 19672
rect 14645 19663 14703 19669
rect 15010 19660 15016 19672
rect 15068 19660 15074 19712
rect 16114 19660 16120 19712
rect 16172 19660 16178 19712
rect 17236 19700 17264 19799
rect 18248 19768 18276 19876
rect 19337 19873 19349 19907
rect 19383 19904 19395 19907
rect 19794 19904 19800 19916
rect 19383 19876 19800 19904
rect 19383 19873 19395 19876
rect 19337 19867 19395 19873
rect 19794 19864 19800 19876
rect 19852 19864 19858 19916
rect 20070 19864 20076 19916
rect 20128 19864 20134 19916
rect 20162 19864 20168 19916
rect 20220 19904 20226 19916
rect 20533 19907 20591 19913
rect 20533 19904 20545 19907
rect 20220 19876 20545 19904
rect 20220 19864 20226 19876
rect 20533 19873 20545 19876
rect 20579 19873 20591 19907
rect 20533 19867 20591 19873
rect 20809 19907 20867 19913
rect 20809 19873 20821 19907
rect 20855 19873 20867 19907
rect 20809 19867 20867 19873
rect 19245 19839 19303 19845
rect 19245 19805 19257 19839
rect 19291 19836 19303 19839
rect 19610 19836 19616 19848
rect 19291 19808 19616 19836
rect 19291 19805 19303 19808
rect 19245 19799 19303 19805
rect 19610 19796 19616 19808
rect 19668 19796 19674 19848
rect 20254 19796 20260 19848
rect 20312 19796 20318 19848
rect 20824 19768 20852 19867
rect 20898 19864 20904 19916
rect 20956 19864 20962 19916
rect 21085 19907 21143 19913
rect 21085 19873 21097 19907
rect 21131 19904 21143 19907
rect 21637 19907 21695 19913
rect 21637 19904 21649 19907
rect 21131 19876 21649 19904
rect 21131 19873 21143 19876
rect 21085 19867 21143 19873
rect 21637 19873 21649 19876
rect 21683 19873 21695 19907
rect 21637 19867 21695 19873
rect 22186 19864 22192 19916
rect 22244 19864 22250 19916
rect 27062 19864 27068 19916
rect 27120 19864 27126 19916
rect 21174 19796 21180 19848
rect 21232 19836 21238 19848
rect 21729 19839 21787 19845
rect 21729 19836 21741 19839
rect 21232 19808 21741 19836
rect 21232 19796 21238 19808
rect 21729 19805 21741 19808
rect 21775 19805 21787 19839
rect 21729 19799 21787 19805
rect 21818 19796 21824 19848
rect 21876 19796 21882 19848
rect 22094 19768 22100 19780
rect 18248 19740 20484 19768
rect 20824 19740 22100 19768
rect 17954 19700 17960 19712
rect 17236 19672 17960 19700
rect 17954 19660 17960 19672
rect 18012 19660 18018 19712
rect 18598 19660 18604 19712
rect 18656 19660 18662 19712
rect 19886 19660 19892 19712
rect 19944 19660 19950 19712
rect 20346 19660 20352 19712
rect 20404 19660 20410 19712
rect 20456 19700 20484 19740
rect 22094 19728 22100 19740
rect 22152 19768 22158 19780
rect 22370 19768 22376 19780
rect 22152 19740 22376 19768
rect 22152 19728 22158 19740
rect 22370 19728 22376 19740
rect 22428 19728 22434 19780
rect 21082 19700 21088 19712
rect 20456 19672 21088 19700
rect 21082 19660 21088 19672
rect 21140 19660 21146 19712
rect 22281 19703 22339 19709
rect 22281 19669 22293 19703
rect 22327 19700 22339 19703
rect 22646 19700 22652 19712
rect 22327 19672 22652 19700
rect 22327 19669 22339 19672
rect 22281 19663 22339 19669
rect 22646 19660 22652 19672
rect 22704 19660 22710 19712
rect 23014 19660 23020 19712
rect 23072 19700 23078 19712
rect 24397 19703 24455 19709
rect 24397 19700 24409 19703
rect 23072 19672 24409 19700
rect 23072 19660 23078 19672
rect 24397 19669 24409 19672
rect 24443 19700 24455 19703
rect 25498 19700 25504 19712
rect 24443 19672 25504 19700
rect 24443 19669 24455 19672
rect 24397 19663 24455 19669
rect 25498 19660 25504 19672
rect 25556 19660 25562 19712
rect 26418 19660 26424 19712
rect 26476 19660 26482 19712
rect 552 19610 27416 19632
rect 552 19558 3756 19610
rect 3808 19558 3820 19610
rect 3872 19558 3884 19610
rect 3936 19558 3948 19610
rect 4000 19558 4012 19610
rect 4064 19558 10472 19610
rect 10524 19558 10536 19610
rect 10588 19558 10600 19610
rect 10652 19558 10664 19610
rect 10716 19558 10728 19610
rect 10780 19558 17188 19610
rect 17240 19558 17252 19610
rect 17304 19558 17316 19610
rect 17368 19558 17380 19610
rect 17432 19558 17444 19610
rect 17496 19558 23904 19610
rect 23956 19558 23968 19610
rect 24020 19558 24032 19610
rect 24084 19558 24096 19610
rect 24148 19558 24160 19610
rect 24212 19558 27416 19610
rect 552 19536 27416 19558
rect 4430 19456 4436 19508
rect 4488 19456 4494 19508
rect 9214 19456 9220 19508
rect 9272 19456 9278 19508
rect 11054 19496 11060 19508
rect 9324 19468 11060 19496
rect 4448 19360 4476 19456
rect 8938 19388 8944 19440
rect 8996 19428 9002 19440
rect 9324 19428 9352 19468
rect 11054 19456 11060 19468
rect 11112 19456 11118 19508
rect 11422 19496 11428 19508
rect 11173 19468 11428 19496
rect 11173 19428 11201 19468
rect 11422 19456 11428 19468
rect 11480 19496 11486 19508
rect 12066 19496 12072 19508
rect 11480 19468 12072 19496
rect 11480 19456 11486 19468
rect 12066 19456 12072 19468
rect 12124 19496 12130 19508
rect 12529 19499 12587 19505
rect 12529 19496 12541 19499
rect 12124 19468 12541 19496
rect 12124 19456 12130 19468
rect 12529 19465 12541 19468
rect 12575 19496 12587 19499
rect 13446 19496 13452 19508
rect 12575 19468 13452 19496
rect 12575 19465 12587 19468
rect 12529 19459 12587 19465
rect 13446 19456 13452 19468
rect 13504 19456 13510 19508
rect 14090 19456 14096 19508
rect 14148 19456 14154 19508
rect 14277 19499 14335 19505
rect 14277 19465 14289 19499
rect 14323 19496 14335 19499
rect 14734 19496 14740 19508
rect 14323 19468 14740 19496
rect 14323 19465 14335 19468
rect 14277 19459 14335 19465
rect 14734 19456 14740 19468
rect 14792 19496 14798 19508
rect 15286 19496 15292 19508
rect 14792 19468 15292 19496
rect 14792 19456 14798 19468
rect 15286 19456 15292 19468
rect 15344 19456 15350 19508
rect 15749 19499 15807 19505
rect 15749 19465 15761 19499
rect 15795 19496 15807 19499
rect 16022 19496 16028 19508
rect 15795 19468 16028 19496
rect 15795 19465 15807 19468
rect 15749 19459 15807 19465
rect 16022 19456 16028 19468
rect 16080 19456 16086 19508
rect 16942 19456 16948 19508
rect 17000 19496 17006 19508
rect 17313 19499 17371 19505
rect 17313 19496 17325 19499
rect 17000 19468 17325 19496
rect 17000 19456 17006 19468
rect 17313 19465 17325 19468
rect 17359 19465 17371 19499
rect 17313 19459 17371 19465
rect 19334 19456 19340 19508
rect 19392 19496 19398 19508
rect 20073 19499 20131 19505
rect 20073 19496 20085 19499
rect 19392 19468 20085 19496
rect 19392 19456 19398 19468
rect 20073 19465 20085 19468
rect 20119 19465 20131 19499
rect 20073 19459 20131 19465
rect 23477 19499 23535 19505
rect 23477 19465 23489 19499
rect 23523 19496 23535 19499
rect 23566 19496 23572 19508
rect 23523 19468 23572 19496
rect 23523 19465 23535 19468
rect 23477 19459 23535 19465
rect 23566 19456 23572 19468
rect 23624 19456 23630 19508
rect 23658 19456 23664 19508
rect 23716 19456 23722 19508
rect 25225 19499 25283 19505
rect 25225 19465 25237 19499
rect 25271 19496 25283 19499
rect 25590 19496 25596 19508
rect 25271 19468 25596 19496
rect 25271 19465 25283 19468
rect 25225 19459 25283 19465
rect 25590 19456 25596 19468
rect 25648 19456 25654 19508
rect 12250 19428 12256 19440
rect 8996 19400 9352 19428
rect 9876 19400 11201 19428
rect 11256 19400 12256 19428
rect 8996 19388 9002 19400
rect 9398 19360 9404 19372
rect 4264 19332 4752 19360
rect 842 19252 848 19304
rect 900 19252 906 19304
rect 1118 19301 1124 19304
rect 1112 19292 1124 19301
rect 1079 19264 1124 19292
rect 1112 19255 1124 19264
rect 1118 19252 1124 19255
rect 1176 19252 1182 19304
rect 2590 19252 2596 19304
rect 2648 19252 2654 19304
rect 2777 19295 2835 19301
rect 2777 19261 2789 19295
rect 2823 19292 2835 19295
rect 2866 19292 2872 19304
rect 2823 19264 2872 19292
rect 2823 19261 2835 19264
rect 2777 19255 2835 19261
rect 2866 19252 2872 19264
rect 2924 19252 2930 19304
rect 3142 19252 3148 19304
rect 3200 19292 3206 19304
rect 3513 19295 3571 19301
rect 3513 19292 3525 19295
rect 3200 19264 3525 19292
rect 3200 19252 3206 19264
rect 3513 19261 3525 19264
rect 3559 19261 3571 19295
rect 3513 19255 3571 19261
rect 4065 19295 4123 19301
rect 4065 19261 4077 19295
rect 4111 19292 4123 19295
rect 4154 19292 4160 19304
rect 4111 19264 4160 19292
rect 4111 19261 4123 19264
rect 4065 19255 4123 19261
rect 4154 19252 4160 19264
rect 4212 19252 4218 19304
rect 3326 19224 3332 19236
rect 2240 19196 3332 19224
rect 1026 19116 1032 19168
rect 1084 19156 1090 19168
rect 2240 19165 2268 19196
rect 3326 19184 3332 19196
rect 3384 19184 3390 19236
rect 4264 19224 4292 19332
rect 4341 19295 4399 19301
rect 4341 19261 4353 19295
rect 4387 19292 4399 19295
rect 4387 19264 4568 19292
rect 4387 19261 4399 19264
rect 4341 19255 4399 19261
rect 3712 19196 4292 19224
rect 4540 19224 4568 19264
rect 4614 19252 4620 19304
rect 4672 19252 4678 19304
rect 4724 19301 4752 19332
rect 8588 19332 9404 19360
rect 4709 19295 4767 19301
rect 4709 19261 4721 19295
rect 4755 19261 4767 19295
rect 5813 19295 5871 19301
rect 4709 19255 4767 19261
rect 4816 19264 5764 19292
rect 4816 19224 4844 19264
rect 4540 19196 4844 19224
rect 2225 19159 2283 19165
rect 2225 19156 2237 19159
rect 1084 19128 2237 19156
rect 1084 19116 1090 19128
rect 2225 19125 2237 19128
rect 2271 19125 2283 19159
rect 2225 19119 2283 19125
rect 2685 19159 2743 19165
rect 2685 19125 2697 19159
rect 2731 19156 2743 19159
rect 2774 19156 2780 19168
rect 2731 19128 2780 19156
rect 2731 19125 2743 19128
rect 2685 19119 2743 19125
rect 2774 19116 2780 19128
rect 2832 19116 2838 19168
rect 3712 19165 3740 19196
rect 4982 19184 4988 19236
rect 5040 19184 5046 19236
rect 5074 19184 5080 19236
rect 5132 19184 5138 19236
rect 3697 19159 3755 19165
rect 3697 19125 3709 19159
rect 3743 19125 3755 19159
rect 3697 19119 3755 19125
rect 4246 19116 4252 19168
rect 4304 19156 4310 19168
rect 4433 19159 4491 19165
rect 4433 19156 4445 19159
rect 4304 19128 4445 19156
rect 4304 19116 4310 19128
rect 4433 19125 4445 19128
rect 4479 19125 4491 19159
rect 5000 19156 5028 19184
rect 5169 19159 5227 19165
rect 5169 19156 5181 19159
rect 5000 19128 5181 19156
rect 4433 19119 4491 19125
rect 5169 19125 5181 19128
rect 5215 19125 5227 19159
rect 5736 19156 5764 19264
rect 5813 19261 5825 19295
rect 5859 19292 5871 19295
rect 6086 19292 6092 19304
rect 5859 19264 6092 19292
rect 5859 19261 5871 19264
rect 5813 19255 5871 19261
rect 6086 19252 6092 19264
rect 6144 19252 6150 19304
rect 6270 19252 6276 19304
rect 6328 19292 6334 19304
rect 7653 19295 7711 19301
rect 7653 19292 7665 19295
rect 6328 19264 7665 19292
rect 6328 19252 6334 19264
rect 7653 19261 7665 19264
rect 7699 19292 7711 19295
rect 8018 19292 8024 19304
rect 7699 19264 8024 19292
rect 7699 19261 7711 19264
rect 7653 19255 7711 19261
rect 8018 19252 8024 19264
rect 8076 19252 8082 19304
rect 8478 19252 8484 19304
rect 8536 19292 8542 19304
rect 8588 19301 8616 19332
rect 9398 19320 9404 19332
rect 9456 19320 9462 19372
rect 8573 19295 8631 19301
rect 8573 19292 8585 19295
rect 8536 19264 8585 19292
rect 8536 19252 8542 19264
rect 8573 19261 8585 19264
rect 8619 19261 8631 19295
rect 8573 19255 8631 19261
rect 8662 19252 8668 19304
rect 8720 19252 8726 19304
rect 8754 19252 8760 19304
rect 8812 19252 8818 19304
rect 8849 19295 8907 19301
rect 8849 19261 8861 19295
rect 8895 19292 8907 19295
rect 8938 19292 8944 19304
rect 8895 19264 8944 19292
rect 8895 19261 8907 19264
rect 8849 19255 8907 19261
rect 8938 19252 8944 19264
rect 8996 19252 9002 19304
rect 9585 19295 9643 19301
rect 9585 19261 9597 19295
rect 9631 19261 9643 19295
rect 9585 19255 9643 19261
rect 9769 19295 9827 19301
rect 9769 19261 9781 19295
rect 9815 19292 9827 19295
rect 9876 19292 9904 19400
rect 11256 19372 11284 19400
rect 12250 19388 12256 19400
rect 12308 19388 12314 19440
rect 15010 19428 15016 19440
rect 13924 19400 15016 19428
rect 11238 19360 11244 19372
rect 10336 19332 11244 19360
rect 9815 19264 9904 19292
rect 9953 19295 10011 19301
rect 9815 19261 9827 19264
rect 9769 19255 9827 19261
rect 9953 19261 9965 19295
rect 9999 19292 10011 19295
rect 10336 19292 10364 19332
rect 11238 19320 11244 19332
rect 11296 19320 11302 19372
rect 13924 19360 13952 19400
rect 15010 19388 15016 19400
rect 15068 19388 15074 19440
rect 15194 19388 15200 19440
rect 15252 19388 15258 19440
rect 18598 19428 18604 19440
rect 18524 19400 18604 19428
rect 12176 19332 12388 19360
rect 9999 19264 10364 19292
rect 9999 19261 10011 19264
rect 9953 19255 10011 19261
rect 5902 19184 5908 19236
rect 5960 19224 5966 19236
rect 9033 19227 9091 19233
rect 5960 19196 8892 19224
rect 5960 19184 5966 19196
rect 8864 19168 8892 19196
rect 9033 19193 9045 19227
rect 9079 19193 9091 19227
rect 9033 19187 9091 19193
rect 8202 19156 8208 19168
rect 5736 19128 8208 19156
rect 5169 19119 5227 19125
rect 8202 19116 8208 19128
rect 8260 19116 8266 19168
rect 8386 19116 8392 19168
rect 8444 19116 8450 19168
rect 8846 19116 8852 19168
rect 8904 19116 8910 19168
rect 8938 19116 8944 19168
rect 8996 19156 9002 19168
rect 9048 19156 9076 19187
rect 8996 19128 9076 19156
rect 8996 19116 9002 19128
rect 9122 19116 9128 19168
rect 9180 19156 9186 19168
rect 9233 19159 9291 19165
rect 9233 19156 9245 19159
rect 9180 19128 9245 19156
rect 9180 19116 9186 19128
rect 9233 19125 9245 19128
rect 9279 19125 9291 19159
rect 9233 19119 9291 19125
rect 9398 19116 9404 19168
rect 9456 19116 9462 19168
rect 9600 19156 9628 19255
rect 10410 19252 10416 19304
rect 10468 19252 10474 19304
rect 10502 19252 10508 19304
rect 10560 19252 10566 19304
rect 10873 19295 10931 19301
rect 10873 19261 10885 19295
rect 10919 19292 10931 19295
rect 11054 19292 11060 19304
rect 10919 19264 11060 19292
rect 10919 19261 10931 19264
rect 10873 19255 10931 19261
rect 11054 19252 11060 19264
rect 11112 19292 11118 19304
rect 11149 19295 11207 19301
rect 11149 19292 11161 19295
rect 11112 19264 11161 19292
rect 11112 19252 11118 19264
rect 11149 19261 11161 19264
rect 11195 19261 11207 19295
rect 11149 19255 11207 19261
rect 11793 19295 11851 19301
rect 11793 19261 11805 19295
rect 11839 19292 11851 19295
rect 11885 19295 11943 19301
rect 11885 19292 11897 19295
rect 11839 19264 11897 19292
rect 11839 19261 11851 19264
rect 11793 19255 11851 19261
rect 11885 19261 11897 19264
rect 11931 19261 11943 19295
rect 12176 19292 12204 19332
rect 11885 19255 11943 19261
rect 11992 19264 12204 19292
rect 9858 19184 9864 19236
rect 9916 19184 9922 19236
rect 11992 19224 12020 19264
rect 12250 19252 12256 19304
rect 12308 19252 12314 19304
rect 12360 19292 12388 19332
rect 13004 19332 13952 19360
rect 12618 19292 12624 19304
rect 12360 19264 12624 19292
rect 12618 19252 12624 19264
rect 12676 19252 12682 19304
rect 12713 19295 12771 19301
rect 12713 19261 12725 19295
rect 12759 19292 12771 19295
rect 12802 19292 12808 19304
rect 12759 19264 12808 19292
rect 12759 19261 12771 19264
rect 12713 19255 12771 19261
rect 12802 19252 12808 19264
rect 12860 19252 12866 19304
rect 13004 19301 13032 19332
rect 12897 19295 12955 19301
rect 12897 19261 12909 19295
rect 12943 19261 12955 19295
rect 12897 19255 12955 19261
rect 12985 19295 13043 19301
rect 12985 19261 12997 19295
rect 13031 19261 13043 19295
rect 12985 19255 13043 19261
rect 10152 19196 12020 19224
rect 9950 19156 9956 19168
rect 9600 19128 9956 19156
rect 9950 19116 9956 19128
rect 10008 19116 10014 19168
rect 10152 19165 10180 19196
rect 12066 19184 12072 19236
rect 12124 19184 12130 19236
rect 12161 19227 12219 19233
rect 12161 19193 12173 19227
rect 12207 19193 12219 19227
rect 12161 19187 12219 19193
rect 10137 19159 10195 19165
rect 10137 19125 10149 19159
rect 10183 19125 10195 19159
rect 10137 19119 10195 19125
rect 10229 19159 10287 19165
rect 10229 19125 10241 19159
rect 10275 19156 10287 19159
rect 10318 19156 10324 19168
rect 10275 19128 10324 19156
rect 10275 19125 10287 19128
rect 10229 19119 10287 19125
rect 10318 19116 10324 19128
rect 10376 19116 10382 19168
rect 11146 19116 11152 19168
rect 11204 19156 11210 19168
rect 11974 19156 11980 19168
rect 11204 19128 11980 19156
rect 11204 19116 11210 19128
rect 11974 19116 11980 19128
rect 12032 19156 12038 19168
rect 12176 19156 12204 19187
rect 12032 19128 12204 19156
rect 12032 19116 12038 19128
rect 12250 19116 12256 19168
rect 12308 19156 12314 19168
rect 12437 19159 12495 19165
rect 12437 19156 12449 19159
rect 12308 19128 12449 19156
rect 12308 19116 12314 19128
rect 12437 19125 12449 19128
rect 12483 19125 12495 19159
rect 12912 19156 12940 19255
rect 13538 19252 13544 19304
rect 13596 19292 13602 19304
rect 13924 19301 13952 19332
rect 14645 19363 14703 19369
rect 14645 19329 14657 19363
rect 14691 19360 14703 19363
rect 14921 19363 14979 19369
rect 14921 19360 14933 19363
rect 14691 19332 14933 19360
rect 14691 19329 14703 19332
rect 14645 19323 14703 19329
rect 14921 19329 14933 19332
rect 14967 19360 14979 19363
rect 15212 19360 15240 19388
rect 14967 19332 15332 19360
rect 14967 19329 14979 19332
rect 14921 19323 14979 19329
rect 13633 19295 13691 19301
rect 13633 19292 13645 19295
rect 13596 19264 13645 19292
rect 13596 19252 13602 19264
rect 13633 19261 13645 19264
rect 13679 19292 13691 19295
rect 13909 19295 13967 19301
rect 13679 19264 13860 19292
rect 13679 19261 13691 19264
rect 13633 19255 13691 19261
rect 13832 19224 13860 19264
rect 13909 19261 13921 19295
rect 13955 19261 13967 19295
rect 13909 19255 13967 19261
rect 15197 19295 15255 19301
rect 15197 19261 15209 19295
rect 15243 19261 15255 19295
rect 15197 19255 15255 19261
rect 14918 19224 14924 19236
rect 13832 19196 14924 19224
rect 14918 19184 14924 19196
rect 14976 19224 14982 19236
rect 15013 19227 15071 19233
rect 15013 19224 15025 19227
rect 14976 19196 15025 19224
rect 14976 19184 14982 19196
rect 15013 19193 15025 19196
rect 15059 19193 15071 19227
rect 15013 19187 15071 19193
rect 13538 19156 13544 19168
rect 12912 19128 13544 19156
rect 12437 19119 12495 19125
rect 13538 19116 13544 19128
rect 13596 19116 13602 19168
rect 13633 19159 13691 19165
rect 13633 19125 13645 19159
rect 13679 19156 13691 19159
rect 13722 19156 13728 19168
rect 13679 19128 13728 19156
rect 13679 19125 13691 19128
rect 13633 19119 13691 19125
rect 13722 19116 13728 19128
rect 13780 19116 13786 19168
rect 14274 19116 14280 19168
rect 14332 19156 14338 19168
rect 15102 19156 15108 19168
rect 14332 19128 15108 19156
rect 14332 19116 14338 19128
rect 15102 19116 15108 19128
rect 15160 19156 15166 19168
rect 15212 19156 15240 19255
rect 15304 19224 15332 19332
rect 15378 19320 15384 19372
rect 15436 19320 15442 19372
rect 15838 19360 15844 19372
rect 15488 19332 15844 19360
rect 15488 19304 15516 19332
rect 15838 19320 15844 19332
rect 15896 19320 15902 19372
rect 17862 19320 17868 19372
rect 17920 19320 17926 19372
rect 18524 19369 18552 19400
rect 18598 19388 18604 19400
rect 18656 19428 18662 19440
rect 22738 19428 22744 19440
rect 18656 19400 22744 19428
rect 18656 19388 18662 19400
rect 22738 19388 22744 19400
rect 22796 19388 22802 19440
rect 25041 19431 25099 19437
rect 25041 19397 25053 19431
rect 25087 19397 25099 19431
rect 25041 19391 25099 19397
rect 18509 19363 18567 19369
rect 18509 19329 18521 19363
rect 18555 19329 18567 19363
rect 18509 19323 18567 19329
rect 19610 19320 19616 19372
rect 19668 19360 19674 19372
rect 21177 19363 21235 19369
rect 21177 19360 21189 19363
rect 19668 19332 21189 19360
rect 19668 19320 19674 19332
rect 21177 19329 21189 19332
rect 21223 19360 21235 19363
rect 21818 19360 21824 19372
rect 21223 19332 21824 19360
rect 21223 19329 21235 19332
rect 21177 19323 21235 19329
rect 21818 19320 21824 19332
rect 21876 19320 21882 19372
rect 22094 19320 22100 19372
rect 22152 19320 22158 19372
rect 24581 19363 24639 19369
rect 24581 19329 24593 19363
rect 24627 19329 24639 19363
rect 24581 19323 24639 19329
rect 15470 19252 15476 19304
rect 15528 19252 15534 19304
rect 15562 19252 15568 19304
rect 15620 19252 15626 19304
rect 16114 19301 16120 19304
rect 16108 19292 16120 19301
rect 16075 19264 16120 19292
rect 16108 19255 16120 19264
rect 16114 19252 16120 19255
rect 16172 19252 16178 19304
rect 17586 19252 17592 19304
rect 17644 19292 17650 19304
rect 17773 19295 17831 19301
rect 17773 19292 17785 19295
rect 17644 19264 17785 19292
rect 17644 19252 17650 19264
rect 17773 19261 17785 19264
rect 17819 19261 17831 19295
rect 17773 19255 17831 19261
rect 18046 19252 18052 19304
rect 18104 19252 18110 19304
rect 18322 19252 18328 19304
rect 18380 19252 18386 19304
rect 19702 19252 19708 19304
rect 19760 19292 19766 19304
rect 21085 19295 21143 19301
rect 21085 19292 21097 19295
rect 19760 19264 21097 19292
rect 19760 19252 19766 19264
rect 21085 19261 21097 19264
rect 21131 19261 21143 19295
rect 21085 19255 21143 19261
rect 22278 19252 22284 19304
rect 22336 19252 22342 19304
rect 22462 19252 22468 19304
rect 22520 19252 22526 19304
rect 22554 19252 22560 19304
rect 22612 19252 22618 19304
rect 22925 19295 22983 19301
rect 22925 19261 22937 19295
rect 22971 19261 22983 19295
rect 22925 19255 22983 19261
rect 23201 19295 23259 19301
rect 23201 19261 23213 19295
rect 23247 19292 23259 19295
rect 24026 19292 24032 19304
rect 23247 19264 24032 19292
rect 23247 19261 23259 19264
rect 23201 19255 23259 19261
rect 17681 19227 17739 19233
rect 15304 19196 16528 19224
rect 16500 19168 16528 19196
rect 17681 19193 17693 19227
rect 17727 19224 17739 19227
rect 18064 19224 18092 19252
rect 18785 19227 18843 19233
rect 18785 19224 18797 19227
rect 17727 19196 17991 19224
rect 18064 19196 18797 19224
rect 17727 19193 17739 19196
rect 17681 19187 17739 19193
rect 15160 19128 15240 19156
rect 15160 19116 15166 19128
rect 16482 19116 16488 19168
rect 16540 19156 16546 19168
rect 17221 19159 17279 19165
rect 17221 19156 17233 19159
rect 16540 19128 17233 19156
rect 16540 19116 16546 19128
rect 17221 19125 17233 19128
rect 17267 19125 17279 19159
rect 17963 19156 17991 19196
rect 18785 19193 18797 19196
rect 18831 19224 18843 19227
rect 19978 19224 19984 19236
rect 18831 19196 19984 19224
rect 18831 19193 18843 19196
rect 18785 19187 18843 19193
rect 19978 19184 19984 19196
rect 20036 19184 20042 19236
rect 22940 19224 22968 19255
rect 24026 19252 24032 19264
rect 24084 19252 24090 19304
rect 24305 19295 24363 19301
rect 24305 19261 24317 19295
rect 24351 19292 24363 19295
rect 24486 19292 24492 19304
rect 24351 19264 24492 19292
rect 24351 19261 24363 19264
rect 24305 19255 24363 19261
rect 24486 19252 24492 19264
rect 24544 19292 24550 19304
rect 24596 19292 24624 19323
rect 24544 19264 24624 19292
rect 24673 19295 24731 19301
rect 24544 19252 24550 19264
rect 24673 19261 24685 19295
rect 24719 19261 24731 19295
rect 25056 19292 25084 19391
rect 25133 19295 25191 19301
rect 25133 19292 25145 19295
rect 25056 19264 25145 19292
rect 24673 19255 24731 19261
rect 25133 19261 25145 19264
rect 25179 19261 25191 19295
rect 25133 19255 25191 19261
rect 23293 19227 23351 19233
rect 22940 19196 23244 19224
rect 18141 19159 18199 19165
rect 18141 19156 18153 19159
rect 17963 19128 18153 19156
rect 17221 19119 17279 19125
rect 18141 19125 18153 19128
rect 18187 19125 18199 19159
rect 18141 19119 18199 19125
rect 20438 19116 20444 19168
rect 20496 19156 20502 19168
rect 20625 19159 20683 19165
rect 20625 19156 20637 19159
rect 20496 19128 20637 19156
rect 20496 19116 20502 19128
rect 20625 19125 20637 19128
rect 20671 19125 20683 19159
rect 20625 19119 20683 19125
rect 20990 19116 20996 19168
rect 21048 19116 21054 19168
rect 22830 19116 22836 19168
rect 22888 19116 22894 19168
rect 23106 19116 23112 19168
rect 23164 19116 23170 19168
rect 23216 19156 23244 19196
rect 23293 19193 23305 19227
rect 23339 19224 23351 19227
rect 23382 19224 23388 19236
rect 23339 19196 23388 19224
rect 23339 19193 23351 19196
rect 23293 19187 23351 19193
rect 23382 19184 23388 19196
rect 23440 19184 23446 19236
rect 23509 19227 23567 19233
rect 23509 19193 23521 19227
rect 23555 19224 23567 19227
rect 23845 19227 23903 19233
rect 23845 19224 23857 19227
rect 23555 19196 23857 19224
rect 23555 19193 23567 19196
rect 23509 19187 23567 19193
rect 23845 19193 23857 19196
rect 23891 19193 23903 19227
rect 24688 19224 24716 19255
rect 25222 19252 25228 19304
rect 25280 19292 25286 19304
rect 25317 19295 25375 19301
rect 25317 19292 25329 19295
rect 25280 19264 25329 19292
rect 25280 19252 25286 19264
rect 25317 19261 25329 19264
rect 25363 19261 25375 19295
rect 25317 19255 25375 19261
rect 25774 19252 25780 19304
rect 25832 19292 25838 19304
rect 26234 19292 26240 19304
rect 25832 19264 26240 19292
rect 25832 19252 25838 19264
rect 26234 19252 26240 19264
rect 26292 19292 26298 19304
rect 26789 19295 26847 19301
rect 26789 19292 26801 19295
rect 26292 19264 26801 19292
rect 26292 19252 26298 19264
rect 26789 19261 26801 19264
rect 26835 19261 26847 19295
rect 26789 19255 26847 19261
rect 24688 19196 25544 19224
rect 23845 19187 23903 19193
rect 24213 19159 24271 19165
rect 24213 19156 24225 19159
rect 23216 19128 24225 19156
rect 24213 19125 24225 19128
rect 24259 19156 24271 19159
rect 24670 19156 24676 19168
rect 24259 19128 24676 19156
rect 24259 19125 24271 19128
rect 24213 19119 24271 19125
rect 24670 19116 24676 19128
rect 24728 19116 24734 19168
rect 24854 19116 24860 19168
rect 24912 19156 24918 19168
rect 25409 19159 25467 19165
rect 25409 19156 25421 19159
rect 24912 19128 25421 19156
rect 24912 19116 24918 19128
rect 25409 19125 25421 19128
rect 25455 19125 25467 19159
rect 25516 19156 25544 19196
rect 25866 19184 25872 19236
rect 25924 19224 25930 19236
rect 26522 19227 26580 19233
rect 26522 19224 26534 19227
rect 25924 19196 26534 19224
rect 25924 19184 25930 19196
rect 26522 19193 26534 19196
rect 26568 19193 26580 19227
rect 26522 19187 26580 19193
rect 26418 19156 26424 19168
rect 25516 19128 26424 19156
rect 25409 19119 25467 19125
rect 26418 19116 26424 19128
rect 26476 19116 26482 19168
rect 552 19066 27576 19088
rect 552 19014 7114 19066
rect 7166 19014 7178 19066
rect 7230 19014 7242 19066
rect 7294 19014 7306 19066
rect 7358 19014 7370 19066
rect 7422 19014 13830 19066
rect 13882 19014 13894 19066
rect 13946 19014 13958 19066
rect 14010 19014 14022 19066
rect 14074 19014 14086 19066
rect 14138 19014 20546 19066
rect 20598 19014 20610 19066
rect 20662 19014 20674 19066
rect 20726 19014 20738 19066
rect 20790 19014 20802 19066
rect 20854 19014 27262 19066
rect 27314 19014 27326 19066
rect 27378 19014 27390 19066
rect 27442 19014 27454 19066
rect 27506 19014 27518 19066
rect 27570 19014 27576 19066
rect 552 18992 27576 19014
rect 1394 18912 1400 18964
rect 1452 18952 1458 18964
rect 1489 18955 1547 18961
rect 1489 18952 1501 18955
rect 1452 18924 1501 18952
rect 1452 18912 1458 18924
rect 1489 18921 1501 18924
rect 1535 18921 1547 18955
rect 1489 18915 1547 18921
rect 1946 18912 1952 18964
rect 2004 18952 2010 18964
rect 2590 18952 2596 18964
rect 2004 18924 2596 18952
rect 2004 18912 2010 18924
rect 2590 18912 2596 18924
rect 2648 18912 2654 18964
rect 5074 18912 5080 18964
rect 5132 18952 5138 18964
rect 5445 18955 5503 18961
rect 5445 18952 5457 18955
rect 5132 18924 5457 18952
rect 5132 18912 5138 18924
rect 5445 18921 5457 18924
rect 5491 18921 5503 18955
rect 5445 18915 5503 18921
rect 7558 18912 7564 18964
rect 7616 18952 7622 18964
rect 8113 18955 8171 18961
rect 8113 18952 8125 18955
rect 7616 18924 8125 18952
rect 7616 18912 7622 18924
rect 8113 18921 8125 18924
rect 8159 18921 8171 18955
rect 8113 18915 8171 18921
rect 8757 18955 8815 18961
rect 8757 18921 8769 18955
rect 8803 18952 8815 18955
rect 9214 18952 9220 18964
rect 8803 18924 9220 18952
rect 8803 18921 8815 18924
rect 8757 18915 8815 18921
rect 2676 18887 2734 18893
rect 860 18856 2452 18884
rect 860 18828 888 18856
rect 842 18776 848 18828
rect 900 18776 906 18828
rect 1026 18776 1032 18828
rect 1084 18776 1090 18828
rect 2133 18819 2191 18825
rect 2133 18785 2145 18819
rect 2179 18816 2191 18819
rect 2222 18816 2228 18828
rect 2179 18788 2228 18816
rect 2179 18785 2191 18788
rect 2133 18779 2191 18785
rect 2222 18776 2228 18788
rect 2280 18776 2286 18828
rect 2424 18825 2452 18856
rect 2676 18853 2688 18887
rect 2722 18884 2734 18887
rect 2774 18884 2780 18896
rect 2722 18856 2780 18884
rect 2722 18853 2734 18856
rect 2676 18847 2734 18853
rect 2774 18844 2780 18856
rect 2832 18844 2838 18896
rect 8128 18884 8156 18915
rect 9214 18912 9220 18924
rect 9272 18912 9278 18964
rect 9398 18912 9404 18964
rect 9456 18912 9462 18964
rect 10321 18955 10379 18961
rect 10321 18952 10333 18955
rect 10152 18924 10333 18952
rect 8662 18884 8668 18896
rect 3988 18856 6224 18884
rect 8128 18856 8668 18884
rect 3988 18825 4016 18856
rect 4246 18825 4252 18828
rect 2409 18819 2467 18825
rect 2409 18785 2421 18819
rect 2455 18785 2467 18819
rect 2409 18779 2467 18785
rect 3973 18819 4031 18825
rect 3973 18785 3985 18819
rect 4019 18785 4031 18819
rect 4240 18816 4252 18825
rect 4207 18788 4252 18816
rect 3973 18779 4031 18785
rect 4240 18779 4252 18788
rect 4246 18776 4252 18779
rect 4304 18776 4310 18828
rect 5442 18776 5448 18828
rect 5500 18776 5506 18828
rect 6196 18825 6224 18856
rect 8662 18844 8668 18856
rect 8720 18844 8726 18896
rect 5629 18819 5687 18825
rect 5629 18785 5641 18819
rect 5675 18785 5687 18819
rect 5629 18779 5687 18785
rect 6181 18819 6239 18825
rect 6181 18785 6193 18819
rect 6227 18816 6239 18819
rect 6270 18816 6276 18828
rect 6227 18788 6276 18816
rect 6227 18785 6239 18788
rect 6181 18779 6239 18785
rect 2317 18751 2375 18757
rect 2317 18717 2329 18751
rect 2363 18717 2375 18751
rect 5644 18748 5672 18779
rect 6270 18776 6276 18788
rect 6328 18776 6334 18828
rect 6454 18825 6460 18828
rect 6448 18816 6460 18825
rect 6415 18788 6460 18816
rect 6448 18779 6460 18788
rect 6454 18776 6460 18779
rect 6512 18776 6518 18828
rect 8021 18819 8079 18825
rect 8021 18785 8033 18819
rect 8067 18785 8079 18819
rect 8021 18779 8079 18785
rect 8205 18819 8263 18825
rect 8205 18785 8217 18819
rect 8251 18785 8263 18819
rect 8205 18779 8263 18785
rect 8481 18819 8539 18825
rect 8481 18785 8493 18819
rect 8527 18816 8539 18819
rect 8570 18816 8576 18828
rect 8527 18788 8576 18816
rect 8527 18785 8539 18788
rect 8481 18779 8539 18785
rect 5644 18720 6224 18748
rect 2317 18711 2375 18717
rect 1394 18640 1400 18692
rect 1452 18640 1458 18692
rect 2332 18612 2360 18711
rect 5810 18680 5816 18692
rect 4908 18652 5816 18680
rect 3602 18612 3608 18624
rect 2332 18584 3608 18612
rect 3602 18572 3608 18584
rect 3660 18612 3666 18624
rect 3789 18615 3847 18621
rect 3789 18612 3801 18615
rect 3660 18584 3801 18612
rect 3660 18572 3666 18584
rect 3789 18581 3801 18584
rect 3835 18581 3847 18615
rect 3789 18575 3847 18581
rect 4154 18572 4160 18624
rect 4212 18612 4218 18624
rect 4908 18612 4936 18652
rect 5810 18640 5816 18652
rect 5868 18640 5874 18692
rect 4212 18584 4936 18612
rect 5353 18615 5411 18621
rect 4212 18572 4218 18584
rect 5353 18581 5365 18615
rect 5399 18612 5411 18615
rect 6086 18612 6092 18624
rect 5399 18584 6092 18612
rect 5399 18581 5411 18584
rect 5353 18575 5411 18581
rect 6086 18572 6092 18584
rect 6144 18572 6150 18624
rect 6196 18612 6224 18720
rect 8036 18680 8064 18779
rect 8220 18748 8248 18779
rect 8570 18776 8576 18788
rect 8628 18776 8634 18828
rect 8754 18776 8760 18828
rect 8812 18816 8818 18828
rect 9416 18816 9444 18912
rect 9984 18887 10042 18893
rect 9984 18853 9996 18887
rect 10030 18884 10042 18887
rect 10152 18884 10180 18924
rect 10321 18921 10333 18924
rect 10367 18921 10379 18955
rect 10321 18915 10379 18921
rect 11054 18912 11060 18964
rect 11112 18912 11118 18964
rect 12342 18912 12348 18964
rect 12400 18952 12406 18964
rect 13722 18952 13728 18964
rect 12400 18924 13728 18952
rect 12400 18912 12406 18924
rect 13722 18912 13728 18924
rect 13780 18912 13786 18964
rect 14274 18912 14280 18964
rect 14332 18952 14338 18964
rect 14645 18955 14703 18961
rect 14645 18952 14657 18955
rect 14332 18924 14657 18952
rect 14332 18912 14338 18924
rect 14645 18921 14657 18924
rect 14691 18921 14703 18955
rect 14645 18915 14703 18921
rect 15562 18912 15568 18964
rect 15620 18952 15626 18964
rect 16117 18955 16175 18961
rect 16117 18952 16129 18955
rect 15620 18924 16129 18952
rect 15620 18912 15626 18924
rect 16117 18921 16129 18924
rect 16163 18921 16175 18955
rect 16117 18915 16175 18921
rect 16482 18912 16488 18964
rect 16540 18952 16546 18964
rect 16577 18955 16635 18961
rect 16577 18952 16589 18955
rect 16540 18924 16589 18952
rect 16540 18912 16546 18924
rect 16577 18921 16589 18924
rect 16623 18921 16635 18955
rect 17586 18952 17592 18964
rect 16577 18915 16635 18921
rect 16684 18924 17592 18952
rect 14553 18887 14611 18893
rect 10030 18856 10180 18884
rect 10244 18856 12480 18884
rect 10030 18853 10042 18856
rect 9984 18847 10042 18853
rect 10244 18828 10272 18856
rect 12452 18828 12480 18856
rect 13740 18856 14320 18884
rect 8812 18788 9168 18816
rect 9416 18788 10180 18816
rect 8812 18776 8818 18788
rect 8772 18748 8800 18776
rect 8220 18720 8800 18748
rect 8202 18680 8208 18692
rect 8036 18652 8208 18680
rect 8202 18640 8208 18652
rect 8260 18640 8266 18692
rect 8294 18640 8300 18692
rect 8352 18680 8358 18692
rect 8389 18683 8447 18689
rect 8389 18680 8401 18683
rect 8352 18652 8401 18680
rect 8352 18640 8358 18652
rect 8389 18649 8401 18652
rect 8435 18680 8447 18683
rect 9030 18680 9036 18692
rect 8435 18652 9036 18680
rect 8435 18649 8447 18652
rect 8389 18643 8447 18649
rect 9030 18640 9036 18652
rect 9088 18640 9094 18692
rect 6914 18612 6920 18624
rect 6196 18584 6920 18612
rect 6914 18572 6920 18584
rect 6972 18572 6978 18624
rect 7834 18572 7840 18624
rect 7892 18572 7898 18624
rect 8849 18615 8907 18621
rect 8849 18581 8861 18615
rect 8895 18612 8907 18615
rect 9140 18612 9168 18788
rect 10152 18748 10180 18788
rect 10226 18776 10232 18828
rect 10284 18776 10290 18828
rect 10505 18819 10563 18825
rect 10505 18785 10517 18819
rect 10551 18785 10563 18819
rect 10505 18779 10563 18785
rect 10520 18748 10548 18779
rect 12158 18776 12164 18828
rect 12216 18825 12222 18828
rect 12216 18819 12239 18825
rect 12227 18785 12239 18819
rect 12216 18779 12239 18785
rect 12216 18776 12222 18779
rect 12434 18776 12440 18828
rect 12492 18776 12498 18828
rect 12526 18776 12532 18828
rect 12584 18776 12590 18828
rect 13740 18825 13768 18856
rect 13725 18819 13783 18825
rect 13725 18785 13737 18819
rect 13771 18785 13783 18819
rect 13725 18779 13783 18785
rect 13909 18819 13967 18825
rect 13909 18785 13921 18819
rect 13955 18816 13967 18819
rect 14292 18816 14320 18856
rect 14553 18853 14565 18887
rect 14599 18884 14611 18887
rect 14918 18884 14924 18896
rect 14599 18856 14924 18884
rect 14599 18853 14611 18856
rect 14553 18847 14611 18853
rect 14918 18844 14924 18856
rect 14976 18884 14982 18896
rect 16684 18884 16712 18924
rect 17586 18912 17592 18924
rect 17644 18912 17650 18964
rect 20438 18912 20444 18964
rect 20496 18912 20502 18964
rect 20717 18955 20775 18961
rect 20717 18921 20729 18955
rect 20763 18952 20775 18955
rect 20990 18952 20996 18964
rect 20763 18924 20996 18952
rect 20763 18921 20775 18924
rect 20717 18915 20775 18921
rect 20990 18912 20996 18924
rect 21048 18912 21054 18964
rect 21910 18912 21916 18964
rect 21968 18952 21974 18964
rect 21968 18924 22324 18952
rect 21968 18912 21974 18924
rect 17954 18884 17960 18896
rect 14976 18856 16712 18884
rect 17328 18856 17960 18884
rect 14976 18844 14982 18856
rect 15378 18816 15384 18828
rect 13955 18788 14228 18816
rect 14292 18788 15384 18816
rect 13955 18785 13967 18788
rect 13909 18779 13967 18785
rect 10152 18720 10548 18748
rect 10226 18640 10232 18692
rect 10284 18680 10290 18692
rect 10410 18680 10416 18692
rect 10284 18652 10416 18680
rect 10284 18640 10290 18652
rect 10410 18640 10416 18652
rect 10468 18680 10474 18692
rect 14200 18689 14228 18788
rect 14568 18760 14596 18788
rect 15378 18776 15384 18788
rect 15436 18776 15442 18828
rect 16485 18819 16543 18825
rect 16485 18785 16497 18819
rect 16531 18816 16543 18819
rect 16531 18788 16988 18816
rect 16531 18785 16543 18788
rect 16485 18779 16543 18785
rect 14550 18708 14556 18760
rect 14608 18708 14614 18760
rect 14642 18708 14648 18760
rect 14700 18748 14706 18760
rect 14737 18751 14795 18757
rect 14737 18748 14749 18751
rect 14700 18720 14749 18748
rect 14700 18708 14706 18720
rect 14737 18717 14749 18720
rect 14783 18748 14795 18751
rect 16669 18751 16727 18757
rect 16669 18748 16681 18751
rect 14783 18720 16681 18748
rect 14783 18717 14795 18720
rect 14737 18711 14795 18717
rect 16669 18717 16681 18720
rect 16715 18717 16727 18751
rect 16669 18711 16727 18717
rect 14185 18683 14243 18689
rect 10468 18652 10824 18680
rect 10468 18640 10474 18652
rect 9306 18612 9312 18624
rect 8895 18584 9312 18612
rect 8895 18581 8907 18584
rect 8849 18575 8907 18581
rect 9306 18572 9312 18584
rect 9364 18612 9370 18624
rect 10502 18612 10508 18624
rect 9364 18584 10508 18612
rect 9364 18572 9370 18584
rect 10502 18572 10508 18584
rect 10560 18572 10566 18624
rect 10796 18612 10824 18652
rect 14185 18649 14197 18683
rect 14231 18649 14243 18683
rect 14185 18643 14243 18649
rect 12621 18615 12679 18621
rect 12621 18612 12633 18615
rect 10796 18584 12633 18612
rect 12621 18581 12633 18584
rect 12667 18581 12679 18615
rect 12621 18575 12679 18581
rect 14093 18615 14151 18621
rect 14093 18581 14105 18615
rect 14139 18612 14151 18615
rect 14274 18612 14280 18624
rect 14139 18584 14280 18612
rect 14139 18581 14151 18584
rect 14093 18575 14151 18581
rect 14274 18572 14280 18584
rect 14332 18572 14338 18624
rect 16960 18612 16988 18788
rect 17034 18776 17040 18828
rect 17092 18776 17098 18828
rect 17328 18825 17356 18856
rect 17954 18844 17960 18856
rect 18012 18884 18018 18896
rect 19334 18884 19340 18896
rect 18012 18856 19340 18884
rect 18012 18844 18018 18856
rect 18984 18825 19012 18856
rect 19334 18844 19340 18856
rect 19392 18844 19398 18896
rect 20346 18844 20352 18896
rect 20404 18844 20410 18896
rect 17313 18819 17371 18825
rect 17313 18785 17325 18819
rect 17359 18785 17371 18819
rect 17569 18819 17627 18825
rect 17569 18816 17581 18819
rect 17313 18779 17371 18785
rect 17420 18788 17581 18816
rect 17420 18748 17448 18788
rect 17569 18785 17581 18788
rect 17615 18785 17627 18819
rect 17569 18779 17627 18785
rect 18969 18819 19027 18825
rect 18969 18785 18981 18819
rect 19015 18785 19027 18819
rect 18969 18779 19027 18785
rect 19236 18819 19294 18825
rect 19236 18785 19248 18819
rect 19282 18816 19294 18819
rect 20364 18816 20392 18844
rect 19282 18788 20392 18816
rect 20456 18816 20484 18912
rect 22296 18884 22324 18924
rect 22554 18912 22560 18964
rect 22612 18912 22618 18964
rect 23106 18912 23112 18964
rect 23164 18912 23170 18964
rect 24026 18912 24032 18964
rect 24084 18952 24090 18964
rect 24305 18955 24363 18961
rect 24305 18952 24317 18955
rect 24084 18924 24317 18952
rect 24084 18912 24090 18924
rect 24305 18921 24317 18924
rect 24351 18952 24363 18955
rect 24581 18955 24639 18961
rect 24581 18952 24593 18955
rect 24351 18924 24593 18952
rect 24351 18921 24363 18924
rect 24305 18915 24363 18921
rect 24581 18921 24593 18924
rect 24627 18921 24639 18955
rect 24581 18915 24639 18921
rect 24670 18912 24676 18964
rect 24728 18952 24734 18964
rect 25593 18955 25651 18961
rect 24728 18924 25544 18952
rect 24728 18912 24734 18924
rect 23124 18884 23152 18912
rect 20824 18856 22140 18884
rect 20625 18819 20683 18825
rect 20625 18816 20637 18819
rect 20456 18788 20637 18816
rect 19282 18785 19294 18788
rect 19236 18779 19294 18785
rect 20625 18785 20637 18788
rect 20671 18785 20683 18819
rect 20625 18779 20683 18785
rect 17236 18720 17448 18748
rect 17236 18689 17264 18720
rect 20254 18708 20260 18760
rect 20312 18748 20318 18760
rect 20824 18748 20852 18856
rect 20898 18776 20904 18828
rect 20956 18776 20962 18828
rect 22112 18825 22140 18856
rect 22296 18856 23152 18884
rect 23192 18887 23250 18893
rect 21913 18819 21971 18825
rect 21913 18785 21925 18819
rect 21959 18785 21971 18819
rect 21913 18779 21971 18785
rect 22097 18819 22155 18825
rect 22097 18785 22109 18819
rect 22143 18785 22155 18819
rect 22097 18779 22155 18785
rect 20312 18720 20852 18748
rect 20312 18708 20318 18720
rect 21082 18708 21088 18760
rect 21140 18708 21146 18760
rect 17221 18683 17279 18689
rect 17221 18649 17233 18683
rect 17267 18649 17279 18683
rect 20272 18680 20300 18708
rect 20349 18683 20407 18689
rect 20349 18680 20361 18683
rect 17221 18643 17279 18649
rect 18248 18652 18828 18680
rect 20272 18652 20361 18680
rect 18248 18624 18276 18652
rect 18230 18612 18236 18624
rect 16960 18584 18236 18612
rect 18230 18572 18236 18584
rect 18288 18572 18294 18624
rect 18690 18572 18696 18624
rect 18748 18572 18754 18624
rect 18800 18612 18828 18652
rect 20349 18649 20361 18652
rect 20395 18649 20407 18683
rect 21928 18680 21956 18779
rect 22186 18776 22192 18828
rect 22244 18776 22250 18828
rect 22296 18825 22324 18856
rect 23192 18853 23204 18887
rect 23238 18884 23250 18887
rect 23474 18884 23480 18896
rect 23238 18856 23480 18884
rect 23238 18853 23250 18856
rect 23192 18847 23250 18853
rect 23474 18844 23480 18856
rect 23532 18844 23538 18896
rect 24854 18844 24860 18896
rect 24912 18844 24918 18896
rect 25409 18887 25467 18893
rect 25409 18853 25421 18887
rect 25455 18853 25467 18887
rect 25409 18847 25467 18853
rect 22281 18819 22339 18825
rect 22281 18785 22293 18819
rect 22327 18785 22339 18819
rect 22281 18779 22339 18785
rect 22925 18819 22983 18825
rect 22925 18785 22937 18819
rect 22971 18816 22983 18819
rect 23014 18816 23020 18828
rect 22971 18788 23020 18816
rect 22971 18785 22983 18788
rect 22925 18779 22983 18785
rect 23014 18776 23020 18788
rect 23072 18776 23078 18828
rect 24302 18776 24308 18828
rect 24360 18816 24366 18828
rect 24765 18819 24823 18825
rect 24596 18816 24777 18819
rect 24360 18791 24777 18816
rect 24360 18788 24624 18791
rect 24360 18776 24366 18788
rect 24765 18785 24777 18791
rect 24811 18785 24823 18819
rect 24765 18779 24823 18785
rect 24397 18751 24455 18757
rect 24397 18717 24409 18751
rect 24443 18748 24455 18751
rect 24486 18748 24492 18760
rect 24443 18720 24492 18748
rect 24443 18717 24455 18720
rect 24397 18711 24455 18717
rect 24486 18708 24492 18720
rect 24544 18748 24550 18760
rect 24872 18748 24900 18844
rect 24544 18720 24900 18748
rect 24544 18708 24550 18720
rect 22830 18680 22836 18692
rect 21928 18652 22836 18680
rect 20349 18643 20407 18649
rect 22830 18640 22836 18652
rect 22888 18640 22894 18692
rect 24854 18640 24860 18692
rect 24912 18680 24918 18692
rect 24949 18683 25007 18689
rect 24949 18680 24961 18683
rect 24912 18652 24961 18680
rect 24912 18640 24918 18652
rect 24949 18649 24961 18652
rect 24995 18680 25007 18683
rect 25041 18683 25099 18689
rect 25041 18680 25053 18683
rect 24995 18652 25053 18680
rect 24995 18649 25007 18652
rect 24949 18643 25007 18649
rect 25041 18649 25053 18652
rect 25087 18649 25099 18683
rect 25424 18680 25452 18847
rect 25516 18748 25544 18924
rect 25593 18921 25605 18955
rect 25639 18921 25651 18955
rect 25593 18915 25651 18921
rect 25608 18816 25636 18915
rect 25866 18912 25872 18964
rect 25924 18912 25930 18964
rect 25685 18819 25743 18825
rect 25685 18816 25697 18819
rect 25608 18788 25697 18816
rect 25685 18785 25697 18788
rect 25731 18785 25743 18819
rect 25685 18779 25743 18785
rect 27062 18748 27068 18760
rect 25516 18720 27068 18748
rect 27062 18708 27068 18720
rect 27120 18708 27126 18760
rect 25041 18643 25099 18649
rect 25128 18652 25452 18680
rect 19702 18612 19708 18624
rect 18800 18584 19708 18612
rect 19702 18572 19708 18584
rect 19760 18572 19766 18624
rect 20438 18572 20444 18624
rect 20496 18572 20502 18624
rect 21174 18572 21180 18624
rect 21232 18612 21238 18624
rect 22186 18612 22192 18624
rect 21232 18584 22192 18612
rect 21232 18572 21238 18584
rect 22186 18572 22192 18584
rect 22244 18572 22250 18624
rect 24762 18572 24768 18624
rect 24820 18612 24826 18624
rect 25128 18612 25156 18652
rect 24820 18584 25156 18612
rect 24820 18572 24826 18584
rect 25406 18572 25412 18624
rect 25464 18572 25470 18624
rect 552 18522 27416 18544
rect 552 18470 3756 18522
rect 3808 18470 3820 18522
rect 3872 18470 3884 18522
rect 3936 18470 3948 18522
rect 4000 18470 4012 18522
rect 4064 18470 10472 18522
rect 10524 18470 10536 18522
rect 10588 18470 10600 18522
rect 10652 18470 10664 18522
rect 10716 18470 10728 18522
rect 10780 18470 17188 18522
rect 17240 18470 17252 18522
rect 17304 18470 17316 18522
rect 17368 18470 17380 18522
rect 17432 18470 17444 18522
rect 17496 18470 23904 18522
rect 23956 18470 23968 18522
rect 24020 18470 24032 18522
rect 24084 18470 24096 18522
rect 24148 18470 24160 18522
rect 24212 18470 27416 18522
rect 552 18448 27416 18470
rect 2777 18411 2835 18417
rect 2777 18377 2789 18411
rect 2823 18408 2835 18411
rect 2866 18408 2872 18420
rect 2823 18380 2872 18408
rect 2823 18377 2835 18380
rect 2777 18371 2835 18377
rect 2866 18368 2872 18380
rect 2924 18368 2930 18420
rect 3160 18380 5212 18408
rect 3160 18352 3188 18380
rect 2406 18300 2412 18352
rect 2464 18300 2470 18352
rect 3050 18340 3056 18352
rect 2700 18312 3056 18340
rect 1946 18232 1952 18284
rect 2004 18232 2010 18284
rect 2424 18272 2452 18300
rect 2700 18281 2728 18312
rect 3050 18300 3056 18312
rect 3108 18300 3114 18352
rect 3142 18300 3148 18352
rect 3200 18300 3206 18352
rect 3418 18300 3424 18352
rect 3476 18340 3482 18352
rect 3602 18340 3608 18352
rect 3476 18312 3608 18340
rect 3476 18300 3482 18312
rect 3602 18300 3608 18312
rect 3660 18340 3666 18352
rect 5184 18349 5212 18380
rect 6454 18368 6460 18420
rect 6512 18408 6518 18420
rect 6549 18411 6607 18417
rect 6549 18408 6561 18411
rect 6512 18380 6561 18408
rect 6512 18368 6518 18380
rect 6549 18377 6561 18380
rect 6595 18377 6607 18411
rect 6549 18371 6607 18377
rect 7285 18411 7343 18417
rect 7285 18377 7297 18411
rect 7331 18408 7343 18411
rect 8386 18408 8392 18420
rect 7331 18380 8392 18408
rect 7331 18377 7343 18380
rect 7285 18371 7343 18377
rect 8386 18368 8392 18380
rect 8444 18368 8450 18420
rect 9950 18368 9956 18420
rect 10008 18408 10014 18420
rect 10413 18411 10471 18417
rect 10413 18408 10425 18411
rect 10008 18380 10425 18408
rect 10008 18368 10014 18380
rect 10413 18377 10425 18380
rect 10459 18377 10471 18411
rect 10413 18371 10471 18377
rect 12434 18368 12440 18420
rect 12492 18368 12498 18420
rect 15102 18368 15108 18420
rect 15160 18368 15166 18420
rect 15841 18411 15899 18417
rect 15841 18377 15853 18411
rect 15887 18408 15899 18411
rect 16206 18408 16212 18420
rect 15887 18380 16212 18408
rect 15887 18377 15899 18380
rect 15841 18371 15899 18377
rect 16206 18368 16212 18380
rect 16264 18368 16270 18420
rect 17034 18368 17040 18420
rect 17092 18408 17098 18420
rect 17773 18411 17831 18417
rect 17773 18408 17785 18411
rect 17092 18380 17785 18408
rect 17092 18368 17098 18380
rect 17773 18377 17785 18380
rect 17819 18377 17831 18411
rect 19702 18408 19708 18420
rect 17773 18371 17831 18377
rect 19260 18380 19708 18408
rect 5169 18343 5227 18349
rect 3660 18312 4016 18340
rect 3660 18300 3666 18312
rect 3988 18281 4016 18312
rect 5169 18309 5181 18343
rect 5215 18309 5227 18343
rect 7653 18343 7711 18349
rect 5169 18303 5227 18309
rect 6012 18312 7052 18340
rect 2674 18275 2732 18281
rect 2674 18272 2686 18275
rect 2424 18244 2686 18272
rect 2674 18241 2686 18244
rect 2720 18241 2732 18275
rect 2674 18235 2732 18241
rect 2869 18275 2927 18281
rect 2869 18241 2881 18275
rect 2915 18272 2927 18275
rect 3973 18275 4031 18281
rect 2915 18244 3648 18272
rect 2915 18241 2927 18244
rect 2869 18235 2927 18241
rect 1394 18164 1400 18216
rect 1452 18164 1458 18216
rect 1857 18207 1915 18213
rect 1857 18173 1869 18207
rect 1903 18204 1915 18207
rect 1964 18204 1992 18232
rect 1903 18176 1992 18204
rect 1903 18173 1915 18176
rect 1857 18167 1915 18173
rect 2222 18164 2228 18216
rect 2280 18204 2286 18216
rect 2280 18176 2443 18204
rect 2280 18164 2286 18176
rect 1412 18136 1440 18164
rect 2415 18136 2443 18176
rect 2884 18136 2912 18235
rect 3620 18216 3648 18244
rect 3973 18241 3985 18275
rect 4019 18241 4031 18275
rect 3973 18235 4031 18241
rect 2961 18207 3019 18213
rect 2961 18173 2973 18207
rect 3007 18204 3019 18207
rect 3421 18207 3479 18213
rect 3421 18204 3433 18207
rect 3007 18176 3433 18204
rect 3007 18173 3019 18176
rect 2961 18167 3019 18173
rect 3421 18173 3433 18176
rect 3467 18173 3479 18207
rect 3421 18167 3479 18173
rect 3602 18164 3608 18216
rect 3660 18164 3666 18216
rect 4893 18207 4951 18213
rect 4893 18173 4905 18207
rect 4939 18204 4951 18207
rect 5074 18204 5080 18216
rect 4939 18176 5080 18204
rect 4939 18173 4951 18176
rect 4893 18167 4951 18173
rect 5074 18164 5080 18176
rect 5132 18164 5138 18216
rect 5810 18164 5816 18216
rect 5868 18204 5874 18216
rect 6012 18204 6040 18312
rect 6089 18275 6147 18281
rect 6089 18241 6101 18275
rect 6135 18272 6147 18275
rect 6914 18272 6920 18284
rect 6135 18244 6920 18272
rect 6135 18241 6147 18244
rect 6089 18235 6147 18241
rect 6914 18232 6920 18244
rect 6972 18232 6978 18284
rect 7024 18272 7052 18312
rect 7653 18309 7665 18343
rect 7699 18340 7711 18343
rect 7834 18340 7840 18352
rect 7699 18312 7840 18340
rect 7699 18309 7711 18312
rect 7653 18303 7711 18309
rect 7834 18300 7840 18312
rect 7892 18300 7898 18352
rect 8938 18340 8944 18352
rect 8680 18312 8944 18340
rect 7024 18244 8524 18272
rect 8496 18216 8524 18244
rect 5868 18176 6040 18204
rect 5868 18164 5874 18176
rect 6362 18164 6368 18216
rect 6420 18204 6426 18216
rect 6457 18207 6515 18213
rect 6457 18204 6469 18207
rect 6420 18176 6469 18204
rect 6420 18164 6426 18176
rect 6457 18173 6469 18176
rect 6503 18173 6515 18207
rect 6457 18167 6515 18173
rect 6641 18207 6699 18213
rect 6641 18173 6653 18207
rect 6687 18204 6699 18207
rect 6730 18204 6736 18216
rect 6687 18176 6736 18204
rect 6687 18173 6699 18176
rect 6641 18167 6699 18173
rect 6730 18164 6736 18176
rect 6788 18164 6794 18216
rect 8478 18164 8484 18216
rect 8536 18164 8542 18216
rect 7285 18139 7343 18145
rect 7285 18136 7297 18139
rect 1412 18108 2360 18136
rect 2415 18108 2912 18136
rect 6932 18108 7297 18136
rect 2332 18080 2360 18108
rect 6932 18080 6960 18108
rect 7285 18105 7297 18108
rect 7331 18136 7343 18139
rect 8680 18136 8708 18312
rect 8938 18300 8944 18312
rect 8996 18300 9002 18352
rect 9030 18300 9036 18352
rect 9088 18340 9094 18352
rect 9582 18340 9588 18352
rect 9088 18312 9588 18340
rect 9088 18300 9094 18312
rect 9582 18300 9588 18312
rect 9640 18300 9646 18352
rect 8757 18275 8815 18281
rect 8757 18241 8769 18275
rect 8803 18272 8815 18275
rect 9674 18272 9680 18284
rect 8803 18244 9680 18272
rect 8803 18241 8815 18244
rect 8757 18235 8815 18241
rect 9674 18232 9680 18244
rect 9732 18232 9738 18284
rect 11054 18272 11060 18284
rect 9968 18244 11060 18272
rect 8938 18164 8944 18216
rect 8996 18164 9002 18216
rect 9030 18164 9036 18216
rect 9088 18164 9094 18216
rect 9401 18207 9459 18213
rect 9401 18173 9413 18207
rect 9447 18204 9459 18207
rect 9968 18204 9996 18244
rect 11054 18232 11060 18244
rect 11112 18232 11118 18284
rect 15010 18232 15016 18284
rect 15068 18272 15074 18284
rect 15068 18244 16160 18272
rect 15068 18232 15074 18244
rect 9447 18176 9996 18204
rect 9447 18173 9459 18176
rect 9401 18167 9459 18173
rect 10042 18164 10048 18216
rect 10100 18164 10106 18216
rect 11149 18207 11207 18213
rect 11149 18173 11161 18207
rect 11195 18204 11207 18207
rect 11606 18204 11612 18216
rect 11195 18176 11612 18204
rect 11195 18173 11207 18176
rect 11149 18167 11207 18173
rect 7331 18108 8708 18136
rect 7331 18105 7343 18108
rect 7285 18099 7343 18105
rect 8846 18096 8852 18148
rect 8904 18136 8910 18148
rect 11164 18136 11192 18167
rect 11606 18164 11612 18176
rect 11664 18164 11670 18216
rect 13262 18164 13268 18216
rect 13320 18204 13326 18216
rect 13725 18207 13783 18213
rect 13725 18204 13737 18207
rect 13320 18176 13737 18204
rect 13320 18164 13326 18176
rect 13725 18173 13737 18176
rect 13771 18204 13783 18207
rect 15470 18204 15476 18216
rect 13771 18176 15476 18204
rect 13771 18173 13783 18176
rect 13725 18167 13783 18173
rect 15470 18164 15476 18176
rect 15528 18164 15534 18216
rect 15565 18207 15623 18213
rect 15565 18173 15577 18207
rect 15611 18204 15623 18207
rect 15657 18207 15715 18213
rect 15657 18204 15669 18207
rect 15611 18176 15669 18204
rect 15611 18173 15623 18176
rect 15565 18167 15623 18173
rect 15657 18173 15669 18176
rect 15703 18173 15715 18207
rect 15657 18167 15715 18173
rect 8904 18108 11192 18136
rect 13992 18139 14050 18145
rect 8904 18096 8910 18108
rect 13992 18105 14004 18139
rect 14038 18136 14050 18139
rect 14182 18136 14188 18148
rect 14038 18108 14188 18136
rect 14038 18105 14050 18108
rect 13992 18099 14050 18105
rect 14182 18096 14188 18108
rect 14240 18096 14246 18148
rect 15102 18096 15108 18148
rect 15160 18096 15166 18148
rect 15194 18096 15200 18148
rect 15252 18096 15258 18148
rect 15381 18139 15439 18145
rect 15381 18105 15393 18139
rect 15427 18105 15439 18139
rect 16132 18136 16160 18244
rect 16224 18204 16252 18368
rect 17497 18275 17555 18281
rect 17497 18241 17509 18275
rect 17543 18272 17555 18275
rect 17862 18272 17868 18284
rect 17543 18244 17868 18272
rect 17543 18241 17555 18244
rect 17497 18235 17555 18241
rect 17862 18232 17868 18244
rect 17920 18272 17926 18284
rect 19260 18281 19288 18380
rect 19702 18368 19708 18380
rect 19760 18368 19766 18420
rect 19797 18411 19855 18417
rect 19797 18377 19809 18411
rect 19843 18408 19855 18411
rect 20162 18408 20168 18420
rect 19843 18380 20168 18408
rect 19843 18377 19855 18380
rect 19797 18371 19855 18377
rect 20162 18368 20168 18380
rect 20220 18368 20226 18420
rect 20990 18408 20996 18420
rect 20272 18380 20996 18408
rect 20272 18340 20300 18380
rect 20990 18368 20996 18380
rect 21048 18368 21054 18420
rect 21082 18368 21088 18420
rect 21140 18408 21146 18420
rect 21729 18411 21787 18417
rect 21729 18408 21741 18411
rect 21140 18380 21741 18408
rect 21140 18368 21146 18380
rect 21729 18377 21741 18380
rect 21775 18377 21787 18411
rect 21729 18371 21787 18377
rect 19352 18312 20300 18340
rect 18417 18275 18475 18281
rect 18417 18272 18429 18275
rect 17920 18244 18429 18272
rect 17920 18232 17926 18244
rect 18417 18241 18429 18244
rect 18463 18272 18475 18275
rect 19245 18275 19303 18281
rect 19245 18272 19257 18275
rect 18463 18244 19257 18272
rect 18463 18241 18475 18244
rect 18417 18235 18475 18241
rect 19245 18241 19257 18244
rect 19291 18241 19303 18275
rect 19245 18235 19303 18241
rect 16761 18207 16819 18213
rect 16761 18204 16773 18207
rect 16224 18176 16773 18204
rect 16761 18173 16773 18176
rect 16807 18204 16819 18207
rect 16850 18204 16856 18216
rect 16807 18176 16856 18204
rect 16807 18173 16819 18176
rect 16761 18167 16819 18173
rect 16850 18164 16856 18176
rect 16908 18164 16914 18216
rect 17221 18207 17279 18213
rect 17221 18173 17233 18207
rect 17267 18173 17279 18207
rect 17221 18167 17279 18173
rect 18233 18207 18291 18213
rect 18233 18173 18245 18207
rect 18279 18204 18291 18207
rect 18506 18204 18512 18216
rect 18279 18176 18512 18204
rect 18279 18173 18291 18176
rect 18233 18167 18291 18173
rect 17236 18136 17264 18167
rect 18506 18164 18512 18176
rect 18564 18164 18570 18216
rect 19352 18145 19380 18312
rect 19426 18232 19432 18284
rect 19484 18272 19490 18284
rect 20349 18275 20407 18281
rect 20349 18272 20361 18275
rect 19484 18244 20361 18272
rect 19484 18232 19490 18244
rect 20349 18241 20361 18244
rect 20395 18241 20407 18275
rect 20349 18235 20407 18241
rect 19886 18164 19892 18216
rect 19944 18164 19950 18216
rect 20438 18164 20444 18216
rect 20496 18204 20502 18216
rect 20605 18207 20663 18213
rect 20605 18204 20617 18207
rect 20496 18176 20617 18204
rect 20496 18164 20502 18176
rect 20605 18173 20617 18176
rect 20651 18173 20663 18207
rect 20605 18167 20663 18173
rect 16132 18108 17264 18136
rect 19337 18139 19395 18145
rect 15381 18099 15439 18105
rect 1670 18028 1676 18080
rect 1728 18028 1734 18080
rect 1762 18028 1768 18080
rect 1820 18028 1826 18080
rect 2314 18028 2320 18080
rect 2372 18028 2378 18080
rect 6914 18028 6920 18080
rect 6972 18028 6978 18080
rect 7006 18028 7012 18080
rect 7064 18068 7070 18080
rect 7101 18071 7159 18077
rect 7101 18068 7113 18071
rect 7064 18040 7113 18068
rect 7064 18028 7070 18040
rect 7101 18037 7113 18040
rect 7147 18037 7159 18071
rect 7101 18031 7159 18037
rect 8662 18028 8668 18080
rect 8720 18068 8726 18080
rect 9214 18068 9220 18080
rect 8720 18040 9220 18068
rect 8720 18028 8726 18040
rect 9214 18028 9220 18040
rect 9272 18028 9278 18080
rect 9490 18028 9496 18080
rect 9548 18028 9554 18080
rect 15120 18068 15148 18096
rect 15396 18068 15424 18099
rect 16776 18080 16804 18108
rect 19337 18105 19349 18139
rect 19383 18105 19395 18139
rect 19337 18099 19395 18105
rect 19429 18139 19487 18145
rect 19429 18105 19441 18139
rect 19475 18136 19487 18139
rect 19904 18136 19932 18164
rect 19475 18108 19932 18136
rect 21744 18136 21772 18371
rect 22278 18368 22284 18420
rect 22336 18368 22342 18420
rect 22462 18368 22468 18420
rect 22520 18408 22526 18420
rect 22557 18411 22615 18417
rect 22557 18408 22569 18411
rect 22520 18380 22569 18408
rect 22520 18368 22526 18380
rect 22557 18377 22569 18380
rect 22603 18377 22615 18411
rect 22557 18371 22615 18377
rect 22738 18368 22744 18420
rect 22796 18368 22802 18420
rect 22830 18368 22836 18420
rect 22888 18408 22894 18420
rect 23293 18411 23351 18417
rect 23293 18408 23305 18411
rect 22888 18380 23305 18408
rect 22888 18368 22894 18380
rect 23293 18377 23305 18380
rect 23339 18377 23351 18411
rect 23293 18371 23351 18377
rect 23566 18368 23572 18420
rect 23624 18408 23630 18420
rect 23661 18411 23719 18417
rect 23661 18408 23673 18411
rect 23624 18380 23673 18408
rect 23624 18368 23630 18380
rect 23661 18377 23673 18380
rect 23707 18408 23719 18411
rect 24118 18408 24124 18420
rect 23707 18380 24124 18408
rect 23707 18377 23719 18380
rect 23661 18371 23719 18377
rect 24118 18368 24124 18380
rect 24176 18368 24182 18420
rect 24213 18411 24271 18417
rect 24213 18377 24225 18411
rect 24259 18408 24271 18411
rect 25406 18408 25412 18420
rect 24259 18380 25412 18408
rect 24259 18377 24271 18380
rect 24213 18371 24271 18377
rect 25406 18368 25412 18380
rect 25464 18368 25470 18420
rect 22296 18340 22324 18368
rect 22649 18343 22707 18349
rect 22649 18340 22661 18343
rect 22296 18312 22661 18340
rect 22649 18309 22661 18312
rect 22695 18309 22707 18343
rect 22756 18340 22784 18368
rect 23109 18343 23167 18349
rect 23109 18340 23121 18343
rect 22756 18312 23121 18340
rect 22649 18303 22707 18309
rect 23109 18309 23121 18312
rect 23155 18309 23167 18343
rect 23109 18303 23167 18309
rect 24302 18300 24308 18352
rect 24360 18300 24366 18352
rect 24486 18300 24492 18352
rect 24544 18300 24550 18352
rect 23385 18275 23443 18281
rect 23385 18272 23397 18275
rect 22296 18244 22968 18272
rect 21910 18164 21916 18216
rect 21968 18204 21974 18216
rect 22296 18213 22324 18244
rect 22940 18213 22968 18244
rect 23124 18244 23397 18272
rect 23124 18216 23152 18244
rect 23385 18241 23397 18244
rect 23431 18241 23443 18275
rect 24320 18272 24348 18300
rect 23385 18235 23443 18241
rect 24044 18244 24348 18272
rect 22005 18207 22063 18213
rect 22005 18204 22017 18207
rect 21968 18176 22017 18204
rect 21968 18164 21974 18176
rect 22005 18173 22017 18176
rect 22051 18173 22063 18207
rect 22005 18167 22063 18173
rect 22281 18207 22339 18213
rect 22281 18173 22293 18207
rect 22327 18173 22339 18207
rect 22281 18167 22339 18173
rect 22373 18207 22431 18213
rect 22373 18173 22385 18207
rect 22419 18204 22431 18207
rect 22833 18207 22891 18213
rect 22833 18204 22845 18207
rect 22419 18176 22845 18204
rect 22419 18173 22431 18176
rect 22373 18167 22431 18173
rect 22833 18173 22845 18176
rect 22879 18173 22891 18207
rect 22833 18167 22891 18173
rect 22925 18207 22983 18213
rect 22925 18173 22937 18207
rect 22971 18173 22983 18207
rect 22925 18167 22983 18173
rect 21744 18108 22140 18136
rect 19475 18105 19487 18108
rect 19429 18099 19487 18105
rect 15120 18040 15424 18068
rect 16758 18028 16764 18080
rect 16816 18028 16822 18080
rect 18138 18028 18144 18080
rect 18196 18028 18202 18080
rect 18690 18028 18696 18080
rect 18748 18068 18754 18080
rect 21174 18068 21180 18080
rect 18748 18040 21180 18068
rect 18748 18028 18754 18040
rect 21174 18028 21180 18040
rect 21232 18028 21238 18080
rect 22112 18068 22140 18108
rect 22186 18096 22192 18148
rect 22244 18096 22250 18148
rect 22388 18068 22416 18167
rect 22940 18136 22968 18167
rect 23106 18164 23112 18216
rect 23164 18164 23170 18216
rect 23198 18164 23204 18216
rect 23256 18164 23262 18216
rect 23290 18164 23296 18216
rect 23348 18204 23354 18216
rect 24044 18213 24072 18244
rect 23937 18207 23995 18213
rect 23937 18204 23949 18207
rect 23348 18176 23949 18204
rect 23348 18164 23354 18176
rect 23937 18173 23949 18176
rect 23983 18173 23995 18207
rect 23937 18167 23995 18173
rect 24029 18207 24087 18213
rect 24029 18173 24041 18207
rect 24075 18173 24087 18207
rect 24029 18167 24087 18173
rect 24118 18164 24124 18216
rect 24176 18164 24182 18216
rect 24305 18207 24363 18213
rect 24305 18173 24317 18207
rect 24351 18173 24363 18207
rect 24504 18204 24532 18300
rect 24581 18207 24639 18213
rect 24581 18204 24593 18207
rect 24504 18176 24593 18204
rect 24305 18167 24363 18173
rect 24581 18173 24593 18176
rect 24627 18173 24639 18207
rect 24581 18167 24639 18173
rect 25685 18207 25743 18213
rect 25685 18173 25697 18207
rect 25731 18204 25743 18207
rect 25774 18204 25780 18216
rect 25731 18176 25780 18204
rect 25731 18173 25743 18176
rect 25685 18167 25743 18173
rect 24320 18136 24348 18167
rect 25774 18164 25780 18176
rect 25832 18164 25838 18216
rect 25958 18145 25964 18148
rect 24489 18139 24547 18145
rect 24489 18136 24501 18139
rect 22940 18108 24501 18136
rect 24489 18105 24501 18108
rect 24535 18105 24547 18139
rect 24489 18099 24547 18105
rect 25952 18099 25964 18145
rect 25958 18096 25964 18099
rect 26016 18096 26022 18148
rect 22112 18040 22416 18068
rect 25038 18028 25044 18080
rect 25096 18068 25102 18080
rect 27065 18071 27123 18077
rect 27065 18068 27077 18071
rect 25096 18040 27077 18068
rect 25096 18028 25102 18040
rect 27065 18037 27077 18040
rect 27111 18037 27123 18071
rect 27065 18031 27123 18037
rect 552 17978 27576 18000
rect 552 17926 7114 17978
rect 7166 17926 7178 17978
rect 7230 17926 7242 17978
rect 7294 17926 7306 17978
rect 7358 17926 7370 17978
rect 7422 17926 13830 17978
rect 13882 17926 13894 17978
rect 13946 17926 13958 17978
rect 14010 17926 14022 17978
rect 14074 17926 14086 17978
rect 14138 17926 20546 17978
rect 20598 17926 20610 17978
rect 20662 17926 20674 17978
rect 20726 17926 20738 17978
rect 20790 17926 20802 17978
rect 20854 17926 27262 17978
rect 27314 17926 27326 17978
rect 27378 17926 27390 17978
rect 27442 17926 27454 17978
rect 27506 17926 27518 17978
rect 27570 17926 27576 17978
rect 552 17904 27576 17926
rect 1762 17824 1768 17876
rect 1820 17864 1826 17876
rect 2317 17867 2375 17873
rect 2317 17864 2329 17867
rect 1820 17836 2329 17864
rect 1820 17824 1826 17836
rect 2317 17833 2329 17836
rect 2363 17833 2375 17867
rect 2317 17827 2375 17833
rect 3436 17836 4016 17864
rect 3436 17808 3464 17836
rect 3418 17756 3424 17808
rect 3476 17756 3482 17808
rect 3510 17756 3516 17808
rect 3568 17796 3574 17808
rect 3881 17799 3939 17805
rect 3881 17796 3893 17799
rect 3568 17768 3893 17796
rect 3568 17756 3574 17768
rect 3881 17765 3893 17768
rect 3927 17765 3939 17799
rect 3881 17759 3939 17765
rect 842 17688 848 17740
rect 900 17688 906 17740
rect 1112 17731 1170 17737
rect 1112 17697 1124 17731
rect 1158 17728 1170 17731
rect 1394 17728 1400 17740
rect 1158 17700 1400 17728
rect 1158 17697 1170 17700
rect 1112 17691 1170 17697
rect 1394 17688 1400 17700
rect 1452 17688 1458 17740
rect 2961 17731 3019 17737
rect 2961 17697 2973 17731
rect 3007 17728 3019 17731
rect 3007 17700 3556 17728
rect 3007 17697 3019 17700
rect 2961 17691 3019 17697
rect 2225 17595 2283 17601
rect 2225 17561 2237 17595
rect 2271 17592 2283 17595
rect 2774 17592 2780 17604
rect 2271 17564 2780 17592
rect 2271 17561 2283 17564
rect 2225 17555 2283 17561
rect 2774 17552 2780 17564
rect 2832 17592 2838 17604
rect 2976 17592 3004 17691
rect 3329 17663 3387 17669
rect 3329 17629 3341 17663
rect 3375 17629 3387 17663
rect 3329 17623 3387 17629
rect 2832 17564 3004 17592
rect 2832 17552 2838 17564
rect 3344 17536 3372 17623
rect 3418 17620 3424 17672
rect 3476 17620 3482 17672
rect 3528 17669 3556 17700
rect 3602 17688 3608 17740
rect 3660 17688 3666 17740
rect 3988 17728 4016 17836
rect 4614 17824 4620 17876
rect 4672 17864 4678 17876
rect 4890 17864 4896 17876
rect 4672 17836 4896 17864
rect 4672 17824 4678 17836
rect 4890 17824 4896 17836
rect 4948 17864 4954 17876
rect 5445 17867 5503 17873
rect 5445 17864 5457 17867
rect 4948 17836 5457 17864
rect 4948 17824 4954 17836
rect 5445 17833 5457 17836
rect 5491 17833 5503 17867
rect 5445 17827 5503 17833
rect 7745 17867 7803 17873
rect 7745 17833 7757 17867
rect 7791 17864 7803 17867
rect 8294 17864 8300 17876
rect 7791 17836 8300 17864
rect 7791 17833 7803 17836
rect 7745 17827 7803 17833
rect 8294 17824 8300 17836
rect 8352 17824 8358 17876
rect 8481 17867 8539 17873
rect 8481 17833 8493 17867
rect 8527 17864 8539 17867
rect 8662 17864 8668 17876
rect 8527 17836 8668 17864
rect 8527 17833 8539 17836
rect 8481 17827 8539 17833
rect 8662 17824 8668 17836
rect 8720 17824 8726 17876
rect 8849 17867 8907 17873
rect 8849 17833 8861 17867
rect 8895 17864 8907 17867
rect 9122 17864 9128 17876
rect 8895 17836 9128 17864
rect 8895 17833 8907 17836
rect 8849 17827 8907 17833
rect 9122 17824 9128 17836
rect 9180 17824 9186 17876
rect 9490 17824 9496 17876
rect 9548 17824 9554 17876
rect 9674 17824 9680 17876
rect 9732 17824 9738 17876
rect 11054 17824 11060 17876
rect 11112 17864 11118 17876
rect 11885 17867 11943 17873
rect 11885 17864 11897 17867
rect 11112 17836 11897 17864
rect 11112 17824 11118 17836
rect 11885 17833 11897 17836
rect 11931 17833 11943 17867
rect 11885 17827 11943 17833
rect 13170 17824 13176 17876
rect 13228 17864 13234 17876
rect 14366 17864 14372 17876
rect 13228 17836 13676 17864
rect 13228 17824 13234 17836
rect 5074 17756 5080 17808
rect 5132 17796 5138 17808
rect 9508 17796 9536 17824
rect 5132 17768 8248 17796
rect 5132 17756 5138 17768
rect 4157 17731 4215 17737
rect 4157 17728 4169 17731
rect 3988 17700 4169 17728
rect 4157 17697 4169 17700
rect 4203 17697 4215 17731
rect 4157 17691 4215 17697
rect 4614 17688 4620 17740
rect 4672 17688 4678 17740
rect 4982 17688 4988 17740
rect 5040 17688 5046 17740
rect 5092 17728 5120 17756
rect 5169 17731 5227 17737
rect 5169 17728 5181 17731
rect 5092 17700 5181 17728
rect 5169 17697 5181 17700
rect 5215 17697 5227 17731
rect 5169 17691 5227 17697
rect 5353 17731 5411 17737
rect 5353 17697 5365 17731
rect 5399 17728 5411 17731
rect 5629 17731 5687 17737
rect 5629 17728 5641 17731
rect 5399 17700 5641 17728
rect 5399 17697 5411 17700
rect 5353 17691 5411 17697
rect 5629 17697 5641 17700
rect 5675 17697 5687 17731
rect 5629 17691 5687 17697
rect 6270 17688 6276 17740
rect 6328 17728 6334 17740
rect 6638 17737 6644 17740
rect 6365 17731 6423 17737
rect 6365 17728 6377 17731
rect 6328 17700 6377 17728
rect 6328 17688 6334 17700
rect 6365 17697 6377 17700
rect 6411 17697 6423 17731
rect 6365 17691 6423 17697
rect 6632 17691 6644 17737
rect 6638 17688 6644 17691
rect 6696 17688 6702 17740
rect 3513 17663 3571 17669
rect 3513 17629 3525 17663
rect 3559 17660 3571 17663
rect 3973 17663 4031 17669
rect 3973 17660 3985 17663
rect 3559 17632 3985 17660
rect 3559 17629 3571 17632
rect 3513 17623 3571 17629
rect 3973 17629 3985 17632
rect 4019 17629 4031 17663
rect 3973 17623 4031 17629
rect 3789 17595 3847 17601
rect 3789 17561 3801 17595
rect 3835 17592 3847 17595
rect 4154 17592 4160 17604
rect 3835 17564 4160 17592
rect 3835 17561 3847 17564
rect 3789 17555 3847 17561
rect 4154 17552 4160 17564
rect 4212 17552 4218 17604
rect 4341 17595 4399 17601
rect 4341 17561 4353 17595
rect 4387 17592 4399 17595
rect 5350 17592 5356 17604
rect 4387 17564 5356 17592
rect 4387 17561 4399 17564
rect 4341 17555 4399 17561
rect 5350 17552 5356 17564
rect 5408 17552 5414 17604
rect 8220 17592 8248 17768
rect 8312 17768 9536 17796
rect 8312 17737 8340 17768
rect 8297 17731 8355 17737
rect 8297 17697 8309 17731
rect 8343 17697 8355 17731
rect 8297 17691 8355 17697
rect 8389 17731 8447 17737
rect 8389 17697 8401 17731
rect 8435 17728 8447 17731
rect 8478 17728 8484 17740
rect 8435 17700 8484 17728
rect 8435 17697 8447 17700
rect 8389 17691 8447 17697
rect 8478 17688 8484 17700
rect 8536 17688 8542 17740
rect 8665 17731 8723 17737
rect 8665 17697 8677 17731
rect 8711 17728 8723 17731
rect 8754 17728 8760 17740
rect 8711 17700 8760 17728
rect 8711 17697 8723 17700
rect 8665 17691 8723 17697
rect 8754 17688 8760 17700
rect 8812 17688 8818 17740
rect 8938 17688 8944 17740
rect 8996 17688 9002 17740
rect 9122 17688 9128 17740
rect 9180 17688 9186 17740
rect 9214 17688 9220 17740
rect 9272 17688 9278 17740
rect 9306 17688 9312 17740
rect 9364 17728 9370 17740
rect 9692 17737 9720 17824
rect 13648 17805 13676 17836
rect 14200 17836 14372 17864
rect 11793 17799 11851 17805
rect 9784 17768 9996 17796
rect 9784 17740 9812 17768
rect 9493 17731 9551 17737
rect 9493 17728 9505 17731
rect 9364 17700 9505 17728
rect 9364 17688 9370 17700
rect 9493 17697 9505 17700
rect 9539 17697 9551 17731
rect 9493 17691 9551 17697
rect 9677 17731 9735 17737
rect 9677 17697 9689 17731
rect 9723 17697 9735 17731
rect 9677 17691 9735 17697
rect 9766 17688 9772 17740
rect 9824 17688 9830 17740
rect 9968 17737 9996 17768
rect 10244 17768 10824 17796
rect 10244 17737 10272 17768
rect 9861 17731 9919 17737
rect 9861 17697 9873 17731
rect 9907 17697 9919 17731
rect 9861 17691 9919 17697
rect 9953 17731 10011 17737
rect 9953 17697 9965 17731
rect 9999 17697 10011 17731
rect 9953 17691 10011 17697
rect 10229 17731 10287 17737
rect 10229 17697 10241 17731
rect 10275 17697 10287 17731
rect 10229 17691 10287 17697
rect 8956 17660 8984 17688
rect 9876 17660 9904 17691
rect 10318 17688 10324 17740
rect 10376 17688 10382 17740
rect 8956 17632 9904 17660
rect 10045 17663 10103 17669
rect 10045 17629 10057 17663
rect 10091 17660 10103 17663
rect 10134 17660 10140 17672
rect 10091 17632 10140 17660
rect 10091 17629 10103 17632
rect 10045 17623 10103 17629
rect 10134 17620 10140 17632
rect 10192 17620 10198 17672
rect 8220 17564 9168 17592
rect 9140 17536 9168 17564
rect 9214 17552 9220 17604
rect 9272 17592 9278 17604
rect 10336 17592 10364 17688
rect 9272 17564 10364 17592
rect 10796 17592 10824 17768
rect 11793 17765 11805 17799
rect 11839 17796 11851 17799
rect 13633 17799 13691 17805
rect 11839 17768 13400 17796
rect 11839 17765 11851 17768
rect 11793 17759 11851 17765
rect 10870 17688 10876 17740
rect 10928 17728 10934 17740
rect 10928 17700 11284 17728
rect 10928 17688 10934 17700
rect 11149 17663 11207 17669
rect 11149 17629 11161 17663
rect 11195 17629 11207 17663
rect 11149 17623 11207 17629
rect 10870 17592 10876 17604
rect 10796 17564 10876 17592
rect 9272 17552 9278 17564
rect 10870 17552 10876 17564
rect 10928 17552 10934 17604
rect 11164 17536 11192 17623
rect 3326 17484 3332 17536
rect 3384 17524 3390 17536
rect 3881 17527 3939 17533
rect 3881 17524 3893 17527
rect 3384 17496 3893 17524
rect 3384 17484 3390 17496
rect 3881 17493 3893 17496
rect 3927 17493 3939 17527
rect 3881 17487 3939 17493
rect 4430 17484 4436 17536
rect 4488 17484 4494 17536
rect 7926 17484 7932 17536
rect 7984 17524 7990 17536
rect 8205 17527 8263 17533
rect 8205 17524 8217 17527
rect 7984 17496 8217 17524
rect 7984 17484 7990 17496
rect 8205 17493 8217 17496
rect 8251 17493 8263 17527
rect 8205 17487 8263 17493
rect 9122 17484 9128 17536
rect 9180 17484 9186 17536
rect 9401 17527 9459 17533
rect 9401 17493 9413 17527
rect 9447 17524 9459 17527
rect 10226 17524 10232 17536
rect 9447 17496 10232 17524
rect 9447 17493 9459 17496
rect 9401 17487 9459 17493
rect 10226 17484 10232 17496
rect 10284 17484 10290 17536
rect 10318 17484 10324 17536
rect 10376 17524 10382 17536
rect 10413 17527 10471 17533
rect 10413 17524 10425 17527
rect 10376 17496 10425 17524
rect 10376 17484 10382 17496
rect 10413 17493 10425 17496
rect 10459 17493 10471 17527
rect 10413 17487 10471 17493
rect 11146 17484 11152 17536
rect 11204 17484 11210 17536
rect 11256 17524 11284 17700
rect 12618 17688 12624 17740
rect 12676 17728 12682 17740
rect 12998 17731 13056 17737
rect 12998 17728 13010 17731
rect 12676 17700 13010 17728
rect 12676 17688 12682 17700
rect 12998 17697 13010 17700
rect 13044 17697 13056 17731
rect 12998 17691 13056 17697
rect 13262 17688 13268 17740
rect 13320 17688 13326 17740
rect 13372 17737 13400 17768
rect 13633 17765 13645 17799
rect 13679 17796 13691 17799
rect 13998 17796 14004 17808
rect 13679 17768 14004 17796
rect 13679 17765 13691 17768
rect 13633 17759 13691 17765
rect 13998 17756 14004 17768
rect 14056 17756 14062 17808
rect 13357 17731 13415 17737
rect 13357 17697 13369 17731
rect 13403 17697 13415 17731
rect 13357 17691 13415 17697
rect 13446 17688 13452 17740
rect 13504 17728 13510 17740
rect 13541 17731 13599 17737
rect 13541 17728 13553 17731
rect 13504 17700 13553 17728
rect 13504 17688 13510 17700
rect 13541 17697 13553 17700
rect 13587 17697 13599 17731
rect 13541 17691 13599 17697
rect 13722 17688 13728 17740
rect 13780 17688 13786 17740
rect 13814 17688 13820 17740
rect 13872 17728 13878 17740
rect 14200 17737 14228 17836
rect 14366 17824 14372 17836
rect 14424 17824 14430 17876
rect 15102 17824 15108 17876
rect 15160 17824 15166 17876
rect 15286 17824 15292 17876
rect 15344 17864 15350 17876
rect 15749 17867 15807 17873
rect 15749 17864 15761 17867
rect 15344 17836 15761 17864
rect 15344 17824 15350 17836
rect 15749 17833 15761 17836
rect 15795 17833 15807 17867
rect 15749 17827 15807 17833
rect 17589 17867 17647 17873
rect 17589 17833 17601 17867
rect 17635 17864 17647 17867
rect 17678 17864 17684 17876
rect 17635 17836 17684 17864
rect 17635 17833 17647 17836
rect 17589 17827 17647 17833
rect 15120 17796 15148 17824
rect 14476 17768 15332 17796
rect 14476 17737 14504 17768
rect 14185 17731 14243 17737
rect 14185 17728 14197 17731
rect 13872 17700 14197 17728
rect 13872 17688 13878 17700
rect 14185 17697 14197 17700
rect 14231 17697 14243 17731
rect 14185 17691 14243 17697
rect 14369 17731 14427 17737
rect 14369 17697 14381 17731
rect 14415 17697 14427 17731
rect 14369 17691 14427 17697
rect 14461 17731 14519 17737
rect 14461 17697 14473 17731
rect 14507 17697 14519 17731
rect 14461 17691 14519 17697
rect 14645 17731 14703 17737
rect 14645 17697 14657 17731
rect 14691 17728 14703 17731
rect 15194 17728 15200 17740
rect 14691 17700 15200 17728
rect 14691 17697 14703 17700
rect 14645 17691 14703 17697
rect 13630 17620 13636 17672
rect 13688 17660 13694 17672
rect 14001 17663 14059 17669
rect 14001 17660 14013 17663
rect 13688 17632 14013 17660
rect 13688 17620 13694 17632
rect 14001 17629 14013 17632
rect 14047 17629 14059 17663
rect 14001 17623 14059 17629
rect 14384 17592 14412 17691
rect 15194 17688 15200 17700
rect 15252 17688 15258 17740
rect 15304 17737 15332 17768
rect 15289 17731 15347 17737
rect 15289 17697 15301 17731
rect 15335 17728 15347 17731
rect 15381 17731 15439 17737
rect 15381 17728 15393 17731
rect 15335 17700 15393 17728
rect 15335 17697 15347 17700
rect 15289 17691 15347 17697
rect 15381 17697 15393 17700
rect 15427 17697 15439 17731
rect 15764 17728 15792 17827
rect 17678 17824 17684 17836
rect 17736 17824 17742 17876
rect 18138 17824 18144 17876
rect 18196 17864 18202 17876
rect 18325 17867 18383 17873
rect 18325 17864 18337 17867
rect 18196 17836 18337 17864
rect 18196 17824 18202 17836
rect 18325 17833 18337 17836
rect 18371 17833 18383 17867
rect 18325 17827 18383 17833
rect 23109 17867 23167 17873
rect 23109 17833 23121 17867
rect 23155 17864 23167 17867
rect 23198 17864 23204 17876
rect 23155 17836 23204 17864
rect 23155 17833 23167 17836
rect 23109 17827 23167 17833
rect 23198 17824 23204 17836
rect 23256 17824 23262 17876
rect 25425 17867 25483 17873
rect 25425 17864 25437 17867
rect 24228 17836 25176 17864
rect 16761 17799 16819 17805
rect 16761 17765 16773 17799
rect 16807 17796 16819 17799
rect 18046 17796 18052 17808
rect 16807 17768 18052 17796
rect 16807 17765 16819 17768
rect 16761 17759 16819 17765
rect 18046 17756 18052 17768
rect 18104 17756 18110 17808
rect 20070 17796 20076 17808
rect 18524 17768 20076 17796
rect 16393 17731 16451 17737
rect 16393 17728 16405 17731
rect 15764 17700 16405 17728
rect 15381 17691 15439 17697
rect 16393 17697 16405 17700
rect 16439 17697 16451 17731
rect 16393 17691 16451 17697
rect 16850 17688 16856 17740
rect 16908 17688 16914 17740
rect 17129 17731 17187 17737
rect 17129 17697 17141 17731
rect 17175 17728 17187 17731
rect 17586 17728 17592 17740
rect 17175 17700 17592 17728
rect 17175 17697 17187 17700
rect 17129 17691 17187 17697
rect 14553 17595 14611 17601
rect 14553 17592 14565 17595
rect 13756 17564 14565 17592
rect 13756 17524 13784 17564
rect 14553 17561 14565 17564
rect 14599 17561 14611 17595
rect 14553 17555 14611 17561
rect 11256 17496 13784 17524
rect 13906 17484 13912 17536
rect 13964 17484 13970 17536
rect 14734 17484 14740 17536
rect 14792 17524 14798 17536
rect 15212 17533 15240 17688
rect 16574 17620 16580 17672
rect 16632 17660 16638 17672
rect 17144 17660 17172 17691
rect 17586 17688 17592 17700
rect 17644 17688 17650 17740
rect 17770 17688 17776 17740
rect 17828 17688 17834 17740
rect 18524 17737 18552 17768
rect 20070 17756 20076 17768
rect 20128 17756 20134 17808
rect 23566 17756 23572 17808
rect 23624 17796 23630 17808
rect 24228 17805 24256 17836
rect 24213 17799 24271 17805
rect 24213 17796 24225 17799
rect 23624 17768 24225 17796
rect 23624 17756 23630 17768
rect 24213 17765 24225 17768
rect 24259 17765 24271 17799
rect 24213 17759 24271 17765
rect 24302 17756 24308 17808
rect 24360 17796 24366 17808
rect 24413 17799 24471 17805
rect 24413 17796 24425 17799
rect 24360 17768 24425 17796
rect 24360 17756 24366 17768
rect 24413 17765 24425 17768
rect 24459 17765 24471 17799
rect 24413 17759 24471 17765
rect 24765 17799 24823 17805
rect 24765 17765 24777 17799
rect 24811 17796 24823 17799
rect 24854 17796 24860 17808
rect 24811 17768 24860 17796
rect 24811 17765 24823 17768
rect 24765 17759 24823 17765
rect 18509 17731 18567 17737
rect 18509 17728 18521 17731
rect 17880 17700 18521 17728
rect 16632 17632 17172 17660
rect 16632 17620 16638 17632
rect 15286 17552 15292 17604
rect 15344 17592 15350 17604
rect 17880 17592 17908 17700
rect 18509 17697 18521 17700
rect 18555 17697 18567 17731
rect 18509 17691 18567 17697
rect 18690 17688 18696 17740
rect 18748 17688 18754 17740
rect 19058 17688 19064 17740
rect 19116 17688 19122 17740
rect 19797 17731 19855 17737
rect 19797 17697 19809 17731
rect 19843 17728 19855 17731
rect 20438 17728 20444 17740
rect 19843 17700 20444 17728
rect 19843 17697 19855 17700
rect 19797 17691 19855 17697
rect 17954 17620 17960 17672
rect 18012 17660 18018 17672
rect 18322 17660 18328 17672
rect 18012 17632 18328 17660
rect 18012 17620 18018 17632
rect 18322 17620 18328 17632
rect 18380 17660 18386 17672
rect 19812 17660 19840 17691
rect 20438 17688 20444 17700
rect 20496 17728 20502 17740
rect 20898 17728 20904 17740
rect 20496 17700 20904 17728
rect 20496 17688 20502 17700
rect 20898 17688 20904 17700
rect 20956 17728 20962 17740
rect 21453 17731 21511 17737
rect 21453 17728 21465 17731
rect 20956 17700 21465 17728
rect 20956 17688 20962 17700
rect 21453 17697 21465 17700
rect 21499 17697 21511 17731
rect 22373 17731 22431 17737
rect 22373 17728 22385 17731
rect 21453 17691 21511 17697
rect 22066 17700 22385 17728
rect 18380 17632 19840 17660
rect 19981 17663 20039 17669
rect 18380 17620 18386 17632
rect 19981 17629 19993 17663
rect 20027 17629 20039 17663
rect 19981 17623 20039 17629
rect 21269 17663 21327 17669
rect 21269 17629 21281 17663
rect 21315 17660 21327 17663
rect 21818 17660 21824 17672
rect 21315 17632 21824 17660
rect 21315 17629 21327 17632
rect 21269 17623 21327 17629
rect 15344 17564 17908 17592
rect 15344 17552 15350 17564
rect 18046 17552 18052 17604
rect 18104 17592 18110 17604
rect 19886 17592 19892 17604
rect 18104 17564 19892 17592
rect 18104 17552 18110 17564
rect 19886 17552 19892 17564
rect 19944 17552 19950 17604
rect 19996 17592 20024 17623
rect 21818 17620 21824 17632
rect 21876 17660 21882 17672
rect 22066 17660 22094 17700
rect 22373 17697 22385 17700
rect 22419 17697 22431 17731
rect 22373 17691 22431 17697
rect 22462 17688 22468 17740
rect 22520 17688 22526 17740
rect 22738 17688 22744 17740
rect 22796 17688 22802 17740
rect 23201 17731 23259 17737
rect 23201 17697 23213 17731
rect 23247 17728 23259 17731
rect 23937 17731 23995 17737
rect 23937 17728 23949 17731
rect 23247 17700 23949 17728
rect 23247 17697 23259 17700
rect 23201 17691 23259 17697
rect 23937 17697 23949 17700
rect 23983 17697 23995 17731
rect 23937 17691 23995 17697
rect 24121 17731 24179 17737
rect 24121 17697 24133 17731
rect 24167 17728 24179 17731
rect 24670 17728 24676 17740
rect 24167 17700 24676 17728
rect 24167 17697 24179 17700
rect 24121 17691 24179 17697
rect 21876 17632 22094 17660
rect 23952 17660 23980 17691
rect 24670 17688 24676 17700
rect 24728 17728 24734 17740
rect 24780 17728 24808 17759
rect 24854 17756 24860 17768
rect 24912 17756 24918 17808
rect 24949 17799 25007 17805
rect 24949 17765 24961 17799
rect 24995 17796 25007 17799
rect 25038 17796 25044 17808
rect 24995 17768 25044 17796
rect 24995 17765 25007 17768
rect 24949 17759 25007 17765
rect 24728 17700 24808 17728
rect 24728 17688 24734 17700
rect 24486 17660 24492 17672
rect 23952 17632 24492 17660
rect 21876 17620 21882 17632
rect 24486 17620 24492 17632
rect 24544 17660 24550 17672
rect 24964 17660 24992 17759
rect 25038 17756 25044 17768
rect 25096 17756 25102 17808
rect 25148 17796 25176 17836
rect 25332 17836 25437 17864
rect 25222 17796 25228 17808
rect 25148 17768 25228 17796
rect 25222 17756 25228 17768
rect 25280 17756 25286 17808
rect 25133 17731 25191 17737
rect 25133 17697 25145 17731
rect 25179 17728 25191 17731
rect 25332 17728 25360 17836
rect 25425 17833 25437 17836
rect 25471 17833 25483 17867
rect 25425 17827 25483 17833
rect 25593 17867 25651 17873
rect 25593 17833 25605 17867
rect 25639 17833 25651 17867
rect 25593 17827 25651 17833
rect 25869 17867 25927 17873
rect 25869 17833 25881 17867
rect 25915 17864 25927 17867
rect 25958 17864 25964 17876
rect 25915 17836 25964 17864
rect 25915 17833 25927 17836
rect 25869 17827 25927 17833
rect 25179 17700 25360 17728
rect 25608 17728 25636 17827
rect 25958 17824 25964 17836
rect 26016 17824 26022 17876
rect 25685 17731 25743 17737
rect 25685 17728 25697 17731
rect 25608 17700 25697 17728
rect 25179 17697 25191 17700
rect 25133 17691 25191 17697
rect 25685 17697 25697 17700
rect 25731 17697 25743 17731
rect 25685 17691 25743 17697
rect 24544 17632 24992 17660
rect 24544 17620 24550 17632
rect 20254 17592 20260 17604
rect 19996 17564 20260 17592
rect 20254 17552 20260 17564
rect 20312 17592 20318 17604
rect 24854 17592 24860 17604
rect 20312 17564 22692 17592
rect 20312 17552 20318 17564
rect 14829 17527 14887 17533
rect 14829 17524 14841 17527
rect 14792 17496 14841 17524
rect 14792 17484 14798 17496
rect 14829 17493 14841 17496
rect 14875 17493 14887 17527
rect 14829 17487 14887 17493
rect 15197 17527 15255 17533
rect 15197 17493 15209 17527
rect 15243 17524 15255 17527
rect 15749 17527 15807 17533
rect 15749 17524 15761 17527
rect 15243 17496 15761 17524
rect 15243 17493 15255 17496
rect 15197 17487 15255 17493
rect 15749 17493 15761 17496
rect 15795 17493 15807 17527
rect 15749 17487 15807 17493
rect 15930 17484 15936 17536
rect 15988 17484 15994 17536
rect 16298 17484 16304 17536
rect 16356 17524 16362 17536
rect 17221 17527 17279 17533
rect 17221 17524 17233 17527
rect 16356 17496 17233 17524
rect 16356 17484 16362 17496
rect 17221 17493 17233 17496
rect 17267 17524 17279 17527
rect 18414 17524 18420 17536
rect 17267 17496 18420 17524
rect 17267 17493 17279 17496
rect 17221 17487 17279 17493
rect 18414 17484 18420 17496
rect 18472 17484 18478 17536
rect 19242 17484 19248 17536
rect 19300 17484 19306 17536
rect 19610 17484 19616 17536
rect 19668 17484 19674 17536
rect 21634 17484 21640 17536
rect 21692 17484 21698 17536
rect 22189 17527 22247 17533
rect 22189 17493 22201 17527
rect 22235 17524 22247 17527
rect 22554 17524 22560 17536
rect 22235 17496 22560 17524
rect 22235 17493 22247 17496
rect 22189 17487 22247 17493
rect 22554 17484 22560 17496
rect 22612 17484 22618 17536
rect 22664 17533 22692 17564
rect 24044 17564 24860 17592
rect 22649 17527 22707 17533
rect 22649 17493 22661 17527
rect 22695 17524 22707 17527
rect 23290 17524 23296 17536
rect 22695 17496 23296 17524
rect 22695 17493 22707 17496
rect 22649 17487 22707 17493
rect 23290 17484 23296 17496
rect 23348 17484 23354 17536
rect 23750 17484 23756 17536
rect 23808 17524 23814 17536
rect 24044 17533 24072 17564
rect 24854 17552 24860 17564
rect 24912 17592 24918 17604
rect 24912 17564 25452 17592
rect 24912 17552 24918 17564
rect 24029 17527 24087 17533
rect 24029 17524 24041 17527
rect 23808 17496 24041 17524
rect 23808 17484 23814 17496
rect 24029 17493 24041 17496
rect 24075 17493 24087 17527
rect 24029 17487 24087 17493
rect 24394 17484 24400 17536
rect 24452 17484 24458 17536
rect 24581 17527 24639 17533
rect 24581 17493 24593 17527
rect 24627 17524 24639 17527
rect 25130 17524 25136 17536
rect 24627 17496 25136 17524
rect 24627 17493 24639 17496
rect 24581 17487 24639 17493
rect 25130 17484 25136 17496
rect 25188 17484 25194 17536
rect 25424 17533 25452 17564
rect 25409 17527 25467 17533
rect 25409 17493 25421 17527
rect 25455 17493 25467 17527
rect 25409 17487 25467 17493
rect 552 17434 27416 17456
rect 552 17382 3756 17434
rect 3808 17382 3820 17434
rect 3872 17382 3884 17434
rect 3936 17382 3948 17434
rect 4000 17382 4012 17434
rect 4064 17382 10472 17434
rect 10524 17382 10536 17434
rect 10588 17382 10600 17434
rect 10652 17382 10664 17434
rect 10716 17382 10728 17434
rect 10780 17382 17188 17434
rect 17240 17382 17252 17434
rect 17304 17382 17316 17434
rect 17368 17382 17380 17434
rect 17432 17382 17444 17434
rect 17496 17382 23904 17434
rect 23956 17382 23968 17434
rect 24020 17382 24032 17434
rect 24084 17382 24096 17434
rect 24148 17382 24160 17434
rect 24212 17382 27416 17434
rect 552 17360 27416 17382
rect 1394 17280 1400 17332
rect 1452 17280 1458 17332
rect 1762 17280 1768 17332
rect 1820 17280 1826 17332
rect 2774 17280 2780 17332
rect 2832 17280 2838 17332
rect 4154 17280 4160 17332
rect 4212 17280 4218 17332
rect 4246 17280 4252 17332
rect 4304 17320 4310 17332
rect 4341 17323 4399 17329
rect 4341 17320 4353 17323
rect 4304 17292 4353 17320
rect 4304 17280 4310 17292
rect 4341 17289 4353 17292
rect 4387 17289 4399 17323
rect 4341 17283 4399 17289
rect 4525 17323 4583 17329
rect 4525 17289 4537 17323
rect 4571 17320 4583 17323
rect 4614 17320 4620 17332
rect 4571 17292 4620 17320
rect 4571 17289 4583 17292
rect 4525 17283 4583 17289
rect 4614 17280 4620 17292
rect 4672 17280 4678 17332
rect 5997 17323 6055 17329
rect 5997 17289 6009 17323
rect 6043 17320 6055 17323
rect 6181 17323 6239 17329
rect 6181 17320 6193 17323
rect 6043 17292 6193 17320
rect 6043 17289 6055 17292
rect 5997 17283 6055 17289
rect 6181 17289 6193 17292
rect 6227 17289 6239 17323
rect 6181 17283 6239 17289
rect 6638 17280 6644 17332
rect 6696 17320 6702 17332
rect 6825 17323 6883 17329
rect 6825 17320 6837 17323
rect 6696 17292 6837 17320
rect 6696 17280 6702 17292
rect 6825 17289 6837 17292
rect 6871 17289 6883 17323
rect 9030 17320 9036 17332
rect 6825 17283 6883 17289
rect 8404 17292 9036 17320
rect 1780 17184 1808 17280
rect 2593 17255 2651 17261
rect 2593 17221 2605 17255
rect 2639 17252 2651 17255
rect 2958 17252 2964 17264
rect 2639 17224 2964 17252
rect 2639 17221 2651 17224
rect 2593 17215 2651 17221
rect 2958 17212 2964 17224
rect 3016 17252 3022 17264
rect 3973 17255 4031 17261
rect 3973 17252 3985 17255
rect 3016 17224 3985 17252
rect 3016 17212 3022 17224
rect 3973 17221 3985 17224
rect 4019 17221 4031 17255
rect 3973 17215 4031 17221
rect 1857 17187 1915 17193
rect 1857 17184 1869 17187
rect 1780 17156 1869 17184
rect 1857 17153 1869 17156
rect 1903 17153 1915 17187
rect 1857 17147 1915 17153
rect 1946 17144 1952 17196
rect 2004 17184 2010 17196
rect 2498 17184 2504 17196
rect 2004 17156 2504 17184
rect 2004 17144 2010 17156
rect 2498 17144 2504 17156
rect 2556 17144 2562 17196
rect 1581 17119 1639 17125
rect 1581 17085 1593 17119
rect 1627 17116 1639 17119
rect 1670 17116 1676 17128
rect 1627 17088 1676 17116
rect 1627 17085 1639 17088
rect 1581 17079 1639 17085
rect 1670 17076 1676 17088
rect 1728 17076 1734 17128
rect 1765 17119 1823 17125
rect 1765 17085 1777 17119
rect 1811 17116 1823 17119
rect 1964 17116 1992 17144
rect 3510 17116 3516 17128
rect 1811 17088 1992 17116
rect 2424 17088 3516 17116
rect 1811 17085 1823 17088
rect 1765 17079 1823 17085
rect 2424 16992 2452 17088
rect 3510 17076 3516 17088
rect 3568 17116 3574 17128
rect 3789 17119 3847 17125
rect 3789 17116 3801 17119
rect 3568 17088 3801 17116
rect 3568 17076 3574 17088
rect 3789 17085 3801 17088
rect 3835 17085 3847 17119
rect 3789 17079 3847 17085
rect 2961 17051 3019 17057
rect 2961 17017 2973 17051
rect 3007 17048 3019 17051
rect 3326 17048 3332 17060
rect 3007 17020 3332 17048
rect 3007 17017 3019 17020
rect 2961 17011 3019 17017
rect 3326 17008 3332 17020
rect 3384 17008 3390 17060
rect 4172 17048 4200 17280
rect 8404 17252 8432 17292
rect 9030 17280 9036 17292
rect 9088 17280 9094 17332
rect 9122 17280 9128 17332
rect 9180 17320 9186 17332
rect 9674 17320 9680 17332
rect 9180 17292 9680 17320
rect 9180 17280 9186 17292
rect 9674 17280 9680 17292
rect 9732 17280 9738 17332
rect 10594 17280 10600 17332
rect 10652 17320 10658 17332
rect 10962 17320 10968 17332
rect 10652 17292 10968 17320
rect 10652 17280 10658 17292
rect 10962 17280 10968 17292
rect 11020 17320 11026 17332
rect 14001 17323 14059 17329
rect 11020 17292 13952 17320
rect 11020 17280 11026 17292
rect 6564 17224 8432 17252
rect 9769 17255 9827 17261
rect 6270 17184 6276 17196
rect 6012 17156 6276 17184
rect 4617 17119 4675 17125
rect 4617 17085 4629 17119
rect 4663 17116 4675 17119
rect 6012 17116 6040 17156
rect 6270 17144 6276 17156
rect 6328 17144 6334 17196
rect 6564 17193 6592 17224
rect 9769 17221 9781 17255
rect 9815 17252 9827 17255
rect 10781 17255 10839 17261
rect 10781 17252 10793 17255
rect 9815 17224 10088 17252
rect 9815 17221 9827 17224
rect 9769 17215 9827 17221
rect 6549 17187 6607 17193
rect 6549 17153 6561 17187
rect 6595 17153 6607 17187
rect 6549 17147 6607 17153
rect 7926 17144 7932 17196
rect 7984 17184 7990 17196
rect 7984 17156 8156 17184
rect 7984 17144 7990 17156
rect 4663 17088 6040 17116
rect 4663 17085 4675 17088
rect 4617 17079 4675 17085
rect 6086 17076 6092 17128
rect 6144 17076 6150 17128
rect 7006 17076 7012 17128
rect 7064 17076 7070 17128
rect 7745 17119 7803 17125
rect 7745 17116 7757 17119
rect 7484 17088 7757 17116
rect 4890 17057 4896 17060
rect 4341 17051 4399 17057
rect 4341 17048 4353 17051
rect 4172 17020 4353 17048
rect 4341 17017 4353 17020
rect 4387 17017 4399 17051
rect 4884 17048 4896 17057
rect 4851 17020 4896 17048
rect 4341 17011 4399 17017
rect 4884 17011 4896 17020
rect 4890 17008 4896 17011
rect 4948 17008 4954 17060
rect 6914 17008 6920 17060
rect 6972 17048 6978 17060
rect 7484 17048 7512 17088
rect 7745 17085 7757 17088
rect 7791 17116 7803 17119
rect 8018 17116 8024 17128
rect 7791 17088 8024 17116
rect 7791 17085 7803 17088
rect 7745 17079 7803 17085
rect 8018 17076 8024 17088
rect 8076 17076 8082 17128
rect 8128 17125 8156 17156
rect 10060 17128 10088 17224
rect 10244 17224 10793 17252
rect 10244 17196 10272 17224
rect 10781 17221 10793 17224
rect 10827 17221 10839 17255
rect 10781 17215 10839 17221
rect 11977 17255 12035 17261
rect 11977 17221 11989 17255
rect 12023 17221 12035 17255
rect 13924 17252 13952 17292
rect 14001 17289 14013 17323
rect 14047 17320 14059 17323
rect 14182 17320 14188 17332
rect 14047 17292 14188 17320
rect 14047 17289 14059 17292
rect 14001 17283 14059 17289
rect 14182 17280 14188 17292
rect 14240 17280 14246 17332
rect 15010 17280 15016 17332
rect 15068 17320 15074 17332
rect 16298 17320 16304 17332
rect 15068 17292 16304 17320
rect 15068 17280 15074 17292
rect 16298 17280 16304 17292
rect 16356 17280 16362 17332
rect 17313 17323 17371 17329
rect 17313 17320 17325 17323
rect 16408 17292 17325 17320
rect 16408 17252 16436 17292
rect 17313 17289 17325 17292
rect 17359 17289 17371 17323
rect 17313 17283 17371 17289
rect 17497 17323 17555 17329
rect 17497 17289 17509 17323
rect 17543 17320 17555 17323
rect 17770 17320 17776 17332
rect 17543 17292 17776 17320
rect 17543 17289 17555 17292
rect 17497 17283 17555 17289
rect 13924 17224 16436 17252
rect 11977 17215 12035 17221
rect 10226 17144 10232 17196
rect 10284 17144 10290 17196
rect 10318 17144 10324 17196
rect 10376 17144 10382 17196
rect 11241 17187 11299 17193
rect 11241 17184 11253 17187
rect 10888 17156 11253 17184
rect 8113 17119 8171 17125
rect 8113 17085 8125 17119
rect 8159 17085 8171 17119
rect 8113 17079 8171 17085
rect 8205 17119 8263 17125
rect 8205 17085 8217 17119
rect 8251 17116 8263 17119
rect 8389 17119 8447 17125
rect 8251 17088 8340 17116
rect 8251 17085 8263 17088
rect 8205 17079 8263 17085
rect 8312 17060 8340 17088
rect 8389 17085 8401 17119
rect 8435 17116 8447 17119
rect 9950 17116 9956 17128
rect 8435 17088 9956 17116
rect 8435 17085 8447 17088
rect 8389 17079 8447 17085
rect 9950 17076 9956 17088
rect 10008 17076 10014 17128
rect 10042 17076 10048 17128
rect 10100 17076 10106 17128
rect 10410 17125 10416 17128
rect 10409 17116 10416 17125
rect 10371 17088 10416 17116
rect 10409 17079 10416 17088
rect 10410 17076 10416 17079
rect 10468 17076 10474 17128
rect 10502 17076 10508 17128
rect 10560 17116 10566 17128
rect 10888 17125 10916 17156
rect 11241 17153 11253 17156
rect 11287 17153 11299 17187
rect 11241 17147 11299 17153
rect 10597 17119 10655 17125
rect 10597 17116 10609 17119
rect 10560 17088 10609 17116
rect 10560 17076 10566 17088
rect 10597 17085 10609 17088
rect 10643 17085 10655 17119
rect 10597 17079 10655 17085
rect 10873 17119 10931 17125
rect 10873 17085 10885 17119
rect 10919 17116 10931 17119
rect 10962 17116 10968 17128
rect 10919 17088 10968 17116
rect 10919 17085 10931 17088
rect 10873 17079 10931 17085
rect 10962 17076 10968 17088
rect 11020 17076 11026 17128
rect 11146 17076 11152 17128
rect 11204 17116 11210 17128
rect 11992 17116 12020 17215
rect 16482 17212 16488 17264
rect 16540 17252 16546 17264
rect 17328 17252 17356 17283
rect 17770 17280 17776 17292
rect 17828 17280 17834 17332
rect 18156 17292 19932 17320
rect 17954 17252 17960 17264
rect 16540 17224 16988 17252
rect 17328 17224 17960 17252
rect 16540 17212 16546 17224
rect 13906 17144 13912 17196
rect 13964 17144 13970 17196
rect 13998 17144 14004 17196
rect 14056 17184 14062 17196
rect 15010 17184 15016 17196
rect 14056 17156 15016 17184
rect 14056 17144 14062 17156
rect 15010 17144 15016 17156
rect 15068 17144 15074 17196
rect 16960 17184 16988 17224
rect 17954 17212 17960 17224
rect 18012 17212 18018 17264
rect 18046 17184 18052 17196
rect 16316 17156 16896 17184
rect 16960 17156 18052 17184
rect 13357 17119 13415 17125
rect 13357 17116 13369 17119
rect 11204 17088 12020 17116
rect 12452 17088 13369 17116
rect 11204 17076 11210 17088
rect 12452 17060 12480 17088
rect 13357 17085 13369 17088
rect 13403 17085 13415 17119
rect 13924 17116 13952 17144
rect 13357 17079 13415 17085
rect 13464 17088 13952 17116
rect 14185 17119 14243 17125
rect 6972 17020 7512 17048
rect 6972 17008 6978 17020
rect 7558 17008 7564 17060
rect 7616 17048 7622 17060
rect 7616 17020 8156 17048
rect 7616 17008 7622 17020
rect 2406 16940 2412 16992
rect 2464 16940 2470 16992
rect 2498 16940 2504 16992
rect 2556 16980 2562 16992
rect 2751 16983 2809 16989
rect 2751 16980 2763 16983
rect 2556 16952 2763 16980
rect 2556 16940 2562 16952
rect 2751 16949 2763 16952
rect 2797 16949 2809 16983
rect 2751 16943 2809 16949
rect 3234 16940 3240 16992
rect 3292 16940 3298 16992
rect 8018 16940 8024 16992
rect 8076 16940 8082 16992
rect 8128 16980 8156 17020
rect 8294 17008 8300 17060
rect 8352 17008 8358 17060
rect 8656 17051 8714 17057
rect 8656 17017 8668 17051
rect 8702 17048 8714 17051
rect 9030 17048 9036 17060
rect 8702 17020 9036 17048
rect 8702 17017 8714 17020
rect 8656 17011 8714 17017
rect 9030 17008 9036 17020
rect 9088 17008 9094 17060
rect 12434 17008 12440 17060
rect 12492 17008 12498 17060
rect 13112 17051 13170 17057
rect 13112 17017 13124 17051
rect 13158 17048 13170 17051
rect 13464 17048 13492 17088
rect 14185 17085 14197 17119
rect 14231 17116 14243 17119
rect 14274 17116 14280 17128
rect 14231 17088 14280 17116
rect 14231 17085 14243 17088
rect 14185 17079 14243 17085
rect 14274 17076 14280 17088
rect 14332 17076 14338 17128
rect 16316 17125 16344 17156
rect 16301 17119 16359 17125
rect 16301 17116 16313 17119
rect 14752 17088 16313 17116
rect 14752 17060 14780 17088
rect 16301 17085 16313 17088
rect 16347 17085 16359 17119
rect 16301 17079 16359 17085
rect 16577 17119 16635 17125
rect 16577 17085 16589 17119
rect 16623 17116 16635 17119
rect 16666 17116 16672 17128
rect 16623 17088 16672 17116
rect 16623 17085 16635 17088
rect 16577 17079 16635 17085
rect 16666 17076 16672 17088
rect 16724 17076 16730 17128
rect 16758 17076 16764 17128
rect 16816 17076 16822 17128
rect 16868 17125 16896 17156
rect 18046 17144 18052 17156
rect 18104 17144 18110 17196
rect 16853 17119 16911 17125
rect 16853 17085 16865 17119
rect 16899 17085 16911 17119
rect 16853 17079 16911 17085
rect 16942 17076 16948 17128
rect 17000 17076 17006 17128
rect 17126 17076 17132 17128
rect 17184 17116 17190 17128
rect 18156 17116 18184 17292
rect 19904 17184 19932 17292
rect 20254 17280 20260 17332
rect 20312 17280 20318 17332
rect 21818 17280 21824 17332
rect 21876 17280 21882 17332
rect 24394 17280 24400 17332
rect 24452 17320 24458 17332
rect 25133 17323 25191 17329
rect 25133 17320 25145 17323
rect 24452 17292 25145 17320
rect 24452 17280 24458 17292
rect 25133 17289 25145 17292
rect 25179 17320 25191 17323
rect 25179 17292 25452 17320
rect 25179 17289 25191 17292
rect 25133 17283 25191 17289
rect 19904 17156 20576 17184
rect 17184 17088 18184 17116
rect 17184 17076 17190 17088
rect 18874 17076 18880 17128
rect 18932 17116 18938 17128
rect 19426 17116 19432 17128
rect 18932 17088 19432 17116
rect 18932 17076 18938 17088
rect 19426 17076 19432 17088
rect 19484 17116 19490 17128
rect 20441 17119 20499 17125
rect 20441 17116 20453 17119
rect 19484 17088 20453 17116
rect 19484 17076 19490 17088
rect 20441 17085 20453 17088
rect 20487 17085 20499 17119
rect 20548 17116 20576 17156
rect 21836 17116 21864 17280
rect 22462 17212 22468 17264
rect 22520 17212 22526 17264
rect 22738 17212 22744 17264
rect 22796 17252 22802 17264
rect 23934 17252 23940 17264
rect 22796 17224 23940 17252
rect 22796 17212 22802 17224
rect 22480 17184 22508 17212
rect 23492 17193 23520 17224
rect 23934 17212 23940 17224
rect 23992 17212 23998 17264
rect 23477 17187 23535 17193
rect 22480 17156 22692 17184
rect 22664 17125 22692 17156
rect 22940 17156 23244 17184
rect 22511 17119 22569 17125
rect 22511 17116 22523 17119
rect 20548 17088 21404 17116
rect 21836 17088 22523 17116
rect 20441 17079 20499 17085
rect 13158 17020 13492 17048
rect 13158 17017 13170 17020
rect 13112 17011 13170 17017
rect 13538 17008 13544 17060
rect 13596 17008 13602 17060
rect 13725 17051 13783 17057
rect 13725 17017 13737 17051
rect 13771 17048 13783 17051
rect 13814 17048 13820 17060
rect 13771 17020 13820 17048
rect 13771 17017 13783 17020
rect 13725 17011 13783 17017
rect 13814 17008 13820 17020
rect 13872 17008 13878 17060
rect 13909 17051 13967 17057
rect 13909 17017 13921 17051
rect 13955 17048 13967 17051
rect 14734 17048 14740 17060
rect 13955 17020 14740 17048
rect 13955 17017 13967 17020
rect 13909 17011 13967 17017
rect 14734 17008 14740 17020
rect 14792 17008 14798 17060
rect 16114 17008 16120 17060
rect 16172 17008 16178 17060
rect 16960 17048 16988 17076
rect 17957 17051 18015 17057
rect 17957 17048 17969 17051
rect 16960 17020 17969 17048
rect 17957 17017 17969 17020
rect 18003 17048 18015 17051
rect 18966 17048 18972 17060
rect 18003 17020 18972 17048
rect 18003 17017 18015 17020
rect 17957 17011 18015 17017
rect 18966 17008 18972 17020
rect 19024 17008 19030 17060
rect 19144 17051 19202 17057
rect 19144 17017 19156 17051
rect 19190 17048 19202 17051
rect 19242 17048 19248 17060
rect 19190 17020 19248 17048
rect 19190 17017 19202 17020
rect 19144 17011 19202 17017
rect 19242 17008 19248 17020
rect 19300 17008 19306 17060
rect 20346 17008 20352 17060
rect 20404 17048 20410 17060
rect 20686 17051 20744 17057
rect 20686 17048 20698 17051
rect 20404 17020 20698 17048
rect 20404 17008 20410 17020
rect 20686 17017 20698 17020
rect 20732 17017 20744 17051
rect 20686 17011 20744 17017
rect 21376 16992 21404 17088
rect 22511 17085 22523 17088
rect 22557 17085 22569 17119
rect 22511 17079 22569 17085
rect 22649 17119 22707 17125
rect 22649 17085 22661 17119
rect 22695 17085 22707 17119
rect 22649 17079 22707 17085
rect 22741 17119 22799 17125
rect 22741 17085 22753 17119
rect 22787 17116 22799 17119
rect 22830 17116 22836 17128
rect 22787 17088 22836 17116
rect 22787 17085 22799 17088
rect 22741 17079 22799 17085
rect 9861 16983 9919 16989
rect 9861 16980 9873 16983
rect 8128 16952 9873 16980
rect 9861 16949 9873 16952
rect 9907 16949 9919 16983
rect 9861 16943 9919 16949
rect 10134 16940 10140 16992
rect 10192 16980 10198 16992
rect 11057 16983 11115 16989
rect 11057 16980 11069 16983
rect 10192 16952 11069 16980
rect 10192 16940 10198 16952
rect 11057 16949 11069 16952
rect 11103 16949 11115 16983
rect 11057 16943 11115 16949
rect 11882 16940 11888 16992
rect 11940 16940 11946 16992
rect 14826 16940 14832 16992
rect 14884 16940 14890 16992
rect 16298 16940 16304 16992
rect 16356 16940 16362 16992
rect 16942 16940 16948 16992
rect 17000 16940 17006 16992
rect 17862 16940 17868 16992
rect 17920 16940 17926 16992
rect 21358 16940 21364 16992
rect 21416 16940 21422 16992
rect 22370 16940 22376 16992
rect 22428 16940 22434 16992
rect 22664 16980 22692 17079
rect 22830 17076 22836 17088
rect 22888 17076 22894 17128
rect 22940 17125 22968 17156
rect 23216 17128 23244 17156
rect 23477 17153 23489 17187
rect 23523 17153 23535 17187
rect 24854 17184 24860 17196
rect 23477 17147 23535 17153
rect 24780 17156 24860 17184
rect 22924 17119 22982 17125
rect 22924 17085 22936 17119
rect 22970 17085 22982 17119
rect 22924 17079 22982 17085
rect 23017 17119 23075 17125
rect 23017 17085 23029 17119
rect 23063 17116 23075 17119
rect 23063 17088 23152 17116
rect 23063 17085 23075 17088
rect 23017 17079 23075 17085
rect 23124 16992 23152 17088
rect 23198 17076 23204 17128
rect 23256 17076 23262 17128
rect 23290 17076 23296 17128
rect 23348 17076 23354 17128
rect 24780 17125 24808 17156
rect 24854 17144 24860 17156
rect 24912 17144 24918 17196
rect 24964 17156 25360 17184
rect 24029 17119 24087 17125
rect 24029 17085 24041 17119
rect 24075 17116 24087 17119
rect 24765 17119 24823 17125
rect 24075 17088 24716 17116
rect 24075 17085 24087 17088
rect 24029 17079 24087 17085
rect 24688 17057 24716 17088
rect 24765 17085 24777 17119
rect 24811 17085 24823 17119
rect 24964 17116 24992 17156
rect 25332 17128 25360 17156
rect 24765 17079 24823 17085
rect 24872 17088 24992 17116
rect 24673 17051 24731 17057
rect 24673 17017 24685 17051
rect 24719 17048 24731 17051
rect 24872 17048 24900 17088
rect 25038 17076 25044 17128
rect 25096 17116 25102 17128
rect 25225 17119 25283 17125
rect 25225 17116 25237 17119
rect 25096 17088 25237 17116
rect 25096 17076 25102 17088
rect 25225 17085 25237 17088
rect 25271 17085 25283 17119
rect 25225 17079 25283 17085
rect 25314 17076 25320 17128
rect 25372 17076 25378 17128
rect 25424 17125 25452 17292
rect 25498 17144 25504 17196
rect 25556 17144 25562 17196
rect 25409 17119 25467 17125
rect 25409 17085 25421 17119
rect 25455 17085 25467 17119
rect 25409 17079 25467 17085
rect 24719 17020 24900 17048
rect 24719 17017 24731 17020
rect 24673 17011 24731 17017
rect 24946 17008 24952 17060
rect 25004 17008 25010 17060
rect 25774 17057 25780 17060
rect 25056 17020 25360 17048
rect 25056 16992 25084 17020
rect 23014 16980 23020 16992
rect 22664 16952 23020 16980
rect 23014 16940 23020 16952
rect 23072 16940 23078 16992
rect 23106 16940 23112 16992
rect 23164 16940 23170 16992
rect 24118 16940 24124 16992
rect 24176 16940 24182 16992
rect 24210 16940 24216 16992
rect 24268 16980 24274 16992
rect 24305 16983 24363 16989
rect 24305 16980 24317 16983
rect 24268 16952 24317 16980
rect 24268 16940 24274 16952
rect 24305 16949 24317 16952
rect 24351 16949 24363 16983
rect 24305 16943 24363 16949
rect 24394 16940 24400 16992
rect 24452 16940 24458 16992
rect 24489 16983 24547 16989
rect 24489 16949 24501 16983
rect 24535 16980 24547 16983
rect 25038 16980 25044 16992
rect 24535 16952 25044 16980
rect 24535 16949 24547 16952
rect 24489 16943 24547 16949
rect 25038 16940 25044 16952
rect 25096 16940 25102 16992
rect 25222 16940 25228 16992
rect 25280 16940 25286 16992
rect 25332 16980 25360 17020
rect 25768 17011 25780 17057
rect 25774 17008 25780 17011
rect 25832 17008 25838 17060
rect 26881 16983 26939 16989
rect 26881 16980 26893 16983
rect 25332 16952 26893 16980
rect 26881 16949 26893 16952
rect 26927 16949 26939 16983
rect 26881 16943 26939 16949
rect 552 16890 27576 16912
rect 552 16838 7114 16890
rect 7166 16838 7178 16890
rect 7230 16838 7242 16890
rect 7294 16838 7306 16890
rect 7358 16838 7370 16890
rect 7422 16838 13830 16890
rect 13882 16838 13894 16890
rect 13946 16838 13958 16890
rect 14010 16838 14022 16890
rect 14074 16838 14086 16890
rect 14138 16838 20546 16890
rect 20598 16838 20610 16890
rect 20662 16838 20674 16890
rect 20726 16838 20738 16890
rect 20790 16838 20802 16890
rect 20854 16838 27262 16890
rect 27314 16838 27326 16890
rect 27378 16838 27390 16890
rect 27442 16838 27454 16890
rect 27506 16838 27518 16890
rect 27570 16838 27576 16890
rect 552 16816 27576 16838
rect 2406 16736 2412 16788
rect 2464 16736 2470 16788
rect 3237 16779 3295 16785
rect 3237 16745 3249 16779
rect 3283 16776 3295 16779
rect 3326 16776 3332 16788
rect 3283 16748 3332 16776
rect 3283 16745 3295 16748
rect 3237 16739 3295 16745
rect 3326 16736 3332 16748
rect 3384 16736 3390 16788
rect 4430 16736 4436 16788
rect 4488 16736 4494 16788
rect 7009 16779 7067 16785
rect 7009 16776 7021 16779
rect 6932 16748 7021 16776
rect 1026 16600 1032 16652
rect 1084 16600 1090 16652
rect 1296 16643 1354 16649
rect 1296 16609 1308 16643
rect 1342 16640 1354 16643
rect 1342 16612 2084 16640
rect 1342 16609 1354 16612
rect 1296 16603 1354 16609
rect 2056 16572 2084 16612
rect 2682 16600 2688 16652
rect 2740 16600 2746 16652
rect 2866 16600 2872 16652
rect 2924 16640 2930 16652
rect 2961 16643 3019 16649
rect 2961 16640 2973 16643
rect 2924 16612 2973 16640
rect 2924 16600 2930 16612
rect 2961 16609 2973 16612
rect 3007 16640 3019 16643
rect 3234 16640 3240 16652
rect 3007 16612 3240 16640
rect 3007 16609 3019 16612
rect 2961 16603 3019 16609
rect 3234 16600 3240 16612
rect 3292 16600 3298 16652
rect 4361 16643 4419 16649
rect 4361 16609 4373 16643
rect 4407 16640 4419 16643
rect 4448 16640 4476 16736
rect 6932 16652 6960 16748
rect 7009 16745 7021 16748
rect 7055 16745 7067 16779
rect 7009 16739 7067 16745
rect 7834 16736 7840 16788
rect 7892 16736 7898 16788
rect 8018 16736 8024 16788
rect 8076 16736 8082 16788
rect 8478 16736 8484 16788
rect 8536 16776 8542 16788
rect 8536 16748 8984 16776
rect 8536 16736 8542 16748
rect 7852 16708 7880 16736
rect 7929 16711 7987 16717
rect 7929 16708 7941 16711
rect 7024 16680 7604 16708
rect 7024 16652 7052 16680
rect 7576 16652 7604 16680
rect 7668 16680 7941 16708
rect 4407 16612 4476 16640
rect 4407 16609 4419 16612
rect 4361 16603 4419 16609
rect 6822 16600 6828 16652
rect 6880 16600 6886 16652
rect 6914 16600 6920 16652
rect 6972 16600 6978 16652
rect 7006 16600 7012 16652
rect 7064 16600 7070 16652
rect 7558 16600 7564 16652
rect 7616 16600 7622 16652
rect 7668 16649 7696 16680
rect 7929 16677 7941 16680
rect 7975 16677 7987 16711
rect 8036 16708 8064 16736
rect 8956 16708 8984 16748
rect 9030 16736 9036 16788
rect 9088 16736 9094 16788
rect 10226 16776 10232 16788
rect 10152 16748 10232 16776
rect 10152 16717 10180 16748
rect 10226 16736 10232 16748
rect 10284 16736 10290 16788
rect 10318 16736 10324 16788
rect 10376 16776 10382 16788
rect 10505 16779 10563 16785
rect 10505 16776 10517 16779
rect 10376 16748 10517 16776
rect 10376 16736 10382 16748
rect 10505 16745 10517 16748
rect 10551 16745 10563 16779
rect 10505 16739 10563 16745
rect 10870 16736 10876 16788
rect 10928 16736 10934 16788
rect 10962 16736 10968 16788
rect 11020 16736 11026 16788
rect 13078 16736 13084 16788
rect 13136 16776 13142 16788
rect 13265 16779 13323 16785
rect 13265 16776 13277 16779
rect 13136 16748 13277 16776
rect 13136 16736 13142 16748
rect 13265 16745 13277 16748
rect 13311 16776 13323 16779
rect 15102 16776 15108 16788
rect 13311 16748 15108 16776
rect 13311 16745 13323 16748
rect 13265 16739 13323 16745
rect 15102 16736 15108 16748
rect 15160 16736 15166 16788
rect 15197 16779 15255 16785
rect 15197 16745 15209 16779
rect 15243 16776 15255 16779
rect 15243 16748 15424 16776
rect 15243 16745 15255 16748
rect 15197 16739 15255 16745
rect 9125 16711 9183 16717
rect 9125 16708 9137 16711
rect 8036 16680 8524 16708
rect 8956 16680 9137 16708
rect 7929 16671 7987 16677
rect 7653 16643 7711 16649
rect 7653 16609 7665 16643
rect 7699 16609 7711 16643
rect 7653 16603 7711 16609
rect 7837 16643 7895 16649
rect 7837 16609 7849 16643
rect 7883 16640 7895 16643
rect 8113 16643 8171 16649
rect 8113 16640 8125 16643
rect 7883 16612 8125 16640
rect 7883 16609 7895 16612
rect 7837 16603 7895 16609
rect 8113 16609 8125 16612
rect 8159 16640 8171 16643
rect 8202 16640 8208 16652
rect 8159 16612 8208 16640
rect 8159 16609 8171 16612
rect 8113 16603 8171 16609
rect 8202 16600 8208 16612
rect 8260 16600 8266 16652
rect 8297 16643 8355 16649
rect 8297 16609 8309 16643
rect 8343 16638 8355 16643
rect 8386 16638 8392 16652
rect 8343 16610 8392 16638
rect 8343 16609 8355 16610
rect 8297 16603 8355 16609
rect 8386 16600 8392 16610
rect 8444 16600 8450 16652
rect 8496 16649 8524 16680
rect 9125 16677 9137 16680
rect 9171 16677 9183 16711
rect 10137 16711 10195 16717
rect 9125 16671 9183 16677
rect 9355 16677 9413 16683
rect 9355 16674 9367 16677
rect 8481 16643 8539 16649
rect 8481 16609 8493 16643
rect 8527 16609 8539 16643
rect 8481 16603 8539 16609
rect 8570 16600 8576 16652
rect 8628 16640 8634 16652
rect 9340 16643 9367 16674
rect 9401 16643 9413 16677
rect 10137 16677 10149 16711
rect 10183 16677 10195 16711
rect 10888 16708 10916 16736
rect 10137 16671 10195 16677
rect 10244 16680 10916 16708
rect 12452 16680 13860 16708
rect 9340 16640 9413 16643
rect 8628 16637 9413 16640
rect 9953 16643 10011 16649
rect 8628 16612 9368 16637
rect 8628 16600 8634 16612
rect 9953 16609 9965 16643
rect 9999 16640 10011 16643
rect 10042 16640 10048 16652
rect 9999 16612 10048 16640
rect 9999 16609 10011 16612
rect 9953 16603 10011 16609
rect 10042 16600 10048 16612
rect 10100 16600 10106 16652
rect 10244 16649 10272 16680
rect 12452 16652 12480 16680
rect 10229 16643 10287 16649
rect 10229 16640 10241 16643
rect 10152 16612 10241 16640
rect 2501 16575 2559 16581
rect 2501 16572 2513 16575
rect 2056 16544 2513 16572
rect 2501 16541 2513 16544
rect 2547 16541 2559 16575
rect 2501 16535 2559 16541
rect 4617 16575 4675 16581
rect 4617 16541 4629 16575
rect 4663 16541 4675 16575
rect 4617 16535 4675 16541
rect 2869 16507 2927 16513
rect 2869 16473 2881 16507
rect 2915 16504 2927 16507
rect 2958 16504 2964 16516
rect 2915 16476 2964 16504
rect 2915 16473 2927 16476
rect 2869 16467 2927 16473
rect 2958 16464 2964 16476
rect 3016 16464 3022 16516
rect 4430 16396 4436 16448
rect 4488 16436 4494 16448
rect 4632 16436 4660 16535
rect 6546 16532 6552 16584
rect 6604 16532 6610 16584
rect 6638 16532 6644 16584
rect 6696 16572 6702 16584
rect 7469 16575 7527 16581
rect 7469 16572 7481 16575
rect 6696 16544 7481 16572
rect 6696 16532 6702 16544
rect 7469 16541 7481 16544
rect 7515 16541 7527 16575
rect 7469 16535 7527 16541
rect 6564 16504 6592 16532
rect 7484 16504 7512 16535
rect 9030 16532 9036 16584
rect 9088 16572 9094 16584
rect 10152 16572 10180 16612
rect 10229 16609 10241 16612
rect 10275 16609 10287 16643
rect 10229 16603 10287 16609
rect 10318 16600 10324 16652
rect 10376 16600 10382 16652
rect 11054 16600 11060 16652
rect 11112 16640 11118 16652
rect 12078 16643 12136 16649
rect 12078 16640 12090 16643
rect 11112 16612 12090 16640
rect 11112 16600 11118 16612
rect 12078 16609 12090 16612
rect 12124 16609 12136 16643
rect 12078 16603 12136 16609
rect 12345 16643 12403 16649
rect 12345 16609 12357 16643
rect 12391 16640 12403 16643
rect 12434 16640 12440 16652
rect 12391 16612 12440 16640
rect 12391 16609 12403 16612
rect 12345 16603 12403 16609
rect 12434 16600 12440 16612
rect 12492 16600 12498 16652
rect 12618 16600 12624 16652
rect 12676 16640 12682 16652
rect 13832 16649 13860 16680
rect 14016 16680 15332 16708
rect 13081 16643 13139 16649
rect 13081 16640 13093 16643
rect 12676 16612 13093 16640
rect 12676 16600 12682 16612
rect 13081 16609 13093 16612
rect 13127 16640 13139 16643
rect 13817 16643 13875 16649
rect 13127 16612 13784 16640
rect 13127 16609 13139 16612
rect 13081 16603 13139 16609
rect 9088 16544 10180 16572
rect 13756 16572 13784 16612
rect 13817 16609 13829 16643
rect 13863 16609 13875 16643
rect 14016 16640 14044 16680
rect 14090 16649 14096 16652
rect 13817 16603 13875 16609
rect 13924 16612 14044 16640
rect 13924 16572 13952 16612
rect 14084 16603 14096 16649
rect 14090 16600 14096 16603
rect 14148 16600 14154 16652
rect 13756 16544 13952 16572
rect 9088 16532 9094 16544
rect 10594 16504 10600 16516
rect 6564 16476 7420 16504
rect 7484 16476 10600 16504
rect 4488 16408 4660 16436
rect 4488 16396 4494 16408
rect 6454 16396 6460 16448
rect 6512 16436 6518 16448
rect 6641 16439 6699 16445
rect 6641 16436 6653 16439
rect 6512 16408 6653 16436
rect 6512 16396 6518 16408
rect 6641 16405 6653 16408
rect 6687 16405 6699 16439
rect 7392 16436 7420 16476
rect 10594 16464 10600 16476
rect 10652 16464 10658 16516
rect 15304 16504 15332 16680
rect 15396 16652 15424 16748
rect 15930 16736 15936 16788
rect 15988 16736 15994 16788
rect 16301 16779 16359 16785
rect 16301 16745 16313 16779
rect 16347 16776 16359 16779
rect 16482 16776 16488 16788
rect 16347 16748 16488 16776
rect 16347 16745 16359 16748
rect 16301 16739 16359 16745
rect 16482 16736 16488 16748
rect 16540 16736 16546 16788
rect 16577 16779 16635 16785
rect 16577 16745 16589 16779
rect 16623 16776 16635 16779
rect 17678 16776 17684 16788
rect 16623 16748 17684 16776
rect 16623 16745 16635 16748
rect 16577 16739 16635 16745
rect 15378 16600 15384 16652
rect 15436 16640 15442 16652
rect 15473 16643 15531 16649
rect 15473 16640 15485 16643
rect 15436 16612 15485 16640
rect 15436 16600 15442 16612
rect 15473 16609 15485 16612
rect 15519 16609 15531 16643
rect 15473 16603 15531 16609
rect 15657 16643 15715 16649
rect 15657 16609 15669 16643
rect 15703 16640 15715 16643
rect 15948 16640 15976 16736
rect 16117 16643 16175 16649
rect 16117 16640 16129 16643
rect 15703 16612 15884 16640
rect 15948 16612 16129 16640
rect 15703 16609 15715 16612
rect 15657 16603 15715 16609
rect 15856 16572 15884 16612
rect 16117 16609 16129 16612
rect 16163 16609 16175 16643
rect 16592 16640 16620 16739
rect 16868 16652 16896 16748
rect 17678 16736 17684 16748
rect 17736 16736 17742 16788
rect 17862 16736 17868 16788
rect 17920 16776 17926 16788
rect 18509 16779 18567 16785
rect 18509 16776 18521 16779
rect 17920 16748 18521 16776
rect 17920 16736 17926 16748
rect 18509 16745 18521 16748
rect 18555 16745 18567 16779
rect 18509 16739 18567 16745
rect 18874 16736 18880 16788
rect 18932 16736 18938 16788
rect 18966 16736 18972 16788
rect 19024 16736 19030 16788
rect 19058 16736 19064 16788
rect 19116 16736 19122 16788
rect 19429 16779 19487 16785
rect 19429 16745 19441 16779
rect 19475 16776 19487 16779
rect 19610 16776 19616 16788
rect 19475 16748 19616 16776
rect 19475 16745 19487 16748
rect 19429 16739 19487 16745
rect 19610 16736 19616 16748
rect 19668 16736 19674 16788
rect 20346 16736 20352 16788
rect 20404 16776 20410 16788
rect 20533 16779 20591 16785
rect 20533 16776 20545 16779
rect 20404 16748 20545 16776
rect 20404 16736 20410 16748
rect 20533 16745 20545 16748
rect 20579 16745 20591 16779
rect 20533 16739 20591 16745
rect 21269 16779 21327 16785
rect 21269 16745 21281 16779
rect 21315 16745 21327 16779
rect 21269 16739 21327 16745
rect 18892 16708 18920 16736
rect 17052 16680 18920 16708
rect 18984 16708 19012 16736
rect 19521 16711 19579 16717
rect 19521 16708 19533 16711
rect 18984 16680 19533 16708
rect 16117 16603 16175 16609
rect 16224 16612 16620 16640
rect 16761 16643 16819 16649
rect 16224 16572 16252 16612
rect 16761 16609 16773 16643
rect 16807 16609 16819 16643
rect 16761 16603 16819 16609
rect 15856 16544 16252 16572
rect 16776 16572 16804 16603
rect 16850 16600 16856 16652
rect 16908 16600 16914 16652
rect 17052 16649 17080 16680
rect 19521 16677 19533 16680
rect 19567 16677 19579 16711
rect 19521 16671 19579 16677
rect 17037 16643 17095 16649
rect 17037 16609 17049 16643
rect 17083 16609 17095 16643
rect 17037 16603 17095 16609
rect 17126 16600 17132 16652
rect 17184 16600 17190 16652
rect 17304 16643 17362 16649
rect 17304 16609 17316 16643
rect 17350 16640 17362 16643
rect 17586 16640 17592 16652
rect 17350 16612 17592 16640
rect 17350 16609 17362 16612
rect 17304 16603 17362 16609
rect 17586 16600 17592 16612
rect 17644 16600 17650 16652
rect 17678 16600 17684 16652
rect 17736 16640 17742 16652
rect 18693 16643 18751 16649
rect 17736 16612 18644 16640
rect 17736 16600 17742 16612
rect 17144 16572 17172 16600
rect 16776 16544 17172 16572
rect 18616 16572 18644 16612
rect 18693 16609 18705 16643
rect 18739 16640 18751 16643
rect 19426 16640 19432 16652
rect 18739 16612 19432 16640
rect 18739 16609 18751 16612
rect 18693 16603 18751 16609
rect 18877 16575 18935 16581
rect 18877 16572 18889 16575
rect 18616 16544 18889 16572
rect 16776 16504 16804 16544
rect 18877 16541 18889 16544
rect 18923 16541 18935 16575
rect 18877 16535 18935 16541
rect 15304 16476 16804 16504
rect 18417 16507 18475 16513
rect 18417 16473 18429 16507
rect 18463 16504 18475 16507
rect 18984 16504 19012 16612
rect 19426 16600 19432 16612
rect 19484 16600 19490 16652
rect 20717 16643 20775 16649
rect 20717 16609 20729 16643
rect 20763 16640 20775 16643
rect 21284 16640 21312 16739
rect 21634 16736 21640 16788
rect 21692 16736 21698 16788
rect 21729 16779 21787 16785
rect 21729 16745 21741 16779
rect 21775 16776 21787 16779
rect 22002 16776 22008 16788
rect 21775 16748 22008 16776
rect 21775 16745 21787 16748
rect 21729 16739 21787 16745
rect 22002 16736 22008 16748
rect 22060 16736 22066 16788
rect 22094 16736 22100 16788
rect 22152 16736 22158 16788
rect 22370 16736 22376 16788
rect 22428 16736 22434 16788
rect 22554 16736 22560 16788
rect 22612 16776 22618 16788
rect 22612 16748 22968 16776
rect 22612 16736 22618 16748
rect 22112 16708 22140 16736
rect 22388 16708 22416 16736
rect 22940 16717 22968 16748
rect 23014 16736 23020 16788
rect 23072 16776 23078 16788
rect 24213 16779 24271 16785
rect 23072 16748 24164 16776
rect 23072 16736 23078 16748
rect 22925 16711 22983 16717
rect 22112 16680 22324 16708
rect 22388 16680 22600 16708
rect 20763 16612 21312 16640
rect 20763 16609 20775 16612
rect 20717 16603 20775 16609
rect 21358 16600 21364 16652
rect 21416 16640 21422 16652
rect 22296 16640 22324 16680
rect 22572 16649 22600 16680
rect 22925 16677 22937 16711
rect 22971 16708 22983 16711
rect 22971 16680 23152 16708
rect 22971 16677 22983 16680
rect 22925 16671 22983 16677
rect 22465 16643 22523 16649
rect 22465 16640 22477 16643
rect 21416 16612 22232 16640
rect 22296 16612 22477 16640
rect 21416 16600 21422 16612
rect 19702 16532 19708 16584
rect 19760 16572 19766 16584
rect 21821 16575 21879 16581
rect 21821 16572 21833 16575
rect 19760 16544 21833 16572
rect 19760 16532 19766 16544
rect 21821 16541 21833 16544
rect 21867 16541 21879 16575
rect 22204 16572 22232 16612
rect 22465 16609 22477 16612
rect 22511 16609 22523 16643
rect 22465 16603 22523 16609
rect 22557 16643 22615 16649
rect 22557 16609 22569 16643
rect 22603 16609 22615 16643
rect 22557 16603 22615 16609
rect 23014 16600 23020 16652
rect 23072 16600 23078 16652
rect 23124 16649 23152 16680
rect 23750 16668 23756 16720
rect 23808 16708 23814 16720
rect 24136 16708 24164 16748
rect 24213 16745 24225 16779
rect 24259 16776 24271 16779
rect 24302 16776 24308 16788
rect 24259 16748 24308 16776
rect 24259 16745 24271 16748
rect 24213 16739 24271 16745
rect 24302 16736 24308 16748
rect 24360 16736 24366 16788
rect 24673 16779 24731 16785
rect 24673 16745 24685 16779
rect 24719 16776 24731 16779
rect 24762 16776 24768 16788
rect 24719 16748 24768 16776
rect 24719 16745 24731 16748
rect 24673 16739 24731 16745
rect 24762 16736 24768 16748
rect 24820 16736 24826 16788
rect 24857 16779 24915 16785
rect 24857 16745 24869 16779
rect 24903 16745 24915 16779
rect 24857 16739 24915 16745
rect 24872 16708 24900 16739
rect 24946 16736 24952 16788
rect 25004 16776 25010 16788
rect 25041 16779 25099 16785
rect 25041 16776 25053 16779
rect 25004 16748 25053 16776
rect 25004 16736 25010 16748
rect 25041 16745 25053 16748
rect 25087 16745 25099 16779
rect 25041 16739 25099 16745
rect 25130 16736 25136 16788
rect 25188 16776 25194 16788
rect 25501 16779 25559 16785
rect 25188 16748 25452 16776
rect 25188 16736 25194 16748
rect 23808 16680 24072 16708
rect 24136 16680 24256 16708
rect 24872 16680 25360 16708
rect 23808 16668 23814 16680
rect 24044 16649 24072 16680
rect 23109 16643 23167 16649
rect 23109 16609 23121 16643
rect 23155 16609 23167 16643
rect 23109 16603 23167 16609
rect 24029 16643 24087 16649
rect 24029 16609 24041 16643
rect 24075 16609 24087 16643
rect 24029 16603 24087 16609
rect 24118 16600 24124 16652
rect 24176 16600 24182 16652
rect 24228 16649 24256 16680
rect 24213 16643 24271 16649
rect 24213 16609 24225 16643
rect 24259 16640 24271 16643
rect 24946 16640 24952 16652
rect 24259 16612 24952 16640
rect 24259 16609 24271 16612
rect 24213 16603 24271 16609
rect 24946 16600 24952 16612
rect 25004 16600 25010 16652
rect 25038 16600 25044 16652
rect 25096 16640 25102 16652
rect 25332 16649 25360 16680
rect 25133 16643 25191 16649
rect 25133 16640 25145 16643
rect 25096 16612 25145 16640
rect 25096 16600 25102 16612
rect 25133 16609 25145 16612
rect 25179 16609 25191 16643
rect 25133 16603 25191 16609
rect 25317 16643 25375 16649
rect 25317 16609 25329 16643
rect 25363 16609 25375 16643
rect 25424 16640 25452 16748
rect 25501 16745 25513 16779
rect 25547 16745 25559 16779
rect 25501 16739 25559 16745
rect 25516 16708 25544 16739
rect 25774 16736 25780 16788
rect 25832 16736 25838 16788
rect 26234 16708 26240 16720
rect 25516 16680 26240 16708
rect 26234 16668 26240 16680
rect 26292 16668 26298 16720
rect 25593 16643 25651 16649
rect 25593 16640 25605 16643
rect 25424 16612 25605 16640
rect 25317 16603 25375 16609
rect 25593 16609 25605 16612
rect 25639 16609 25651 16643
rect 25593 16603 25651 16609
rect 24136 16572 24164 16600
rect 24302 16572 24308 16584
rect 22204 16544 23520 16572
rect 24136 16544 24308 16572
rect 21821 16535 21879 16541
rect 23014 16504 23020 16516
rect 18463 16476 19012 16504
rect 22848 16476 23020 16504
rect 18463 16473 18475 16476
rect 18417 16467 18475 16473
rect 7558 16436 7564 16448
rect 7392 16408 7564 16436
rect 6641 16399 6699 16405
rect 7558 16396 7564 16408
rect 7616 16396 7622 16448
rect 7745 16439 7803 16445
rect 7745 16405 7757 16439
rect 7791 16436 7803 16439
rect 8294 16436 8300 16448
rect 7791 16408 8300 16436
rect 7791 16405 7803 16408
rect 7745 16399 7803 16405
rect 8294 16396 8300 16408
rect 8352 16436 8358 16448
rect 9309 16439 9367 16445
rect 9309 16436 9321 16439
rect 8352 16408 9321 16436
rect 8352 16396 8358 16408
rect 9309 16405 9321 16408
rect 9355 16405 9367 16439
rect 9309 16399 9367 16405
rect 9493 16439 9551 16445
rect 9493 16405 9505 16439
rect 9539 16436 9551 16439
rect 10870 16436 10876 16448
rect 9539 16408 10876 16436
rect 9539 16405 9551 16408
rect 9493 16399 9551 16405
rect 10870 16396 10876 16408
rect 10928 16396 10934 16448
rect 11238 16396 11244 16448
rect 11296 16436 11302 16448
rect 13722 16436 13728 16448
rect 11296 16408 13728 16436
rect 11296 16396 11302 16408
rect 13722 16396 13728 16408
rect 13780 16396 13786 16448
rect 15286 16396 15292 16448
rect 15344 16396 15350 16448
rect 22281 16439 22339 16445
rect 22281 16405 22293 16439
rect 22327 16436 22339 16439
rect 22370 16436 22376 16448
rect 22327 16408 22376 16436
rect 22327 16405 22339 16408
rect 22281 16399 22339 16405
rect 22370 16396 22376 16408
rect 22428 16396 22434 16448
rect 22848 16445 22876 16476
rect 23014 16464 23020 16476
rect 23072 16504 23078 16516
rect 23492 16504 23520 16544
rect 24302 16532 24308 16544
rect 24360 16532 24366 16584
rect 24578 16532 24584 16584
rect 24636 16532 24642 16584
rect 24596 16504 24624 16532
rect 23072 16476 23336 16504
rect 23492 16476 24624 16504
rect 24688 16476 25268 16504
rect 23072 16464 23078 16476
rect 23308 16448 23336 16476
rect 22833 16439 22891 16445
rect 22833 16405 22845 16439
rect 22879 16405 22891 16439
rect 22833 16399 22891 16405
rect 23106 16396 23112 16448
rect 23164 16396 23170 16448
rect 23290 16396 23296 16448
rect 23348 16396 23354 16448
rect 23382 16396 23388 16448
rect 23440 16396 23446 16448
rect 24688 16445 24716 16476
rect 25240 16448 25268 16476
rect 24673 16439 24731 16445
rect 24673 16405 24685 16439
rect 24719 16405 24731 16439
rect 24673 16399 24731 16405
rect 25222 16396 25228 16448
rect 25280 16396 25286 16448
rect 552 16346 27416 16368
rect 552 16294 3756 16346
rect 3808 16294 3820 16346
rect 3872 16294 3884 16346
rect 3936 16294 3948 16346
rect 4000 16294 4012 16346
rect 4064 16294 10472 16346
rect 10524 16294 10536 16346
rect 10588 16294 10600 16346
rect 10652 16294 10664 16346
rect 10716 16294 10728 16346
rect 10780 16294 17188 16346
rect 17240 16294 17252 16346
rect 17304 16294 17316 16346
rect 17368 16294 17380 16346
rect 17432 16294 17444 16346
rect 17496 16294 23904 16346
rect 23956 16294 23968 16346
rect 24020 16294 24032 16346
rect 24084 16294 24096 16346
rect 24148 16294 24160 16346
rect 24212 16294 27416 16346
rect 552 16272 27416 16294
rect 2682 16192 2688 16244
rect 2740 16192 2746 16244
rect 5905 16235 5963 16241
rect 5905 16201 5917 16235
rect 5951 16232 5963 16235
rect 6178 16232 6184 16244
rect 5951 16204 6184 16232
rect 5951 16201 5963 16204
rect 5905 16195 5963 16201
rect 6178 16192 6184 16204
rect 6236 16192 6242 16244
rect 8846 16192 8852 16244
rect 8904 16192 8910 16244
rect 9398 16192 9404 16244
rect 9456 16192 9462 16244
rect 11054 16192 11060 16244
rect 11112 16192 11118 16244
rect 11146 16192 11152 16244
rect 11204 16232 11210 16244
rect 11422 16232 11428 16244
rect 11204 16204 11428 16232
rect 11204 16192 11210 16204
rect 11422 16192 11428 16204
rect 11480 16232 11486 16244
rect 12161 16235 12219 16241
rect 12161 16232 12173 16235
rect 11480 16204 12173 16232
rect 11480 16192 11486 16204
rect 12161 16201 12173 16204
rect 12207 16201 12219 16235
rect 12161 16195 12219 16201
rect 14090 16192 14096 16244
rect 14148 16232 14154 16244
rect 14277 16235 14335 16241
rect 14277 16232 14289 16235
rect 14148 16204 14289 16232
rect 14148 16192 14154 16204
rect 14277 16201 14289 16204
rect 14323 16201 14335 16235
rect 15562 16232 15568 16244
rect 14277 16195 14335 16201
rect 15304 16204 15568 16232
rect 7377 16167 7435 16173
rect 7377 16133 7389 16167
rect 7423 16133 7435 16167
rect 9416 16164 9444 16192
rect 11330 16164 11336 16176
rect 9416 16136 11336 16164
rect 7377 16127 7435 16133
rect 2590 16096 2596 16108
rect 2056 16068 2596 16096
rect 2056 16037 2084 16068
rect 2590 16056 2596 16068
rect 2648 16096 2654 16108
rect 7392 16096 7420 16127
rect 11330 16124 11336 16136
rect 11388 16164 11394 16176
rect 12894 16164 12900 16176
rect 11388 16136 12900 16164
rect 11388 16124 11394 16136
rect 12894 16124 12900 16136
rect 12952 16124 12958 16176
rect 8021 16099 8079 16105
rect 8021 16096 8033 16099
rect 2648 16068 3464 16096
rect 7392 16068 8033 16096
rect 2648 16056 2654 16068
rect 2041 16031 2099 16037
rect 2041 15997 2053 16031
rect 2087 15997 2099 16031
rect 2041 15991 2099 15997
rect 2130 15988 2136 16040
rect 2188 15988 2194 16040
rect 2225 16031 2283 16037
rect 2225 15997 2237 16031
rect 2271 15997 2283 16031
rect 2225 15991 2283 15997
rect 1670 15920 1676 15972
rect 1728 15960 1734 15972
rect 1728 15932 1900 15960
rect 1728 15920 1734 15932
rect 1762 15852 1768 15904
rect 1820 15852 1826 15904
rect 1872 15892 1900 15932
rect 1946 15920 1952 15972
rect 2004 15960 2010 15972
rect 2240 15960 2268 15991
rect 2406 15988 2412 16040
rect 2464 15988 2470 16040
rect 2501 16031 2559 16037
rect 2501 15997 2513 16031
rect 2547 15997 2559 16031
rect 2501 15991 2559 15997
rect 2004 15932 2268 15960
rect 2004 15920 2010 15932
rect 2314 15920 2320 15972
rect 2372 15960 2378 15972
rect 2516 15960 2544 15991
rect 2866 15988 2872 16040
rect 2924 15988 2930 16040
rect 2958 15988 2964 16040
rect 3016 15988 3022 16040
rect 3436 16037 3464 16068
rect 8021 16065 8033 16068
rect 8067 16065 8079 16099
rect 8021 16059 8079 16065
rect 8202 16056 8208 16108
rect 8260 16096 8266 16108
rect 9030 16096 9036 16108
rect 8260 16068 9036 16096
rect 8260 16056 8266 16068
rect 9030 16056 9036 16068
rect 9088 16056 9094 16108
rect 10152 16068 14872 16096
rect 3421 16031 3479 16037
rect 3421 15997 3433 16031
rect 3467 15997 3479 16031
rect 3421 15991 3479 15997
rect 4430 15988 4436 16040
rect 4488 16028 4494 16040
rect 4525 16031 4583 16037
rect 4525 16028 4537 16031
rect 4488 16000 4537 16028
rect 4488 15988 4494 16000
rect 4525 15997 4537 16000
rect 4571 16028 4583 16031
rect 5997 16031 6055 16037
rect 5997 16028 6009 16031
rect 4571 16000 6009 16028
rect 4571 15997 4583 16000
rect 4525 15991 4583 15997
rect 5997 15997 6009 16000
rect 6043 15997 6055 16031
rect 5997 15991 6055 15997
rect 6086 15988 6092 16040
rect 6144 16028 6150 16040
rect 10152 16037 10180 16068
rect 10137 16031 10195 16037
rect 6144 16000 7604 16028
rect 6144 15988 6150 16000
rect 2372 15932 2544 15960
rect 2746 15932 3280 15960
rect 2372 15920 2378 15932
rect 2746 15892 2774 15932
rect 3252 15901 3280 15932
rect 3326 15920 3332 15972
rect 3384 15960 3390 15972
rect 3605 15963 3663 15969
rect 3605 15960 3617 15963
rect 3384 15932 3617 15960
rect 3384 15920 3390 15932
rect 3605 15929 3617 15932
rect 3651 15929 3663 15963
rect 3605 15923 3663 15929
rect 4792 15963 4850 15969
rect 4792 15929 4804 15963
rect 4838 15960 4850 15963
rect 6264 15963 6322 15969
rect 4838 15932 6040 15960
rect 4838 15929 4850 15932
rect 4792 15923 4850 15929
rect 1872 15864 2774 15892
rect 3237 15895 3295 15901
rect 3237 15861 3249 15895
rect 3283 15861 3295 15895
rect 6012 15892 6040 15932
rect 6264 15929 6276 15963
rect 6310 15960 6322 15963
rect 6546 15960 6552 15972
rect 6310 15932 6552 15960
rect 6310 15929 6322 15932
rect 6264 15923 6322 15929
rect 6546 15920 6552 15932
rect 6604 15920 6610 15972
rect 6454 15892 6460 15904
rect 6012 15864 6460 15892
rect 3237 15855 3295 15861
rect 6454 15852 6460 15864
rect 6512 15852 6518 15904
rect 7466 15852 7472 15904
rect 7524 15852 7530 15904
rect 7576 15892 7604 16000
rect 10137 15997 10149 16031
rect 10183 15997 10195 16031
rect 10137 15991 10195 15997
rect 10965 16031 11023 16037
rect 10965 15997 10977 16031
rect 11011 16028 11023 16031
rect 11011 16000 11192 16028
rect 11011 15997 11023 16000
rect 10965 15991 11023 15997
rect 7650 15920 7656 15972
rect 7708 15960 7714 15972
rect 9950 15960 9956 15972
rect 7708 15932 9956 15960
rect 7708 15920 7714 15932
rect 9950 15920 9956 15932
rect 10008 15960 10014 15972
rect 10686 15960 10692 15972
rect 10008 15932 10692 15960
rect 10008 15920 10014 15932
rect 10686 15920 10692 15932
rect 10744 15920 10750 15972
rect 11054 15920 11060 15972
rect 11112 15920 11118 15972
rect 11072 15892 11100 15920
rect 7576 15864 11100 15892
rect 11164 15892 11192 16000
rect 11238 15988 11244 16040
rect 11296 15988 11302 16040
rect 11330 15988 11336 16040
rect 11388 15988 11394 16040
rect 11609 16031 11667 16037
rect 11609 15997 11621 16031
rect 11655 16028 11667 16031
rect 11882 16028 11888 16040
rect 11655 16000 11888 16028
rect 11655 15997 11667 16000
rect 11609 15991 11667 15997
rect 11882 15988 11888 16000
rect 11940 15988 11946 16040
rect 13446 16028 13452 16040
rect 11992 16000 13452 16028
rect 11425 15963 11483 15969
rect 11425 15929 11437 15963
rect 11471 15960 11483 15963
rect 11992 15960 12020 16000
rect 13446 15988 13452 16000
rect 13504 15988 13510 16040
rect 14461 16031 14519 16037
rect 14461 15997 14473 16031
rect 14507 16028 14519 16031
rect 14507 16000 14688 16028
rect 14507 15997 14519 16000
rect 14461 15991 14519 15997
rect 11471 15932 12020 15960
rect 12069 15963 12127 15969
rect 11471 15929 11483 15932
rect 11425 15923 11483 15929
rect 12069 15929 12081 15963
rect 12115 15929 12127 15963
rect 12069 15923 12127 15929
rect 11698 15892 11704 15904
rect 11164 15864 11704 15892
rect 11698 15852 11704 15864
rect 11756 15892 11762 15904
rect 12084 15892 12112 15923
rect 14660 15901 14688 16000
rect 14844 15972 14872 16068
rect 14918 16056 14924 16108
rect 14976 16096 14982 16108
rect 15105 16099 15163 16105
rect 15105 16096 15117 16099
rect 14976 16068 15117 16096
rect 14976 16056 14982 16068
rect 15105 16065 15117 16068
rect 15151 16065 15163 16099
rect 15105 16059 15163 16065
rect 15197 16099 15255 16105
rect 15197 16065 15209 16099
rect 15243 16096 15255 16099
rect 15304 16096 15332 16204
rect 15562 16192 15568 16204
rect 15620 16232 15626 16244
rect 16482 16232 16488 16244
rect 15620 16204 16488 16232
rect 15620 16192 15626 16204
rect 16482 16192 16488 16204
rect 16540 16192 16546 16244
rect 19702 16232 19708 16244
rect 16592 16204 19708 16232
rect 16592 16164 16620 16204
rect 19702 16192 19708 16204
rect 19760 16192 19766 16244
rect 19978 16192 19984 16244
rect 20036 16192 20042 16244
rect 25314 16192 25320 16244
rect 25372 16232 25378 16244
rect 25409 16235 25467 16241
rect 25409 16232 25421 16235
rect 25372 16204 25421 16232
rect 25372 16192 25378 16204
rect 25409 16201 25421 16204
rect 25455 16201 25467 16235
rect 25409 16195 25467 16201
rect 20717 16167 20775 16173
rect 20717 16164 20729 16167
rect 15243 16068 15332 16096
rect 15488 16136 16620 16164
rect 18432 16136 20729 16164
rect 15243 16065 15255 16068
rect 15197 16059 15255 16065
rect 15488 16040 15516 16136
rect 15746 16056 15752 16108
rect 15804 16056 15810 16108
rect 18432 16040 18460 16136
rect 20717 16133 20729 16136
rect 20763 16133 20775 16167
rect 20717 16127 20775 16133
rect 15013 16031 15071 16037
rect 15013 15997 15025 16031
rect 15059 16028 15071 16031
rect 15286 16028 15292 16040
rect 15059 16000 15292 16028
rect 15059 15997 15071 16000
rect 15013 15991 15071 15997
rect 15286 15988 15292 16000
rect 15344 15988 15350 16040
rect 15470 15988 15476 16040
rect 15528 15988 15534 16040
rect 15841 16031 15899 16037
rect 15841 15997 15853 16031
rect 15887 16028 15899 16031
rect 16117 16031 16175 16037
rect 16117 16028 16129 16031
rect 15887 16000 16129 16028
rect 15887 15997 15899 16000
rect 15841 15991 15899 15997
rect 16117 15997 16129 16000
rect 16163 15997 16175 16031
rect 16117 15991 16175 15997
rect 16206 15988 16212 16040
rect 16264 16028 16270 16040
rect 16669 16031 16727 16037
rect 16669 16028 16681 16031
rect 16264 16000 16681 16028
rect 16264 15988 16270 16000
rect 16669 15997 16681 16000
rect 16715 15997 16727 16031
rect 16669 15991 16727 15997
rect 17497 16031 17555 16037
rect 17497 15997 17509 16031
rect 17543 16028 17555 16031
rect 17770 16028 17776 16040
rect 17543 16000 17776 16028
rect 17543 15997 17555 16000
rect 17497 15991 17555 15997
rect 17770 15988 17776 16000
rect 17828 15988 17834 16040
rect 18322 15988 18328 16040
rect 18380 15988 18386 16040
rect 18414 15988 18420 16040
rect 18472 15988 18478 16040
rect 20438 15988 20444 16040
rect 20496 16028 20502 16040
rect 20533 16031 20591 16037
rect 20533 16028 20545 16031
rect 20496 16000 20545 16028
rect 20496 15988 20502 16000
rect 20533 15997 20545 16000
rect 20579 15997 20591 16031
rect 20533 15991 20591 15997
rect 20901 16031 20959 16037
rect 20901 15997 20913 16031
rect 20947 15997 20959 16031
rect 20901 15991 20959 15997
rect 14826 15920 14832 15972
rect 14884 15960 14890 15972
rect 18693 15963 18751 15969
rect 18693 15960 18705 15963
rect 14884 15932 18705 15960
rect 14884 15920 14890 15932
rect 18693 15929 18705 15932
rect 18739 15929 18751 15963
rect 18693 15923 18751 15929
rect 18782 15920 18788 15972
rect 18840 15960 18846 15972
rect 20916 15960 20944 15991
rect 21082 15988 21088 16040
rect 21140 15988 21146 16040
rect 22646 15988 22652 16040
rect 22704 16028 22710 16040
rect 23750 16028 23756 16040
rect 22704 16000 23756 16028
rect 22704 15988 22710 16000
rect 23750 15988 23756 16000
rect 23808 15988 23814 16040
rect 24118 15988 24124 16040
rect 24176 16028 24182 16040
rect 24762 16028 24768 16040
rect 24176 16000 24768 16028
rect 24176 15988 24182 16000
rect 24762 15988 24768 16000
rect 24820 15988 24826 16040
rect 26234 15988 26240 16040
rect 26292 16028 26298 16040
rect 26522 16031 26580 16037
rect 26522 16028 26534 16031
rect 26292 16000 26534 16028
rect 26292 15988 26298 16000
rect 26522 15997 26534 16000
rect 26568 15997 26580 16031
rect 26522 15991 26580 15997
rect 26789 16031 26847 16037
rect 26789 15997 26801 16031
rect 26835 16028 26847 16031
rect 26878 16028 26884 16040
rect 26835 16000 26884 16028
rect 26835 15997 26847 16000
rect 26789 15991 26847 15997
rect 26878 15988 26884 16000
rect 26936 15988 26942 16040
rect 18840 15932 21496 15960
rect 18840 15920 18846 15932
rect 21468 15904 21496 15932
rect 11756 15864 12112 15892
rect 14645 15895 14703 15901
rect 11756 15852 11762 15864
rect 14645 15861 14657 15895
rect 14691 15861 14703 15895
rect 14645 15855 14703 15861
rect 15470 15852 15476 15904
rect 15528 15852 15534 15904
rect 17678 15852 17684 15904
rect 17736 15852 17742 15904
rect 17954 15852 17960 15904
rect 18012 15892 18018 15904
rect 18141 15895 18199 15901
rect 18141 15892 18153 15895
rect 18012 15864 18153 15892
rect 18012 15852 18018 15864
rect 18141 15861 18153 15864
rect 18187 15861 18199 15895
rect 18141 15855 18199 15861
rect 20898 15852 20904 15904
rect 20956 15852 20962 15904
rect 21450 15852 21456 15904
rect 21508 15852 21514 15904
rect 23566 15852 23572 15904
rect 23624 15892 23630 15904
rect 24213 15895 24271 15901
rect 24213 15892 24225 15895
rect 23624 15864 24225 15892
rect 23624 15852 23630 15864
rect 24213 15861 24225 15864
rect 24259 15892 24271 15895
rect 24670 15892 24676 15904
rect 24259 15864 24676 15892
rect 24259 15861 24271 15864
rect 24213 15855 24271 15861
rect 24670 15852 24676 15864
rect 24728 15852 24734 15904
rect 552 15802 27576 15824
rect 552 15750 7114 15802
rect 7166 15750 7178 15802
rect 7230 15750 7242 15802
rect 7294 15750 7306 15802
rect 7358 15750 7370 15802
rect 7422 15750 13830 15802
rect 13882 15750 13894 15802
rect 13946 15750 13958 15802
rect 14010 15750 14022 15802
rect 14074 15750 14086 15802
rect 14138 15750 20546 15802
rect 20598 15750 20610 15802
rect 20662 15750 20674 15802
rect 20726 15750 20738 15802
rect 20790 15750 20802 15802
rect 20854 15750 27262 15802
rect 27314 15750 27326 15802
rect 27378 15750 27390 15802
rect 27442 15750 27454 15802
rect 27506 15750 27518 15802
rect 27570 15750 27576 15802
rect 552 15728 27576 15750
rect 1670 15648 1676 15700
rect 1728 15648 1734 15700
rect 1762 15648 1768 15700
rect 1820 15648 1826 15700
rect 2501 15691 2559 15697
rect 2501 15657 2513 15691
rect 2547 15688 2559 15691
rect 2590 15688 2596 15700
rect 2547 15660 2596 15688
rect 2547 15657 2559 15660
rect 2501 15651 2559 15657
rect 2590 15648 2596 15660
rect 2648 15648 2654 15700
rect 6733 15691 6791 15697
rect 6733 15657 6745 15691
rect 6779 15688 6791 15691
rect 6822 15688 6828 15700
rect 6779 15660 6828 15688
rect 6779 15657 6791 15660
rect 6733 15651 6791 15657
rect 6822 15648 6828 15660
rect 6880 15648 6886 15700
rect 7466 15648 7472 15700
rect 7524 15648 7530 15700
rect 7558 15648 7564 15700
rect 7616 15688 7622 15700
rect 8478 15688 8484 15700
rect 7616 15660 8484 15688
rect 7616 15648 7622 15660
rect 1688 15620 1716 15648
rect 1412 15592 1716 15620
rect 934 15512 940 15564
rect 992 15552 998 15564
rect 1412 15561 1440 15592
rect 1780 15561 1808 15648
rect 4430 15620 4436 15632
rect 3252 15592 4436 15620
rect 1213 15555 1271 15561
rect 1213 15552 1225 15555
rect 992 15524 1225 15552
rect 992 15512 998 15524
rect 1213 15521 1225 15524
rect 1259 15521 1271 15555
rect 1213 15515 1271 15521
rect 1305 15555 1363 15561
rect 1305 15521 1317 15555
rect 1351 15521 1363 15555
rect 1305 15515 1363 15521
rect 1397 15555 1455 15561
rect 1397 15521 1409 15555
rect 1443 15521 1455 15555
rect 1397 15515 1455 15521
rect 1581 15555 1639 15561
rect 1581 15521 1593 15555
rect 1627 15521 1639 15555
rect 1581 15515 1639 15521
rect 1765 15555 1823 15561
rect 1765 15521 1777 15555
rect 1811 15521 1823 15555
rect 1765 15515 1823 15521
rect 1320 15416 1348 15515
rect 1596 15484 1624 15515
rect 2406 15512 2412 15564
rect 2464 15512 2470 15564
rect 2424 15484 2452 15512
rect 1596 15456 2452 15484
rect 3142 15444 3148 15496
rect 3200 15444 3206 15496
rect 3252 15493 3280 15592
rect 4430 15580 4436 15592
rect 4488 15580 4494 15632
rect 7484 15620 7512 15648
rect 7852 15629 7880 15660
rect 8478 15648 8484 15660
rect 8536 15648 8542 15700
rect 9030 15648 9036 15700
rect 9088 15648 9094 15700
rect 10505 15691 10563 15697
rect 10505 15657 10517 15691
rect 10551 15657 10563 15691
rect 10505 15651 10563 15657
rect 5644 15592 7512 15620
rect 7837 15623 7895 15629
rect 3510 15561 3516 15564
rect 3504 15515 3516 15561
rect 3510 15512 3516 15515
rect 3568 15512 3574 15564
rect 4246 15512 4252 15564
rect 4304 15552 4310 15564
rect 5644 15561 5672 15592
rect 5629 15555 5687 15561
rect 4304 15524 5396 15552
rect 4304 15512 4310 15524
rect 3237 15487 3295 15493
rect 3237 15453 3249 15487
rect 3283 15453 3295 15487
rect 3237 15447 3295 15453
rect 5261 15487 5319 15493
rect 5261 15453 5273 15487
rect 5307 15453 5319 15487
rect 5368 15484 5396 15524
rect 5629 15521 5641 15555
rect 5675 15521 5687 15555
rect 5629 15515 5687 15521
rect 5905 15555 5963 15561
rect 5905 15521 5917 15555
rect 5951 15552 5963 15555
rect 6086 15552 6092 15564
rect 5951 15524 6092 15552
rect 5951 15521 5963 15524
rect 5905 15515 5963 15521
rect 5920 15484 5948 15515
rect 6086 15512 6092 15524
rect 6144 15512 6150 15564
rect 6178 15512 6184 15564
rect 6236 15512 6242 15564
rect 6472 15561 6500 15592
rect 7837 15589 7849 15623
rect 7883 15589 7895 15623
rect 7837 15583 7895 15589
rect 8018 15580 8024 15632
rect 8076 15629 8082 15632
rect 8076 15623 8095 15629
rect 8083 15589 8095 15623
rect 8076 15583 8095 15589
rect 10168 15623 10226 15629
rect 10168 15589 10180 15623
rect 10214 15620 10226 15623
rect 10520 15620 10548 15651
rect 10870 15648 10876 15700
rect 10928 15648 10934 15700
rect 15289 15691 15347 15697
rect 15289 15657 15301 15691
rect 15335 15688 15347 15691
rect 15654 15688 15660 15700
rect 15335 15660 15660 15688
rect 15335 15657 15347 15660
rect 15289 15651 15347 15657
rect 15654 15648 15660 15660
rect 15712 15688 15718 15700
rect 15930 15688 15936 15700
rect 15712 15660 15936 15688
rect 15712 15648 15718 15660
rect 15930 15648 15936 15660
rect 15988 15648 15994 15700
rect 16117 15691 16175 15697
rect 16117 15657 16129 15691
rect 16163 15688 16175 15691
rect 16206 15688 16212 15700
rect 16163 15660 16212 15688
rect 16163 15657 16175 15660
rect 16117 15651 16175 15657
rect 16206 15648 16212 15660
rect 16264 15648 16270 15700
rect 17678 15648 17684 15700
rect 17736 15648 17742 15700
rect 18322 15648 18328 15700
rect 18380 15688 18386 15700
rect 18969 15691 19027 15697
rect 18969 15688 18981 15691
rect 18380 15660 18981 15688
rect 18380 15648 18386 15660
rect 18969 15657 18981 15660
rect 19015 15657 19027 15691
rect 18969 15651 19027 15657
rect 20993 15691 21051 15697
rect 20993 15657 21005 15691
rect 21039 15688 21051 15691
rect 21266 15688 21272 15700
rect 21039 15660 21272 15688
rect 21039 15657 21051 15660
rect 20993 15651 21051 15657
rect 10214 15592 10548 15620
rect 10214 15589 10226 15592
rect 10168 15583 10226 15589
rect 8076 15580 8082 15583
rect 6457 15555 6515 15561
rect 6457 15521 6469 15555
rect 6503 15521 6515 15555
rect 6457 15515 6515 15521
rect 6549 15555 6607 15561
rect 6549 15521 6561 15555
rect 6595 15552 6607 15555
rect 6638 15552 6644 15564
rect 6595 15524 6644 15552
rect 6595 15521 6607 15524
rect 6549 15515 6607 15521
rect 6638 15512 6644 15524
rect 6696 15512 6702 15564
rect 6730 15512 6736 15564
rect 6788 15552 6794 15564
rect 6825 15555 6883 15561
rect 6825 15552 6837 15555
rect 6788 15524 6837 15552
rect 6788 15512 6794 15524
rect 6825 15521 6837 15524
rect 6871 15521 6883 15555
rect 6825 15515 6883 15521
rect 7285 15555 7343 15561
rect 7285 15521 7297 15555
rect 7331 15521 7343 15555
rect 7285 15515 7343 15521
rect 7392 15524 8984 15552
rect 5368 15456 5948 15484
rect 6196 15484 6224 15512
rect 7300 15484 7328 15515
rect 6196 15456 7328 15484
rect 5261 15447 5319 15453
rect 2130 15416 2136 15428
rect 1320 15388 2136 15416
rect 2130 15376 2136 15388
rect 2188 15376 2194 15428
rect 3252 15416 3280 15447
rect 2792 15388 3280 15416
rect 4617 15419 4675 15425
rect 2792 15360 2820 15388
rect 4617 15385 4629 15419
rect 4663 15416 4675 15419
rect 5276 15416 5304 15447
rect 4663 15388 5304 15416
rect 4663 15385 4675 15388
rect 4617 15379 4675 15385
rect 937 15351 995 15357
rect 937 15317 949 15351
rect 983 15348 995 15351
rect 1118 15348 1124 15360
rect 983 15320 1124 15348
rect 983 15317 995 15320
rect 937 15311 995 15317
rect 1118 15308 1124 15320
rect 1176 15308 1182 15360
rect 1578 15308 1584 15360
rect 1636 15348 1642 15360
rect 2314 15348 2320 15360
rect 1636 15320 2320 15348
rect 1636 15308 1642 15320
rect 2314 15308 2320 15320
rect 2372 15308 2378 15360
rect 2406 15308 2412 15360
rect 2464 15308 2470 15360
rect 2774 15308 2780 15360
rect 2832 15308 2838 15360
rect 4154 15308 4160 15360
rect 4212 15348 4218 15360
rect 4632 15348 4660 15379
rect 5718 15376 5724 15428
rect 5776 15416 5782 15428
rect 6181 15419 6239 15425
rect 6181 15416 6193 15419
rect 5776 15388 6193 15416
rect 5776 15376 5782 15388
rect 6181 15385 6193 15388
rect 6227 15416 6239 15419
rect 7392 15416 7420 15524
rect 7466 15444 7472 15496
rect 7524 15444 7530 15496
rect 8386 15444 8392 15496
rect 8444 15484 8450 15496
rect 8849 15487 8907 15493
rect 8849 15484 8861 15487
rect 8444 15456 8861 15484
rect 8444 15444 8450 15456
rect 8849 15453 8861 15456
rect 8895 15453 8907 15487
rect 8849 15447 8907 15453
rect 8297 15419 8355 15425
rect 8297 15416 8309 15419
rect 6227 15388 7420 15416
rect 8036 15388 8309 15416
rect 6227 15385 6239 15388
rect 6181 15379 6239 15385
rect 4212 15320 4660 15348
rect 4212 15308 4218 15320
rect 4706 15308 4712 15360
rect 4764 15308 4770 15360
rect 5534 15308 5540 15360
rect 5592 15308 5598 15360
rect 8036 15357 8064 15388
rect 8297 15385 8309 15388
rect 8343 15385 8355 15419
rect 8297 15379 8355 15385
rect 8021 15351 8079 15357
rect 8021 15317 8033 15351
rect 8067 15317 8079 15351
rect 8021 15311 8079 15317
rect 8205 15351 8263 15357
rect 8205 15317 8217 15351
rect 8251 15348 8263 15351
rect 8662 15348 8668 15360
rect 8251 15320 8668 15348
rect 8251 15317 8263 15320
rect 8205 15311 8263 15317
rect 8662 15308 8668 15320
rect 8720 15308 8726 15360
rect 8956 15348 8984 15524
rect 10318 15512 10324 15564
rect 10376 15552 10382 15564
rect 10413 15555 10471 15561
rect 10413 15552 10425 15555
rect 10376 15524 10425 15552
rect 10376 15512 10382 15524
rect 10413 15521 10425 15524
rect 10459 15521 10471 15555
rect 10413 15515 10471 15521
rect 10689 15555 10747 15561
rect 10689 15521 10701 15555
rect 10735 15552 10747 15555
rect 10888 15552 10916 15648
rect 13538 15580 13544 15632
rect 13596 15620 13602 15632
rect 13596 15592 14504 15620
rect 13596 15580 13602 15592
rect 11238 15561 11244 15564
rect 11232 15552 11244 15561
rect 10735 15524 10916 15552
rect 11199 15524 11244 15552
rect 10735 15521 10747 15524
rect 10689 15515 10747 15521
rect 11232 15515 11244 15524
rect 10428 15484 10456 15515
rect 11238 15512 11244 15515
rect 11296 15512 11302 15564
rect 12434 15512 12440 15564
rect 12492 15512 12498 15564
rect 12710 15561 12716 15564
rect 12704 15515 12716 15561
rect 12710 15512 12716 15515
rect 12768 15512 12774 15564
rect 12986 15512 12992 15564
rect 13044 15552 13050 15564
rect 14274 15552 14280 15564
rect 13044 15524 14280 15552
rect 13044 15512 13050 15524
rect 14274 15512 14280 15524
rect 14332 15512 14338 15564
rect 10965 15487 11023 15493
rect 10965 15484 10977 15487
rect 10428 15456 10977 15484
rect 10965 15453 10977 15456
rect 11011 15453 11023 15487
rect 10965 15447 11023 15453
rect 13814 15444 13820 15496
rect 13872 15484 13878 15496
rect 14476 15493 14504 15592
rect 15470 15580 15476 15632
rect 15528 15580 15534 15632
rect 15841 15623 15899 15629
rect 15841 15589 15853 15623
rect 15887 15620 15899 15623
rect 17230 15623 17288 15629
rect 17230 15620 17242 15623
rect 15887 15592 17242 15620
rect 15887 15589 15899 15592
rect 15841 15583 15899 15589
rect 17230 15589 17242 15592
rect 17276 15589 17288 15623
rect 17696 15620 17724 15648
rect 17834 15623 17892 15629
rect 17834 15620 17846 15623
rect 17696 15592 17846 15620
rect 17230 15583 17288 15589
rect 17834 15589 17846 15592
rect 17880 15589 17892 15623
rect 17834 15583 17892 15589
rect 18782 15580 18788 15632
rect 18840 15580 18846 15632
rect 18984 15620 19012 15651
rect 21266 15648 21272 15660
rect 21324 15648 21330 15700
rect 22833 15691 22891 15697
rect 22833 15657 22845 15691
rect 22879 15688 22891 15691
rect 23201 15691 23259 15697
rect 22879 15660 23060 15688
rect 22879 15657 22891 15660
rect 22833 15651 22891 15657
rect 22189 15623 22247 15629
rect 18984 15592 19932 15620
rect 15194 15512 15200 15564
rect 15252 15512 15258 15564
rect 15488 15552 15516 15580
rect 15749 15555 15807 15561
rect 15749 15552 15761 15555
rect 15488 15524 15761 15552
rect 15749 15521 15761 15524
rect 15795 15521 15807 15555
rect 15749 15515 15807 15521
rect 15933 15555 15991 15561
rect 15933 15521 15945 15555
rect 15979 15552 15991 15555
rect 18800 15552 18828 15580
rect 15979 15524 18828 15552
rect 19337 15555 19395 15561
rect 15979 15521 15991 15524
rect 15933 15515 15991 15521
rect 19337 15521 19349 15555
rect 19383 15552 19395 15555
rect 19610 15552 19616 15564
rect 19383 15524 19616 15552
rect 19383 15521 19395 15524
rect 19337 15515 19395 15521
rect 14369 15487 14427 15493
rect 14369 15484 14381 15487
rect 13872 15456 14381 15484
rect 13872 15444 13878 15456
rect 14369 15453 14381 15456
rect 14415 15453 14427 15487
rect 14369 15447 14427 15453
rect 14461 15487 14519 15493
rect 14461 15453 14473 15487
rect 14507 15453 14519 15487
rect 14461 15447 14519 15453
rect 15473 15487 15531 15493
rect 15473 15453 15485 15487
rect 15519 15484 15531 15487
rect 15562 15484 15568 15496
rect 15519 15456 15568 15484
rect 15519 15453 15531 15456
rect 15473 15447 15531 15453
rect 15562 15444 15568 15456
rect 15620 15444 15626 15496
rect 15948 15416 15976 15515
rect 19610 15512 19616 15524
rect 19668 15512 19674 15564
rect 19904 15561 19932 15592
rect 22189 15589 22201 15623
rect 22235 15620 22247 15623
rect 23032 15620 23060 15660
rect 23201 15657 23213 15691
rect 23247 15688 23259 15691
rect 23290 15688 23296 15700
rect 23247 15660 23296 15688
rect 23247 15657 23259 15660
rect 23201 15651 23259 15657
rect 23290 15648 23296 15660
rect 23348 15648 23354 15700
rect 23584 15660 24624 15688
rect 23584 15620 23612 15660
rect 24596 15632 24624 15660
rect 24029 15623 24087 15629
rect 22235 15592 22968 15620
rect 23032 15592 23612 15620
rect 22235 15589 22247 15592
rect 22189 15583 22247 15589
rect 19889 15555 19947 15561
rect 19889 15521 19901 15555
rect 19935 15521 19947 15555
rect 19889 15515 19947 15521
rect 20717 15555 20775 15561
rect 20717 15521 20729 15555
rect 20763 15552 20775 15555
rect 20990 15552 20996 15564
rect 20763 15524 20996 15552
rect 20763 15521 20775 15524
rect 20717 15515 20775 15521
rect 20990 15512 20996 15524
rect 21048 15512 21054 15564
rect 22097 15555 22155 15561
rect 22097 15521 22109 15555
rect 22143 15521 22155 15555
rect 22097 15515 22155 15521
rect 22281 15555 22339 15561
rect 22281 15521 22293 15555
rect 22327 15552 22339 15555
rect 22327 15524 22416 15552
rect 22327 15521 22339 15524
rect 22281 15515 22339 15521
rect 17497 15487 17555 15493
rect 17497 15453 17509 15487
rect 17543 15484 17555 15487
rect 17586 15484 17592 15496
rect 17543 15456 17592 15484
rect 17543 15453 17555 15456
rect 17497 15447 17555 15453
rect 17586 15444 17592 15456
rect 17644 15444 17650 15496
rect 19426 15444 19432 15496
rect 19484 15444 19490 15496
rect 20254 15444 20260 15496
rect 20312 15484 20318 15496
rect 21269 15487 21327 15493
rect 21269 15484 21281 15487
rect 20312 15456 21281 15484
rect 20312 15444 20318 15456
rect 21269 15453 21281 15456
rect 21315 15453 21327 15487
rect 21269 15447 21327 15453
rect 11900 15388 12480 15416
rect 11900 15348 11928 15388
rect 8956 15320 11928 15348
rect 12342 15308 12348 15360
rect 12400 15308 12406 15360
rect 12452 15348 12480 15388
rect 13372 15388 15976 15416
rect 13372 15348 13400 15388
rect 19334 15376 19340 15428
rect 19392 15376 19398 15428
rect 22112 15416 22140 15515
rect 22388 15493 22416 15524
rect 22646 15512 22652 15564
rect 22704 15552 22710 15564
rect 22836 15555 22894 15561
rect 22836 15552 22848 15555
rect 22704 15524 22848 15552
rect 22704 15512 22710 15524
rect 22836 15521 22848 15524
rect 22882 15521 22894 15555
rect 22940 15552 22968 15592
rect 23201 15555 23259 15561
rect 23201 15552 23213 15555
rect 22940 15524 23213 15552
rect 22836 15515 22894 15521
rect 23201 15521 23213 15524
rect 23247 15552 23259 15555
rect 23474 15552 23480 15564
rect 23247 15524 23480 15552
rect 23247 15521 23259 15524
rect 23201 15515 23259 15521
rect 23474 15512 23480 15524
rect 23532 15512 23538 15564
rect 23584 15561 23612 15592
rect 23676 15592 23980 15620
rect 23676 15561 23704 15592
rect 23569 15555 23627 15561
rect 23569 15521 23581 15555
rect 23615 15521 23627 15555
rect 23569 15515 23627 15521
rect 23661 15555 23719 15561
rect 23661 15521 23673 15555
rect 23707 15521 23719 15555
rect 23661 15515 23719 15521
rect 23750 15512 23756 15564
rect 23808 15512 23814 15564
rect 23845 15555 23903 15561
rect 23845 15521 23857 15555
rect 23891 15521 23903 15555
rect 23952 15552 23980 15592
rect 24029 15589 24041 15623
rect 24075 15620 24087 15623
rect 24118 15620 24124 15632
rect 24075 15592 24124 15620
rect 24075 15589 24087 15592
rect 24029 15583 24087 15589
rect 24118 15580 24124 15592
rect 24176 15580 24182 15632
rect 24302 15580 24308 15632
rect 24360 15620 24366 15632
rect 24397 15623 24455 15629
rect 24397 15620 24409 15623
rect 24360 15592 24409 15620
rect 24360 15580 24366 15592
rect 24397 15589 24409 15592
rect 24443 15589 24455 15623
rect 24397 15583 24455 15589
rect 24578 15580 24584 15632
rect 24636 15580 24642 15632
rect 24486 15552 24492 15564
rect 23952 15524 24492 15552
rect 23845 15515 23903 15521
rect 22373 15487 22431 15493
rect 22373 15453 22385 15487
rect 22419 15484 22431 15487
rect 22922 15484 22928 15496
rect 22419 15456 22928 15484
rect 22419 15453 22431 15456
rect 22373 15447 22431 15453
rect 22922 15444 22928 15456
rect 22980 15444 22986 15496
rect 23290 15484 23296 15496
rect 23032 15456 23296 15484
rect 22278 15416 22284 15428
rect 22112 15388 22284 15416
rect 22278 15376 22284 15388
rect 22336 15416 22342 15428
rect 22465 15419 22523 15425
rect 22465 15416 22477 15419
rect 22336 15388 22477 15416
rect 22336 15376 22342 15388
rect 22465 15385 22477 15388
rect 22511 15385 22523 15419
rect 22465 15379 22523 15385
rect 12452 15320 13400 15348
rect 13446 15308 13452 15360
rect 13504 15348 13510 15360
rect 13817 15351 13875 15357
rect 13817 15348 13829 15351
rect 13504 15320 13829 15348
rect 13504 15308 13510 15320
rect 13817 15317 13829 15320
rect 13863 15317 13875 15351
rect 13817 15311 13875 15317
rect 13906 15308 13912 15360
rect 13964 15308 13970 15360
rect 14826 15308 14832 15360
rect 14884 15308 14890 15360
rect 21910 15308 21916 15360
rect 21968 15308 21974 15360
rect 23032 15357 23060 15456
rect 23290 15444 23296 15456
rect 23348 15444 23354 15496
rect 23477 15419 23535 15425
rect 23477 15385 23489 15419
rect 23523 15416 23535 15419
rect 23768 15416 23796 15512
rect 23523 15388 23796 15416
rect 23523 15385 23535 15388
rect 23477 15379 23535 15385
rect 23017 15351 23075 15357
rect 23017 15317 23029 15351
rect 23063 15317 23075 15351
rect 23017 15311 23075 15317
rect 23566 15308 23572 15360
rect 23624 15348 23630 15360
rect 23860 15348 23888 15515
rect 24486 15512 24492 15524
rect 24544 15512 24550 15564
rect 25406 15512 25412 15564
rect 25464 15512 25470 15564
rect 23624 15320 23888 15348
rect 23624 15308 23630 15320
rect 24762 15308 24768 15360
rect 24820 15308 24826 15360
rect 25593 15351 25651 15357
rect 25593 15317 25605 15351
rect 25639 15348 25651 15351
rect 26234 15348 26240 15360
rect 25639 15320 26240 15348
rect 25639 15317 25651 15320
rect 25593 15311 25651 15317
rect 26234 15308 26240 15320
rect 26292 15308 26298 15360
rect 552 15258 27416 15280
rect 552 15206 3756 15258
rect 3808 15206 3820 15258
rect 3872 15206 3884 15258
rect 3936 15206 3948 15258
rect 4000 15206 4012 15258
rect 4064 15206 10472 15258
rect 10524 15206 10536 15258
rect 10588 15206 10600 15258
rect 10652 15206 10664 15258
rect 10716 15206 10728 15258
rect 10780 15206 17188 15258
rect 17240 15206 17252 15258
rect 17304 15206 17316 15258
rect 17368 15206 17380 15258
rect 17432 15206 17444 15258
rect 17496 15206 23904 15258
rect 23956 15206 23968 15258
rect 24020 15206 24032 15258
rect 24084 15206 24096 15258
rect 24148 15206 24160 15258
rect 24212 15206 27416 15258
rect 552 15184 27416 15206
rect 934 15104 940 15156
rect 992 15104 998 15156
rect 2038 15144 2044 15156
rect 1688 15116 2044 15144
rect 1026 14968 1032 15020
rect 1084 15008 1090 15020
rect 1688 15017 1716 15116
rect 2038 15104 2044 15116
rect 2096 15144 2102 15156
rect 2682 15144 2688 15156
rect 2096 15116 2688 15144
rect 2096 15104 2102 15116
rect 2682 15104 2688 15116
rect 2740 15104 2746 15156
rect 3510 15104 3516 15156
rect 3568 15144 3574 15156
rect 3881 15147 3939 15153
rect 3881 15144 3893 15147
rect 3568 15116 3893 15144
rect 3568 15104 3574 15116
rect 3881 15113 3893 15116
rect 3927 15113 3939 15147
rect 3881 15107 3939 15113
rect 4430 15104 4436 15156
rect 4488 15144 4494 15156
rect 5353 15147 5411 15153
rect 5353 15144 5365 15147
rect 4488 15116 5365 15144
rect 4488 15104 4494 15116
rect 5353 15113 5365 15116
rect 5399 15113 5411 15147
rect 5353 15107 5411 15113
rect 4522 15076 4528 15088
rect 3528 15048 4528 15076
rect 1673 15011 1731 15017
rect 1673 15008 1685 15011
rect 1084 14980 1685 15008
rect 1084 14968 1090 14980
rect 1673 14977 1685 14980
rect 1719 14977 1731 15011
rect 1673 14971 1731 14977
rect 1581 14943 1639 14949
rect 1581 14909 1593 14943
rect 1627 14909 1639 14943
rect 1581 14903 1639 14909
rect 1940 14943 1998 14949
rect 1940 14909 1952 14943
rect 1986 14940 1998 14943
rect 2406 14940 2412 14952
rect 1986 14912 2412 14940
rect 1986 14909 1998 14912
rect 1940 14903 1998 14909
rect 1596 14872 1624 14903
rect 2406 14900 2412 14912
rect 2464 14900 2470 14952
rect 2498 14900 2504 14952
rect 2556 14940 2562 14952
rect 3528 14949 3556 15048
rect 4522 15036 4528 15048
rect 4580 15036 4586 15088
rect 4706 15036 4712 15088
rect 4764 15036 4770 15088
rect 5368 15076 5396 15107
rect 6546 15104 6552 15156
rect 6604 15104 6610 15156
rect 6641 15147 6699 15153
rect 6641 15113 6653 15147
rect 6687 15144 6699 15147
rect 7006 15144 7012 15156
rect 6687 15116 7012 15144
rect 6687 15113 6699 15116
rect 6641 15107 6699 15113
rect 7006 15104 7012 15116
rect 7064 15104 7070 15156
rect 8205 15147 8263 15153
rect 8205 15113 8217 15147
rect 8251 15144 8263 15147
rect 8386 15144 8392 15156
rect 8251 15116 8392 15144
rect 8251 15113 8263 15116
rect 8205 15107 8263 15113
rect 8386 15104 8392 15116
rect 8444 15104 8450 15156
rect 10226 15104 10232 15156
rect 10284 15144 10290 15156
rect 12986 15144 12992 15156
rect 10284 15116 12992 15144
rect 10284 15104 10290 15116
rect 12986 15104 12992 15116
rect 13044 15104 13050 15156
rect 13357 15147 13415 15153
rect 13357 15113 13369 15147
rect 13403 15144 13415 15147
rect 13814 15144 13820 15156
rect 13403 15116 13820 15144
rect 13403 15113 13415 15116
rect 13357 15107 13415 15113
rect 13814 15104 13820 15116
rect 13872 15104 13878 15156
rect 14734 15104 14740 15156
rect 14792 15144 14798 15156
rect 15194 15144 15200 15156
rect 14792 15116 15200 15144
rect 14792 15104 14798 15116
rect 15194 15104 15200 15116
rect 15252 15104 15258 15156
rect 17589 15147 17647 15153
rect 17589 15113 17601 15147
rect 17635 15144 17647 15147
rect 17770 15144 17776 15156
rect 17635 15116 17776 15144
rect 17635 15113 17647 15116
rect 17589 15107 17647 15113
rect 17770 15104 17776 15116
rect 17828 15104 17834 15156
rect 19613 15147 19671 15153
rect 19613 15113 19625 15147
rect 19659 15144 19671 15147
rect 20254 15144 20260 15156
rect 19659 15116 20260 15144
rect 19659 15113 19671 15116
rect 19613 15107 19671 15113
rect 20254 15104 20260 15116
rect 20312 15104 20318 15156
rect 21082 15104 21088 15156
rect 21140 15144 21146 15156
rect 21361 15147 21419 15153
rect 21361 15144 21373 15147
rect 21140 15116 21373 15144
rect 21140 15104 21146 15116
rect 21361 15113 21373 15116
rect 21407 15113 21419 15147
rect 21361 15107 21419 15113
rect 23290 15104 23296 15156
rect 23348 15104 23354 15156
rect 24762 15104 24768 15156
rect 24820 15144 24826 15156
rect 24857 15147 24915 15153
rect 24857 15144 24869 15147
rect 24820 15116 24869 15144
rect 24820 15104 24826 15116
rect 24857 15113 24869 15116
rect 24903 15113 24915 15147
rect 24857 15107 24915 15113
rect 25041 15147 25099 15153
rect 25041 15113 25053 15147
rect 25087 15144 25099 15147
rect 25406 15144 25412 15156
rect 25087 15116 25412 15144
rect 25087 15113 25099 15116
rect 25041 15107 25099 15113
rect 25406 15104 25412 15116
rect 25464 15104 25470 15156
rect 10413 15079 10471 15085
rect 5368 15048 6868 15076
rect 4724 15008 4752 15036
rect 6840 15020 6868 15048
rect 10413 15045 10425 15079
rect 10459 15076 10471 15079
rect 12253 15079 12311 15085
rect 10459 15048 10916 15076
rect 10459 15045 10471 15048
rect 10413 15039 10471 15045
rect 3620 14980 4752 15008
rect 5905 15011 5963 15017
rect 3620 14949 3648 14980
rect 5905 14977 5917 15011
rect 5951 15008 5963 15011
rect 6270 15008 6276 15020
rect 5951 14980 6276 15008
rect 5951 14977 5963 14980
rect 5905 14971 5963 14977
rect 6270 14968 6276 14980
rect 6328 14968 6334 15020
rect 6454 14968 6460 15020
rect 6512 15008 6518 15020
rect 6549 15011 6607 15017
rect 6549 15008 6561 15011
rect 6512 14980 6561 15008
rect 6512 14968 6518 14980
rect 6549 14977 6561 14980
rect 6595 14977 6607 15011
rect 6549 14971 6607 14977
rect 6822 14968 6828 15020
rect 6880 14968 6886 15020
rect 10888 15008 10916 15048
rect 12253 15045 12265 15079
rect 12299 15076 12311 15079
rect 12618 15076 12624 15088
rect 12299 15048 12624 15076
rect 12299 15045 12311 15048
rect 12253 15039 12311 15045
rect 12618 15036 12624 15048
rect 12676 15036 12682 15088
rect 12710 15036 12716 15088
rect 12768 15036 12774 15088
rect 14090 15036 14096 15088
rect 14148 15076 14154 15088
rect 14550 15076 14556 15088
rect 14148 15048 14556 15076
rect 14148 15036 14154 15048
rect 14550 15036 14556 15048
rect 14608 15036 14614 15088
rect 15562 15036 15568 15088
rect 15620 15036 15626 15088
rect 22922 15036 22928 15088
rect 22980 15076 22986 15088
rect 23937 15079 23995 15085
rect 23937 15076 23949 15079
rect 22980 15048 23949 15076
rect 22980 15036 22986 15048
rect 23937 15045 23949 15048
rect 23983 15076 23995 15079
rect 23983 15048 25360 15076
rect 23983 15045 23995 15048
rect 23937 15039 23995 15045
rect 11057 15011 11115 15017
rect 11057 15008 11069 15011
rect 7852 14980 8892 15008
rect 3237 14943 3295 14949
rect 3237 14940 3249 14943
rect 2556 14912 3249 14940
rect 2556 14900 2562 14912
rect 3237 14909 3249 14912
rect 3283 14909 3295 14943
rect 3237 14903 3295 14909
rect 3421 14943 3479 14949
rect 3421 14909 3433 14943
rect 3467 14909 3479 14943
rect 3421 14903 3479 14909
rect 3513 14943 3571 14949
rect 3513 14909 3525 14943
rect 3559 14909 3571 14943
rect 3513 14903 3571 14909
rect 3605 14943 3663 14949
rect 3605 14909 3617 14943
rect 3651 14909 3663 14943
rect 3605 14903 3663 14909
rect 3436 14872 3464 14903
rect 3694 14900 3700 14952
rect 3752 14940 3758 14952
rect 4065 14943 4123 14949
rect 4065 14940 4077 14943
rect 3752 14912 4077 14940
rect 3752 14900 3758 14912
rect 4065 14909 4077 14912
rect 4111 14940 4123 14943
rect 4111 14912 6684 14940
rect 4111 14909 4123 14912
rect 4065 14903 4123 14909
rect 5074 14872 5080 14884
rect 1596 14844 2360 14872
rect 3436 14844 5080 14872
rect 2332 14816 2360 14844
rect 5074 14832 5080 14844
rect 5132 14832 5138 14884
rect 5534 14832 5540 14884
rect 5592 14832 5598 14884
rect 6089 14875 6147 14881
rect 6089 14841 6101 14875
rect 6135 14841 6147 14875
rect 6089 14835 6147 14841
rect 2314 14764 2320 14816
rect 2372 14764 2378 14816
rect 3053 14807 3111 14813
rect 3053 14773 3065 14807
rect 3099 14804 3111 14807
rect 3142 14804 3148 14816
rect 3099 14776 3148 14804
rect 3099 14773 3111 14776
rect 3053 14767 3111 14773
rect 3142 14764 3148 14776
rect 3200 14804 3206 14816
rect 3418 14804 3424 14816
rect 3200 14776 3424 14804
rect 3200 14764 3206 14776
rect 3418 14764 3424 14776
rect 3476 14764 3482 14816
rect 5552 14804 5580 14832
rect 6104 14804 6132 14835
rect 6178 14832 6184 14884
rect 6236 14872 6242 14884
rect 6273 14875 6331 14881
rect 6273 14872 6285 14875
rect 6236 14844 6285 14872
rect 6236 14832 6242 14844
rect 6273 14841 6285 14844
rect 6319 14841 6331 14875
rect 6273 14835 6331 14841
rect 6362 14832 6368 14884
rect 6420 14832 6426 14884
rect 6656 14872 6684 14912
rect 6730 14900 6736 14952
rect 6788 14900 6794 14952
rect 7852 14940 7880 14980
rect 8864 14952 8892 14980
rect 8956 14980 9168 15008
rect 8481 14943 8539 14949
rect 8481 14940 8493 14943
rect 7024 14912 7880 14940
rect 7944 14912 8493 14940
rect 7024 14872 7052 14912
rect 6656 14844 7052 14872
rect 7092 14875 7150 14881
rect 7092 14841 7104 14875
rect 7138 14872 7150 14875
rect 7944 14872 7972 14912
rect 8481 14909 8493 14912
rect 8527 14909 8539 14943
rect 8481 14903 8539 14909
rect 8662 14900 8668 14952
rect 8720 14900 8726 14952
rect 8846 14900 8852 14952
rect 8904 14900 8910 14952
rect 8956 14949 8984 14980
rect 8941 14943 8999 14949
rect 8941 14909 8953 14943
rect 8987 14909 8999 14943
rect 8941 14903 8999 14909
rect 9033 14943 9091 14949
rect 9033 14909 9045 14943
rect 9079 14909 9091 14943
rect 9033 14903 9091 14909
rect 9048 14872 9076 14903
rect 9140 14884 9168 14980
rect 10888 14980 11069 15008
rect 10888 14952 10916 14980
rect 11057 14977 11069 14980
rect 11103 14977 11115 15011
rect 13906 15008 13912 15020
rect 11057 14971 11115 14977
rect 12912 14980 13912 15008
rect 9674 14900 9680 14952
rect 9732 14940 9738 14952
rect 9732 14912 10456 14940
rect 9732 14900 9738 14912
rect 7138 14844 7972 14872
rect 8312 14844 9076 14872
rect 7138 14841 7150 14844
rect 7092 14835 7150 14841
rect 8312 14816 8340 14844
rect 9122 14832 9128 14884
rect 9180 14832 9186 14884
rect 9300 14875 9358 14881
rect 9300 14841 9312 14875
rect 9346 14872 9358 14875
rect 9398 14872 9404 14884
rect 9346 14844 9404 14872
rect 9346 14841 9358 14844
rect 9300 14835 9358 14841
rect 9398 14832 9404 14844
rect 9456 14832 9462 14884
rect 10428 14872 10456 14912
rect 10870 14900 10876 14952
rect 10928 14900 10934 14952
rect 11793 14943 11851 14949
rect 11793 14909 11805 14943
rect 11839 14940 11851 14943
rect 12342 14940 12348 14952
rect 11839 14912 12348 14940
rect 11839 14909 11851 14912
rect 11793 14903 11851 14909
rect 12342 14900 12348 14912
rect 12400 14900 12406 14952
rect 12912 14949 12940 14980
rect 13906 14968 13912 14980
rect 13964 14968 13970 15020
rect 15197 15011 15255 15017
rect 14384 14980 14964 15008
rect 14384 14952 14412 14980
rect 14936 14952 14964 14980
rect 15197 14977 15209 15011
rect 15243 15008 15255 15011
rect 15378 15008 15384 15020
rect 15243 14980 15384 15008
rect 15243 14977 15255 14980
rect 15197 14971 15255 14977
rect 15378 14968 15384 14980
rect 15436 14968 15442 15020
rect 15933 15011 15991 15017
rect 15933 14977 15945 15011
rect 15979 15008 15991 15011
rect 16206 15008 16212 15020
rect 15979 14980 16212 15008
rect 15979 14977 15991 14980
rect 15933 14971 15991 14977
rect 16206 14968 16212 14980
rect 16264 14968 16270 15020
rect 18046 14968 18052 15020
rect 18104 15008 18110 15020
rect 18141 15011 18199 15017
rect 18141 15008 18153 15011
rect 18104 14980 18153 15008
rect 18104 14968 18110 14980
rect 18141 14977 18153 14980
rect 18187 14977 18199 15011
rect 18141 14971 18199 14977
rect 21729 15011 21787 15017
rect 21729 14977 21741 15011
rect 21775 15008 21787 15011
rect 23658 15008 23664 15020
rect 21775 14980 23664 15008
rect 21775 14977 21787 14980
rect 21729 14971 21787 14977
rect 23658 14968 23664 14980
rect 23716 14968 23722 15020
rect 12897 14943 12955 14949
rect 12897 14909 12909 14943
rect 12943 14909 12955 14943
rect 12897 14903 12955 14909
rect 13078 14900 13084 14952
rect 13136 14900 13142 14952
rect 13170 14900 13176 14952
rect 13228 14940 13234 14952
rect 13446 14940 13452 14952
rect 13228 14912 13452 14940
rect 13228 14900 13234 14912
rect 13446 14900 13452 14912
rect 13504 14900 13510 14952
rect 14277 14943 14335 14949
rect 14277 14940 14289 14943
rect 13648 14912 14289 14940
rect 10428 14844 10640 14872
rect 6730 14804 6736 14816
rect 5552 14776 6736 14804
rect 6730 14764 6736 14776
rect 6788 14764 6794 14816
rect 8294 14764 8300 14816
rect 8352 14764 8358 14816
rect 8849 14807 8907 14813
rect 8849 14773 8861 14807
rect 8895 14804 8907 14807
rect 10226 14804 10232 14816
rect 8895 14776 10232 14804
rect 8895 14773 8907 14776
rect 8849 14767 8907 14773
rect 10226 14764 10232 14776
rect 10284 14764 10290 14816
rect 10502 14764 10508 14816
rect 10560 14764 10566 14816
rect 10612 14804 10640 14844
rect 11698 14832 11704 14884
rect 11756 14872 11762 14884
rect 13648 14881 13676 14912
rect 14277 14909 14289 14912
rect 14323 14909 14335 14943
rect 14277 14903 14335 14909
rect 13633 14875 13691 14881
rect 13633 14872 13645 14875
rect 11756 14844 13645 14872
rect 11756 14832 11762 14844
rect 13633 14841 13645 14844
rect 13679 14841 13691 14875
rect 13633 14835 13691 14841
rect 14001 14875 14059 14881
rect 14001 14841 14013 14875
rect 14047 14872 14059 14875
rect 14090 14872 14096 14884
rect 14047 14844 14096 14872
rect 14047 14841 14059 14844
rect 14001 14835 14059 14841
rect 14090 14832 14096 14844
rect 14148 14832 14154 14884
rect 11793 14807 11851 14813
rect 11793 14804 11805 14807
rect 10612 14776 11805 14804
rect 11793 14773 11805 14776
rect 11839 14773 11851 14807
rect 11793 14767 11851 14773
rect 12066 14764 12072 14816
rect 12124 14804 12130 14816
rect 13538 14804 13544 14816
rect 12124 14776 13544 14804
rect 12124 14764 12130 14776
rect 13538 14764 13544 14776
rect 13596 14764 13602 14816
rect 14292 14804 14320 14903
rect 14366 14900 14372 14952
rect 14424 14900 14430 14952
rect 14461 14943 14519 14949
rect 14461 14909 14473 14943
rect 14507 14909 14519 14943
rect 14461 14903 14519 14909
rect 14645 14943 14703 14949
rect 14645 14909 14657 14943
rect 14691 14940 14703 14943
rect 14734 14940 14740 14952
rect 14691 14912 14740 14940
rect 14691 14909 14703 14912
rect 14645 14903 14703 14909
rect 14476 14872 14504 14903
rect 14734 14900 14740 14912
rect 14792 14900 14798 14952
rect 14918 14900 14924 14952
rect 14976 14900 14982 14952
rect 15565 14943 15623 14949
rect 15565 14909 15577 14943
rect 15611 14909 15623 14943
rect 15565 14903 15623 14909
rect 15286 14872 15292 14884
rect 14476 14844 15292 14872
rect 15286 14832 15292 14844
rect 15344 14872 15350 14884
rect 15580 14872 15608 14903
rect 17954 14900 17960 14952
rect 18012 14900 18018 14952
rect 20737 14943 20795 14949
rect 20737 14909 20749 14943
rect 20783 14940 20795 14943
rect 20783 14912 20852 14940
rect 20783 14909 20795 14912
rect 20737 14903 20795 14909
rect 18414 14872 18420 14884
rect 15344 14844 15608 14872
rect 17788 14844 18420 14872
rect 15344 14832 15350 14844
rect 17788 14804 17816 14844
rect 18414 14832 18420 14844
rect 18472 14872 18478 14884
rect 19242 14872 19248 14884
rect 18472 14844 19248 14872
rect 18472 14832 18478 14844
rect 19242 14832 19248 14844
rect 19300 14872 19306 14884
rect 19429 14875 19487 14881
rect 19429 14872 19441 14875
rect 19300 14844 19441 14872
rect 19300 14832 19306 14844
rect 19429 14841 19441 14844
rect 19475 14841 19487 14875
rect 19429 14835 19487 14841
rect 20824 14816 20852 14912
rect 20898 14900 20904 14952
rect 20956 14940 20962 14952
rect 20993 14943 21051 14949
rect 20993 14940 21005 14943
rect 20956 14912 21005 14940
rect 20956 14900 20962 14912
rect 20993 14909 21005 14912
rect 21039 14909 21051 14943
rect 20993 14903 21051 14909
rect 21637 14943 21695 14949
rect 21637 14909 21649 14943
rect 21683 14940 21695 14943
rect 21910 14940 21916 14952
rect 21683 14912 21916 14940
rect 21683 14909 21695 14912
rect 21637 14903 21695 14909
rect 21910 14900 21916 14912
rect 21968 14900 21974 14952
rect 22830 14900 22836 14952
rect 22888 14900 22894 14952
rect 23474 14900 23480 14952
rect 23532 14900 23538 14952
rect 24029 14943 24087 14949
rect 24029 14909 24041 14943
rect 24075 14909 24087 14943
rect 24029 14903 24087 14909
rect 24121 14943 24179 14949
rect 24121 14909 24133 14943
rect 24167 14940 24179 14943
rect 24228 14940 24256 15048
rect 24167 14912 24256 14940
rect 24305 14943 24363 14949
rect 24167 14909 24179 14912
rect 24121 14903 24179 14909
rect 24305 14909 24317 14943
rect 24351 14909 24363 14943
rect 24305 14903 24363 14909
rect 24044 14872 24072 14903
rect 24320 14872 24348 14903
rect 24394 14900 24400 14952
rect 24452 14900 24458 14952
rect 24578 14900 24584 14952
rect 24636 14940 24642 14952
rect 25332 14949 25360 15048
rect 25317 14943 25375 14949
rect 24636 14912 25268 14940
rect 24636 14900 24642 14912
rect 24044 14844 24256 14872
rect 24320 14844 24624 14872
rect 14292 14776 17816 14804
rect 18049 14807 18107 14813
rect 18049 14773 18061 14807
rect 18095 14804 18107 14807
rect 18230 14804 18236 14816
rect 18095 14776 18236 14804
rect 18095 14773 18107 14776
rect 18049 14767 18107 14773
rect 18230 14764 18236 14776
rect 18288 14764 18294 14816
rect 18322 14764 18328 14816
rect 18380 14804 18386 14816
rect 19153 14807 19211 14813
rect 19153 14804 19165 14807
rect 18380 14776 19165 14804
rect 18380 14764 18386 14776
rect 19153 14773 19165 14776
rect 19199 14773 19211 14807
rect 19153 14767 19211 14773
rect 20806 14764 20812 14816
rect 20864 14764 20870 14816
rect 22278 14764 22284 14816
rect 22336 14764 22342 14816
rect 23014 14764 23020 14816
rect 23072 14764 23078 14816
rect 24118 14764 24124 14816
rect 24176 14764 24182 14816
rect 24228 14804 24256 14844
rect 24394 14804 24400 14816
rect 24228 14776 24400 14804
rect 24394 14764 24400 14776
rect 24452 14764 24458 14816
rect 24596 14813 24624 14844
rect 24670 14832 24676 14884
rect 24728 14832 24734 14884
rect 24889 14875 24947 14881
rect 24889 14872 24901 14875
rect 24780 14844 24901 14872
rect 24581 14807 24639 14813
rect 24581 14773 24593 14807
rect 24627 14804 24639 14807
rect 24780 14804 24808 14844
rect 24889 14841 24901 14844
rect 24935 14872 24947 14875
rect 25133 14875 25191 14881
rect 25133 14872 25145 14875
rect 24935 14844 25145 14872
rect 24935 14841 24947 14844
rect 24889 14835 24947 14841
rect 25133 14841 25145 14844
rect 25179 14841 25191 14875
rect 25240 14872 25268 14912
rect 25317 14909 25329 14943
rect 25363 14909 25375 14943
rect 25317 14903 25375 14909
rect 26234 14900 26240 14952
rect 26292 14940 26298 14952
rect 26706 14943 26764 14949
rect 26706 14940 26718 14943
rect 26292 14912 26718 14940
rect 26292 14900 26298 14912
rect 26706 14909 26718 14912
rect 26752 14909 26764 14943
rect 26706 14903 26764 14909
rect 26878 14900 26884 14952
rect 26936 14940 26942 14952
rect 26973 14943 27031 14949
rect 26973 14940 26985 14943
rect 26936 14912 26985 14940
rect 26936 14900 26942 14912
rect 26973 14909 26985 14912
rect 27019 14909 27031 14943
rect 26973 14903 27031 14909
rect 25240 14844 25636 14872
rect 25133 14835 25191 14841
rect 24627 14776 24808 14804
rect 24627 14773 24639 14776
rect 24581 14767 24639 14773
rect 25222 14764 25228 14816
rect 25280 14804 25286 14816
rect 25608 14813 25636 14844
rect 25501 14807 25559 14813
rect 25501 14804 25513 14807
rect 25280 14776 25513 14804
rect 25280 14764 25286 14776
rect 25501 14773 25513 14776
rect 25547 14773 25559 14807
rect 25501 14767 25559 14773
rect 25593 14807 25651 14813
rect 25593 14773 25605 14807
rect 25639 14773 25651 14807
rect 25593 14767 25651 14773
rect 552 14714 27576 14736
rect 552 14662 7114 14714
rect 7166 14662 7178 14714
rect 7230 14662 7242 14714
rect 7294 14662 7306 14714
rect 7358 14662 7370 14714
rect 7422 14662 13830 14714
rect 13882 14662 13894 14714
rect 13946 14662 13958 14714
rect 14010 14662 14022 14714
rect 14074 14662 14086 14714
rect 14138 14662 20546 14714
rect 20598 14662 20610 14714
rect 20662 14662 20674 14714
rect 20726 14662 20738 14714
rect 20790 14662 20802 14714
rect 20854 14662 27262 14714
rect 27314 14662 27326 14714
rect 27378 14662 27390 14714
rect 27442 14662 27454 14714
rect 27506 14662 27518 14714
rect 27570 14662 27576 14714
rect 552 14640 27576 14662
rect 1026 14560 1032 14612
rect 1084 14560 1090 14612
rect 4522 14600 4528 14612
rect 2746 14572 4528 14600
rect 845 14467 903 14473
rect 845 14433 857 14467
rect 891 14464 903 14467
rect 1044 14464 1072 14560
rect 2746 14544 2774 14572
rect 4522 14560 4528 14572
rect 4580 14560 4586 14612
rect 6362 14560 6368 14612
rect 6420 14600 6426 14612
rect 6914 14600 6920 14612
rect 6420 14572 6920 14600
rect 6420 14560 6426 14572
rect 6914 14560 6920 14572
rect 6972 14560 6978 14612
rect 7466 14560 7472 14612
rect 7524 14560 7530 14612
rect 8018 14560 8024 14612
rect 8076 14560 8082 14612
rect 8110 14560 8116 14612
rect 8168 14600 8174 14612
rect 8168 14572 9168 14600
rect 8168 14560 8174 14572
rect 1118 14541 1124 14544
rect 1112 14495 1124 14541
rect 1176 14532 1182 14544
rect 1176 14504 1212 14532
rect 1118 14492 1124 14495
rect 1176 14492 1182 14504
rect 1762 14492 1768 14544
rect 1820 14532 1826 14544
rect 2130 14532 2136 14544
rect 1820 14504 2136 14532
rect 1820 14492 1826 14504
rect 2130 14492 2136 14504
rect 2188 14532 2194 14544
rect 2682 14532 2688 14544
rect 2188 14504 2688 14532
rect 2188 14492 2194 14504
rect 2682 14492 2688 14504
rect 2740 14532 2774 14544
rect 2740 14504 2912 14532
rect 2740 14492 2746 14504
rect 891 14436 1072 14464
rect 891 14433 903 14436
rect 845 14427 903 14433
rect 2498 14424 2504 14476
rect 2556 14464 2562 14476
rect 2593 14467 2651 14473
rect 2593 14464 2605 14467
rect 2556 14436 2605 14464
rect 2556 14424 2562 14436
rect 2593 14433 2605 14436
rect 2639 14433 2651 14467
rect 2593 14427 2651 14433
rect 2774 14424 2780 14476
rect 2832 14424 2838 14476
rect 2884 14473 2912 14504
rect 3326 14492 3332 14544
rect 3384 14532 3390 14544
rect 6270 14532 6276 14544
rect 3384 14504 6276 14532
rect 3384 14492 3390 14504
rect 6270 14492 6276 14504
rect 6328 14492 6334 14544
rect 7484 14532 7512 14560
rect 6380 14504 7512 14532
rect 8036 14532 8064 14560
rect 9030 14541 9036 14544
rect 9001 14535 9036 14541
rect 9001 14532 9013 14535
rect 8036 14504 9013 14532
rect 2869 14467 2927 14473
rect 2869 14433 2881 14467
rect 2915 14433 2927 14467
rect 2869 14427 2927 14433
rect 2961 14467 3019 14473
rect 2961 14433 2973 14467
rect 3007 14464 3019 14467
rect 4065 14467 4123 14473
rect 4065 14464 4077 14467
rect 3007 14436 4077 14464
rect 3007 14433 3019 14436
rect 2961 14427 3019 14433
rect 4065 14433 4077 14436
rect 4111 14433 4123 14467
rect 4065 14427 4123 14433
rect 4522 14424 4528 14476
rect 4580 14464 4586 14476
rect 6380 14464 6408 14504
rect 9001 14501 9013 14504
rect 9001 14495 9036 14501
rect 9030 14492 9036 14495
rect 9088 14492 9094 14544
rect 9140 14532 9168 14572
rect 9398 14560 9404 14612
rect 9456 14560 9462 14612
rect 9490 14560 9496 14612
rect 9548 14600 9554 14612
rect 10121 14603 10179 14609
rect 10121 14600 10133 14603
rect 9548 14572 10133 14600
rect 9548 14560 9554 14572
rect 10121 14569 10133 14572
rect 10167 14600 10179 14603
rect 11882 14600 11888 14612
rect 10167 14572 11888 14600
rect 10167 14569 10179 14572
rect 10121 14563 10179 14569
rect 9217 14535 9275 14541
rect 9217 14532 9229 14535
rect 9140 14504 9229 14532
rect 9217 14501 9229 14504
rect 9263 14501 9275 14535
rect 9217 14495 9275 14501
rect 9315 14504 9904 14532
rect 4580 14436 6408 14464
rect 6733 14467 6791 14473
rect 4580 14424 4586 14436
rect 6733 14433 6745 14467
rect 6779 14464 6791 14467
rect 6822 14464 6828 14476
rect 6779 14436 6828 14464
rect 6779 14433 6791 14436
rect 6733 14427 6791 14433
rect 6822 14424 6828 14436
rect 6880 14424 6886 14476
rect 7000 14467 7058 14473
rect 7000 14433 7012 14467
rect 7046 14464 7058 14467
rect 8297 14467 8355 14473
rect 8297 14464 8309 14467
rect 7046 14436 8309 14464
rect 7046 14433 7058 14436
rect 7000 14427 7058 14433
rect 8297 14433 8309 14436
rect 8343 14433 8355 14467
rect 8297 14427 8355 14433
rect 8481 14467 8539 14473
rect 8481 14433 8493 14467
rect 8527 14433 8539 14467
rect 8481 14427 8539 14433
rect 3237 14399 3295 14405
rect 3237 14365 3249 14399
rect 3283 14396 3295 14399
rect 3329 14399 3387 14405
rect 3329 14396 3341 14399
rect 3283 14368 3341 14396
rect 3283 14365 3295 14368
rect 3237 14359 3295 14365
rect 3329 14365 3341 14368
rect 3375 14365 3387 14399
rect 3329 14359 3387 14365
rect 3510 14356 3516 14408
rect 3568 14396 3574 14408
rect 4617 14399 4675 14405
rect 4617 14396 4629 14399
rect 3568 14368 4629 14396
rect 3568 14356 3574 14368
rect 4617 14365 4629 14368
rect 4663 14365 4675 14399
rect 4617 14359 4675 14365
rect 4798 14356 4804 14408
rect 4856 14396 4862 14408
rect 4985 14399 5043 14405
rect 4985 14396 4997 14399
rect 4856 14368 4997 14396
rect 4856 14356 4862 14368
rect 4985 14365 4997 14368
rect 5031 14365 5043 14399
rect 4985 14359 5043 14365
rect 6549 14399 6607 14405
rect 6549 14365 6561 14399
rect 6595 14365 6607 14399
rect 8496 14396 8524 14427
rect 8662 14424 8668 14476
rect 8720 14424 8726 14476
rect 8757 14467 8815 14473
rect 8757 14433 8769 14467
rect 8803 14464 8815 14467
rect 8803 14436 8984 14464
rect 8803 14433 8815 14436
rect 8757 14427 8815 14433
rect 8956 14396 8984 14436
rect 9122 14396 9128 14408
rect 8496 14368 8892 14396
rect 8956 14368 9128 14396
rect 6549 14359 6607 14365
rect 3973 14331 4031 14337
rect 3973 14297 3985 14331
rect 4019 14328 4031 14331
rect 4338 14328 4344 14340
rect 4019 14300 4344 14328
rect 4019 14297 4031 14300
rect 3973 14291 4031 14297
rect 4338 14288 4344 14300
rect 4396 14288 4402 14340
rect 5629 14331 5687 14337
rect 5629 14297 5641 14331
rect 5675 14328 5687 14331
rect 6362 14328 6368 14340
rect 5675 14300 6368 14328
rect 5675 14297 5687 14300
rect 5629 14291 5687 14297
rect 6362 14288 6368 14300
rect 6420 14288 6426 14340
rect 2225 14263 2283 14269
rect 2225 14229 2237 14263
rect 2271 14260 2283 14263
rect 2314 14260 2320 14272
rect 2271 14232 2320 14260
rect 2271 14229 2283 14232
rect 2225 14223 2283 14229
rect 2314 14220 2320 14232
rect 2372 14220 2378 14272
rect 5902 14220 5908 14272
rect 5960 14220 5966 14272
rect 6564 14260 6592 14359
rect 8864 14337 8892 14368
rect 9122 14356 9128 14368
rect 9180 14396 9186 14408
rect 9315 14396 9343 14504
rect 9582 14424 9588 14476
rect 9640 14424 9646 14476
rect 9766 14424 9772 14476
rect 9824 14424 9830 14476
rect 9876 14473 9904 14504
rect 10226 14492 10232 14544
rect 10284 14532 10290 14544
rect 10321 14535 10379 14541
rect 10321 14532 10333 14535
rect 10284 14504 10333 14532
rect 10284 14492 10290 14504
rect 10321 14501 10333 14504
rect 10367 14501 10379 14535
rect 10321 14495 10379 14501
rect 10428 14473 10456 14572
rect 11882 14560 11888 14572
rect 11940 14600 11946 14612
rect 13630 14600 13636 14612
rect 11940 14572 13636 14600
rect 11940 14560 11946 14572
rect 13630 14560 13636 14572
rect 13688 14560 13694 14612
rect 13817 14603 13875 14609
rect 13817 14569 13829 14603
rect 13863 14569 13875 14603
rect 13817 14563 13875 14569
rect 11054 14492 11060 14544
rect 11112 14532 11118 14544
rect 11974 14532 11980 14544
rect 11112 14504 11980 14532
rect 11112 14492 11118 14504
rect 11974 14492 11980 14504
rect 12032 14532 12038 14544
rect 12253 14535 12311 14541
rect 12253 14532 12265 14535
rect 12032 14504 12265 14532
rect 12032 14492 12038 14504
rect 12253 14501 12265 14504
rect 12299 14501 12311 14535
rect 13832 14532 13860 14563
rect 14826 14560 14832 14612
rect 14884 14560 14890 14612
rect 15286 14560 15292 14612
rect 15344 14560 15350 14612
rect 19242 14560 19248 14612
rect 19300 14600 19306 14612
rect 22278 14600 22284 14612
rect 19300 14572 21772 14600
rect 19300 14560 19306 14572
rect 14154 14535 14212 14541
rect 14154 14532 14166 14535
rect 13832 14504 14166 14532
rect 12253 14495 12311 14501
rect 14154 14501 14166 14504
rect 14200 14501 14212 14535
rect 14154 14495 14212 14501
rect 9861 14467 9919 14473
rect 9861 14433 9873 14467
rect 9907 14464 9919 14467
rect 10413 14467 10471 14473
rect 9907 14436 10180 14464
rect 9907 14433 9919 14436
rect 9861 14427 9919 14433
rect 9180 14368 9343 14396
rect 10152 14396 10180 14436
rect 10413 14433 10425 14467
rect 10459 14433 10471 14467
rect 10413 14427 10471 14433
rect 13633 14467 13691 14473
rect 13633 14433 13645 14467
rect 13679 14464 13691 14467
rect 14844 14464 14872 14560
rect 19610 14532 19616 14544
rect 14936 14504 19616 14532
rect 14936 14476 14964 14504
rect 13679 14436 14872 14464
rect 13679 14433 13691 14436
rect 13633 14427 13691 14433
rect 14918 14424 14924 14476
rect 14976 14424 14982 14476
rect 17696 14473 17724 14504
rect 19610 14492 19616 14504
rect 19668 14492 19674 14544
rect 19886 14492 19892 14544
rect 19944 14532 19950 14544
rect 20456 14541 20484 14572
rect 20441 14535 20499 14541
rect 19944 14504 20392 14532
rect 19944 14492 19950 14504
rect 20364 14476 20392 14504
rect 20441 14501 20453 14535
rect 20487 14501 20499 14535
rect 20441 14495 20499 14501
rect 21266 14492 21272 14544
rect 21324 14532 21330 14544
rect 21545 14535 21603 14541
rect 21545 14532 21557 14535
rect 21324 14504 21557 14532
rect 21324 14492 21330 14504
rect 21545 14501 21557 14504
rect 21591 14501 21603 14535
rect 21545 14495 21603 14501
rect 16669 14467 16727 14473
rect 16669 14433 16681 14467
rect 16715 14464 16727 14467
rect 17681 14467 17739 14473
rect 16715 14436 16988 14464
rect 16715 14433 16727 14436
rect 16669 14427 16727 14433
rect 10505 14399 10563 14405
rect 10505 14396 10517 14399
rect 10152 14368 10517 14396
rect 9180 14356 9186 14368
rect 10505 14365 10517 14368
rect 10551 14365 10563 14399
rect 10505 14359 10563 14365
rect 8849 14331 8907 14337
rect 8849 14297 8861 14331
rect 8895 14297 8907 14331
rect 8849 14291 8907 14297
rect 9582 14288 9588 14340
rect 9640 14328 9646 14340
rect 9953 14331 10011 14337
rect 9953 14328 9965 14331
rect 9640 14300 9965 14328
rect 9640 14288 9646 14300
rect 9953 14297 9965 14300
rect 9999 14297 10011 14331
rect 10410 14328 10416 14340
rect 9953 14291 10011 14297
rect 10152 14300 10416 14328
rect 7006 14260 7012 14272
rect 6564 14232 7012 14260
rect 7006 14220 7012 14232
rect 7064 14220 7070 14272
rect 8478 14220 8484 14272
rect 8536 14260 8542 14272
rect 9033 14263 9091 14269
rect 9033 14260 9045 14263
rect 8536 14232 9045 14260
rect 8536 14220 8542 14232
rect 9033 14229 9045 14232
rect 9079 14260 9091 14263
rect 9858 14260 9864 14272
rect 9079 14232 9864 14260
rect 9079 14229 9091 14232
rect 9033 14223 9091 14229
rect 9858 14220 9864 14232
rect 9916 14220 9922 14272
rect 10152 14269 10180 14300
rect 10410 14288 10416 14300
rect 10468 14288 10474 14340
rect 10520 14328 10548 14359
rect 10962 14356 10968 14408
rect 11020 14356 11026 14408
rect 12066 14356 12072 14408
rect 12124 14356 12130 14408
rect 12158 14356 12164 14408
rect 12216 14356 12222 14408
rect 13909 14399 13967 14405
rect 13909 14365 13921 14399
rect 13955 14365 13967 14399
rect 13909 14359 13967 14365
rect 11238 14328 11244 14340
rect 10520 14300 11244 14328
rect 11238 14288 11244 14300
rect 11296 14328 11302 14340
rect 11296 14300 11836 14328
rect 11296 14288 11302 14300
rect 11808 14272 11836 14300
rect 10137 14263 10195 14269
rect 10137 14229 10149 14263
rect 10183 14229 10195 14263
rect 10137 14223 10195 14229
rect 11606 14220 11612 14272
rect 11664 14220 11670 14272
rect 11790 14220 11796 14272
rect 11848 14220 11854 14272
rect 12618 14220 12624 14272
rect 12676 14220 12682 14272
rect 13924 14260 13952 14359
rect 16850 14356 16856 14408
rect 16908 14356 16914 14408
rect 16960 14396 16988 14436
rect 17681 14433 17693 14467
rect 17727 14433 17739 14467
rect 17681 14427 17739 14433
rect 18414 14424 18420 14476
rect 18472 14424 18478 14476
rect 18598 14424 18604 14476
rect 18656 14464 18662 14476
rect 18656 14436 18828 14464
rect 18656 14424 18662 14436
rect 17034 14396 17040 14408
rect 16960 14368 17040 14396
rect 17034 14356 17040 14368
rect 17092 14396 17098 14408
rect 17589 14399 17647 14405
rect 17589 14396 17601 14399
rect 17092 14368 17601 14396
rect 17092 14356 17098 14368
rect 17589 14365 17601 14368
rect 17635 14365 17647 14399
rect 17589 14359 17647 14365
rect 18138 14356 18144 14408
rect 18196 14356 18202 14408
rect 18690 14356 18696 14408
rect 18748 14356 18754 14408
rect 18800 14396 18828 14436
rect 18874 14424 18880 14476
rect 18932 14464 18938 14476
rect 19521 14467 19579 14473
rect 19521 14464 19533 14467
rect 18932 14436 19533 14464
rect 18932 14424 18938 14436
rect 19521 14433 19533 14436
rect 19567 14433 19579 14467
rect 19981 14467 20039 14473
rect 19981 14464 19993 14467
rect 19521 14427 19579 14433
rect 19628 14436 19993 14464
rect 19628 14396 19656 14436
rect 19981 14433 19993 14436
rect 20027 14433 20039 14467
rect 19981 14427 20039 14433
rect 20346 14424 20352 14476
rect 20404 14464 20410 14476
rect 20625 14467 20683 14473
rect 20625 14464 20637 14467
rect 20404 14436 20637 14464
rect 20404 14424 20410 14436
rect 20625 14433 20637 14436
rect 20671 14464 20683 14467
rect 21453 14467 21511 14473
rect 21453 14464 21465 14467
rect 20671 14436 21465 14464
rect 20671 14433 20683 14436
rect 20625 14427 20683 14433
rect 21453 14433 21465 14436
rect 21499 14433 21511 14467
rect 21453 14427 21511 14433
rect 21637 14467 21695 14473
rect 21637 14433 21649 14467
rect 21683 14433 21695 14467
rect 21637 14427 21695 14433
rect 18800 14368 19656 14396
rect 19702 14356 19708 14408
rect 19760 14396 19766 14408
rect 19797 14399 19855 14405
rect 19797 14396 19809 14399
rect 19760 14368 19809 14396
rect 19760 14356 19766 14368
rect 19797 14365 19809 14368
rect 19843 14396 19855 14399
rect 19886 14396 19892 14408
rect 19843 14368 19892 14396
rect 19843 14365 19855 14368
rect 19797 14359 19855 14365
rect 19886 14356 19892 14368
rect 19944 14356 19950 14408
rect 16868 14328 16896 14356
rect 18708 14328 18736 14356
rect 21652 14328 21680 14427
rect 21744 14396 21772 14572
rect 22066 14572 22284 14600
rect 22066 14532 22094 14572
rect 22278 14560 22284 14572
rect 22336 14560 22342 14612
rect 22370 14560 22376 14612
rect 22428 14560 22434 14612
rect 23014 14600 23020 14612
rect 22848 14572 23020 14600
rect 21836 14504 22094 14532
rect 21836 14473 21864 14504
rect 21821 14467 21879 14473
rect 21821 14433 21833 14467
rect 21867 14433 21879 14467
rect 21821 14427 21879 14433
rect 22005 14467 22063 14473
rect 22005 14433 22017 14467
rect 22051 14433 22063 14467
rect 22388 14464 22416 14560
rect 22848 14541 22876 14572
rect 23014 14560 23020 14572
rect 23072 14560 23078 14612
rect 23124 14572 23428 14600
rect 22833 14535 22891 14541
rect 22833 14501 22845 14535
rect 22879 14501 22891 14535
rect 23124 14532 23152 14572
rect 23400 14544 23428 14572
rect 24118 14560 24124 14612
rect 24176 14560 24182 14612
rect 24302 14560 24308 14612
rect 24360 14600 24366 14612
rect 24489 14603 24547 14609
rect 24489 14600 24501 14603
rect 24360 14572 24501 14600
rect 24360 14560 24366 14572
rect 24489 14569 24501 14572
rect 24535 14569 24547 14603
rect 24489 14563 24547 14569
rect 24578 14560 24584 14612
rect 24636 14560 24642 14612
rect 24670 14560 24676 14612
rect 24728 14600 24734 14612
rect 24728 14572 25176 14600
rect 24728 14560 24734 14572
rect 22833 14495 22891 14501
rect 22940 14504 23152 14532
rect 22649 14467 22707 14473
rect 22649 14464 22661 14467
rect 22388 14436 22661 14464
rect 22005 14427 22063 14433
rect 22649 14433 22661 14436
rect 22695 14433 22707 14467
rect 22649 14427 22707 14433
rect 22741 14467 22799 14473
rect 22741 14433 22753 14467
rect 22787 14464 22799 14467
rect 22940 14464 22968 14504
rect 23382 14492 23388 14544
rect 23440 14492 23446 14544
rect 22787 14436 22968 14464
rect 22787 14433 22799 14436
rect 22741 14427 22799 14433
rect 22020 14396 22048 14427
rect 23014 14424 23020 14476
rect 23072 14424 23078 14476
rect 23107 14457 23165 14463
rect 23107 14423 23119 14457
rect 23153 14423 23165 14457
rect 23198 14424 23204 14476
rect 23256 14473 23262 14476
rect 23256 14467 23283 14473
rect 23271 14433 23283 14467
rect 23256 14427 23283 14433
rect 23256 14424 23262 14427
rect 23107 14417 23165 14423
rect 21744 14368 22048 14396
rect 16868 14300 18736 14328
rect 21008 14300 21680 14328
rect 23124 14328 23152 14417
rect 24136 14396 24164 14560
rect 24394 14492 24400 14544
rect 24452 14532 24458 14544
rect 24452 14504 24716 14532
rect 24452 14492 24458 14504
rect 24688 14473 24716 14504
rect 24673 14467 24731 14473
rect 24673 14433 24685 14467
rect 24719 14464 24731 14467
rect 25038 14464 25044 14476
rect 24719 14436 25044 14464
rect 24719 14433 24731 14436
rect 24673 14427 24731 14433
rect 25038 14424 25044 14436
rect 25096 14424 25102 14476
rect 25148 14464 25176 14572
rect 25222 14560 25228 14612
rect 25280 14600 25286 14612
rect 25793 14603 25851 14609
rect 25793 14600 25805 14603
rect 25280 14572 25805 14600
rect 25280 14560 25286 14572
rect 25793 14569 25805 14572
rect 25839 14569 25851 14603
rect 25793 14563 25851 14569
rect 25961 14603 26019 14609
rect 25961 14569 25973 14603
rect 26007 14569 26019 14603
rect 25961 14563 26019 14569
rect 25317 14535 25375 14541
rect 25317 14501 25329 14535
rect 25363 14532 25375 14535
rect 25498 14532 25504 14544
rect 25363 14504 25504 14532
rect 25363 14501 25375 14504
rect 25317 14495 25375 14501
rect 25498 14492 25504 14504
rect 25556 14492 25562 14544
rect 25593 14535 25651 14541
rect 25593 14501 25605 14535
rect 25639 14501 25651 14535
rect 25593 14495 25651 14501
rect 25406 14464 25412 14476
rect 25148 14436 25412 14464
rect 25406 14424 25412 14436
rect 25464 14464 25470 14476
rect 25608 14464 25636 14495
rect 25464 14436 25636 14464
rect 25976 14464 26004 14563
rect 26053 14467 26111 14473
rect 26053 14464 26065 14467
rect 25976 14436 26065 14464
rect 25464 14424 25470 14436
rect 26053 14433 26065 14436
rect 26099 14433 26111 14467
rect 26053 14427 26111 14433
rect 26605 14467 26663 14473
rect 26605 14433 26617 14467
rect 26651 14433 26663 14467
rect 26605 14427 26663 14433
rect 26620 14396 26648 14427
rect 24136 14368 25452 14396
rect 24762 14328 24768 14340
rect 23124 14300 24768 14328
rect 21008 14272 21036 14300
rect 24762 14288 24768 14300
rect 24820 14288 24826 14340
rect 24854 14288 24860 14340
rect 24912 14288 24918 14340
rect 24949 14331 25007 14337
rect 24949 14297 24961 14331
rect 24995 14328 25007 14331
rect 25130 14328 25136 14340
rect 24995 14300 25136 14328
rect 24995 14297 25007 14300
rect 24949 14291 25007 14297
rect 14642 14260 14648 14272
rect 13924 14232 14648 14260
rect 14642 14220 14648 14232
rect 14700 14220 14706 14272
rect 16482 14220 16488 14272
rect 16540 14220 16546 14272
rect 19518 14220 19524 14272
rect 19576 14260 19582 14272
rect 19613 14263 19671 14269
rect 19613 14260 19625 14263
rect 19576 14232 19625 14260
rect 19576 14220 19582 14232
rect 19613 14229 19625 14232
rect 19659 14229 19671 14263
rect 19613 14223 19671 14229
rect 19702 14220 19708 14272
rect 19760 14220 19766 14272
rect 19794 14220 19800 14272
rect 19852 14260 19858 14272
rect 20073 14263 20131 14269
rect 20073 14260 20085 14263
rect 19852 14232 20085 14260
rect 19852 14220 19858 14232
rect 20073 14229 20085 14232
rect 20119 14260 20131 14263
rect 20254 14260 20260 14272
rect 20119 14232 20260 14260
rect 20119 14229 20131 14232
rect 20073 14223 20131 14229
rect 20254 14220 20260 14232
rect 20312 14220 20318 14272
rect 20809 14263 20867 14269
rect 20809 14229 20821 14263
rect 20855 14260 20867 14263
rect 20990 14260 20996 14272
rect 20855 14232 20996 14260
rect 20855 14229 20867 14232
rect 20809 14223 20867 14229
rect 20990 14220 20996 14232
rect 21048 14220 21054 14272
rect 21269 14263 21327 14269
rect 21269 14229 21281 14263
rect 21315 14260 21327 14263
rect 21542 14260 21548 14272
rect 21315 14232 21548 14260
rect 21315 14229 21327 14232
rect 21269 14223 21327 14229
rect 21542 14220 21548 14232
rect 21600 14220 21606 14272
rect 22278 14220 22284 14272
rect 22336 14220 22342 14272
rect 22462 14220 22468 14272
rect 22520 14220 22526 14272
rect 23293 14263 23351 14269
rect 23293 14229 23305 14263
rect 23339 14260 23351 14263
rect 23750 14260 23756 14272
rect 23339 14232 23756 14260
rect 23339 14229 23351 14232
rect 23293 14223 23351 14229
rect 23750 14220 23756 14232
rect 23808 14220 23814 14272
rect 24305 14263 24363 14269
rect 24305 14229 24317 14263
rect 24351 14260 24363 14263
rect 24964 14260 24992 14291
rect 25130 14288 25136 14300
rect 25188 14288 25194 14340
rect 24351 14232 24992 14260
rect 24351 14229 24363 14232
rect 24305 14223 24363 14229
rect 25314 14220 25320 14272
rect 25372 14220 25378 14272
rect 25424 14260 25452 14368
rect 25516 14368 26648 14396
rect 25516 14337 25544 14368
rect 25501 14331 25559 14337
rect 25501 14297 25513 14331
rect 25547 14297 25559 14331
rect 25501 14291 25559 14297
rect 26142 14288 26148 14340
rect 26200 14328 26206 14340
rect 26421 14331 26479 14337
rect 26421 14328 26433 14331
rect 26200 14300 26433 14328
rect 26200 14288 26206 14300
rect 26421 14297 26433 14300
rect 26467 14297 26479 14331
rect 26421 14291 26479 14297
rect 25777 14263 25835 14269
rect 25777 14260 25789 14263
rect 25424 14232 25789 14260
rect 25777 14229 25789 14232
rect 25823 14229 25835 14263
rect 25777 14223 25835 14229
rect 26234 14220 26240 14272
rect 26292 14220 26298 14272
rect 552 14170 27416 14192
rect 552 14118 3756 14170
rect 3808 14118 3820 14170
rect 3872 14118 3884 14170
rect 3936 14118 3948 14170
rect 4000 14118 4012 14170
rect 4064 14118 10472 14170
rect 10524 14118 10536 14170
rect 10588 14118 10600 14170
rect 10652 14118 10664 14170
rect 10716 14118 10728 14170
rect 10780 14118 17188 14170
rect 17240 14118 17252 14170
rect 17304 14118 17316 14170
rect 17368 14118 17380 14170
rect 17432 14118 17444 14170
rect 17496 14118 23904 14170
rect 23956 14118 23968 14170
rect 24020 14118 24032 14170
rect 24084 14118 24096 14170
rect 24148 14118 24160 14170
rect 24212 14118 27416 14170
rect 552 14096 27416 14118
rect 1397 14059 1455 14065
rect 1397 14025 1409 14059
rect 1443 14056 1455 14059
rect 2774 14056 2780 14068
rect 1443 14028 2780 14056
rect 1443 14025 1455 14028
rect 1397 14019 1455 14025
rect 2774 14016 2780 14028
rect 2832 14016 2838 14068
rect 3237 14059 3295 14065
rect 3237 14025 3249 14059
rect 3283 14056 3295 14059
rect 3510 14056 3516 14068
rect 3283 14028 3516 14056
rect 3283 14025 3295 14028
rect 3237 14019 3295 14025
rect 3510 14016 3516 14028
rect 3568 14016 3574 14068
rect 4430 14016 4436 14068
rect 4488 14056 4494 14068
rect 4488 14028 4660 14056
rect 4488 14016 4494 14028
rect 4632 13929 4660 14028
rect 5074 14016 5080 14068
rect 5132 14056 5138 14068
rect 6641 14059 6699 14065
rect 6641 14056 6653 14059
rect 5132 14028 6653 14056
rect 5132 14016 5138 14028
rect 6641 14025 6653 14028
rect 6687 14025 6699 14059
rect 6641 14019 6699 14025
rect 6822 14016 6828 14068
rect 6880 14016 6886 14068
rect 7006 14016 7012 14068
rect 7064 14016 7070 14068
rect 7193 14059 7251 14065
rect 7193 14025 7205 14059
rect 7239 14056 7251 14059
rect 7466 14056 7472 14068
rect 7239 14028 7472 14056
rect 7239 14025 7251 14028
rect 7193 14019 7251 14025
rect 4617 13923 4675 13929
rect 1228 13892 2636 13920
rect 1228 13861 1256 13892
rect 1213 13855 1271 13861
rect 1213 13821 1225 13855
rect 1259 13821 1271 13855
rect 1213 13815 1271 13821
rect 1489 13855 1547 13861
rect 1489 13821 1501 13855
rect 1535 13821 1547 13855
rect 2608 13852 2636 13892
rect 2746 13892 3004 13920
rect 2746 13852 2774 13892
rect 2608 13824 2774 13852
rect 1489 13815 1547 13821
rect 1029 13787 1087 13793
rect 1029 13753 1041 13787
rect 1075 13753 1087 13787
rect 1029 13747 1087 13753
rect 1044 13716 1072 13747
rect 1302 13744 1308 13796
rect 1360 13784 1366 13796
rect 1504 13784 1532 13815
rect 2866 13812 2872 13864
rect 2924 13812 2930 13864
rect 2976 13852 3004 13892
rect 4617 13889 4629 13923
rect 4663 13889 4675 13923
rect 4617 13883 4675 13889
rect 6178 13880 6184 13932
rect 6236 13920 6242 13932
rect 6840 13920 6868 14016
rect 7208 13988 7236 14019
rect 7466 14016 7472 14028
rect 7524 14016 7530 14068
rect 8662 14016 8668 14068
rect 8720 14056 8726 14068
rect 11054 14056 11060 14068
rect 8720 14028 11060 14056
rect 8720 14016 8726 14028
rect 11054 14016 11060 14028
rect 11112 14016 11118 14068
rect 12158 14016 12164 14068
rect 12216 14056 12222 14068
rect 12713 14059 12771 14065
rect 12713 14056 12725 14059
rect 12216 14028 12725 14056
rect 12216 14016 12222 14028
rect 12713 14025 12725 14028
rect 12759 14025 12771 14059
rect 12713 14019 12771 14025
rect 17034 14016 17040 14068
rect 17092 14056 17098 14068
rect 17129 14059 17187 14065
rect 17129 14056 17141 14059
rect 17092 14028 17141 14056
rect 17092 14016 17098 14028
rect 17129 14025 17141 14028
rect 17175 14025 17187 14059
rect 17129 14019 17187 14025
rect 19886 14016 19892 14068
rect 19944 14056 19950 14068
rect 22738 14056 22744 14068
rect 19944 14028 22744 14056
rect 19944 14016 19950 14028
rect 22738 14016 22744 14028
rect 22796 14016 22802 14068
rect 24210 14016 24216 14068
rect 24268 14056 24274 14068
rect 24268 14028 24900 14056
rect 24268 14016 24274 14028
rect 6236 13892 6868 13920
rect 6932 13960 7236 13988
rect 7285 13991 7343 13997
rect 6236 13880 6242 13892
rect 4062 13852 4068 13864
rect 2976 13824 4068 13852
rect 4062 13812 4068 13824
rect 4120 13812 4126 13864
rect 4338 13812 4344 13864
rect 4396 13861 4402 13864
rect 4396 13852 4408 13861
rect 4396 13824 4441 13852
rect 4396 13815 4408 13824
rect 4396 13812 4402 13815
rect 5902 13812 5908 13864
rect 5960 13861 5966 13864
rect 5960 13852 5972 13861
rect 5960 13824 6005 13852
rect 5960 13815 5972 13824
rect 5960 13812 5966 13815
rect 6086 13812 6092 13864
rect 6144 13852 6150 13864
rect 6733 13855 6791 13861
rect 6733 13852 6745 13855
rect 6144 13824 6745 13852
rect 6144 13812 6150 13824
rect 6733 13821 6745 13824
rect 6779 13821 6791 13855
rect 6733 13815 6791 13821
rect 6825 13855 6883 13861
rect 6825 13821 6837 13855
rect 6871 13852 6883 13855
rect 6932 13852 6960 13960
rect 7285 13957 7297 13991
rect 7331 13957 7343 13991
rect 14826 13988 14832 14000
rect 7285 13951 7343 13957
rect 13096 13960 14832 13988
rect 7300 13920 7328 13951
rect 13096 13932 13124 13960
rect 7024 13892 7328 13920
rect 7377 13923 7435 13929
rect 7024 13861 7052 13892
rect 7377 13889 7389 13923
rect 7423 13920 7435 13923
rect 7650 13920 7656 13932
rect 7423 13892 7656 13920
rect 7423 13889 7435 13892
rect 7377 13883 7435 13889
rect 6871 13824 6960 13852
rect 7009 13855 7067 13861
rect 6871 13821 6883 13824
rect 6825 13815 6883 13821
rect 7009 13821 7021 13855
rect 7055 13821 7067 13855
rect 7009 13815 7067 13821
rect 7101 13855 7159 13861
rect 7101 13821 7113 13855
rect 7147 13821 7159 13855
rect 7392 13852 7420 13883
rect 7650 13880 7656 13892
rect 7708 13880 7714 13932
rect 9048 13892 11376 13920
rect 7101 13815 7159 13821
rect 7309 13824 7420 13852
rect 3326 13784 3332 13796
rect 1360 13756 1532 13784
rect 1596 13756 3332 13784
rect 1360 13744 1366 13756
rect 1118 13716 1124 13728
rect 1044 13688 1124 13716
rect 1118 13676 1124 13688
rect 1176 13716 1182 13728
rect 1596 13716 1624 13756
rect 3326 13744 3332 13756
rect 3384 13744 3390 13796
rect 4724 13756 6224 13784
rect 1176 13688 1624 13716
rect 1176 13676 1182 13688
rect 2130 13676 2136 13728
rect 2188 13676 2194 13728
rect 2222 13676 2228 13728
rect 2280 13676 2286 13728
rect 3050 13676 3056 13728
rect 3108 13716 3114 13728
rect 4724 13716 4752 13756
rect 3108 13688 4752 13716
rect 3108 13676 3114 13688
rect 4798 13676 4804 13728
rect 4856 13676 4862 13728
rect 6196 13716 6224 13756
rect 6270 13744 6276 13796
rect 6328 13744 6334 13796
rect 6362 13744 6368 13796
rect 6420 13784 6426 13796
rect 6457 13787 6515 13793
rect 6457 13784 6469 13787
rect 6420 13756 6469 13784
rect 6420 13744 6426 13756
rect 6457 13753 6469 13756
rect 6503 13784 6515 13787
rect 7116 13784 7144 13815
rect 6503 13756 7144 13784
rect 6503 13753 6515 13756
rect 6457 13747 6515 13753
rect 7309 13716 7337 13824
rect 8846 13812 8852 13864
rect 8904 13852 8910 13864
rect 9048 13861 9076 13892
rect 11348 13864 11376 13892
rect 13078 13880 13084 13932
rect 13136 13880 13142 13932
rect 14366 13920 14372 13932
rect 13464 13892 14372 13920
rect 9033 13855 9091 13861
rect 9033 13852 9045 13855
rect 8904 13824 9045 13852
rect 8904 13812 8910 13824
rect 9033 13821 9045 13824
rect 9079 13821 9091 13855
rect 11241 13855 11299 13861
rect 11241 13852 11253 13855
rect 9033 13815 9091 13821
rect 10796 13824 11253 13852
rect 8202 13744 8208 13796
rect 8260 13744 8266 13796
rect 6196 13688 7337 13716
rect 8220 13716 8248 13744
rect 10796 13728 10824 13824
rect 11241 13821 11253 13824
rect 11287 13821 11299 13855
rect 11241 13815 11299 13821
rect 11330 13812 11336 13864
rect 11388 13812 11394 13864
rect 12710 13812 12716 13864
rect 12768 13852 12774 13864
rect 12897 13855 12955 13861
rect 12897 13852 12909 13855
rect 12768 13824 12909 13852
rect 12768 13812 12774 13824
rect 12897 13821 12909 13824
rect 12943 13821 12955 13855
rect 12897 13815 12955 13821
rect 11508 13787 11566 13793
rect 11508 13753 11520 13787
rect 11554 13784 11566 13787
rect 12250 13784 12256 13796
rect 11554 13756 12256 13784
rect 11554 13753 11566 13756
rect 11508 13747 11566 13753
rect 12250 13744 12256 13756
rect 12308 13744 12314 13796
rect 13464 13784 13492 13892
rect 14366 13880 14372 13892
rect 14424 13880 14430 13932
rect 14660 13929 14688 13960
rect 14826 13948 14832 13960
rect 14884 13948 14890 14000
rect 17497 13991 17555 13997
rect 17497 13957 17509 13991
rect 17543 13957 17555 13991
rect 17497 13951 17555 13957
rect 22833 13991 22891 13997
rect 22833 13957 22845 13991
rect 22879 13988 22891 13991
rect 23198 13988 23204 14000
rect 22879 13960 23204 13988
rect 22879 13957 22891 13960
rect 22833 13951 22891 13957
rect 14645 13923 14703 13929
rect 14645 13889 14657 13923
rect 14691 13889 14703 13923
rect 14645 13883 14703 13889
rect 14734 13880 14740 13932
rect 14792 13920 14798 13932
rect 15749 13923 15807 13929
rect 15749 13920 15761 13923
rect 14792 13892 15761 13920
rect 14792 13880 14798 13892
rect 15749 13889 15761 13892
rect 15795 13889 15807 13923
rect 15749 13883 15807 13889
rect 13541 13855 13599 13861
rect 13541 13821 13553 13855
rect 13587 13821 13599 13855
rect 13725 13855 13783 13861
rect 13725 13852 13737 13855
rect 13541 13815 13599 13821
rect 13648 13824 13737 13852
rect 12406 13756 13492 13784
rect 10318 13716 10324 13728
rect 8220 13688 10324 13716
rect 10318 13676 10324 13688
rect 10376 13716 10382 13728
rect 10778 13716 10784 13728
rect 10376 13688 10784 13716
rect 10376 13676 10382 13688
rect 10778 13676 10784 13688
rect 10836 13676 10842 13728
rect 11054 13676 11060 13728
rect 11112 13716 11118 13728
rect 12406 13716 12434 13756
rect 11112 13688 12434 13716
rect 12621 13719 12679 13725
rect 11112 13676 11118 13688
rect 12621 13685 12633 13719
rect 12667 13716 12679 13719
rect 12710 13716 12716 13728
rect 12667 13688 12716 13716
rect 12667 13685 12679 13688
rect 12621 13679 12679 13685
rect 12710 13676 12716 13688
rect 12768 13676 12774 13728
rect 13078 13676 13084 13728
rect 13136 13716 13142 13728
rect 13556 13716 13584 13815
rect 13648 13728 13676 13824
rect 13725 13821 13737 13824
rect 13771 13821 13783 13855
rect 13725 13815 13783 13821
rect 14550 13812 14556 13864
rect 14608 13812 14614 13864
rect 14829 13855 14887 13861
rect 14829 13821 14841 13855
rect 14875 13821 14887 13855
rect 14829 13815 14887 13821
rect 14844 13784 14872 13815
rect 15470 13812 15476 13864
rect 15528 13812 15534 13864
rect 16005 13855 16063 13861
rect 16005 13852 16017 13855
rect 15672 13824 16017 13852
rect 14476 13756 14872 13784
rect 14476 13728 14504 13756
rect 13136 13688 13584 13716
rect 13136 13676 13142 13688
rect 13630 13676 13636 13728
rect 13688 13676 13694 13728
rect 13909 13719 13967 13725
rect 13909 13685 13921 13719
rect 13955 13716 13967 13719
rect 14182 13716 14188 13728
rect 13955 13688 14188 13716
rect 13955 13685 13967 13688
rect 13909 13679 13967 13685
rect 14182 13676 14188 13688
rect 14240 13676 14246 13728
rect 14274 13676 14280 13728
rect 14332 13716 14338 13728
rect 14369 13719 14427 13725
rect 14369 13716 14381 13719
rect 14332 13688 14381 13716
rect 14332 13676 14338 13688
rect 14369 13685 14381 13688
rect 14415 13685 14427 13719
rect 14369 13679 14427 13685
rect 14458 13676 14464 13728
rect 14516 13676 14522 13728
rect 15010 13676 15016 13728
rect 15068 13676 15074 13728
rect 15672 13725 15700 13824
rect 16005 13821 16017 13824
rect 16051 13821 16063 13855
rect 16005 13815 16063 13821
rect 17405 13855 17463 13861
rect 17405 13821 17417 13855
rect 17451 13852 17463 13855
rect 17512 13852 17540 13951
rect 23198 13948 23204 13960
rect 23256 13988 23262 14000
rect 23256 13960 23520 13988
rect 23256 13948 23262 13960
rect 18046 13920 18052 13932
rect 17451 13824 17540 13852
rect 17584 13892 18052 13920
rect 17451 13821 17463 13824
rect 17405 13815 17463 13821
rect 16666 13744 16672 13796
rect 16724 13784 16730 13796
rect 17584 13784 17612 13892
rect 18046 13880 18052 13892
rect 18104 13880 18110 13932
rect 18598 13880 18604 13932
rect 18656 13880 18662 13932
rect 23492 13929 23520 13960
rect 23842 13948 23848 14000
rect 23900 13988 23906 14000
rect 24872 13988 24900 14028
rect 24946 14016 24952 14068
rect 25004 14016 25010 14068
rect 25038 14016 25044 14068
rect 25096 14056 25102 14068
rect 25593 14059 25651 14065
rect 25593 14056 25605 14059
rect 25096 14028 25605 14056
rect 25096 14016 25102 14028
rect 25593 14025 25605 14028
rect 25639 14025 25651 14059
rect 25593 14019 25651 14025
rect 25317 13991 25375 13997
rect 25317 13988 25329 13991
rect 23900 13960 24624 13988
rect 24872 13960 25329 13988
rect 23900 13948 23906 13960
rect 23477 13923 23535 13929
rect 23477 13889 23489 13923
rect 23523 13889 23535 13923
rect 23477 13883 23535 13889
rect 23750 13880 23756 13932
rect 23808 13920 23814 13932
rect 24397 13923 24455 13929
rect 24397 13920 24409 13923
rect 23808 13892 24409 13920
rect 23808 13880 23814 13892
rect 24397 13889 24409 13892
rect 24443 13889 24455 13923
rect 24397 13883 24455 13889
rect 17770 13812 17776 13864
rect 17828 13852 17834 13864
rect 17957 13855 18015 13861
rect 17957 13852 17969 13855
rect 17828 13824 17969 13852
rect 17828 13812 17834 13824
rect 17957 13821 17969 13824
rect 18003 13852 18015 13855
rect 18616 13852 18644 13880
rect 18003 13824 18644 13852
rect 19613 13855 19671 13861
rect 18003 13821 18015 13824
rect 17957 13815 18015 13821
rect 19613 13821 19625 13855
rect 19659 13852 19671 13855
rect 19978 13852 19984 13864
rect 19659 13824 19984 13852
rect 19659 13821 19671 13824
rect 19613 13815 19671 13821
rect 19978 13812 19984 13824
rect 20036 13852 20042 13864
rect 20438 13852 20444 13864
rect 20036 13824 20444 13852
rect 20036 13812 20042 13824
rect 20438 13812 20444 13824
rect 20496 13812 20502 13864
rect 21453 13855 21511 13861
rect 21453 13852 21465 13855
rect 20916 13824 21465 13852
rect 16724 13756 17612 13784
rect 16724 13744 16730 13756
rect 20916 13728 20944 13824
rect 21453 13821 21465 13824
rect 21499 13821 21511 13855
rect 21453 13815 21511 13821
rect 22830 13812 22836 13864
rect 22888 13852 22894 13864
rect 24029 13855 24087 13861
rect 24029 13852 24041 13855
rect 22888 13824 24041 13852
rect 22888 13812 22894 13824
rect 24029 13821 24041 13824
rect 24075 13821 24087 13855
rect 24029 13815 24087 13821
rect 24121 13855 24179 13861
rect 24121 13821 24133 13855
rect 24167 13852 24179 13855
rect 24210 13852 24216 13864
rect 24167 13824 24216 13852
rect 24167 13821 24179 13824
rect 24121 13815 24179 13821
rect 21082 13744 21088 13796
rect 21140 13784 21146 13796
rect 21698 13787 21756 13793
rect 21698 13784 21710 13787
rect 21140 13756 21710 13784
rect 21140 13744 21146 13756
rect 21698 13753 21710 13756
rect 21744 13753 21756 13787
rect 21698 13747 21756 13753
rect 23658 13744 23664 13796
rect 23716 13784 23722 13796
rect 24136 13784 24164 13815
rect 24210 13812 24216 13824
rect 24268 13812 24274 13864
rect 23716 13756 24164 13784
rect 23716 13744 23722 13756
rect 24394 13744 24400 13796
rect 24452 13784 24458 13796
rect 24489 13787 24547 13793
rect 24489 13784 24501 13787
rect 24452 13756 24501 13784
rect 24452 13744 24458 13756
rect 24489 13753 24501 13756
rect 24535 13753 24547 13787
rect 24596 13784 24624 13960
rect 25317 13957 25329 13960
rect 25363 13957 25375 13991
rect 25317 13951 25375 13957
rect 24762 13880 24768 13932
rect 24820 13920 24826 13932
rect 24857 13923 24915 13929
rect 24857 13920 24869 13923
rect 24820 13892 24869 13920
rect 24820 13880 24826 13892
rect 24857 13889 24869 13892
rect 24903 13889 24915 13923
rect 24857 13883 24915 13889
rect 25133 13855 25191 13861
rect 25133 13852 25145 13855
rect 24964 13824 25145 13852
rect 24964 13784 24992 13824
rect 25133 13821 25145 13824
rect 25179 13821 25191 13855
rect 25133 13815 25191 13821
rect 25225 13855 25283 13861
rect 25225 13821 25237 13855
rect 25271 13821 25283 13855
rect 25225 13815 25283 13821
rect 25240 13784 25268 13815
rect 26234 13812 26240 13864
rect 26292 13852 26298 13864
rect 26706 13855 26764 13861
rect 26706 13852 26718 13855
rect 26292 13824 26718 13852
rect 26292 13812 26298 13824
rect 26706 13821 26718 13824
rect 26752 13821 26764 13855
rect 26706 13815 26764 13821
rect 26878 13812 26884 13864
rect 26936 13852 26942 13864
rect 26973 13855 27031 13861
rect 26973 13852 26985 13855
rect 26936 13824 26985 13852
rect 26936 13812 26942 13824
rect 26973 13821 26985 13824
rect 27019 13821 27031 13855
rect 26973 13815 27031 13821
rect 24596 13756 24992 13784
rect 25148 13756 25268 13784
rect 24489 13747 24547 13753
rect 15657 13719 15715 13725
rect 15657 13685 15669 13719
rect 15703 13685 15715 13719
rect 15657 13679 15715 13685
rect 17221 13719 17279 13725
rect 17221 13685 17233 13719
rect 17267 13716 17279 13719
rect 17310 13716 17316 13728
rect 17267 13688 17316 13716
rect 17267 13685 17279 13688
rect 17221 13679 17279 13685
rect 17310 13676 17316 13688
rect 17368 13676 17374 13728
rect 17862 13676 17868 13728
rect 17920 13676 17926 13728
rect 20898 13676 20904 13728
rect 20956 13676 20962 13728
rect 22922 13676 22928 13728
rect 22980 13676 22986 13728
rect 23474 13676 23480 13728
rect 23532 13716 23538 13728
rect 24581 13719 24639 13725
rect 24581 13716 24593 13719
rect 23532 13688 24593 13716
rect 23532 13676 23538 13688
rect 24581 13685 24593 13688
rect 24627 13685 24639 13719
rect 24581 13679 24639 13685
rect 24854 13676 24860 13728
rect 24912 13716 24918 13728
rect 25148 13716 25176 13756
rect 24912 13688 25176 13716
rect 24912 13676 24918 13688
rect 552 13626 27576 13648
rect 552 13574 7114 13626
rect 7166 13574 7178 13626
rect 7230 13574 7242 13626
rect 7294 13574 7306 13626
rect 7358 13574 7370 13626
rect 7422 13574 13830 13626
rect 13882 13574 13894 13626
rect 13946 13574 13958 13626
rect 14010 13574 14022 13626
rect 14074 13574 14086 13626
rect 14138 13574 20546 13626
rect 20598 13574 20610 13626
rect 20662 13574 20674 13626
rect 20726 13574 20738 13626
rect 20790 13574 20802 13626
rect 20854 13574 27262 13626
rect 27314 13574 27326 13626
rect 27378 13574 27390 13626
rect 27442 13574 27454 13626
rect 27506 13574 27518 13626
rect 27570 13574 27576 13626
rect 552 13552 27576 13574
rect 2222 13512 2228 13524
rect 2148 13484 2228 13512
rect 1980 13447 2038 13453
rect 1980 13413 1992 13447
rect 2026 13444 2038 13447
rect 2148 13444 2176 13484
rect 2222 13472 2228 13484
rect 2280 13472 2286 13524
rect 2498 13472 2504 13524
rect 2556 13472 2562 13524
rect 2682 13472 2688 13524
rect 2740 13472 2746 13524
rect 2866 13472 2872 13524
rect 2924 13512 2930 13524
rect 2961 13515 3019 13521
rect 2961 13512 2973 13515
rect 2924 13484 2973 13512
rect 2924 13472 2930 13484
rect 2961 13481 2973 13484
rect 3007 13481 3019 13515
rect 4798 13512 4804 13524
rect 2961 13475 3019 13481
rect 3712 13484 4804 13512
rect 2516 13444 2544 13472
rect 2700 13444 2728 13472
rect 2026 13416 2176 13444
rect 2332 13416 2544 13444
rect 2608 13416 2728 13444
rect 3237 13447 3295 13453
rect 2026 13413 2038 13416
rect 1980 13407 2038 13413
rect 2130 13336 2136 13388
rect 2188 13336 2194 13388
rect 2222 13336 2228 13388
rect 2280 13336 2286 13388
rect 2332 13385 2360 13416
rect 2317 13379 2375 13385
rect 2317 13345 2329 13379
rect 2363 13345 2375 13379
rect 2317 13339 2375 13345
rect 2406 13336 2412 13388
rect 2464 13376 2470 13388
rect 2608 13385 2636 13416
rect 3237 13413 3249 13447
rect 3283 13444 3295 13447
rect 3326 13444 3332 13456
rect 3283 13416 3332 13444
rect 3283 13413 3295 13416
rect 3237 13407 3295 13413
rect 3326 13404 3332 13416
rect 3384 13404 3390 13456
rect 3418 13404 3424 13456
rect 3476 13404 3482 13456
rect 2501 13379 2559 13385
rect 2501 13376 2513 13379
rect 2464 13348 2513 13376
rect 2464 13336 2470 13348
rect 2501 13345 2513 13348
rect 2547 13345 2559 13379
rect 2501 13339 2559 13345
rect 2593 13379 2651 13385
rect 2593 13345 2605 13379
rect 2639 13345 2651 13379
rect 2593 13339 2651 13345
rect 2685 13379 2743 13385
rect 2685 13345 2697 13379
rect 2731 13345 2743 13379
rect 2685 13339 2743 13345
rect 2148 13308 2176 13336
rect 2700 13308 2728 13339
rect 3510 13336 3516 13388
rect 3568 13376 3574 13388
rect 3712 13385 3740 13484
rect 4798 13472 4804 13484
rect 4856 13472 4862 13524
rect 5353 13515 5411 13521
rect 5353 13481 5365 13515
rect 5399 13512 5411 13515
rect 6086 13512 6092 13524
rect 5399 13484 6092 13512
rect 5399 13481 5411 13484
rect 5353 13475 5411 13481
rect 6086 13472 6092 13484
rect 6144 13472 6150 13524
rect 9401 13515 9459 13521
rect 9401 13481 9413 13515
rect 9447 13512 9459 13515
rect 9766 13512 9772 13524
rect 9447 13484 9772 13512
rect 9447 13481 9459 13484
rect 9401 13475 9459 13481
rect 9766 13472 9772 13484
rect 9824 13512 9830 13524
rect 10962 13512 10968 13524
rect 9824 13484 10968 13512
rect 9824 13472 9830 13484
rect 10962 13472 10968 13484
rect 11020 13472 11026 13524
rect 12250 13472 12256 13524
rect 12308 13472 12314 13524
rect 12618 13512 12624 13524
rect 12452 13484 12624 13512
rect 3973 13447 4031 13453
rect 3973 13413 3985 13447
rect 4019 13444 4031 13447
rect 4985 13447 5043 13453
rect 4985 13444 4997 13447
rect 4019 13416 4997 13444
rect 4019 13413 4031 13416
rect 3973 13407 4031 13413
rect 4985 13413 4997 13416
rect 5031 13413 5043 13447
rect 5994 13444 6000 13456
rect 4985 13407 5043 13413
rect 5920 13416 6000 13444
rect 3605 13379 3663 13385
rect 3605 13376 3617 13379
rect 3568 13348 3617 13376
rect 3568 13336 3574 13348
rect 3605 13345 3617 13348
rect 3651 13345 3663 13379
rect 3605 13339 3663 13345
rect 3697 13379 3755 13385
rect 3697 13345 3709 13379
rect 3743 13345 3755 13379
rect 3697 13339 3755 13345
rect 4154 13336 4160 13388
rect 4212 13336 4218 13388
rect 5920 13385 5948 13416
rect 5994 13404 6000 13416
rect 6052 13404 6058 13456
rect 6172 13447 6230 13453
rect 6172 13413 6184 13447
rect 6218 13444 6230 13447
rect 6270 13444 6276 13456
rect 6218 13416 6276 13444
rect 6218 13413 6230 13416
rect 6172 13407 6230 13413
rect 6270 13404 6276 13416
rect 6328 13404 6334 13456
rect 10536 13447 10594 13453
rect 10536 13413 10548 13447
rect 10582 13444 10594 13447
rect 11701 13447 11759 13453
rect 11701 13444 11713 13447
rect 10582 13416 11713 13444
rect 10582 13413 10594 13416
rect 10536 13407 10594 13413
rect 11701 13413 11713 13416
rect 11747 13413 11759 13447
rect 11701 13407 11759 13413
rect 11790 13404 11796 13456
rect 11848 13444 11854 13456
rect 11848 13416 12204 13444
rect 11848 13404 11854 13416
rect 4433 13379 4491 13385
rect 4433 13345 4445 13379
rect 4479 13345 4491 13379
rect 4433 13339 4491 13345
rect 5905 13379 5963 13385
rect 5905 13345 5917 13379
rect 5951 13345 5963 13379
rect 5905 13339 5963 13345
rect 6012 13348 7328 13376
rect 2148 13280 2728 13308
rect 3881 13243 3939 13249
rect 3881 13209 3893 13243
rect 3927 13240 3939 13243
rect 4249 13243 4307 13249
rect 4249 13240 4261 13243
rect 3927 13212 4261 13240
rect 3927 13209 3939 13212
rect 3881 13203 3939 13209
rect 4249 13209 4261 13212
rect 4295 13209 4307 13243
rect 4249 13203 4307 13209
rect 4341 13243 4399 13249
rect 4341 13209 4353 13243
rect 4387 13209 4399 13243
rect 4448 13240 4476 13339
rect 4798 13268 4804 13320
rect 4856 13268 4862 13320
rect 4893 13311 4951 13317
rect 4893 13277 4905 13311
rect 4939 13308 4951 13311
rect 6012 13308 6040 13348
rect 4939 13280 6040 13308
rect 7300 13308 7328 13348
rect 8110 13336 8116 13388
rect 8168 13376 8174 13388
rect 8297 13379 8355 13385
rect 8297 13376 8309 13379
rect 8168 13348 8309 13376
rect 8168 13336 8174 13348
rect 8297 13345 8309 13348
rect 8343 13345 8355 13379
rect 11054 13376 11060 13388
rect 8297 13339 8355 13345
rect 8496 13348 11060 13376
rect 7650 13308 7656 13320
rect 7300 13280 7656 13308
rect 4939 13277 4951 13280
rect 4893 13271 4951 13277
rect 5902 13240 5908 13252
rect 4448 13212 5908 13240
rect 4341 13203 4399 13209
rect 845 13175 903 13181
rect 845 13141 857 13175
rect 891 13172 903 13175
rect 1210 13172 1216 13184
rect 891 13144 1216 13172
rect 891 13141 903 13144
rect 845 13135 903 13141
rect 1210 13132 1216 13144
rect 1268 13132 1274 13184
rect 3142 13132 3148 13184
rect 3200 13132 3206 13184
rect 3697 13175 3755 13181
rect 3697 13141 3709 13175
rect 3743 13172 3755 13175
rect 4062 13172 4068 13184
rect 3743 13144 4068 13172
rect 3743 13141 3755 13144
rect 3697 13135 3755 13141
rect 4062 13132 4068 13144
rect 4120 13132 4126 13184
rect 4356 13172 4384 13203
rect 5902 13200 5908 13212
rect 5960 13200 5966 13252
rect 7300 13249 7328 13280
rect 7650 13268 7656 13280
rect 7708 13308 7714 13320
rect 7929 13311 7987 13317
rect 7929 13308 7941 13311
rect 7708 13280 7941 13308
rect 7708 13268 7714 13280
rect 7929 13277 7941 13280
rect 7975 13277 7987 13311
rect 7929 13271 7987 13277
rect 8386 13268 8392 13320
rect 8444 13268 8450 13320
rect 7285 13243 7343 13249
rect 7285 13209 7297 13243
rect 7331 13209 7343 13243
rect 7285 13203 7343 13209
rect 7742 13200 7748 13252
rect 7800 13240 7806 13252
rect 8496 13240 8524 13348
rect 11054 13336 11060 13348
rect 11112 13336 11118 13388
rect 11882 13336 11888 13388
rect 11940 13336 11946 13388
rect 12176 13385 12204 13416
rect 12452 13385 12480 13484
rect 12618 13472 12624 13484
rect 12676 13472 12682 13524
rect 14458 13472 14464 13524
rect 14516 13512 14522 13524
rect 15381 13515 15439 13521
rect 15381 13512 15393 13515
rect 14516 13484 15393 13512
rect 14516 13472 14522 13484
rect 15381 13481 15393 13484
rect 15427 13481 15439 13515
rect 15381 13475 15439 13481
rect 15470 13472 15476 13524
rect 15528 13512 15534 13524
rect 16117 13515 16175 13521
rect 16117 13512 16129 13515
rect 15528 13484 16129 13512
rect 15528 13472 15534 13484
rect 16117 13481 16129 13484
rect 16163 13481 16175 13515
rect 16117 13475 16175 13481
rect 16482 13472 16488 13524
rect 16540 13472 16546 13524
rect 18414 13472 18420 13524
rect 18472 13472 18478 13524
rect 18785 13515 18843 13521
rect 18785 13481 18797 13515
rect 18831 13512 18843 13515
rect 18874 13512 18880 13524
rect 18831 13484 18880 13512
rect 18831 13481 18843 13484
rect 18785 13475 18843 13481
rect 18874 13472 18880 13484
rect 18932 13472 18938 13524
rect 20441 13515 20499 13521
rect 20441 13481 20453 13515
rect 20487 13512 20499 13515
rect 21082 13512 21088 13524
rect 20487 13484 21088 13512
rect 20487 13481 20499 13484
rect 20441 13475 20499 13481
rect 21082 13472 21088 13484
rect 21140 13472 21146 13524
rect 22649 13515 22707 13521
rect 22649 13481 22661 13515
rect 22695 13512 22707 13515
rect 22830 13512 22836 13524
rect 22695 13484 22836 13512
rect 22695 13481 22707 13484
rect 22649 13475 22707 13481
rect 22830 13472 22836 13484
rect 22888 13472 22894 13524
rect 23014 13472 23020 13524
rect 23072 13512 23078 13524
rect 23385 13515 23443 13521
rect 23385 13512 23397 13515
rect 23072 13484 23397 13512
rect 23072 13472 23078 13484
rect 23385 13481 23397 13484
rect 23431 13481 23443 13515
rect 24121 13515 24179 13521
rect 24121 13512 24133 13515
rect 23385 13475 23443 13481
rect 23952 13484 24133 13512
rect 16577 13447 16635 13453
rect 16577 13444 16589 13447
rect 12544 13416 14780 13444
rect 12544 13385 12572 13416
rect 12802 13385 12808 13388
rect 12069 13379 12127 13385
rect 12069 13345 12081 13379
rect 12115 13345 12127 13379
rect 12069 13339 12127 13345
rect 12161 13379 12219 13385
rect 12161 13345 12173 13379
rect 12207 13345 12219 13379
rect 12161 13339 12219 13345
rect 12437 13379 12495 13385
rect 12437 13345 12449 13379
rect 12483 13345 12495 13379
rect 12437 13339 12495 13345
rect 12529 13379 12587 13385
rect 12529 13345 12541 13379
rect 12575 13345 12587 13379
rect 12529 13339 12587 13345
rect 12796 13339 12808 13385
rect 10778 13268 10784 13320
rect 10836 13268 10842 13320
rect 10870 13268 10876 13320
rect 10928 13308 10934 13320
rect 11517 13311 11575 13317
rect 11517 13308 11529 13311
rect 10928 13280 11529 13308
rect 10928 13268 10934 13280
rect 11517 13277 11529 13280
rect 11563 13277 11575 13311
rect 11517 13271 11575 13277
rect 7800 13212 8524 13240
rect 12084 13240 12112 13339
rect 12802 13336 12808 13339
rect 12860 13336 12866 13388
rect 14016 13385 14044 13416
rect 14752 13388 14780 13416
rect 15212 13416 16589 13444
rect 14274 13385 14280 13388
rect 14001 13379 14059 13385
rect 14001 13345 14013 13379
rect 14047 13345 14059 13379
rect 14268 13376 14280 13385
rect 14235 13348 14280 13376
rect 14001 13339 14059 13345
rect 14268 13339 14280 13348
rect 14274 13336 14280 13339
rect 14332 13336 14338 13388
rect 14734 13336 14740 13388
rect 14792 13336 14798 13388
rect 15212 13320 15240 13416
rect 16577 13413 16589 13416
rect 16623 13444 16635 13447
rect 20898 13444 20904 13456
rect 16623 13416 16804 13444
rect 16623 13413 16635 13416
rect 16577 13407 16635 13413
rect 13906 13268 13912 13320
rect 13964 13268 13970 13320
rect 15194 13268 15200 13320
rect 15252 13268 15258 13320
rect 16666 13268 16672 13320
rect 16724 13268 16730 13320
rect 13924 13240 13952 13268
rect 12084 13212 12434 13240
rect 7800 13200 7806 13212
rect 6914 13172 6920 13184
rect 4356 13144 6920 13172
rect 6914 13132 6920 13144
rect 6972 13132 6978 13184
rect 7374 13132 7380 13184
rect 7432 13132 7438 13184
rect 8570 13132 8576 13184
rect 8628 13132 8634 13184
rect 10962 13132 10968 13184
rect 11020 13132 11026 13184
rect 12406 13172 12434 13212
rect 13556 13212 13952 13240
rect 13556 13172 13584 13212
rect 12406 13144 13584 13172
rect 13630 13132 13636 13184
rect 13688 13172 13694 13184
rect 13909 13175 13967 13181
rect 13909 13172 13921 13175
rect 13688 13144 13921 13172
rect 13688 13132 13694 13144
rect 13909 13141 13921 13144
rect 13955 13141 13967 13175
rect 16776 13172 16804 13416
rect 17052 13416 20904 13444
rect 17052 13385 17080 13416
rect 17604 13388 17632 13416
rect 17310 13385 17316 13388
rect 17037 13379 17095 13385
rect 17037 13345 17049 13379
rect 17083 13345 17095 13379
rect 17304 13376 17316 13385
rect 17271 13348 17316 13376
rect 17037 13339 17095 13345
rect 17304 13339 17316 13348
rect 17310 13336 17316 13339
rect 17368 13336 17374 13388
rect 17586 13336 17592 13388
rect 17644 13336 17650 13388
rect 19886 13336 19892 13388
rect 19944 13385 19950 13388
rect 20180 13385 20208 13416
rect 20898 13404 20904 13416
rect 20956 13444 20962 13456
rect 22922 13444 22928 13456
rect 20956 13416 21312 13444
rect 20956 13404 20962 13416
rect 21284 13388 21312 13416
rect 21376 13416 22928 13444
rect 19944 13339 19956 13385
rect 20165 13379 20223 13385
rect 20165 13345 20177 13379
rect 20211 13345 20223 13379
rect 20165 13339 20223 13345
rect 19944 13336 19950 13339
rect 20254 13336 20260 13388
rect 20312 13336 20318 13388
rect 20346 13336 20352 13388
rect 20404 13376 20410 13388
rect 20530 13376 20536 13388
rect 20404 13348 20536 13376
rect 20404 13336 20410 13348
rect 20530 13336 20536 13348
rect 20588 13376 20594 13388
rect 20625 13379 20683 13385
rect 20625 13376 20637 13379
rect 20588 13348 20637 13376
rect 20588 13336 20594 13348
rect 20625 13345 20637 13348
rect 20671 13345 20683 13379
rect 20625 13339 20683 13345
rect 20717 13379 20775 13385
rect 20717 13345 20729 13379
rect 20763 13345 20775 13379
rect 20717 13339 20775 13345
rect 20809 13379 20867 13385
rect 20809 13345 20821 13379
rect 20855 13345 20867 13379
rect 20809 13339 20867 13345
rect 20993 13379 21051 13385
rect 20993 13345 21005 13379
rect 21039 13345 21051 13379
rect 20993 13339 21051 13345
rect 20272 13308 20300 13336
rect 20732 13308 20760 13339
rect 20272 13280 20760 13308
rect 20824 13240 20852 13339
rect 21008 13308 21036 13339
rect 21266 13336 21272 13388
rect 21324 13336 21330 13388
rect 21376 13308 21404 13416
rect 22922 13404 22928 13416
rect 22980 13404 22986 13456
rect 23032 13416 23520 13444
rect 21542 13385 21548 13388
rect 21536 13376 21548 13385
rect 21503 13348 21548 13376
rect 21536 13339 21548 13348
rect 21542 13336 21548 13339
rect 21600 13336 21606 13388
rect 22462 13336 22468 13388
rect 22520 13336 22526 13388
rect 23032 13385 23060 13416
rect 23492 13388 23520 13416
rect 23017 13379 23075 13385
rect 23017 13345 23029 13379
rect 23063 13345 23075 13379
rect 23017 13339 23075 13345
rect 23201 13379 23259 13385
rect 23201 13345 23213 13379
rect 23247 13376 23259 13379
rect 23290 13376 23296 13388
rect 23247 13348 23296 13376
rect 23247 13345 23259 13348
rect 23201 13339 23259 13345
rect 23290 13336 23296 13348
rect 23348 13336 23354 13388
rect 23474 13336 23480 13388
rect 23532 13336 23538 13388
rect 23569 13379 23627 13385
rect 23569 13345 23581 13379
rect 23615 13345 23627 13379
rect 23569 13339 23627 13345
rect 21008 13280 21404 13308
rect 22480 13308 22508 13336
rect 22925 13311 22983 13317
rect 22925 13308 22937 13311
rect 22480 13280 22937 13308
rect 22925 13277 22937 13280
rect 22971 13277 22983 13311
rect 22925 13271 22983 13277
rect 23106 13268 23112 13320
rect 23164 13268 23170 13320
rect 21082 13240 21088 13252
rect 20824 13212 21088 13240
rect 21082 13200 21088 13212
rect 21140 13200 21146 13252
rect 22830 13200 22836 13252
rect 22888 13240 22894 13252
rect 23584 13240 23612 13339
rect 23658 13336 23664 13388
rect 23716 13336 23722 13388
rect 23750 13336 23756 13388
rect 23808 13336 23814 13388
rect 23842 13336 23848 13388
rect 23900 13336 23906 13388
rect 23952 13385 23980 13484
rect 24121 13481 24133 13484
rect 24167 13512 24179 13515
rect 24167 13484 24716 13512
rect 24167 13481 24179 13484
rect 24121 13475 24179 13481
rect 24688 13444 24716 13484
rect 24854 13472 24860 13524
rect 24912 13472 24918 13524
rect 24946 13472 24952 13524
rect 25004 13472 25010 13524
rect 24964 13444 24992 13472
rect 24688 13416 24992 13444
rect 25992 13447 26050 13453
rect 25992 13413 26004 13447
rect 26038 13444 26050 13447
rect 26142 13444 26148 13456
rect 26038 13416 26148 13444
rect 26038 13413 26050 13416
rect 25992 13407 26050 13413
rect 26142 13404 26148 13416
rect 26200 13404 26206 13456
rect 23937 13379 23995 13385
rect 23937 13345 23949 13379
rect 23983 13345 23995 13379
rect 23937 13339 23995 13345
rect 24029 13379 24087 13385
rect 24029 13345 24041 13379
rect 24075 13345 24087 13379
rect 24029 13339 24087 13345
rect 24213 13379 24271 13385
rect 24213 13345 24225 13379
rect 24259 13345 24271 13379
rect 24213 13339 24271 13345
rect 24489 13379 24547 13385
rect 24489 13345 24501 13379
rect 24535 13376 24547 13379
rect 26237 13379 26295 13385
rect 24535 13348 25176 13376
rect 24535 13345 24547 13348
rect 24489 13339 24547 13345
rect 23768 13308 23796 13336
rect 24044 13308 24072 13339
rect 23768 13280 24072 13308
rect 22888 13212 23612 13240
rect 24228 13240 24256 13339
rect 25148 13320 25176 13348
rect 26237 13345 26249 13379
rect 26283 13376 26295 13379
rect 26878 13376 26884 13388
rect 26283 13348 26884 13376
rect 26283 13345 26295 13348
rect 26237 13339 26295 13345
rect 26878 13336 26884 13348
rect 26936 13336 26942 13388
rect 24673 13311 24731 13317
rect 24673 13277 24685 13311
rect 24719 13308 24731 13311
rect 25038 13308 25044 13320
rect 24719 13280 25044 13308
rect 24719 13277 24731 13280
rect 24673 13271 24731 13277
rect 24394 13240 24400 13252
rect 24228 13212 24400 13240
rect 22888 13200 22894 13212
rect 24394 13200 24400 13212
rect 24452 13240 24458 13252
rect 24688 13240 24716 13271
rect 25038 13268 25044 13280
rect 25096 13268 25102 13320
rect 25130 13268 25136 13320
rect 25188 13268 25194 13320
rect 24452 13212 24716 13240
rect 24452 13200 24458 13212
rect 20254 13172 20260 13184
rect 16776 13144 20260 13172
rect 13909 13135 13967 13141
rect 20254 13132 20260 13144
rect 20312 13132 20318 13184
rect 20622 13132 20628 13184
rect 20680 13172 20686 13184
rect 22741 13175 22799 13181
rect 22741 13172 22753 13175
rect 20680 13144 22753 13172
rect 20680 13132 20686 13144
rect 22741 13141 22753 13144
rect 22787 13172 22799 13175
rect 23566 13172 23572 13184
rect 22787 13144 23572 13172
rect 22787 13141 22799 13144
rect 22741 13135 22799 13141
rect 23566 13132 23572 13144
rect 23624 13132 23630 13184
rect 24302 13132 24308 13184
rect 24360 13132 24366 13184
rect 552 13082 27416 13104
rect 552 13030 3756 13082
rect 3808 13030 3820 13082
rect 3872 13030 3884 13082
rect 3936 13030 3948 13082
rect 4000 13030 4012 13082
rect 4064 13030 10472 13082
rect 10524 13030 10536 13082
rect 10588 13030 10600 13082
rect 10652 13030 10664 13082
rect 10716 13030 10728 13082
rect 10780 13030 17188 13082
rect 17240 13030 17252 13082
rect 17304 13030 17316 13082
rect 17368 13030 17380 13082
rect 17432 13030 17444 13082
rect 17496 13030 23904 13082
rect 23956 13030 23968 13082
rect 24020 13030 24032 13082
rect 24084 13030 24096 13082
rect 24148 13030 24160 13082
rect 24212 13030 27416 13082
rect 552 13008 27416 13030
rect 1581 12971 1639 12977
rect 1581 12937 1593 12971
rect 1627 12968 1639 12971
rect 2406 12968 2412 12980
rect 1627 12940 2412 12968
rect 1627 12937 1639 12940
rect 1581 12931 1639 12937
rect 2406 12928 2412 12940
rect 2464 12928 2470 12980
rect 6270 12928 6276 12980
rect 6328 12928 6334 12980
rect 7374 12928 7380 12980
rect 7432 12928 7438 12980
rect 7929 12971 7987 12977
rect 7929 12937 7941 12971
rect 7975 12968 7987 12971
rect 8110 12968 8116 12980
rect 7975 12940 8116 12968
rect 7975 12937 7987 12940
rect 7929 12931 7987 12937
rect 8110 12928 8116 12940
rect 8168 12928 8174 12980
rect 8570 12928 8576 12980
rect 8628 12928 8634 12980
rect 10962 12928 10968 12980
rect 11020 12928 11026 12980
rect 11698 12928 11704 12980
rect 11756 12928 11762 12980
rect 11882 12928 11888 12980
rect 11940 12928 11946 12980
rect 12802 12928 12808 12980
rect 12860 12928 12866 12980
rect 13464 12940 14044 12968
rect 5074 12900 5080 12912
rect 4356 12872 5080 12900
rect 1118 12724 1124 12776
rect 1176 12764 1182 12776
rect 1213 12767 1271 12773
rect 1213 12764 1225 12767
rect 1176 12736 1225 12764
rect 1176 12724 1182 12736
rect 1213 12733 1225 12736
rect 1259 12733 1271 12767
rect 1213 12727 1271 12733
rect 2222 12724 2228 12776
rect 2280 12764 2286 12776
rect 4356 12773 4384 12872
rect 5074 12860 5080 12872
rect 5132 12860 5138 12912
rect 7101 12903 7159 12909
rect 7101 12900 7113 12903
rect 5828 12872 7113 12900
rect 4632 12804 5396 12832
rect 3053 12767 3111 12773
rect 3053 12764 3065 12767
rect 2280 12736 3065 12764
rect 2280 12724 2286 12736
rect 3053 12733 3065 12736
rect 3099 12733 3111 12767
rect 3053 12727 3111 12733
rect 3789 12767 3847 12773
rect 3789 12733 3801 12767
rect 3835 12733 3847 12767
rect 3789 12727 3847 12733
rect 4249 12767 4307 12773
rect 4249 12733 4261 12767
rect 4295 12733 4307 12767
rect 4249 12727 4307 12733
rect 4341 12767 4399 12773
rect 4341 12733 4353 12767
rect 4387 12733 4399 12767
rect 4341 12727 4399 12733
rect 1397 12699 1455 12705
rect 1397 12665 1409 12699
rect 1443 12696 1455 12699
rect 2314 12696 2320 12708
rect 1443 12668 2320 12696
rect 1443 12665 1455 12668
rect 1397 12659 1455 12665
rect 2314 12656 2320 12668
rect 2372 12696 2378 12708
rect 2682 12696 2688 12708
rect 2372 12668 2688 12696
rect 2372 12656 2378 12668
rect 2682 12656 2688 12668
rect 2740 12656 2746 12708
rect 2774 12656 2780 12708
rect 2832 12705 2838 12708
rect 2832 12659 2844 12705
rect 3804 12696 3832 12727
rect 3160 12668 3832 12696
rect 4264 12696 4292 12727
rect 4430 12724 4436 12776
rect 4488 12724 4494 12776
rect 4632 12773 4660 12804
rect 4617 12767 4675 12773
rect 4617 12733 4629 12767
rect 4663 12733 4675 12767
rect 4617 12727 4675 12733
rect 4798 12724 4804 12776
rect 4856 12764 4862 12776
rect 5261 12767 5319 12773
rect 5261 12764 5273 12767
rect 4856 12736 5273 12764
rect 4856 12724 4862 12736
rect 5261 12733 5273 12736
rect 5307 12733 5319 12767
rect 5261 12727 5319 12733
rect 5368 12764 5396 12804
rect 5629 12767 5687 12773
rect 5629 12764 5641 12767
rect 5368 12736 5641 12764
rect 4709 12699 4767 12705
rect 4709 12696 4721 12699
rect 4264 12668 4721 12696
rect 2832 12656 2838 12659
rect 3160 12640 3188 12668
rect 4709 12665 4721 12668
rect 4755 12665 4767 12699
rect 4709 12659 4767 12665
rect 4982 12656 4988 12708
rect 5040 12696 5046 12708
rect 5368 12696 5396 12736
rect 5629 12733 5641 12736
rect 5675 12764 5687 12767
rect 5718 12764 5724 12776
rect 5675 12736 5724 12764
rect 5675 12733 5687 12736
rect 5629 12727 5687 12733
rect 5718 12724 5724 12736
rect 5776 12724 5782 12776
rect 5828 12773 5856 12872
rect 7101 12869 7113 12872
rect 7147 12869 7159 12903
rect 7101 12863 7159 12869
rect 7392 12832 7420 12928
rect 6012 12804 7420 12832
rect 6012 12773 6040 12804
rect 7742 12792 7748 12844
rect 7800 12792 7806 12844
rect 8588 12832 8616 12928
rect 9677 12835 9735 12841
rect 9677 12832 9689 12835
rect 8588 12804 9689 12832
rect 9677 12801 9689 12804
rect 9723 12801 9735 12835
rect 9677 12795 9735 12801
rect 9766 12792 9772 12844
rect 9824 12792 9830 12844
rect 5813 12767 5871 12773
rect 5813 12733 5825 12767
rect 5859 12733 5871 12767
rect 5813 12727 5871 12733
rect 5905 12767 5963 12773
rect 5905 12733 5917 12767
rect 5951 12733 5963 12767
rect 5905 12727 5963 12733
rect 5997 12767 6055 12773
rect 5997 12733 6009 12767
rect 6043 12733 6055 12767
rect 5997 12727 6055 12733
rect 5920 12696 5948 12727
rect 6454 12724 6460 12776
rect 6512 12724 6518 12776
rect 7760 12764 7788 12792
rect 6564 12736 7788 12764
rect 8021 12767 8079 12773
rect 5040 12668 5396 12696
rect 5828 12668 5948 12696
rect 5040 12656 5046 12668
rect 1302 12588 1308 12640
rect 1360 12628 1366 12640
rect 1673 12631 1731 12637
rect 1673 12628 1685 12631
rect 1360 12600 1685 12628
rect 1360 12588 1366 12600
rect 1673 12597 1685 12600
rect 1719 12628 1731 12631
rect 3142 12628 3148 12640
rect 1719 12600 3148 12628
rect 1719 12597 1731 12600
rect 1673 12591 1731 12597
rect 3142 12588 3148 12600
rect 3200 12588 3206 12640
rect 3234 12588 3240 12640
rect 3292 12588 3298 12640
rect 3970 12588 3976 12640
rect 4028 12588 4034 12640
rect 5074 12588 5080 12640
rect 5132 12628 5138 12640
rect 5828 12628 5856 12668
rect 5132 12600 5856 12628
rect 5132 12588 5138 12600
rect 5902 12588 5908 12640
rect 5960 12628 5966 12640
rect 6564 12628 6592 12736
rect 8021 12733 8033 12767
rect 8067 12764 8079 12767
rect 9784 12764 9812 12792
rect 8067 12736 9812 12764
rect 10229 12767 10287 12773
rect 8067 12733 8079 12736
rect 8021 12727 8079 12733
rect 10229 12733 10241 12767
rect 10275 12764 10287 12767
rect 10980 12764 11008 12928
rect 12066 12860 12072 12912
rect 12124 12900 12130 12912
rect 13464 12900 13492 12940
rect 12124 12872 13492 12900
rect 13541 12903 13599 12909
rect 12124 12860 12130 12872
rect 13541 12869 13553 12903
rect 13587 12869 13599 12903
rect 14016 12900 14044 12940
rect 14550 12928 14556 12980
rect 14608 12928 14614 12980
rect 17862 12928 17868 12980
rect 17920 12968 17926 12980
rect 18141 12971 18199 12977
rect 18141 12968 18153 12971
rect 17920 12940 18153 12968
rect 17920 12928 17926 12940
rect 18141 12937 18153 12940
rect 18187 12937 18199 12971
rect 18141 12931 18199 12937
rect 19886 12928 19892 12980
rect 19944 12968 19950 12980
rect 19981 12971 20039 12977
rect 19981 12968 19993 12971
rect 19944 12940 19993 12968
rect 19944 12928 19950 12940
rect 19981 12937 19993 12940
rect 20027 12937 20039 12971
rect 19981 12931 20039 12937
rect 20272 12940 22876 12968
rect 18782 12900 18788 12912
rect 14016 12872 18788 12900
rect 13541 12863 13599 12869
rect 12713 12835 12771 12841
rect 12713 12801 12725 12835
rect 12759 12832 12771 12835
rect 13078 12832 13084 12844
rect 12759 12804 13084 12832
rect 12759 12801 12771 12804
rect 12713 12795 12771 12801
rect 13078 12792 13084 12804
rect 13136 12792 13142 12844
rect 11974 12764 11980 12776
rect 10275 12736 11008 12764
rect 11748 12739 11980 12764
rect 11747 12736 11980 12739
rect 10275 12733 10287 12736
rect 10229 12727 10287 12733
rect 11747 12733 11805 12736
rect 7006 12656 7012 12708
rect 7064 12696 7070 12708
rect 7285 12699 7343 12705
rect 7285 12696 7297 12699
rect 7064 12668 7297 12696
rect 7064 12656 7070 12668
rect 7285 12665 7297 12668
rect 7331 12665 7343 12699
rect 7285 12659 7343 12665
rect 7466 12656 7472 12708
rect 7524 12656 7530 12708
rect 9585 12699 9643 12705
rect 9585 12665 9597 12699
rect 9631 12696 9643 12699
rect 10870 12696 10876 12708
rect 9631 12668 10876 12696
rect 9631 12665 9643 12668
rect 9585 12659 9643 12665
rect 10870 12656 10876 12668
rect 10928 12656 10934 12708
rect 11517 12699 11575 12705
rect 11517 12665 11529 12699
rect 11563 12696 11575 12699
rect 11606 12696 11612 12708
rect 11563 12668 11612 12696
rect 11563 12665 11575 12668
rect 11517 12659 11575 12665
rect 11606 12656 11612 12668
rect 11664 12656 11670 12708
rect 11747 12699 11759 12733
rect 11793 12699 11805 12733
rect 11974 12724 11980 12736
rect 12032 12724 12038 12776
rect 12161 12767 12219 12773
rect 12161 12733 12173 12767
rect 12207 12764 12219 12767
rect 12434 12764 12440 12776
rect 12207 12736 12440 12764
rect 12207 12733 12219 12736
rect 12161 12727 12219 12733
rect 12434 12724 12440 12736
rect 12492 12724 12498 12776
rect 12529 12767 12587 12773
rect 12529 12733 12541 12767
rect 12575 12733 12587 12767
rect 12529 12727 12587 12733
rect 12989 12767 13047 12773
rect 12989 12733 13001 12767
rect 13035 12764 13047 12767
rect 13556 12764 13584 12863
rect 18782 12860 18788 12872
rect 18840 12900 18846 12912
rect 19150 12900 19156 12912
rect 18840 12872 19156 12900
rect 18840 12860 18846 12872
rect 19150 12860 19156 12872
rect 19208 12900 19214 12912
rect 20272 12900 20300 12940
rect 19208 12872 20300 12900
rect 19208 12860 19214 12872
rect 20346 12860 20352 12912
rect 20404 12900 20410 12912
rect 20533 12903 20591 12909
rect 20533 12900 20545 12903
rect 20404 12872 20545 12900
rect 20404 12860 20410 12872
rect 20533 12869 20545 12872
rect 20579 12869 20591 12903
rect 20533 12863 20591 12869
rect 13814 12792 13820 12844
rect 13872 12832 13878 12844
rect 14093 12835 14151 12841
rect 14093 12832 14105 12835
rect 13872 12804 14105 12832
rect 13872 12792 13878 12804
rect 14093 12801 14105 12804
rect 14139 12801 14151 12835
rect 14093 12795 14151 12801
rect 14182 12792 14188 12844
rect 14240 12792 14246 12844
rect 15197 12835 15255 12841
rect 15197 12801 15209 12835
rect 15243 12832 15255 12835
rect 15746 12832 15752 12844
rect 15243 12804 15752 12832
rect 15243 12801 15255 12804
rect 15197 12795 15255 12801
rect 15746 12792 15752 12804
rect 15804 12832 15810 12844
rect 16298 12832 16304 12844
rect 15804 12804 16304 12832
rect 15804 12792 15810 12804
rect 16298 12792 16304 12804
rect 16356 12832 16362 12844
rect 16393 12835 16451 12841
rect 16393 12832 16405 12835
rect 16356 12804 16405 12832
rect 16356 12792 16362 12804
rect 16393 12801 16405 12804
rect 16439 12801 16451 12835
rect 16393 12795 16451 12801
rect 18506 12792 18512 12844
rect 18564 12792 18570 12844
rect 18874 12792 18880 12844
rect 18932 12832 18938 12844
rect 19245 12835 19303 12841
rect 19245 12832 19257 12835
rect 18932 12804 19257 12832
rect 18932 12792 18938 12804
rect 19245 12801 19257 12804
rect 19291 12801 19303 12835
rect 19245 12795 19303 12801
rect 19518 12792 19524 12844
rect 19576 12832 19582 12844
rect 20622 12832 20628 12844
rect 19576 12804 20628 12832
rect 19576 12792 19582 12804
rect 13035 12736 13584 12764
rect 14001 12767 14059 12773
rect 13035 12733 13047 12736
rect 12989 12727 13047 12733
rect 14001 12733 14013 12767
rect 14047 12764 14059 12767
rect 14200 12764 14228 12792
rect 14047 12736 14228 12764
rect 14921 12767 14979 12773
rect 14047 12733 14059 12736
rect 14001 12727 14059 12733
rect 14921 12733 14933 12767
rect 14967 12764 14979 12767
rect 15010 12764 15016 12776
rect 14967 12736 15016 12764
rect 14967 12733 14979 12736
rect 14921 12727 14979 12733
rect 11747 12693 11805 12699
rect 12544 12640 12572 12727
rect 15010 12724 15016 12736
rect 15068 12724 15074 12776
rect 16206 12724 16212 12776
rect 16264 12724 16270 12776
rect 18230 12724 18236 12776
rect 18288 12724 18294 12776
rect 18325 12767 18383 12773
rect 18325 12733 18337 12767
rect 18371 12764 18383 12767
rect 18414 12764 18420 12776
rect 18371 12736 18420 12764
rect 18371 12733 18383 12736
rect 18325 12727 18383 12733
rect 18414 12724 18420 12736
rect 18472 12724 18478 12776
rect 18693 12767 18751 12773
rect 18693 12733 18705 12767
rect 18739 12764 18751 12767
rect 19610 12764 19616 12776
rect 18739 12736 19616 12764
rect 18739 12733 18751 12736
rect 18693 12727 18751 12733
rect 13906 12656 13912 12708
rect 13964 12696 13970 12708
rect 15102 12696 15108 12708
rect 13964 12668 15108 12696
rect 13964 12656 13970 12668
rect 15102 12656 15108 12668
rect 15160 12696 15166 12708
rect 16301 12699 16359 12705
rect 15160 12668 16252 12696
rect 15160 12656 15166 12668
rect 5960 12600 6592 12628
rect 7561 12631 7619 12637
rect 5960 12588 5966 12600
rect 7561 12597 7573 12631
rect 7607 12628 7619 12631
rect 8294 12628 8300 12640
rect 7607 12600 8300 12628
rect 7607 12597 7619 12600
rect 7561 12591 7619 12597
rect 8294 12588 8300 12600
rect 8352 12588 8358 12640
rect 9214 12588 9220 12640
rect 9272 12588 9278 12640
rect 10134 12588 10140 12640
rect 10192 12588 10198 12640
rect 11974 12588 11980 12640
rect 12032 12588 12038 12640
rect 12342 12588 12348 12640
rect 12400 12588 12406 12640
rect 12526 12588 12532 12640
rect 12584 12588 12590 12640
rect 12894 12588 12900 12640
rect 12952 12628 12958 12640
rect 15013 12631 15071 12637
rect 15013 12628 15025 12631
rect 12952 12600 15025 12628
rect 12952 12588 12958 12600
rect 15013 12597 15025 12600
rect 15059 12628 15071 12631
rect 15194 12628 15200 12640
rect 15059 12600 15200 12628
rect 15059 12597 15071 12600
rect 15013 12591 15071 12597
rect 15194 12588 15200 12600
rect 15252 12588 15258 12640
rect 15838 12588 15844 12640
rect 15896 12588 15902 12640
rect 16224 12628 16252 12668
rect 16301 12665 16313 12699
rect 16347 12696 16359 12699
rect 18248 12696 18276 12724
rect 18708 12696 18736 12727
rect 19610 12724 19616 12736
rect 19668 12724 19674 12776
rect 19702 12724 19708 12776
rect 19760 12764 19766 12776
rect 20456 12773 20484 12804
rect 20622 12792 20628 12804
rect 20680 12792 20686 12844
rect 21821 12835 21879 12841
rect 21821 12832 21833 12835
rect 20916 12804 21833 12832
rect 20165 12767 20223 12773
rect 20165 12764 20177 12767
rect 19760 12736 20177 12764
rect 19760 12724 19766 12736
rect 20165 12733 20177 12736
rect 20211 12733 20223 12767
rect 20165 12727 20223 12733
rect 20441 12767 20499 12773
rect 20441 12733 20453 12767
rect 20487 12733 20499 12767
rect 20441 12727 20499 12733
rect 20530 12724 20536 12776
rect 20588 12724 20594 12776
rect 20714 12724 20720 12776
rect 20772 12724 20778 12776
rect 20916 12773 20944 12804
rect 21821 12801 21833 12804
rect 21867 12801 21879 12835
rect 21821 12795 21879 12801
rect 22066 12804 22784 12832
rect 20901 12767 20959 12773
rect 20901 12733 20913 12767
rect 20947 12733 20959 12767
rect 21269 12767 21327 12773
rect 21269 12764 21281 12767
rect 20901 12727 20959 12733
rect 21008 12736 21281 12764
rect 16347 12668 18736 12696
rect 16347 12665 16359 12668
rect 16301 12659 16359 12665
rect 18782 12656 18788 12708
rect 18840 12696 18846 12708
rect 18969 12699 19027 12705
rect 18969 12696 18981 12699
rect 18840 12668 18981 12696
rect 18840 12656 18846 12668
rect 18969 12665 18981 12668
rect 19015 12665 19027 12699
rect 20548 12696 20576 12724
rect 21008 12696 21036 12736
rect 21269 12733 21281 12736
rect 21315 12764 21327 12767
rect 22066 12764 22094 12804
rect 21315 12736 22094 12764
rect 21315 12733 21327 12736
rect 21269 12727 21327 12733
rect 22462 12724 22468 12776
rect 22520 12724 22526 12776
rect 22756 12773 22784 12804
rect 22848 12773 22876 12940
rect 23106 12928 23112 12980
rect 23164 12968 23170 12980
rect 23201 12971 23259 12977
rect 23201 12968 23213 12971
rect 23164 12940 23213 12968
rect 23164 12928 23170 12940
rect 23201 12937 23213 12940
rect 23247 12937 23259 12971
rect 23201 12931 23259 12937
rect 23842 12928 23848 12980
rect 23900 12968 23906 12980
rect 24489 12971 24547 12977
rect 24489 12968 24501 12971
rect 23900 12940 24501 12968
rect 23900 12928 23906 12940
rect 24489 12937 24501 12940
rect 24535 12937 24547 12971
rect 24489 12931 24547 12937
rect 24121 12903 24179 12909
rect 24121 12869 24133 12903
rect 24167 12900 24179 12903
rect 24302 12900 24308 12912
rect 24167 12872 24308 12900
rect 24167 12869 24179 12872
rect 24121 12863 24179 12869
rect 24302 12860 24308 12872
rect 24360 12860 24366 12912
rect 24504 12900 24532 12931
rect 24670 12928 24676 12980
rect 24728 12968 24734 12980
rect 26234 12968 26240 12980
rect 24728 12940 26240 12968
rect 24728 12928 24734 12940
rect 26234 12928 26240 12940
rect 26292 12928 26298 12980
rect 25314 12900 25320 12912
rect 24504 12872 25320 12900
rect 25314 12860 25320 12872
rect 25372 12860 25378 12912
rect 23937 12835 23995 12841
rect 23937 12801 23949 12835
rect 23983 12832 23995 12835
rect 25498 12832 25504 12844
rect 23983 12804 25504 12832
rect 23983 12801 23995 12804
rect 23937 12795 23995 12801
rect 25498 12792 25504 12804
rect 25556 12792 25562 12844
rect 26878 12792 26884 12844
rect 26936 12792 26942 12844
rect 22741 12767 22799 12773
rect 22741 12733 22753 12767
rect 22787 12733 22799 12767
rect 22741 12727 22799 12733
rect 22833 12767 22891 12773
rect 22833 12733 22845 12767
rect 22879 12733 22891 12767
rect 22833 12727 22891 12733
rect 23106 12724 23112 12776
rect 23164 12724 23170 12776
rect 23658 12724 23664 12776
rect 23716 12764 23722 12776
rect 23845 12767 23903 12773
rect 23845 12764 23857 12767
rect 23716 12736 23857 12764
rect 23716 12724 23722 12736
rect 23845 12733 23857 12736
rect 23891 12733 23903 12767
rect 23845 12727 23903 12733
rect 24029 12767 24087 12773
rect 24029 12733 24041 12767
rect 24075 12764 24087 12767
rect 25222 12764 25228 12776
rect 24075 12736 25228 12764
rect 24075 12733 24087 12736
rect 24029 12727 24087 12733
rect 25222 12724 25228 12736
rect 25280 12724 25286 12776
rect 25314 12724 25320 12776
rect 25372 12724 25378 12776
rect 18969 12659 19027 12665
rect 19812 12668 20484 12696
rect 20548 12668 21036 12696
rect 19812 12628 19840 12668
rect 16224 12600 19840 12628
rect 19889 12631 19947 12637
rect 19889 12597 19901 12631
rect 19935 12628 19947 12631
rect 20349 12631 20407 12637
rect 20349 12628 20361 12631
rect 19935 12600 20361 12628
rect 19935 12597 19947 12600
rect 19889 12591 19947 12597
rect 20349 12597 20361 12600
rect 20395 12597 20407 12631
rect 20456 12628 20484 12668
rect 21082 12656 21088 12708
rect 21140 12656 21146 12708
rect 21174 12656 21180 12708
rect 21232 12656 21238 12708
rect 22925 12699 22983 12705
rect 21284 12668 22692 12696
rect 20990 12628 20996 12640
rect 20456 12600 20996 12628
rect 20349 12591 20407 12597
rect 20990 12588 20996 12600
rect 21048 12588 21054 12640
rect 21100 12628 21128 12656
rect 21284 12628 21312 12668
rect 21100 12600 21312 12628
rect 21450 12588 21456 12640
rect 21508 12588 21514 12640
rect 22554 12588 22560 12640
rect 22612 12588 22618 12640
rect 22664 12628 22692 12668
rect 22925 12665 22937 12699
rect 22971 12665 22983 12699
rect 22925 12659 22983 12665
rect 22940 12628 22968 12659
rect 23382 12656 23388 12708
rect 23440 12656 23446 12708
rect 23566 12656 23572 12708
rect 23624 12656 23630 12708
rect 24946 12696 24952 12708
rect 24504 12668 24952 12696
rect 24504 12637 24532 12668
rect 24946 12656 24952 12668
rect 25004 12656 25010 12708
rect 26602 12656 26608 12708
rect 26660 12705 26666 12708
rect 26660 12659 26672 12705
rect 26660 12656 26666 12659
rect 22664 12600 22968 12628
rect 24489 12631 24547 12637
rect 24489 12597 24501 12631
rect 24535 12597 24547 12631
rect 24489 12591 24547 12597
rect 24670 12588 24676 12640
rect 24728 12588 24734 12640
rect 24762 12588 24768 12640
rect 24820 12588 24826 12640
rect 25038 12588 25044 12640
rect 25096 12628 25102 12640
rect 25501 12631 25559 12637
rect 25501 12628 25513 12631
rect 25096 12600 25513 12628
rect 25096 12588 25102 12600
rect 25501 12597 25513 12600
rect 25547 12597 25559 12631
rect 25501 12591 25559 12597
rect 552 12538 27576 12560
rect 552 12486 7114 12538
rect 7166 12486 7178 12538
rect 7230 12486 7242 12538
rect 7294 12486 7306 12538
rect 7358 12486 7370 12538
rect 7422 12486 13830 12538
rect 13882 12486 13894 12538
rect 13946 12486 13958 12538
rect 14010 12486 14022 12538
rect 14074 12486 14086 12538
rect 14138 12486 20546 12538
rect 20598 12486 20610 12538
rect 20662 12486 20674 12538
rect 20726 12486 20738 12538
rect 20790 12486 20802 12538
rect 20854 12486 27262 12538
rect 27314 12486 27326 12538
rect 27378 12486 27390 12538
rect 27442 12486 27454 12538
rect 27506 12486 27518 12538
rect 27570 12486 27576 12538
rect 552 12464 27576 12486
rect 1397 12427 1455 12433
rect 1397 12393 1409 12427
rect 1443 12424 1455 12427
rect 1946 12424 1952 12436
rect 1443 12396 1952 12424
rect 1443 12393 1455 12396
rect 1397 12387 1455 12393
rect 1946 12384 1952 12396
rect 2004 12384 2010 12436
rect 2774 12384 2780 12436
rect 2832 12424 2838 12436
rect 2869 12427 2927 12433
rect 2869 12424 2881 12427
rect 2832 12396 2881 12424
rect 2832 12384 2838 12396
rect 2869 12393 2881 12396
rect 2915 12393 2927 12427
rect 2869 12387 2927 12393
rect 3234 12384 3240 12436
rect 3292 12384 3298 12436
rect 3421 12427 3479 12433
rect 3421 12393 3433 12427
rect 3467 12424 3479 12427
rect 4154 12424 4160 12436
rect 3467 12396 4160 12424
rect 3467 12393 3479 12396
rect 3421 12387 3479 12393
rect 4154 12384 4160 12396
rect 4212 12384 4218 12436
rect 7742 12384 7748 12436
rect 7800 12384 7806 12436
rect 10134 12384 10140 12436
rect 10192 12384 10198 12436
rect 11974 12424 11980 12436
rect 11440 12396 11980 12424
rect 3252 12356 3280 12384
rect 1872 12328 3280 12356
rect 1026 12248 1032 12300
rect 1084 12248 1090 12300
rect 1213 12291 1271 12297
rect 1213 12257 1225 12291
rect 1259 12257 1271 12291
rect 1213 12251 1271 12257
rect 1489 12291 1547 12297
rect 1489 12257 1501 12291
rect 1535 12257 1547 12291
rect 1489 12251 1547 12257
rect 1228 12152 1256 12251
rect 1504 12220 1532 12251
rect 1670 12248 1676 12300
rect 1728 12248 1734 12300
rect 1762 12248 1768 12300
rect 1820 12248 1826 12300
rect 1872 12297 1900 12328
rect 3510 12316 3516 12368
rect 3568 12316 3574 12368
rect 3780 12359 3838 12365
rect 3780 12325 3792 12359
rect 3826 12356 3838 12359
rect 3970 12356 3976 12368
rect 3826 12328 3976 12356
rect 3826 12325 3838 12328
rect 3780 12319 3838 12325
rect 3970 12316 3976 12328
rect 4028 12316 4034 12368
rect 5629 12359 5687 12365
rect 5092 12328 5304 12356
rect 1857 12291 1915 12297
rect 1857 12257 1869 12291
rect 1903 12257 1915 12291
rect 2498 12288 2504 12300
rect 1857 12251 1915 12257
rect 1964 12260 2504 12288
rect 1964 12220 1992 12260
rect 2498 12248 2504 12260
rect 2556 12248 2562 12300
rect 2958 12248 2964 12300
rect 3016 12248 3022 12300
rect 3142 12248 3148 12300
rect 3200 12248 3206 12300
rect 3237 12291 3295 12297
rect 3237 12257 3249 12291
rect 3283 12257 3295 12291
rect 3528 12288 3556 12316
rect 5092 12300 5120 12328
rect 3237 12251 3295 12257
rect 3344 12260 3556 12288
rect 1504 12192 1992 12220
rect 2133 12223 2191 12229
rect 2133 12189 2145 12223
rect 2179 12220 2191 12223
rect 2225 12223 2283 12229
rect 2225 12220 2237 12223
rect 2179 12192 2237 12220
rect 2179 12189 2191 12192
rect 2133 12183 2191 12189
rect 2225 12189 2237 12192
rect 2271 12189 2283 12223
rect 2225 12183 2283 12189
rect 2774 12180 2780 12232
rect 2832 12220 2838 12232
rect 3252 12220 3280 12251
rect 2832 12192 3280 12220
rect 2832 12180 2838 12192
rect 3344 12152 3372 12260
rect 4982 12248 4988 12300
rect 5040 12248 5046 12300
rect 5074 12248 5080 12300
rect 5132 12248 5138 12300
rect 5276 12297 5304 12328
rect 5629 12325 5641 12359
rect 5675 12356 5687 12359
rect 7294 12359 7352 12365
rect 7294 12356 7306 12359
rect 5675 12328 7306 12356
rect 5675 12325 5687 12328
rect 5629 12319 5687 12325
rect 7294 12325 7306 12328
rect 7340 12325 7352 12359
rect 7294 12319 7352 12325
rect 8757 12359 8815 12365
rect 8757 12325 8769 12359
rect 8803 12356 8815 12359
rect 8938 12356 8944 12368
rect 8803 12328 8944 12356
rect 8803 12325 8815 12328
rect 8757 12319 8815 12325
rect 8938 12316 8944 12328
rect 8996 12316 9002 12368
rect 9674 12356 9680 12368
rect 9140 12328 9680 12356
rect 9140 12300 9168 12328
rect 9674 12316 9680 12328
rect 9732 12316 9738 12368
rect 11324 12359 11382 12365
rect 11324 12325 11336 12359
rect 11370 12356 11382 12359
rect 11440 12356 11468 12396
rect 11974 12384 11980 12396
rect 12032 12384 12038 12436
rect 14734 12384 14740 12436
rect 14792 12384 14798 12436
rect 15473 12427 15531 12433
rect 15473 12393 15485 12427
rect 15519 12393 15531 12427
rect 15473 12387 15531 12393
rect 11370 12328 11468 12356
rect 11370 12325 11382 12328
rect 11324 12319 11382 12325
rect 11514 12316 11520 12368
rect 11572 12356 11578 12368
rect 12713 12359 12771 12365
rect 12713 12356 12725 12359
rect 11572 12328 12725 12356
rect 11572 12316 11578 12328
rect 12713 12325 12725 12328
rect 12759 12325 12771 12359
rect 12713 12319 12771 12325
rect 14461 12359 14519 12365
rect 14461 12325 14473 12359
rect 14507 12356 14519 12359
rect 14752 12356 14780 12384
rect 14507 12328 14780 12356
rect 15488 12356 15516 12387
rect 15654 12384 15660 12436
rect 15712 12424 15718 12436
rect 15838 12424 15844 12436
rect 15712 12396 15844 12424
rect 15712 12384 15718 12396
rect 15838 12384 15844 12396
rect 15896 12384 15902 12436
rect 15933 12427 15991 12433
rect 15933 12393 15945 12427
rect 15979 12424 15991 12427
rect 16206 12424 16212 12436
rect 15979 12396 16212 12424
rect 15979 12393 15991 12396
rect 15933 12387 15991 12393
rect 16206 12384 16212 12396
rect 16264 12384 16270 12436
rect 19610 12384 19616 12436
rect 19668 12384 19674 12436
rect 20717 12427 20775 12433
rect 20717 12393 20729 12427
rect 20763 12424 20775 12427
rect 20898 12424 20904 12436
rect 20763 12396 20904 12424
rect 20763 12393 20775 12396
rect 20717 12387 20775 12393
rect 20898 12384 20904 12396
rect 20956 12384 20962 12436
rect 22002 12424 22008 12436
rect 21008 12396 22008 12424
rect 17230 12359 17288 12365
rect 17230 12356 17242 12359
rect 15488 12328 17242 12356
rect 14507 12325 14519 12328
rect 14461 12319 14519 12325
rect 17230 12325 17242 12328
rect 17276 12325 17288 12359
rect 17230 12319 17288 12325
rect 5169 12291 5227 12297
rect 5169 12257 5181 12291
rect 5215 12257 5227 12291
rect 5169 12251 5227 12257
rect 5261 12291 5319 12297
rect 5261 12257 5273 12291
rect 5307 12257 5319 12291
rect 5261 12251 5319 12257
rect 5353 12291 5411 12297
rect 5353 12257 5365 12291
rect 5399 12288 5411 12291
rect 7006 12288 7012 12300
rect 5399 12260 7012 12288
rect 5399 12257 5411 12260
rect 5353 12251 5411 12257
rect 3513 12223 3571 12229
rect 3513 12189 3525 12223
rect 3559 12189 3571 12223
rect 3513 12183 3571 12189
rect 1228 12124 3372 12152
rect 1118 12044 1124 12096
rect 1176 12084 1182 12096
rect 2961 12087 3019 12093
rect 2961 12084 2973 12087
rect 1176 12056 2973 12084
rect 1176 12044 1182 12056
rect 2961 12053 2973 12056
rect 3007 12053 3019 12087
rect 3528 12084 3556 12183
rect 5000 12152 5028 12248
rect 5184 12220 5212 12251
rect 7006 12248 7012 12260
rect 7064 12248 7070 12300
rect 7650 12248 7656 12300
rect 7708 12248 7714 12300
rect 8202 12248 8208 12300
rect 8260 12248 8266 12300
rect 8294 12248 8300 12300
rect 8352 12248 8358 12300
rect 8478 12248 8484 12300
rect 8536 12248 8542 12300
rect 8662 12248 8668 12300
rect 8720 12288 8726 12300
rect 8849 12291 8907 12297
rect 8849 12288 8861 12291
rect 8720 12260 8861 12288
rect 8720 12248 8726 12260
rect 8849 12257 8861 12260
rect 8895 12257 8907 12291
rect 8849 12251 8907 12257
rect 9033 12291 9091 12297
rect 9033 12257 9045 12291
rect 9079 12257 9091 12291
rect 9033 12251 9091 12257
rect 6546 12220 6552 12232
rect 5184 12192 6552 12220
rect 6546 12180 6552 12192
rect 6604 12180 6610 12232
rect 7558 12180 7564 12232
rect 7616 12220 7622 12232
rect 8220 12220 8248 12248
rect 7616 12192 8248 12220
rect 7616 12180 7622 12192
rect 5000 12124 5488 12152
rect 5460 12096 5488 12124
rect 4430 12084 4436 12096
rect 3528 12056 4436 12084
rect 2961 12047 3019 12053
rect 4430 12044 4436 12056
rect 4488 12044 4494 12096
rect 4798 12044 4804 12096
rect 4856 12084 4862 12096
rect 4893 12087 4951 12093
rect 4893 12084 4905 12087
rect 4856 12056 4905 12084
rect 4856 12044 4862 12056
rect 4893 12053 4905 12056
rect 4939 12053 4951 12087
rect 4893 12047 4951 12053
rect 5442 12044 5448 12096
rect 5500 12044 5506 12096
rect 6181 12087 6239 12093
rect 6181 12053 6193 12087
rect 6227 12084 6239 12087
rect 6454 12084 6460 12096
rect 6227 12056 6460 12084
rect 6227 12053 6239 12056
rect 6181 12047 6239 12053
rect 6454 12044 6460 12056
rect 6512 12084 6518 12096
rect 6822 12084 6828 12096
rect 6512 12056 6828 12084
rect 6512 12044 6518 12056
rect 6822 12044 6828 12056
rect 6880 12044 6886 12096
rect 8864 12084 8892 12251
rect 9048 12220 9076 12251
rect 9122 12248 9128 12300
rect 9180 12248 9186 12300
rect 9306 12248 9312 12300
rect 9364 12248 9370 12300
rect 9692 12220 9720 12316
rect 10781 12291 10839 12297
rect 10781 12288 10793 12291
rect 10520 12260 10793 12288
rect 9861 12223 9919 12229
rect 9861 12220 9873 12223
rect 9048 12192 9352 12220
rect 9692 12192 9873 12220
rect 9324 12096 9352 12192
rect 9861 12189 9873 12192
rect 9907 12189 9919 12223
rect 9861 12183 9919 12189
rect 10042 12180 10048 12232
rect 10100 12180 10106 12232
rect 10520 12161 10548 12260
rect 10781 12257 10793 12260
rect 10827 12257 10839 12291
rect 10781 12251 10839 12257
rect 11054 12248 11060 12300
rect 11112 12288 11118 12300
rect 11882 12288 11888 12300
rect 11112 12260 11888 12288
rect 11112 12248 11118 12260
rect 11882 12248 11888 12260
rect 11940 12288 11946 12300
rect 14476 12288 14504 12319
rect 20254 12316 20260 12368
rect 20312 12356 20318 12368
rect 21008 12356 21036 12396
rect 22002 12384 22008 12396
rect 22060 12384 22066 12436
rect 22462 12384 22468 12436
rect 22520 12424 22526 12436
rect 22649 12427 22707 12433
rect 22649 12424 22661 12427
rect 22520 12396 22661 12424
rect 22520 12384 22526 12396
rect 22649 12393 22661 12396
rect 22695 12424 22707 12427
rect 22922 12424 22928 12436
rect 22695 12396 22928 12424
rect 22695 12393 22707 12396
rect 22649 12387 22707 12393
rect 22922 12384 22928 12396
rect 22980 12384 22986 12436
rect 23106 12384 23112 12436
rect 23164 12424 23170 12436
rect 23385 12427 23443 12433
rect 23385 12424 23397 12427
rect 23164 12396 23397 12424
rect 23164 12384 23170 12396
rect 23385 12393 23397 12396
rect 23431 12393 23443 12427
rect 23845 12427 23903 12433
rect 23845 12424 23857 12427
rect 23385 12387 23443 12393
rect 23584 12396 23857 12424
rect 21542 12365 21548 12368
rect 20312 12328 21036 12356
rect 21514 12359 21548 12365
rect 20312 12316 20318 12328
rect 21514 12325 21526 12359
rect 21514 12319 21548 12325
rect 21542 12316 21548 12319
rect 21600 12316 21606 12368
rect 23584 12356 23612 12396
rect 23845 12393 23857 12396
rect 23891 12393 23903 12427
rect 23845 12387 23903 12393
rect 25314 12384 25320 12436
rect 25372 12424 25378 12436
rect 26237 12427 26295 12433
rect 26237 12424 26249 12427
rect 25372 12396 26249 12424
rect 25372 12384 25378 12396
rect 26237 12393 26249 12396
rect 26283 12393 26295 12427
rect 26237 12387 26295 12393
rect 26602 12384 26608 12436
rect 26660 12384 26666 12436
rect 23400 12328 23612 12356
rect 11940 12260 14504 12288
rect 11940 12248 11946 12260
rect 14550 12248 14556 12300
rect 14608 12248 14614 12300
rect 14737 12291 14795 12297
rect 14737 12257 14749 12291
rect 14783 12257 14795 12291
rect 14737 12251 14795 12257
rect 10505 12155 10563 12161
rect 10505 12121 10517 12155
rect 10551 12121 10563 12155
rect 14752 12152 14780 12251
rect 14826 12248 14832 12300
rect 14884 12248 14890 12300
rect 15289 12291 15347 12297
rect 15289 12257 15301 12291
rect 15335 12288 15347 12291
rect 15654 12288 15660 12300
rect 15335 12260 15660 12288
rect 15335 12257 15347 12260
rect 15289 12251 15347 12257
rect 15654 12248 15660 12260
rect 15712 12248 15718 12300
rect 15749 12291 15807 12297
rect 15749 12257 15761 12291
rect 15795 12257 15807 12291
rect 15749 12251 15807 12257
rect 14844 12220 14872 12248
rect 15565 12223 15623 12229
rect 15565 12220 15577 12223
rect 14844 12192 15577 12220
rect 15565 12189 15577 12192
rect 15611 12189 15623 12223
rect 15565 12183 15623 12189
rect 15764 12152 15792 12251
rect 16666 12248 16672 12300
rect 16724 12288 16730 12300
rect 17954 12297 17960 12300
rect 16724 12260 17540 12288
rect 16724 12248 16730 12260
rect 17512 12229 17540 12260
rect 17948 12251 17960 12297
rect 17954 12248 17960 12251
rect 18012 12248 18018 12300
rect 19518 12248 19524 12300
rect 19576 12248 19582 12300
rect 19794 12248 19800 12300
rect 19852 12288 19858 12300
rect 20349 12291 20407 12297
rect 20349 12288 20361 12291
rect 19852 12260 20361 12288
rect 19852 12248 19858 12260
rect 20349 12257 20361 12260
rect 20395 12257 20407 12291
rect 20349 12251 20407 12257
rect 21266 12248 21272 12300
rect 21324 12248 21330 12300
rect 17497 12223 17555 12229
rect 17497 12189 17509 12223
rect 17543 12220 17555 12223
rect 17681 12223 17739 12229
rect 17681 12220 17693 12223
rect 17543 12192 17693 12220
rect 17543 12189 17555 12192
rect 17497 12183 17555 12189
rect 17681 12189 17693 12192
rect 17727 12189 17739 12223
rect 19705 12223 19763 12229
rect 19705 12220 19717 12223
rect 17681 12183 17739 12189
rect 18708 12192 19717 12220
rect 16117 12155 16175 12161
rect 16117 12152 16129 12155
rect 14752 12124 16129 12152
rect 10505 12115 10563 12121
rect 16117 12121 16129 12124
rect 16163 12121 16175 12155
rect 16117 12115 16175 12121
rect 9125 12087 9183 12093
rect 9125 12084 9137 12087
rect 8864 12056 9137 12084
rect 9125 12053 9137 12056
rect 9171 12053 9183 12087
rect 9125 12047 9183 12053
rect 9306 12044 9312 12096
rect 9364 12044 9370 12096
rect 9582 12044 9588 12096
rect 9640 12044 9646 12096
rect 10318 12044 10324 12096
rect 10376 12084 10382 12096
rect 10597 12087 10655 12093
rect 10597 12084 10609 12087
rect 10376 12056 10609 12084
rect 10376 12044 10382 12056
rect 10597 12053 10609 12056
rect 10643 12053 10655 12087
rect 10597 12047 10655 12053
rect 12437 12087 12495 12093
rect 12437 12053 12449 12087
rect 12483 12084 12495 12087
rect 12526 12084 12532 12096
rect 12483 12056 12532 12084
rect 12483 12053 12495 12056
rect 12437 12047 12495 12053
rect 12526 12044 12532 12056
rect 12584 12084 12590 12096
rect 13354 12084 13360 12096
rect 12584 12056 13360 12084
rect 12584 12044 12590 12056
rect 13354 12044 13360 12056
rect 13412 12044 13418 12096
rect 14366 12044 14372 12096
rect 14424 12084 14430 12096
rect 14553 12087 14611 12093
rect 14553 12084 14565 12087
rect 14424 12056 14565 12084
rect 14424 12044 14430 12056
rect 14553 12053 14565 12056
rect 14599 12053 14611 12087
rect 14553 12047 14611 12053
rect 17678 12044 17684 12096
rect 17736 12084 17742 12096
rect 18708 12084 18736 12192
rect 19705 12189 19717 12192
rect 19751 12220 19763 12223
rect 19978 12220 19984 12232
rect 19751 12192 19984 12220
rect 19751 12189 19763 12192
rect 19705 12183 19763 12189
rect 19978 12180 19984 12192
rect 20036 12220 20042 12232
rect 20073 12223 20131 12229
rect 20073 12220 20085 12223
rect 20036 12192 20085 12220
rect 20036 12180 20042 12192
rect 20073 12189 20085 12192
rect 20119 12189 20131 12223
rect 20073 12183 20131 12189
rect 22830 12180 22836 12232
rect 22888 12180 22894 12232
rect 23400 12096 23428 12328
rect 23658 12316 23664 12368
rect 23716 12356 23722 12368
rect 25958 12356 25964 12368
rect 23716 12328 25964 12356
rect 23716 12316 23722 12328
rect 23842 12288 23848 12300
rect 23584 12260 23848 12288
rect 23584 12232 23612 12260
rect 23842 12248 23848 12260
rect 23900 12248 23906 12300
rect 24872 12297 24900 12328
rect 25958 12316 25964 12328
rect 26016 12356 26022 12368
rect 26878 12356 26884 12368
rect 26016 12328 26884 12356
rect 26016 12316 26022 12328
rect 26878 12316 26884 12328
rect 26936 12316 26942 12368
rect 23937 12291 23995 12297
rect 23937 12257 23949 12291
rect 23983 12288 23995 12291
rect 24857 12291 24915 12297
rect 23983 12260 24716 12288
rect 23983 12257 23995 12260
rect 23937 12251 23995 12257
rect 23477 12223 23535 12229
rect 23477 12189 23489 12223
rect 23523 12220 23535 12223
rect 23566 12220 23572 12232
rect 23523 12192 23572 12220
rect 23523 12189 23535 12192
rect 23477 12183 23535 12189
rect 23566 12180 23572 12192
rect 23624 12180 23630 12232
rect 23661 12223 23719 12229
rect 23661 12189 23673 12223
rect 23707 12220 23719 12223
rect 24581 12223 24639 12229
rect 24581 12220 24593 12223
rect 23707 12192 24593 12220
rect 23707 12189 23719 12192
rect 23661 12183 23719 12189
rect 24581 12189 24593 12192
rect 24627 12189 24639 12223
rect 24581 12183 24639 12189
rect 24688 12152 24716 12260
rect 24857 12257 24869 12291
rect 24903 12257 24915 12291
rect 25113 12291 25171 12297
rect 25113 12288 25125 12291
rect 24857 12251 24915 12257
rect 24964 12260 25125 12288
rect 24762 12180 24768 12232
rect 24820 12220 24826 12232
rect 24964 12220 24992 12260
rect 25113 12257 25125 12260
rect 25159 12257 25171 12291
rect 25113 12251 25171 12257
rect 26418 12248 26424 12300
rect 26476 12248 26482 12300
rect 24820 12192 24992 12220
rect 24820 12180 24826 12192
rect 24688 12124 24900 12152
rect 24872 12096 24900 12124
rect 17736 12056 18736 12084
rect 17736 12044 17742 12056
rect 19058 12044 19064 12096
rect 19116 12044 19122 12096
rect 19150 12044 19156 12096
rect 19208 12044 19214 12096
rect 23382 12044 23388 12096
rect 23440 12044 23446 12096
rect 23750 12044 23756 12096
rect 23808 12084 23814 12096
rect 24029 12087 24087 12093
rect 24029 12084 24041 12087
rect 23808 12056 24041 12084
rect 23808 12044 23814 12056
rect 24029 12053 24041 12056
rect 24075 12053 24087 12087
rect 24029 12047 24087 12053
rect 24854 12044 24860 12096
rect 24912 12044 24918 12096
rect 552 11994 27416 12016
rect 552 11942 3756 11994
rect 3808 11942 3820 11994
rect 3872 11942 3884 11994
rect 3936 11942 3948 11994
rect 4000 11942 4012 11994
rect 4064 11942 10472 11994
rect 10524 11942 10536 11994
rect 10588 11942 10600 11994
rect 10652 11942 10664 11994
rect 10716 11942 10728 11994
rect 10780 11942 17188 11994
rect 17240 11942 17252 11994
rect 17304 11942 17316 11994
rect 17368 11942 17380 11994
rect 17432 11942 17444 11994
rect 17496 11942 23904 11994
rect 23956 11942 23968 11994
rect 24020 11942 24032 11994
rect 24084 11942 24096 11994
rect 24148 11942 24160 11994
rect 24212 11942 27416 11994
rect 552 11920 27416 11942
rect 3326 11880 3332 11892
rect 1412 11852 3332 11880
rect 1210 11636 1216 11688
rect 1268 11636 1274 11688
rect 1412 11685 1440 11852
rect 3326 11840 3332 11852
rect 3384 11880 3390 11892
rect 4062 11880 4068 11892
rect 3384 11852 4068 11880
rect 3384 11840 3390 11852
rect 4062 11840 4068 11852
rect 4120 11880 4126 11892
rect 7466 11880 7472 11892
rect 4120 11852 7472 11880
rect 4120 11840 4126 11852
rect 7466 11840 7472 11852
rect 7524 11840 7530 11892
rect 8478 11840 8484 11892
rect 8536 11880 8542 11892
rect 9125 11883 9183 11889
rect 9125 11880 9137 11883
rect 8536 11852 9137 11880
rect 8536 11840 8542 11852
rect 9125 11849 9137 11852
rect 9171 11849 9183 11883
rect 9125 11843 9183 11849
rect 12434 11840 12440 11892
rect 12492 11840 12498 11892
rect 13722 11840 13728 11892
rect 13780 11840 13786 11892
rect 17954 11840 17960 11892
rect 18012 11840 18018 11892
rect 19061 11883 19119 11889
rect 19061 11849 19073 11883
rect 19107 11880 19119 11883
rect 19518 11880 19524 11892
rect 19107 11852 19524 11880
rect 19107 11849 19119 11852
rect 19061 11843 19119 11849
rect 19518 11840 19524 11852
rect 19576 11840 19582 11892
rect 21266 11880 21272 11892
rect 21100 11852 21272 11880
rect 2682 11812 2688 11824
rect 1872 11784 2688 11812
rect 1397 11679 1455 11685
rect 1397 11645 1409 11679
rect 1443 11645 1455 11679
rect 1397 11639 1455 11645
rect 1762 11636 1768 11688
rect 1820 11636 1826 11688
rect 1872 11685 1900 11784
rect 2682 11772 2688 11784
rect 2740 11772 2746 11824
rect 2958 11772 2964 11824
rect 3016 11772 3022 11824
rect 4341 11815 4399 11821
rect 4341 11812 4353 11815
rect 4080 11784 4353 11812
rect 2869 11747 2927 11753
rect 2869 11713 2881 11747
rect 2915 11744 2927 11747
rect 2976 11744 3004 11772
rect 2915 11716 3004 11744
rect 2915 11713 2927 11716
rect 2869 11707 2927 11713
rect 1857 11679 1915 11685
rect 1857 11645 1869 11679
rect 1903 11645 1915 11679
rect 1857 11639 1915 11645
rect 1949 11679 2007 11685
rect 1949 11645 1961 11679
rect 1995 11676 2007 11679
rect 2133 11679 2191 11685
rect 1995 11648 2084 11676
rect 1995 11645 2007 11648
rect 1949 11639 2007 11645
rect 1029 11611 1087 11617
rect 1029 11577 1041 11611
rect 1075 11608 1087 11611
rect 1075 11580 1900 11608
rect 1075 11577 1087 11580
rect 1029 11571 1087 11577
rect 1486 11500 1492 11552
rect 1544 11500 1550 11552
rect 1872 11540 1900 11580
rect 2056 11540 2084 11648
rect 2133 11645 2145 11679
rect 2179 11676 2191 11679
rect 2498 11676 2504 11688
rect 2179 11648 2504 11676
rect 2179 11645 2191 11648
rect 2133 11639 2191 11645
rect 2498 11636 2504 11648
rect 2556 11636 2562 11688
rect 2682 11636 2688 11688
rect 2740 11676 2746 11688
rect 4080 11676 4108 11784
rect 4341 11781 4353 11784
rect 4387 11812 4399 11815
rect 4982 11812 4988 11824
rect 4387 11784 4988 11812
rect 4387 11781 4399 11784
rect 4341 11775 4399 11781
rect 4982 11772 4988 11784
rect 5040 11772 5046 11824
rect 8205 11815 8263 11821
rect 8205 11781 8217 11815
rect 8251 11812 8263 11815
rect 8251 11784 9720 11812
rect 8251 11781 8263 11784
rect 8205 11775 8263 11781
rect 4430 11704 4436 11756
rect 4488 11744 4494 11756
rect 4890 11744 4896 11756
rect 4488 11716 4896 11744
rect 4488 11704 4494 11716
rect 4890 11704 4896 11716
rect 4948 11744 4954 11756
rect 9692 11753 9720 11784
rect 11900 11784 13216 11812
rect 5353 11747 5411 11753
rect 5353 11744 5365 11747
rect 4948 11716 5365 11744
rect 4948 11704 4954 11716
rect 5353 11713 5365 11716
rect 5399 11713 5411 11747
rect 5353 11707 5411 11713
rect 9677 11747 9735 11753
rect 9677 11713 9689 11747
rect 9723 11713 9735 11747
rect 9677 11707 9735 11713
rect 11054 11704 11060 11756
rect 11112 11704 11118 11756
rect 11900 11753 11928 11784
rect 11885 11747 11943 11753
rect 11885 11713 11897 11747
rect 11931 11713 11943 11747
rect 11885 11707 11943 11713
rect 11977 11747 12035 11753
rect 11977 11713 11989 11747
rect 12023 11744 12035 11747
rect 12342 11744 12348 11756
rect 12023 11716 12348 11744
rect 12023 11713 12035 11716
rect 11977 11707 12035 11713
rect 12342 11704 12348 11716
rect 12400 11704 12406 11756
rect 13188 11753 13216 11784
rect 13173 11747 13231 11753
rect 13173 11713 13185 11747
rect 13219 11744 13231 11747
rect 13740 11744 13768 11840
rect 15197 11815 15255 11821
rect 15197 11781 15209 11815
rect 15243 11781 15255 11815
rect 19150 11812 19156 11824
rect 15197 11775 15255 11781
rect 18156 11784 19156 11812
rect 13219 11716 13768 11744
rect 13219 11713 13231 11716
rect 13173 11707 13231 11713
rect 14734 11704 14740 11756
rect 14792 11704 14798 11756
rect 2740 11648 4108 11676
rect 4157 11679 4215 11685
rect 2740 11636 2746 11648
rect 4157 11645 4169 11679
rect 4203 11645 4215 11679
rect 4157 11639 4215 11645
rect 4172 11552 4200 11639
rect 4522 11636 4528 11688
rect 4580 11636 4586 11688
rect 4614 11636 4620 11688
rect 4672 11636 4678 11688
rect 6825 11679 6883 11685
rect 6825 11645 6837 11679
rect 6871 11676 6883 11679
rect 7558 11676 7564 11688
rect 6871 11648 7564 11676
rect 6871 11645 6883 11648
rect 6825 11639 6883 11645
rect 7558 11636 7564 11648
rect 7616 11636 7622 11688
rect 8665 11679 8723 11685
rect 8665 11645 8677 11679
rect 8711 11645 8723 11679
rect 8665 11639 8723 11645
rect 5261 11611 5319 11617
rect 5261 11577 5273 11611
rect 5307 11608 5319 11611
rect 5598 11611 5656 11617
rect 5598 11608 5610 11611
rect 5307 11580 5610 11608
rect 5307 11577 5319 11580
rect 5261 11571 5319 11577
rect 5598 11577 5610 11580
rect 5644 11577 5656 11611
rect 5598 11571 5656 11577
rect 7092 11611 7150 11617
rect 7092 11577 7104 11611
rect 7138 11608 7150 11611
rect 7742 11608 7748 11620
rect 7138 11580 7748 11608
rect 7138 11577 7150 11580
rect 7092 11571 7150 11577
rect 7742 11568 7748 11580
rect 7800 11568 7806 11620
rect 8680 11608 8708 11639
rect 8754 11636 8760 11688
rect 8812 11636 8818 11688
rect 8846 11636 8852 11688
rect 8904 11636 8910 11688
rect 9033 11679 9091 11685
rect 9033 11645 9045 11679
rect 9079 11676 9091 11679
rect 9122 11676 9128 11688
rect 9079 11648 9128 11676
rect 9079 11645 9091 11648
rect 9033 11639 9091 11645
rect 9122 11636 9128 11648
rect 9180 11636 9186 11688
rect 9306 11636 9312 11688
rect 9364 11636 9370 11688
rect 9953 11679 10011 11685
rect 9953 11645 9965 11679
rect 9999 11676 10011 11679
rect 11072 11676 11100 11704
rect 9999 11648 11100 11676
rect 11425 11679 11483 11685
rect 9999 11645 10011 11648
rect 9953 11639 10011 11645
rect 11425 11645 11437 11679
rect 11471 11645 11483 11679
rect 11425 11639 11483 11645
rect 9324 11608 9352 11636
rect 8680 11580 9352 11608
rect 10220 11611 10278 11617
rect 10220 11577 10232 11611
rect 10266 11608 10278 11611
rect 10318 11608 10324 11620
rect 10266 11580 10324 11608
rect 10266 11577 10278 11580
rect 10220 11571 10278 11577
rect 10318 11568 10324 11580
rect 10376 11568 10382 11620
rect 11440 11608 11468 11639
rect 12066 11636 12072 11688
rect 12124 11636 12130 11688
rect 12894 11636 12900 11688
rect 12952 11636 12958 11688
rect 13725 11679 13783 11685
rect 13725 11645 13737 11679
rect 13771 11676 13783 11679
rect 14458 11676 14464 11688
rect 13771 11648 14464 11676
rect 13771 11645 13783 11648
rect 13725 11639 13783 11645
rect 14458 11636 14464 11648
rect 14516 11676 14522 11688
rect 14752 11676 14780 11704
rect 15212 11676 15240 11775
rect 15746 11704 15752 11756
rect 15804 11704 15810 11756
rect 16942 11704 16948 11756
rect 17000 11744 17006 11756
rect 17589 11747 17647 11753
rect 17589 11744 17601 11747
rect 17000 11716 17601 11744
rect 17000 11704 17006 11716
rect 17589 11713 17601 11716
rect 17635 11744 17647 11747
rect 17678 11744 17684 11756
rect 17635 11716 17684 11744
rect 17635 11713 17647 11716
rect 17589 11707 17647 11713
rect 17678 11704 17684 11716
rect 17736 11704 17742 11756
rect 14516 11648 14780 11676
rect 14844 11648 15240 11676
rect 15657 11679 15715 11685
rect 14516 11636 14522 11648
rect 13992 11611 14050 11617
rect 11440 11580 12434 11608
rect 1872 11512 2084 11540
rect 2130 11500 2136 11552
rect 2188 11540 2194 11552
rect 2225 11543 2283 11549
rect 2225 11540 2237 11543
rect 2188 11512 2237 11540
rect 2188 11500 2194 11512
rect 2225 11509 2237 11512
rect 2271 11540 2283 11543
rect 2774 11540 2780 11552
rect 2271 11512 2780 11540
rect 2271 11509 2283 11512
rect 2225 11503 2283 11509
rect 2774 11500 2780 11512
rect 2832 11500 2838 11552
rect 3234 11500 3240 11552
rect 3292 11540 3298 11552
rect 3513 11543 3571 11549
rect 3513 11540 3525 11543
rect 3292 11512 3525 11540
rect 3292 11500 3298 11512
rect 3513 11509 3525 11512
rect 3559 11509 3571 11543
rect 3513 11503 3571 11509
rect 4154 11500 4160 11552
rect 4212 11500 4218 11552
rect 6546 11500 6552 11552
rect 6604 11540 6610 11552
rect 6733 11543 6791 11549
rect 6733 11540 6745 11543
rect 6604 11512 6745 11540
rect 6604 11500 6610 11512
rect 6733 11509 6745 11512
rect 6779 11509 6791 11543
rect 6733 11503 6791 11509
rect 8386 11500 8392 11552
rect 8444 11500 8450 11552
rect 11238 11500 11244 11552
rect 11296 11540 11302 11552
rect 11333 11543 11391 11549
rect 11333 11540 11345 11543
rect 11296 11512 11345 11540
rect 11296 11500 11302 11512
rect 11333 11509 11345 11512
rect 11379 11509 11391 11543
rect 11333 11503 11391 11509
rect 11606 11500 11612 11552
rect 11664 11500 11670 11552
rect 12406 11540 12434 11580
rect 13992 11577 14004 11611
rect 14038 11608 14050 11611
rect 14182 11608 14188 11620
rect 14038 11580 14188 11608
rect 14038 11577 14050 11580
rect 13992 11571 14050 11577
rect 14182 11568 14188 11580
rect 14240 11568 14246 11620
rect 14274 11568 14280 11620
rect 14332 11608 14338 11620
rect 14844 11608 14872 11648
rect 15657 11645 15669 11679
rect 15703 11676 15715 11679
rect 16574 11676 16580 11688
rect 15703 11648 16580 11676
rect 15703 11645 15715 11648
rect 15657 11639 15715 11645
rect 16574 11636 16580 11648
rect 16632 11676 16638 11688
rect 18156 11685 18184 11784
rect 19150 11772 19156 11784
rect 19208 11772 19214 11824
rect 19058 11704 19064 11756
rect 19116 11704 19122 11756
rect 21100 11753 21128 11852
rect 21266 11840 21272 11852
rect 21324 11840 21330 11892
rect 22830 11840 22836 11892
rect 22888 11840 22894 11892
rect 22922 11840 22928 11892
rect 22980 11880 22986 11892
rect 23109 11883 23167 11889
rect 23109 11880 23121 11883
rect 22980 11852 23121 11880
rect 22980 11840 22986 11852
rect 23109 11849 23121 11852
rect 23155 11849 23167 11883
rect 23109 11843 23167 11849
rect 23293 11883 23351 11889
rect 23293 11849 23305 11883
rect 23339 11880 23351 11883
rect 23474 11880 23480 11892
rect 23339 11852 23480 11880
rect 23339 11849 23351 11852
rect 23293 11843 23351 11849
rect 22465 11815 22523 11821
rect 22465 11781 22477 11815
rect 22511 11812 22523 11815
rect 22848 11812 22876 11840
rect 22511 11784 22876 11812
rect 22511 11781 22523 11784
rect 22465 11775 22523 11781
rect 20625 11747 20683 11753
rect 20625 11713 20637 11747
rect 20671 11744 20683 11747
rect 21085 11747 21143 11753
rect 21085 11744 21097 11747
rect 20671 11716 21097 11744
rect 20671 11713 20683 11716
rect 20625 11707 20683 11713
rect 21085 11713 21097 11716
rect 21131 11713 21143 11747
rect 21085 11707 21143 11713
rect 17497 11679 17555 11685
rect 17497 11676 17509 11679
rect 16632 11648 17509 11676
rect 16632 11636 16638 11648
rect 17497 11645 17509 11648
rect 17543 11645 17555 11679
rect 17497 11639 17555 11645
rect 18141 11679 18199 11685
rect 18141 11645 18153 11679
rect 18187 11645 18199 11679
rect 18141 11639 18199 11645
rect 18230 11636 18236 11688
rect 18288 11676 18294 11688
rect 18690 11676 18696 11688
rect 18288 11648 18696 11676
rect 18288 11636 18294 11648
rect 18690 11636 18696 11648
rect 18748 11636 18754 11688
rect 18877 11679 18935 11685
rect 18877 11645 18889 11679
rect 18923 11676 18935 11679
rect 19076 11676 19104 11704
rect 18923 11648 19104 11676
rect 18923 11645 18935 11648
rect 18877 11639 18935 11645
rect 20346 11636 20352 11688
rect 20404 11685 20410 11688
rect 20404 11639 20416 11685
rect 21352 11679 21410 11685
rect 21352 11645 21364 11679
rect 21398 11676 21410 11679
rect 22554 11676 22560 11688
rect 21398 11648 22560 11676
rect 21398 11645 21410 11648
rect 21352 11639 21410 11645
rect 20404 11636 20410 11639
rect 22554 11636 22560 11648
rect 22612 11636 22618 11688
rect 22848 11685 22876 11784
rect 22833 11679 22891 11685
rect 22833 11645 22845 11679
rect 22879 11645 22891 11679
rect 22833 11639 22891 11645
rect 22925 11679 22983 11685
rect 22925 11645 22937 11679
rect 22971 11676 22983 11679
rect 22971 11648 23060 11676
rect 22971 11645 22983 11648
rect 22925 11639 22983 11645
rect 23032 11620 23060 11648
rect 14332 11580 14872 11608
rect 14332 11568 14338 11580
rect 15010 11568 15016 11620
rect 15068 11608 15074 11620
rect 15565 11611 15623 11617
rect 15565 11608 15577 11611
rect 15068 11580 15577 11608
rect 15068 11568 15074 11580
rect 15565 11577 15577 11580
rect 15611 11577 15623 11611
rect 15565 11571 15623 11577
rect 23014 11568 23020 11620
rect 23072 11568 23078 11620
rect 23124 11608 23152 11843
rect 23474 11840 23480 11852
rect 23532 11840 23538 11892
rect 23937 11883 23995 11889
rect 23937 11849 23949 11883
rect 23983 11880 23995 11883
rect 24578 11880 24584 11892
rect 23983 11852 24584 11880
rect 23983 11849 23995 11852
rect 23937 11843 23995 11849
rect 24578 11840 24584 11852
rect 24636 11840 24642 11892
rect 24762 11840 24768 11892
rect 24820 11840 24826 11892
rect 24857 11883 24915 11889
rect 24857 11849 24869 11883
rect 24903 11880 24915 11883
rect 24946 11880 24952 11892
rect 24903 11852 24952 11880
rect 24903 11849 24915 11852
rect 24857 11843 24915 11849
rect 24946 11840 24952 11852
rect 25004 11840 25010 11892
rect 26789 11883 26847 11889
rect 26789 11849 26801 11883
rect 26835 11880 26847 11883
rect 26878 11880 26884 11892
rect 26835 11852 26884 11880
rect 26835 11849 26847 11852
rect 26789 11843 26847 11849
rect 26878 11840 26884 11852
rect 26936 11840 26942 11892
rect 23566 11772 23572 11824
rect 23624 11812 23630 11824
rect 23624 11784 23704 11812
rect 23624 11772 23630 11784
rect 23382 11744 23388 11756
rect 23216 11716 23388 11744
rect 23216 11685 23244 11716
rect 23382 11704 23388 11716
rect 23440 11744 23446 11756
rect 23676 11744 23704 11784
rect 24946 11744 24952 11756
rect 23440 11716 23612 11744
rect 23676 11716 24164 11744
rect 23440 11704 23446 11716
rect 23584 11688 23612 11716
rect 23201 11679 23259 11685
rect 23201 11645 23213 11679
rect 23247 11645 23259 11679
rect 23477 11679 23535 11685
rect 23477 11676 23489 11679
rect 23201 11639 23259 11645
rect 23308 11648 23489 11676
rect 23308 11608 23336 11648
rect 23477 11645 23489 11648
rect 23523 11645 23535 11679
rect 23477 11639 23535 11645
rect 23566 11636 23572 11688
rect 23624 11636 23630 11688
rect 24136 11685 24164 11716
rect 24320 11716 24952 11744
rect 24320 11685 24348 11716
rect 24946 11704 24952 11716
rect 25004 11704 25010 11756
rect 23845 11679 23903 11685
rect 23845 11645 23857 11679
rect 23891 11645 23903 11679
rect 24029 11679 24087 11685
rect 24029 11676 24041 11679
rect 23845 11639 23903 11645
rect 23952 11648 24041 11676
rect 23124 11580 23336 11608
rect 23382 11568 23388 11620
rect 23440 11608 23446 11620
rect 23860 11608 23888 11639
rect 23440 11580 23888 11608
rect 23440 11568 23446 11580
rect 12529 11543 12587 11549
rect 12529 11540 12541 11543
rect 12406 11512 12541 11540
rect 12529 11509 12541 11512
rect 12575 11509 12587 11543
rect 12529 11503 12587 11509
rect 12986 11500 12992 11552
rect 13044 11500 13050 11552
rect 15102 11500 15108 11552
rect 15160 11500 15166 11552
rect 16574 11500 16580 11552
rect 16632 11540 16638 11552
rect 17037 11543 17095 11549
rect 17037 11540 17049 11543
rect 16632 11512 17049 11540
rect 16632 11500 16638 11512
rect 17037 11509 17049 11512
rect 17083 11509 17095 11543
rect 17037 11503 17095 11509
rect 17402 11500 17408 11552
rect 17460 11500 17466 11552
rect 19242 11500 19248 11552
rect 19300 11500 19306 11552
rect 22649 11543 22707 11549
rect 22649 11509 22661 11543
rect 22695 11540 22707 11543
rect 23290 11540 23296 11552
rect 22695 11512 23296 11540
rect 22695 11509 22707 11512
rect 22649 11503 22707 11509
rect 23290 11500 23296 11512
rect 23348 11540 23354 11552
rect 23952 11540 23980 11648
rect 24029 11645 24041 11648
rect 24075 11645 24087 11679
rect 24029 11639 24087 11645
rect 24121 11679 24179 11685
rect 24121 11645 24133 11679
rect 24167 11645 24179 11679
rect 24121 11639 24179 11645
rect 24305 11679 24363 11685
rect 24305 11645 24317 11679
rect 24351 11645 24363 11679
rect 24305 11639 24363 11645
rect 24397 11679 24455 11685
rect 24397 11645 24409 11679
rect 24443 11645 24455 11679
rect 24397 11639 24455 11645
rect 24489 11679 24547 11685
rect 24489 11645 24501 11679
rect 24535 11645 24547 11679
rect 24489 11639 24547 11645
rect 23348 11512 23980 11540
rect 24412 11540 24440 11639
rect 24504 11608 24532 11639
rect 25130 11636 25136 11688
rect 25188 11676 25194 11688
rect 25225 11679 25283 11685
rect 25225 11676 25237 11679
rect 25188 11648 25237 11676
rect 25188 11636 25194 11648
rect 25225 11645 25237 11648
rect 25271 11645 25283 11679
rect 25225 11639 25283 11645
rect 24504 11580 24716 11608
rect 24688 11552 24716 11580
rect 25038 11568 25044 11620
rect 25096 11568 25102 11620
rect 25317 11611 25375 11617
rect 25317 11577 25329 11611
rect 25363 11577 25375 11611
rect 25317 11571 25375 11577
rect 24486 11540 24492 11552
rect 24412 11512 24492 11540
rect 23348 11500 23354 11512
rect 24486 11500 24492 11512
rect 24544 11500 24550 11552
rect 24670 11500 24676 11552
rect 24728 11500 24734 11552
rect 24762 11500 24768 11552
rect 24820 11540 24826 11552
rect 25332 11540 25360 11571
rect 24820 11512 25360 11540
rect 24820 11500 24826 11512
rect 552 11450 27576 11472
rect 552 11398 7114 11450
rect 7166 11398 7178 11450
rect 7230 11398 7242 11450
rect 7294 11398 7306 11450
rect 7358 11398 7370 11450
rect 7422 11398 13830 11450
rect 13882 11398 13894 11450
rect 13946 11398 13958 11450
rect 14010 11398 14022 11450
rect 14074 11398 14086 11450
rect 14138 11398 20546 11450
rect 20598 11398 20610 11450
rect 20662 11398 20674 11450
rect 20726 11398 20738 11450
rect 20790 11398 20802 11450
rect 20854 11398 27262 11450
rect 27314 11398 27326 11450
rect 27378 11398 27390 11450
rect 27442 11398 27454 11450
rect 27506 11398 27518 11450
rect 27570 11398 27576 11450
rect 552 11376 27576 11398
rect 1762 11296 1768 11348
rect 1820 11336 1826 11348
rect 2130 11336 2136 11348
rect 1820 11308 2136 11336
rect 1820 11296 1826 11308
rect 2130 11296 2136 11308
rect 2188 11296 2194 11348
rect 2225 11339 2283 11345
rect 2225 11305 2237 11339
rect 2271 11336 2283 11339
rect 2958 11336 2964 11348
rect 2271 11308 2964 11336
rect 2271 11305 2283 11308
rect 2225 11299 2283 11305
rect 2958 11296 2964 11308
rect 3016 11296 3022 11348
rect 4614 11296 4620 11348
rect 4672 11296 4678 11348
rect 6914 11296 6920 11348
rect 6972 11336 6978 11348
rect 7101 11339 7159 11345
rect 7101 11336 7113 11339
rect 6972 11308 7113 11336
rect 6972 11296 6978 11308
rect 7101 11305 7113 11308
rect 7147 11305 7159 11339
rect 7101 11299 7159 11305
rect 7742 11296 7748 11348
rect 7800 11296 7806 11348
rect 8386 11296 8392 11348
rect 8444 11296 8450 11348
rect 8754 11296 8760 11348
rect 8812 11296 8818 11348
rect 8846 11296 8852 11348
rect 8904 11336 8910 11348
rect 8941 11339 8999 11345
rect 8941 11336 8953 11339
rect 8904 11308 8953 11336
rect 8904 11296 8910 11308
rect 8941 11305 8953 11308
rect 8987 11305 8999 11339
rect 8941 11299 8999 11305
rect 9582 11296 9588 11348
rect 9640 11296 9646 11348
rect 9861 11339 9919 11345
rect 9861 11305 9873 11339
rect 9907 11336 9919 11339
rect 10042 11336 10048 11348
rect 9907 11308 10048 11336
rect 9907 11305 9919 11308
rect 9861 11299 9919 11305
rect 10042 11296 10048 11308
rect 10100 11296 10106 11348
rect 12986 11296 12992 11348
rect 13044 11336 13050 11348
rect 13449 11339 13507 11345
rect 13449 11336 13461 11339
rect 13044 11308 13461 11336
rect 13044 11296 13050 11308
rect 13449 11305 13461 11308
rect 13495 11305 13507 11339
rect 13449 11299 13507 11305
rect 14093 11339 14151 11345
rect 14093 11305 14105 11339
rect 14139 11336 14151 11339
rect 14182 11336 14188 11348
rect 14139 11308 14188 11336
rect 14139 11305 14151 11308
rect 14093 11299 14151 11305
rect 14182 11296 14188 11308
rect 14240 11296 14246 11348
rect 14550 11336 14556 11348
rect 14476 11308 14556 11336
rect 4341 11271 4399 11277
rect 2746 11240 4292 11268
rect 1118 11209 1124 11212
rect 1112 11163 1124 11209
rect 1118 11160 1124 11163
rect 1176 11160 1182 11212
rect 2593 11203 2651 11209
rect 2593 11169 2605 11203
rect 2639 11200 2651 11203
rect 2746 11200 2774 11240
rect 4264 11212 4292 11240
rect 4341 11237 4353 11271
rect 4387 11268 4399 11271
rect 4798 11268 4804 11280
rect 4387 11240 4804 11268
rect 4387 11237 4399 11240
rect 4341 11231 4399 11237
rect 4798 11228 4804 11240
rect 4856 11228 4862 11280
rect 5905 11271 5963 11277
rect 5905 11268 5917 11271
rect 4908 11240 5917 11268
rect 2958 11209 2964 11212
rect 2639 11172 2774 11200
rect 2639 11169 2651 11172
rect 2593 11163 2651 11169
rect 2952 11163 2964 11209
rect 2958 11160 2964 11163
rect 3016 11160 3022 11212
rect 4062 11160 4068 11212
rect 4120 11200 4126 11212
rect 4157 11203 4215 11209
rect 4157 11200 4169 11203
rect 4120 11172 4169 11200
rect 4120 11160 4126 11172
rect 4157 11169 4169 11172
rect 4203 11169 4215 11203
rect 4157 11163 4215 11169
rect 4246 11160 4252 11212
rect 4304 11160 4310 11212
rect 4908 11209 4936 11240
rect 5905 11237 5917 11240
rect 5951 11268 5963 11271
rect 7377 11271 7435 11277
rect 7377 11268 7389 11271
rect 5951 11240 7389 11268
rect 5951 11237 5963 11240
rect 5905 11231 5963 11237
rect 7377 11237 7389 11240
rect 7423 11237 7435 11271
rect 7377 11231 7435 11237
rect 7466 11228 7472 11280
rect 7524 11268 7530 11280
rect 7561 11271 7619 11277
rect 7561 11268 7573 11271
rect 7524 11240 7573 11268
rect 7524 11228 7530 11240
rect 7561 11237 7573 11240
rect 7607 11237 7619 11271
rect 7561 11231 7619 11237
rect 4893 11203 4951 11209
rect 4893 11169 4905 11203
rect 4939 11169 4951 11203
rect 4893 11163 4951 11169
rect 4982 11160 4988 11212
rect 5040 11160 5046 11212
rect 5077 11203 5135 11209
rect 5077 11169 5089 11203
rect 5123 11169 5135 11203
rect 5077 11163 5135 11169
rect 5261 11203 5319 11209
rect 5261 11169 5273 11203
rect 5307 11200 5319 11203
rect 5442 11200 5448 11212
rect 5307 11172 5448 11200
rect 5307 11169 5319 11172
rect 5261 11163 5319 11169
rect 845 11135 903 11141
rect 845 11101 857 11135
rect 891 11101 903 11135
rect 2685 11135 2743 11141
rect 2685 11132 2697 11135
rect 845 11095 903 11101
rect 2148 11104 2697 11132
rect 860 10996 888 11095
rect 2148 11008 2176 11104
rect 2685 11101 2697 11104
rect 2731 11101 2743 11135
rect 2685 11095 2743 11101
rect 4525 11135 4583 11141
rect 4525 11101 4537 11135
rect 4571 11132 4583 11135
rect 5092 11132 5120 11163
rect 5442 11160 5448 11172
rect 5500 11160 5506 11212
rect 6546 11160 6552 11212
rect 6604 11160 6610 11212
rect 6638 11160 6644 11212
rect 6696 11160 6702 11212
rect 6730 11160 6736 11212
rect 6788 11160 6794 11212
rect 6822 11160 6828 11212
rect 6880 11160 6886 11212
rect 6914 11160 6920 11212
rect 6972 11160 6978 11212
rect 8404 11209 8432 11296
rect 8772 11268 8800 11296
rect 9125 11271 9183 11277
rect 9125 11268 9137 11271
rect 8772 11240 9137 11268
rect 9125 11237 9137 11240
rect 9171 11237 9183 11271
rect 9125 11231 9183 11237
rect 8389 11203 8447 11209
rect 8389 11169 8401 11203
rect 8435 11169 8447 11203
rect 8389 11163 8447 11169
rect 8481 11203 8539 11209
rect 8481 11169 8493 11203
rect 8527 11200 8539 11203
rect 8662 11200 8668 11212
rect 8527 11172 8668 11200
rect 8527 11169 8539 11172
rect 8481 11163 8539 11169
rect 8662 11160 8668 11172
rect 8720 11160 8726 11212
rect 8938 11160 8944 11212
rect 8996 11200 9002 11212
rect 9033 11203 9091 11209
rect 9033 11200 9045 11203
rect 8996 11172 9045 11200
rect 8996 11160 9002 11172
rect 9033 11169 9045 11172
rect 9079 11169 9091 11203
rect 9033 11163 9091 11169
rect 9493 11203 9551 11209
rect 9493 11169 9505 11203
rect 9539 11169 9551 11203
rect 9493 11163 9551 11169
rect 4571 11104 5120 11132
rect 4571 11101 4583 11104
rect 4525 11095 4583 11101
rect 2409 11067 2467 11073
rect 2409 11033 2421 11067
rect 2455 11064 2467 11067
rect 2498 11064 2504 11076
rect 2455 11036 2504 11064
rect 2455 11033 2467 11036
rect 2409 11027 2467 11033
rect 2498 11024 2504 11036
rect 2556 11024 2562 11076
rect 4065 11067 4123 11073
rect 4065 11033 4077 11067
rect 4111 11064 4123 11067
rect 4154 11064 4160 11076
rect 4111 11036 4160 11064
rect 4111 11033 4123 11036
rect 4065 11027 4123 11033
rect 4154 11024 4160 11036
rect 4212 11064 4218 11076
rect 4212 11036 6132 11064
rect 4212 11024 4218 11036
rect 6104 11008 6132 11036
rect 2130 10996 2136 11008
rect 860 10968 2136 10996
rect 2130 10956 2136 10968
rect 2188 10956 2194 11008
rect 6086 10956 6092 11008
rect 6144 10956 6150 11008
rect 6564 10996 6592 11160
rect 6748 11132 6776 11160
rect 7193 11135 7251 11141
rect 7193 11132 7205 11135
rect 6748 11104 7205 11132
rect 7193 11101 7205 11104
rect 7239 11101 7251 11135
rect 7193 11095 7251 11101
rect 9508 11064 9536 11163
rect 9600 11141 9628 11296
rect 9674 11228 9680 11280
rect 9732 11268 9738 11280
rect 10229 11271 10287 11277
rect 10229 11268 10241 11271
rect 9732 11240 10241 11268
rect 9732 11228 9738 11240
rect 10229 11237 10241 11240
rect 10275 11237 10287 11271
rect 10229 11231 10287 11237
rect 11606 11228 11612 11280
rect 11664 11268 11670 11280
rect 12130 11271 12188 11277
rect 12130 11268 12142 11271
rect 11664 11240 12142 11268
rect 11664 11228 11670 11240
rect 12130 11237 12142 11240
rect 12176 11237 12188 11271
rect 14476 11268 14504 11308
rect 14550 11296 14556 11308
rect 14608 11296 14614 11348
rect 15010 11296 15016 11348
rect 15068 11296 15074 11348
rect 15102 11296 15108 11348
rect 15160 11296 15166 11348
rect 16574 11296 16580 11348
rect 16632 11296 16638 11348
rect 16669 11339 16727 11345
rect 16669 11305 16681 11339
rect 16715 11305 16727 11339
rect 16669 11299 16727 11305
rect 12130 11231 12188 11237
rect 14200 11240 14504 11268
rect 14200 11212 14228 11240
rect 9766 11160 9772 11212
rect 9824 11200 9830 11212
rect 9953 11203 10011 11209
rect 9953 11200 9965 11203
rect 9824 11172 9965 11200
rect 9824 11160 9830 11172
rect 9953 11169 9965 11172
rect 9999 11169 10011 11203
rect 9953 11163 10011 11169
rect 10042 11160 10048 11212
rect 10100 11160 10106 11212
rect 11149 11203 11207 11209
rect 11149 11169 11161 11203
rect 11195 11200 11207 11203
rect 11238 11200 11244 11212
rect 11195 11172 11244 11200
rect 11195 11169 11207 11172
rect 11149 11163 11207 11169
rect 11238 11160 11244 11172
rect 11296 11160 11302 11212
rect 11882 11160 11888 11212
rect 11940 11209 11946 11212
rect 11940 11200 11950 11209
rect 13633 11203 13691 11209
rect 13633 11200 13645 11203
rect 11940 11172 11985 11200
rect 13280 11172 13645 11200
rect 11940 11163 11950 11172
rect 11940 11160 11946 11163
rect 9585 11135 9643 11141
rect 9585 11101 9597 11135
rect 9631 11101 9643 11135
rect 9585 11095 9643 11101
rect 11333 11135 11391 11141
rect 11333 11101 11345 11135
rect 11379 11101 11391 11135
rect 11333 11095 11391 11101
rect 11054 11064 11060 11076
rect 9508 11036 11060 11064
rect 11054 11024 11060 11036
rect 11112 11064 11118 11076
rect 11348 11064 11376 11095
rect 11112 11036 11376 11064
rect 11112 11024 11118 11036
rect 6641 10999 6699 11005
rect 6641 10996 6653 10999
rect 6564 10968 6653 10996
rect 6641 10965 6653 10968
rect 6687 10965 6699 10999
rect 6641 10959 6699 10965
rect 8478 10956 8484 11008
rect 8536 10996 8542 11008
rect 8573 10999 8631 11005
rect 8573 10996 8585 10999
rect 8536 10968 8585 10996
rect 8536 10956 8542 10968
rect 8573 10965 8585 10968
rect 8619 10965 8631 10999
rect 8573 10959 8631 10965
rect 9398 10956 9404 11008
rect 9456 10996 9462 11008
rect 9766 10996 9772 11008
rect 9456 10968 9772 10996
rect 9456 10956 9462 10968
rect 9766 10956 9772 10968
rect 9824 10956 9830 11008
rect 10226 10956 10232 11008
rect 10284 10956 10290 11008
rect 12986 10956 12992 11008
rect 13044 10996 13050 11008
rect 13280 11005 13308 11172
rect 13633 11169 13645 11172
rect 13679 11169 13691 11203
rect 13633 11163 13691 11169
rect 13817 11203 13875 11209
rect 13817 11169 13829 11203
rect 13863 11169 13875 11203
rect 13817 11163 13875 11169
rect 13832 11064 13860 11163
rect 14182 11160 14188 11212
rect 14240 11160 14246 11212
rect 14274 11160 14280 11212
rect 14332 11160 14338 11212
rect 14369 11203 14427 11209
rect 14369 11169 14381 11203
rect 14415 11200 14427 11203
rect 14476 11200 14504 11240
rect 14415 11172 14504 11200
rect 14553 11203 14611 11209
rect 14415 11169 14427 11172
rect 14369 11163 14427 11169
rect 14553 11169 14565 11203
rect 14599 11200 14611 11203
rect 14829 11203 14887 11209
rect 14829 11200 14841 11203
rect 14599 11172 14841 11200
rect 14599 11169 14611 11172
rect 14553 11163 14611 11169
rect 14829 11169 14841 11172
rect 14875 11200 14887 11203
rect 15120 11200 15148 11296
rect 14875 11172 15148 11200
rect 16485 11203 16543 11209
rect 14875 11169 14887 11172
rect 14829 11163 14887 11169
rect 16485 11169 16497 11203
rect 16531 11200 16543 11203
rect 16592 11200 16620 11296
rect 16684 11268 16712 11299
rect 17402 11296 17408 11348
rect 17460 11336 17466 11348
rect 18233 11339 18291 11345
rect 18233 11336 18245 11339
rect 17460 11308 18245 11336
rect 17460 11296 17466 11308
rect 18233 11305 18245 11308
rect 18279 11305 18291 11339
rect 18233 11299 18291 11305
rect 19794 11296 19800 11348
rect 19852 11296 19858 11348
rect 22830 11296 22836 11348
rect 22888 11296 22894 11348
rect 23566 11296 23572 11348
rect 23624 11336 23630 11348
rect 25961 11339 26019 11345
rect 25961 11336 25973 11339
rect 23624 11308 25973 11336
rect 23624 11296 23630 11308
rect 25961 11305 25973 11308
rect 26007 11305 26019 11339
rect 25961 11299 26019 11305
rect 17006 11271 17064 11277
rect 17006 11268 17018 11271
rect 16684 11240 17018 11268
rect 17006 11237 17018 11240
rect 17052 11237 17064 11271
rect 17006 11231 17064 11237
rect 19242 11228 19248 11280
rect 19300 11268 19306 11280
rect 22848 11268 22876 11296
rect 19300 11240 19656 11268
rect 19300 11228 19306 11240
rect 18414 11200 18420 11212
rect 16531 11172 16620 11200
rect 18156 11172 18420 11200
rect 16531 11169 16543 11172
rect 16485 11163 16543 11169
rect 14645 11135 14703 11141
rect 14645 11101 14657 11135
rect 14691 11132 14703 11135
rect 14691 11104 14872 11132
rect 14691 11101 14703 11104
rect 14645 11095 14703 11101
rect 14844 11076 14872 11104
rect 16666 11092 16672 11144
rect 16724 11132 16730 11144
rect 16761 11135 16819 11141
rect 16761 11132 16773 11135
rect 16724 11104 16773 11132
rect 16724 11092 16730 11104
rect 16761 11101 16773 11104
rect 16807 11101 16819 11135
rect 16761 11095 16819 11101
rect 14826 11064 14832 11076
rect 13832 11036 14832 11064
rect 14826 11024 14832 11036
rect 14884 11024 14890 11076
rect 18156 11073 18184 11172
rect 18414 11160 18420 11172
rect 18472 11160 18478 11212
rect 19628 11209 19656 11240
rect 22664 11240 22876 11268
rect 22925 11271 22983 11277
rect 22664 11209 22692 11240
rect 22925 11237 22937 11271
rect 22971 11268 22983 11271
rect 23474 11268 23480 11280
rect 22971 11240 23480 11268
rect 22971 11237 22983 11240
rect 22925 11231 22983 11237
rect 23474 11228 23480 11240
rect 23532 11228 23538 11280
rect 23750 11228 23756 11280
rect 23808 11268 23814 11280
rect 23906 11271 23964 11277
rect 23906 11268 23918 11271
rect 23808 11240 23918 11268
rect 23808 11228 23814 11240
rect 23906 11237 23918 11240
rect 23952 11237 23964 11271
rect 23906 11231 23964 11237
rect 19613 11203 19671 11209
rect 19613 11169 19625 11203
rect 19659 11169 19671 11203
rect 19613 11163 19671 11169
rect 22649 11203 22707 11209
rect 22649 11169 22661 11203
rect 22695 11169 22707 11203
rect 22649 11163 22707 11169
rect 22741 11203 22799 11209
rect 22741 11169 22753 11203
rect 22787 11200 22799 11203
rect 23014 11200 23020 11212
rect 22787 11172 23020 11200
rect 22787 11169 22799 11172
rect 22741 11163 22799 11169
rect 23014 11160 23020 11172
rect 23072 11200 23078 11212
rect 23569 11203 23627 11209
rect 23072 11172 23520 11200
rect 23072 11160 23078 11172
rect 18230 11092 18236 11144
rect 18288 11132 18294 11144
rect 18601 11135 18659 11141
rect 18601 11132 18613 11135
rect 18288 11104 18613 11132
rect 18288 11092 18294 11104
rect 18601 11101 18613 11104
rect 18647 11132 18659 11135
rect 19426 11132 19432 11144
rect 18647 11104 19432 11132
rect 18647 11101 18659 11104
rect 18601 11095 18659 11101
rect 19426 11092 19432 11104
rect 19484 11092 19490 11144
rect 23492 11141 23520 11172
rect 23569 11169 23581 11203
rect 23615 11200 23627 11203
rect 25314 11200 25320 11212
rect 23615 11172 25320 11200
rect 23615 11169 23627 11172
rect 23569 11163 23627 11169
rect 25314 11160 25320 11172
rect 25372 11160 25378 11212
rect 25777 11203 25835 11209
rect 25777 11169 25789 11203
rect 25823 11200 25835 11203
rect 25869 11203 25927 11209
rect 25869 11200 25881 11203
rect 25823 11172 25881 11200
rect 25823 11169 25835 11172
rect 25777 11163 25835 11169
rect 25869 11169 25881 11172
rect 25915 11169 25927 11203
rect 25869 11163 25927 11169
rect 23477 11135 23535 11141
rect 23477 11101 23489 11135
rect 23523 11101 23535 11135
rect 23477 11095 23535 11101
rect 23658 11092 23664 11144
rect 23716 11092 23722 11144
rect 25133 11135 25191 11141
rect 25133 11101 25145 11135
rect 25179 11101 25191 11135
rect 25133 11095 25191 11101
rect 18141 11067 18199 11073
rect 18141 11033 18153 11067
rect 18187 11033 18199 11067
rect 18141 11027 18199 11033
rect 22925 11067 22983 11073
rect 22925 11033 22937 11067
rect 22971 11064 22983 11067
rect 23382 11064 23388 11076
rect 22971 11036 23388 11064
rect 22971 11033 22983 11036
rect 22925 11027 22983 11033
rect 23382 11024 23388 11036
rect 23440 11024 23446 11076
rect 25041 11067 25099 11073
rect 25041 11033 25053 11067
rect 25087 11064 25099 11067
rect 25148 11064 25176 11095
rect 25087 11036 25176 11064
rect 25087 11033 25099 11036
rect 25041 11027 25099 11033
rect 13265 10999 13323 11005
rect 13265 10996 13277 10999
rect 13044 10968 13277 10996
rect 13044 10956 13050 10968
rect 13265 10965 13277 10968
rect 13311 10965 13323 10999
rect 13265 10959 13323 10965
rect 14274 10956 14280 11008
rect 14332 10996 14338 11008
rect 14553 10999 14611 11005
rect 14553 10996 14565 10999
rect 14332 10968 14565 10996
rect 14332 10956 14338 10968
rect 14553 10965 14565 10968
rect 14599 10965 14611 10999
rect 14553 10959 14611 10965
rect 552 10906 27416 10928
rect 552 10854 3756 10906
rect 3808 10854 3820 10906
rect 3872 10854 3884 10906
rect 3936 10854 3948 10906
rect 4000 10854 4012 10906
rect 4064 10854 10472 10906
rect 10524 10854 10536 10906
rect 10588 10854 10600 10906
rect 10652 10854 10664 10906
rect 10716 10854 10728 10906
rect 10780 10854 17188 10906
rect 17240 10854 17252 10906
rect 17304 10854 17316 10906
rect 17368 10854 17380 10906
rect 17432 10854 17444 10906
rect 17496 10854 23904 10906
rect 23956 10854 23968 10906
rect 24020 10854 24032 10906
rect 24084 10854 24096 10906
rect 24148 10854 24160 10906
rect 24212 10854 27416 10906
rect 552 10832 27416 10854
rect 1118 10752 1124 10804
rect 1176 10792 1182 10804
rect 1489 10795 1547 10801
rect 1489 10792 1501 10795
rect 1176 10764 1501 10792
rect 1176 10752 1182 10764
rect 1489 10761 1501 10764
rect 1535 10761 1547 10795
rect 1489 10755 1547 10761
rect 1670 10752 1676 10804
rect 1728 10752 1734 10804
rect 4982 10752 4988 10804
rect 5040 10792 5046 10804
rect 6730 10792 6736 10804
rect 5040 10764 6736 10792
rect 5040 10752 5046 10764
rect 6730 10752 6736 10764
rect 6788 10752 6794 10804
rect 6822 10752 6828 10804
rect 6880 10792 6886 10804
rect 7929 10795 7987 10801
rect 7929 10792 7941 10795
rect 6880 10764 7941 10792
rect 6880 10752 6886 10764
rect 7929 10761 7941 10764
rect 7975 10761 7987 10795
rect 7929 10755 7987 10761
rect 9585 10795 9643 10801
rect 9585 10761 9597 10795
rect 9631 10792 9643 10795
rect 10042 10792 10048 10804
rect 9631 10764 10048 10792
rect 9631 10761 9643 10764
rect 9585 10755 9643 10761
rect 1397 10727 1455 10733
rect 1397 10693 1409 10727
rect 1443 10724 1455 10727
rect 1688 10724 1716 10752
rect 5534 10724 5540 10736
rect 1443 10696 1716 10724
rect 3252 10696 5540 10724
rect 1443 10693 1455 10696
rect 1397 10687 1455 10693
rect 1486 10616 1492 10668
rect 1544 10656 1550 10668
rect 2041 10659 2099 10665
rect 2041 10656 2053 10659
rect 1544 10628 2053 10656
rect 1544 10616 1550 10628
rect 2041 10625 2053 10628
rect 2087 10625 2099 10659
rect 2041 10619 2099 10625
rect 1026 10548 1032 10600
rect 1084 10548 1090 10600
rect 1210 10548 1216 10600
rect 1268 10548 1274 10600
rect 3053 10591 3111 10597
rect 3053 10557 3065 10591
rect 3099 10557 3111 10591
rect 3252 10588 3280 10696
rect 5534 10684 5540 10696
rect 5592 10684 5598 10736
rect 5810 10724 5816 10736
rect 5736 10696 5816 10724
rect 3326 10616 3332 10668
rect 3384 10656 3390 10668
rect 5736 10665 5764 10696
rect 5810 10684 5816 10696
rect 5868 10684 5874 10736
rect 6270 10684 6276 10736
rect 6328 10724 6334 10736
rect 6328 10696 7788 10724
rect 6328 10684 6334 10696
rect 4249 10659 4307 10665
rect 3384 10628 3648 10656
rect 3384 10616 3390 10628
rect 3620 10597 3648 10628
rect 4249 10625 4261 10659
rect 4295 10656 4307 10659
rect 4893 10659 4951 10665
rect 4893 10656 4905 10659
rect 4295 10628 4905 10656
rect 4295 10625 4307 10628
rect 4249 10619 4307 10625
rect 4893 10625 4905 10628
rect 4939 10625 4951 10659
rect 4893 10619 4951 10625
rect 5721 10659 5779 10665
rect 5721 10625 5733 10659
rect 5767 10625 5779 10659
rect 6748 10656 7052 10664
rect 5721 10619 5779 10625
rect 6380 10636 7052 10656
rect 6380 10628 6776 10636
rect 3421 10591 3479 10597
rect 3421 10588 3433 10591
rect 3252 10560 3433 10588
rect 3053 10551 3111 10557
rect 3421 10557 3433 10560
rect 3467 10557 3479 10591
rect 3421 10551 3479 10557
rect 3605 10591 3663 10597
rect 3605 10557 3617 10591
rect 3651 10557 3663 10591
rect 3605 10551 3663 10557
rect 3068 10464 3096 10551
rect 3694 10548 3700 10600
rect 3752 10548 3758 10600
rect 3789 10591 3847 10597
rect 3789 10557 3801 10591
rect 3835 10557 3847 10591
rect 3789 10551 3847 10557
rect 3510 10480 3516 10532
rect 3568 10520 3574 10532
rect 3804 10520 3832 10551
rect 4982 10548 4988 10600
rect 5040 10548 5046 10600
rect 5166 10548 5172 10600
rect 5224 10548 5230 10600
rect 5261 10591 5319 10597
rect 5261 10557 5273 10591
rect 5307 10557 5319 10591
rect 5261 10551 5319 10557
rect 5353 10591 5411 10597
rect 5353 10557 5365 10591
rect 5399 10557 5411 10591
rect 5353 10551 5411 10557
rect 3568 10492 3832 10520
rect 5000 10520 5028 10548
rect 5276 10520 5304 10551
rect 5000 10492 5304 10520
rect 5368 10520 5396 10551
rect 5534 10548 5540 10600
rect 5592 10588 5598 10600
rect 6380 10588 6408 10628
rect 5592 10560 6408 10588
rect 5592 10548 5598 10560
rect 6546 10548 6552 10600
rect 6604 10588 6610 10600
rect 6641 10591 6699 10597
rect 6641 10588 6653 10591
rect 6604 10560 6653 10588
rect 6604 10548 6610 10560
rect 6641 10557 6653 10560
rect 6687 10557 6699 10591
rect 6641 10551 6699 10557
rect 6730 10548 6736 10600
rect 6788 10548 6794 10600
rect 6822 10548 6828 10600
rect 6880 10548 6886 10600
rect 7024 10597 7052 10636
rect 7009 10591 7067 10597
rect 7009 10557 7021 10591
rect 7055 10557 7067 10591
rect 7009 10551 7067 10557
rect 7466 10548 7472 10600
rect 7524 10588 7530 10600
rect 7760 10597 7788 10696
rect 9217 10659 9275 10665
rect 9217 10656 9229 10659
rect 9140 10628 9229 10656
rect 9140 10600 9168 10628
rect 9217 10625 9229 10628
rect 9263 10625 9275 10659
rect 9217 10619 9275 10625
rect 7561 10591 7619 10597
rect 7561 10588 7573 10591
rect 7524 10560 7573 10588
rect 7524 10548 7530 10560
rect 7561 10557 7573 10560
rect 7607 10557 7619 10591
rect 7561 10551 7619 10557
rect 7745 10591 7803 10597
rect 7745 10557 7757 10591
rect 7791 10557 7803 10591
rect 7745 10551 7803 10557
rect 8202 10548 8208 10600
rect 8260 10548 8266 10600
rect 9122 10548 9128 10600
rect 9180 10548 9186 10600
rect 9398 10548 9404 10600
rect 9456 10548 9462 10600
rect 9493 10591 9551 10597
rect 9493 10557 9505 10591
rect 9539 10588 9551 10591
rect 9600 10588 9628 10755
rect 10042 10752 10048 10764
rect 10100 10752 10106 10804
rect 24946 10752 24952 10804
rect 25004 10752 25010 10804
rect 13078 10684 13084 10736
rect 13136 10724 13142 10736
rect 18138 10724 18144 10736
rect 13136 10696 18144 10724
rect 13136 10684 13142 10696
rect 18138 10684 18144 10696
rect 18196 10684 18202 10736
rect 10226 10616 10232 10668
rect 10284 10656 10290 10668
rect 10321 10659 10379 10665
rect 10321 10656 10333 10659
rect 10284 10628 10333 10656
rect 10284 10616 10290 10628
rect 10321 10625 10333 10628
rect 10367 10625 10379 10659
rect 10321 10619 10379 10625
rect 12268 10628 13032 10656
rect 9539 10560 9628 10588
rect 9539 10557 9551 10560
rect 9493 10551 9551 10557
rect 10134 10548 10140 10600
rect 10192 10588 10198 10600
rect 10870 10588 10876 10600
rect 10192 10560 10876 10588
rect 10192 10548 10198 10560
rect 10870 10548 10876 10560
rect 10928 10548 10934 10600
rect 12158 10548 12164 10600
rect 12216 10548 12222 10600
rect 12268 10597 12296 10628
rect 13004 10600 13032 10628
rect 19426 10616 19432 10668
rect 19484 10656 19490 10668
rect 19521 10659 19579 10665
rect 19521 10656 19533 10659
rect 19484 10628 19533 10656
rect 19484 10616 19490 10628
rect 19521 10625 19533 10628
rect 19567 10625 19579 10659
rect 21085 10659 21143 10665
rect 21085 10656 21097 10659
rect 19521 10619 19579 10625
rect 20732 10628 21097 10656
rect 12253 10591 12311 10597
rect 12253 10557 12265 10591
rect 12299 10557 12311 10591
rect 12253 10551 12311 10557
rect 12437 10591 12495 10597
rect 12437 10557 12449 10591
rect 12483 10557 12495 10591
rect 12437 10551 12495 10557
rect 12529 10591 12587 10597
rect 12529 10557 12541 10591
rect 12575 10557 12587 10591
rect 12529 10551 12587 10557
rect 7101 10523 7159 10529
rect 7101 10520 7113 10523
rect 5368 10492 7113 10520
rect 3568 10480 3574 10492
rect 7101 10489 7113 10492
rect 7147 10489 7159 10523
rect 7101 10483 7159 10489
rect 7285 10523 7343 10529
rect 7285 10489 7297 10523
rect 7331 10489 7343 10523
rect 7285 10483 7343 10489
rect 9217 10523 9275 10529
rect 9217 10489 9229 10523
rect 9263 10520 9275 10523
rect 9674 10520 9680 10532
rect 9263 10492 9680 10520
rect 9263 10489 9275 10492
rect 9217 10483 9275 10489
rect 2314 10412 2320 10464
rect 2372 10452 2378 10464
rect 2409 10455 2467 10461
rect 2409 10452 2421 10455
rect 2372 10424 2421 10452
rect 2372 10412 2378 10424
rect 2409 10421 2421 10424
rect 2455 10421 2467 10455
rect 2409 10415 2467 10421
rect 3050 10412 3056 10464
rect 3108 10412 3114 10464
rect 4065 10455 4123 10461
rect 4065 10421 4077 10455
rect 4111 10452 4123 10455
rect 4154 10452 4160 10464
rect 4111 10424 4160 10452
rect 4111 10421 4123 10424
rect 4065 10415 4123 10421
rect 4154 10412 4160 10424
rect 4212 10412 4218 10464
rect 4798 10412 4804 10464
rect 4856 10412 4862 10464
rect 5166 10412 5172 10464
rect 5224 10452 5230 10464
rect 6270 10452 6276 10464
rect 5224 10424 6276 10452
rect 5224 10412 5230 10424
rect 6270 10412 6276 10424
rect 6328 10412 6334 10464
rect 6362 10412 6368 10464
rect 6420 10412 6426 10464
rect 6454 10412 6460 10464
rect 6512 10452 6518 10464
rect 7300 10452 7328 10483
rect 9674 10480 9680 10492
rect 9732 10480 9738 10532
rect 6512 10424 7328 10452
rect 6512 10412 6518 10424
rect 8018 10412 8024 10464
rect 8076 10412 8082 10464
rect 10778 10412 10784 10464
rect 10836 10452 10842 10464
rect 10965 10455 11023 10461
rect 10965 10452 10977 10455
rect 10836 10424 10977 10452
rect 10836 10412 10842 10424
rect 10965 10421 10977 10424
rect 11011 10421 11023 10455
rect 10965 10415 11023 10421
rect 11974 10412 11980 10464
rect 12032 10412 12038 10464
rect 12452 10452 12480 10551
rect 12544 10520 12572 10551
rect 12986 10548 12992 10600
rect 13044 10588 13050 10600
rect 13173 10591 13231 10597
rect 13173 10588 13185 10591
rect 13044 10560 13185 10588
rect 13044 10548 13050 10560
rect 13173 10557 13185 10560
rect 13219 10557 13231 10591
rect 13173 10551 13231 10557
rect 13357 10591 13415 10597
rect 13357 10557 13369 10591
rect 13403 10588 13415 10591
rect 13630 10588 13636 10600
rect 13403 10560 13636 10588
rect 13403 10557 13415 10560
rect 13357 10551 13415 10557
rect 13630 10548 13636 10560
rect 13688 10548 13694 10600
rect 14918 10548 14924 10600
rect 14976 10548 14982 10600
rect 15381 10591 15439 10597
rect 15381 10557 15393 10591
rect 15427 10588 15439 10591
rect 15565 10591 15623 10597
rect 15427 10560 15516 10588
rect 15427 10557 15439 10560
rect 15381 10551 15439 10557
rect 13446 10520 13452 10532
rect 12544 10492 13452 10520
rect 13446 10480 13452 10492
rect 13504 10480 13510 10532
rect 15488 10464 15516 10560
rect 15565 10557 15577 10591
rect 15611 10588 15623 10591
rect 15654 10588 15660 10600
rect 15611 10560 15660 10588
rect 15611 10557 15623 10560
rect 15565 10551 15623 10557
rect 15654 10548 15660 10560
rect 15712 10548 15718 10600
rect 16022 10548 16028 10600
rect 16080 10548 16086 10600
rect 18414 10548 18420 10600
rect 18472 10588 18478 10600
rect 18693 10591 18751 10597
rect 18693 10588 18705 10591
rect 18472 10560 18705 10588
rect 18472 10548 18478 10560
rect 18693 10557 18705 10560
rect 18739 10557 18751 10591
rect 18693 10551 18751 10557
rect 18877 10591 18935 10597
rect 18877 10557 18889 10591
rect 18923 10557 18935 10591
rect 18877 10551 18935 10557
rect 18969 10591 19027 10597
rect 18969 10557 18981 10591
rect 19015 10588 19027 10591
rect 19058 10588 19064 10600
rect 19015 10560 19064 10588
rect 19015 10557 19027 10560
rect 18969 10551 19027 10557
rect 18598 10480 18604 10532
rect 18656 10520 18662 10532
rect 18892 10520 18920 10551
rect 19058 10548 19064 10560
rect 19116 10548 19122 10600
rect 19153 10591 19211 10597
rect 19153 10557 19165 10591
rect 19199 10588 19211 10591
rect 19242 10588 19248 10600
rect 19199 10560 19248 10588
rect 19199 10557 19211 10560
rect 19153 10551 19211 10557
rect 19168 10520 19196 10551
rect 19242 10548 19248 10560
rect 19300 10548 19306 10600
rect 19702 10548 19708 10600
rect 19760 10548 19766 10600
rect 20732 10597 20760 10628
rect 21085 10625 21097 10628
rect 21131 10625 21143 10659
rect 21085 10619 21143 10625
rect 21266 10616 21272 10668
rect 21324 10656 21330 10668
rect 21637 10659 21695 10665
rect 21637 10656 21649 10659
rect 21324 10628 21649 10656
rect 21324 10616 21330 10628
rect 21637 10625 21649 10628
rect 21683 10625 21695 10659
rect 21637 10619 21695 10625
rect 22278 10616 22284 10668
rect 22336 10616 22342 10668
rect 24486 10616 24492 10668
rect 24544 10656 24550 10668
rect 24544 10628 25084 10656
rect 24544 10616 24550 10628
rect 20625 10591 20683 10597
rect 20625 10557 20637 10591
rect 20671 10557 20683 10591
rect 20625 10551 20683 10557
rect 20717 10591 20775 10597
rect 20717 10557 20729 10591
rect 20763 10557 20775 10591
rect 20717 10551 20775 10557
rect 20809 10591 20867 10597
rect 20809 10557 20821 10591
rect 20855 10588 20867 10591
rect 20898 10588 20904 10600
rect 20855 10560 20904 10588
rect 20855 10557 20867 10560
rect 20809 10551 20867 10557
rect 18656 10492 19196 10520
rect 18656 10480 18662 10492
rect 20346 10480 20352 10532
rect 20404 10480 20410 10532
rect 20640 10520 20668 10551
rect 20898 10548 20904 10560
rect 20956 10548 20962 10600
rect 20993 10591 21051 10597
rect 20993 10557 21005 10591
rect 21039 10588 21051 10591
rect 21542 10588 21548 10600
rect 21039 10560 21548 10588
rect 21039 10557 21051 10560
rect 20993 10551 21051 10557
rect 21542 10548 21548 10560
rect 21600 10548 21606 10600
rect 21821 10591 21879 10597
rect 21821 10557 21833 10591
rect 21867 10588 21879 10591
rect 21910 10588 21916 10600
rect 21867 10560 21916 10588
rect 21867 10557 21879 10560
rect 21821 10551 21879 10557
rect 21910 10548 21916 10560
rect 21968 10548 21974 10600
rect 22097 10591 22155 10597
rect 22097 10557 22109 10591
rect 22143 10588 22155 10591
rect 22186 10588 22192 10600
rect 22143 10560 22192 10588
rect 22143 10557 22155 10560
rect 22097 10551 22155 10557
rect 22186 10548 22192 10560
rect 22244 10548 22250 10600
rect 24670 10548 24676 10600
rect 24728 10588 24734 10600
rect 25056 10597 25084 10628
rect 24857 10591 24915 10597
rect 24857 10588 24869 10591
rect 24728 10560 24869 10588
rect 24728 10548 24734 10560
rect 24857 10557 24869 10560
rect 24903 10557 24915 10591
rect 24857 10551 24915 10557
rect 25041 10591 25099 10597
rect 25041 10557 25053 10591
rect 25087 10557 25099 10591
rect 25041 10551 25099 10557
rect 20640 10492 21036 10520
rect 21008 10464 21036 10492
rect 12894 10452 12900 10464
rect 12452 10424 12900 10452
rect 12894 10412 12900 10424
rect 12952 10452 12958 10464
rect 13078 10452 13084 10464
rect 12952 10424 13084 10452
rect 12952 10412 12958 10424
rect 13078 10412 13084 10424
rect 13136 10412 13142 10464
rect 13262 10412 13268 10464
rect 13320 10412 13326 10464
rect 14734 10412 14740 10464
rect 14792 10412 14798 10464
rect 15194 10412 15200 10464
rect 15252 10412 15258 10464
rect 15470 10412 15476 10464
rect 15528 10412 15534 10464
rect 16209 10455 16267 10461
rect 16209 10421 16221 10455
rect 16255 10452 16267 10455
rect 16758 10452 16764 10464
rect 16255 10424 16764 10452
rect 16255 10421 16267 10424
rect 16209 10415 16267 10421
rect 16758 10412 16764 10424
rect 16816 10412 16822 10464
rect 18782 10412 18788 10464
rect 18840 10412 18846 10464
rect 18874 10412 18880 10464
rect 18932 10452 18938 10464
rect 19061 10455 19119 10461
rect 19061 10452 19073 10455
rect 18932 10424 19073 10452
rect 18932 10412 18938 10424
rect 19061 10421 19073 10424
rect 19107 10421 19119 10455
rect 19061 10415 19119 10421
rect 19886 10412 19892 10464
rect 19944 10412 19950 10464
rect 20990 10412 20996 10464
rect 21048 10412 21054 10464
rect 21082 10412 21088 10464
rect 21140 10452 21146 10464
rect 21913 10455 21971 10461
rect 21913 10452 21925 10455
rect 21140 10424 21925 10452
rect 21140 10412 21146 10424
rect 21913 10421 21925 10424
rect 21959 10421 21971 10455
rect 21913 10415 21971 10421
rect 552 10362 27576 10384
rect 552 10310 7114 10362
rect 7166 10310 7178 10362
rect 7230 10310 7242 10362
rect 7294 10310 7306 10362
rect 7358 10310 7370 10362
rect 7422 10310 13830 10362
rect 13882 10310 13894 10362
rect 13946 10310 13958 10362
rect 14010 10310 14022 10362
rect 14074 10310 14086 10362
rect 14138 10310 20546 10362
rect 20598 10310 20610 10362
rect 20662 10310 20674 10362
rect 20726 10310 20738 10362
rect 20790 10310 20802 10362
rect 20854 10310 27262 10362
rect 27314 10310 27326 10362
rect 27378 10310 27390 10362
rect 27442 10310 27454 10362
rect 27506 10310 27518 10362
rect 27570 10310 27576 10362
rect 552 10288 27576 10310
rect 1854 10208 1860 10260
rect 1912 10208 1918 10260
rect 2682 10208 2688 10260
rect 2740 10248 2746 10260
rect 3694 10248 3700 10260
rect 2740 10220 3700 10248
rect 2740 10208 2746 10220
rect 3694 10208 3700 10220
rect 3752 10208 3758 10260
rect 4890 10208 4896 10260
rect 4948 10208 4954 10260
rect 6273 10251 6331 10257
rect 6273 10217 6285 10251
rect 6319 10248 6331 10251
rect 6638 10248 6644 10260
rect 6319 10220 6644 10248
rect 6319 10217 6331 10220
rect 6273 10211 6331 10217
rect 6638 10208 6644 10220
rect 6696 10208 6702 10260
rect 7558 10208 7564 10260
rect 7616 10208 7622 10260
rect 8018 10208 8024 10260
rect 8076 10208 8082 10260
rect 8938 10208 8944 10260
rect 8996 10208 9002 10260
rect 9401 10251 9459 10257
rect 9401 10217 9413 10251
rect 9447 10248 9459 10251
rect 10134 10248 10140 10260
rect 9447 10220 10140 10248
rect 9447 10217 9459 10220
rect 9401 10211 9459 10217
rect 10134 10208 10140 10220
rect 10192 10208 10198 10260
rect 10778 10208 10784 10260
rect 10836 10208 10842 10260
rect 13446 10208 13452 10260
rect 13504 10208 13510 10260
rect 13817 10251 13875 10257
rect 13817 10217 13829 10251
rect 13863 10248 13875 10251
rect 14550 10248 14556 10260
rect 13863 10220 14556 10248
rect 13863 10217 13875 10220
rect 13817 10211 13875 10217
rect 14550 10208 14556 10220
rect 14608 10208 14614 10260
rect 15930 10208 15936 10260
rect 15988 10208 15994 10260
rect 16022 10208 16028 10260
rect 16080 10248 16086 10260
rect 16117 10251 16175 10257
rect 16117 10248 16129 10251
rect 16080 10220 16129 10248
rect 16080 10208 16086 10220
rect 16117 10217 16129 10220
rect 16163 10217 16175 10251
rect 17865 10251 17923 10257
rect 17865 10248 17877 10251
rect 16117 10211 16175 10217
rect 16408 10220 17877 10248
rect 3142 10180 3148 10192
rect 1412 10152 3148 10180
rect 1412 10121 1440 10152
rect 3142 10140 3148 10152
rect 3200 10140 3206 10192
rect 3602 10140 3608 10192
rect 3660 10140 3666 10192
rect 5810 10140 5816 10192
rect 5868 10140 5874 10192
rect 7576 10180 7604 10208
rect 7208 10152 7604 10180
rect 1213 10115 1271 10121
rect 1213 10081 1225 10115
rect 1259 10081 1271 10115
rect 1213 10075 1271 10081
rect 1397 10115 1455 10121
rect 1397 10081 1409 10115
rect 1443 10081 1455 10115
rect 1397 10075 1455 10081
rect 1489 10115 1547 10121
rect 1489 10081 1501 10115
rect 1535 10081 1547 10115
rect 1489 10075 1547 10081
rect 1581 10115 1639 10121
rect 1581 10081 1593 10115
rect 1627 10112 1639 10115
rect 1854 10112 1860 10124
rect 1627 10084 1860 10112
rect 1627 10081 1639 10084
rect 1581 10075 1639 10081
rect 1228 9908 1256 10075
rect 1302 10004 1308 10056
rect 1360 10044 1366 10056
rect 1504 10044 1532 10075
rect 1854 10072 1860 10084
rect 1912 10072 1918 10124
rect 2406 10121 2412 10124
rect 2400 10075 2412 10121
rect 2406 10072 2412 10075
rect 2464 10072 2470 10124
rect 6086 10072 6092 10124
rect 6144 10072 6150 10124
rect 6454 10072 6460 10124
rect 6512 10072 6518 10124
rect 6914 10072 6920 10124
rect 6972 10112 6978 10124
rect 7208 10121 7236 10152
rect 7009 10115 7067 10121
rect 7009 10112 7021 10115
rect 6972 10084 7021 10112
rect 6972 10072 6978 10084
rect 7009 10081 7021 10084
rect 7055 10081 7067 10115
rect 7009 10075 7067 10081
rect 7193 10115 7251 10121
rect 7193 10081 7205 10115
rect 7239 10081 7251 10115
rect 7193 10075 7251 10081
rect 7460 10115 7518 10121
rect 7460 10081 7472 10115
rect 7506 10112 7518 10115
rect 8036 10112 8064 10208
rect 8956 10180 8984 10208
rect 9125 10183 9183 10189
rect 9125 10180 9137 10183
rect 8956 10152 9137 10180
rect 9125 10149 9137 10152
rect 9171 10149 9183 10183
rect 9125 10143 9183 10149
rect 10536 10183 10594 10189
rect 10536 10149 10548 10183
rect 10582 10180 10594 10183
rect 10796 10180 10824 10208
rect 10582 10152 10824 10180
rect 10582 10149 10594 10152
rect 10536 10143 10594 10149
rect 10870 10140 10876 10192
rect 10928 10180 10934 10192
rect 14734 10189 14740 10192
rect 14717 10183 14740 10189
rect 10928 10152 11284 10180
rect 10928 10140 10934 10152
rect 7506 10084 8064 10112
rect 8941 10115 8999 10121
rect 7506 10081 7518 10084
rect 7460 10075 7518 10081
rect 8941 10081 8953 10115
rect 8987 10112 8999 10115
rect 9490 10112 9496 10124
rect 8987 10084 9496 10112
rect 8987 10081 8999 10084
rect 8941 10075 8999 10081
rect 1360 10016 1532 10044
rect 1360 10004 1366 10016
rect 2130 10004 2136 10056
rect 2188 10004 2194 10056
rect 5994 10004 6000 10056
rect 6052 10044 6058 10056
rect 6472 10044 6500 10072
rect 6052 10016 6500 10044
rect 6052 10004 6058 10016
rect 8573 9979 8631 9985
rect 8573 9945 8585 9979
rect 8619 9976 8631 9979
rect 8956 9976 8984 10075
rect 9490 10072 9496 10084
rect 9548 10072 9554 10124
rect 10781 10115 10839 10121
rect 10781 10081 10793 10115
rect 10827 10112 10839 10115
rect 10962 10112 10968 10124
rect 10827 10084 10968 10112
rect 10827 10081 10839 10084
rect 10781 10075 10839 10081
rect 10962 10072 10968 10084
rect 11020 10072 11026 10124
rect 11054 10072 11060 10124
rect 11112 10072 11118 10124
rect 11256 10121 11284 10152
rect 13004 10152 13584 10180
rect 13004 10124 13032 10152
rect 11241 10115 11299 10121
rect 11241 10081 11253 10115
rect 11287 10081 11299 10115
rect 11241 10075 11299 10081
rect 12069 10115 12127 10121
rect 12069 10081 12081 10115
rect 12115 10112 12127 10115
rect 12897 10115 12955 10121
rect 12897 10112 12909 10115
rect 12115 10084 12909 10112
rect 12115 10081 12127 10084
rect 12069 10075 12127 10081
rect 12897 10081 12909 10084
rect 12943 10081 12955 10115
rect 12897 10075 12955 10081
rect 12912 10044 12940 10075
rect 12986 10072 12992 10124
rect 13044 10072 13050 10124
rect 13078 10072 13084 10124
rect 13136 10112 13142 10124
rect 13173 10115 13231 10121
rect 13173 10112 13185 10115
rect 13136 10084 13185 10112
rect 13136 10072 13142 10084
rect 13173 10081 13185 10084
rect 13219 10081 13231 10115
rect 13173 10075 13231 10081
rect 13262 10072 13268 10124
rect 13320 10072 13326 10124
rect 13354 10072 13360 10124
rect 13412 10072 13418 10124
rect 13556 10121 13584 10152
rect 14016 10152 14504 10180
rect 14016 10121 14044 10152
rect 13541 10115 13599 10121
rect 13541 10081 13553 10115
rect 13587 10081 13599 10115
rect 13541 10075 13599 10081
rect 14001 10115 14059 10121
rect 14001 10081 14013 10115
rect 14047 10081 14059 10115
rect 14001 10075 14059 10081
rect 14093 10115 14151 10121
rect 14093 10081 14105 10115
rect 14139 10112 14151 10115
rect 14182 10112 14188 10124
rect 14139 10084 14188 10112
rect 14139 10081 14151 10084
rect 14093 10075 14151 10081
rect 14016 10044 14044 10075
rect 14182 10072 14188 10084
rect 14240 10072 14246 10124
rect 14274 10072 14280 10124
rect 14332 10072 14338 10124
rect 14369 10115 14427 10121
rect 14369 10081 14381 10115
rect 14415 10081 14427 10115
rect 14476 10112 14504 10152
rect 14717 10149 14729 10183
rect 14717 10143 14740 10149
rect 14734 10140 14740 10143
rect 14792 10140 14798 10192
rect 15948 10180 15976 10208
rect 16408 10180 16436 10220
rect 17865 10217 17877 10220
rect 17911 10217 17923 10251
rect 17865 10211 17923 10217
rect 18782 10208 18788 10260
rect 18840 10208 18846 10260
rect 19337 10251 19395 10257
rect 19337 10217 19349 10251
rect 19383 10217 19395 10251
rect 19337 10211 19395 10217
rect 19705 10251 19763 10257
rect 19705 10217 19717 10251
rect 19751 10248 19763 10251
rect 19886 10248 19892 10260
rect 19751 10220 19892 10248
rect 19751 10217 19763 10220
rect 19705 10211 19763 10217
rect 15948 10152 16436 10180
rect 16485 10183 16543 10189
rect 16485 10149 16497 10183
rect 16531 10180 16543 10183
rect 16574 10180 16580 10192
rect 16531 10152 16580 10180
rect 16531 10149 16543 10152
rect 16485 10143 16543 10149
rect 16574 10140 16580 10152
rect 16632 10140 16638 10192
rect 18800 10180 18828 10208
rect 16868 10152 18552 10180
rect 18800 10152 18920 10180
rect 16868 10112 16896 10152
rect 14476 10084 16896 10112
rect 14369 10075 14427 10081
rect 12912 10016 14044 10044
rect 8619 9948 8984 9976
rect 8619 9945 8631 9948
rect 8573 9939 8631 9945
rect 2038 9908 2044 9920
rect 1228 9880 2044 9908
rect 2038 9868 2044 9880
rect 2096 9908 2102 9920
rect 2498 9908 2504 9920
rect 2096 9880 2504 9908
rect 2096 9868 2102 9880
rect 2498 9868 2504 9880
rect 2556 9868 2562 9920
rect 3050 9868 3056 9920
rect 3108 9908 3114 9920
rect 3513 9911 3571 9917
rect 3513 9908 3525 9911
rect 3108 9880 3525 9908
rect 3108 9868 3114 9880
rect 3513 9877 3525 9880
rect 3559 9908 3571 9911
rect 5813 9911 5871 9917
rect 5813 9908 5825 9911
rect 3559 9880 5825 9908
rect 3559 9877 3571 9880
rect 3513 9871 3571 9877
rect 5813 9877 5825 9880
rect 5859 9877 5871 9911
rect 5813 9871 5871 9877
rect 6454 9868 6460 9920
rect 6512 9868 6518 9920
rect 8662 9868 8668 9920
rect 8720 9908 8726 9920
rect 8757 9911 8815 9917
rect 8757 9908 8769 9911
rect 8720 9880 8769 9908
rect 8720 9868 8726 9880
rect 8757 9877 8769 9880
rect 8803 9877 8815 9911
rect 8757 9871 8815 9877
rect 12713 9911 12771 9917
rect 12713 9877 12725 9911
rect 12759 9908 12771 9911
rect 13078 9908 13084 9920
rect 12759 9880 13084 9908
rect 12759 9877 12771 9880
rect 12713 9871 12771 9877
rect 13078 9868 13084 9880
rect 13136 9868 13142 9920
rect 14384 9908 14412 10075
rect 17770 10072 17776 10124
rect 17828 10072 17834 10124
rect 18524 10121 18552 10152
rect 18509 10115 18567 10121
rect 18509 10081 18521 10115
rect 18555 10081 18567 10115
rect 18509 10075 18567 10081
rect 18598 10072 18604 10124
rect 18656 10072 18662 10124
rect 18892 10121 18920 10152
rect 18785 10115 18843 10121
rect 18785 10112 18797 10115
rect 18708 10084 18797 10112
rect 18708 10056 18736 10084
rect 18785 10081 18797 10084
rect 18831 10081 18843 10115
rect 18785 10075 18843 10081
rect 18877 10115 18935 10121
rect 18877 10081 18889 10115
rect 18923 10081 18935 10115
rect 18877 10075 18935 10081
rect 19245 10115 19303 10121
rect 19245 10081 19257 10115
rect 19291 10112 19303 10115
rect 19352 10112 19380 10211
rect 19886 10208 19892 10220
rect 19944 10208 19950 10260
rect 21266 10208 21272 10260
rect 21324 10208 21330 10260
rect 21174 10180 21180 10192
rect 19291 10084 19380 10112
rect 20640 10152 21180 10180
rect 19291 10081 19303 10084
rect 19245 10075 19303 10081
rect 14458 10004 14464 10056
rect 14516 10004 14522 10056
rect 15562 10004 15568 10056
rect 15620 10004 15626 10056
rect 15746 10004 15752 10056
rect 15804 10004 15810 10056
rect 15930 10004 15936 10056
rect 15988 10044 15994 10056
rect 16577 10047 16635 10053
rect 16577 10044 16589 10047
rect 15988 10016 16589 10044
rect 15988 10004 15994 10016
rect 16577 10013 16589 10016
rect 16623 10013 16635 10047
rect 16577 10007 16635 10013
rect 16669 10047 16727 10053
rect 16669 10013 16681 10047
rect 16715 10013 16727 10047
rect 16669 10007 16727 10013
rect 17957 10047 18015 10053
rect 17957 10013 17969 10047
rect 18003 10013 18015 10047
rect 17957 10007 18015 10013
rect 15580 9976 15608 10004
rect 15396 9948 15608 9976
rect 15764 9976 15792 10004
rect 16684 9976 16712 10007
rect 15764 9948 16712 9976
rect 14458 9908 14464 9920
rect 14384 9880 14464 9908
rect 14458 9868 14464 9880
rect 14516 9908 14522 9920
rect 15396 9908 15424 9948
rect 17678 9936 17684 9988
rect 17736 9976 17742 9988
rect 17972 9976 18000 10007
rect 18690 10004 18696 10056
rect 18748 10044 18754 10056
rect 19150 10044 19156 10056
rect 18748 10016 19156 10044
rect 18748 10004 18754 10016
rect 19150 10004 19156 10016
rect 19208 10004 19214 10056
rect 19334 10004 19340 10056
rect 19392 10044 19398 10056
rect 19797 10047 19855 10053
rect 19797 10044 19809 10047
rect 19392 10016 19809 10044
rect 19392 10004 19398 10016
rect 19797 10013 19809 10016
rect 19843 10013 19855 10047
rect 19797 10007 19855 10013
rect 19978 10004 19984 10056
rect 20036 10004 20042 10056
rect 17736 9948 18000 9976
rect 18325 9979 18383 9985
rect 17736 9936 17742 9948
rect 18325 9945 18337 9979
rect 18371 9976 18383 9979
rect 20640 9976 20668 10152
rect 21174 10140 21180 10152
rect 21232 10140 21238 10192
rect 20717 10115 20775 10121
rect 20717 10081 20729 10115
rect 20763 10081 20775 10115
rect 21284 10112 21312 10208
rect 20717 10075 20775 10081
rect 20824 10084 21312 10112
rect 18371 9948 20668 9976
rect 20732 9976 20760 10075
rect 20824 10053 20852 10084
rect 22094 10072 22100 10124
rect 22152 10112 22158 10124
rect 22382 10115 22440 10121
rect 22382 10112 22394 10115
rect 22152 10084 22394 10112
rect 22152 10072 22158 10084
rect 22382 10081 22394 10084
rect 22428 10081 22440 10115
rect 22382 10075 22440 10081
rect 22649 10115 22707 10121
rect 22649 10081 22661 10115
rect 22695 10112 22707 10115
rect 23658 10112 23664 10124
rect 22695 10084 23664 10112
rect 22695 10081 22707 10084
rect 22649 10075 22707 10081
rect 23658 10072 23664 10084
rect 23716 10072 23722 10124
rect 24670 10072 24676 10124
rect 24728 10072 24734 10124
rect 20809 10047 20867 10053
rect 20809 10013 20821 10047
rect 20855 10013 20867 10047
rect 20809 10007 20867 10013
rect 21082 10004 21088 10056
rect 21140 10004 21146 10056
rect 20732 9948 21036 9976
rect 18371 9945 18383 9948
rect 18325 9939 18383 9945
rect 21008 9920 21036 9948
rect 14516 9880 15424 9908
rect 14516 9868 14522 9880
rect 15470 9868 15476 9920
rect 15528 9908 15534 9920
rect 15841 9911 15899 9917
rect 15841 9908 15853 9911
rect 15528 9880 15853 9908
rect 15528 9868 15534 9880
rect 15841 9877 15853 9880
rect 15887 9877 15899 9911
rect 15841 9871 15899 9877
rect 17405 9911 17463 9917
rect 17405 9877 17417 9911
rect 17451 9908 17463 9911
rect 17586 9908 17592 9920
rect 17451 9880 17592 9908
rect 17451 9877 17463 9880
rect 17405 9871 17463 9877
rect 17586 9868 17592 9880
rect 17644 9868 17650 9920
rect 19058 9868 19064 9920
rect 19116 9868 19122 9920
rect 20990 9868 20996 9920
rect 21048 9868 21054 9920
rect 24854 9868 24860 9920
rect 24912 9868 24918 9920
rect 552 9818 27416 9840
rect 552 9766 3756 9818
rect 3808 9766 3820 9818
rect 3872 9766 3884 9818
rect 3936 9766 3948 9818
rect 4000 9766 4012 9818
rect 4064 9766 10472 9818
rect 10524 9766 10536 9818
rect 10588 9766 10600 9818
rect 10652 9766 10664 9818
rect 10716 9766 10728 9818
rect 10780 9766 17188 9818
rect 17240 9766 17252 9818
rect 17304 9766 17316 9818
rect 17368 9766 17380 9818
rect 17432 9766 17444 9818
rect 17496 9766 23904 9818
rect 23956 9766 23968 9818
rect 24020 9766 24032 9818
rect 24084 9766 24096 9818
rect 24148 9766 24160 9818
rect 24212 9766 27416 9818
rect 552 9744 27416 9766
rect 2222 9664 2228 9716
rect 2280 9704 2286 9716
rect 2682 9704 2688 9716
rect 2280 9676 2688 9704
rect 2280 9664 2286 9676
rect 2682 9664 2688 9676
rect 2740 9664 2746 9716
rect 3510 9664 3516 9716
rect 3568 9704 3574 9716
rect 3789 9707 3847 9713
rect 3789 9704 3801 9707
rect 3568 9676 3801 9704
rect 3568 9664 3574 9676
rect 3789 9673 3801 9676
rect 3835 9673 3847 9707
rect 4890 9704 4896 9716
rect 3789 9667 3847 9673
rect 4540 9676 4896 9704
rect 2958 9596 2964 9648
rect 3016 9636 3022 9648
rect 3053 9639 3111 9645
rect 3053 9636 3065 9639
rect 3016 9608 3065 9636
rect 3016 9596 3022 9608
rect 3053 9605 3065 9608
rect 3099 9605 3111 9639
rect 3053 9599 3111 9605
rect 3697 9639 3755 9645
rect 3697 9605 3709 9639
rect 3743 9636 3755 9639
rect 4338 9636 4344 9648
rect 3743 9608 4344 9636
rect 3743 9605 3755 9608
rect 3697 9599 3755 9605
rect 4338 9596 4344 9608
rect 4396 9596 4402 9648
rect 4540 9577 4568 9676
rect 4890 9664 4896 9676
rect 4948 9704 4954 9716
rect 4948 9676 5488 9704
rect 4948 9664 4954 9676
rect 5460 9636 5488 9676
rect 5810 9664 5816 9716
rect 5868 9704 5874 9716
rect 5905 9707 5963 9713
rect 5905 9704 5917 9707
rect 5868 9676 5917 9704
rect 5868 9664 5874 9676
rect 5905 9673 5917 9676
rect 5951 9673 5963 9707
rect 5905 9667 5963 9673
rect 6914 9664 6920 9716
rect 6972 9704 6978 9716
rect 7377 9707 7435 9713
rect 7377 9704 7389 9707
rect 6972 9676 7389 9704
rect 6972 9664 6978 9676
rect 7377 9673 7389 9676
rect 7423 9673 7435 9707
rect 7377 9667 7435 9673
rect 7466 9664 7472 9716
rect 7524 9704 7530 9716
rect 8021 9707 8079 9713
rect 8021 9704 8033 9707
rect 7524 9676 8033 9704
rect 7524 9664 7530 9676
rect 8021 9673 8033 9676
rect 8067 9673 8079 9707
rect 8021 9667 8079 9673
rect 8202 9664 8208 9716
rect 8260 9664 8266 9716
rect 10137 9707 10195 9713
rect 10137 9673 10149 9707
rect 10183 9704 10195 9707
rect 10962 9704 10968 9716
rect 10183 9676 10968 9704
rect 10183 9673 10195 9676
rect 10137 9667 10195 9673
rect 5460 9608 6040 9636
rect 6012 9577 6040 9608
rect 8864 9608 9168 9636
rect 8864 9580 8892 9608
rect 4525 9571 4583 9577
rect 4525 9568 4537 9571
rect 3896 9540 4537 9568
rect 3896 9512 3924 9540
rect 4525 9537 4537 9540
rect 4571 9537 4583 9571
rect 4525 9531 4583 9537
rect 5997 9571 6055 9577
rect 5997 9537 6009 9571
rect 6043 9537 6055 9571
rect 5997 9531 6055 9537
rect 8846 9528 8852 9580
rect 8904 9528 8910 9580
rect 9030 9528 9036 9580
rect 9088 9528 9094 9580
rect 9140 9568 9168 9608
rect 9306 9596 9312 9648
rect 9364 9596 9370 9648
rect 10152 9636 10180 9667
rect 10962 9664 10968 9676
rect 11020 9664 11026 9716
rect 11054 9664 11060 9716
rect 11112 9664 11118 9716
rect 14918 9664 14924 9716
rect 14976 9664 14982 9716
rect 16316 9676 17264 9704
rect 9692 9608 10180 9636
rect 9692 9568 9720 9608
rect 9140 9540 9720 9568
rect 2130 9460 2136 9512
rect 2188 9500 2194 9512
rect 2225 9503 2283 9509
rect 2225 9500 2237 9503
rect 2188 9472 2237 9500
rect 2188 9460 2194 9472
rect 2225 9469 2237 9472
rect 2271 9469 2283 9503
rect 2225 9463 2283 9469
rect 2409 9503 2467 9509
rect 2409 9469 2421 9503
rect 2455 9500 2467 9503
rect 2498 9500 2504 9512
rect 2455 9472 2504 9500
rect 2455 9469 2467 9472
rect 2409 9463 2467 9469
rect 1946 9392 1952 9444
rect 2004 9441 2010 9444
rect 2004 9395 2016 9441
rect 2240 9432 2268 9463
rect 2498 9460 2504 9472
rect 2556 9460 2562 9512
rect 2590 9460 2596 9512
rect 2648 9460 2654 9512
rect 2682 9460 2688 9512
rect 2740 9460 2746 9512
rect 2777 9503 2835 9509
rect 2777 9469 2789 9503
rect 2823 9500 2835 9503
rect 3234 9500 3240 9512
rect 2823 9472 3240 9500
rect 2823 9469 2835 9472
rect 2777 9463 2835 9469
rect 3234 9460 3240 9472
rect 3292 9460 3298 9512
rect 3329 9503 3387 9509
rect 3329 9469 3341 9503
rect 3375 9500 3387 9503
rect 3418 9500 3424 9512
rect 3375 9472 3424 9500
rect 3375 9469 3387 9472
rect 3329 9463 3387 9469
rect 3418 9460 3424 9472
rect 3476 9460 3482 9512
rect 3878 9460 3884 9512
rect 3936 9460 3942 9512
rect 4798 9509 4804 9512
rect 4433 9503 4491 9509
rect 4433 9469 4445 9503
rect 4479 9469 4491 9503
rect 4792 9500 4804 9509
rect 4759 9472 4804 9500
rect 4433 9463 4491 9469
rect 4792 9463 4804 9472
rect 3513 9435 3571 9441
rect 2240 9404 3004 9432
rect 2004 9392 2010 9395
rect 2976 9376 3004 9404
rect 3513 9401 3525 9435
rect 3559 9401 3571 9435
rect 4448 9432 4476 9463
rect 4798 9460 4804 9463
rect 4856 9460 4862 9512
rect 7653 9503 7711 9509
rect 7653 9469 7665 9503
rect 7699 9500 7711 9503
rect 7926 9500 7932 9512
rect 7699 9472 7932 9500
rect 7699 9469 7711 9472
rect 7653 9463 7711 9469
rect 7926 9460 7932 9472
rect 7984 9460 7990 9512
rect 8757 9503 8815 9509
rect 8757 9469 8769 9503
rect 8803 9469 8815 9503
rect 8757 9463 8815 9469
rect 8941 9503 8999 9509
rect 8941 9469 8953 9503
rect 8987 9500 8999 9503
rect 9490 9500 9496 9512
rect 8987 9472 9496 9500
rect 8987 9469 8999 9472
rect 8941 9463 8999 9469
rect 5994 9432 6000 9444
rect 4448 9404 6000 9432
rect 3513 9395 3571 9401
rect 842 9324 848 9376
rect 900 9324 906 9376
rect 2314 9324 2320 9376
rect 2372 9364 2378 9376
rect 2498 9364 2504 9376
rect 2372 9336 2504 9364
rect 2372 9324 2378 9336
rect 2498 9324 2504 9336
rect 2556 9324 2562 9376
rect 2958 9324 2964 9376
rect 3016 9324 3022 9376
rect 3528 9364 3556 9395
rect 5994 9392 6000 9404
rect 6052 9392 6058 9444
rect 6264 9435 6322 9441
rect 6264 9401 6276 9435
rect 6310 9432 6322 9435
rect 6362 9432 6368 9444
rect 6310 9404 6368 9432
rect 6310 9401 6322 9404
rect 6264 9395 6322 9401
rect 6362 9392 6368 9404
rect 6420 9392 6426 9444
rect 8021 9435 8079 9441
rect 8021 9401 8033 9435
rect 8067 9432 8079 9435
rect 8662 9432 8668 9444
rect 8067 9404 8668 9432
rect 8067 9401 8079 9404
rect 8021 9395 8079 9401
rect 8662 9392 8668 9404
rect 8720 9392 8726 9444
rect 8772 9432 8800 9463
rect 9490 9460 9496 9472
rect 9548 9460 9554 9512
rect 9585 9503 9643 9509
rect 9585 9469 9597 9503
rect 9631 9500 9643 9503
rect 9692 9500 9720 9540
rect 9861 9571 9919 9577
rect 9861 9537 9873 9571
rect 9907 9568 9919 9571
rect 10134 9568 10140 9580
rect 9907 9540 10140 9568
rect 9907 9537 9919 9540
rect 9861 9531 9919 9537
rect 10134 9528 10140 9540
rect 10192 9528 10198 9580
rect 11072 9568 11100 9664
rect 12802 9596 12808 9648
rect 12860 9636 12866 9648
rect 13173 9639 13231 9645
rect 13173 9636 13185 9639
rect 12860 9608 13185 9636
rect 12860 9596 12866 9608
rect 13173 9605 13185 9608
rect 13219 9605 13231 9639
rect 16316 9636 16344 9676
rect 13173 9599 13231 9605
rect 15396 9608 16344 9636
rect 17236 9636 17264 9676
rect 17770 9664 17776 9716
rect 17828 9704 17834 9716
rect 17865 9707 17923 9713
rect 17865 9704 17877 9707
rect 17828 9676 17877 9704
rect 17828 9664 17834 9676
rect 17865 9673 17877 9676
rect 17911 9673 17923 9707
rect 19334 9704 19340 9716
rect 17865 9667 17923 9673
rect 18984 9676 19340 9704
rect 17678 9636 17684 9648
rect 17236 9608 17684 9636
rect 11149 9571 11207 9577
rect 11149 9568 11161 9571
rect 11072 9540 11161 9568
rect 11149 9537 11161 9540
rect 11195 9537 11207 9571
rect 11149 9531 11207 9537
rect 11885 9571 11943 9577
rect 11885 9537 11897 9571
rect 11931 9568 11943 9571
rect 12158 9568 12164 9580
rect 11931 9540 12164 9568
rect 11931 9537 11943 9540
rect 11885 9531 11943 9537
rect 12158 9528 12164 9540
rect 12216 9568 12222 9580
rect 15396 9577 15424 9608
rect 17678 9596 17684 9608
rect 17736 9636 17742 9648
rect 18984 9636 19012 9676
rect 19334 9664 19340 9676
rect 19392 9664 19398 9716
rect 19702 9664 19708 9716
rect 19760 9704 19766 9716
rect 20254 9704 20260 9716
rect 19760 9676 20260 9704
rect 19760 9664 19766 9676
rect 20254 9664 20260 9676
rect 20312 9704 20318 9716
rect 20349 9707 20407 9713
rect 20349 9704 20361 9707
rect 20312 9676 20361 9704
rect 20312 9664 20318 9676
rect 20349 9673 20361 9676
rect 20395 9673 20407 9707
rect 20349 9667 20407 9673
rect 20898 9664 20904 9716
rect 20956 9664 20962 9716
rect 21082 9664 21088 9716
rect 21140 9664 21146 9716
rect 17736 9608 19012 9636
rect 20625 9639 20683 9645
rect 17736 9596 17742 9608
rect 20625 9605 20637 9639
rect 20671 9636 20683 9639
rect 20916 9636 20944 9664
rect 20671 9608 20944 9636
rect 20671 9605 20683 9608
rect 20625 9599 20683 9605
rect 15381 9571 15439 9577
rect 12216 9540 14136 9568
rect 12216 9528 12222 9540
rect 9631 9472 9720 9500
rect 11057 9503 11115 9509
rect 9631 9469 9643 9472
rect 9585 9463 9643 9469
rect 11057 9469 11069 9503
rect 11103 9469 11115 9503
rect 11057 9463 11115 9469
rect 9677 9435 9735 9441
rect 9677 9432 9689 9435
rect 8772 9404 9689 9432
rect 9677 9401 9689 9404
rect 9723 9432 9735 9435
rect 10318 9432 10324 9444
rect 9723 9404 10324 9432
rect 9723 9401 9735 9404
rect 9677 9395 9735 9401
rect 10318 9392 10324 9404
rect 10376 9432 10382 9444
rect 11072 9432 11100 9463
rect 12342 9460 12348 9512
rect 12400 9500 12406 9512
rect 12437 9503 12495 9509
rect 12437 9500 12449 9503
rect 12400 9472 12449 9500
rect 12400 9460 12406 9472
rect 12437 9469 12449 9472
rect 12483 9469 12495 9503
rect 12437 9463 12495 9469
rect 10376 9404 11100 9432
rect 12452 9432 12480 9463
rect 12618 9460 12624 9512
rect 12676 9460 12682 9512
rect 13170 9460 13176 9512
rect 13228 9460 13234 9512
rect 14108 9509 14136 9540
rect 15381 9537 15393 9571
rect 15427 9537 15439 9571
rect 15381 9531 15439 9537
rect 15565 9571 15623 9577
rect 15565 9537 15577 9571
rect 15611 9568 15623 9571
rect 15746 9568 15752 9580
rect 15611 9540 15752 9568
rect 15611 9537 15623 9540
rect 15565 9531 15623 9537
rect 15746 9528 15752 9540
rect 15804 9528 15810 9580
rect 18969 9571 19027 9577
rect 18969 9568 18981 9571
rect 17236 9540 18981 9568
rect 13357 9503 13415 9509
rect 13357 9469 13369 9503
rect 13403 9469 13415 9503
rect 13357 9463 13415 9469
rect 14093 9503 14151 9509
rect 14093 9469 14105 9503
rect 14139 9469 14151 9503
rect 14093 9463 14151 9469
rect 12986 9432 12992 9444
rect 12452 9404 12992 9432
rect 10376 9392 10382 9404
rect 12986 9392 12992 9404
rect 13044 9432 13050 9444
rect 13372 9432 13400 9463
rect 13044 9404 13400 9432
rect 14108 9432 14136 9463
rect 14182 9460 14188 9512
rect 14240 9460 14246 9512
rect 14366 9460 14372 9512
rect 14424 9460 14430 9512
rect 14458 9460 14464 9512
rect 14516 9460 14522 9512
rect 15194 9460 15200 9512
rect 15252 9500 15258 9512
rect 15289 9503 15347 9509
rect 15289 9500 15301 9503
rect 15252 9472 15301 9500
rect 15252 9460 15258 9472
rect 15289 9469 15301 9472
rect 15335 9469 15347 9503
rect 15289 9463 15347 9469
rect 16666 9460 16672 9512
rect 16724 9500 16730 9512
rect 17126 9500 17132 9512
rect 16724 9472 17132 9500
rect 16724 9460 16730 9472
rect 17126 9460 17132 9472
rect 17184 9500 17190 9512
rect 17236 9509 17264 9540
rect 18969 9537 18981 9540
rect 19015 9537 19027 9571
rect 21100 9568 21128 9664
rect 21729 9639 21787 9645
rect 21729 9605 21741 9639
rect 21775 9636 21787 9639
rect 22094 9636 22100 9648
rect 21775 9608 22100 9636
rect 21775 9605 21787 9608
rect 21729 9599 21787 9605
rect 22094 9596 22100 9608
rect 22152 9596 22158 9648
rect 23474 9636 23480 9648
rect 22848 9608 23480 9636
rect 22848 9577 22876 9608
rect 23474 9596 23480 9608
rect 23532 9636 23538 9648
rect 24581 9639 24639 9645
rect 24581 9636 24593 9639
rect 23532 9608 24593 9636
rect 23532 9596 23538 9608
rect 24581 9605 24593 9608
rect 24627 9605 24639 9639
rect 24581 9599 24639 9605
rect 21269 9571 21327 9577
rect 21269 9568 21281 9571
rect 21100 9540 21281 9568
rect 18969 9531 19027 9537
rect 21269 9537 21281 9540
rect 21315 9537 21327 9571
rect 21269 9531 21327 9537
rect 22833 9571 22891 9577
rect 22833 9537 22845 9571
rect 22879 9537 22891 9571
rect 22833 9531 22891 9537
rect 24121 9571 24179 9577
rect 24121 9537 24133 9571
rect 24167 9568 24179 9571
rect 24302 9568 24308 9580
rect 24167 9540 24308 9568
rect 24167 9537 24179 9540
rect 24121 9531 24179 9537
rect 24302 9528 24308 9540
rect 24360 9528 24366 9580
rect 25958 9528 25964 9580
rect 26016 9528 26022 9580
rect 17221 9503 17279 9509
rect 17221 9500 17233 9503
rect 17184 9472 17233 9500
rect 17184 9460 17190 9472
rect 17221 9469 17233 9472
rect 17267 9469 17279 9503
rect 17221 9463 17279 9469
rect 17586 9460 17592 9512
rect 17644 9460 17650 9512
rect 18046 9460 18052 9512
rect 18104 9460 18110 9512
rect 18138 9460 18144 9512
rect 18196 9460 18202 9512
rect 19058 9460 19064 9512
rect 19116 9500 19122 9512
rect 19225 9503 19283 9509
rect 19225 9500 19237 9503
rect 19116 9472 19237 9500
rect 19116 9460 19122 9472
rect 19225 9469 19237 9472
rect 19271 9469 19283 9503
rect 19225 9463 19283 9469
rect 20809 9503 20867 9509
rect 20809 9469 20821 9503
rect 20855 9469 20867 9503
rect 20809 9463 20867 9469
rect 21085 9503 21143 9509
rect 21085 9469 21097 9503
rect 21131 9500 21143 9503
rect 21361 9503 21419 9509
rect 21131 9472 21312 9500
rect 21131 9469 21143 9472
rect 21085 9463 21143 9469
rect 14108 9404 15976 9432
rect 13044 9392 13050 9404
rect 6454 9364 6460 9376
rect 3528 9336 6460 9364
rect 6454 9324 6460 9336
rect 6512 9324 6518 9376
rect 9214 9324 9220 9376
rect 9272 9324 9278 9376
rect 9490 9324 9496 9376
rect 9548 9324 9554 9376
rect 9950 9324 9956 9376
rect 10008 9324 10014 9376
rect 10134 9373 10140 9376
rect 10121 9367 10140 9373
rect 10121 9333 10133 9367
rect 10121 9327 10140 9333
rect 10134 9324 10140 9327
rect 10192 9324 10198 9376
rect 12526 9324 12532 9376
rect 12584 9324 12590 9376
rect 13909 9367 13967 9373
rect 13909 9333 13921 9367
rect 13955 9364 13967 9367
rect 14642 9364 14648 9376
rect 13955 9336 14648 9364
rect 13955 9333 13967 9336
rect 13909 9327 13967 9333
rect 14642 9324 14648 9336
rect 14700 9324 14706 9376
rect 15378 9324 15384 9376
rect 15436 9364 15442 9376
rect 15838 9364 15844 9376
rect 15436 9336 15844 9364
rect 15436 9324 15442 9336
rect 15838 9324 15844 9336
rect 15896 9324 15902 9376
rect 15948 9364 15976 9404
rect 16758 9392 16764 9444
rect 16816 9432 16822 9444
rect 16954 9435 17012 9441
rect 16954 9432 16966 9435
rect 16816 9404 16966 9432
rect 16816 9392 16822 9404
rect 16954 9401 16966 9404
rect 17000 9401 17012 9435
rect 20824 9432 20852 9463
rect 21284 9444 21312 9472
rect 21361 9469 21373 9503
rect 21407 9469 21419 9503
rect 21361 9463 21419 9469
rect 21545 9503 21603 9509
rect 21545 9469 21557 9503
rect 21591 9500 21603 9503
rect 22186 9500 22192 9512
rect 21591 9472 22192 9500
rect 21591 9469 21603 9472
rect 21545 9463 21603 9469
rect 16954 9395 17012 9401
rect 17052 9404 19012 9432
rect 20824 9404 21128 9432
rect 17052 9364 17080 9404
rect 18984 9376 19012 9404
rect 15948 9336 17080 9364
rect 17402 9324 17408 9376
rect 17460 9324 17466 9376
rect 18966 9324 18972 9376
rect 19024 9324 19030 9376
rect 20990 9324 20996 9376
rect 21048 9324 21054 9376
rect 21100 9364 21128 9404
rect 21266 9392 21272 9444
rect 21324 9392 21330 9444
rect 21376 9432 21404 9463
rect 22186 9460 22192 9472
rect 22244 9460 22250 9512
rect 22741 9503 22799 9509
rect 22741 9469 22753 9503
rect 22787 9500 22799 9503
rect 23014 9500 23020 9512
rect 22787 9472 23020 9500
rect 22787 9469 22799 9472
rect 22741 9463 22799 9469
rect 23014 9460 23020 9472
rect 23072 9460 23078 9512
rect 24029 9503 24087 9509
rect 24029 9469 24041 9503
rect 24075 9469 24087 9503
rect 24029 9463 24087 9469
rect 21910 9432 21916 9444
rect 21376 9404 21916 9432
rect 21376 9364 21404 9404
rect 21910 9392 21916 9404
rect 21968 9392 21974 9444
rect 21100 9336 21404 9364
rect 23106 9324 23112 9376
rect 23164 9364 23170 9376
rect 24044 9364 24072 9463
rect 24854 9460 24860 9512
rect 24912 9500 24918 9512
rect 25694 9503 25752 9509
rect 25694 9500 25706 9503
rect 24912 9472 25706 9500
rect 24912 9460 24918 9472
rect 25694 9469 25706 9472
rect 25740 9469 25752 9503
rect 25694 9463 25752 9469
rect 23164 9336 24072 9364
rect 23164 9324 23170 9336
rect 24394 9324 24400 9376
rect 24452 9324 24458 9376
rect 552 9274 27576 9296
rect 552 9222 7114 9274
rect 7166 9222 7178 9274
rect 7230 9222 7242 9274
rect 7294 9222 7306 9274
rect 7358 9222 7370 9274
rect 7422 9222 13830 9274
rect 13882 9222 13894 9274
rect 13946 9222 13958 9274
rect 14010 9222 14022 9274
rect 14074 9222 14086 9274
rect 14138 9222 20546 9274
rect 20598 9222 20610 9274
rect 20662 9222 20674 9274
rect 20726 9222 20738 9274
rect 20790 9222 20802 9274
rect 20854 9222 27262 9274
rect 27314 9222 27326 9274
rect 27378 9222 27390 9274
rect 27442 9222 27454 9274
rect 27506 9222 27518 9274
rect 27570 9222 27576 9274
rect 552 9200 27576 9222
rect 1213 9163 1271 9169
rect 1213 9129 1225 9163
rect 1259 9160 1271 9163
rect 1302 9160 1308 9172
rect 1259 9132 1308 9160
rect 1259 9129 1271 9132
rect 1213 9123 1271 9129
rect 1302 9120 1308 9132
rect 1360 9120 1366 9172
rect 2777 9163 2835 9169
rect 2777 9160 2789 9163
rect 1872 9132 2789 9160
rect 1872 9036 1900 9132
rect 2777 9129 2789 9132
rect 2823 9129 2835 9163
rect 2777 9123 2835 9129
rect 3142 9120 3148 9172
rect 3200 9120 3206 9172
rect 3326 9120 3332 9172
rect 3384 9160 3390 9172
rect 3421 9163 3479 9169
rect 3421 9160 3433 9163
rect 3384 9132 3433 9160
rect 3384 9120 3390 9132
rect 3421 9129 3433 9132
rect 3467 9129 3479 9163
rect 3421 9123 3479 9129
rect 5261 9163 5319 9169
rect 5261 9129 5273 9163
rect 5307 9160 5319 9163
rect 5994 9160 6000 9172
rect 5307 9132 6000 9160
rect 5307 9129 5319 9132
rect 5261 9123 5319 9129
rect 5994 9120 6000 9132
rect 6052 9120 6058 9172
rect 7837 9163 7895 9169
rect 7837 9129 7849 9163
rect 7883 9160 7895 9163
rect 7883 9132 8524 9160
rect 7883 9129 7895 9132
rect 7837 9123 7895 9129
rect 2498 9092 2504 9104
rect 2332 9064 2504 9092
rect 842 8984 848 9036
rect 900 9024 906 9036
rect 1670 9024 1676 9036
rect 900 8996 1676 9024
rect 900 8984 906 8996
rect 1670 8984 1676 8996
rect 1728 9024 1734 9036
rect 1765 9027 1823 9033
rect 1765 9024 1777 9027
rect 1728 8996 1777 9024
rect 1728 8984 1734 8996
rect 1765 8993 1777 8996
rect 1811 8993 1823 9027
rect 1765 8987 1823 8993
rect 1780 8820 1808 8987
rect 1854 8984 1860 9036
rect 1912 8984 1918 9036
rect 1949 9027 2007 9033
rect 1949 8993 1961 9027
rect 1995 9024 2007 9027
rect 2038 9024 2044 9036
rect 1995 8996 2044 9024
rect 1995 8993 2007 8996
rect 1949 8987 2007 8993
rect 2038 8984 2044 8996
rect 2096 8984 2102 9036
rect 2130 8984 2136 9036
rect 2188 8984 2194 9036
rect 2222 8984 2228 9036
rect 2280 8984 2286 9036
rect 2332 9033 2360 9064
rect 2498 9052 2504 9064
rect 2556 9092 2562 9104
rect 3605 9095 3663 9101
rect 3605 9092 3617 9095
rect 2556 9064 3617 9092
rect 2556 9052 2562 9064
rect 3605 9061 3617 9064
rect 3651 9061 3663 9095
rect 8496 9092 8524 9132
rect 8846 9120 8852 9172
rect 8904 9120 8910 9172
rect 9030 9120 9036 9172
rect 9088 9120 9094 9172
rect 9214 9120 9220 9172
rect 9272 9160 9278 9172
rect 9401 9163 9459 9169
rect 9401 9160 9413 9163
rect 9272 9132 9413 9160
rect 9272 9120 9278 9132
rect 9401 9129 9413 9132
rect 9447 9129 9459 9163
rect 9401 9123 9459 9129
rect 12802 9120 12808 9172
rect 12860 9120 12866 9172
rect 12894 9120 12900 9172
rect 12952 9120 12958 9172
rect 14090 9160 14096 9172
rect 13372 9132 14096 9160
rect 8864 9092 8892 9120
rect 9048 9092 9076 9120
rect 3605 9055 3663 9061
rect 8128 9064 8432 9092
rect 2317 9027 2375 9033
rect 2317 8993 2329 9027
rect 2363 8993 2375 9027
rect 2317 8987 2375 8993
rect 2685 9027 2743 9033
rect 2685 8993 2697 9027
rect 2731 8993 2743 9027
rect 2685 8987 2743 8993
rect 2961 9027 3019 9033
rect 2961 8993 2973 9027
rect 3007 8993 3019 9027
rect 2961 8987 3019 8993
rect 2406 8916 2412 8968
rect 2464 8956 2470 8968
rect 2593 8959 2651 8965
rect 2593 8956 2605 8959
rect 2464 8928 2605 8956
rect 2464 8916 2470 8928
rect 2593 8925 2605 8928
rect 2639 8925 2651 8959
rect 2700 8956 2728 8987
rect 2700 8928 2774 8956
rect 2593 8919 2651 8925
rect 2746 8820 2774 8928
rect 2866 8916 2872 8968
rect 2924 8956 2930 8968
rect 2976 8956 3004 8987
rect 3050 8984 3056 9036
rect 3108 9024 3114 9036
rect 3418 9024 3424 9036
rect 3108 8996 3424 9024
rect 3108 8984 3114 8996
rect 3418 8984 3424 8996
rect 3476 9024 3482 9036
rect 4154 9033 4160 9036
rect 3789 9027 3847 9033
rect 3789 9024 3801 9027
rect 3476 8996 3801 9024
rect 3476 8984 3482 8996
rect 3789 8993 3801 8996
rect 3835 8993 3847 9027
rect 4148 9024 4160 9033
rect 4115 8996 4160 9024
rect 3789 8987 3847 8993
rect 4148 8987 4160 8996
rect 4154 8984 4160 8987
rect 4212 8984 4218 9036
rect 7466 8984 7472 9036
rect 7524 8984 7530 9036
rect 7926 8984 7932 9036
rect 7984 9033 7990 9036
rect 7984 9024 7992 9033
rect 8128 9024 8156 9064
rect 7984 8996 8156 9024
rect 8205 9027 8263 9033
rect 7984 8987 7992 8996
rect 8205 8993 8217 9027
rect 8251 8993 8263 9027
rect 8205 8987 8263 8993
rect 7984 8984 7990 8987
rect 2924 8928 3004 8956
rect 2924 8916 2930 8928
rect 3878 8916 3884 8968
rect 3936 8916 3942 8968
rect 2958 8848 2964 8900
rect 3016 8888 3022 8900
rect 3896 8888 3924 8916
rect 3016 8860 3924 8888
rect 7484 8888 7512 8984
rect 7653 8959 7711 8965
rect 7653 8925 7665 8959
rect 7699 8956 7711 8959
rect 8220 8956 8248 8987
rect 7699 8928 8248 8956
rect 7699 8925 7711 8928
rect 7653 8919 7711 8925
rect 8404 8897 8432 9064
rect 8496 9064 8892 9092
rect 8956 9064 9076 9092
rect 8496 9033 8524 9064
rect 8481 9027 8539 9033
rect 8481 8993 8493 9027
rect 8527 8993 8539 9027
rect 8481 8987 8539 8993
rect 8757 9027 8815 9033
rect 8757 8993 8769 9027
rect 8803 9024 8815 9027
rect 8956 9024 8984 9064
rect 9490 9052 9496 9104
rect 9548 9092 9554 9104
rect 9548 9064 11468 9092
rect 9548 9052 9554 9064
rect 8803 8996 8984 9024
rect 9033 9027 9091 9033
rect 8803 8993 8815 8996
rect 8757 8987 8815 8993
rect 9033 8993 9045 9027
rect 9079 9024 9091 9027
rect 9398 9024 9404 9036
rect 9079 8996 9404 9024
rect 9079 8993 9091 8996
rect 9033 8987 9091 8993
rect 9398 8984 9404 8996
rect 9456 9024 9462 9036
rect 9950 9024 9956 9036
rect 9456 8996 9956 9024
rect 9456 8984 9462 8996
rect 9950 8984 9956 8996
rect 10008 8984 10014 9036
rect 10134 8984 10140 9036
rect 10192 8984 10198 9036
rect 11054 8984 11060 9036
rect 11112 8984 11118 9036
rect 11440 9033 11468 9064
rect 11425 9027 11483 9033
rect 11425 8993 11437 9027
rect 11471 8993 11483 9027
rect 12820 9024 12848 9120
rect 12912 9092 12940 9120
rect 12912 9064 13124 9092
rect 13096 9033 13124 9064
rect 13372 9036 13400 9132
rect 14090 9120 14096 9132
rect 14148 9160 14154 9172
rect 14148 9132 15608 9160
rect 14148 9120 14154 9132
rect 14200 9064 14964 9092
rect 14200 9036 14228 9064
rect 12989 9027 13047 9033
rect 12989 9024 13001 9027
rect 12820 8996 13001 9024
rect 11425 8987 11483 8993
rect 12989 8993 13001 8996
rect 13035 8993 13047 9027
rect 12989 8987 13047 8993
rect 13081 9027 13139 9033
rect 13081 8993 13093 9027
rect 13127 8993 13139 9027
rect 13081 8987 13139 8993
rect 13170 8984 13176 9036
rect 13228 9024 13234 9036
rect 13265 9027 13323 9033
rect 13265 9024 13277 9027
rect 13228 8996 13277 9024
rect 13228 8984 13234 8996
rect 13265 8993 13277 8996
rect 13311 8993 13323 9027
rect 13265 8987 13323 8993
rect 13354 8984 13360 9036
rect 13412 8984 13418 9036
rect 13722 8984 13728 9036
rect 13780 9024 13786 9036
rect 14001 9027 14059 9033
rect 14001 9024 14013 9027
rect 13780 8996 14013 9024
rect 13780 8984 13786 8996
rect 14001 8993 14013 8996
rect 14047 8993 14059 9027
rect 14001 8987 14059 8993
rect 14093 9027 14151 9033
rect 14093 8993 14105 9027
rect 14139 9024 14151 9027
rect 14182 9024 14188 9036
rect 14139 8996 14188 9024
rect 14139 8993 14151 8996
rect 14093 8987 14151 8993
rect 14182 8984 14188 8996
rect 14240 8984 14246 9036
rect 14277 9027 14335 9033
rect 14277 8993 14289 9027
rect 14323 8993 14335 9027
rect 14277 8987 14335 8993
rect 14369 9027 14427 9033
rect 14369 8993 14381 9027
rect 14415 9024 14427 9027
rect 14458 9024 14464 9036
rect 14415 8996 14464 9024
rect 14415 8993 14427 8996
rect 14369 8987 14427 8993
rect 8941 8959 8999 8965
rect 8941 8925 8953 8959
rect 8987 8956 8999 8959
rect 9490 8956 9496 8968
rect 8987 8928 9496 8956
rect 8987 8925 8999 8928
rect 8941 8919 8999 8925
rect 9490 8916 9496 8928
rect 9548 8916 9554 8968
rect 8389 8891 8447 8897
rect 7484 8860 8340 8888
rect 3016 8848 3022 8860
rect 1780 8792 2774 8820
rect 8018 8780 8024 8832
rect 8076 8780 8082 8832
rect 8312 8820 8340 8860
rect 8389 8857 8401 8891
rect 8435 8888 8447 8891
rect 8573 8891 8631 8897
rect 8573 8888 8585 8891
rect 8435 8860 8585 8888
rect 8435 8857 8447 8860
rect 8389 8851 8447 8857
rect 8573 8857 8585 8860
rect 8619 8888 8631 8891
rect 10152 8888 10180 8984
rect 12434 8916 12440 8968
rect 12492 8956 12498 8968
rect 12897 8959 12955 8965
rect 12897 8956 12909 8959
rect 12492 8928 12909 8956
rect 12492 8916 12498 8928
rect 12897 8925 12909 8928
rect 12943 8956 12955 8959
rect 13740 8956 13768 8984
rect 12943 8928 13768 8956
rect 14292 8956 14320 8987
rect 14458 8984 14464 8996
rect 14516 8984 14522 9036
rect 14660 9033 14688 9064
rect 14936 9036 14964 9064
rect 14645 9027 14703 9033
rect 14645 8993 14657 9027
rect 14691 8993 14703 9027
rect 14645 8987 14703 8993
rect 14829 9027 14887 9033
rect 14829 8993 14841 9027
rect 14875 8993 14887 9027
rect 14829 8987 14887 8993
rect 14844 8956 14872 8987
rect 14918 8984 14924 9036
rect 14976 8984 14982 9036
rect 15105 9027 15163 9033
rect 15105 8993 15117 9027
rect 15151 9024 15163 9027
rect 15470 9024 15476 9036
rect 15151 8996 15476 9024
rect 15151 8993 15163 8996
rect 15105 8987 15163 8993
rect 15470 8984 15476 8996
rect 15528 8984 15534 9036
rect 15378 8956 15384 8968
rect 14292 8928 14780 8956
rect 14844 8928 15384 8956
rect 12943 8925 12955 8928
rect 12897 8919 12955 8925
rect 8619 8860 10180 8888
rect 8619 8857 8631 8860
rect 8573 8851 8631 8857
rect 14752 8832 14780 8928
rect 15378 8916 15384 8928
rect 15436 8916 15442 8968
rect 9122 8820 9128 8832
rect 8312 8792 9128 8820
rect 9122 8780 9128 8792
rect 9180 8820 9186 8832
rect 9401 8823 9459 8829
rect 9401 8820 9413 8823
rect 9180 8792 9413 8820
rect 9180 8780 9186 8792
rect 9401 8789 9413 8792
rect 9447 8789 9459 8823
rect 9401 8783 9459 8789
rect 9585 8823 9643 8829
rect 9585 8789 9597 8823
rect 9631 8820 9643 8823
rect 9674 8820 9680 8832
rect 9631 8792 9680 8820
rect 9631 8789 9643 8792
rect 9585 8783 9643 8789
rect 9674 8780 9680 8792
rect 9732 8780 9738 8832
rect 13538 8780 13544 8832
rect 13596 8780 13602 8832
rect 13817 8823 13875 8829
rect 13817 8789 13829 8823
rect 13863 8820 13875 8823
rect 14274 8820 14280 8832
rect 13863 8792 14280 8820
rect 13863 8789 13875 8792
rect 13817 8783 13875 8789
rect 14274 8780 14280 8792
rect 14332 8780 14338 8832
rect 14734 8780 14740 8832
rect 14792 8820 14798 8832
rect 14829 8823 14887 8829
rect 14829 8820 14841 8823
rect 14792 8792 14841 8820
rect 14792 8780 14798 8792
rect 14829 8789 14841 8792
rect 14875 8789 14887 8823
rect 14829 8783 14887 8789
rect 15102 8780 15108 8832
rect 15160 8780 15166 8832
rect 15580 8820 15608 9132
rect 15838 9120 15844 9172
rect 15896 9120 15902 9172
rect 16574 9120 16580 9172
rect 16632 9120 16638 9172
rect 18046 9120 18052 9172
rect 18104 9160 18110 9172
rect 18509 9163 18567 9169
rect 18509 9160 18521 9163
rect 18104 9132 18521 9160
rect 18104 9120 18110 9132
rect 18509 9129 18521 9132
rect 18555 9129 18567 9163
rect 18509 9123 18567 9129
rect 18874 9120 18880 9172
rect 18932 9120 18938 9172
rect 19334 9160 19340 9172
rect 19076 9132 19340 9160
rect 15856 9092 15884 9120
rect 17402 9101 17408 9104
rect 17385 9095 17408 9101
rect 15856 9064 16436 9092
rect 15654 8984 15660 9036
rect 15712 9024 15718 9036
rect 16408 9033 16436 9064
rect 17385 9061 17397 9095
rect 17385 9055 17408 9061
rect 17402 9052 17408 9055
rect 17460 9052 17466 9104
rect 18892 9092 18920 9120
rect 18616 9064 18920 9092
rect 16209 9027 16267 9033
rect 16209 9024 16221 9027
rect 15712 8996 16221 9024
rect 15712 8984 15718 8996
rect 16209 8993 16221 8996
rect 16255 8993 16267 9027
rect 16209 8987 16267 8993
rect 16393 9027 16451 9033
rect 16393 8993 16405 9027
rect 16439 8993 16451 9027
rect 18138 9024 18144 9036
rect 16393 8987 16451 8993
rect 16960 8996 18144 9024
rect 16224 8956 16252 8987
rect 16960 8956 16988 8996
rect 18138 8984 18144 8996
rect 18196 8984 18202 9036
rect 18616 9033 18644 9064
rect 18601 9027 18659 9033
rect 18601 8993 18613 9027
rect 18647 8993 18659 9027
rect 18601 8987 18659 8993
rect 18693 9027 18751 9033
rect 18693 8993 18705 9027
rect 18739 9024 18751 9027
rect 18782 9024 18788 9036
rect 18739 8996 18788 9024
rect 18739 8993 18751 8996
rect 18693 8987 18751 8993
rect 18782 8984 18788 8996
rect 18840 8984 18846 9036
rect 18877 9027 18935 9033
rect 18877 8993 18889 9027
rect 18923 8993 18935 9027
rect 18877 8987 18935 8993
rect 16224 8928 16988 8956
rect 17034 8916 17040 8968
rect 17092 8956 17098 8968
rect 17129 8959 17187 8965
rect 17129 8956 17141 8959
rect 17092 8928 17141 8956
rect 17092 8916 17098 8928
rect 17129 8925 17141 8928
rect 17175 8925 17187 8959
rect 18892 8956 18920 8987
rect 18966 8984 18972 9036
rect 19024 8984 19030 9036
rect 19076 8956 19104 9132
rect 19334 9120 19340 9132
rect 19392 9160 19398 9172
rect 19392 9132 19748 9160
rect 19392 9120 19398 9132
rect 19153 9095 19211 9101
rect 19153 9061 19165 9095
rect 19199 9092 19211 9095
rect 19518 9092 19524 9104
rect 19199 9064 19524 9092
rect 19199 9061 19211 9064
rect 19153 9055 19211 9061
rect 19518 9052 19524 9064
rect 19576 9052 19582 9104
rect 19720 9092 19748 9132
rect 23106 9120 23112 9172
rect 23164 9120 23170 9172
rect 23474 9120 23480 9172
rect 23532 9120 23538 9172
rect 24394 9120 24400 9172
rect 24452 9120 24458 9172
rect 24670 9120 24676 9172
rect 24728 9160 24734 9172
rect 24765 9163 24823 9169
rect 24765 9160 24777 9163
rect 24728 9132 24777 9160
rect 24728 9120 24734 9132
rect 24765 9129 24777 9132
rect 24811 9129 24823 9163
rect 24765 9123 24823 9129
rect 23124 9092 23152 9120
rect 19720 9064 20116 9092
rect 19720 9033 19748 9064
rect 20088 9033 20116 9064
rect 22848 9064 23152 9092
rect 19613 9027 19671 9033
rect 17129 8919 17187 8925
rect 18616 8928 19104 8956
rect 19168 8996 19334 9024
rect 18616 8900 18644 8928
rect 18598 8848 18604 8900
rect 18656 8848 18662 8900
rect 19168 8820 19196 8996
rect 19306 8956 19334 8996
rect 19613 8993 19625 9027
rect 19659 8993 19671 9027
rect 19613 8987 19671 8993
rect 19705 9027 19763 9033
rect 19705 8993 19717 9027
rect 19751 8993 19763 9027
rect 19705 8987 19763 8993
rect 19889 9027 19947 9033
rect 19889 8993 19901 9027
rect 19935 8993 19947 9027
rect 19889 8987 19947 8993
rect 19981 9027 20039 9033
rect 19981 8993 19993 9027
rect 20027 8993 20039 9027
rect 19981 8987 20039 8993
rect 20073 9027 20131 9033
rect 20073 8993 20085 9027
rect 20119 8993 20131 9027
rect 20073 8987 20131 8993
rect 19628 8956 19656 8987
rect 19306 8928 19656 8956
rect 19242 8848 19248 8900
rect 19300 8888 19306 8900
rect 19904 8888 19932 8987
rect 19996 8956 20024 8987
rect 20254 8984 20260 9036
rect 20312 8984 20318 9036
rect 22646 8984 22652 9036
rect 22704 8984 22710 9036
rect 22848 9033 22876 9064
rect 22833 9027 22891 9033
rect 22833 8993 22845 9027
rect 22879 8993 22891 9027
rect 22833 8987 22891 8993
rect 22925 9027 22983 9033
rect 22925 8993 22937 9027
rect 22971 8993 22983 9027
rect 22925 8987 22983 8993
rect 20165 8959 20223 8965
rect 20165 8956 20177 8959
rect 19996 8928 20177 8956
rect 20165 8925 20177 8928
rect 20211 8925 20223 8959
rect 20165 8919 20223 8925
rect 20622 8916 20628 8968
rect 20680 8956 20686 8968
rect 22278 8956 22284 8968
rect 20680 8928 22284 8956
rect 20680 8916 20686 8928
rect 22278 8916 22284 8928
rect 22336 8916 22342 8968
rect 19300 8860 19932 8888
rect 22741 8891 22799 8897
rect 19300 8848 19306 8860
rect 22741 8857 22753 8891
rect 22787 8888 22799 8891
rect 22830 8888 22836 8900
rect 22787 8860 22836 8888
rect 22787 8857 22799 8860
rect 22741 8851 22799 8857
rect 22830 8848 22836 8860
rect 22888 8848 22894 8900
rect 22940 8832 22968 8987
rect 23106 8984 23112 9036
rect 23164 9024 23170 9036
rect 23492 9033 23520 9120
rect 23385 9027 23443 9033
rect 23385 9024 23397 9027
rect 23164 8996 23397 9024
rect 23164 8984 23170 8996
rect 23385 8993 23397 8996
rect 23431 8993 23443 9027
rect 23385 8987 23443 8993
rect 23477 9027 23535 9033
rect 23477 8993 23489 9027
rect 23523 8993 23535 9027
rect 23477 8987 23535 8993
rect 23566 8984 23572 9036
rect 23624 8984 23630 9036
rect 23753 9027 23811 9033
rect 23753 8993 23765 9027
rect 23799 8993 23811 9027
rect 24412 9024 24440 9120
rect 24581 9027 24639 9033
rect 24581 9024 24593 9027
rect 24412 8996 24593 9024
rect 23753 8987 23811 8993
rect 24581 8993 24593 8996
rect 24627 8993 24639 9027
rect 24581 8987 24639 8993
rect 23474 8848 23480 8900
rect 23532 8888 23538 8900
rect 23768 8888 23796 8987
rect 24394 8916 24400 8968
rect 24452 8916 24458 8968
rect 23532 8860 23796 8888
rect 23532 8848 23538 8860
rect 15580 8792 19196 8820
rect 19429 8823 19487 8829
rect 19429 8789 19441 8823
rect 19475 8820 19487 8823
rect 21082 8820 21088 8832
rect 19475 8792 21088 8820
rect 19475 8789 19487 8792
rect 19429 8783 19487 8789
rect 21082 8780 21088 8792
rect 21140 8780 21146 8832
rect 22002 8780 22008 8832
rect 22060 8820 22066 8832
rect 22465 8823 22523 8829
rect 22465 8820 22477 8823
rect 22060 8792 22477 8820
rect 22060 8780 22066 8792
rect 22465 8789 22477 8792
rect 22511 8789 22523 8823
rect 22465 8783 22523 8789
rect 22922 8780 22928 8832
rect 22980 8780 22986 8832
rect 23014 8780 23020 8832
rect 23072 8820 23078 8832
rect 23109 8823 23167 8829
rect 23109 8820 23121 8823
rect 23072 8792 23121 8820
rect 23072 8780 23078 8792
rect 23109 8789 23121 8792
rect 23155 8789 23167 8823
rect 23109 8783 23167 8789
rect 552 8730 27416 8752
rect 552 8678 3756 8730
rect 3808 8678 3820 8730
rect 3872 8678 3884 8730
rect 3936 8678 3948 8730
rect 4000 8678 4012 8730
rect 4064 8678 10472 8730
rect 10524 8678 10536 8730
rect 10588 8678 10600 8730
rect 10652 8678 10664 8730
rect 10716 8678 10728 8730
rect 10780 8678 17188 8730
rect 17240 8678 17252 8730
rect 17304 8678 17316 8730
rect 17368 8678 17380 8730
rect 17432 8678 17444 8730
rect 17496 8678 23904 8730
rect 23956 8678 23968 8730
rect 24020 8678 24032 8730
rect 24084 8678 24096 8730
rect 24148 8678 24160 8730
rect 24212 8678 27416 8730
rect 552 8656 27416 8678
rect 1397 8619 1455 8625
rect 1397 8616 1409 8619
rect 768 8588 1409 8616
rect 768 8412 796 8588
rect 1397 8585 1409 8588
rect 1443 8616 1455 8619
rect 1443 8588 2360 8616
rect 1443 8585 1455 8588
rect 1397 8579 1455 8585
rect 1029 8551 1087 8557
rect 1029 8517 1041 8551
rect 1075 8548 1087 8551
rect 1075 8520 2176 8548
rect 1075 8517 1087 8520
rect 1029 8511 1087 8517
rect 845 8483 903 8489
rect 845 8449 857 8483
rect 891 8480 903 8483
rect 1578 8480 1584 8492
rect 891 8452 1584 8480
rect 891 8449 903 8452
rect 845 8443 903 8449
rect 1578 8440 1584 8452
rect 1636 8440 1642 8492
rect 1670 8440 1676 8492
rect 1728 8440 1734 8492
rect 1946 8440 1952 8492
rect 2004 8480 2010 8492
rect 2041 8483 2099 8489
rect 2041 8480 2053 8483
rect 2004 8452 2053 8480
rect 2004 8440 2010 8452
rect 2041 8449 2053 8452
rect 2087 8449 2099 8483
rect 2041 8443 2099 8449
rect 1213 8415 1271 8421
rect 1213 8412 1225 8415
rect 768 8384 1225 8412
rect 1213 8381 1225 8384
rect 1259 8381 1271 8415
rect 1213 8375 1271 8381
rect 1305 8415 1363 8421
rect 1305 8381 1317 8415
rect 1351 8381 1363 8415
rect 1305 8375 1363 8381
rect 1765 8415 1823 8421
rect 1765 8381 1777 8415
rect 1811 8412 1823 8415
rect 1854 8412 1860 8424
rect 1811 8384 1860 8412
rect 1811 8381 1823 8384
rect 1765 8375 1823 8381
rect 1320 8276 1348 8375
rect 1854 8372 1860 8384
rect 1912 8372 1918 8424
rect 2148 8412 2176 8520
rect 2332 8480 2360 8588
rect 2590 8576 2596 8628
rect 2648 8576 2654 8628
rect 8113 8619 8171 8625
rect 8113 8585 8125 8619
rect 8159 8616 8171 8619
rect 8846 8616 8852 8628
rect 8159 8588 8852 8616
rect 8159 8585 8171 8588
rect 8113 8579 8171 8585
rect 8846 8576 8852 8588
rect 8904 8576 8910 8628
rect 10318 8576 10324 8628
rect 10376 8616 10382 8628
rect 10597 8619 10655 8625
rect 10597 8616 10609 8619
rect 10376 8588 10609 8616
rect 10376 8576 10382 8588
rect 10597 8585 10609 8588
rect 10643 8585 10655 8619
rect 10597 8579 10655 8585
rect 18046 8576 18052 8628
rect 18104 8616 18110 8628
rect 21729 8619 21787 8625
rect 18104 8588 18368 8616
rect 18104 8576 18110 8588
rect 2406 8508 2412 8560
rect 2464 8548 2470 8560
rect 2866 8548 2872 8560
rect 2464 8520 2872 8548
rect 2464 8508 2470 8520
rect 2866 8508 2872 8520
rect 2924 8508 2930 8560
rect 12894 8508 12900 8560
rect 12952 8508 12958 8560
rect 14093 8551 14151 8557
rect 14093 8517 14105 8551
rect 14139 8548 14151 8551
rect 14366 8548 14372 8560
rect 14139 8520 14372 8548
rect 14139 8517 14151 8520
rect 14093 8511 14151 8517
rect 14366 8508 14372 8520
rect 14424 8508 14430 8560
rect 16393 8551 16451 8557
rect 16393 8517 16405 8551
rect 16439 8548 16451 8551
rect 16850 8548 16856 8560
rect 16439 8520 16856 8548
rect 16439 8517 16451 8520
rect 16393 8511 16451 8517
rect 16850 8508 16856 8520
rect 16908 8508 16914 8560
rect 17589 8551 17647 8557
rect 17589 8517 17601 8551
rect 17635 8548 17647 8551
rect 18138 8548 18144 8560
rect 17635 8520 18144 8548
rect 17635 8517 17647 8520
rect 17589 8511 17647 8517
rect 18138 8508 18144 8520
rect 18196 8508 18202 8560
rect 2501 8483 2559 8489
rect 2501 8480 2513 8483
rect 2332 8452 2513 8480
rect 2501 8449 2513 8452
rect 2547 8449 2559 8483
rect 2501 8443 2559 8449
rect 11054 8440 11060 8492
rect 11112 8440 11118 8492
rect 12437 8483 12495 8489
rect 12437 8449 12449 8483
rect 12483 8480 12495 8483
rect 12526 8480 12532 8492
rect 12483 8452 12532 8480
rect 12483 8449 12495 8452
rect 12437 8443 12495 8449
rect 12526 8440 12532 8452
rect 12584 8440 12590 8492
rect 12618 8440 12624 8492
rect 12676 8480 12682 8492
rect 12912 8480 12940 8508
rect 12676 8452 12940 8480
rect 14740 8492 14792 8498
rect 12676 8440 12682 8452
rect 14740 8434 14792 8440
rect 2225 8415 2283 8421
rect 2225 8412 2237 8415
rect 2148 8384 2237 8412
rect 2225 8381 2237 8384
rect 2271 8381 2283 8415
rect 2225 8375 2283 8381
rect 2406 8372 2412 8424
rect 2464 8372 2470 8424
rect 2866 8372 2872 8424
rect 2924 8412 2930 8424
rect 3237 8415 3295 8421
rect 3237 8412 3249 8415
rect 2924 8384 3249 8412
rect 2924 8372 2930 8384
rect 3237 8381 3249 8384
rect 3283 8412 3295 8415
rect 5261 8415 5319 8421
rect 5261 8412 5273 8415
rect 3283 8384 5273 8412
rect 3283 8381 3295 8384
rect 3237 8375 3295 8381
rect 5261 8381 5273 8384
rect 5307 8381 5319 8415
rect 5261 8375 5319 8381
rect 6086 8372 6092 8424
rect 6144 8412 6150 8424
rect 6733 8415 6791 8421
rect 6733 8412 6745 8415
rect 6144 8384 6745 8412
rect 6144 8372 6150 8384
rect 6733 8381 6745 8384
rect 6779 8412 6791 8415
rect 9214 8412 9220 8424
rect 6779 8384 9220 8412
rect 6779 8381 6791 8384
rect 6733 8375 6791 8381
rect 9214 8372 9220 8384
rect 9272 8372 9278 8424
rect 10962 8372 10968 8424
rect 11020 8372 11026 8424
rect 12342 8372 12348 8424
rect 12400 8412 12406 8424
rect 12897 8415 12955 8421
rect 12897 8412 12909 8415
rect 12400 8384 12909 8412
rect 12400 8372 12406 8384
rect 12897 8381 12909 8384
rect 12943 8412 12955 8415
rect 13170 8412 13176 8424
rect 12943 8384 13176 8412
rect 12943 8381 12955 8384
rect 12897 8375 12955 8381
rect 13170 8372 13176 8384
rect 13228 8372 13234 8424
rect 13265 8415 13323 8421
rect 13265 8381 13277 8415
rect 13311 8381 13323 8415
rect 13265 8375 13323 8381
rect 2774 8304 2780 8356
rect 2832 8304 2838 8356
rect 2961 8347 3019 8353
rect 2961 8313 2973 8347
rect 3007 8344 3019 8347
rect 3050 8344 3056 8356
rect 3007 8316 3056 8344
rect 3007 8313 3019 8316
rect 2961 8307 3019 8313
rect 3050 8304 3056 8316
rect 3108 8304 3114 8356
rect 3142 8304 3148 8356
rect 3200 8344 3206 8356
rect 3482 8347 3540 8353
rect 3482 8344 3494 8347
rect 3200 8316 3494 8344
rect 3200 8304 3206 8316
rect 3482 8313 3494 8316
rect 3528 8313 3540 8347
rect 3482 8307 3540 8313
rect 5528 8347 5586 8353
rect 5528 8313 5540 8347
rect 5574 8344 5586 8347
rect 6362 8344 6368 8356
rect 5574 8316 6368 8344
rect 5574 8313 5586 8316
rect 5528 8307 5586 8313
rect 6362 8304 6368 8316
rect 6420 8304 6426 8356
rect 7000 8347 7058 8353
rect 7000 8313 7012 8347
rect 7046 8344 7058 8347
rect 8018 8344 8024 8356
rect 7046 8316 8024 8344
rect 7046 8313 7058 8316
rect 7000 8307 7058 8313
rect 8018 8304 8024 8316
rect 8076 8304 8082 8356
rect 9490 8353 9496 8356
rect 9484 8307 9496 8353
rect 9490 8304 9496 8307
rect 9548 8304 9554 8356
rect 12802 8304 12808 8356
rect 12860 8304 12866 8356
rect 13280 8344 13308 8375
rect 14458 8372 14464 8424
rect 14516 8372 14522 8424
rect 14918 8372 14924 8424
rect 14976 8372 14982 8424
rect 15473 8415 15531 8421
rect 15473 8381 15485 8415
rect 15519 8381 15531 8415
rect 15473 8375 15531 8381
rect 13722 8344 13728 8356
rect 13280 8316 13728 8344
rect 13722 8304 13728 8316
rect 13780 8344 13786 8356
rect 15488 8344 15516 8375
rect 16206 8372 16212 8424
rect 16264 8372 16270 8424
rect 17405 8415 17463 8421
rect 17405 8381 17417 8415
rect 17451 8412 17463 8415
rect 17586 8412 17592 8424
rect 17451 8384 17592 8412
rect 17451 8381 17463 8384
rect 17405 8375 17463 8381
rect 17586 8372 17592 8384
rect 17644 8372 17650 8424
rect 18340 8421 18368 8588
rect 21729 8585 21741 8619
rect 21775 8616 21787 8619
rect 21818 8616 21824 8628
rect 21775 8588 21824 8616
rect 21775 8585 21787 8588
rect 21729 8579 21787 8585
rect 21818 8576 21824 8588
rect 21876 8616 21882 8628
rect 22097 8619 22155 8625
rect 22097 8616 22109 8619
rect 21876 8588 22109 8616
rect 21876 8576 21882 8588
rect 22097 8585 22109 8588
rect 22143 8585 22155 8619
rect 22097 8579 22155 8585
rect 22922 8576 22928 8628
rect 22980 8576 22986 8628
rect 23937 8619 23995 8625
rect 23937 8616 23949 8619
rect 23400 8588 23949 8616
rect 22002 8548 22008 8560
rect 21100 8520 22008 8548
rect 19610 8440 19616 8492
rect 19668 8480 19674 8492
rect 20622 8480 20628 8492
rect 19668 8452 20628 8480
rect 19668 8440 19674 8452
rect 20622 8440 20628 8452
rect 20680 8440 20686 8492
rect 21100 8480 21128 8520
rect 22002 8508 22008 8520
rect 22060 8508 22066 8560
rect 23400 8548 23428 8588
rect 23937 8585 23949 8588
rect 23983 8585 23995 8619
rect 23937 8579 23995 8585
rect 24029 8619 24087 8625
rect 24029 8585 24041 8619
rect 24075 8616 24087 8619
rect 24210 8616 24216 8628
rect 24075 8588 24216 8616
rect 24075 8585 24087 8588
rect 24029 8579 24087 8585
rect 22848 8520 23428 8548
rect 23569 8551 23627 8557
rect 22848 8492 22876 8520
rect 23569 8517 23581 8551
rect 23615 8517 23627 8551
rect 23952 8548 23980 8579
rect 24210 8576 24216 8588
rect 24268 8576 24274 8628
rect 24394 8576 24400 8628
rect 24452 8616 24458 8628
rect 24452 8588 25452 8616
rect 24452 8576 24458 8588
rect 24305 8551 24363 8557
rect 24305 8548 24317 8551
rect 23952 8520 24317 8548
rect 23569 8511 23627 8517
rect 24305 8517 24317 8520
rect 24351 8517 24363 8551
rect 24305 8511 24363 8517
rect 21913 8483 21971 8489
rect 21913 8480 21925 8483
rect 21008 8452 21128 8480
rect 21836 8452 21925 8480
rect 18325 8415 18383 8421
rect 18325 8381 18337 8415
rect 18371 8381 18383 8415
rect 18325 8375 18383 8381
rect 18509 8415 18567 8421
rect 18509 8381 18521 8415
rect 18555 8412 18567 8415
rect 18598 8412 18604 8424
rect 18555 8384 18604 8412
rect 18555 8381 18567 8384
rect 18509 8375 18567 8381
rect 18598 8372 18604 8384
rect 18656 8372 18662 8424
rect 19150 8372 19156 8424
rect 19208 8372 19214 8424
rect 20438 8372 20444 8424
rect 20496 8372 20502 8424
rect 21008 8421 21036 8452
rect 20993 8415 21051 8421
rect 20993 8381 21005 8415
rect 21039 8381 21051 8415
rect 20993 8375 21051 8381
rect 21085 8415 21143 8421
rect 21085 8381 21097 8415
rect 21131 8412 21143 8415
rect 21634 8412 21640 8424
rect 21131 8384 21640 8412
rect 21131 8381 21143 8384
rect 21085 8375 21143 8381
rect 21634 8372 21640 8384
rect 21692 8372 21698 8424
rect 21836 8421 21864 8452
rect 21913 8449 21925 8452
rect 21959 8480 21971 8483
rect 22094 8480 22100 8492
rect 21959 8452 22100 8480
rect 21959 8449 21971 8452
rect 21913 8443 21971 8449
rect 22094 8440 22100 8452
rect 22152 8440 22158 8492
rect 22830 8440 22836 8492
rect 22888 8440 22894 8492
rect 23382 8480 23388 8492
rect 23216 8452 23388 8480
rect 21821 8415 21879 8421
rect 21821 8381 21833 8415
rect 21867 8381 21879 8415
rect 21821 8375 21879 8381
rect 22002 8372 22008 8424
rect 22060 8412 22066 8424
rect 22189 8415 22247 8421
rect 22189 8412 22201 8415
rect 22060 8384 22201 8412
rect 22060 8372 22066 8384
rect 22189 8381 22201 8384
rect 22235 8381 22247 8415
rect 22189 8375 22247 8381
rect 22848 8384 23060 8412
rect 19168 8344 19196 8372
rect 13780 8316 19196 8344
rect 20456 8344 20484 8372
rect 22848 8344 22876 8384
rect 20456 8316 22876 8344
rect 13780 8304 13786 8316
rect 22922 8304 22928 8356
rect 22980 8304 22986 8356
rect 23032 8344 23060 8384
rect 23106 8372 23112 8424
rect 23164 8372 23170 8424
rect 23216 8421 23244 8452
rect 23382 8440 23388 8452
rect 23440 8440 23446 8492
rect 23584 8480 23612 8511
rect 25130 8508 25136 8560
rect 25188 8508 25194 8560
rect 24121 8483 24179 8489
rect 24121 8480 24133 8483
rect 23584 8452 24133 8480
rect 24121 8449 24133 8452
rect 24167 8480 24179 8483
rect 24167 8452 24440 8480
rect 24167 8449 24179 8452
rect 24121 8443 24179 8449
rect 23201 8415 23259 8421
rect 23201 8381 23213 8415
rect 23247 8381 23259 8415
rect 23201 8375 23259 8381
rect 23474 8372 23480 8424
rect 23532 8372 23538 8424
rect 23566 8372 23572 8424
rect 23624 8412 23630 8424
rect 23661 8415 23719 8421
rect 23661 8412 23673 8415
rect 23624 8384 23673 8412
rect 23624 8372 23630 8384
rect 23661 8381 23673 8384
rect 23707 8381 23719 8415
rect 23661 8375 23719 8381
rect 23750 8372 23756 8424
rect 23808 8412 23814 8424
rect 23845 8415 23903 8421
rect 23845 8412 23857 8415
rect 23808 8384 23857 8412
rect 23808 8372 23814 8384
rect 23845 8381 23857 8384
rect 23891 8381 23903 8415
rect 23845 8375 23903 8381
rect 24210 8372 24216 8424
rect 24268 8372 24274 8424
rect 24412 8421 24440 8452
rect 24762 8440 24768 8492
rect 24820 8440 24826 8492
rect 25424 8489 25452 8588
rect 25409 8483 25467 8489
rect 25409 8449 25421 8483
rect 25455 8449 25467 8483
rect 25409 8443 25467 8449
rect 24397 8415 24455 8421
rect 24397 8381 24409 8415
rect 24443 8381 24455 8415
rect 24780 8412 24808 8440
rect 24397 8375 24455 8381
rect 24596 8384 24808 8412
rect 24596 8356 24624 8384
rect 25590 8372 25596 8424
rect 25648 8372 25654 8424
rect 24578 8344 24584 8356
rect 23032 8316 24584 8344
rect 24578 8304 24584 8316
rect 24636 8304 24642 8356
rect 24762 8304 24768 8356
rect 24820 8304 24826 8356
rect 25777 8347 25835 8353
rect 25777 8313 25789 8347
rect 25823 8344 25835 8347
rect 26234 8344 26240 8356
rect 25823 8316 26240 8344
rect 25823 8313 25835 8316
rect 25777 8307 25835 8313
rect 26234 8304 26240 8316
rect 26292 8304 26298 8356
rect 2406 8276 2412 8288
rect 1320 8248 2412 8276
rect 2406 8236 2412 8248
rect 2464 8236 2470 8288
rect 4154 8236 4160 8288
rect 4212 8276 4218 8288
rect 4614 8276 4620 8288
rect 4212 8248 4620 8276
rect 4212 8236 4218 8248
rect 4614 8236 4620 8248
rect 4672 8236 4678 8288
rect 6638 8236 6644 8288
rect 6696 8236 6702 8288
rect 11793 8279 11851 8285
rect 11793 8245 11805 8279
rect 11839 8276 11851 8279
rect 13354 8276 13360 8288
rect 11839 8248 13360 8276
rect 11839 8245 11851 8248
rect 11793 8239 11851 8245
rect 13354 8236 13360 8248
rect 13412 8236 13418 8288
rect 13630 8236 13636 8288
rect 13688 8276 13694 8288
rect 15010 8276 15016 8288
rect 13688 8248 15016 8276
rect 13688 8236 13694 8248
rect 15010 8236 15016 8248
rect 15068 8276 15074 8288
rect 18046 8276 18052 8288
rect 15068 8248 18052 8276
rect 15068 8236 15074 8248
rect 18046 8236 18052 8248
rect 18104 8236 18110 8288
rect 18414 8236 18420 8288
rect 18472 8236 18478 8288
rect 19153 8279 19211 8285
rect 19153 8245 19165 8279
rect 19199 8276 19211 8279
rect 19426 8276 19432 8288
rect 19199 8248 19432 8276
rect 19199 8245 19211 8248
rect 19153 8239 19211 8245
rect 19426 8236 19432 8248
rect 19484 8236 19490 8288
rect 20898 8236 20904 8288
rect 20956 8236 20962 8288
rect 21361 8279 21419 8285
rect 21361 8245 21373 8279
rect 21407 8276 21419 8279
rect 21634 8276 21640 8288
rect 21407 8248 21640 8276
rect 21407 8245 21419 8248
rect 21361 8239 21419 8245
rect 21634 8236 21640 8248
rect 21692 8236 21698 8288
rect 21910 8236 21916 8288
rect 21968 8236 21974 8288
rect 25222 8236 25228 8288
rect 25280 8236 25286 8288
rect 552 8186 27576 8208
rect 552 8134 7114 8186
rect 7166 8134 7178 8186
rect 7230 8134 7242 8186
rect 7294 8134 7306 8186
rect 7358 8134 7370 8186
rect 7422 8134 13830 8186
rect 13882 8134 13894 8186
rect 13946 8134 13958 8186
rect 14010 8134 14022 8186
rect 14074 8134 14086 8186
rect 14138 8134 20546 8186
rect 20598 8134 20610 8186
rect 20662 8134 20674 8186
rect 20726 8134 20738 8186
rect 20790 8134 20802 8186
rect 20854 8134 27262 8186
rect 27314 8134 27326 8186
rect 27378 8134 27390 8186
rect 27442 8134 27454 8186
rect 27506 8134 27518 8186
rect 27570 8134 27576 8186
rect 552 8112 27576 8134
rect 2130 8032 2136 8084
rect 2188 8072 2194 8084
rect 3237 8075 3295 8081
rect 3237 8072 3249 8075
rect 2188 8044 3249 8072
rect 2188 8032 2194 8044
rect 3237 8041 3249 8044
rect 3283 8041 3295 8075
rect 4801 8075 4859 8081
rect 3237 8035 3295 8041
rect 3804 8044 4752 8072
rect 2501 8007 2559 8013
rect 2501 7973 2513 8007
rect 2547 8004 2559 8007
rect 2869 8007 2927 8013
rect 2869 8004 2881 8007
rect 2547 7976 2881 8004
rect 2547 7973 2559 7976
rect 2501 7967 2559 7973
rect 2869 7973 2881 7976
rect 2915 7973 2927 8007
rect 2869 7967 2927 7973
rect 3050 7964 3056 8016
rect 3108 7964 3114 8016
rect 3326 7964 3332 8016
rect 3384 8004 3390 8016
rect 3421 8007 3479 8013
rect 3421 8004 3433 8007
rect 3384 7976 3433 8004
rect 3384 7964 3390 7976
rect 3421 7973 3433 7976
rect 3467 7973 3479 8007
rect 3421 7967 3479 7973
rect 3510 7964 3516 8016
rect 3568 8004 3574 8016
rect 3804 8013 3832 8044
rect 3605 8007 3663 8013
rect 3605 8004 3617 8007
rect 3568 7976 3617 8004
rect 3568 7964 3574 7976
rect 3605 7973 3617 7976
rect 3651 7973 3663 8007
rect 3605 7967 3663 7973
rect 3789 8007 3847 8013
rect 3789 7973 3801 8007
rect 3835 7973 3847 8007
rect 3789 7967 3847 7973
rect 3896 7976 4492 8004
rect 2777 7939 2835 7945
rect 2777 7905 2789 7939
rect 2823 7936 2835 7939
rect 3068 7936 3096 7964
rect 2823 7908 3096 7936
rect 3145 7939 3203 7945
rect 2823 7905 2835 7908
rect 2777 7899 2835 7905
rect 3145 7905 3157 7939
rect 3191 7936 3203 7939
rect 3234 7936 3240 7948
rect 3191 7908 3240 7936
rect 3191 7905 3203 7908
rect 3145 7899 3203 7905
rect 3234 7896 3240 7908
rect 3292 7896 3298 7948
rect 2501 7871 2559 7877
rect 2501 7837 2513 7871
rect 2547 7868 2559 7871
rect 2958 7868 2964 7880
rect 2547 7840 2964 7868
rect 2547 7837 2559 7840
rect 2501 7831 2559 7837
rect 2958 7828 2964 7840
rect 3016 7828 3022 7880
rect 2869 7803 2927 7809
rect 2869 7769 2881 7803
rect 2915 7800 2927 7803
rect 3142 7800 3148 7812
rect 2915 7772 3148 7800
rect 2915 7769 2927 7772
rect 2869 7763 2927 7769
rect 3142 7760 3148 7772
rect 3200 7760 3206 7812
rect 2685 7735 2743 7741
rect 2685 7701 2697 7735
rect 2731 7732 2743 7735
rect 3252 7732 3280 7896
rect 3602 7828 3608 7880
rect 3660 7868 3666 7880
rect 3896 7868 3924 7976
rect 3973 7939 4031 7945
rect 3973 7905 3985 7939
rect 4019 7905 4031 7939
rect 3973 7899 4031 7905
rect 3660 7840 3924 7868
rect 3660 7828 3666 7840
rect 3988 7800 4016 7899
rect 4154 7896 4160 7948
rect 4212 7896 4218 7948
rect 4464 7945 4492 7976
rect 4433 7939 4492 7945
rect 4433 7905 4445 7939
rect 4479 7912 4492 7939
rect 4724 7936 4752 8044
rect 4801 8041 4813 8075
rect 4847 8041 4859 8075
rect 4801 8035 4859 8041
rect 4816 8004 4844 8035
rect 6362 8032 6368 8084
rect 6420 8032 6426 8084
rect 9490 8032 9496 8084
rect 9548 8032 9554 8084
rect 9674 8032 9680 8084
rect 9732 8032 9738 8084
rect 12526 8032 12532 8084
rect 12584 8032 12590 8084
rect 14182 8032 14188 8084
rect 14240 8032 14246 8084
rect 14918 8072 14924 8084
rect 14292 8044 14924 8072
rect 4816 7976 5396 8004
rect 4893 7939 4951 7945
rect 4893 7936 4905 7939
rect 4479 7905 4491 7912
rect 4724 7908 4905 7936
rect 4433 7899 4491 7905
rect 4893 7905 4905 7908
rect 4939 7905 4951 7939
rect 4893 7899 4951 7905
rect 5074 7896 5080 7948
rect 5132 7896 5138 7948
rect 5368 7945 5396 7976
rect 5353 7939 5411 7945
rect 5353 7905 5365 7939
rect 5399 7905 5411 7939
rect 5353 7899 5411 7905
rect 6549 7939 6607 7945
rect 6549 7905 6561 7939
rect 6595 7936 6607 7939
rect 6641 7939 6699 7945
rect 6641 7936 6653 7939
rect 6595 7908 6653 7936
rect 6595 7905 6607 7908
rect 6549 7899 6607 7905
rect 6641 7905 6653 7908
rect 6687 7905 6699 7939
rect 6641 7899 6699 7905
rect 6822 7896 6828 7948
rect 6880 7896 6886 7948
rect 9692 7945 9720 8032
rect 12434 8004 12440 8016
rect 12268 7976 12440 8004
rect 9677 7939 9735 7945
rect 9677 7905 9689 7939
rect 9723 7905 9735 7939
rect 9677 7899 9735 7905
rect 11882 7896 11888 7948
rect 11940 7896 11946 7948
rect 12268 7945 12296 7976
rect 12434 7964 12440 7976
rect 12492 7964 12498 8016
rect 12544 8004 12572 8032
rect 12544 7976 12664 8004
rect 11977 7939 12035 7945
rect 11977 7905 11989 7939
rect 12023 7905 12035 7939
rect 11977 7899 12035 7905
rect 12253 7939 12311 7945
rect 12253 7905 12265 7939
rect 12299 7905 12311 7939
rect 12253 7899 12311 7905
rect 4338 7828 4344 7880
rect 4396 7828 4402 7880
rect 5537 7871 5595 7877
rect 5537 7837 5549 7871
rect 5583 7868 5595 7871
rect 7009 7871 7067 7877
rect 7009 7868 7021 7871
rect 5583 7840 7021 7868
rect 5583 7837 5595 7840
rect 5537 7831 5595 7837
rect 7009 7837 7021 7840
rect 7055 7868 7067 7871
rect 8846 7868 8852 7880
rect 7055 7840 8852 7868
rect 7055 7837 7067 7840
rect 7009 7831 7067 7837
rect 8846 7828 8852 7840
rect 8904 7828 8910 7880
rect 11517 7871 11575 7877
rect 11517 7837 11529 7871
rect 11563 7837 11575 7871
rect 11992 7868 12020 7899
rect 12342 7896 12348 7948
rect 12400 7896 12406 7948
rect 12526 7896 12532 7948
rect 12584 7896 12590 7948
rect 12636 7945 12664 7976
rect 14200 7945 14228 8032
rect 14292 7945 14320 8044
rect 14918 8032 14924 8044
rect 14976 8032 14982 8084
rect 18414 8032 18420 8084
rect 18472 8072 18478 8084
rect 18472 8044 19104 8072
rect 18472 8032 18478 8044
rect 14476 7976 15148 8004
rect 14476 7945 14504 7976
rect 15120 7948 15148 7976
rect 16850 7964 16856 8016
rect 16908 7964 16914 8016
rect 17034 7964 17040 8016
rect 17092 8004 17098 8016
rect 17092 7976 19012 8004
rect 17092 7964 17098 7976
rect 12621 7939 12679 7945
rect 12621 7905 12633 7939
rect 12667 7905 12679 7939
rect 12621 7899 12679 7905
rect 14185 7939 14243 7945
rect 14185 7905 14197 7939
rect 14231 7905 14243 7939
rect 14185 7899 14243 7905
rect 14277 7939 14335 7945
rect 14277 7905 14289 7939
rect 14323 7905 14335 7939
rect 14277 7899 14335 7905
rect 14461 7939 14519 7945
rect 14461 7905 14473 7939
rect 14507 7905 14519 7939
rect 14461 7899 14519 7905
rect 14550 7896 14556 7948
rect 14608 7896 14614 7948
rect 14826 7896 14832 7948
rect 14884 7896 14890 7948
rect 15102 7896 15108 7948
rect 15160 7896 15166 7948
rect 15194 7896 15200 7948
rect 15252 7936 15258 7948
rect 15473 7939 15531 7945
rect 15473 7936 15485 7939
rect 15252 7908 15485 7936
rect 15252 7896 15258 7908
rect 15473 7905 15485 7908
rect 15519 7905 15531 7939
rect 16868 7936 16896 7964
rect 17512 7945 17540 7976
rect 17230 7939 17288 7945
rect 17230 7936 17242 7939
rect 16868 7908 17242 7936
rect 15473 7899 15531 7905
rect 17230 7905 17242 7908
rect 17276 7905 17288 7939
rect 17230 7899 17288 7905
rect 17497 7939 17555 7945
rect 17497 7905 17509 7939
rect 17543 7905 17555 7939
rect 17497 7899 17555 7905
rect 18138 7896 18144 7948
rect 18196 7936 18202 7948
rect 18702 7939 18760 7945
rect 18702 7936 18714 7939
rect 18196 7908 18714 7936
rect 18196 7896 18202 7908
rect 18702 7905 18714 7908
rect 18748 7905 18760 7939
rect 18702 7899 18760 7905
rect 12158 7868 12164 7880
rect 11992 7840 12164 7868
rect 11517 7831 11575 7837
rect 4430 7800 4436 7812
rect 3988 7772 4436 7800
rect 4430 7760 4436 7772
rect 4488 7760 4494 7812
rect 11532 7800 11560 7831
rect 12158 7828 12164 7840
rect 12216 7868 12222 7880
rect 12894 7868 12900 7880
rect 12216 7840 12900 7868
rect 12216 7828 12222 7840
rect 12894 7828 12900 7840
rect 12952 7828 12958 7880
rect 14921 7871 14979 7877
rect 14921 7837 14933 7871
rect 14967 7837 14979 7871
rect 14921 7831 14979 7837
rect 14550 7800 14556 7812
rect 4908 7772 14556 7800
rect 2731 7704 3280 7732
rect 2731 7701 2743 7704
rect 2685 7695 2743 7701
rect 4246 7692 4252 7744
rect 4304 7732 4310 7744
rect 4908 7732 4936 7772
rect 14550 7760 14556 7772
rect 14608 7760 14614 7812
rect 14936 7800 14964 7831
rect 15378 7828 15384 7880
rect 15436 7828 15442 7880
rect 18984 7877 19012 7976
rect 19076 7948 19104 8044
rect 19150 8032 19156 8084
rect 19208 8032 19214 8084
rect 20898 8032 20904 8084
rect 20956 8032 20962 8084
rect 21818 8032 21824 8084
rect 21876 8072 21882 8084
rect 21913 8075 21971 8081
rect 21913 8072 21925 8075
rect 21876 8044 21925 8072
rect 21876 8032 21882 8044
rect 21913 8041 21925 8044
rect 21959 8041 21971 8075
rect 21913 8035 21971 8041
rect 22094 8032 22100 8084
rect 22152 8072 22158 8084
rect 22189 8075 22247 8081
rect 22189 8072 22201 8075
rect 22152 8044 22201 8072
rect 22152 8032 22158 8044
rect 22189 8041 22201 8044
rect 22235 8041 22247 8075
rect 22189 8035 22247 8041
rect 22646 8032 22652 8084
rect 22704 8072 22710 8084
rect 22741 8075 22799 8081
rect 22741 8072 22753 8075
rect 22704 8044 22753 8072
rect 22704 8032 22710 8044
rect 22741 8041 22753 8044
rect 22787 8072 22799 8075
rect 23750 8072 23756 8084
rect 22787 8044 23756 8072
rect 22787 8041 22799 8044
rect 22741 8035 22799 8041
rect 19168 8004 19196 8032
rect 20916 8004 20944 8032
rect 22557 8007 22615 8013
rect 19168 7976 19472 8004
rect 20916 7976 21496 8004
rect 19058 7896 19064 7948
rect 19116 7896 19122 7948
rect 19153 7939 19211 7945
rect 19153 7905 19165 7939
rect 19199 7936 19211 7939
rect 19242 7936 19248 7948
rect 19199 7908 19248 7936
rect 19199 7905 19211 7908
rect 19153 7899 19211 7905
rect 19242 7896 19248 7908
rect 19300 7896 19306 7948
rect 19334 7896 19340 7948
rect 19392 7896 19398 7948
rect 19444 7945 19472 7976
rect 21468 7945 21496 7976
rect 21744 7976 21956 8004
rect 19429 7939 19487 7945
rect 19429 7905 19441 7939
rect 19475 7905 19487 7939
rect 19429 7899 19487 7905
rect 19972 7939 20030 7945
rect 19972 7905 19984 7939
rect 20018 7936 20030 7939
rect 21269 7939 21327 7945
rect 21269 7936 21281 7939
rect 20018 7908 21281 7936
rect 20018 7905 20030 7908
rect 19972 7899 20030 7905
rect 21269 7905 21281 7908
rect 21315 7905 21327 7939
rect 21269 7899 21327 7905
rect 21453 7939 21511 7945
rect 21453 7905 21465 7939
rect 21499 7905 21511 7939
rect 21453 7899 21511 7905
rect 21634 7896 21640 7948
rect 21692 7896 21698 7948
rect 21744 7945 21772 7976
rect 21928 7948 21956 7976
rect 22020 7976 22324 8004
rect 21729 7939 21787 7945
rect 21729 7905 21741 7939
rect 21775 7905 21787 7939
rect 21729 7899 21787 7905
rect 21821 7939 21879 7945
rect 21821 7905 21833 7939
rect 21867 7905 21879 7939
rect 21821 7899 21879 7905
rect 18969 7871 19027 7877
rect 18969 7837 18981 7871
rect 19015 7868 19027 7871
rect 19705 7871 19763 7877
rect 19705 7868 19717 7871
rect 19015 7840 19717 7868
rect 19015 7837 19027 7840
rect 18969 7831 19027 7837
rect 19444 7812 19472 7840
rect 19705 7837 19717 7840
rect 19751 7837 19763 7871
rect 19705 7831 19763 7837
rect 21836 7868 21864 7899
rect 21910 7896 21916 7948
rect 21968 7896 21974 7948
rect 22020 7945 22048 7976
rect 22296 7945 22324 7976
rect 22557 7973 22569 8007
rect 22603 8004 22615 8007
rect 22925 8007 22983 8013
rect 22925 8004 22937 8007
rect 22603 7976 22937 8004
rect 22603 7973 22615 7976
rect 22557 7967 22615 7973
rect 22925 7973 22937 7976
rect 22971 7973 22983 8007
rect 23124 8004 23152 8044
rect 23750 8032 23756 8044
rect 23808 8032 23814 8084
rect 23845 8075 23903 8081
rect 23845 8041 23857 8075
rect 23891 8072 23903 8075
rect 24210 8072 24216 8084
rect 23891 8044 24216 8072
rect 23891 8041 23903 8044
rect 23845 8035 23903 8041
rect 24210 8032 24216 8044
rect 24268 8032 24274 8084
rect 25958 8032 25964 8084
rect 26016 8032 26022 8084
rect 26234 8032 26240 8084
rect 26292 8072 26298 8084
rect 26292 8044 26648 8072
rect 26292 8032 26298 8044
rect 23124 7976 23244 8004
rect 22925 7967 22983 7973
rect 22005 7939 22063 7945
rect 22005 7905 22017 7939
rect 22051 7905 22063 7939
rect 22005 7899 22063 7905
rect 22097 7939 22155 7945
rect 22097 7905 22109 7939
rect 22143 7905 22155 7939
rect 22097 7899 22155 7905
rect 22281 7939 22339 7945
rect 22281 7905 22293 7939
rect 22327 7936 22339 7939
rect 22462 7936 22468 7948
rect 22327 7908 22468 7936
rect 22327 7905 22339 7908
rect 22281 7899 22339 7905
rect 22112 7868 22140 7899
rect 22462 7896 22468 7908
rect 22520 7896 22526 7948
rect 22738 7896 22744 7948
rect 22796 7896 22802 7948
rect 22830 7896 22836 7948
rect 22888 7936 22894 7948
rect 23216 7945 23244 7976
rect 23474 7964 23480 8016
rect 23532 7964 23538 8016
rect 23109 7939 23167 7945
rect 23109 7936 23121 7939
rect 22888 7908 23121 7936
rect 22888 7896 22894 7908
rect 23109 7905 23121 7908
rect 23155 7905 23167 7939
rect 23109 7899 23167 7905
rect 23201 7939 23259 7945
rect 23201 7905 23213 7939
rect 23247 7905 23259 7939
rect 23201 7899 23259 7905
rect 23566 7896 23572 7948
rect 23624 7936 23630 7948
rect 23661 7939 23719 7945
rect 23661 7936 23673 7939
rect 23624 7908 23673 7936
rect 23624 7896 23630 7908
rect 23661 7905 23673 7908
rect 23707 7905 23719 7939
rect 23661 7899 23719 7905
rect 21836 7840 22140 7868
rect 22756 7868 22784 7896
rect 22925 7871 22983 7877
rect 22925 7868 22937 7871
rect 22756 7840 22937 7868
rect 15010 7800 15016 7812
rect 14936 7772 15016 7800
rect 15010 7760 15016 7772
rect 15068 7800 15074 7812
rect 16117 7803 16175 7809
rect 16117 7800 16129 7803
rect 15068 7772 16129 7800
rect 15068 7760 15074 7772
rect 16117 7769 16129 7772
rect 16163 7769 16175 7803
rect 16117 7763 16175 7769
rect 19426 7760 19432 7812
rect 19484 7760 19490 7812
rect 21085 7803 21143 7809
rect 21085 7769 21097 7803
rect 21131 7800 21143 7803
rect 21836 7800 21864 7840
rect 22925 7837 22937 7840
rect 22971 7837 22983 7871
rect 22925 7831 22983 7837
rect 21131 7772 21864 7800
rect 21131 7769 21143 7772
rect 21085 7763 21143 7769
rect 4304 7704 4936 7732
rect 4304 7692 4310 7704
rect 4982 7692 4988 7744
rect 5040 7692 5046 7744
rect 5166 7692 5172 7744
rect 5224 7692 5230 7744
rect 11698 7692 11704 7744
rect 11756 7692 11762 7744
rect 12069 7735 12127 7741
rect 12069 7701 12081 7735
rect 12115 7732 12127 7735
rect 12342 7732 12348 7744
rect 12115 7704 12348 7732
rect 12115 7701 12127 7704
rect 12069 7695 12127 7701
rect 12342 7692 12348 7704
rect 12400 7692 12406 7744
rect 14001 7735 14059 7741
rect 14001 7701 14013 7735
rect 14047 7732 14059 7735
rect 14182 7732 14188 7744
rect 14047 7704 14188 7732
rect 14047 7701 14059 7704
rect 14001 7695 14059 7701
rect 14182 7692 14188 7704
rect 14240 7692 14246 7744
rect 15105 7735 15163 7741
rect 15105 7701 15117 7735
rect 15151 7732 15163 7735
rect 15194 7732 15200 7744
rect 15151 7704 15200 7732
rect 15151 7701 15163 7704
rect 15105 7695 15163 7701
rect 15194 7692 15200 7704
rect 15252 7692 15258 7744
rect 15746 7692 15752 7744
rect 15804 7692 15810 7744
rect 16850 7692 16856 7744
rect 16908 7732 16914 7744
rect 17589 7735 17647 7741
rect 17589 7732 17601 7735
rect 16908 7704 17601 7732
rect 16908 7692 16914 7704
rect 17589 7701 17601 7704
rect 17635 7701 17647 7735
rect 17589 7695 17647 7701
rect 19613 7735 19671 7741
rect 19613 7701 19625 7735
rect 19659 7732 19671 7735
rect 20438 7732 20444 7744
rect 19659 7704 20444 7732
rect 19659 7701 19671 7704
rect 19613 7695 19671 7701
rect 20438 7692 20444 7704
rect 20496 7692 20502 7744
rect 22554 7692 22560 7744
rect 22612 7692 22618 7744
rect 23768 7732 23796 8032
rect 24121 8007 24179 8013
rect 24121 7973 24133 8007
rect 24167 8004 24179 8007
rect 24762 8004 24768 8016
rect 24167 7976 24768 8004
rect 24167 7973 24179 7976
rect 24121 7967 24179 7973
rect 24762 7964 24768 7976
rect 24820 7964 24826 8016
rect 25976 8004 26004 8032
rect 25976 7976 26280 8004
rect 24029 7939 24087 7945
rect 24029 7905 24041 7939
rect 24075 7905 24087 7939
rect 24029 7899 24087 7905
rect 24213 7939 24271 7945
rect 24213 7905 24225 7939
rect 24259 7936 24271 7939
rect 24489 7939 24547 7945
rect 24259 7908 24440 7936
rect 24259 7905 24271 7908
rect 24213 7899 24271 7905
rect 24044 7868 24072 7899
rect 24302 7868 24308 7880
rect 24044 7840 24308 7868
rect 24302 7828 24308 7840
rect 24360 7828 24366 7880
rect 24412 7800 24440 7908
rect 24489 7905 24501 7939
rect 24535 7936 24547 7939
rect 25130 7936 25136 7948
rect 24535 7908 25136 7936
rect 24535 7905 24547 7908
rect 24489 7899 24547 7905
rect 25130 7896 25136 7908
rect 25188 7936 25194 7948
rect 25498 7936 25504 7948
rect 25188 7908 25504 7936
rect 25188 7896 25194 7908
rect 25498 7896 25504 7908
rect 25556 7896 25562 7948
rect 26252 7945 26280 7976
rect 26620 7945 26648 8044
rect 25981 7939 26039 7945
rect 25981 7905 25993 7939
rect 26027 7936 26039 7939
rect 26237 7939 26295 7945
rect 26027 7908 26188 7936
rect 26027 7905 26039 7908
rect 25981 7899 26039 7905
rect 24765 7871 24823 7877
rect 24765 7837 24777 7871
rect 24811 7868 24823 7871
rect 25038 7868 25044 7880
rect 24811 7840 25044 7868
rect 24811 7837 24823 7840
rect 24765 7831 24823 7837
rect 25038 7828 25044 7840
rect 25096 7828 25102 7880
rect 26160 7868 26188 7908
rect 26237 7905 26249 7939
rect 26283 7905 26295 7939
rect 26237 7899 26295 7905
rect 26605 7939 26663 7945
rect 26605 7905 26617 7939
rect 26651 7905 26663 7939
rect 26605 7899 26663 7905
rect 26160 7840 26464 7868
rect 26436 7809 26464 7840
rect 26421 7803 26479 7809
rect 24412 7772 24900 7800
rect 24305 7735 24363 7741
rect 24305 7732 24317 7735
rect 23768 7704 24317 7732
rect 24305 7701 24317 7704
rect 24351 7701 24363 7735
rect 24305 7695 24363 7701
rect 24673 7735 24731 7741
rect 24673 7701 24685 7735
rect 24719 7732 24731 7735
rect 24762 7732 24768 7744
rect 24719 7704 24768 7732
rect 24719 7701 24731 7704
rect 24673 7695 24731 7701
rect 24762 7692 24768 7704
rect 24820 7692 24826 7744
rect 24872 7741 24900 7772
rect 26421 7769 26433 7803
rect 26467 7769 26479 7803
rect 26421 7763 26479 7769
rect 24857 7735 24915 7741
rect 24857 7701 24869 7735
rect 24903 7732 24915 7735
rect 25314 7732 25320 7744
rect 24903 7704 25320 7732
rect 24903 7701 24915 7704
rect 24857 7695 24915 7701
rect 25314 7692 25320 7704
rect 25372 7692 25378 7744
rect 552 7642 27416 7664
rect 552 7590 3756 7642
rect 3808 7590 3820 7642
rect 3872 7590 3884 7642
rect 3936 7590 3948 7642
rect 4000 7590 4012 7642
rect 4064 7590 10472 7642
rect 10524 7590 10536 7642
rect 10588 7590 10600 7642
rect 10652 7590 10664 7642
rect 10716 7590 10728 7642
rect 10780 7590 17188 7642
rect 17240 7590 17252 7642
rect 17304 7590 17316 7642
rect 17368 7590 17380 7642
rect 17432 7590 17444 7642
rect 17496 7590 23904 7642
rect 23956 7590 23968 7642
rect 24020 7590 24032 7642
rect 24084 7590 24096 7642
rect 24148 7590 24160 7642
rect 24212 7590 27416 7642
rect 552 7568 27416 7590
rect 2406 7488 2412 7540
rect 2464 7488 2470 7540
rect 3234 7488 3240 7540
rect 3292 7528 3298 7540
rect 4249 7531 4307 7537
rect 3292 7500 4200 7528
rect 3292 7488 3298 7500
rect 3528 7469 3556 7500
rect 4172 7472 4200 7500
rect 4249 7497 4261 7531
rect 4295 7528 4307 7531
rect 4338 7528 4344 7540
rect 4295 7500 4344 7528
rect 4295 7497 4307 7500
rect 4249 7491 4307 7497
rect 4338 7488 4344 7500
rect 4396 7488 4402 7540
rect 4525 7531 4583 7537
rect 4525 7497 4537 7531
rect 4571 7528 4583 7531
rect 5074 7528 5080 7540
rect 4571 7500 5080 7528
rect 4571 7497 4583 7500
rect 4525 7491 4583 7497
rect 3513 7463 3571 7469
rect 3513 7429 3525 7463
rect 3559 7429 3571 7463
rect 3513 7423 3571 7429
rect 3602 7420 3608 7472
rect 3660 7420 3666 7472
rect 4154 7420 4160 7472
rect 4212 7420 4218 7472
rect 1397 7395 1455 7401
rect 1397 7361 1409 7395
rect 1443 7392 1455 7395
rect 1578 7392 1584 7404
rect 1443 7364 1584 7392
rect 1443 7361 1455 7364
rect 1397 7355 1455 7361
rect 1578 7352 1584 7364
rect 1636 7392 1642 7404
rect 4246 7392 4252 7404
rect 1636 7364 4252 7392
rect 1636 7352 1642 7364
rect 4246 7352 4252 7364
rect 4304 7352 4310 7404
rect 4341 7395 4399 7401
rect 4341 7361 4353 7395
rect 4387 7392 4399 7395
rect 4540 7392 4568 7491
rect 5074 7488 5080 7500
rect 5132 7488 5138 7540
rect 5166 7488 5172 7540
rect 5224 7488 5230 7540
rect 6641 7531 6699 7537
rect 6641 7497 6653 7531
rect 6687 7528 6699 7531
rect 6822 7528 6828 7540
rect 6687 7500 6828 7528
rect 6687 7497 6699 7500
rect 6641 7491 6699 7497
rect 6822 7488 6828 7500
rect 6880 7488 6886 7540
rect 11698 7488 11704 7540
rect 11756 7528 11762 7540
rect 11756 7500 12756 7528
rect 11756 7488 11762 7500
rect 4614 7420 4620 7472
rect 4672 7420 4678 7472
rect 4387 7364 4568 7392
rect 4387 7361 4399 7364
rect 4341 7355 4399 7361
rect 1854 7284 1860 7336
rect 1912 7284 1918 7336
rect 2130 7284 2136 7336
rect 2188 7284 2194 7336
rect 2317 7327 2375 7333
rect 2317 7293 2329 7327
rect 2363 7324 2375 7327
rect 3237 7327 3295 7333
rect 3237 7324 3249 7327
rect 2363 7296 3249 7324
rect 2363 7293 2375 7296
rect 2317 7287 2375 7293
rect 3237 7293 3249 7296
rect 3283 7293 3295 7327
rect 3237 7287 3295 7293
rect 3421 7327 3479 7333
rect 3421 7293 3433 7327
rect 3467 7293 3479 7327
rect 3421 7287 3479 7293
rect 1762 7216 1768 7268
rect 1820 7256 1826 7268
rect 2332 7256 2360 7287
rect 1820 7228 2360 7256
rect 1820 7216 1826 7228
rect 2498 7216 2504 7268
rect 2556 7216 2562 7268
rect 3050 7216 3056 7268
rect 3108 7256 3114 7268
rect 3436 7256 3464 7287
rect 3694 7284 3700 7336
rect 3752 7284 3758 7336
rect 4065 7327 4123 7333
rect 4065 7293 4077 7327
rect 4111 7293 4123 7327
rect 4065 7287 4123 7293
rect 4080 7256 4108 7287
rect 4154 7284 4160 7336
rect 4212 7284 4218 7336
rect 4433 7327 4491 7333
rect 4433 7293 4445 7327
rect 4479 7324 4491 7327
rect 4522 7324 4528 7336
rect 4479 7296 4528 7324
rect 4479 7293 4491 7296
rect 4433 7287 4491 7293
rect 4522 7284 4528 7296
rect 4580 7284 4586 7336
rect 4632 7333 4660 7420
rect 4617 7327 4675 7333
rect 4617 7293 4629 7327
rect 4663 7293 4675 7327
rect 5184 7324 5212 7488
rect 7006 7352 7012 7404
rect 7064 7352 7070 7404
rect 8846 7352 8852 7404
rect 8904 7392 8910 7404
rect 12618 7392 12624 7404
rect 8904 7364 10456 7392
rect 8904 7352 8910 7364
rect 5261 7327 5319 7333
rect 5261 7324 5273 7327
rect 5184 7296 5273 7324
rect 4617 7287 4675 7293
rect 5261 7293 5273 7296
rect 5307 7293 5319 7327
rect 5261 7287 5319 7293
rect 6914 7284 6920 7336
rect 6972 7284 6978 7336
rect 8662 7284 8668 7336
rect 8720 7284 8726 7336
rect 10134 7284 10140 7336
rect 10192 7284 10198 7336
rect 10229 7327 10287 7333
rect 10229 7293 10241 7327
rect 10275 7293 10287 7327
rect 10229 7287 10287 7293
rect 7466 7256 7472 7268
rect 3108 7228 7472 7256
rect 3108 7216 3114 7228
rect 7466 7216 7472 7228
rect 7524 7216 7530 7268
rect 9858 7216 9864 7268
rect 9916 7216 9922 7268
rect 1670 7148 1676 7200
rect 1728 7148 1734 7200
rect 4154 7148 4160 7200
rect 4212 7188 4218 7200
rect 4982 7188 4988 7200
rect 4212 7160 4988 7188
rect 4212 7148 4218 7160
rect 4982 7148 4988 7160
rect 5040 7148 5046 7200
rect 5350 7148 5356 7200
rect 5408 7188 5414 7200
rect 5445 7191 5503 7197
rect 5445 7188 5457 7191
rect 5408 7160 5457 7188
rect 5408 7148 5414 7160
rect 5445 7157 5457 7160
rect 5491 7157 5503 7191
rect 5445 7151 5503 7157
rect 8478 7148 8484 7200
rect 8536 7148 8542 7200
rect 9674 7148 9680 7200
rect 9732 7188 9738 7200
rect 10244 7188 10272 7287
rect 10318 7284 10324 7336
rect 10376 7284 10382 7336
rect 10428 7256 10456 7364
rect 12360 7364 12624 7392
rect 10502 7284 10508 7336
rect 10560 7324 10566 7336
rect 12360 7324 12388 7364
rect 12618 7352 12624 7364
rect 12676 7352 12682 7404
rect 10560 7296 12388 7324
rect 10560 7284 10566 7296
rect 12434 7284 12440 7336
rect 12492 7284 12498 7336
rect 12728 7333 12756 7500
rect 12894 7488 12900 7540
rect 12952 7488 12958 7540
rect 13630 7488 13636 7540
rect 13688 7488 13694 7540
rect 14550 7488 14556 7540
rect 14608 7488 14614 7540
rect 15746 7488 15752 7540
rect 15804 7488 15810 7540
rect 16206 7488 16212 7540
rect 16264 7528 16270 7540
rect 16301 7531 16359 7537
rect 16301 7528 16313 7531
rect 16264 7500 16313 7528
rect 16264 7488 16270 7500
rect 16301 7497 16313 7500
rect 16347 7497 16359 7531
rect 16301 7491 16359 7497
rect 17586 7488 17592 7540
rect 17644 7488 17650 7540
rect 18046 7488 18052 7540
rect 18104 7528 18110 7540
rect 18104 7500 23428 7528
rect 18104 7488 18110 7500
rect 13648 7392 13676 7488
rect 12912 7364 13676 7392
rect 12713 7327 12771 7333
rect 12713 7293 12725 7327
rect 12759 7293 12771 7327
rect 12713 7287 12771 7293
rect 12192 7259 12250 7265
rect 10428 7228 11192 7256
rect 9732 7160 10272 7188
rect 9732 7148 9738 7160
rect 11054 7148 11060 7200
rect 11112 7148 11118 7200
rect 11164 7188 11192 7228
rect 12192 7225 12204 7259
rect 12238 7256 12250 7259
rect 12529 7259 12587 7265
rect 12529 7256 12541 7259
rect 12238 7228 12541 7256
rect 12238 7225 12250 7228
rect 12192 7219 12250 7225
rect 12529 7225 12541 7228
rect 12575 7225 12587 7259
rect 12529 7219 12587 7225
rect 12912 7188 12940 7364
rect 12986 7284 12992 7336
rect 13044 7324 13050 7336
rect 14458 7324 14464 7336
rect 13044 7296 14464 7324
rect 13044 7284 13050 7296
rect 14458 7284 14464 7296
rect 14516 7284 14522 7336
rect 14568 7324 14596 7488
rect 15764 7392 15792 7488
rect 19610 7460 19616 7472
rect 17236 7432 19616 7460
rect 15764 7364 16160 7392
rect 16132 7333 16160 7364
rect 17236 7333 17264 7432
rect 19610 7420 19616 7432
rect 19668 7420 19674 7472
rect 23400 7460 23428 7500
rect 23474 7488 23480 7540
rect 23532 7528 23538 7540
rect 23661 7531 23719 7537
rect 23661 7528 23673 7531
rect 23532 7500 23673 7528
rect 23532 7488 23538 7500
rect 23661 7497 23673 7500
rect 23707 7497 23719 7531
rect 23661 7491 23719 7497
rect 25317 7531 25375 7537
rect 25317 7497 25329 7531
rect 25363 7528 25375 7531
rect 25590 7528 25596 7540
rect 25363 7500 25596 7528
rect 25363 7497 25375 7500
rect 25317 7491 25375 7497
rect 25590 7488 25596 7500
rect 25648 7488 25654 7540
rect 24394 7460 24400 7472
rect 23400 7432 24400 7460
rect 24394 7420 24400 7432
rect 24452 7420 24458 7472
rect 19058 7352 19064 7404
rect 19116 7392 19122 7404
rect 19797 7395 19855 7401
rect 19797 7392 19809 7395
rect 19116 7364 19809 7392
rect 19116 7352 19122 7364
rect 19797 7361 19809 7364
rect 19843 7361 19855 7395
rect 19797 7355 19855 7361
rect 24302 7352 24308 7404
rect 24360 7352 24366 7404
rect 25133 7395 25191 7401
rect 25133 7361 25145 7395
rect 25179 7392 25191 7395
rect 25222 7392 25228 7404
rect 25179 7364 25228 7392
rect 25179 7361 25191 7364
rect 25133 7355 25191 7361
rect 25222 7352 25228 7364
rect 25280 7352 25286 7404
rect 25314 7352 25320 7404
rect 25372 7392 25378 7404
rect 25372 7364 25728 7392
rect 25372 7352 25378 7364
rect 15933 7327 15991 7333
rect 15933 7324 15945 7327
rect 14568 7296 15945 7324
rect 15933 7293 15945 7296
rect 15979 7293 15991 7327
rect 15933 7287 15991 7293
rect 16117 7327 16175 7333
rect 16117 7293 16129 7327
rect 16163 7293 16175 7327
rect 17221 7327 17279 7333
rect 17221 7324 17233 7327
rect 16117 7287 16175 7293
rect 16960 7296 17233 7324
rect 15948 7256 15976 7287
rect 16960 7256 16988 7296
rect 17221 7293 17233 7296
rect 17267 7293 17279 7327
rect 17221 7287 17279 7293
rect 17405 7327 17463 7333
rect 17405 7293 17417 7327
rect 17451 7293 17463 7327
rect 17405 7287 17463 7293
rect 18969 7327 19027 7333
rect 18969 7293 18981 7327
rect 19015 7324 19027 7327
rect 19150 7324 19156 7336
rect 19015 7296 19156 7324
rect 19015 7293 19027 7296
rect 18969 7287 19027 7293
rect 15948 7228 16988 7256
rect 17034 7216 17040 7268
rect 17092 7256 17098 7268
rect 17420 7256 17448 7287
rect 19150 7284 19156 7296
rect 19208 7284 19214 7336
rect 19334 7284 19340 7336
rect 19392 7284 19398 7336
rect 19521 7327 19579 7333
rect 19521 7293 19533 7327
rect 19567 7293 19579 7327
rect 19521 7287 19579 7293
rect 17092 7228 17448 7256
rect 17092 7216 17098 7228
rect 19242 7216 19248 7268
rect 19300 7256 19306 7268
rect 19536 7256 19564 7287
rect 21634 7284 21640 7336
rect 21692 7284 21698 7336
rect 22281 7327 22339 7333
rect 22281 7293 22293 7327
rect 22327 7324 22339 7327
rect 23750 7324 23756 7336
rect 22327 7296 23756 7324
rect 22327 7293 22339 7296
rect 22281 7287 22339 7293
rect 23750 7284 23756 7296
rect 23808 7284 23814 7336
rect 22554 7265 22560 7268
rect 22548 7256 22560 7265
rect 19300 7228 19564 7256
rect 22515 7228 22560 7256
rect 19300 7216 19306 7228
rect 22548 7219 22560 7228
rect 22554 7216 22560 7219
rect 22612 7216 22618 7268
rect 24320 7256 24348 7352
rect 25038 7284 25044 7336
rect 25096 7324 25102 7336
rect 25406 7324 25412 7336
rect 25096 7296 25412 7324
rect 25096 7284 25102 7296
rect 25406 7284 25412 7296
rect 25464 7284 25470 7336
rect 25700 7333 25728 7364
rect 25501 7327 25559 7333
rect 25501 7293 25513 7327
rect 25547 7293 25559 7327
rect 25501 7287 25559 7293
rect 25685 7327 25743 7333
rect 25685 7293 25697 7327
rect 25731 7293 25743 7327
rect 25685 7287 25743 7293
rect 25516 7256 25544 7287
rect 24320 7228 25544 7256
rect 11164 7160 12940 7188
rect 19705 7191 19763 7197
rect 19705 7157 19717 7191
rect 19751 7188 19763 7191
rect 20346 7188 20352 7200
rect 19751 7160 20352 7188
rect 19751 7157 19763 7160
rect 19705 7151 19763 7157
rect 20346 7148 20352 7160
rect 20404 7148 20410 7200
rect 25498 7148 25504 7200
rect 25556 7148 25562 7200
rect 552 7098 27576 7120
rect 552 7046 7114 7098
rect 7166 7046 7178 7098
rect 7230 7046 7242 7098
rect 7294 7046 7306 7098
rect 7358 7046 7370 7098
rect 7422 7046 13830 7098
rect 13882 7046 13894 7098
rect 13946 7046 13958 7098
rect 14010 7046 14022 7098
rect 14074 7046 14086 7098
rect 14138 7046 20546 7098
rect 20598 7046 20610 7098
rect 20662 7046 20674 7098
rect 20726 7046 20738 7098
rect 20790 7046 20802 7098
rect 20854 7046 27262 7098
rect 27314 7046 27326 7098
rect 27378 7046 27390 7098
rect 27442 7046 27454 7098
rect 27506 7046 27518 7098
rect 27570 7046 27576 7098
rect 552 7024 27576 7046
rect 1854 6944 1860 6996
rect 1912 6984 1918 6996
rect 2317 6987 2375 6993
rect 2317 6984 2329 6987
rect 1912 6956 2329 6984
rect 1912 6944 1918 6956
rect 2317 6953 2329 6956
rect 2363 6953 2375 6987
rect 2317 6947 2375 6953
rect 2958 6944 2964 6996
rect 3016 6984 3022 6996
rect 6917 6987 6975 6993
rect 3016 6956 6868 6984
rect 3016 6944 3022 6956
rect 2866 6916 2872 6928
rect 860 6888 2872 6916
rect 860 6857 888 6888
rect 2866 6876 2872 6888
rect 2924 6876 2930 6928
rect 4522 6916 4528 6928
rect 3344 6888 3648 6916
rect 1118 6857 1124 6860
rect 845 6851 903 6857
rect 845 6817 857 6851
rect 891 6817 903 6851
rect 845 6811 903 6817
rect 1112 6811 1124 6857
rect 1118 6808 1124 6811
rect 1176 6808 1182 6860
rect 2498 6808 2504 6860
rect 2556 6848 2562 6860
rect 2777 6851 2835 6857
rect 2777 6848 2789 6851
rect 2556 6820 2789 6848
rect 2556 6808 2562 6820
rect 2777 6817 2789 6820
rect 2823 6817 2835 6851
rect 2777 6811 2835 6817
rect 3145 6851 3203 6857
rect 3145 6817 3157 6851
rect 3191 6817 3203 6851
rect 3145 6811 3203 6817
rect 3237 6851 3295 6857
rect 3237 6817 3249 6851
rect 3283 6848 3295 6851
rect 3344 6848 3372 6888
rect 3620 6860 3648 6888
rect 3988 6888 4528 6916
rect 3283 6820 3372 6848
rect 3421 6851 3479 6857
rect 3283 6817 3295 6820
rect 3237 6811 3295 6817
rect 3421 6817 3433 6851
rect 3467 6848 3479 6851
rect 3467 6820 3556 6848
rect 3467 6817 3479 6820
rect 3421 6811 3479 6817
rect 3160 6780 3188 6811
rect 3528 6789 3556 6820
rect 3602 6808 3608 6860
rect 3660 6848 3666 6860
rect 3988 6857 4016 6888
rect 4522 6876 4528 6888
rect 4580 6876 4586 6928
rect 5350 6916 5356 6928
rect 5408 6925 5414 6928
rect 5320 6888 5356 6916
rect 5350 6876 5356 6888
rect 5408 6879 5420 6925
rect 6840 6916 6868 6956
rect 6917 6953 6929 6987
rect 6963 6984 6975 6987
rect 7006 6984 7012 6996
rect 6963 6956 7012 6984
rect 6963 6953 6975 6956
rect 6917 6947 6975 6953
rect 7006 6944 7012 6956
rect 7064 6944 7070 6996
rect 7466 6944 7472 6996
rect 7524 6944 7530 6996
rect 10042 6944 10048 6996
rect 10100 6944 10106 6996
rect 10318 6944 10324 6996
rect 10376 6984 10382 6996
rect 10413 6987 10471 6993
rect 10413 6984 10425 6987
rect 10376 6956 10425 6984
rect 10376 6944 10382 6956
rect 10413 6953 10425 6956
rect 10459 6953 10471 6987
rect 10413 6947 10471 6953
rect 11882 6944 11888 6996
rect 11940 6944 11946 6996
rect 12158 6944 12164 6996
rect 12216 6984 12222 6996
rect 12437 6987 12495 6993
rect 12437 6984 12449 6987
rect 12216 6956 12449 6984
rect 12216 6944 12222 6956
rect 12437 6953 12449 6956
rect 12483 6953 12495 6987
rect 12437 6947 12495 6953
rect 12798 6987 12856 6993
rect 12798 6953 12810 6987
rect 12844 6984 12856 6987
rect 12844 6956 13288 6984
rect 12844 6953 12856 6956
rect 12798 6947 12856 6953
rect 10060 6916 10088 6944
rect 10502 6916 10508 6928
rect 6840 6888 10508 6916
rect 5408 6876 5414 6879
rect 10502 6876 10508 6888
rect 10560 6876 10566 6928
rect 11054 6876 11060 6928
rect 11112 6916 11118 6928
rect 11112 6888 11560 6916
rect 11112 6876 11118 6888
rect 3789 6851 3847 6857
rect 3789 6848 3801 6851
rect 3660 6820 3801 6848
rect 3660 6808 3666 6820
rect 3789 6817 3801 6820
rect 3835 6817 3847 6851
rect 3789 6811 3847 6817
rect 3881 6851 3939 6857
rect 3881 6817 3893 6851
rect 3927 6817 3939 6851
rect 3881 6811 3939 6817
rect 3973 6851 4031 6857
rect 3973 6817 3985 6851
rect 4019 6817 4031 6851
rect 3973 6811 4031 6817
rect 4157 6851 4215 6857
rect 4157 6817 4169 6851
rect 4203 6848 4215 6851
rect 4614 6848 4620 6860
rect 4203 6820 4620 6848
rect 4203 6817 4215 6820
rect 4157 6811 4215 6817
rect 3513 6783 3571 6789
rect 3160 6752 3280 6780
rect 2148 6684 2544 6712
rect 2148 6656 2176 6684
rect 2130 6604 2136 6656
rect 2188 6604 2194 6656
rect 2222 6604 2228 6656
rect 2280 6604 2286 6656
rect 2516 6653 2544 6684
rect 2501 6647 2559 6653
rect 2501 6613 2513 6647
rect 2547 6613 2559 6647
rect 3252 6644 3280 6752
rect 3513 6749 3525 6783
rect 3559 6749 3571 6783
rect 3513 6743 3571 6749
rect 3694 6740 3700 6792
rect 3752 6740 3758 6792
rect 3896 6780 3924 6811
rect 4614 6808 4620 6820
rect 4672 6808 4678 6860
rect 5629 6851 5687 6857
rect 5629 6817 5641 6851
rect 5675 6848 5687 6851
rect 6086 6848 6092 6860
rect 5675 6820 6092 6848
rect 5675 6817 5687 6820
rect 5629 6811 5687 6817
rect 6086 6808 6092 6820
rect 6144 6808 6150 6860
rect 6178 6808 6184 6860
rect 6236 6808 6242 6860
rect 6365 6851 6423 6857
rect 6365 6817 6377 6851
rect 6411 6848 6423 6851
rect 6638 6848 6644 6860
rect 6411 6820 6644 6848
rect 6411 6817 6423 6820
rect 6365 6811 6423 6817
rect 6638 6808 6644 6820
rect 6696 6808 6702 6860
rect 6914 6808 6920 6860
rect 6972 6848 6978 6860
rect 7009 6851 7067 6857
rect 7009 6848 7021 6851
rect 6972 6820 7021 6848
rect 6972 6808 6978 6820
rect 7009 6817 7021 6820
rect 7055 6817 7067 6851
rect 7009 6811 7067 6817
rect 7285 6851 7343 6857
rect 7285 6817 7297 6851
rect 7331 6817 7343 6851
rect 7285 6811 7343 6817
rect 7653 6851 7711 6857
rect 7653 6817 7665 6851
rect 7699 6848 7711 6851
rect 8478 6848 8484 6860
rect 7699 6820 8484 6848
rect 7699 6817 7711 6820
rect 7653 6811 7711 6817
rect 6273 6783 6331 6789
rect 3896 6752 4292 6780
rect 3421 6715 3479 6721
rect 3421 6681 3433 6715
rect 3467 6712 3479 6715
rect 3712 6712 3740 6740
rect 3467 6684 3740 6712
rect 3467 6681 3479 6684
rect 3421 6675 3479 6681
rect 3896 6644 3924 6752
rect 4264 6724 4292 6752
rect 6273 6749 6285 6783
rect 6319 6780 6331 6783
rect 6457 6783 6515 6789
rect 6457 6780 6469 6783
rect 6319 6752 6469 6780
rect 6319 6749 6331 6752
rect 6273 6743 6331 6749
rect 6457 6749 6469 6752
rect 6503 6780 6515 6783
rect 7101 6783 7159 6789
rect 7101 6780 7113 6783
rect 6503 6752 7113 6780
rect 6503 6749 6515 6752
rect 6457 6743 6515 6749
rect 7101 6749 7113 6752
rect 7147 6749 7159 6783
rect 7101 6743 7159 6749
rect 4246 6672 4252 6724
rect 4304 6672 4310 6724
rect 6733 6715 6791 6721
rect 6733 6712 6745 6715
rect 6656 6684 6745 6712
rect 6656 6656 6684 6684
rect 6733 6681 6745 6684
rect 6779 6712 6791 6715
rect 7300 6712 7328 6811
rect 8478 6808 8484 6820
rect 8536 6808 8542 6860
rect 8570 6808 8576 6860
rect 8628 6848 8634 6860
rect 9042 6851 9100 6857
rect 9042 6848 9054 6851
rect 8628 6820 9054 6848
rect 8628 6808 8634 6820
rect 9042 6817 9054 6820
rect 9088 6817 9100 6851
rect 9042 6811 9100 6817
rect 9214 6808 9220 6860
rect 9272 6848 9278 6860
rect 9309 6851 9367 6857
rect 9309 6848 9321 6851
rect 9272 6820 9321 6848
rect 9272 6808 9278 6820
rect 9309 6817 9321 6820
rect 9355 6817 9367 6851
rect 9953 6851 10011 6857
rect 9953 6848 9965 6851
rect 9309 6811 9367 6817
rect 9692 6820 9965 6848
rect 9692 6792 9720 6820
rect 9953 6817 9965 6820
rect 9999 6817 10011 6851
rect 9953 6811 10011 6817
rect 10045 6851 10103 6857
rect 10045 6817 10057 6851
rect 10091 6848 10103 6851
rect 10134 6848 10140 6860
rect 10091 6820 10140 6848
rect 10091 6817 10103 6820
rect 10045 6811 10103 6817
rect 10134 6808 10140 6820
rect 10192 6808 10198 6860
rect 10226 6808 10232 6860
rect 10284 6808 10290 6860
rect 11532 6857 11560 6888
rect 11333 6851 11391 6857
rect 11333 6817 11345 6851
rect 11379 6817 11391 6851
rect 11333 6811 11391 6817
rect 11517 6851 11575 6857
rect 11517 6817 11529 6851
rect 11563 6848 11575 6851
rect 11790 6848 11796 6860
rect 11563 6820 11796 6848
rect 11563 6817 11575 6820
rect 11517 6811 11575 6817
rect 9674 6740 9680 6792
rect 9732 6740 9738 6792
rect 6779 6684 7328 6712
rect 7837 6715 7895 6721
rect 6779 6681 6791 6684
rect 6733 6675 6791 6681
rect 7837 6681 7849 6715
rect 7883 6712 7895 6715
rect 7883 6684 8432 6712
rect 7883 6681 7895 6684
rect 7837 6675 7895 6681
rect 3252 6616 3924 6644
rect 2501 6607 2559 6613
rect 6638 6604 6644 6656
rect 6696 6604 6702 6656
rect 7926 6604 7932 6656
rect 7984 6604 7990 6656
rect 8404 6644 8432 6684
rect 8570 6644 8576 6656
rect 8404 6616 8576 6644
rect 8570 6604 8576 6616
rect 8628 6604 8634 6656
rect 10244 6644 10272 6808
rect 11238 6740 11244 6792
rect 11296 6780 11302 6792
rect 11348 6780 11376 6811
rect 11790 6808 11796 6820
rect 11848 6808 11854 6860
rect 11900 6857 11928 6944
rect 12894 6876 12900 6928
rect 12952 6876 12958 6928
rect 11885 6851 11943 6857
rect 11885 6817 11897 6851
rect 11931 6817 11943 6851
rect 11885 6811 11943 6817
rect 11977 6851 12035 6857
rect 11977 6817 11989 6851
rect 12023 6817 12035 6851
rect 11977 6811 12035 6817
rect 11296 6752 11376 6780
rect 11425 6783 11483 6789
rect 11296 6740 11302 6752
rect 11425 6749 11437 6783
rect 11471 6780 11483 6783
rect 11609 6783 11667 6789
rect 11609 6780 11621 6783
rect 11471 6752 11621 6780
rect 11471 6749 11483 6752
rect 11425 6743 11483 6749
rect 11609 6749 11621 6752
rect 11655 6780 11667 6783
rect 11992 6780 12020 6811
rect 12526 6808 12532 6860
rect 12584 6848 12590 6860
rect 12621 6851 12679 6857
rect 12621 6848 12633 6851
rect 12584 6820 12633 6848
rect 12584 6808 12590 6820
rect 12621 6817 12633 6820
rect 12667 6817 12679 6851
rect 12621 6811 12679 6817
rect 12710 6808 12716 6860
rect 12768 6808 12774 6860
rect 13260 6857 13288 6956
rect 14458 6944 14464 6996
rect 14516 6944 14522 6996
rect 15105 6987 15163 6993
rect 15105 6953 15117 6987
rect 15151 6984 15163 6987
rect 15378 6984 15384 6996
rect 15151 6956 15384 6984
rect 15151 6953 15163 6956
rect 15105 6947 15163 6953
rect 15378 6944 15384 6956
rect 15436 6944 15442 6996
rect 22738 6944 22744 6996
rect 22796 6944 22802 6996
rect 14844 6888 15056 6916
rect 12989 6851 13047 6857
rect 12989 6846 13001 6851
rect 12820 6818 13001 6846
rect 12820 6780 12848 6818
rect 12989 6817 13001 6818
rect 13035 6817 13047 6851
rect 12989 6811 13047 6817
rect 13245 6851 13303 6857
rect 13245 6817 13257 6851
rect 13291 6817 13303 6851
rect 14645 6851 14703 6857
rect 14645 6848 14657 6851
rect 13245 6811 13303 6817
rect 14568 6820 14657 6848
rect 14568 6780 14596 6820
rect 14645 6817 14657 6820
rect 14691 6848 14703 6851
rect 14844 6848 14872 6888
rect 14691 6820 14872 6848
rect 14921 6851 14979 6857
rect 14691 6817 14703 6820
rect 14645 6811 14703 6817
rect 14921 6817 14933 6851
rect 14967 6817 14979 6851
rect 15028 6848 15056 6888
rect 16850 6876 16856 6928
rect 16908 6876 16914 6928
rect 19886 6876 19892 6928
rect 19944 6916 19950 6928
rect 20438 6916 20444 6928
rect 19944 6888 20444 6916
rect 19944 6876 19950 6888
rect 20438 6876 20444 6888
rect 20496 6916 20502 6928
rect 22756 6916 22784 6944
rect 20496 6888 20760 6916
rect 20496 6876 20502 6888
rect 15378 6848 15384 6860
rect 15028 6820 15384 6848
rect 14921 6811 14979 6817
rect 14936 6780 14964 6811
rect 15378 6808 15384 6820
rect 15436 6808 15442 6860
rect 16574 6808 16580 6860
rect 16632 6808 16638 6860
rect 16761 6851 16819 6857
rect 16761 6817 16773 6851
rect 16807 6848 16819 6851
rect 16868 6848 16896 6876
rect 16807 6820 16896 6848
rect 16807 6817 16819 6820
rect 16761 6811 16819 6817
rect 18046 6808 18052 6860
rect 18104 6848 18110 6860
rect 18877 6851 18935 6857
rect 18877 6848 18889 6851
rect 18104 6820 18889 6848
rect 18104 6808 18110 6820
rect 18877 6817 18889 6820
rect 18923 6817 18935 6851
rect 18877 6811 18935 6817
rect 19058 6808 19064 6860
rect 19116 6808 19122 6860
rect 19245 6851 19303 6857
rect 19245 6817 19257 6851
rect 19291 6848 19303 6851
rect 19337 6851 19395 6857
rect 19337 6848 19349 6851
rect 19291 6820 19349 6848
rect 19291 6817 19303 6820
rect 19245 6811 19303 6817
rect 19337 6817 19349 6820
rect 19383 6817 19395 6851
rect 19337 6811 19395 6817
rect 19518 6808 19524 6860
rect 19576 6848 19582 6860
rect 19794 6848 19800 6860
rect 19576 6820 19800 6848
rect 19576 6808 19582 6820
rect 19794 6808 19800 6820
rect 19852 6848 19858 6860
rect 20732 6857 20760 6888
rect 21376 6888 21772 6916
rect 22756 6888 23980 6916
rect 21376 6857 21404 6888
rect 20625 6851 20683 6857
rect 20625 6848 20637 6851
rect 19852 6820 20637 6848
rect 19852 6808 19858 6820
rect 20625 6817 20637 6820
rect 20671 6817 20683 6851
rect 20625 6811 20683 6817
rect 20717 6851 20775 6857
rect 20717 6817 20729 6851
rect 20763 6817 20775 6851
rect 20717 6811 20775 6817
rect 20901 6851 20959 6857
rect 20901 6817 20913 6851
rect 20947 6817 20959 6851
rect 20901 6811 20959 6817
rect 21085 6851 21143 6857
rect 21085 6817 21097 6851
rect 21131 6848 21143 6851
rect 21269 6851 21327 6857
rect 21269 6848 21281 6851
rect 21131 6820 21281 6848
rect 21131 6817 21143 6820
rect 21085 6811 21143 6817
rect 21269 6817 21281 6820
rect 21315 6817 21327 6851
rect 21269 6811 21327 6817
rect 21361 6851 21419 6857
rect 21361 6817 21373 6851
rect 21407 6817 21419 6851
rect 21361 6811 21419 6817
rect 21453 6851 21511 6857
rect 21453 6817 21465 6851
rect 21499 6817 21511 6851
rect 21453 6811 21511 6817
rect 11655 6752 12020 6780
rect 12452 6752 12848 6780
rect 14292 6752 14596 6780
rect 14660 6752 14964 6780
rect 11655 6749 11667 6752
rect 11609 6743 11667 6749
rect 12452 6724 12480 6752
rect 10318 6672 10324 6724
rect 10376 6712 10382 6724
rect 12434 6712 12440 6724
rect 10376 6684 12440 6712
rect 10376 6672 10382 6684
rect 12434 6672 12440 6684
rect 12492 6672 12498 6724
rect 12710 6672 12716 6724
rect 12768 6672 12774 6724
rect 11698 6644 11704 6656
rect 10244 6616 11704 6644
rect 11698 6604 11704 6616
rect 11756 6604 11762 6656
rect 11793 6647 11851 6653
rect 11793 6613 11805 6647
rect 11839 6644 11851 6647
rect 12066 6644 12072 6656
rect 11839 6616 12072 6644
rect 11839 6613 11851 6616
rect 11793 6607 11851 6613
rect 12066 6604 12072 6616
rect 12124 6604 12130 6656
rect 12728 6644 12756 6672
rect 14292 6644 14320 6752
rect 14660 6656 14688 6752
rect 15102 6740 15108 6792
rect 15160 6740 15166 6792
rect 17954 6740 17960 6792
rect 18012 6740 18018 6792
rect 20916 6780 20944 6811
rect 20916 6752 21128 6780
rect 21100 6724 21128 6752
rect 21174 6740 21180 6792
rect 21232 6780 21238 6792
rect 21468 6780 21496 6811
rect 21634 6808 21640 6860
rect 21692 6808 21698 6860
rect 21744 6848 21772 6888
rect 23952 6857 23980 6888
rect 25516 6888 25912 6916
rect 21913 6851 21971 6857
rect 21913 6848 21925 6851
rect 21744 6820 21925 6848
rect 21913 6817 21925 6820
rect 21959 6817 21971 6851
rect 21913 6811 21971 6817
rect 23937 6851 23995 6857
rect 23937 6817 23949 6851
rect 23983 6817 23995 6851
rect 23937 6811 23995 6817
rect 24121 6851 24179 6857
rect 24121 6817 24133 6851
rect 24167 6817 24179 6851
rect 24121 6811 24179 6817
rect 24305 6851 24363 6857
rect 24305 6817 24317 6851
rect 24351 6848 24363 6851
rect 24397 6851 24455 6857
rect 24397 6848 24409 6851
rect 24351 6820 24409 6848
rect 24351 6817 24363 6820
rect 24305 6811 24363 6817
rect 24397 6817 24409 6820
rect 24443 6817 24455 6851
rect 24397 6811 24455 6817
rect 21542 6780 21548 6792
rect 21232 6752 21548 6780
rect 21232 6740 21238 6752
rect 21542 6740 21548 6752
rect 21600 6740 21606 6792
rect 24136 6780 24164 6811
rect 25038 6808 25044 6860
rect 25096 6848 25102 6860
rect 25516 6857 25544 6888
rect 25501 6851 25559 6857
rect 25501 6848 25513 6851
rect 25096 6820 25513 6848
rect 25096 6808 25102 6820
rect 25501 6817 25513 6820
rect 25547 6817 25559 6851
rect 25685 6851 25743 6857
rect 25685 6848 25697 6851
rect 25501 6811 25559 6817
rect 25608 6820 25697 6848
rect 24946 6780 24952 6792
rect 24136 6752 24952 6780
rect 24946 6740 24952 6752
rect 25004 6740 25010 6792
rect 14737 6715 14795 6721
rect 14737 6681 14749 6715
rect 14783 6681 14795 6715
rect 14737 6675 14795 6681
rect 14829 6715 14887 6721
rect 14829 6681 14841 6715
rect 14875 6712 14887 6715
rect 15194 6712 15200 6724
rect 14875 6684 15200 6712
rect 14875 6681 14887 6684
rect 14829 6675 14887 6681
rect 12728 6616 14320 6644
rect 14366 6604 14372 6656
rect 14424 6604 14430 6656
rect 14642 6604 14648 6656
rect 14700 6604 14706 6656
rect 14752 6644 14780 6675
rect 15194 6672 15200 6684
rect 15252 6672 15258 6724
rect 18322 6672 18328 6724
rect 18380 6672 18386 6724
rect 21082 6672 21088 6724
rect 21140 6672 21146 6724
rect 22649 6715 22707 6721
rect 22649 6681 22661 6715
rect 22695 6712 22707 6715
rect 23106 6712 23112 6724
rect 22695 6684 23112 6712
rect 22695 6681 22707 6684
rect 22649 6675 22707 6681
rect 23106 6672 23112 6684
rect 23164 6672 23170 6724
rect 25608 6656 25636 6820
rect 25685 6817 25697 6820
rect 25731 6848 25743 6851
rect 25777 6851 25835 6857
rect 25777 6848 25789 6851
rect 25731 6820 25789 6848
rect 25731 6817 25743 6820
rect 25685 6811 25743 6817
rect 25777 6817 25789 6820
rect 25823 6817 25835 6851
rect 25884 6848 25912 6888
rect 25961 6851 26019 6857
rect 25961 6848 25973 6851
rect 25884 6820 25973 6848
rect 25777 6811 25835 6817
rect 25961 6817 25973 6820
rect 26007 6817 26019 6851
rect 25961 6811 26019 6817
rect 15286 6644 15292 6656
rect 14752 6616 15292 6644
rect 15286 6604 15292 6616
rect 15344 6604 15350 6656
rect 16666 6604 16672 6656
rect 16724 6604 16730 6656
rect 18414 6604 18420 6656
rect 18472 6604 18478 6656
rect 19518 6604 19524 6656
rect 19576 6604 19582 6656
rect 19978 6604 19984 6656
rect 20036 6604 20042 6656
rect 24486 6604 24492 6656
rect 24544 6644 24550 6656
rect 24581 6647 24639 6653
rect 24581 6644 24593 6647
rect 24544 6616 24593 6644
rect 24544 6604 24550 6616
rect 24581 6613 24593 6616
rect 24627 6613 24639 6647
rect 24581 6607 24639 6613
rect 25590 6604 25596 6656
rect 25648 6604 25654 6656
rect 25682 6604 25688 6656
rect 25740 6604 25746 6656
rect 25774 6604 25780 6656
rect 25832 6644 25838 6656
rect 25869 6647 25927 6653
rect 25869 6644 25881 6647
rect 25832 6616 25881 6644
rect 25832 6604 25838 6616
rect 25869 6613 25881 6616
rect 25915 6613 25927 6647
rect 25869 6607 25927 6613
rect 552 6554 27416 6576
rect 552 6502 3756 6554
rect 3808 6502 3820 6554
rect 3872 6502 3884 6554
rect 3936 6502 3948 6554
rect 4000 6502 4012 6554
rect 4064 6502 10472 6554
rect 10524 6502 10536 6554
rect 10588 6502 10600 6554
rect 10652 6502 10664 6554
rect 10716 6502 10728 6554
rect 10780 6502 17188 6554
rect 17240 6502 17252 6554
rect 17304 6502 17316 6554
rect 17368 6502 17380 6554
rect 17432 6502 17444 6554
rect 17496 6502 23904 6554
rect 23956 6502 23968 6554
rect 24020 6502 24032 6554
rect 24084 6502 24096 6554
rect 24148 6502 24160 6554
rect 24212 6502 27416 6554
rect 552 6480 27416 6502
rect 1118 6400 1124 6452
rect 1176 6440 1182 6452
rect 1397 6443 1455 6449
rect 1397 6440 1409 6443
rect 1176 6412 1409 6440
rect 1176 6400 1182 6412
rect 1397 6409 1409 6412
rect 1443 6409 1455 6443
rect 1397 6403 1455 6409
rect 1765 6443 1823 6449
rect 1765 6409 1777 6443
rect 1811 6440 1823 6443
rect 1854 6440 1860 6452
rect 1811 6412 1860 6440
rect 1811 6409 1823 6412
rect 1765 6403 1823 6409
rect 1854 6400 1860 6412
rect 1912 6400 1918 6452
rect 2130 6400 2136 6452
rect 2188 6400 2194 6452
rect 2222 6400 2228 6452
rect 2280 6400 2286 6452
rect 2317 6443 2375 6449
rect 2317 6409 2329 6443
rect 2363 6440 2375 6443
rect 2498 6440 2504 6452
rect 2363 6412 2504 6440
rect 2363 6409 2375 6412
rect 2317 6403 2375 6409
rect 2498 6400 2504 6412
rect 2556 6400 2562 6452
rect 3602 6400 3608 6452
rect 3660 6400 3666 6452
rect 4246 6400 4252 6452
rect 4304 6400 4310 6452
rect 6178 6400 6184 6452
rect 6236 6400 6242 6452
rect 6638 6400 6644 6452
rect 6696 6400 6702 6452
rect 6914 6400 6920 6452
rect 6972 6440 6978 6452
rect 7193 6443 7251 6449
rect 7193 6440 7205 6443
rect 6972 6412 7205 6440
rect 6972 6400 6978 6412
rect 7193 6409 7205 6412
rect 7239 6409 7251 6443
rect 7193 6403 7251 6409
rect 8662 6400 8668 6452
rect 8720 6440 8726 6452
rect 8849 6443 8907 6449
rect 8849 6440 8861 6443
rect 8720 6412 8861 6440
rect 8720 6400 8726 6412
rect 8849 6409 8861 6412
rect 8895 6409 8907 6443
rect 8849 6403 8907 6409
rect 9214 6400 9220 6452
rect 9272 6440 9278 6452
rect 10318 6440 10324 6452
rect 9272 6412 10324 6440
rect 9272 6400 9278 6412
rect 10318 6400 10324 6412
rect 10376 6400 10382 6452
rect 11698 6400 11704 6452
rect 11756 6400 11762 6452
rect 12066 6400 12072 6452
rect 12124 6440 12130 6452
rect 12345 6443 12403 6449
rect 12345 6440 12357 6443
rect 12124 6412 12357 6440
rect 12124 6400 12130 6412
rect 12345 6409 12357 6412
rect 12391 6409 12403 6443
rect 12345 6403 12403 6409
rect 12894 6400 12900 6452
rect 12952 6440 12958 6452
rect 13633 6443 13691 6449
rect 13633 6440 13645 6443
rect 12952 6412 13645 6440
rect 12952 6400 12958 6412
rect 13633 6409 13645 6412
rect 13679 6409 13691 6443
rect 13633 6403 13691 6409
rect 14090 6400 14096 6452
rect 14148 6440 14154 6452
rect 14185 6443 14243 6449
rect 14185 6440 14197 6443
rect 14148 6412 14197 6440
rect 14148 6400 14154 6412
rect 14185 6409 14197 6412
rect 14231 6409 14243 6443
rect 14185 6403 14243 6409
rect 14366 6400 14372 6452
rect 14424 6400 14430 6452
rect 14642 6400 14648 6452
rect 14700 6400 14706 6452
rect 15010 6400 15016 6452
rect 15068 6400 15074 6452
rect 15378 6400 15384 6452
rect 15436 6440 15442 6452
rect 16025 6443 16083 6449
rect 16025 6440 16037 6443
rect 15436 6412 16037 6440
rect 15436 6400 15442 6412
rect 16025 6409 16037 6412
rect 16071 6409 16083 6443
rect 16025 6403 16083 6409
rect 17034 6400 17040 6452
rect 17092 6400 17098 6452
rect 18414 6400 18420 6452
rect 18472 6400 18478 6452
rect 19058 6400 19064 6452
rect 19116 6400 19122 6452
rect 19978 6400 19984 6452
rect 20036 6440 20042 6452
rect 20036 6412 20392 6440
rect 20036 6400 20042 6412
rect 1762 6264 1768 6316
rect 1820 6304 1826 6316
rect 1857 6307 1915 6313
rect 1857 6304 1869 6307
rect 1820 6276 1869 6304
rect 1820 6264 1826 6276
rect 1857 6273 1869 6276
rect 1903 6273 1915 6307
rect 1857 6267 1915 6273
rect 1581 6239 1639 6245
rect 1581 6205 1593 6239
rect 1627 6236 1639 6239
rect 1670 6236 1676 6248
rect 1627 6208 1676 6236
rect 1627 6205 1639 6208
rect 1581 6199 1639 6205
rect 1670 6196 1676 6208
rect 1728 6196 1734 6248
rect 2240 6245 2268 6400
rect 1949 6239 2007 6245
rect 1949 6205 1961 6239
rect 1995 6205 2007 6239
rect 1949 6199 2007 6205
rect 2133 6239 2191 6245
rect 2133 6205 2145 6239
rect 2179 6236 2191 6239
rect 2225 6239 2283 6245
rect 2225 6236 2237 6239
rect 2179 6208 2237 6236
rect 2179 6205 2191 6208
rect 2133 6199 2191 6205
rect 2225 6205 2237 6208
rect 2271 6205 2283 6239
rect 2225 6199 2283 6205
rect 2409 6239 2467 6245
rect 2409 6205 2421 6239
rect 2455 6205 2467 6239
rect 2409 6199 2467 6205
rect 1964 6168 1992 6199
rect 2424 6168 2452 6199
rect 2682 6196 2688 6248
rect 2740 6196 2746 6248
rect 3510 6196 3516 6248
rect 3568 6196 3574 6248
rect 3620 6245 3648 6400
rect 3697 6307 3755 6313
rect 3697 6273 3709 6307
rect 3743 6304 3755 6307
rect 4264 6304 4292 6400
rect 3743 6276 4292 6304
rect 6196 6304 6224 6400
rect 8110 6372 8116 6384
rect 7484 6344 8116 6372
rect 6196 6276 6776 6304
rect 3743 6273 3755 6276
rect 3697 6267 3755 6273
rect 6748 6248 6776 6276
rect 3605 6239 3663 6245
rect 3605 6205 3617 6239
rect 3651 6205 3663 6239
rect 3605 6199 3663 6205
rect 4798 6196 4804 6248
rect 4856 6196 4862 6248
rect 5810 6196 5816 6248
rect 5868 6196 5874 6248
rect 6546 6196 6552 6248
rect 6604 6196 6610 6248
rect 6730 6196 6736 6248
rect 6788 6196 6794 6248
rect 7377 6239 7435 6245
rect 7377 6205 7389 6239
rect 7423 6236 7435 6239
rect 7484 6236 7512 6344
rect 8110 6332 8116 6344
rect 8168 6332 8174 6384
rect 8294 6332 8300 6384
rect 8352 6372 8358 6384
rect 14384 6372 14412 6400
rect 8352 6344 12480 6372
rect 8352 6332 8358 6344
rect 7561 6307 7619 6313
rect 7561 6273 7573 6307
rect 7607 6304 7619 6307
rect 7742 6304 7748 6316
rect 7607 6276 7748 6304
rect 7607 6273 7619 6276
rect 7561 6267 7619 6273
rect 7742 6264 7748 6276
rect 7800 6264 7806 6316
rect 8205 6307 8263 6313
rect 8205 6273 8217 6307
rect 8251 6304 8263 6307
rect 8481 6307 8539 6313
rect 8481 6304 8493 6307
rect 8251 6276 8493 6304
rect 8251 6273 8263 6276
rect 8205 6267 8263 6273
rect 8481 6273 8493 6276
rect 8527 6273 8539 6307
rect 8481 6267 8539 6273
rect 11256 6276 12204 6304
rect 11256 6248 11284 6276
rect 7423 6208 7512 6236
rect 7653 6239 7711 6245
rect 7423 6205 7435 6208
rect 7377 6199 7435 6205
rect 7653 6205 7665 6239
rect 7699 6236 7711 6239
rect 8573 6239 8631 6245
rect 8573 6236 8585 6239
rect 7699 6208 8585 6236
rect 7699 6205 7711 6208
rect 7653 6199 7711 6205
rect 1964 6140 2452 6168
rect 2240 6112 2268 6140
rect 2222 6060 2228 6112
rect 2280 6060 2286 6112
rect 3528 6100 3556 6196
rect 8220 6112 8248 6208
rect 8573 6205 8585 6208
rect 8619 6205 8631 6239
rect 8573 6199 8631 6205
rect 11238 6196 11244 6248
rect 11296 6196 11302 6248
rect 11514 6196 11520 6248
rect 11572 6196 11578 6248
rect 11609 6239 11667 6245
rect 11609 6205 11621 6239
rect 11655 6205 11667 6239
rect 11609 6199 11667 6205
rect 11624 6168 11652 6199
rect 11790 6196 11796 6248
rect 11848 6196 11854 6248
rect 11882 6196 11888 6248
rect 11940 6196 11946 6248
rect 12176 6245 12204 6276
rect 12161 6239 12219 6245
rect 12161 6205 12173 6239
rect 12207 6205 12219 6239
rect 12161 6199 12219 6205
rect 12345 6239 12403 6245
rect 12345 6205 12357 6239
rect 12391 6205 12403 6239
rect 12345 6199 12403 6205
rect 11532 6140 11652 6168
rect 11808 6168 11836 6196
rect 12360 6168 12388 6199
rect 11808 6140 12388 6168
rect 11532 6112 11560 6140
rect 3973 6103 4031 6109
rect 3973 6100 3985 6103
rect 3528 6072 3985 6100
rect 3973 6069 3985 6072
rect 4019 6069 4031 6103
rect 3973 6063 4031 6069
rect 8202 6060 8208 6112
rect 8260 6060 8266 6112
rect 10229 6103 10287 6109
rect 10229 6069 10241 6103
rect 10275 6100 10287 6103
rect 10318 6100 10324 6112
rect 10275 6072 10324 6100
rect 10275 6069 10287 6072
rect 10229 6063 10287 6069
rect 10318 6060 10324 6072
rect 10376 6060 10382 6112
rect 11514 6060 11520 6112
rect 11572 6060 11578 6112
rect 11606 6060 11612 6112
rect 11664 6100 11670 6112
rect 12069 6103 12127 6109
rect 12069 6100 12081 6103
rect 11664 6072 12081 6100
rect 11664 6060 11670 6072
rect 12069 6069 12081 6072
rect 12115 6069 12127 6103
rect 12452 6100 12480 6344
rect 14108 6344 14412 6372
rect 12526 6264 12532 6316
rect 12584 6264 12590 6316
rect 12618 6264 12624 6316
rect 12676 6304 12682 6316
rect 13541 6307 13599 6313
rect 13541 6304 13553 6307
rect 12676 6276 13553 6304
rect 12676 6264 12682 6276
rect 13541 6273 13553 6276
rect 13587 6273 13599 6307
rect 13541 6267 13599 6273
rect 12544 6236 12572 6264
rect 13722 6236 13728 6248
rect 12544 6208 13728 6236
rect 13722 6196 13728 6208
rect 13780 6196 13786 6248
rect 14108 6245 14136 6344
rect 15028 6304 15056 6400
rect 15194 6332 15200 6384
rect 15252 6372 15258 6384
rect 16666 6372 16672 6384
rect 15252 6344 15516 6372
rect 15252 6332 15258 6344
rect 14384 6276 15148 6304
rect 14384 6245 14412 6276
rect 13817 6239 13875 6245
rect 13817 6205 13829 6239
rect 13863 6205 13875 6239
rect 13817 6199 13875 6205
rect 14093 6239 14151 6245
rect 14093 6205 14105 6239
rect 14139 6205 14151 6239
rect 14093 6199 14151 6205
rect 14277 6239 14335 6245
rect 14277 6205 14289 6239
rect 14323 6205 14335 6239
rect 14277 6199 14335 6205
rect 14369 6239 14427 6245
rect 14369 6205 14381 6239
rect 14415 6205 14427 6239
rect 14369 6199 14427 6205
rect 12710 6128 12716 6180
rect 12768 6168 12774 6180
rect 13832 6168 13860 6199
rect 12768 6140 13860 6168
rect 14292 6168 14320 6199
rect 15010 6196 15016 6248
rect 15068 6196 15074 6248
rect 15120 6245 15148 6276
rect 15488 6245 15516 6344
rect 16224 6344 16672 6372
rect 16224 6245 16252 6344
rect 16666 6332 16672 6344
rect 16724 6372 16730 6384
rect 17313 6375 17371 6381
rect 17313 6372 17325 6375
rect 16724 6344 17325 6372
rect 16724 6332 16730 6344
rect 17313 6341 17325 6344
rect 17359 6341 17371 6375
rect 17313 6335 17371 6341
rect 16853 6307 16911 6313
rect 16853 6273 16865 6307
rect 16899 6304 16911 6307
rect 17221 6307 17279 6313
rect 17221 6304 17233 6307
rect 16899 6276 17233 6304
rect 16899 6273 16911 6276
rect 16853 6267 16911 6273
rect 17221 6273 17233 6276
rect 17267 6273 17279 6307
rect 17221 6267 17279 6273
rect 18233 6307 18291 6313
rect 18233 6273 18245 6307
rect 18279 6304 18291 6307
rect 18432 6304 18460 6400
rect 18509 6375 18567 6381
rect 18509 6341 18521 6375
rect 18555 6372 18567 6375
rect 19076 6372 19104 6400
rect 18555 6344 19104 6372
rect 18555 6341 18567 6344
rect 18509 6335 18567 6341
rect 20364 6313 20392 6412
rect 20990 6400 20996 6452
rect 21048 6440 21054 6452
rect 21361 6443 21419 6449
rect 21361 6440 21373 6443
rect 21048 6412 21373 6440
rect 21048 6400 21054 6412
rect 21361 6409 21373 6412
rect 21407 6409 21419 6443
rect 21361 6403 21419 6409
rect 22462 6400 22468 6452
rect 22520 6400 22526 6452
rect 23566 6400 23572 6452
rect 23624 6400 23630 6452
rect 24946 6400 24952 6452
rect 25004 6440 25010 6452
rect 25004 6412 25176 6440
rect 25004 6400 25010 6412
rect 25148 6372 25176 6412
rect 25590 6400 25596 6452
rect 25648 6400 25654 6452
rect 25961 6443 26019 6449
rect 25961 6440 25973 6443
rect 25700 6412 25973 6440
rect 25700 6372 25728 6412
rect 25961 6409 25973 6412
rect 26007 6409 26019 6443
rect 25961 6403 26019 6409
rect 25148 6344 25728 6372
rect 25774 6332 25780 6384
rect 25832 6372 25838 6384
rect 26605 6375 26663 6381
rect 26605 6372 26617 6375
rect 25832 6344 26617 6372
rect 25832 6332 25838 6344
rect 26605 6341 26617 6344
rect 26651 6341 26663 6375
rect 26605 6335 26663 6341
rect 18279 6276 18460 6304
rect 20349 6307 20407 6313
rect 18279 6273 18291 6276
rect 18233 6267 18291 6273
rect 20349 6273 20361 6307
rect 20395 6273 20407 6307
rect 20349 6267 20407 6273
rect 23750 6264 23756 6316
rect 23808 6304 23814 6316
rect 24213 6307 24271 6313
rect 24213 6304 24225 6307
rect 23808 6276 24225 6304
rect 23808 6264 23814 6276
rect 24213 6273 24225 6276
rect 24259 6273 24271 6307
rect 24213 6267 24271 6273
rect 26329 6307 26387 6313
rect 26329 6273 26341 6307
rect 26375 6304 26387 6307
rect 26513 6307 26571 6313
rect 26513 6304 26525 6307
rect 26375 6276 26525 6304
rect 26375 6273 26387 6276
rect 26329 6267 26387 6273
rect 26513 6273 26525 6276
rect 26559 6273 26571 6307
rect 26513 6267 26571 6273
rect 15105 6239 15163 6245
rect 15105 6205 15117 6239
rect 15151 6205 15163 6239
rect 15105 6199 15163 6205
rect 15197 6239 15255 6245
rect 15197 6205 15209 6239
rect 15243 6205 15255 6239
rect 15197 6199 15255 6205
rect 15381 6239 15439 6245
rect 15381 6205 15393 6239
rect 15427 6236 15439 6239
rect 15473 6239 15531 6245
rect 15473 6236 15485 6239
rect 15427 6208 15485 6236
rect 15427 6205 15439 6208
rect 15381 6199 15439 6205
rect 15473 6205 15485 6208
rect 15519 6205 15531 6239
rect 15473 6199 15531 6205
rect 16209 6239 16267 6245
rect 16209 6205 16221 6239
rect 16255 6205 16267 6239
rect 16209 6199 16267 6205
rect 16393 6239 16451 6245
rect 16393 6205 16405 6239
rect 16439 6205 16451 6239
rect 16393 6199 16451 6205
rect 16485 6239 16543 6245
rect 16485 6205 16497 6239
rect 16531 6236 16543 6239
rect 16761 6239 16819 6245
rect 16761 6236 16773 6239
rect 16531 6208 16773 6236
rect 16531 6205 16543 6208
rect 16485 6199 16543 6205
rect 16761 6205 16773 6208
rect 16807 6236 16819 6239
rect 17586 6236 17592 6248
rect 16807 6208 17592 6236
rect 16807 6205 16819 6208
rect 16761 6199 16819 6205
rect 14645 6171 14703 6177
rect 14292 6140 14596 6168
rect 12768 6128 12774 6140
rect 14274 6100 14280 6112
rect 12452 6072 14280 6100
rect 12069 6063 12127 6069
rect 14274 6060 14280 6072
rect 14332 6060 14338 6112
rect 14458 6060 14464 6112
rect 14516 6060 14522 6112
rect 14568 6100 14596 6140
rect 14645 6137 14657 6171
rect 14691 6168 14703 6171
rect 14737 6171 14795 6177
rect 14737 6168 14749 6171
rect 14691 6140 14749 6168
rect 14691 6137 14703 6140
rect 14645 6131 14703 6137
rect 14737 6137 14749 6140
rect 14783 6137 14795 6171
rect 14737 6131 14795 6137
rect 15212 6168 15240 6199
rect 15657 6171 15715 6177
rect 15657 6168 15669 6171
rect 15212 6140 15669 6168
rect 15212 6112 15240 6140
rect 15657 6137 15669 6140
rect 15703 6137 15715 6171
rect 16408 6168 16436 6199
rect 17586 6196 17592 6208
rect 17644 6196 17650 6248
rect 18046 6196 18052 6248
rect 18104 6236 18110 6248
rect 18141 6239 18199 6245
rect 18141 6236 18153 6239
rect 18104 6208 18153 6236
rect 18104 6196 18110 6208
rect 18141 6205 18153 6208
rect 18187 6205 18199 6239
rect 18141 6199 18199 6205
rect 19426 6196 19432 6248
rect 19484 6236 19490 6248
rect 20257 6239 20315 6245
rect 20257 6236 20269 6239
rect 19484 6208 20269 6236
rect 19484 6196 19490 6208
rect 20257 6205 20269 6208
rect 20303 6205 20315 6239
rect 20625 6239 20683 6245
rect 20625 6236 20637 6239
rect 20257 6199 20315 6205
rect 20456 6208 20637 6236
rect 17678 6168 17684 6180
rect 16408 6140 17684 6168
rect 15657 6131 15715 6137
rect 17678 6128 17684 6140
rect 17736 6128 17742 6180
rect 19518 6128 19524 6180
rect 19576 6168 19582 6180
rect 19990 6171 20048 6177
rect 19990 6168 20002 6171
rect 19576 6140 20002 6168
rect 19576 6128 19582 6140
rect 19990 6137 20002 6140
rect 20036 6137 20048 6171
rect 19990 6131 20048 6137
rect 20456 6112 20484 6208
rect 20625 6205 20637 6208
rect 20671 6205 20683 6239
rect 20625 6199 20683 6205
rect 21450 6196 21456 6248
rect 21508 6196 21514 6248
rect 21729 6239 21787 6245
rect 21729 6205 21741 6239
rect 21775 6205 21787 6239
rect 21729 6199 21787 6205
rect 21744 6112 21772 6199
rect 22554 6196 22560 6248
rect 22612 6196 22618 6248
rect 22830 6196 22836 6248
rect 22888 6196 22894 6248
rect 23474 6196 23480 6248
rect 23532 6236 23538 6248
rect 24486 6245 24492 6248
rect 23845 6239 23903 6245
rect 23845 6236 23857 6239
rect 23532 6208 23857 6236
rect 23532 6196 23538 6208
rect 23845 6205 23857 6208
rect 23891 6205 23903 6239
rect 24480 6236 24492 6245
rect 24447 6208 24492 6236
rect 23845 6199 23903 6205
rect 24480 6199 24492 6208
rect 24486 6196 24492 6199
rect 24544 6196 24550 6248
rect 26142 6196 26148 6248
rect 26200 6236 26206 6248
rect 26237 6239 26295 6245
rect 26237 6236 26249 6239
rect 26200 6208 26249 6236
rect 26200 6196 26206 6208
rect 26237 6205 26249 6208
rect 26283 6205 26295 6239
rect 26237 6199 26295 6205
rect 25682 6128 25688 6180
rect 25740 6168 25746 6180
rect 26973 6171 27031 6177
rect 26973 6168 26985 6171
rect 25740 6140 26985 6168
rect 25740 6128 25746 6140
rect 26973 6137 26985 6140
rect 27019 6137 27031 6171
rect 26973 6131 27031 6137
rect 15194 6100 15200 6112
rect 14568 6072 15200 6100
rect 15194 6060 15200 6072
rect 15252 6060 15258 6112
rect 15838 6060 15844 6112
rect 15896 6060 15902 6112
rect 18874 6060 18880 6112
rect 18932 6060 18938 6112
rect 20438 6060 20444 6112
rect 20496 6060 20502 6112
rect 21726 6060 21732 6112
rect 21784 6060 21790 6112
rect 552 6010 27576 6032
rect 552 5958 7114 6010
rect 7166 5958 7178 6010
rect 7230 5958 7242 6010
rect 7294 5958 7306 6010
rect 7358 5958 7370 6010
rect 7422 5958 13830 6010
rect 13882 5958 13894 6010
rect 13946 5958 13958 6010
rect 14010 5958 14022 6010
rect 14074 5958 14086 6010
rect 14138 5958 20546 6010
rect 20598 5958 20610 6010
rect 20662 5958 20674 6010
rect 20726 5958 20738 6010
rect 20790 5958 20802 6010
rect 20854 5958 27262 6010
rect 27314 5958 27326 6010
rect 27378 5958 27390 6010
rect 27442 5958 27454 6010
rect 27506 5958 27518 6010
rect 27570 5958 27576 6010
rect 552 5936 27576 5958
rect 2682 5856 2688 5908
rect 2740 5856 2746 5908
rect 3602 5856 3608 5908
rect 3660 5896 3666 5908
rect 3697 5899 3755 5905
rect 3697 5896 3709 5899
rect 3660 5868 3709 5896
rect 3660 5856 3666 5868
rect 3697 5865 3709 5868
rect 3743 5865 3755 5899
rect 3697 5859 3755 5865
rect 4522 5856 4528 5908
rect 4580 5856 4586 5908
rect 4798 5856 4804 5908
rect 4856 5856 4862 5908
rect 5810 5856 5816 5908
rect 5868 5856 5874 5908
rect 6730 5856 6736 5908
rect 6788 5896 6794 5908
rect 6825 5899 6883 5905
rect 6825 5896 6837 5899
rect 6788 5868 6837 5896
rect 6788 5856 6794 5868
rect 6825 5865 6837 5868
rect 6871 5865 6883 5899
rect 6825 5859 6883 5865
rect 7742 5856 7748 5908
rect 7800 5896 7806 5908
rect 7837 5899 7895 5905
rect 7837 5896 7849 5899
rect 7800 5868 7849 5896
rect 7800 5856 7806 5868
rect 7837 5865 7849 5868
rect 7883 5865 7895 5899
rect 7837 5859 7895 5865
rect 8110 5856 8116 5908
rect 8168 5856 8174 5908
rect 9125 5899 9183 5905
rect 9125 5865 9137 5899
rect 9171 5896 9183 5899
rect 9674 5896 9680 5908
rect 9171 5868 9680 5896
rect 9171 5865 9183 5868
rect 9125 5859 9183 5865
rect 9674 5856 9680 5868
rect 9732 5856 9738 5908
rect 14182 5896 14188 5908
rect 9784 5868 14188 5896
rect 2314 5720 2320 5772
rect 2372 5720 2378 5772
rect 2700 5769 2728 5856
rect 4816 5828 4844 5856
rect 4816 5800 5580 5828
rect 2685 5763 2743 5769
rect 2685 5729 2697 5763
rect 2731 5729 2743 5763
rect 2685 5723 2743 5729
rect 2958 5720 2964 5772
rect 3016 5720 3022 5772
rect 5258 5720 5264 5772
rect 5316 5720 5322 5772
rect 5552 5769 5580 5800
rect 5828 5769 5856 5856
rect 7760 5800 8064 5828
rect 5537 5763 5595 5769
rect 5537 5729 5549 5763
rect 5583 5729 5595 5763
rect 5537 5723 5595 5729
rect 5813 5763 5871 5769
rect 5813 5729 5825 5763
rect 5859 5729 5871 5763
rect 5813 5723 5871 5729
rect 6086 5720 6092 5772
rect 6144 5720 6150 5772
rect 7650 5720 7656 5772
rect 7708 5760 7714 5772
rect 7760 5769 7788 5800
rect 7745 5763 7803 5769
rect 7745 5760 7757 5763
rect 7708 5732 7757 5760
rect 7708 5720 7714 5732
rect 7745 5729 7757 5732
rect 7791 5729 7803 5763
rect 7745 5723 7803 5729
rect 7926 5720 7932 5772
rect 7984 5720 7990 5772
rect 8036 5769 8064 5800
rect 9490 5788 9496 5840
rect 9548 5828 9554 5840
rect 9784 5828 9812 5868
rect 14182 5856 14188 5868
rect 14240 5856 14246 5908
rect 15013 5899 15071 5905
rect 15013 5896 15025 5899
rect 14844 5868 15025 5896
rect 9548 5800 9812 5828
rect 10260 5831 10318 5837
rect 9548 5788 9554 5800
rect 10260 5797 10272 5831
rect 10306 5828 10318 5831
rect 11606 5828 11612 5840
rect 10306 5800 11612 5828
rect 10306 5797 10318 5800
rect 10260 5791 10318 5797
rect 11606 5788 11612 5800
rect 11664 5788 11670 5840
rect 13538 5828 13544 5840
rect 12544 5800 13544 5828
rect 12544 5772 12572 5800
rect 13538 5788 13544 5800
rect 13596 5788 13602 5840
rect 13722 5788 13728 5840
rect 13780 5828 13786 5840
rect 14844 5828 14872 5868
rect 15013 5865 15025 5868
rect 15059 5865 15071 5899
rect 15013 5859 15071 5865
rect 15102 5856 15108 5908
rect 15160 5856 15166 5908
rect 15838 5856 15844 5908
rect 15896 5856 15902 5908
rect 17586 5856 17592 5908
rect 17644 5856 17650 5908
rect 17678 5856 17684 5908
rect 17736 5856 17742 5908
rect 18322 5896 18328 5908
rect 17880 5868 18328 5896
rect 15120 5828 15148 5856
rect 13780 5800 14872 5828
rect 13780 5788 13786 5800
rect 8021 5763 8079 5769
rect 8021 5729 8033 5763
rect 8067 5729 8079 5763
rect 8021 5723 8079 5729
rect 8205 5763 8263 5769
rect 8205 5729 8217 5763
rect 8251 5729 8263 5763
rect 8205 5723 8263 5729
rect 2590 5652 2596 5704
rect 2648 5652 2654 5704
rect 7944 5692 7972 5720
rect 8220 5692 8248 5723
rect 8294 5720 8300 5772
rect 8352 5720 8358 5772
rect 9674 5720 9680 5772
rect 9732 5760 9738 5772
rect 11149 5763 11207 5769
rect 9732 5732 11100 5760
rect 9732 5720 9738 5732
rect 7944 5664 8248 5692
rect 8312 5624 8340 5720
rect 10502 5652 10508 5704
rect 10560 5652 10566 5704
rect 11072 5701 11100 5732
rect 11149 5729 11161 5763
rect 11195 5729 11207 5763
rect 11149 5723 11207 5729
rect 11057 5695 11115 5701
rect 11057 5661 11069 5695
rect 11103 5661 11115 5695
rect 11057 5655 11115 5661
rect 6380 5596 8340 5624
rect 1210 5516 1216 5568
rect 1268 5556 1274 5568
rect 1305 5559 1363 5565
rect 1305 5556 1317 5559
rect 1268 5528 1317 5556
rect 1268 5516 1274 5528
rect 1305 5525 1317 5528
rect 1351 5525 1363 5559
rect 1305 5519 1363 5525
rect 2130 5516 2136 5568
rect 2188 5516 2194 5568
rect 2501 5559 2559 5565
rect 2501 5525 2513 5559
rect 2547 5556 2559 5559
rect 3234 5556 3240 5568
rect 2547 5528 3240 5556
rect 2547 5525 2559 5528
rect 2501 5519 2559 5525
rect 3234 5516 3240 5528
rect 3292 5556 3298 5568
rect 6380 5556 6408 5596
rect 3292 5528 6408 5556
rect 3292 5516 3298 5528
rect 6914 5516 6920 5568
rect 6972 5516 6978 5568
rect 9766 5516 9772 5568
rect 9824 5556 9830 5568
rect 10134 5556 10140 5568
rect 9824 5528 10140 5556
rect 9824 5516 9830 5528
rect 10134 5516 10140 5528
rect 10192 5556 10198 5568
rect 11164 5556 11192 5723
rect 11790 5720 11796 5772
rect 11848 5760 11854 5772
rect 11974 5760 11980 5772
rect 11848 5732 11980 5760
rect 11848 5720 11854 5732
rect 11974 5720 11980 5732
rect 12032 5760 12038 5772
rect 12250 5760 12256 5772
rect 12032 5732 12256 5760
rect 12032 5720 12038 5732
rect 12250 5720 12256 5732
rect 12308 5720 12314 5772
rect 12342 5720 12348 5772
rect 12400 5720 12406 5772
rect 12526 5720 12532 5772
rect 12584 5720 12590 5772
rect 12894 5720 12900 5772
rect 12952 5760 12958 5772
rect 13265 5763 13323 5769
rect 13265 5760 13277 5763
rect 12952 5732 13277 5760
rect 12952 5720 12958 5732
rect 13265 5729 13277 5732
rect 13311 5729 13323 5763
rect 13265 5723 13323 5729
rect 12986 5652 12992 5704
rect 13044 5652 13050 5704
rect 14844 5692 14872 5800
rect 14936 5800 15148 5828
rect 14936 5769 14964 5800
rect 14921 5763 14979 5769
rect 14921 5729 14933 5763
rect 14967 5729 14979 5763
rect 14921 5723 14979 5729
rect 15105 5763 15163 5769
rect 15105 5729 15117 5763
rect 15151 5760 15163 5763
rect 15856 5760 15884 5856
rect 16669 5831 16727 5837
rect 16669 5797 16681 5831
rect 16715 5828 16727 5831
rect 17696 5828 17724 5856
rect 16715 5800 17724 5828
rect 16715 5797 16727 5800
rect 16669 5791 16727 5797
rect 15151 5732 15884 5760
rect 15151 5729 15163 5732
rect 15105 5723 15163 5729
rect 16574 5720 16580 5772
rect 16632 5720 16638 5772
rect 16761 5763 16819 5769
rect 16761 5729 16773 5763
rect 16807 5760 16819 5763
rect 16850 5760 16856 5772
rect 16807 5732 16856 5760
rect 16807 5729 16819 5732
rect 16761 5723 16819 5729
rect 16850 5720 16856 5732
rect 16908 5720 16914 5772
rect 17773 5763 17831 5769
rect 17773 5729 17785 5763
rect 17819 5760 17831 5763
rect 17880 5760 17908 5868
rect 18322 5856 18328 5868
rect 18380 5896 18386 5908
rect 18417 5899 18475 5905
rect 18417 5896 18429 5899
rect 18380 5868 18429 5896
rect 18380 5856 18386 5868
rect 18417 5865 18429 5868
rect 18463 5865 18475 5899
rect 18417 5859 18475 5865
rect 18874 5856 18880 5908
rect 18932 5856 18938 5908
rect 21450 5856 21456 5908
rect 21508 5856 21514 5908
rect 22554 5856 22560 5908
rect 22612 5856 22618 5908
rect 22830 5856 22836 5908
rect 22888 5856 22894 5908
rect 23385 5899 23443 5905
rect 23385 5865 23397 5899
rect 23431 5865 23443 5899
rect 23385 5859 23443 5865
rect 18340 5800 18644 5828
rect 17819 5732 17908 5760
rect 17819 5729 17831 5732
rect 17773 5723 17831 5729
rect 17954 5720 17960 5772
rect 18012 5720 18018 5772
rect 18046 5720 18052 5772
rect 18104 5720 18110 5772
rect 18138 5720 18144 5772
rect 18196 5720 18202 5772
rect 18340 5769 18368 5800
rect 18616 5769 18644 5800
rect 18325 5763 18383 5769
rect 18325 5729 18337 5763
rect 18371 5729 18383 5763
rect 18325 5723 18383 5729
rect 18417 5763 18475 5769
rect 18417 5729 18429 5763
rect 18463 5729 18475 5763
rect 18417 5723 18475 5729
rect 18601 5763 18659 5769
rect 18601 5729 18613 5763
rect 18647 5760 18659 5763
rect 18892 5760 18920 5856
rect 18647 5732 18920 5760
rect 20993 5763 21051 5769
rect 18647 5729 18659 5732
rect 18601 5723 18659 5729
rect 20993 5729 21005 5763
rect 21039 5760 21051 5763
rect 21468 5760 21496 5856
rect 22572 5769 22600 5856
rect 21039 5732 21496 5760
rect 22557 5763 22615 5769
rect 21039 5729 21051 5732
rect 20993 5723 21051 5729
rect 22557 5729 22569 5763
rect 22603 5729 22615 5763
rect 22557 5723 22615 5729
rect 15286 5692 15292 5704
rect 14844 5664 15292 5692
rect 15286 5652 15292 5664
rect 15344 5652 15350 5704
rect 17972 5692 18000 5720
rect 18233 5695 18291 5701
rect 18233 5692 18245 5695
rect 17972 5664 18245 5692
rect 18233 5661 18245 5664
rect 18279 5661 18291 5695
rect 18233 5655 18291 5661
rect 14001 5627 14059 5633
rect 14001 5593 14013 5627
rect 14047 5624 14059 5627
rect 14458 5624 14464 5636
rect 14047 5596 14464 5624
rect 14047 5593 14059 5596
rect 14001 5587 14059 5593
rect 14458 5584 14464 5596
rect 14516 5624 14522 5636
rect 15010 5624 15016 5636
rect 14516 5596 15016 5624
rect 14516 5584 14522 5596
rect 15010 5584 15016 5596
rect 15068 5584 15074 5636
rect 18138 5584 18144 5636
rect 18196 5624 18202 5636
rect 18432 5624 18460 5723
rect 23014 5720 23020 5772
rect 23072 5720 23078 5772
rect 23198 5720 23204 5772
rect 23256 5720 23262 5772
rect 23400 5760 23428 5859
rect 24302 5856 24308 5908
rect 24360 5896 24366 5908
rect 24489 5899 24547 5905
rect 24489 5896 24501 5899
rect 24360 5868 24501 5896
rect 24360 5856 24366 5868
rect 24489 5865 24501 5868
rect 24535 5865 24547 5899
rect 24489 5859 24547 5865
rect 25406 5856 25412 5908
rect 25464 5856 25470 5908
rect 23753 5763 23811 5769
rect 23753 5760 23765 5763
rect 23400 5732 23765 5760
rect 23753 5729 23765 5732
rect 23799 5729 23811 5763
rect 23753 5723 23811 5729
rect 25593 5763 25651 5769
rect 25593 5729 25605 5763
rect 25639 5760 25651 5763
rect 25774 5760 25780 5772
rect 25639 5732 25780 5760
rect 25639 5729 25651 5732
rect 25593 5723 25651 5729
rect 25774 5720 25780 5732
rect 25832 5720 25838 5772
rect 23474 5652 23480 5704
rect 23532 5652 23538 5704
rect 25682 5652 25688 5704
rect 25740 5652 25746 5704
rect 25869 5695 25927 5701
rect 25869 5661 25881 5695
rect 25915 5692 25927 5695
rect 26142 5692 26148 5704
rect 25915 5664 26148 5692
rect 25915 5661 25927 5664
rect 25869 5655 25927 5661
rect 26142 5652 26148 5664
rect 26200 5652 26206 5704
rect 18196 5596 18460 5624
rect 18196 5584 18202 5596
rect 24302 5584 24308 5636
rect 24360 5624 24366 5636
rect 24581 5627 24639 5633
rect 24581 5624 24593 5627
rect 24360 5596 24593 5624
rect 24360 5584 24366 5596
rect 24581 5593 24593 5596
rect 24627 5593 24639 5627
rect 25700 5624 25728 5652
rect 25777 5627 25835 5633
rect 25777 5624 25789 5627
rect 25700 5596 25789 5624
rect 24581 5587 24639 5593
rect 25777 5593 25789 5596
rect 25823 5593 25835 5627
rect 25777 5587 25835 5593
rect 10192 5528 11192 5556
rect 10192 5516 10198 5528
rect 11514 5516 11520 5568
rect 11572 5516 11578 5568
rect 11793 5559 11851 5565
rect 11793 5525 11805 5559
rect 11839 5556 11851 5559
rect 12066 5556 12072 5568
rect 11839 5528 12072 5556
rect 11839 5525 11851 5528
rect 11793 5519 11851 5525
rect 12066 5516 12072 5528
rect 12124 5516 12130 5568
rect 12710 5516 12716 5568
rect 12768 5516 12774 5568
rect 14182 5516 14188 5568
rect 14240 5516 14246 5568
rect 15562 5516 15568 5568
rect 15620 5556 15626 5568
rect 15657 5559 15715 5565
rect 15657 5556 15669 5559
rect 15620 5528 15669 5556
rect 15620 5516 15626 5528
rect 15657 5525 15669 5528
rect 15703 5525 15715 5559
rect 15657 5519 15715 5525
rect 20714 5516 20720 5568
rect 20772 5556 20778 5568
rect 21542 5556 21548 5568
rect 20772 5528 21548 5556
rect 20772 5516 20778 5528
rect 21542 5516 21548 5528
rect 21600 5516 21606 5568
rect 552 5466 27416 5488
rect 552 5414 3756 5466
rect 3808 5414 3820 5466
rect 3872 5414 3884 5466
rect 3936 5414 3948 5466
rect 4000 5414 4012 5466
rect 4064 5414 10472 5466
rect 10524 5414 10536 5466
rect 10588 5414 10600 5466
rect 10652 5414 10664 5466
rect 10716 5414 10728 5466
rect 10780 5414 17188 5466
rect 17240 5414 17252 5466
rect 17304 5414 17316 5466
rect 17368 5414 17380 5466
rect 17432 5414 17444 5466
rect 17496 5414 23904 5466
rect 23956 5414 23968 5466
rect 24020 5414 24032 5466
rect 24084 5414 24096 5466
rect 24148 5414 24160 5466
rect 24212 5414 27416 5466
rect 552 5392 27416 5414
rect 2222 5312 2228 5364
rect 2280 5312 2286 5364
rect 2685 5355 2743 5361
rect 2685 5321 2697 5355
rect 2731 5352 2743 5355
rect 2958 5352 2964 5364
rect 2731 5324 2964 5352
rect 2731 5321 2743 5324
rect 2685 5315 2743 5321
rect 2958 5312 2964 5324
rect 3016 5312 3022 5364
rect 5077 5355 5135 5361
rect 5077 5321 5089 5355
rect 5123 5352 5135 5355
rect 5258 5352 5264 5364
rect 5123 5324 5264 5352
rect 5123 5321 5135 5324
rect 5077 5315 5135 5321
rect 5258 5312 5264 5324
rect 5316 5312 5322 5364
rect 5905 5355 5963 5361
rect 5905 5321 5917 5355
rect 5951 5352 5963 5355
rect 6086 5352 6092 5364
rect 5951 5324 6092 5352
rect 5951 5321 5963 5324
rect 5905 5315 5963 5321
rect 6086 5312 6092 5324
rect 6144 5312 6150 5364
rect 6914 5352 6920 5364
rect 6656 5324 6920 5352
rect 6656 5225 6684 5324
rect 6914 5312 6920 5324
rect 6972 5312 6978 5364
rect 7650 5312 7656 5364
rect 7708 5312 7714 5364
rect 10229 5355 10287 5361
rect 10229 5321 10241 5355
rect 10275 5352 10287 5355
rect 11882 5352 11888 5364
rect 10275 5324 11888 5352
rect 10275 5321 10287 5324
rect 10229 5315 10287 5321
rect 11882 5312 11888 5324
rect 11940 5312 11946 5364
rect 11974 5312 11980 5364
rect 12032 5352 12038 5364
rect 12713 5355 12771 5361
rect 12032 5324 12434 5352
rect 12032 5312 12038 5324
rect 11238 5244 11244 5296
rect 11296 5244 11302 5296
rect 12406 5284 12434 5324
rect 12713 5321 12725 5355
rect 12759 5352 12771 5355
rect 12894 5352 12900 5364
rect 12759 5324 12900 5352
rect 12759 5321 12771 5324
rect 12713 5315 12771 5321
rect 12894 5312 12900 5324
rect 12952 5312 12958 5364
rect 12986 5312 12992 5364
rect 13044 5312 13050 5364
rect 14292 5324 15148 5352
rect 14292 5284 14320 5324
rect 12406 5256 14320 5284
rect 15120 5284 15148 5324
rect 15194 5312 15200 5364
rect 15252 5312 15258 5364
rect 15672 5324 16528 5352
rect 15672 5284 15700 5324
rect 15120 5256 15700 5284
rect 16500 5284 16528 5324
rect 16574 5312 16580 5364
rect 16632 5312 16638 5364
rect 19978 5352 19984 5364
rect 19628 5324 19984 5352
rect 18690 5284 18696 5296
rect 16500 5256 18696 5284
rect 18690 5244 18696 5256
rect 18748 5244 18754 5296
rect 6641 5219 6699 5225
rect 6641 5185 6653 5219
rect 6687 5185 6699 5219
rect 6641 5179 6699 5185
rect 8757 5219 8815 5225
rect 8757 5185 8769 5219
rect 8803 5216 8815 5219
rect 8846 5216 8852 5228
rect 8803 5188 8852 5216
rect 8803 5185 8815 5188
rect 8757 5179 8815 5185
rect 8846 5176 8852 5188
rect 8904 5176 8910 5228
rect 14182 5176 14188 5228
rect 14240 5176 14246 5228
rect 1118 5108 1124 5160
rect 1176 5108 1182 5160
rect 1210 5108 1216 5160
rect 1268 5108 1274 5160
rect 1489 5151 1547 5157
rect 1489 5117 1501 5151
rect 1535 5117 1547 5151
rect 1489 5111 1547 5117
rect 1504 5080 1532 5111
rect 2130 5108 2136 5160
rect 2188 5148 2194 5160
rect 2685 5151 2743 5157
rect 2685 5148 2697 5151
rect 2188 5120 2697 5148
rect 2188 5108 2194 5120
rect 2685 5117 2697 5120
rect 2731 5117 2743 5151
rect 2685 5111 2743 5117
rect 2869 5151 2927 5157
rect 2869 5117 2881 5151
rect 2915 5148 2927 5151
rect 3326 5148 3332 5160
rect 2915 5120 3332 5148
rect 2915 5117 2927 5120
rect 2869 5111 2927 5117
rect 3326 5108 3332 5120
rect 3384 5108 3390 5160
rect 4893 5151 4951 5157
rect 4893 5117 4905 5151
rect 4939 5148 4951 5151
rect 5074 5148 5080 5160
rect 4939 5120 5080 5148
rect 4939 5117 4951 5120
rect 4893 5111 4951 5117
rect 5074 5108 5080 5120
rect 5132 5108 5138 5160
rect 5718 5108 5724 5160
rect 5776 5108 5782 5160
rect 6362 5108 6368 5160
rect 6420 5108 6426 5160
rect 6917 5151 6975 5157
rect 6917 5117 6929 5151
rect 6963 5117 6975 5151
rect 6917 5111 6975 5117
rect 8481 5151 8539 5157
rect 8481 5117 8493 5151
rect 8527 5117 8539 5151
rect 8481 5111 8539 5117
rect 6932 5080 6960 5111
rect 1504 5052 2774 5080
rect 2746 5012 2774 5052
rect 6564 5052 6960 5080
rect 3418 5012 3424 5024
rect 2746 4984 3424 5012
rect 3418 4972 3424 4984
rect 3476 4972 3482 5024
rect 6564 5021 6592 5052
rect 8496 5024 8524 5111
rect 8570 5108 8576 5160
rect 8628 5108 8634 5160
rect 10045 5151 10103 5157
rect 10045 5117 10057 5151
rect 10091 5117 10103 5151
rect 10045 5111 10103 5117
rect 6549 5015 6607 5021
rect 6549 4981 6561 5015
rect 6595 4981 6607 5015
rect 6549 4975 6607 4981
rect 8478 4972 8484 5024
rect 8536 4972 8542 5024
rect 8754 4972 8760 5024
rect 8812 4972 8818 5024
rect 9582 4972 9588 5024
rect 9640 5012 9646 5024
rect 10060 5012 10088 5111
rect 10226 5108 10232 5160
rect 10284 5148 10290 5160
rect 10505 5151 10563 5157
rect 10505 5148 10517 5151
rect 10284 5120 10517 5148
rect 10284 5108 10290 5120
rect 10505 5117 10517 5120
rect 10551 5117 10563 5151
rect 10505 5111 10563 5117
rect 10778 5108 10784 5160
rect 10836 5108 10842 5160
rect 11977 5151 12035 5157
rect 11977 5117 11989 5151
rect 12023 5117 12035 5151
rect 11977 5111 12035 5117
rect 10413 5083 10471 5089
rect 10413 5049 10425 5083
rect 10459 5080 10471 5083
rect 11514 5080 11520 5092
rect 10459 5052 11520 5080
rect 10459 5049 10471 5052
rect 10413 5043 10471 5049
rect 11514 5040 11520 5052
rect 11572 5040 11578 5092
rect 11992 5080 12020 5111
rect 12066 5108 12072 5160
rect 12124 5148 12130 5160
rect 12253 5151 12311 5157
rect 12253 5148 12265 5151
rect 12124 5120 12265 5148
rect 12124 5108 12130 5120
rect 12253 5117 12265 5120
rect 12299 5117 12311 5151
rect 12253 5111 12311 5117
rect 12529 5151 12587 5157
rect 12529 5117 12541 5151
rect 12575 5117 12587 5151
rect 12529 5111 12587 5117
rect 11992 5052 12112 5080
rect 12084 5024 12112 5052
rect 12158 5040 12164 5092
rect 12216 5080 12222 5092
rect 12544 5080 12572 5111
rect 12710 5108 12716 5160
rect 12768 5108 12774 5160
rect 13078 5108 13084 5160
rect 13136 5108 13142 5160
rect 14458 5108 14464 5160
rect 14516 5108 14522 5160
rect 15286 5108 15292 5160
rect 15344 5108 15350 5160
rect 15562 5108 15568 5160
rect 15620 5108 15626 5160
rect 19628 5157 19656 5324
rect 19978 5312 19984 5324
rect 20036 5352 20042 5364
rect 20714 5352 20720 5364
rect 20036 5324 20720 5352
rect 20036 5312 20042 5324
rect 20714 5312 20720 5324
rect 20772 5312 20778 5364
rect 20993 5355 21051 5361
rect 20993 5321 21005 5355
rect 21039 5352 21051 5355
rect 21726 5352 21732 5364
rect 21039 5324 21732 5352
rect 21039 5321 21051 5324
rect 20993 5315 21051 5321
rect 21726 5312 21732 5324
rect 21784 5352 21790 5364
rect 22741 5355 22799 5361
rect 22741 5352 22753 5355
rect 21784 5324 22753 5352
rect 21784 5312 21790 5324
rect 22741 5321 22753 5324
rect 22787 5321 22799 5355
rect 22741 5315 22799 5321
rect 23109 5355 23167 5361
rect 23109 5321 23121 5355
rect 23155 5352 23167 5355
rect 23198 5352 23204 5364
rect 23155 5324 23204 5352
rect 23155 5321 23167 5324
rect 23109 5315 23167 5321
rect 23198 5312 23204 5324
rect 23256 5312 23262 5364
rect 23750 5312 23756 5364
rect 23808 5352 23814 5364
rect 24486 5352 24492 5364
rect 23808 5324 24492 5352
rect 23808 5312 23814 5324
rect 24486 5312 24492 5324
rect 24544 5352 24550 5364
rect 25869 5355 25927 5361
rect 25869 5352 25881 5355
rect 24544 5324 25881 5352
rect 24544 5312 24550 5324
rect 25869 5321 25881 5324
rect 25915 5352 25927 5355
rect 26326 5352 26332 5364
rect 25915 5324 26332 5352
rect 25915 5321 25927 5324
rect 25869 5315 25927 5321
rect 26326 5312 26332 5324
rect 26384 5312 26390 5364
rect 26421 5355 26479 5361
rect 26421 5321 26433 5355
rect 26467 5321 26479 5355
rect 26421 5315 26479 5321
rect 19812 5256 21220 5284
rect 19812 5160 19840 5256
rect 21192 5228 21220 5256
rect 21542 5244 21548 5296
rect 21600 5244 21606 5296
rect 25774 5244 25780 5296
rect 25832 5284 25838 5296
rect 26436 5284 26464 5315
rect 25832 5256 26464 5284
rect 25832 5244 25838 5256
rect 20272 5188 20852 5216
rect 15841 5151 15899 5157
rect 15841 5117 15853 5151
rect 15887 5117 15899 5151
rect 15841 5111 15899 5117
rect 19613 5151 19671 5157
rect 19613 5117 19625 5151
rect 19659 5117 19671 5151
rect 19613 5111 19671 5117
rect 13096 5080 13124 5108
rect 15856 5080 15884 5111
rect 19794 5108 19800 5160
rect 19852 5108 19858 5160
rect 20272 5089 20300 5188
rect 20346 5108 20352 5160
rect 20404 5148 20410 5160
rect 20533 5151 20591 5157
rect 20533 5148 20545 5151
rect 20404 5120 20545 5148
rect 20404 5108 20410 5120
rect 20533 5117 20545 5120
rect 20579 5117 20591 5151
rect 20533 5111 20591 5117
rect 20714 5108 20720 5160
rect 20772 5108 20778 5160
rect 20824 5157 20852 5188
rect 21174 5176 21180 5228
rect 21232 5176 21238 5228
rect 21637 5219 21695 5225
rect 21637 5185 21649 5219
rect 21683 5216 21695 5219
rect 26513 5219 26571 5225
rect 26513 5216 26525 5219
rect 21683 5188 22048 5216
rect 21683 5185 21695 5188
rect 21637 5179 21695 5185
rect 20809 5151 20867 5157
rect 20809 5117 20821 5151
rect 20855 5117 20867 5151
rect 20993 5151 21051 5157
rect 20993 5148 21005 5151
rect 20809 5111 20867 5117
rect 20916 5120 21005 5148
rect 20916 5092 20944 5120
rect 20993 5117 21005 5120
rect 21039 5148 21051 5151
rect 21450 5148 21456 5160
rect 21039 5120 21456 5148
rect 21039 5117 21051 5120
rect 20993 5111 21051 5117
rect 21450 5108 21456 5120
rect 21508 5148 21514 5160
rect 21729 5151 21787 5157
rect 21729 5148 21741 5151
rect 21508 5120 21741 5148
rect 21508 5108 21514 5120
rect 21729 5117 21741 5120
rect 21775 5117 21787 5151
rect 21729 5111 21787 5117
rect 21913 5151 21971 5157
rect 21913 5117 21925 5151
rect 21959 5148 21971 5151
rect 22020 5148 22048 5188
rect 25608 5188 26525 5216
rect 25608 5160 25636 5188
rect 26513 5185 26525 5188
rect 26559 5185 26571 5219
rect 26513 5179 26571 5185
rect 22189 5151 22247 5157
rect 22189 5148 22201 5151
rect 21959 5120 22201 5148
rect 21959 5117 21971 5120
rect 21913 5111 21971 5117
rect 22189 5117 22201 5120
rect 22235 5117 22247 5151
rect 22189 5111 22247 5117
rect 22738 5108 22744 5160
rect 22796 5108 22802 5160
rect 22922 5108 22928 5160
rect 22980 5108 22986 5160
rect 23750 5108 23756 5160
rect 23808 5148 23814 5160
rect 24121 5151 24179 5157
rect 24121 5148 24133 5151
rect 23808 5120 24133 5148
rect 23808 5108 23814 5120
rect 24121 5117 24133 5120
rect 24167 5117 24179 5151
rect 24121 5111 24179 5117
rect 24578 5108 24584 5160
rect 24636 5108 24642 5160
rect 25590 5108 25596 5160
rect 25648 5108 25654 5160
rect 26050 5108 26056 5160
rect 26108 5148 26114 5160
rect 26421 5151 26479 5157
rect 26421 5148 26433 5151
rect 26108 5120 26433 5148
rect 26108 5108 26114 5120
rect 26421 5117 26433 5120
rect 26467 5117 26479 5151
rect 26421 5111 26479 5117
rect 12216 5052 13124 5080
rect 15488 5052 15884 5080
rect 19981 5083 20039 5089
rect 12216 5040 12222 5052
rect 11330 5012 11336 5024
rect 9640 4984 11336 5012
rect 9640 4972 9646 4984
rect 11330 4972 11336 4984
rect 11388 5012 11394 5024
rect 11882 5012 11888 5024
rect 11388 4984 11888 5012
rect 11388 4972 11394 4984
rect 11882 4972 11888 4984
rect 11940 4972 11946 5024
rect 12066 4972 12072 5024
rect 12124 4972 12130 5024
rect 15488 5021 15516 5052
rect 19981 5049 19993 5083
rect 20027 5080 20039 5083
rect 20257 5083 20315 5089
rect 20257 5080 20269 5083
rect 20027 5052 20269 5080
rect 20027 5049 20039 5052
rect 19981 5043 20039 5049
rect 20257 5049 20269 5052
rect 20303 5049 20315 5083
rect 20257 5043 20315 5049
rect 20441 5083 20499 5089
rect 20441 5049 20453 5083
rect 20487 5049 20499 5083
rect 20441 5043 20499 5049
rect 20625 5083 20683 5089
rect 20625 5049 20637 5083
rect 20671 5080 20683 5083
rect 20898 5080 20904 5092
rect 20671 5052 20904 5080
rect 20671 5049 20683 5052
rect 20625 5043 20683 5049
rect 15473 5015 15531 5021
rect 15473 4981 15485 5015
rect 15519 4981 15531 5015
rect 15473 4975 15531 4981
rect 20070 4972 20076 5024
rect 20128 4972 20134 5024
rect 20162 4972 20168 5024
rect 20220 5012 20226 5024
rect 20456 5012 20484 5043
rect 20898 5040 20904 5052
rect 20956 5040 20962 5092
rect 21082 5040 21088 5092
rect 21140 5040 21146 5092
rect 20714 5012 20720 5024
rect 20220 4984 20720 5012
rect 20220 4972 20226 4984
rect 20714 4972 20720 4984
rect 20772 5012 20778 5024
rect 21100 5012 21128 5040
rect 20772 4984 21128 5012
rect 20772 4972 20778 4984
rect 22094 4972 22100 5024
rect 22152 4972 22158 5024
rect 22186 4972 22192 5024
rect 22244 5012 22250 5024
rect 22281 5015 22339 5021
rect 22281 5012 22293 5015
rect 22244 4984 22293 5012
rect 22244 4972 22250 4984
rect 22281 4981 22293 4984
rect 22327 4981 22339 5015
rect 22281 4975 22339 4981
rect 26786 4972 26792 5024
rect 26844 4972 26850 5024
rect 552 4922 27576 4944
rect 552 4870 7114 4922
rect 7166 4870 7178 4922
rect 7230 4870 7242 4922
rect 7294 4870 7306 4922
rect 7358 4870 7370 4922
rect 7422 4870 13830 4922
rect 13882 4870 13894 4922
rect 13946 4870 13958 4922
rect 14010 4870 14022 4922
rect 14074 4870 14086 4922
rect 14138 4870 20546 4922
rect 20598 4870 20610 4922
rect 20662 4870 20674 4922
rect 20726 4870 20738 4922
rect 20790 4870 20802 4922
rect 20854 4870 27262 4922
rect 27314 4870 27326 4922
rect 27378 4870 27390 4922
rect 27442 4870 27454 4922
rect 27506 4870 27518 4922
rect 27570 4870 27576 4922
rect 552 4848 27576 4870
rect 1118 4768 1124 4820
rect 1176 4768 1182 4820
rect 1946 4768 1952 4820
rect 2004 4808 2010 4820
rect 2225 4811 2283 4817
rect 2225 4808 2237 4811
rect 2004 4780 2237 4808
rect 2004 4768 2010 4780
rect 2225 4777 2237 4780
rect 2271 4777 2283 4811
rect 2225 4771 2283 4777
rect 5718 4768 5724 4820
rect 5776 4808 5782 4820
rect 5813 4811 5871 4817
rect 5813 4808 5825 4811
rect 5776 4780 5825 4808
rect 5776 4768 5782 4780
rect 5813 4777 5825 4780
rect 5859 4777 5871 4811
rect 5813 4771 5871 4777
rect 8202 4768 8208 4820
rect 8260 4768 8266 4820
rect 8754 4768 8760 4820
rect 8812 4808 8818 4820
rect 9141 4811 9199 4817
rect 9141 4808 9153 4811
rect 8812 4780 9153 4808
rect 8812 4768 8818 4780
rect 9141 4777 9153 4780
rect 9187 4777 9199 4811
rect 9141 4771 9199 4777
rect 9766 4768 9772 4820
rect 9824 4768 9830 4820
rect 10778 4768 10784 4820
rect 10836 4768 10842 4820
rect 12250 4768 12256 4820
rect 12308 4808 12314 4820
rect 14369 4811 14427 4817
rect 12308 4780 12756 4808
rect 12308 4768 12314 4780
rect 1136 4672 1164 4768
rect 2590 4700 2596 4752
rect 2648 4740 2654 4752
rect 3145 4743 3203 4749
rect 2648 4712 3004 4740
rect 2648 4700 2654 4712
rect 1213 4675 1271 4681
rect 1213 4672 1225 4675
rect 1136 4644 1225 4672
rect 1213 4641 1225 4644
rect 1259 4641 1271 4675
rect 1213 4635 1271 4641
rect 1489 4675 1547 4681
rect 1489 4641 1501 4675
rect 1535 4672 1547 4675
rect 2130 4672 2136 4684
rect 1535 4644 2136 4672
rect 1535 4641 1547 4644
rect 1489 4635 1547 4641
rect 2130 4632 2136 4644
rect 2188 4632 2194 4684
rect 2976 4681 3004 4712
rect 3145 4709 3157 4743
rect 3191 4740 3203 4743
rect 4154 4740 4160 4752
rect 3191 4712 3372 4740
rect 3191 4709 3203 4712
rect 3145 4703 3203 4709
rect 3344 4684 3372 4712
rect 3436 4712 4160 4740
rect 2961 4675 3019 4681
rect 2961 4641 2973 4675
rect 3007 4672 3019 4675
rect 3050 4672 3056 4684
rect 3007 4644 3056 4672
rect 3007 4641 3019 4644
rect 2961 4635 3019 4641
rect 3050 4632 3056 4644
rect 3108 4632 3114 4684
rect 3237 4675 3295 4681
rect 3237 4641 3249 4675
rect 3283 4641 3295 4675
rect 3237 4635 3295 4641
rect 2590 4564 2596 4616
rect 2648 4604 2654 4616
rect 2777 4607 2835 4613
rect 2777 4604 2789 4607
rect 2648 4576 2789 4604
rect 2648 4564 2654 4576
rect 2777 4573 2789 4576
rect 2823 4604 2835 4607
rect 3252 4604 3280 4635
rect 3326 4632 3332 4684
rect 3384 4632 3390 4684
rect 3436 4681 3464 4712
rect 4154 4700 4160 4712
rect 4212 4740 4218 4752
rect 8294 4740 8300 4752
rect 4212 4712 5028 4740
rect 4212 4700 4218 4712
rect 3421 4675 3479 4681
rect 3421 4641 3433 4675
rect 3467 4641 3479 4675
rect 3421 4635 3479 4641
rect 2823 4576 3280 4604
rect 3436 4604 3464 4635
rect 3510 4632 3516 4684
rect 3568 4632 3574 4684
rect 3697 4675 3755 4681
rect 3697 4641 3709 4675
rect 3743 4672 3755 4675
rect 4338 4672 4344 4684
rect 3743 4644 4344 4672
rect 3743 4641 3755 4644
rect 3697 4635 3755 4641
rect 4338 4632 4344 4644
rect 4396 4632 4402 4684
rect 4798 4672 4804 4684
rect 4632 4644 4804 4672
rect 3605 4607 3663 4613
rect 3605 4604 3617 4607
rect 3436 4576 3617 4604
rect 2823 4573 2835 4576
rect 2777 4567 2835 4573
rect 3605 4573 3617 4576
rect 3651 4573 3663 4607
rect 3605 4567 3663 4573
rect 4157 4607 4215 4613
rect 4157 4573 4169 4607
rect 4203 4604 4215 4607
rect 4246 4604 4252 4616
rect 4203 4576 4252 4604
rect 4203 4573 4215 4576
rect 4157 4567 4215 4573
rect 4246 4564 4252 4576
rect 4304 4564 4310 4616
rect 4632 4613 4660 4644
rect 4798 4632 4804 4644
rect 4856 4672 4862 4684
rect 4893 4675 4951 4681
rect 4893 4672 4905 4675
rect 4856 4644 4905 4672
rect 4856 4632 4862 4644
rect 4893 4641 4905 4644
rect 4939 4641 4951 4675
rect 4893 4635 4951 4641
rect 4617 4607 4675 4613
rect 4617 4573 4629 4607
rect 4663 4573 4675 4607
rect 4617 4567 4675 4573
rect 4709 4607 4767 4613
rect 4709 4573 4721 4607
rect 4755 4604 4767 4607
rect 5000 4604 5028 4712
rect 7944 4712 8300 4740
rect 5077 4675 5135 4681
rect 5077 4641 5089 4675
rect 5123 4672 5135 4675
rect 5169 4675 5227 4681
rect 5169 4672 5181 4675
rect 5123 4644 5181 4672
rect 5123 4641 5135 4644
rect 5077 4635 5135 4641
rect 5169 4641 5181 4644
rect 5215 4641 5227 4675
rect 5169 4635 5227 4641
rect 5534 4632 5540 4684
rect 5592 4672 5598 4684
rect 7944 4681 7972 4712
rect 8294 4700 8300 4712
rect 8352 4700 8358 4752
rect 8570 4740 8576 4752
rect 8404 4712 8576 4740
rect 8404 4681 8432 4712
rect 8570 4700 8576 4712
rect 8628 4700 8634 4752
rect 8941 4743 8999 4749
rect 8941 4709 8953 4743
rect 8987 4740 8999 4743
rect 9030 4740 9036 4752
rect 8987 4712 9036 4740
rect 8987 4709 8999 4712
rect 8941 4703 8999 4709
rect 9030 4700 9036 4712
rect 9088 4740 9094 4752
rect 9582 4740 9588 4752
rect 9088 4712 9588 4740
rect 9088 4700 9094 4712
rect 9582 4700 9588 4712
rect 9640 4700 9646 4752
rect 10686 4700 10692 4752
rect 10744 4700 10750 4752
rect 6181 4675 6239 4681
rect 6181 4672 6193 4675
rect 5592 4644 6193 4672
rect 5592 4632 5598 4644
rect 6181 4641 6193 4644
rect 6227 4641 6239 4675
rect 6181 4635 6239 4641
rect 7469 4675 7527 4681
rect 7469 4641 7481 4675
rect 7515 4641 7527 4675
rect 7469 4635 7527 4641
rect 7653 4675 7711 4681
rect 7653 4641 7665 4675
rect 7699 4672 7711 4675
rect 7929 4675 7987 4681
rect 7929 4672 7941 4675
rect 7699 4644 7941 4672
rect 7699 4641 7711 4644
rect 7653 4635 7711 4641
rect 7929 4641 7941 4644
rect 7975 4641 7987 4675
rect 7929 4635 7987 4641
rect 8113 4675 8171 4681
rect 8113 4641 8125 4675
rect 8159 4672 8171 4675
rect 8389 4675 8447 4681
rect 8389 4672 8401 4675
rect 8159 4644 8401 4672
rect 8159 4641 8171 4644
rect 8113 4635 8171 4641
rect 8389 4641 8401 4644
rect 8435 4641 8447 4675
rect 8665 4675 8723 4681
rect 8665 4672 8677 4675
rect 8389 4635 8447 4641
rect 8496 4644 8677 4672
rect 4755 4576 5028 4604
rect 4755 4573 4767 4576
rect 4709 4567 4767 4573
rect 5994 4564 6000 4616
rect 6052 4604 6058 4616
rect 6089 4607 6147 4613
rect 6089 4604 6101 4607
rect 6052 4576 6101 4604
rect 6052 4564 6058 4576
rect 6089 4573 6101 4576
rect 6135 4573 6147 4607
rect 7484 4604 7512 4635
rect 7745 4607 7803 4613
rect 7745 4604 7757 4607
rect 7484 4576 7757 4604
rect 6089 4567 6147 4573
rect 7745 4573 7757 4576
rect 7791 4604 7803 4607
rect 8018 4604 8024 4616
rect 7791 4576 8024 4604
rect 7791 4573 7803 4576
rect 7745 4567 7803 4573
rect 8018 4564 8024 4576
rect 8076 4564 8082 4616
rect 8496 4548 8524 4644
rect 8665 4641 8677 4644
rect 8711 4641 8723 4675
rect 8665 4635 8723 4641
rect 8846 4632 8852 4684
rect 8904 4632 8910 4684
rect 9401 4675 9459 4681
rect 9401 4672 9413 4675
rect 9324 4644 9413 4672
rect 3418 4496 3424 4548
rect 3476 4536 3482 4548
rect 3476 4508 4108 4536
rect 3476 4496 3482 4508
rect 4080 4468 4108 4508
rect 4430 4496 4436 4548
rect 4488 4496 4494 4548
rect 7653 4539 7711 4545
rect 4540 4508 6040 4536
rect 4540 4468 4568 4508
rect 4080 4440 4568 4468
rect 5353 4471 5411 4477
rect 5353 4437 5365 4471
rect 5399 4468 5411 4471
rect 5442 4468 5448 4480
rect 5399 4440 5448 4468
rect 5399 4437 5411 4440
rect 5353 4431 5411 4437
rect 5442 4428 5448 4440
rect 5500 4428 5506 4480
rect 6012 4477 6040 4508
rect 7653 4505 7665 4539
rect 7699 4536 7711 4539
rect 8478 4536 8484 4548
rect 7699 4508 8484 4536
rect 7699 4505 7711 4508
rect 7653 4499 7711 4505
rect 8478 4496 8484 4508
rect 8536 4496 8542 4548
rect 9324 4545 9352 4644
rect 9401 4641 9413 4644
rect 9447 4641 9459 4675
rect 9401 4635 9459 4641
rect 10505 4675 10563 4681
rect 10505 4641 10517 4675
rect 10551 4672 10563 4675
rect 10704 4672 10732 4700
rect 10796 4681 10824 4768
rect 11149 4743 11207 4749
rect 11149 4709 11161 4743
rect 11195 4740 11207 4743
rect 11517 4743 11575 4749
rect 11517 4740 11529 4743
rect 11195 4712 11529 4740
rect 11195 4709 11207 4712
rect 11149 4703 11207 4709
rect 11517 4709 11529 4712
rect 11563 4740 11575 4743
rect 11563 4712 12020 4740
rect 11563 4709 11575 4712
rect 11517 4703 11575 4709
rect 10551 4644 10732 4672
rect 10781 4675 10839 4681
rect 10551 4641 10563 4644
rect 10505 4635 10563 4641
rect 10781 4641 10793 4675
rect 10827 4641 10839 4675
rect 10781 4635 10839 4641
rect 11238 4632 11244 4684
rect 11296 4672 11302 4684
rect 11333 4675 11391 4681
rect 11333 4672 11345 4675
rect 11296 4644 11345 4672
rect 11296 4632 11302 4644
rect 11333 4641 11345 4644
rect 11379 4641 11391 4675
rect 11333 4635 11391 4641
rect 11701 4675 11759 4681
rect 11701 4641 11713 4675
rect 11747 4672 11759 4675
rect 11790 4672 11796 4684
rect 11747 4644 11796 4672
rect 11747 4641 11759 4644
rect 11701 4635 11759 4641
rect 11790 4632 11796 4644
rect 11848 4632 11854 4684
rect 11992 4681 12020 4712
rect 12066 4700 12072 4752
rect 12124 4740 12130 4752
rect 12728 4749 12756 4780
rect 14369 4777 14381 4811
rect 14415 4808 14427 4811
rect 14458 4808 14464 4820
rect 14415 4780 14464 4808
rect 14415 4777 14427 4780
rect 14369 4771 14427 4777
rect 14458 4768 14464 4780
rect 14516 4768 14522 4820
rect 15105 4811 15163 4817
rect 15105 4777 15117 4811
rect 15151 4808 15163 4811
rect 15286 4808 15292 4820
rect 15151 4780 15292 4808
rect 15151 4777 15163 4780
rect 15105 4771 15163 4777
rect 15286 4768 15292 4780
rect 15344 4768 15350 4820
rect 18046 4768 18052 4820
rect 18104 4808 18110 4820
rect 18141 4811 18199 4817
rect 18141 4808 18153 4811
rect 18104 4780 18153 4808
rect 18104 4768 18110 4780
rect 18141 4777 18153 4780
rect 18187 4777 18199 4811
rect 18141 4771 18199 4777
rect 21450 4768 21456 4820
rect 21508 4817 21514 4820
rect 21508 4811 21527 4817
rect 21515 4777 21527 4811
rect 21508 4771 21527 4777
rect 21508 4768 21514 4771
rect 22094 4768 22100 4820
rect 22152 4768 22158 4820
rect 23477 4811 23535 4817
rect 23477 4777 23489 4811
rect 23523 4777 23535 4811
rect 23477 4771 23535 4777
rect 23937 4811 23995 4817
rect 23937 4777 23949 4811
rect 23983 4777 23995 4811
rect 23937 4771 23995 4777
rect 12713 4743 12771 4749
rect 12124 4712 12664 4740
rect 12124 4700 12130 4712
rect 11885 4675 11943 4681
rect 11885 4641 11897 4675
rect 11931 4641 11943 4675
rect 11885 4635 11943 4641
rect 11977 4675 12035 4681
rect 11977 4641 11989 4675
rect 12023 4641 12035 4675
rect 11977 4635 12035 4641
rect 12161 4675 12219 4681
rect 12161 4641 12173 4675
rect 12207 4641 12219 4675
rect 12161 4635 12219 4641
rect 12253 4675 12311 4681
rect 12253 4641 12265 4675
rect 12299 4641 12311 4675
rect 12253 4635 12311 4641
rect 12437 4675 12495 4681
rect 12437 4641 12449 4675
rect 12483 4672 12495 4675
rect 12526 4672 12532 4684
rect 12483 4644 12532 4672
rect 12483 4641 12495 4644
rect 12437 4635 12495 4641
rect 11900 4604 11928 4635
rect 12066 4604 12072 4616
rect 11900 4576 12072 4604
rect 12066 4564 12072 4576
rect 12124 4564 12130 4616
rect 9309 4539 9367 4545
rect 9309 4505 9321 4539
rect 9355 4505 9367 4539
rect 12176 4536 12204 4635
rect 12268 4604 12296 4635
rect 12526 4632 12532 4644
rect 12584 4632 12590 4684
rect 12636 4672 12664 4712
rect 12713 4709 12725 4743
rect 12759 4709 12771 4743
rect 20070 4740 20076 4752
rect 12713 4703 12771 4709
rect 12993 4712 13584 4740
rect 12993 4672 13021 4712
rect 13446 4672 13452 4684
rect 12636 4644 13021 4672
rect 13188 4644 13452 4672
rect 12802 4604 12808 4616
rect 12268 4576 12808 4604
rect 12802 4564 12808 4576
rect 12860 4564 12866 4616
rect 13188 4613 13216 4644
rect 13446 4632 13452 4644
rect 13504 4632 13510 4684
rect 13173 4607 13231 4613
rect 13173 4573 13185 4607
rect 13219 4573 13231 4607
rect 13173 4567 13231 4573
rect 13265 4607 13323 4613
rect 13265 4573 13277 4607
rect 13311 4573 13323 4607
rect 13556 4604 13584 4712
rect 19904 4712 20076 4740
rect 13633 4675 13691 4681
rect 13633 4641 13645 4675
rect 13679 4672 13691 4675
rect 13725 4675 13783 4681
rect 13725 4672 13737 4675
rect 13679 4644 13737 4672
rect 13679 4641 13691 4644
rect 13633 4635 13691 4641
rect 13725 4641 13737 4644
rect 13771 4641 13783 4675
rect 13725 4635 13783 4641
rect 14182 4632 14188 4684
rect 14240 4632 14246 4684
rect 14734 4632 14740 4684
rect 14792 4632 14798 4684
rect 14918 4632 14924 4684
rect 14976 4632 14982 4684
rect 16574 4632 16580 4684
rect 16632 4632 16638 4684
rect 17497 4675 17555 4681
rect 17497 4641 17509 4675
rect 17543 4672 17555 4675
rect 17586 4672 17592 4684
rect 17543 4644 17592 4672
rect 17543 4641 17555 4644
rect 17497 4635 17555 4641
rect 17586 4632 17592 4644
rect 17644 4632 17650 4684
rect 17678 4632 17684 4684
rect 17736 4632 17742 4684
rect 17957 4675 18015 4681
rect 17957 4672 17969 4675
rect 17880 4644 17969 4672
rect 17880 4616 17908 4644
rect 17957 4641 17969 4644
rect 18003 4641 18015 4675
rect 17957 4635 18015 4641
rect 19334 4632 19340 4684
rect 19392 4681 19398 4684
rect 19392 4635 19404 4681
rect 19392 4632 19398 4635
rect 19702 4632 19708 4684
rect 19760 4672 19766 4684
rect 19904 4681 19932 4712
rect 20070 4700 20076 4712
rect 20128 4700 20134 4752
rect 21174 4700 21180 4752
rect 21232 4740 21238 4752
rect 21269 4743 21327 4749
rect 21269 4740 21281 4743
rect 21232 4712 21281 4740
rect 21232 4700 21238 4712
rect 21269 4709 21281 4712
rect 21315 4709 21327 4743
rect 22112 4740 22140 4768
rect 21269 4703 21327 4709
rect 22020 4712 22140 4740
rect 23017 4743 23075 4749
rect 22020 4681 22048 4712
rect 23017 4709 23029 4743
rect 23063 4740 23075 4743
rect 23063 4712 23428 4740
rect 23063 4709 23075 4712
rect 23017 4703 23075 4709
rect 23400 4684 23428 4712
rect 19889 4675 19947 4681
rect 19889 4672 19901 4675
rect 19760 4644 19901 4672
rect 19760 4632 19766 4644
rect 19889 4641 19901 4644
rect 19935 4641 19947 4675
rect 19889 4635 19947 4641
rect 21997 4675 22055 4681
rect 21997 4641 22009 4675
rect 22043 4641 22055 4675
rect 21997 4635 22055 4641
rect 22281 4675 22339 4681
rect 22281 4641 22293 4675
rect 22327 4641 22339 4675
rect 22281 4635 22339 4641
rect 23293 4675 23351 4681
rect 23293 4641 23305 4675
rect 23339 4641 23351 4675
rect 23293 4635 23351 4641
rect 15933 4607 15991 4613
rect 13556 4576 14780 4604
rect 13265 4567 13323 4573
rect 12253 4539 12311 4545
rect 12253 4536 12265 4539
rect 12176 4508 12265 4536
rect 9309 4499 9367 4505
rect 12253 4505 12265 4508
rect 12299 4505 12311 4539
rect 12253 4499 12311 4505
rect 5997 4471 6055 4477
rect 5997 4437 6009 4471
rect 6043 4437 6055 4471
rect 5997 4431 6055 4437
rect 7006 4428 7012 4480
rect 7064 4468 7070 4480
rect 7101 4471 7159 4477
rect 7101 4468 7113 4471
rect 7064 4440 7113 4468
rect 7064 4428 7070 4440
rect 7101 4437 7113 4440
rect 7147 4437 7159 4471
rect 7101 4431 7159 4437
rect 9122 4428 9128 4480
rect 9180 4428 9186 4480
rect 9585 4471 9643 4477
rect 9585 4437 9597 4471
rect 9631 4468 9643 4471
rect 9674 4468 9680 4480
rect 9631 4440 9680 4468
rect 9631 4437 9643 4440
rect 9585 4431 9643 4437
rect 9674 4428 9680 4440
rect 9732 4428 9738 4480
rect 10962 4428 10968 4480
rect 11020 4428 11026 4480
rect 12268 4468 12296 4499
rect 13078 4496 13084 4548
rect 13136 4496 13142 4548
rect 12802 4468 12808 4480
rect 12268 4440 12808 4468
rect 12802 4428 12808 4440
rect 12860 4468 12866 4480
rect 13170 4468 13176 4480
rect 12860 4440 13176 4468
rect 12860 4428 12866 4440
rect 13170 4428 13176 4440
rect 13228 4468 13234 4480
rect 13280 4468 13308 4567
rect 13228 4440 13308 4468
rect 13909 4471 13967 4477
rect 13228 4428 13234 4440
rect 13909 4437 13921 4471
rect 13955 4468 13967 4471
rect 14274 4468 14280 4480
rect 13955 4440 14280 4468
rect 13955 4437 13967 4440
rect 13909 4431 13967 4437
rect 14274 4428 14280 4440
rect 14332 4428 14338 4480
rect 14752 4477 14780 4576
rect 15933 4573 15945 4607
rect 15979 4604 15991 4607
rect 16301 4607 16359 4613
rect 16301 4604 16313 4607
rect 15979 4576 16313 4604
rect 15979 4573 15991 4576
rect 15933 4567 15991 4573
rect 16301 4573 16313 4576
rect 16347 4573 16359 4607
rect 16301 4567 16359 4573
rect 17862 4564 17868 4616
rect 17920 4564 17926 4616
rect 19613 4607 19671 4613
rect 19613 4573 19625 4607
rect 19659 4573 19671 4607
rect 22296 4604 22324 4635
rect 19613 4567 19671 4573
rect 21652 4576 22324 4604
rect 17313 4539 17371 4545
rect 17313 4505 17325 4539
rect 17359 4536 17371 4539
rect 18138 4536 18144 4548
rect 17359 4508 18144 4536
rect 17359 4505 17371 4508
rect 17313 4499 17371 4505
rect 18138 4496 18144 4508
rect 18196 4496 18202 4548
rect 14737 4471 14795 4477
rect 14737 4437 14749 4471
rect 14783 4437 14795 4471
rect 14737 4431 14795 4437
rect 18230 4428 18236 4480
rect 18288 4428 18294 4480
rect 19426 4428 19432 4480
rect 19484 4468 19490 4480
rect 19628 4468 19656 4567
rect 19981 4539 20039 4545
rect 19981 4505 19993 4539
rect 20027 4536 20039 4539
rect 20438 4536 20444 4548
rect 20027 4508 20444 4536
rect 20027 4505 20039 4508
rect 19981 4499 20039 4505
rect 20438 4496 20444 4508
rect 20496 4536 20502 4548
rect 21652 4545 21680 4576
rect 22554 4564 22560 4616
rect 22612 4604 22618 4616
rect 23109 4607 23167 4613
rect 23109 4604 23121 4607
rect 22612 4576 23121 4604
rect 22612 4564 22618 4576
rect 23109 4573 23121 4576
rect 23155 4573 23167 4607
rect 23109 4567 23167 4573
rect 21637 4539 21695 4545
rect 20496 4508 21588 4536
rect 20496 4496 20502 4508
rect 19484 4440 19656 4468
rect 19484 4428 19490 4440
rect 21358 4428 21364 4480
rect 21416 4468 21422 4480
rect 21453 4471 21511 4477
rect 21453 4468 21465 4471
rect 21416 4440 21465 4468
rect 21416 4428 21422 4440
rect 21453 4437 21465 4440
rect 21499 4437 21511 4471
rect 21560 4468 21588 4508
rect 21637 4505 21649 4539
rect 21683 4505 21695 4539
rect 23308 4536 23336 4635
rect 23382 4632 23388 4684
rect 23440 4632 23446 4684
rect 23492 4672 23520 4771
rect 23753 4675 23811 4681
rect 23753 4672 23765 4675
rect 23492 4644 23765 4672
rect 23753 4641 23765 4644
rect 23799 4641 23811 4675
rect 23952 4672 23980 4771
rect 25038 4768 25044 4820
rect 25096 4768 25102 4820
rect 25774 4808 25780 4820
rect 25148 4780 25780 4808
rect 25148 4681 25176 4780
rect 25774 4768 25780 4780
rect 25832 4768 25838 4820
rect 26142 4768 26148 4820
rect 26200 4768 26206 4820
rect 26621 4811 26679 4817
rect 26621 4808 26633 4811
rect 26252 4780 26633 4808
rect 25409 4743 25467 4749
rect 25409 4709 25421 4743
rect 25455 4740 25467 4743
rect 26252 4740 26280 4780
rect 26621 4777 26633 4780
rect 26667 4777 26679 4811
rect 26621 4771 26679 4777
rect 26789 4811 26847 4817
rect 26789 4777 26801 4811
rect 26835 4777 26847 4811
rect 26789 4771 26847 4777
rect 25455 4712 26280 4740
rect 25455 4709 25467 4712
rect 25409 4703 25467 4709
rect 26418 4700 26424 4752
rect 26476 4700 26482 4752
rect 24305 4675 24363 4681
rect 24305 4672 24317 4675
rect 23952 4644 24317 4672
rect 23753 4635 23811 4641
rect 24305 4641 24317 4644
rect 24351 4641 24363 4675
rect 24305 4635 24363 4641
rect 25133 4675 25191 4681
rect 25133 4641 25145 4675
rect 25179 4641 25191 4675
rect 25501 4675 25559 4681
rect 25501 4672 25513 4675
rect 25133 4635 25191 4641
rect 25424 4644 25513 4672
rect 25424 4613 25452 4644
rect 25501 4641 25513 4644
rect 25547 4672 25559 4675
rect 25590 4672 25596 4684
rect 25547 4644 25596 4672
rect 25547 4641 25559 4644
rect 25501 4635 25559 4641
rect 25590 4632 25596 4644
rect 25648 4632 25654 4684
rect 25685 4675 25743 4681
rect 25685 4641 25697 4675
rect 25731 4672 25743 4675
rect 25774 4672 25780 4684
rect 25731 4644 25780 4672
rect 25731 4641 25743 4644
rect 25685 4635 25743 4641
rect 25774 4632 25780 4644
rect 25832 4632 25838 4684
rect 25961 4675 26019 4681
rect 25961 4641 25973 4675
rect 26007 4672 26019 4675
rect 26050 4672 26056 4684
rect 26007 4644 26056 4672
rect 26007 4641 26019 4644
rect 25961 4635 26019 4641
rect 24029 4607 24087 4613
rect 24029 4573 24041 4607
rect 24075 4573 24087 4607
rect 24029 4567 24087 4573
rect 25409 4607 25467 4613
rect 25409 4573 25421 4607
rect 25455 4573 25467 4607
rect 25409 4567 25467 4573
rect 21637 4499 21695 4505
rect 22066 4508 23336 4536
rect 22066 4468 22094 4508
rect 21560 4440 22094 4468
rect 22189 4471 22247 4477
rect 21453 4431 21511 4437
rect 22189 4437 22201 4471
rect 22235 4468 22247 4471
rect 22278 4468 22284 4480
rect 22235 4440 22284 4468
rect 22235 4437 22247 4440
rect 22189 4431 22247 4437
rect 22278 4428 22284 4440
rect 22336 4428 22342 4480
rect 22462 4428 22468 4480
rect 22520 4428 22526 4480
rect 23106 4428 23112 4480
rect 23164 4428 23170 4480
rect 24044 4468 24072 4567
rect 25225 4539 25283 4545
rect 25225 4505 25237 4539
rect 25271 4536 25283 4539
rect 25498 4536 25504 4548
rect 25271 4508 25504 4536
rect 25271 4505 25283 4508
rect 25225 4499 25283 4505
rect 25498 4496 25504 4508
rect 25556 4536 25562 4548
rect 25976 4536 26004 4635
rect 26050 4632 26056 4644
rect 26108 4632 26114 4684
rect 26804 4672 26832 4771
rect 27065 4675 27123 4681
rect 27065 4672 27077 4675
rect 26804 4644 27077 4672
rect 27065 4641 27077 4644
rect 27111 4641 27123 4675
rect 27065 4635 27123 4641
rect 26786 4564 26792 4616
rect 26844 4564 26850 4616
rect 25556 4508 26004 4536
rect 25556 4496 25562 4508
rect 24302 4468 24308 4480
rect 24044 4440 24308 4468
rect 24302 4428 24308 4440
rect 24360 4428 24366 4480
rect 26605 4471 26663 4477
rect 26605 4437 26617 4471
rect 26651 4468 26663 4471
rect 26804 4468 26832 4564
rect 26651 4440 26832 4468
rect 26651 4437 26663 4440
rect 26605 4431 26663 4437
rect 26878 4428 26884 4480
rect 26936 4428 26942 4480
rect 552 4378 27416 4400
rect 552 4326 3756 4378
rect 3808 4326 3820 4378
rect 3872 4326 3884 4378
rect 3936 4326 3948 4378
rect 4000 4326 4012 4378
rect 4064 4326 10472 4378
rect 10524 4326 10536 4378
rect 10588 4326 10600 4378
rect 10652 4326 10664 4378
rect 10716 4326 10728 4378
rect 10780 4326 17188 4378
rect 17240 4326 17252 4378
rect 17304 4326 17316 4378
rect 17368 4326 17380 4378
rect 17432 4326 17444 4378
rect 17496 4326 23904 4378
rect 23956 4326 23968 4378
rect 24020 4326 24032 4378
rect 24084 4326 24096 4378
rect 24148 4326 24160 4378
rect 24212 4326 27416 4378
rect 552 4304 27416 4326
rect 4246 4264 4252 4276
rect 3528 4236 4252 4264
rect 3050 4156 3056 4208
rect 3108 4196 3114 4208
rect 3418 4196 3424 4208
rect 3108 4168 3424 4196
rect 3108 4156 3114 4168
rect 3418 4156 3424 4168
rect 3476 4196 3482 4208
rect 3528 4205 3556 4236
rect 4246 4224 4252 4236
rect 4304 4224 4310 4276
rect 4430 4224 4436 4276
rect 4488 4224 4494 4276
rect 4617 4267 4675 4273
rect 4617 4233 4629 4267
rect 4663 4264 4675 4267
rect 4890 4264 4896 4276
rect 4663 4236 4896 4264
rect 4663 4233 4675 4236
rect 4617 4227 4675 4233
rect 4890 4224 4896 4236
rect 4948 4224 4954 4276
rect 6273 4267 6331 4273
rect 6273 4233 6285 4267
rect 6319 4233 6331 4267
rect 6273 4227 6331 4233
rect 3513 4199 3571 4205
rect 3513 4196 3525 4199
rect 3476 4168 3525 4196
rect 3476 4156 3482 4168
rect 3513 4165 3525 4168
rect 3559 4165 3571 4199
rect 4448 4196 4476 4224
rect 4982 4196 4988 4208
rect 3513 4159 3571 4165
rect 3620 4168 4988 4196
rect 3237 4131 3295 4137
rect 3237 4097 3249 4131
rect 3283 4128 3295 4131
rect 3326 4128 3332 4140
rect 3283 4100 3332 4128
rect 3283 4097 3295 4100
rect 3237 4091 3295 4097
rect 3326 4088 3332 4100
rect 3384 4128 3390 4140
rect 3620 4128 3648 4168
rect 4982 4156 4988 4168
rect 5040 4156 5046 4208
rect 6288 4196 6316 4227
rect 6362 4224 6368 4276
rect 6420 4264 6426 4276
rect 6549 4267 6607 4273
rect 6549 4264 6561 4267
rect 6420 4236 6561 4264
rect 6420 4224 6426 4236
rect 6549 4233 6561 4236
rect 6595 4233 6607 4267
rect 6549 4227 6607 4233
rect 8018 4224 8024 4276
rect 8076 4224 8082 4276
rect 8478 4224 8484 4276
rect 8536 4264 8542 4276
rect 8573 4267 8631 4273
rect 8573 4264 8585 4267
rect 8536 4236 8585 4264
rect 8536 4224 8542 4236
rect 8573 4233 8585 4236
rect 8619 4233 8631 4267
rect 8573 4227 8631 4233
rect 8941 4267 8999 4273
rect 8941 4233 8953 4267
rect 8987 4264 8999 4267
rect 9122 4264 9128 4276
rect 8987 4236 9128 4264
rect 8987 4233 8999 4236
rect 8941 4227 8999 4233
rect 9122 4224 9128 4236
rect 9180 4224 9186 4276
rect 13078 4224 13084 4276
rect 13136 4224 13142 4276
rect 17497 4267 17555 4273
rect 17497 4233 17509 4267
rect 17543 4264 17555 4267
rect 17678 4264 17684 4276
rect 17543 4236 17684 4264
rect 17543 4233 17555 4236
rect 17497 4227 17555 4233
rect 17678 4224 17684 4236
rect 17736 4264 17742 4276
rect 18049 4267 18107 4273
rect 18049 4264 18061 4267
rect 17736 4236 18061 4264
rect 17736 4224 17742 4236
rect 18049 4233 18061 4236
rect 18095 4233 18107 4267
rect 18049 4227 18107 4233
rect 18417 4267 18475 4273
rect 18417 4233 18429 4267
rect 18463 4264 18475 4267
rect 18877 4267 18935 4273
rect 18877 4264 18889 4267
rect 18463 4236 18889 4264
rect 18463 4233 18475 4236
rect 18417 4227 18475 4233
rect 18877 4233 18889 4236
rect 18923 4233 18935 4267
rect 18877 4227 18935 4233
rect 19334 4224 19340 4276
rect 19392 4224 19398 4276
rect 22554 4264 22560 4276
rect 21284 4236 22560 4264
rect 6454 4196 6460 4208
rect 6288 4168 6460 4196
rect 6454 4156 6460 4168
rect 6512 4156 6518 4208
rect 10689 4199 10747 4205
rect 10689 4165 10701 4199
rect 10735 4196 10747 4199
rect 10870 4196 10876 4208
rect 10735 4168 10876 4196
rect 10735 4165 10747 4168
rect 10689 4159 10747 4165
rect 10870 4156 10876 4168
rect 10928 4196 10934 4208
rect 15010 4196 15016 4208
rect 10928 4168 15016 4196
rect 10928 4156 10934 4168
rect 15010 4156 15016 4168
rect 15068 4156 15074 4208
rect 18230 4156 18236 4208
rect 18288 4156 18294 4208
rect 20441 4199 20499 4205
rect 20441 4165 20453 4199
rect 20487 4196 20499 4199
rect 21174 4196 21180 4208
rect 20487 4168 21180 4196
rect 20487 4165 20499 4168
rect 20441 4159 20499 4165
rect 3384 4100 3648 4128
rect 3697 4131 3755 4137
rect 3384 4088 3390 4100
rect 3697 4097 3709 4131
rect 3743 4128 3755 4131
rect 6181 4131 6239 4137
rect 6181 4128 6193 4131
rect 3743 4100 6193 4128
rect 3743 4097 3755 4100
rect 3697 4091 3755 4097
rect 2041 4063 2099 4069
rect 2041 4029 2053 4063
rect 2087 4060 2099 4063
rect 2222 4060 2228 4072
rect 2087 4032 2228 4060
rect 2087 4029 2099 4032
rect 2041 4023 2099 4029
rect 2222 4020 2228 4032
rect 2280 4060 2286 4072
rect 2409 4063 2467 4069
rect 2409 4060 2421 4063
rect 2280 4032 2421 4060
rect 2280 4020 2286 4032
rect 2409 4029 2421 4032
rect 2455 4029 2467 4063
rect 2409 4023 2467 4029
rect 2590 4020 2596 4072
rect 2648 4020 2654 4072
rect 3510 4020 3516 4072
rect 3568 4060 3574 4072
rect 3988 4069 4016 4100
rect 3789 4063 3847 4069
rect 3789 4060 3801 4063
rect 3568 4032 3801 4060
rect 3568 4020 3574 4032
rect 3789 4029 3801 4032
rect 3835 4029 3847 4063
rect 3789 4023 3847 4029
rect 3973 4063 4031 4069
rect 3973 4029 3985 4063
rect 4019 4029 4031 4063
rect 3973 4023 4031 4029
rect 4154 4020 4160 4072
rect 4212 4060 4218 4072
rect 4212 4032 4384 4060
rect 4212 4020 4218 4032
rect 4356 4004 4384 4032
rect 4798 4020 4804 4072
rect 4856 4020 4862 4072
rect 4890 4020 4896 4072
rect 4948 4060 4954 4072
rect 5368 4069 5396 4100
rect 6181 4097 6193 4100
rect 6227 4097 6239 4131
rect 10962 4128 10968 4140
rect 6181 4091 6239 4097
rect 10612 4100 10968 4128
rect 10612 4072 10640 4100
rect 10962 4088 10968 4100
rect 11020 4088 11026 4140
rect 17589 4131 17647 4137
rect 17589 4128 17601 4131
rect 17328 4100 17601 4128
rect 5077 4063 5135 4069
rect 5077 4060 5089 4063
rect 4948 4032 5089 4060
rect 4948 4020 4954 4032
rect 5077 4029 5089 4032
rect 5123 4029 5135 4063
rect 5077 4023 5135 4029
rect 5353 4063 5411 4069
rect 5353 4029 5365 4063
rect 5399 4029 5411 4063
rect 5353 4023 5411 4029
rect 5442 4020 5448 4072
rect 5500 4060 5506 4072
rect 5629 4063 5687 4069
rect 5629 4060 5641 4063
rect 5500 4032 5641 4060
rect 5500 4020 5506 4032
rect 5629 4029 5641 4032
rect 5675 4060 5687 4063
rect 5810 4060 5816 4072
rect 5675 4032 5816 4060
rect 5675 4029 5687 4032
rect 5629 4023 5687 4029
rect 5810 4020 5816 4032
rect 5868 4020 5874 4072
rect 6365 4063 6423 4069
rect 6365 4060 6377 4063
rect 5920 4032 6377 4060
rect 2314 3952 2320 4004
rect 2372 3992 2378 4004
rect 2774 3992 2780 4004
rect 2372 3964 2780 3992
rect 2372 3952 2378 3964
rect 2774 3952 2780 3964
rect 2832 3992 2838 4004
rect 4062 3992 4068 4004
rect 2832 3964 4068 3992
rect 2832 3952 2838 3964
rect 4062 3952 4068 3964
rect 4120 3952 4126 4004
rect 4246 3952 4252 4004
rect 4304 3952 4310 4004
rect 4338 3952 4344 4004
rect 4396 3992 4402 4004
rect 4449 3995 4507 4001
rect 4449 3992 4461 3995
rect 4396 3964 4461 3992
rect 4396 3952 4402 3964
rect 4449 3961 4461 3964
rect 4495 3961 4507 3995
rect 5920 3992 5948 4032
rect 6365 4029 6377 4032
rect 6411 4029 6423 4063
rect 6365 4023 6423 4029
rect 6730 4020 6736 4072
rect 6788 4020 6794 4072
rect 7006 4020 7012 4072
rect 7064 4020 7070 4072
rect 7285 4063 7343 4069
rect 7285 4029 7297 4063
rect 7331 4029 7343 4063
rect 7285 4023 7343 4029
rect 4449 3955 4507 3961
rect 4540 3964 5948 3992
rect 6089 3995 6147 4001
rect 2130 3884 2136 3936
rect 2188 3924 2194 3936
rect 4540 3924 4568 3964
rect 6089 3961 6101 3995
rect 6135 3992 6147 3995
rect 6178 3992 6184 4004
rect 6135 3964 6184 3992
rect 6135 3961 6147 3964
rect 6089 3955 6147 3961
rect 6178 3952 6184 3964
rect 6236 3952 6242 4004
rect 7300 3992 7328 4023
rect 8570 4020 8576 4072
rect 8628 4020 8634 4072
rect 8757 4063 8815 4069
rect 8757 4029 8769 4063
rect 8803 4060 8815 4063
rect 8846 4060 8852 4072
rect 8803 4032 8852 4060
rect 8803 4029 8815 4032
rect 8757 4023 8815 4029
rect 8846 4020 8852 4032
rect 8904 4060 8910 4072
rect 9122 4060 9128 4072
rect 8904 4032 9128 4060
rect 8904 4020 8910 4032
rect 9122 4020 9128 4032
rect 9180 4020 9186 4072
rect 9674 4020 9680 4072
rect 9732 4060 9738 4072
rect 10238 4063 10296 4069
rect 10238 4060 10250 4063
rect 9732 4032 10250 4060
rect 9732 4020 9738 4032
rect 10238 4029 10250 4032
rect 10284 4029 10296 4063
rect 10238 4023 10296 4029
rect 10505 4063 10563 4069
rect 10505 4029 10517 4063
rect 10551 4029 10563 4063
rect 10505 4023 10563 4029
rect 6932 3964 7328 3992
rect 2188 3896 4568 3924
rect 2188 3884 2194 3896
rect 4890 3884 4896 3936
rect 4948 3884 4954 3936
rect 5258 3884 5264 3936
rect 5316 3884 5322 3936
rect 5442 3884 5448 3936
rect 5500 3884 5506 3936
rect 5813 3927 5871 3933
rect 5813 3893 5825 3927
rect 5859 3924 5871 3927
rect 5994 3924 6000 3936
rect 5859 3896 6000 3924
rect 5859 3893 5871 3896
rect 5813 3887 5871 3893
rect 5994 3884 6000 3896
rect 6052 3924 6058 3936
rect 6638 3924 6644 3936
rect 6052 3896 6644 3924
rect 6052 3884 6058 3896
rect 6638 3884 6644 3896
rect 6696 3884 6702 3936
rect 6932 3933 6960 3964
rect 9950 3952 9956 4004
rect 10008 3992 10014 4004
rect 10318 3992 10324 4004
rect 10008 3964 10324 3992
rect 10008 3952 10014 3964
rect 10318 3952 10324 3964
rect 10376 3992 10382 4004
rect 10520 3992 10548 4023
rect 10594 4020 10600 4072
rect 10652 4020 10658 4072
rect 11701 4063 11759 4069
rect 11701 4029 11713 4063
rect 11747 4060 11759 4063
rect 11790 4060 11796 4072
rect 11747 4032 11796 4060
rect 11747 4029 11759 4032
rect 11701 4023 11759 4029
rect 11790 4020 11796 4032
rect 11848 4020 11854 4072
rect 11885 4063 11943 4069
rect 11885 4029 11897 4063
rect 11931 4060 11943 4063
rect 12066 4060 12072 4072
rect 11931 4032 12072 4060
rect 11931 4029 11943 4032
rect 11885 4023 11943 4029
rect 12066 4020 12072 4032
rect 12124 4020 12130 4072
rect 13354 4060 13360 4072
rect 12912 4032 13360 4060
rect 10376 3964 10548 3992
rect 11808 3992 11836 4020
rect 12912 4001 12940 4032
rect 13354 4020 13360 4032
rect 13412 4020 13418 4072
rect 13446 4020 13452 4072
rect 13504 4060 13510 4072
rect 13541 4063 13599 4069
rect 13541 4060 13553 4063
rect 13504 4032 13553 4060
rect 13504 4020 13510 4032
rect 13541 4029 13553 4032
rect 13587 4029 13599 4063
rect 13541 4023 13599 4029
rect 13909 4063 13967 4069
rect 13909 4029 13921 4063
rect 13955 4029 13967 4063
rect 13909 4023 13967 4029
rect 13170 4001 13176 4004
rect 12897 3995 12955 4001
rect 12897 3992 12909 3995
rect 11808 3964 12909 3992
rect 10376 3952 10382 3964
rect 12897 3961 12909 3964
rect 12943 3961 12955 3995
rect 12897 3955 12955 3961
rect 13113 3995 13176 4001
rect 13113 3961 13125 3995
rect 13159 3961 13176 3995
rect 13113 3955 13176 3961
rect 13170 3952 13176 3955
rect 13228 3952 13234 4004
rect 13924 3992 13952 4023
rect 15286 4020 15292 4072
rect 15344 4020 15350 4072
rect 15562 4020 15568 4072
rect 15620 4020 15626 4072
rect 16025 4063 16083 4069
rect 16025 4029 16037 4063
rect 16071 4060 16083 4063
rect 16117 4063 16175 4069
rect 16117 4060 16129 4063
rect 16071 4032 16129 4060
rect 16071 4029 16083 4032
rect 16025 4023 16083 4029
rect 16117 4029 16129 4032
rect 16163 4029 16175 4063
rect 16117 4023 16175 4029
rect 16393 4063 16451 4069
rect 16393 4029 16405 4063
rect 16439 4029 16451 4063
rect 16393 4023 16451 4029
rect 16408 3992 16436 4023
rect 16574 4020 16580 4072
rect 16632 4020 16638 4072
rect 17328 4069 17356 4100
rect 17589 4097 17601 4100
rect 17635 4097 17647 4131
rect 18248 4128 18276 4156
rect 20456 4128 20484 4159
rect 21174 4156 21180 4168
rect 21232 4156 21238 4208
rect 17589 4091 17647 4097
rect 17788 4100 18276 4128
rect 19720 4100 20484 4128
rect 20533 4131 20591 4137
rect 17788 4069 17816 4100
rect 17313 4063 17371 4069
rect 17313 4060 17325 4063
rect 17144 4032 17325 4060
rect 13280 3964 13952 3992
rect 15488 3964 16436 3992
rect 6917 3927 6975 3933
rect 6917 3893 6929 3927
rect 6963 3893 6975 3927
rect 6917 3887 6975 3893
rect 8294 3884 8300 3936
rect 8352 3924 8358 3936
rect 9125 3927 9183 3933
rect 9125 3924 9137 3927
rect 8352 3896 9137 3924
rect 8352 3884 8358 3896
rect 9125 3893 9137 3896
rect 9171 3893 9183 3927
rect 9125 3887 9183 3893
rect 11054 3884 11060 3936
rect 11112 3924 11118 3936
rect 11793 3927 11851 3933
rect 11793 3924 11805 3927
rect 11112 3896 11805 3924
rect 11112 3884 11118 3896
rect 11793 3893 11805 3896
rect 11839 3924 11851 3927
rect 12986 3924 12992 3936
rect 11839 3896 12992 3924
rect 11839 3893 11851 3896
rect 11793 3887 11851 3893
rect 12986 3884 12992 3896
rect 13044 3884 13050 3936
rect 13280 3933 13308 3964
rect 13265 3927 13323 3933
rect 13265 3893 13277 3927
rect 13311 3893 13323 3927
rect 13265 3887 13323 3893
rect 13630 3884 13636 3936
rect 13688 3884 13694 3936
rect 14093 3927 14151 3933
rect 14093 3893 14105 3927
rect 14139 3924 14151 3927
rect 15378 3924 15384 3936
rect 14139 3896 15384 3924
rect 14139 3893 14151 3896
rect 14093 3887 14151 3893
rect 15378 3884 15384 3896
rect 15436 3884 15442 3936
rect 15488 3933 15516 3964
rect 15473 3927 15531 3933
rect 15473 3893 15485 3927
rect 15519 3893 15531 3927
rect 15473 3887 15531 3893
rect 15749 3927 15807 3933
rect 15749 3893 15761 3927
rect 15795 3924 15807 3927
rect 16592 3924 16620 4020
rect 17144 3933 17172 4032
rect 17313 4029 17325 4032
rect 17359 4029 17371 4063
rect 17313 4023 17371 4029
rect 17497 4063 17555 4069
rect 17497 4029 17509 4063
rect 17543 4060 17555 4063
rect 17773 4063 17831 4069
rect 17773 4060 17785 4063
rect 17543 4032 17785 4060
rect 17543 4029 17555 4032
rect 17497 4023 17555 4029
rect 17773 4029 17785 4032
rect 17819 4029 17831 4063
rect 17773 4023 17831 4029
rect 17862 4020 17868 4072
rect 17920 4060 17926 4072
rect 19720 4069 19748 4100
rect 20533 4097 20545 4131
rect 20579 4128 20591 4131
rect 21284 4128 21312 4236
rect 22554 4224 22560 4236
rect 22612 4224 22618 4276
rect 22922 4224 22928 4276
rect 22980 4224 22986 4276
rect 23198 4224 23204 4276
rect 23256 4224 23262 4276
rect 25409 4267 25467 4273
rect 25409 4233 25421 4267
rect 25455 4264 25467 4267
rect 25498 4264 25504 4276
rect 25455 4236 25504 4264
rect 25455 4233 25467 4236
rect 25409 4227 25467 4233
rect 25498 4224 25504 4236
rect 25556 4224 25562 4276
rect 26326 4224 26332 4276
rect 26384 4264 26390 4276
rect 26384 4236 27108 4264
rect 26384 4224 26390 4236
rect 21358 4156 21364 4208
rect 21416 4196 21422 4208
rect 22278 4196 22284 4208
rect 21416 4168 21496 4196
rect 21416 4156 21422 4168
rect 20579 4100 21312 4128
rect 20579 4097 20591 4100
rect 20533 4091 20591 4097
rect 18049 4063 18107 4069
rect 18049 4060 18061 4063
rect 17920 4032 18061 4060
rect 17920 4020 17926 4032
rect 18049 4029 18061 4032
rect 18095 4029 18107 4063
rect 18049 4023 18107 4029
rect 18141 4063 18199 4069
rect 18141 4029 18153 4063
rect 18187 4029 18199 4063
rect 19153 4063 19211 4069
rect 19153 4060 19165 4063
rect 18141 4023 18199 4029
rect 19076 4032 19165 4060
rect 17586 3952 17592 4004
rect 17644 3992 17650 4004
rect 18156 3992 18184 4023
rect 17644 3964 18184 3992
rect 17644 3952 17650 3964
rect 18690 3952 18696 4004
rect 18748 3952 18754 4004
rect 15795 3896 16620 3924
rect 17129 3927 17187 3933
rect 15795 3893 15807 3896
rect 15749 3887 15807 3893
rect 17129 3893 17141 3927
rect 17175 3893 17187 3927
rect 17129 3887 17187 3893
rect 17862 3884 17868 3936
rect 17920 3924 17926 3936
rect 17957 3927 18015 3933
rect 17957 3924 17969 3927
rect 17920 3896 17969 3924
rect 17920 3884 17926 3896
rect 17957 3893 17969 3896
rect 18003 3893 18015 3927
rect 17957 3887 18015 3893
rect 18046 3884 18052 3936
rect 18104 3924 18110 3936
rect 19076 3933 19104 4032
rect 19153 4029 19165 4032
rect 19199 4029 19211 4063
rect 19153 4023 19211 4029
rect 19705 4063 19763 4069
rect 19705 4029 19717 4063
rect 19751 4029 19763 4063
rect 19705 4023 19763 4029
rect 19889 4063 19947 4069
rect 19889 4029 19901 4063
rect 19935 4060 19947 4063
rect 19978 4060 19984 4072
rect 19935 4032 19984 4060
rect 19935 4029 19947 4032
rect 19889 4023 19947 4029
rect 19978 4020 19984 4032
rect 20036 4060 20042 4072
rect 20073 4063 20131 4069
rect 20073 4060 20085 4063
rect 20036 4032 20085 4060
rect 20036 4020 20042 4032
rect 20073 4029 20085 4032
rect 20119 4029 20131 4063
rect 20073 4023 20131 4029
rect 20254 4020 20260 4072
rect 20312 4060 20318 4072
rect 20824 4069 20852 4100
rect 20625 4063 20683 4069
rect 20625 4060 20637 4063
rect 20312 4032 20637 4060
rect 20312 4020 20318 4032
rect 20625 4029 20637 4032
rect 20671 4029 20683 4063
rect 20625 4023 20683 4029
rect 20809 4063 20867 4069
rect 20809 4029 20821 4063
rect 20855 4029 20867 4063
rect 20809 4023 20867 4029
rect 20898 4020 20904 4072
rect 20956 4020 20962 4072
rect 21174 4020 21180 4072
rect 21232 4060 21238 4072
rect 21468 4069 21496 4168
rect 22112 4168 22284 4196
rect 21637 4131 21695 4137
rect 21637 4097 21649 4131
rect 21683 4128 21695 4131
rect 21683 4100 22048 4128
rect 21683 4097 21695 4100
rect 21637 4091 21695 4097
rect 21299 4063 21357 4069
rect 21299 4060 21311 4063
rect 21232 4032 21311 4060
rect 21232 4020 21238 4032
rect 21299 4029 21311 4032
rect 21345 4029 21357 4063
rect 21299 4023 21357 4029
rect 21453 4063 21511 4069
rect 21453 4029 21465 4063
rect 21499 4029 21511 4063
rect 21453 4023 21511 4029
rect 21545 4063 21603 4069
rect 21545 4029 21557 4063
rect 21591 4029 21603 4063
rect 21545 4023 21603 4029
rect 21729 4063 21787 4069
rect 21729 4029 21741 4063
rect 21775 4029 21787 4063
rect 21729 4023 21787 4029
rect 21560 3992 21588 4023
rect 21192 3964 21588 3992
rect 21192 3936 21220 3964
rect 18893 3927 18951 3933
rect 18893 3924 18905 3927
rect 18104 3896 18905 3924
rect 18104 3884 18110 3896
rect 18893 3893 18905 3896
rect 18939 3893 18951 3927
rect 18893 3887 18951 3893
rect 19061 3927 19119 3933
rect 19061 3893 19073 3927
rect 19107 3893 19119 3927
rect 19061 3887 19119 3893
rect 19794 3884 19800 3936
rect 19852 3884 19858 3936
rect 21085 3927 21143 3933
rect 21085 3893 21097 3927
rect 21131 3924 21143 3927
rect 21174 3924 21180 3936
rect 21131 3896 21180 3924
rect 21131 3893 21143 3896
rect 21085 3887 21143 3893
rect 21174 3884 21180 3896
rect 21232 3884 21238 3936
rect 21450 3884 21456 3936
rect 21508 3924 21514 3936
rect 21744 3924 21772 4023
rect 21818 4020 21824 4072
rect 21876 4020 21882 4072
rect 22020 4004 22048 4100
rect 22112 4069 22140 4168
rect 22278 4156 22284 4168
rect 22336 4196 22342 4208
rect 22646 4196 22652 4208
rect 22336 4168 22652 4196
rect 22336 4156 22342 4168
rect 22646 4156 22652 4168
rect 22704 4156 22710 4208
rect 23109 4131 23167 4137
rect 23109 4128 23121 4131
rect 22388 4100 23121 4128
rect 22097 4063 22155 4069
rect 22097 4029 22109 4063
rect 22143 4029 22155 4063
rect 22388 4060 22416 4100
rect 23109 4097 23121 4100
rect 23155 4097 23167 4131
rect 23109 4091 23167 4097
rect 23750 4088 23756 4140
rect 23808 4128 23814 4140
rect 23937 4131 23995 4137
rect 23937 4128 23949 4131
rect 23808 4100 23949 4128
rect 23808 4088 23814 4100
rect 23937 4097 23949 4100
rect 23983 4097 23995 4131
rect 23937 4091 23995 4097
rect 22097 4023 22155 4029
rect 22204 4032 22416 4060
rect 22465 4063 22523 4069
rect 22002 3952 22008 4004
rect 22060 3992 22066 4004
rect 22204 3992 22232 4032
rect 22465 4029 22477 4063
rect 22511 4060 22523 4063
rect 22554 4060 22560 4072
rect 22511 4032 22560 4060
rect 22511 4029 22523 4032
rect 22465 4023 22523 4029
rect 22554 4020 22560 4032
rect 22612 4020 22618 4072
rect 22646 4020 22652 4072
rect 22704 4060 22710 4072
rect 22741 4063 22799 4069
rect 22741 4060 22753 4063
rect 22704 4032 22753 4060
rect 22704 4020 22710 4032
rect 22741 4029 22753 4032
rect 22787 4029 22799 4063
rect 22741 4023 22799 4029
rect 23290 4020 23296 4072
rect 23348 4020 23354 4072
rect 24210 4020 24216 4072
rect 24268 4020 24274 4072
rect 27080 4069 27108 4236
rect 25041 4063 25099 4069
rect 25041 4060 25053 4063
rect 24964 4032 25053 4060
rect 22060 3964 22232 3992
rect 22281 3995 22339 4001
rect 22060 3952 22066 3964
rect 22281 3961 22293 3995
rect 22327 3992 22339 3995
rect 23017 3995 23075 4001
rect 23017 3992 23029 3995
rect 22327 3964 23029 3992
rect 22327 3961 22339 3964
rect 22281 3955 22339 3961
rect 23017 3961 23029 3964
rect 23063 3961 23075 3995
rect 23017 3955 23075 3961
rect 24964 3936 24992 4032
rect 25041 4029 25053 4032
rect 25087 4029 25099 4063
rect 25041 4023 25099 4029
rect 25225 4063 25283 4069
rect 25225 4029 25237 4063
rect 25271 4060 25283 4063
rect 26798 4063 26856 4069
rect 25271 4032 25728 4060
rect 25271 4029 25283 4032
rect 25225 4023 25283 4029
rect 25700 3936 25728 4032
rect 26798 4029 26810 4063
rect 26844 4029 26856 4063
rect 26798 4023 26856 4029
rect 27065 4063 27123 4069
rect 27065 4029 27077 4063
rect 27111 4029 27123 4063
rect 27065 4023 27123 4029
rect 26804 3992 26832 4023
rect 26878 3992 26884 4004
rect 26804 3964 26884 3992
rect 26878 3952 26884 3964
rect 26936 3952 26942 4004
rect 21508 3896 21772 3924
rect 21508 3884 21514 3896
rect 21818 3884 21824 3936
rect 21876 3924 21882 3936
rect 21913 3927 21971 3933
rect 21913 3924 21925 3927
rect 21876 3896 21925 3924
rect 21876 3884 21882 3896
rect 21913 3893 21925 3896
rect 21959 3893 21971 3927
rect 21913 3887 21971 3893
rect 22554 3884 22560 3936
rect 22612 3884 22618 3936
rect 23474 3884 23480 3936
rect 23532 3884 23538 3936
rect 24946 3884 24952 3936
rect 25004 3884 25010 3936
rect 25682 3884 25688 3936
rect 25740 3884 25746 3936
rect 552 3834 27576 3856
rect 552 3782 7114 3834
rect 7166 3782 7178 3834
rect 7230 3782 7242 3834
rect 7294 3782 7306 3834
rect 7358 3782 7370 3834
rect 7422 3782 13830 3834
rect 13882 3782 13894 3834
rect 13946 3782 13958 3834
rect 14010 3782 14022 3834
rect 14074 3782 14086 3834
rect 14138 3782 20546 3834
rect 20598 3782 20610 3834
rect 20662 3782 20674 3834
rect 20726 3782 20738 3834
rect 20790 3782 20802 3834
rect 20854 3782 27262 3834
rect 27314 3782 27326 3834
rect 27378 3782 27390 3834
rect 27442 3782 27454 3834
rect 27506 3782 27518 3834
rect 27570 3782 27576 3834
rect 552 3760 27576 3782
rect 2958 3720 2964 3732
rect 2746 3692 2964 3720
rect 2038 3408 2044 3460
rect 2096 3448 2102 3460
rect 2746 3448 2774 3692
rect 2958 3680 2964 3692
rect 3016 3680 3022 3732
rect 3050 3680 3056 3732
rect 3108 3720 3114 3732
rect 3108 3692 4936 3720
rect 3108 3680 3114 3692
rect 3697 3655 3755 3661
rect 2976 3624 3372 3652
rect 2976 3593 3004 3624
rect 3344 3596 3372 3624
rect 3697 3621 3709 3655
rect 3743 3652 3755 3655
rect 4908 3652 4936 3692
rect 5074 3680 5080 3732
rect 5132 3680 5138 3732
rect 6549 3723 6607 3729
rect 6549 3689 6561 3723
rect 6595 3720 6607 3723
rect 6730 3720 6736 3732
rect 6595 3692 6736 3720
rect 6595 3689 6607 3692
rect 6549 3683 6607 3689
rect 6730 3680 6736 3692
rect 6788 3680 6794 3732
rect 9766 3680 9772 3732
rect 9824 3720 9830 3732
rect 10689 3723 10747 3729
rect 10689 3720 10701 3723
rect 9824 3692 10701 3720
rect 9824 3680 9830 3692
rect 10689 3689 10701 3692
rect 10735 3720 10747 3723
rect 10778 3720 10784 3732
rect 10735 3692 10784 3720
rect 10735 3689 10747 3692
rect 10689 3683 10747 3689
rect 10778 3680 10784 3692
rect 10836 3680 10842 3732
rect 12066 3720 12072 3732
rect 11716 3692 12072 3720
rect 11716 3661 11744 3692
rect 12066 3680 12072 3692
rect 12124 3680 12130 3732
rect 12802 3680 12808 3732
rect 12860 3680 12866 3732
rect 12986 3680 12992 3732
rect 13044 3720 13050 3732
rect 13633 3723 13691 3729
rect 13633 3720 13645 3723
rect 13044 3692 13645 3720
rect 13044 3680 13050 3692
rect 13633 3689 13645 3692
rect 13679 3720 13691 3723
rect 13722 3720 13728 3732
rect 13679 3692 13728 3720
rect 13679 3689 13691 3692
rect 13633 3683 13691 3689
rect 13722 3680 13728 3692
rect 13780 3680 13786 3732
rect 14918 3680 14924 3732
rect 14976 3720 14982 3732
rect 14976 3692 15240 3720
rect 14976 3680 14982 3692
rect 5261 3655 5319 3661
rect 5261 3652 5273 3655
rect 3743 3624 4568 3652
rect 3743 3621 3755 3624
rect 3697 3615 3755 3621
rect 4540 3596 4568 3624
rect 4908 3624 5273 3652
rect 2961 3587 3019 3593
rect 2961 3553 2973 3587
rect 3007 3553 3019 3587
rect 2961 3547 3019 3553
rect 3145 3587 3203 3593
rect 3145 3553 3157 3587
rect 3191 3553 3203 3587
rect 3145 3547 3203 3553
rect 3160 3516 3188 3547
rect 3326 3544 3332 3596
rect 3384 3544 3390 3596
rect 3418 3544 3424 3596
rect 3476 3584 3482 3596
rect 4065 3587 4123 3593
rect 4065 3584 4077 3587
rect 3476 3556 3521 3584
rect 3988 3556 4077 3584
rect 3476 3544 3482 3556
rect 3436 3516 3464 3544
rect 3160 3488 3464 3516
rect 2096 3420 2774 3448
rect 2096 3408 2102 3420
rect 3234 3408 3240 3460
rect 3292 3448 3298 3460
rect 3988 3448 4016 3556
rect 4065 3553 4077 3556
rect 4111 3553 4123 3587
rect 4065 3547 4123 3553
rect 4154 3544 4160 3596
rect 4212 3584 4218 3596
rect 4249 3587 4307 3593
rect 4249 3584 4261 3587
rect 4212 3556 4261 3584
rect 4212 3544 4218 3556
rect 4249 3553 4261 3556
rect 4295 3553 4307 3587
rect 4249 3547 4307 3553
rect 4264 3516 4292 3547
rect 4338 3544 4344 3596
rect 4396 3544 4402 3596
rect 4522 3544 4528 3596
rect 4580 3544 4586 3596
rect 4706 3544 4712 3596
rect 4764 3544 4770 3596
rect 4908 3593 4936 3624
rect 5261 3621 5273 3624
rect 5307 3621 5319 3655
rect 11701 3655 11759 3661
rect 11701 3652 11713 3655
rect 5261 3615 5319 3621
rect 5368 3624 6868 3652
rect 4893 3587 4951 3593
rect 4893 3553 4905 3587
rect 4939 3553 4951 3587
rect 4893 3547 4951 3553
rect 5169 3587 5227 3593
rect 5169 3553 5181 3587
rect 5215 3584 5227 3587
rect 5368 3584 5396 3624
rect 6840 3596 6868 3624
rect 8680 3624 9352 3652
rect 5215 3556 5396 3584
rect 5445 3587 5503 3593
rect 5215 3553 5227 3556
rect 5169 3547 5227 3553
rect 5445 3553 5457 3587
rect 5491 3553 5503 3587
rect 5445 3547 5503 3553
rect 5629 3587 5687 3593
rect 5629 3553 5641 3587
rect 5675 3584 5687 3587
rect 6089 3587 6147 3593
rect 6089 3584 6101 3587
rect 5675 3556 6101 3584
rect 5675 3553 5687 3556
rect 5629 3547 5687 3553
rect 6089 3553 6101 3556
rect 6135 3553 6147 3587
rect 6089 3547 6147 3553
rect 6365 3587 6423 3593
rect 6365 3553 6377 3587
rect 6411 3553 6423 3587
rect 6365 3547 6423 3553
rect 4430 3516 4436 3528
rect 4264 3488 4436 3516
rect 4430 3476 4436 3488
rect 4488 3516 4494 3528
rect 5184 3516 5212 3547
rect 4488 3488 5212 3516
rect 5460 3516 5488 3547
rect 5810 3516 5816 3528
rect 5460 3488 5816 3516
rect 4488 3476 4494 3488
rect 5810 3476 5816 3488
rect 5868 3476 5874 3528
rect 6181 3519 6239 3525
rect 6181 3516 6193 3519
rect 5920 3488 6193 3516
rect 3292 3420 4016 3448
rect 4525 3451 4583 3457
rect 3292 3408 3298 3420
rect 4525 3417 4537 3451
rect 4571 3448 4583 3451
rect 5920 3448 5948 3488
rect 6181 3485 6193 3488
rect 6227 3485 6239 3519
rect 6181 3479 6239 3485
rect 6270 3476 6276 3528
rect 6328 3516 6334 3528
rect 6380 3516 6408 3547
rect 6638 3544 6644 3596
rect 6696 3544 6702 3596
rect 6822 3544 6828 3596
rect 6880 3544 6886 3596
rect 7101 3587 7159 3593
rect 7101 3584 7113 3587
rect 7024 3556 7113 3584
rect 6733 3519 6791 3525
rect 6733 3516 6745 3519
rect 6328 3488 6745 3516
rect 6328 3476 6334 3488
rect 6733 3485 6745 3488
rect 6779 3485 6791 3519
rect 6733 3479 6791 3485
rect 7024 3457 7052 3556
rect 7101 3553 7113 3556
rect 7147 3553 7159 3587
rect 7101 3547 7159 3553
rect 8570 3544 8576 3596
rect 8628 3584 8634 3596
rect 8680 3593 8708 3624
rect 9324 3593 9352 3624
rect 11624 3624 11713 3652
rect 8665 3587 8723 3593
rect 8665 3584 8677 3587
rect 8628 3556 8677 3584
rect 8628 3544 8634 3556
rect 8665 3553 8677 3556
rect 8711 3553 8723 3587
rect 8665 3547 8723 3553
rect 8849 3587 8907 3593
rect 8849 3553 8861 3587
rect 8895 3584 8907 3587
rect 9125 3587 9183 3593
rect 9125 3584 9137 3587
rect 8895 3556 9137 3584
rect 8895 3553 8907 3556
rect 8849 3547 8907 3553
rect 9125 3553 9137 3556
rect 9171 3553 9183 3587
rect 9125 3547 9183 3553
rect 9309 3587 9367 3593
rect 9309 3553 9321 3587
rect 9355 3553 9367 3587
rect 9309 3547 9367 3553
rect 8202 3476 8208 3528
rect 8260 3516 8266 3528
rect 8864 3516 8892 3547
rect 10226 3544 10232 3596
rect 10284 3584 10290 3596
rect 10594 3584 10600 3596
rect 10284 3556 10600 3584
rect 10284 3544 10290 3556
rect 10594 3544 10600 3556
rect 10652 3544 10658 3596
rect 11624 3593 11652 3624
rect 11701 3621 11713 3624
rect 11747 3621 11759 3655
rect 12820 3652 12848 3680
rect 12820 3624 13124 3652
rect 11701 3615 11759 3621
rect 10781 3587 10839 3593
rect 10781 3553 10793 3587
rect 10827 3553 10839 3587
rect 10781 3547 10839 3553
rect 11516 3587 11574 3593
rect 11516 3553 11528 3587
rect 11562 3553 11574 3587
rect 11516 3547 11574 3553
rect 11609 3587 11667 3593
rect 11609 3553 11621 3587
rect 11655 3553 11667 3587
rect 11609 3547 11667 3553
rect 12437 3587 12495 3593
rect 12437 3553 12449 3587
rect 12483 3553 12495 3587
rect 12437 3547 12495 3553
rect 8260 3488 8892 3516
rect 10796 3516 10824 3547
rect 11330 3516 11336 3528
rect 10796 3488 11336 3516
rect 8260 3476 8266 3488
rect 11330 3476 11336 3488
rect 11388 3476 11394 3528
rect 11532 3516 11560 3547
rect 12161 3519 12219 3525
rect 11532 3488 11836 3516
rect 11808 3460 11836 3488
rect 12161 3485 12173 3519
rect 12207 3516 12219 3519
rect 12452 3516 12480 3547
rect 12526 3544 12532 3596
rect 12584 3584 12590 3596
rect 13096 3593 13124 3624
rect 13262 3612 13268 3664
rect 13320 3612 13326 3664
rect 13538 3612 13544 3664
rect 13596 3615 13602 3664
rect 14001 3655 14059 3661
rect 14001 3621 14013 3655
rect 14047 3652 14059 3655
rect 15013 3655 15071 3661
rect 15013 3652 15025 3655
rect 14047 3624 15025 3652
rect 14047 3621 14059 3624
rect 14001 3615 14059 3621
rect 15013 3621 15025 3624
rect 15059 3621 15071 3655
rect 15212 3652 15240 3692
rect 15286 3680 15292 3732
rect 15344 3720 15350 3732
rect 15473 3723 15531 3729
rect 15473 3720 15485 3723
rect 15344 3692 15485 3720
rect 15344 3680 15350 3692
rect 15473 3689 15485 3692
rect 15519 3689 15531 3723
rect 15473 3683 15531 3689
rect 17678 3680 17684 3732
rect 17736 3680 17742 3732
rect 18046 3680 18052 3732
rect 18104 3680 18110 3732
rect 19334 3680 19340 3732
rect 19392 3720 19398 3732
rect 19702 3720 19708 3732
rect 19392 3692 19708 3720
rect 19392 3680 19398 3692
rect 19702 3680 19708 3692
rect 19760 3680 19766 3732
rect 19794 3680 19800 3732
rect 19852 3680 19858 3732
rect 21818 3680 21824 3732
rect 21876 3680 21882 3732
rect 21910 3680 21916 3732
rect 21968 3720 21974 3732
rect 22554 3720 22560 3732
rect 21968 3692 22560 3720
rect 21968 3680 21974 3692
rect 22554 3680 22560 3692
rect 22612 3680 22618 3732
rect 22922 3680 22928 3732
rect 22980 3680 22986 3732
rect 23290 3680 23296 3732
rect 23348 3680 23354 3732
rect 23474 3680 23480 3732
rect 23532 3680 23538 3732
rect 23845 3723 23903 3729
rect 23845 3689 23857 3723
rect 23891 3720 23903 3723
rect 24210 3720 24216 3732
rect 23891 3692 24216 3720
rect 23891 3689 23903 3692
rect 23845 3683 23903 3689
rect 24210 3680 24216 3692
rect 24268 3680 24274 3732
rect 24946 3680 24952 3732
rect 25004 3680 25010 3732
rect 25682 3680 25688 3732
rect 25740 3680 25746 3732
rect 15212 3624 16160 3652
rect 15013 3615 15071 3621
rect 13596 3612 13615 3615
rect 13557 3609 13615 3612
rect 12897 3587 12955 3593
rect 12897 3584 12909 3587
rect 12584 3556 12909 3584
rect 12584 3544 12590 3556
rect 12897 3553 12909 3556
rect 12943 3553 12955 3587
rect 12897 3547 12955 3553
rect 13081 3587 13139 3593
rect 13081 3553 13093 3587
rect 13127 3553 13139 3587
rect 13081 3547 13139 3553
rect 13170 3544 13176 3596
rect 13228 3544 13234 3596
rect 13354 3544 13360 3596
rect 13412 3544 13418 3596
rect 13557 3575 13569 3609
rect 13603 3575 13615 3609
rect 13557 3569 13615 3575
rect 13817 3587 13875 3593
rect 13817 3553 13829 3587
rect 13863 3584 13875 3587
rect 13863 3556 14228 3584
rect 13863 3553 13875 3556
rect 13817 3547 13875 3553
rect 12621 3519 12679 3525
rect 12207 3488 12572 3516
rect 12207 3485 12219 3488
rect 12161 3479 12219 3485
rect 4571 3420 5948 3448
rect 7009 3451 7067 3457
rect 4571 3417 4583 3420
rect 4525 3411 4583 3417
rect 4157 3383 4215 3389
rect 4157 3349 4169 3383
rect 4203 3380 4215 3383
rect 4430 3380 4436 3392
rect 4203 3352 4436 3380
rect 4203 3349 4215 3352
rect 4157 3343 4215 3349
rect 4430 3340 4436 3352
rect 4488 3340 4494 3392
rect 4908 3389 4936 3420
rect 7009 3417 7021 3451
rect 7055 3417 7067 3451
rect 7009 3411 7067 3417
rect 7116 3420 11560 3448
rect 4893 3383 4951 3389
rect 4893 3349 4905 3383
rect 4939 3349 4951 3383
rect 4893 3343 4951 3349
rect 6362 3340 6368 3392
rect 6420 3340 6426 3392
rect 6454 3340 6460 3392
rect 6512 3380 6518 3392
rect 6641 3383 6699 3389
rect 6641 3380 6653 3383
rect 6512 3352 6653 3380
rect 6512 3340 6518 3352
rect 6641 3349 6653 3352
rect 6687 3349 6699 3383
rect 6641 3343 6699 3349
rect 6914 3340 6920 3392
rect 6972 3380 6978 3392
rect 7116 3380 7144 3420
rect 6972 3352 7144 3380
rect 7285 3383 7343 3389
rect 6972 3340 6978 3352
rect 7285 3349 7297 3383
rect 7331 3380 7343 3383
rect 7374 3380 7380 3392
rect 7331 3352 7380 3380
rect 7331 3349 7343 3352
rect 7285 3343 7343 3349
rect 7374 3340 7380 3352
rect 7432 3340 7438 3392
rect 7466 3340 7472 3392
rect 7524 3340 7530 3392
rect 8846 3340 8852 3392
rect 8904 3380 8910 3392
rect 9033 3383 9091 3389
rect 9033 3380 9045 3383
rect 8904 3352 9045 3380
rect 8904 3340 8910 3352
rect 9033 3349 9045 3352
rect 9079 3349 9091 3383
rect 9033 3343 9091 3349
rect 9122 3340 9128 3392
rect 9180 3380 9186 3392
rect 9217 3383 9275 3389
rect 9217 3380 9229 3383
rect 9180 3352 9229 3380
rect 9180 3340 9186 3352
rect 9217 3349 9229 3352
rect 9263 3349 9275 3383
rect 9217 3343 9275 3349
rect 11422 3340 11428 3392
rect 11480 3340 11486 3392
rect 11532 3380 11560 3420
rect 11790 3408 11796 3460
rect 11848 3448 11854 3460
rect 11977 3451 12035 3457
rect 11977 3448 11989 3451
rect 11848 3420 11989 3448
rect 11848 3408 11854 3420
rect 11977 3417 11989 3420
rect 12023 3417 12035 3451
rect 12544 3448 12572 3488
rect 12621 3485 12633 3519
rect 12667 3516 12679 3519
rect 12802 3516 12808 3528
rect 12667 3488 12808 3516
rect 12667 3485 12679 3488
rect 12621 3479 12679 3485
rect 12802 3476 12808 3488
rect 12860 3476 12866 3528
rect 12989 3519 13047 3525
rect 12989 3485 13001 3519
rect 13035 3516 13047 3519
rect 13906 3516 13912 3528
rect 13035 3488 13912 3516
rect 13035 3485 13047 3488
rect 12989 3479 13047 3485
rect 13906 3476 13912 3488
rect 13964 3476 13970 3528
rect 14200 3516 14228 3556
rect 14366 3544 14372 3596
rect 14424 3584 14430 3596
rect 14461 3587 14519 3593
rect 14461 3584 14473 3587
rect 14424 3556 14473 3584
rect 14424 3544 14430 3556
rect 14461 3553 14473 3556
rect 14507 3553 14519 3587
rect 14461 3547 14519 3553
rect 14550 3544 14556 3596
rect 14608 3544 14614 3596
rect 14737 3587 14795 3593
rect 14737 3553 14749 3587
rect 14783 3584 14795 3587
rect 14826 3584 14832 3596
rect 14783 3556 14832 3584
rect 14783 3553 14795 3556
rect 14737 3547 14795 3553
rect 14274 3516 14280 3528
rect 14200 3488 14280 3516
rect 14274 3476 14280 3488
rect 14332 3516 14338 3528
rect 14752 3516 14780 3547
rect 14826 3544 14832 3556
rect 14884 3544 14890 3596
rect 15289 3587 15347 3593
rect 15289 3553 15301 3587
rect 15335 3553 15347 3587
rect 15289 3547 15347 3553
rect 14332 3488 14780 3516
rect 14332 3476 14338 3488
rect 14918 3476 14924 3528
rect 14976 3516 14982 3528
rect 15105 3519 15163 3525
rect 15105 3516 15117 3519
rect 14976 3488 15117 3516
rect 14976 3476 14982 3488
rect 15105 3485 15117 3488
rect 15151 3485 15163 3519
rect 15304 3516 15332 3547
rect 15378 3544 15384 3596
rect 15436 3584 15442 3596
rect 15565 3587 15623 3593
rect 15565 3584 15577 3587
rect 15436 3556 15577 3584
rect 15436 3544 15442 3556
rect 15565 3553 15577 3556
rect 15611 3584 15623 3587
rect 15654 3584 15660 3596
rect 15611 3556 15660 3584
rect 15611 3553 15623 3556
rect 15565 3547 15623 3553
rect 15654 3544 15660 3556
rect 15712 3544 15718 3596
rect 15746 3544 15752 3596
rect 15804 3544 15810 3596
rect 16132 3593 16160 3624
rect 16117 3587 16175 3593
rect 16117 3553 16129 3587
rect 16163 3553 16175 3587
rect 17696 3584 17724 3680
rect 19812 3652 19840 3680
rect 21836 3652 21864 3680
rect 19812 3624 22232 3652
rect 17773 3587 17831 3593
rect 17773 3584 17785 3587
rect 17696 3556 17785 3584
rect 16117 3547 16175 3553
rect 17773 3553 17785 3556
rect 17819 3553 17831 3587
rect 17773 3547 17831 3553
rect 17862 3544 17868 3596
rect 17920 3544 17926 3596
rect 19521 3587 19579 3593
rect 19521 3553 19533 3587
rect 19567 3553 19579 3587
rect 19521 3547 19579 3553
rect 19705 3587 19763 3593
rect 19705 3553 19717 3587
rect 19751 3584 19763 3587
rect 19812 3584 19840 3624
rect 19751 3556 19840 3584
rect 19751 3553 19763 3556
rect 19705 3547 19763 3553
rect 15933 3519 15991 3525
rect 15933 3516 15945 3519
rect 15304 3488 15945 3516
rect 15105 3479 15163 3485
rect 15933 3485 15945 3488
rect 15979 3516 15991 3519
rect 16209 3519 16267 3525
rect 16209 3516 16221 3519
rect 15979 3488 16221 3516
rect 15979 3485 15991 3488
rect 15933 3479 15991 3485
rect 16209 3485 16221 3488
rect 16255 3485 16267 3519
rect 16209 3479 16267 3485
rect 17586 3476 17592 3528
rect 17644 3516 17650 3528
rect 18049 3519 18107 3525
rect 18049 3516 18061 3519
rect 17644 3488 18061 3516
rect 17644 3476 17650 3488
rect 18049 3485 18061 3488
rect 18095 3485 18107 3519
rect 19536 3516 19564 3547
rect 20162 3544 20168 3596
rect 20220 3544 20226 3596
rect 21266 3544 21272 3596
rect 21324 3584 21330 3596
rect 21361 3587 21419 3593
rect 21361 3584 21373 3587
rect 21324 3556 21373 3584
rect 21324 3544 21330 3556
rect 21361 3553 21373 3556
rect 21407 3553 21419 3587
rect 21361 3547 21419 3553
rect 21450 3544 21456 3596
rect 21508 3584 21514 3596
rect 21545 3587 21603 3593
rect 21545 3584 21557 3587
rect 21508 3556 21557 3584
rect 21508 3544 21514 3556
rect 21545 3553 21557 3556
rect 21591 3553 21603 3587
rect 21545 3547 21603 3553
rect 21637 3587 21695 3593
rect 21637 3553 21649 3587
rect 21683 3553 21695 3587
rect 21821 3587 21879 3593
rect 21821 3584 21833 3587
rect 21637 3547 21695 3553
rect 21744 3556 21833 3584
rect 20180 3516 20208 3544
rect 19536 3488 20208 3516
rect 18049 3479 18107 3485
rect 21082 3476 21088 3528
rect 21140 3516 21146 3528
rect 21652 3516 21680 3547
rect 21744 3528 21772 3556
rect 21821 3553 21833 3556
rect 21867 3553 21879 3587
rect 21821 3547 21879 3553
rect 22094 3544 22100 3596
rect 22152 3544 22158 3596
rect 22204 3593 22232 3624
rect 22189 3587 22247 3593
rect 22189 3553 22201 3587
rect 22235 3553 22247 3587
rect 22189 3547 22247 3553
rect 22462 3544 22468 3596
rect 22520 3584 22526 3596
rect 22649 3587 22707 3593
rect 22649 3584 22661 3587
rect 22520 3556 22661 3584
rect 22520 3544 22526 3556
rect 22649 3553 22661 3556
rect 22695 3584 22707 3587
rect 22738 3584 22744 3596
rect 22695 3556 22744 3584
rect 22695 3553 22707 3556
rect 22649 3547 22707 3553
rect 22738 3544 22744 3556
rect 22796 3544 22802 3596
rect 22833 3587 22891 3593
rect 22833 3553 22845 3587
rect 22879 3553 22891 3587
rect 22940 3584 22968 3680
rect 23017 3655 23075 3661
rect 23017 3621 23029 3655
rect 23063 3652 23075 3655
rect 23308 3652 23336 3680
rect 23063 3624 23336 3652
rect 23063 3621 23075 3624
rect 23017 3615 23075 3621
rect 23308 3593 23336 3624
rect 23109 3587 23167 3593
rect 23109 3584 23121 3587
rect 22940 3556 23121 3584
rect 22833 3547 22891 3553
rect 23109 3553 23121 3556
rect 23155 3553 23167 3587
rect 23109 3547 23167 3553
rect 23293 3587 23351 3593
rect 23293 3553 23305 3587
rect 23339 3553 23351 3587
rect 23492 3584 23520 3680
rect 23661 3587 23719 3593
rect 23661 3584 23673 3587
rect 23492 3556 23673 3584
rect 23293 3547 23351 3553
rect 23661 3553 23673 3556
rect 23707 3553 23719 3587
rect 23661 3547 23719 3553
rect 23937 3587 23995 3593
rect 23937 3553 23949 3587
rect 23983 3553 23995 3587
rect 24964 3584 24992 3680
rect 25409 3587 25467 3593
rect 25409 3584 25421 3587
rect 24964 3556 25421 3584
rect 23937 3547 23995 3553
rect 25409 3553 25421 3556
rect 25455 3553 25467 3587
rect 25409 3547 25467 3553
rect 25593 3587 25651 3593
rect 25593 3553 25605 3587
rect 25639 3584 25651 3587
rect 25700 3584 25728 3680
rect 25639 3556 25728 3584
rect 25639 3553 25651 3556
rect 25593 3547 25651 3553
rect 21140 3488 21680 3516
rect 21140 3476 21146 3488
rect 21726 3476 21732 3528
rect 21784 3476 21790 3528
rect 14366 3448 14372 3460
rect 11977 3411 12035 3417
rect 12084 3420 12434 3448
rect 12544 3420 14372 3448
rect 12084 3380 12112 3420
rect 11532 3352 12112 3380
rect 12250 3340 12256 3392
rect 12308 3340 12314 3392
rect 12406 3380 12434 3420
rect 14366 3408 14372 3420
rect 14424 3408 14430 3460
rect 15120 3420 17080 3448
rect 15120 3392 15148 3420
rect 17052 3392 17080 3420
rect 19518 3408 19524 3460
rect 19576 3448 19582 3460
rect 22848 3448 22876 3547
rect 23014 3476 23020 3528
rect 23072 3476 23078 3528
rect 23952 3516 23980 3547
rect 25501 3519 25559 3525
rect 23492 3488 23980 3516
rect 24044 3488 25452 3516
rect 19576 3420 22876 3448
rect 19576 3408 19582 3420
rect 14458 3380 14464 3392
rect 12406 3352 14464 3380
rect 14458 3340 14464 3352
rect 14516 3340 14522 3392
rect 15102 3340 15108 3392
rect 15160 3340 15166 3392
rect 15470 3340 15476 3392
rect 15528 3380 15534 3392
rect 16117 3383 16175 3389
rect 16117 3380 16129 3383
rect 15528 3352 16129 3380
rect 15528 3340 15534 3352
rect 16117 3349 16129 3352
rect 16163 3349 16175 3383
rect 16117 3343 16175 3349
rect 16482 3340 16488 3392
rect 16540 3340 16546 3392
rect 17034 3340 17040 3392
rect 17092 3340 17098 3392
rect 17678 3340 17684 3392
rect 17736 3380 17742 3392
rect 19426 3380 19432 3392
rect 17736 3352 19432 3380
rect 17736 3340 17742 3352
rect 19426 3340 19432 3352
rect 19484 3340 19490 3392
rect 19613 3383 19671 3389
rect 19613 3349 19625 3383
rect 19659 3380 19671 3383
rect 19702 3380 19708 3392
rect 19659 3352 19708 3380
rect 19659 3349 19671 3352
rect 19613 3343 19671 3349
rect 19702 3340 19708 3352
rect 19760 3340 19766 3392
rect 21450 3340 21456 3392
rect 21508 3340 21514 3392
rect 21729 3383 21787 3389
rect 21729 3349 21741 3383
rect 21775 3380 21787 3383
rect 21818 3380 21824 3392
rect 21775 3352 21824 3380
rect 21775 3349 21787 3352
rect 21729 3343 21787 3349
rect 21818 3340 21824 3352
rect 21876 3340 21882 3392
rect 22002 3340 22008 3392
rect 22060 3380 22066 3392
rect 22097 3383 22155 3389
rect 22097 3380 22109 3383
rect 22060 3352 22109 3380
rect 22060 3340 22066 3352
rect 22097 3349 22109 3352
rect 22143 3349 22155 3383
rect 22097 3343 22155 3349
rect 22465 3383 22523 3389
rect 22465 3349 22477 3383
rect 22511 3380 22523 3383
rect 23032 3380 23060 3476
rect 23492 3457 23520 3488
rect 23477 3451 23535 3457
rect 23477 3417 23489 3451
rect 23523 3417 23535 3451
rect 24044 3448 24072 3488
rect 23477 3411 23535 3417
rect 23768 3420 24072 3448
rect 24121 3451 24179 3457
rect 23768 3392 23796 3420
rect 24121 3417 24133 3451
rect 24167 3448 24179 3451
rect 24302 3448 24308 3460
rect 24167 3420 24308 3448
rect 24167 3417 24179 3420
rect 24121 3411 24179 3417
rect 24302 3408 24308 3420
rect 24360 3408 24366 3460
rect 25424 3448 25452 3488
rect 25501 3485 25513 3519
rect 25547 3516 25559 3519
rect 25774 3516 25780 3528
rect 25547 3488 25780 3516
rect 25547 3485 25559 3488
rect 25501 3479 25559 3485
rect 25774 3476 25780 3488
rect 25832 3476 25838 3528
rect 25682 3448 25688 3460
rect 25424 3420 25688 3448
rect 25682 3408 25688 3420
rect 25740 3448 25746 3460
rect 26418 3448 26424 3460
rect 25740 3420 26424 3448
rect 25740 3408 25746 3420
rect 26418 3408 26424 3420
rect 26476 3408 26482 3460
rect 22511 3352 23060 3380
rect 22511 3349 22523 3352
rect 22465 3343 22523 3349
rect 23106 3340 23112 3392
rect 23164 3340 23170 3392
rect 23750 3340 23756 3392
rect 23808 3340 23814 3392
rect 24213 3383 24271 3389
rect 24213 3349 24225 3383
rect 24259 3380 24271 3383
rect 24578 3380 24584 3392
rect 24259 3352 24584 3380
rect 24259 3349 24271 3352
rect 24213 3343 24271 3349
rect 24578 3340 24584 3352
rect 24636 3340 24642 3392
rect 552 3290 27416 3312
rect 552 3238 3756 3290
rect 3808 3238 3820 3290
rect 3872 3238 3884 3290
rect 3936 3238 3948 3290
rect 4000 3238 4012 3290
rect 4064 3238 10472 3290
rect 10524 3238 10536 3290
rect 10588 3238 10600 3290
rect 10652 3238 10664 3290
rect 10716 3238 10728 3290
rect 10780 3238 17188 3290
rect 17240 3238 17252 3290
rect 17304 3238 17316 3290
rect 17368 3238 17380 3290
rect 17432 3238 17444 3290
rect 17496 3238 23904 3290
rect 23956 3238 23968 3290
rect 24020 3238 24032 3290
rect 24084 3238 24096 3290
rect 24148 3238 24160 3290
rect 24212 3238 27416 3290
rect 552 3216 27416 3238
rect 2222 3136 2228 3188
rect 2280 3136 2286 3188
rect 5997 3179 6055 3185
rect 5997 3145 6009 3179
rect 6043 3176 6055 3179
rect 6270 3176 6276 3188
rect 6043 3148 6276 3176
rect 6043 3145 6055 3148
rect 5997 3139 6055 3145
rect 6270 3136 6276 3148
rect 6328 3136 6334 3188
rect 7006 3176 7012 3188
rect 6840 3148 7012 3176
rect 2240 3040 2268 3136
rect 1872 3012 2268 3040
rect 1872 2981 1900 3012
rect 1673 2975 1731 2981
rect 1673 2941 1685 2975
rect 1719 2941 1731 2975
rect 1673 2935 1731 2941
rect 1857 2975 1915 2981
rect 1857 2941 1869 2975
rect 1903 2941 1915 2975
rect 1857 2935 1915 2941
rect 1949 2975 2007 2981
rect 1949 2941 1961 2975
rect 1995 2972 2007 2975
rect 2038 2972 2044 2984
rect 1995 2944 2044 2972
rect 1995 2941 2007 2944
rect 1949 2935 2007 2941
rect 1688 2904 1716 2935
rect 1964 2904 1992 2935
rect 2038 2932 2044 2944
rect 2096 2932 2102 2984
rect 2240 2981 2268 3012
rect 2424 3080 3280 3108
rect 2424 2984 2452 3080
rect 2774 3000 2780 3052
rect 2832 3000 2838 3052
rect 3050 3040 3056 3052
rect 2884 3012 3056 3040
rect 2133 2975 2191 2981
rect 2133 2941 2145 2975
rect 2179 2941 2191 2975
rect 2133 2935 2191 2941
rect 2225 2975 2283 2981
rect 2225 2941 2237 2975
rect 2271 2941 2283 2975
rect 2225 2935 2283 2941
rect 1688 2876 1992 2904
rect 1302 2796 1308 2848
rect 1360 2836 1366 2848
rect 1765 2839 1823 2845
rect 1765 2836 1777 2839
rect 1360 2808 1777 2836
rect 1360 2796 1366 2808
rect 1765 2805 1777 2808
rect 1811 2805 1823 2839
rect 1765 2799 1823 2805
rect 2038 2796 2044 2848
rect 2096 2796 2102 2848
rect 2148 2836 2176 2935
rect 2406 2932 2412 2984
rect 2464 2932 2470 2984
rect 2685 2975 2743 2981
rect 2685 2941 2697 2975
rect 2731 2972 2743 2975
rect 2792 2972 2820 3000
rect 2884 2981 2912 3012
rect 3050 3000 3056 3012
rect 3108 3000 3114 3052
rect 3252 2984 3280 3080
rect 5258 3068 5264 3120
rect 5316 3108 5322 3120
rect 6840 3108 6868 3148
rect 7006 3136 7012 3148
rect 7064 3136 7070 3188
rect 7466 3176 7472 3188
rect 7208 3148 7472 3176
rect 5316 3080 6868 3108
rect 5316 3068 5322 3080
rect 6914 3068 6920 3120
rect 6972 3068 6978 3120
rect 3786 3000 3792 3052
rect 3844 3040 3850 3052
rect 6932 3040 6960 3068
rect 7208 3049 7236 3148
rect 7466 3136 7472 3148
rect 7524 3136 7530 3188
rect 8202 3136 8208 3188
rect 8260 3136 8266 3188
rect 8570 3136 8576 3188
rect 8628 3136 8634 3188
rect 10226 3136 10232 3188
rect 10284 3136 10290 3188
rect 10612 3148 10824 3176
rect 10244 3108 10272 3136
rect 10244 3080 10456 3108
rect 3844 3012 6224 3040
rect 3844 3000 3850 3012
rect 2731 2944 2820 2972
rect 2869 2975 2927 2981
rect 2731 2941 2743 2944
rect 2685 2935 2743 2941
rect 2869 2941 2881 2975
rect 2915 2941 2927 2975
rect 2869 2935 2927 2941
rect 3234 2932 3240 2984
rect 3292 2972 3298 2984
rect 6196 2981 6224 3012
rect 6279 3012 6960 3040
rect 7193 3043 7251 3049
rect 3421 2975 3479 2981
rect 3421 2972 3433 2975
rect 3292 2944 3433 2972
rect 3292 2932 3298 2944
rect 3421 2941 3433 2944
rect 3467 2941 3479 2975
rect 6181 2975 6239 2981
rect 3421 2935 3479 2941
rect 3528 2944 5856 2972
rect 2317 2907 2375 2913
rect 2317 2873 2329 2907
rect 2363 2904 2375 2907
rect 2498 2904 2504 2916
rect 2363 2876 2504 2904
rect 2363 2873 2375 2876
rect 2317 2867 2375 2873
rect 2498 2864 2504 2876
rect 2556 2904 2562 2916
rect 3528 2904 3556 2944
rect 2556 2876 3556 2904
rect 3605 2907 3663 2913
rect 2556 2864 2562 2876
rect 3605 2873 3617 2907
rect 3651 2904 3663 2907
rect 4338 2904 4344 2916
rect 3651 2876 4344 2904
rect 3651 2873 3663 2876
rect 3605 2867 3663 2873
rect 4338 2864 4344 2876
rect 4396 2864 4402 2916
rect 5258 2864 5264 2916
rect 5316 2904 5322 2916
rect 5828 2913 5856 2944
rect 6181 2941 6193 2975
rect 6227 2941 6239 2975
rect 6181 2935 6239 2941
rect 5629 2907 5687 2913
rect 5629 2904 5641 2907
rect 5316 2876 5641 2904
rect 5316 2864 5322 2876
rect 5629 2873 5641 2876
rect 5675 2873 5687 2907
rect 5629 2867 5687 2873
rect 5813 2907 5871 2913
rect 5813 2873 5825 2907
rect 5859 2873 5871 2907
rect 6279 2904 6307 3012
rect 6365 2975 6423 2981
rect 6365 2941 6377 2975
rect 6411 2972 6423 2975
rect 6457 2975 6515 2981
rect 6457 2972 6469 2975
rect 6411 2944 6469 2972
rect 6411 2941 6423 2944
rect 6365 2935 6423 2941
rect 6457 2941 6469 2944
rect 6503 2941 6515 2975
rect 6457 2935 6515 2941
rect 5813 2867 5871 2873
rect 5920 2876 6307 2904
rect 6472 2904 6500 2935
rect 6638 2932 6644 2984
rect 6696 2932 6702 2984
rect 6748 2981 6776 3012
rect 7193 3009 7205 3043
rect 7239 3009 7251 3043
rect 7193 3003 7251 3009
rect 9950 3000 9956 3052
rect 10008 3000 10014 3052
rect 6733 2975 6791 2981
rect 6733 2941 6745 2975
rect 6779 2941 6791 2975
rect 6733 2935 6791 2941
rect 6917 2975 6975 2981
rect 6917 2941 6929 2975
rect 6963 2941 6975 2975
rect 6917 2935 6975 2941
rect 6825 2907 6883 2913
rect 6825 2904 6837 2907
rect 6472 2876 6837 2904
rect 2682 2836 2688 2848
rect 2148 2808 2688 2836
rect 2682 2796 2688 2808
rect 2740 2836 2746 2848
rect 2777 2839 2835 2845
rect 2777 2836 2789 2839
rect 2740 2808 2789 2836
rect 2740 2796 2746 2808
rect 2777 2805 2789 2808
rect 2823 2805 2835 2839
rect 2777 2799 2835 2805
rect 4246 2796 4252 2848
rect 4304 2836 4310 2848
rect 5920 2836 5948 2876
rect 6825 2873 6837 2876
rect 6871 2873 6883 2907
rect 6932 2904 6960 2935
rect 7374 2932 7380 2984
rect 7432 2972 7438 2984
rect 10428 2981 10456 3080
rect 7469 2975 7527 2981
rect 7469 2972 7481 2975
rect 7432 2944 7481 2972
rect 7432 2932 7438 2944
rect 7469 2941 7481 2944
rect 7515 2941 7527 2975
rect 7469 2935 7527 2941
rect 10229 2975 10287 2981
rect 10229 2941 10241 2975
rect 10275 2941 10287 2975
rect 10229 2935 10287 2941
rect 10413 2975 10471 2981
rect 10413 2941 10425 2975
rect 10459 2941 10471 2975
rect 10413 2935 10471 2941
rect 10505 2975 10563 2981
rect 10505 2941 10517 2975
rect 10551 2972 10563 2975
rect 10612 2972 10640 3148
rect 10686 3068 10692 3120
rect 10744 3068 10750 3120
rect 10796 3108 10824 3148
rect 11882 3136 11888 3188
rect 11940 3176 11946 3188
rect 11940 3148 13021 3176
rect 11940 3136 11946 3148
rect 12894 3108 12900 3120
rect 10796 3080 12900 3108
rect 12894 3068 12900 3080
rect 12952 3068 12958 3120
rect 12993 3108 13021 3148
rect 13814 3136 13820 3188
rect 13872 3136 13878 3188
rect 14182 3136 14188 3188
rect 14240 3136 14246 3188
rect 14277 3179 14335 3185
rect 14277 3145 14289 3179
rect 14323 3176 14335 3179
rect 15102 3176 15108 3188
rect 14323 3148 15108 3176
rect 14323 3145 14335 3148
rect 14277 3139 14335 3145
rect 15102 3136 15108 3148
rect 15160 3136 15166 3188
rect 15470 3136 15476 3188
rect 15528 3136 15534 3188
rect 15562 3136 15568 3188
rect 15620 3176 15626 3188
rect 15657 3179 15715 3185
rect 15657 3176 15669 3179
rect 15620 3148 15669 3176
rect 15620 3136 15626 3148
rect 15657 3145 15669 3148
rect 15703 3145 15715 3179
rect 16482 3176 16488 3188
rect 15657 3139 15715 3145
rect 15948 3148 16488 3176
rect 14090 3108 14096 3120
rect 12993 3080 14096 3108
rect 14090 3068 14096 3080
rect 14148 3068 14154 3120
rect 14366 3068 14372 3120
rect 14424 3108 14430 3120
rect 14424 3080 15332 3108
rect 14424 3068 14430 3080
rect 11149 3043 11207 3049
rect 11149 3040 11161 3043
rect 10704 3012 11161 3040
rect 10704 2981 10732 3012
rect 10551 2944 10640 2972
rect 10689 2975 10747 2981
rect 10551 2941 10563 2944
rect 10505 2935 10563 2941
rect 10689 2941 10701 2975
rect 10735 2941 10747 2975
rect 10689 2935 10747 2941
rect 7190 2904 7196 2916
rect 6932 2876 7196 2904
rect 6825 2867 6883 2873
rect 7190 2864 7196 2876
rect 7248 2864 7254 2916
rect 9674 2864 9680 2916
rect 9732 2913 9738 2916
rect 9732 2867 9744 2913
rect 10244 2904 10272 2935
rect 10520 2904 10548 2935
rect 10778 2932 10784 2984
rect 10836 2932 10842 2984
rect 10888 2974 10916 3012
rect 11149 3009 11161 3012
rect 11195 3009 11207 3043
rect 11149 3003 11207 3009
rect 11716 3012 13032 3040
rect 10965 2975 11023 2981
rect 10965 2974 10977 2975
rect 10888 2946 10977 2974
rect 10965 2941 10977 2946
rect 11011 2941 11023 2975
rect 10965 2935 11023 2941
rect 11054 2932 11060 2984
rect 11112 2932 11118 2984
rect 11238 2932 11244 2984
rect 11296 2972 11302 2984
rect 11716 2981 11744 3012
rect 11701 2975 11759 2981
rect 11701 2972 11713 2975
rect 11296 2944 11713 2972
rect 11296 2932 11302 2944
rect 11701 2941 11713 2944
rect 11747 2941 11759 2975
rect 11701 2935 11759 2941
rect 12342 2932 12348 2984
rect 12400 2972 12406 2984
rect 12728 2981 12756 3012
rect 12529 2975 12587 2981
rect 12529 2972 12541 2975
rect 12400 2944 12541 2972
rect 12400 2932 12406 2944
rect 12529 2941 12541 2944
rect 12575 2941 12587 2975
rect 12529 2935 12587 2941
rect 12713 2975 12771 2981
rect 12713 2941 12725 2975
rect 12759 2941 12771 2975
rect 12713 2935 12771 2941
rect 12805 2975 12863 2981
rect 12805 2941 12817 2975
rect 12851 2972 12863 2975
rect 12894 2972 12900 2984
rect 12851 2944 12900 2972
rect 12851 2941 12863 2944
rect 12805 2935 12863 2941
rect 12894 2932 12900 2944
rect 12952 2932 12958 2984
rect 13004 2981 13032 3012
rect 13262 3000 13268 3052
rect 13320 3040 13326 3052
rect 15304 3049 15332 3080
rect 15289 3043 15347 3049
rect 13320 3012 14504 3040
rect 13320 3000 13326 3012
rect 12989 2975 13047 2981
rect 12989 2941 13001 2975
rect 13035 2972 13047 2975
rect 13538 2972 13544 2984
rect 13035 2944 13544 2972
rect 13035 2941 13047 2944
rect 12989 2935 13047 2941
rect 13538 2932 13544 2944
rect 13596 2932 13602 2984
rect 13722 2932 13728 2984
rect 13780 2932 13786 2984
rect 13814 2932 13820 2984
rect 13872 2932 13878 2984
rect 13909 2975 13967 2981
rect 13909 2941 13921 2975
rect 13955 2941 13967 2975
rect 13909 2935 13967 2941
rect 10244 2876 10548 2904
rect 9732 2864 9738 2867
rect 11330 2864 11336 2916
rect 11388 2904 11394 2916
rect 11517 2907 11575 2913
rect 11517 2904 11529 2907
rect 11388 2876 11529 2904
rect 11388 2864 11394 2876
rect 11517 2873 11529 2876
rect 11563 2904 11575 2907
rect 12360 2904 12388 2932
rect 11563 2876 12388 2904
rect 13740 2904 13768 2932
rect 13924 2904 13952 2935
rect 14274 2932 14280 2984
rect 14332 2932 14338 2984
rect 14476 2981 14504 3012
rect 15289 3009 15301 3043
rect 15335 3009 15347 3043
rect 15289 3003 15347 3009
rect 14461 2975 14519 2981
rect 14461 2941 14473 2975
rect 14507 2972 14519 2975
rect 14553 2975 14611 2981
rect 14553 2972 14565 2975
rect 14507 2944 14565 2972
rect 14507 2941 14519 2944
rect 14461 2935 14519 2941
rect 14553 2941 14565 2944
rect 14599 2941 14611 2975
rect 14553 2935 14611 2941
rect 14737 2975 14795 2981
rect 14737 2941 14749 2975
rect 14783 2941 14795 2975
rect 14737 2935 14795 2941
rect 13740 2876 13952 2904
rect 11563 2873 11575 2876
rect 11517 2867 11575 2873
rect 14182 2864 14188 2916
rect 14240 2904 14246 2916
rect 14752 2904 14780 2935
rect 15010 2932 15016 2984
rect 15068 2972 15074 2984
rect 15948 2981 15976 3148
rect 16482 3136 16488 3148
rect 16540 3136 16546 3188
rect 17586 3136 17592 3188
rect 17644 3176 17650 3188
rect 17865 3179 17923 3185
rect 17865 3176 17877 3179
rect 17644 3148 17877 3176
rect 17644 3136 17650 3148
rect 17865 3145 17877 3148
rect 17911 3176 17923 3179
rect 18233 3179 18291 3185
rect 18233 3176 18245 3179
rect 17911 3148 18245 3176
rect 17911 3145 17923 3148
rect 17865 3139 17923 3145
rect 18233 3145 18245 3148
rect 18279 3145 18291 3179
rect 18233 3139 18291 3145
rect 18690 3136 18696 3188
rect 18748 3176 18754 3188
rect 23750 3176 23756 3188
rect 18748 3148 23756 3176
rect 18748 3136 18754 3148
rect 23750 3136 23756 3148
rect 23808 3136 23814 3188
rect 24578 3176 24584 3188
rect 23952 3148 24584 3176
rect 17221 3111 17279 3117
rect 17221 3077 17233 3111
rect 17267 3077 17279 3111
rect 17221 3071 17279 3077
rect 15473 2975 15531 2981
rect 15473 2972 15485 2975
rect 15068 2944 15485 2972
rect 15068 2932 15074 2944
rect 15473 2941 15485 2944
rect 15519 2941 15531 2975
rect 15473 2935 15531 2941
rect 15933 2975 15991 2981
rect 15933 2941 15945 2975
rect 15979 2941 15991 2975
rect 15933 2935 15991 2941
rect 16206 2932 16212 2984
rect 16264 2932 16270 2984
rect 16485 2975 16543 2981
rect 16485 2941 16497 2975
rect 16531 2941 16543 2975
rect 17236 2972 17264 3071
rect 19242 3068 19248 3120
rect 19300 3068 19306 3120
rect 19334 3068 19340 3120
rect 19392 3108 19398 3120
rect 19392 3080 19472 3108
rect 19392 3068 19398 3080
rect 18138 2972 18144 2984
rect 17236 2944 18144 2972
rect 16485 2935 16543 2941
rect 14240 2876 14780 2904
rect 15197 2907 15255 2913
rect 14240 2864 14246 2876
rect 15197 2873 15209 2907
rect 15243 2904 15255 2907
rect 15838 2904 15844 2916
rect 15243 2876 15844 2904
rect 15243 2873 15255 2876
rect 15197 2867 15255 2873
rect 4304 2808 5948 2836
rect 4304 2796 4310 2808
rect 6270 2796 6276 2848
rect 6328 2796 6334 2848
rect 6362 2796 6368 2848
rect 6420 2836 6426 2848
rect 6549 2839 6607 2845
rect 6549 2836 6561 2839
rect 6420 2808 6561 2836
rect 6420 2796 6426 2808
rect 6549 2805 6561 2808
rect 6595 2836 6607 2839
rect 8294 2836 8300 2848
rect 6595 2808 8300 2836
rect 6595 2805 6607 2808
rect 6549 2799 6607 2805
rect 8294 2796 8300 2808
rect 8352 2796 8358 2848
rect 10042 2796 10048 2848
rect 10100 2836 10106 2848
rect 10321 2839 10379 2845
rect 10321 2836 10333 2839
rect 10100 2808 10333 2836
rect 10100 2796 10106 2808
rect 10321 2805 10333 2808
rect 10367 2805 10379 2839
rect 10321 2799 10379 2805
rect 10873 2839 10931 2845
rect 10873 2805 10885 2839
rect 10919 2836 10931 2839
rect 10962 2836 10968 2848
rect 10919 2808 10968 2836
rect 10919 2805 10931 2808
rect 10873 2799 10931 2805
rect 10962 2796 10968 2808
rect 11020 2796 11026 2848
rect 12710 2796 12716 2848
rect 12768 2796 12774 2848
rect 12894 2796 12900 2848
rect 12952 2796 12958 2848
rect 14645 2839 14703 2845
rect 14645 2805 14657 2839
rect 14691 2836 14703 2839
rect 15212 2836 15240 2867
rect 15838 2864 15844 2876
rect 15896 2864 15902 2916
rect 16500 2904 16528 2935
rect 18138 2932 18144 2944
rect 18196 2932 18202 2984
rect 18322 2932 18328 2984
rect 18380 2932 18386 2984
rect 19260 2981 19288 3068
rect 19444 3049 19472 3080
rect 19886 3068 19892 3120
rect 19944 3108 19950 3120
rect 21082 3108 21088 3120
rect 19944 3080 21088 3108
rect 19944 3068 19950 3080
rect 21082 3068 21088 3080
rect 21140 3068 21146 3120
rect 21450 3068 21456 3120
rect 21508 3108 21514 3120
rect 21508 3080 22508 3108
rect 21508 3068 21514 3080
rect 19429 3043 19487 3049
rect 19429 3009 19441 3043
rect 19475 3009 19487 3043
rect 19904 3040 19932 3068
rect 19429 3003 19487 3009
rect 19628 3012 19932 3040
rect 20441 3043 20499 3049
rect 19628 2981 19656 3012
rect 20441 3009 20453 3043
rect 20487 3040 20499 3043
rect 20990 3040 20996 3052
rect 20487 3012 20996 3040
rect 20487 3009 20499 3012
rect 20441 3003 20499 3009
rect 20990 3000 20996 3012
rect 21048 3000 21054 3052
rect 19061 2975 19119 2981
rect 19061 2941 19073 2975
rect 19107 2941 19119 2975
rect 19061 2935 19119 2941
rect 19245 2975 19303 2981
rect 19245 2941 19257 2975
rect 19291 2972 19303 2975
rect 19337 2975 19395 2981
rect 19337 2972 19349 2975
rect 19291 2944 19349 2972
rect 19291 2941 19303 2944
rect 19245 2935 19303 2941
rect 19337 2941 19349 2944
rect 19383 2941 19395 2975
rect 19337 2935 19395 2941
rect 19521 2975 19579 2981
rect 19521 2941 19533 2975
rect 19567 2974 19579 2975
rect 19613 2975 19671 2981
rect 19613 2974 19625 2975
rect 19567 2946 19625 2974
rect 19567 2941 19579 2946
rect 19521 2935 19579 2941
rect 19613 2941 19625 2946
rect 19659 2941 19671 2975
rect 19613 2935 19671 2941
rect 16132 2876 16528 2904
rect 18049 2907 18107 2913
rect 16132 2845 16160 2876
rect 18049 2873 18061 2907
rect 18095 2904 18107 2907
rect 18690 2904 18696 2916
rect 18095 2876 18696 2904
rect 18095 2873 18107 2876
rect 18049 2867 18107 2873
rect 18690 2864 18696 2876
rect 18748 2864 18754 2916
rect 19076 2904 19104 2935
rect 19702 2932 19708 2984
rect 19760 2972 19766 2984
rect 19797 2975 19855 2981
rect 19797 2972 19809 2975
rect 19760 2944 19809 2972
rect 19760 2932 19766 2944
rect 19797 2941 19809 2944
rect 19843 2972 19855 2975
rect 19889 2975 19947 2981
rect 19889 2972 19901 2975
rect 19843 2944 19901 2972
rect 19843 2941 19855 2944
rect 19797 2935 19855 2941
rect 19889 2941 19901 2944
rect 19935 2941 19947 2975
rect 19889 2935 19947 2941
rect 20073 2975 20131 2981
rect 20073 2941 20085 2975
rect 20119 2972 20131 2975
rect 20346 2972 20352 2984
rect 20404 2981 20410 2984
rect 21100 2981 21128 3068
rect 22094 3000 22100 3052
rect 22152 3000 22158 3052
rect 20119 2944 20352 2972
rect 20119 2941 20131 2944
rect 20073 2935 20131 2941
rect 20088 2904 20116 2935
rect 20346 2932 20352 2944
rect 20404 2972 20413 2981
rect 20533 2975 20591 2981
rect 20404 2944 20449 2972
rect 20404 2935 20413 2944
rect 20533 2941 20545 2975
rect 20579 2941 20591 2975
rect 20533 2935 20591 2941
rect 21085 2975 21143 2981
rect 21085 2941 21097 2975
rect 21131 2941 21143 2975
rect 21085 2935 21143 2941
rect 22005 2975 22063 2981
rect 22005 2941 22017 2975
rect 22051 2972 22063 2975
rect 22051 2944 22085 2972
rect 22051 2941 22063 2944
rect 22005 2935 22063 2941
rect 20404 2932 20410 2935
rect 19076 2876 20116 2904
rect 20162 2864 20168 2916
rect 20220 2904 20226 2916
rect 20548 2904 20576 2935
rect 20901 2907 20959 2913
rect 20901 2904 20913 2907
rect 20220 2876 20913 2904
rect 20220 2864 20226 2876
rect 20901 2873 20913 2876
rect 20947 2904 20959 2907
rect 21726 2904 21732 2916
rect 20947 2876 21732 2904
rect 20947 2873 20959 2876
rect 20901 2867 20959 2873
rect 21726 2864 21732 2876
rect 21784 2864 21790 2916
rect 22020 2904 22048 2935
rect 22186 2932 22192 2984
rect 22244 2932 22250 2984
rect 22480 2981 22508 3080
rect 22554 3068 22560 3120
rect 22612 3108 22618 3120
rect 22612 3080 22692 3108
rect 22612 3068 22618 3080
rect 22664 3040 22692 3080
rect 22738 3068 22744 3120
rect 22796 3108 22802 3120
rect 22796 3080 23704 3108
rect 22796 3068 22802 3080
rect 22664 3012 22784 3040
rect 22756 2981 22784 3012
rect 22281 2975 22339 2981
rect 22281 2941 22293 2975
rect 22327 2941 22339 2975
rect 22281 2935 22339 2941
rect 22465 2975 22523 2981
rect 22465 2941 22477 2975
rect 22511 2972 22523 2975
rect 22557 2975 22615 2981
rect 22557 2972 22569 2975
rect 22511 2944 22569 2972
rect 22511 2941 22523 2944
rect 22465 2935 22523 2941
rect 22557 2941 22569 2944
rect 22603 2941 22615 2975
rect 22557 2935 22615 2941
rect 22741 2975 22799 2981
rect 22741 2941 22753 2975
rect 22787 2941 22799 2975
rect 22741 2935 22799 2941
rect 22296 2904 22324 2935
rect 23382 2932 23388 2984
rect 23440 2932 23446 2984
rect 22020 2876 22324 2904
rect 22373 2907 22431 2913
rect 14691 2808 15240 2836
rect 16117 2839 16175 2845
rect 14691 2805 14703 2808
rect 14645 2799 14703 2805
rect 16117 2805 16129 2839
rect 16163 2805 16175 2839
rect 16117 2799 16175 2805
rect 17678 2796 17684 2848
rect 17736 2796 17742 2848
rect 17849 2839 17907 2845
rect 17849 2805 17861 2839
rect 17895 2836 17907 2839
rect 18138 2836 18144 2848
rect 17895 2808 18144 2836
rect 17895 2805 17907 2808
rect 17849 2799 17907 2805
rect 18138 2796 18144 2808
rect 18196 2796 18202 2848
rect 19150 2796 19156 2848
rect 19208 2796 19214 2848
rect 19702 2796 19708 2848
rect 19760 2796 19766 2848
rect 19978 2796 19984 2848
rect 20036 2796 20042 2848
rect 20714 2796 20720 2848
rect 20772 2836 20778 2848
rect 22020 2836 22048 2876
rect 22373 2873 22385 2907
rect 22419 2904 22431 2907
rect 23566 2904 23572 2916
rect 22419 2876 23572 2904
rect 22419 2873 22431 2876
rect 22373 2867 22431 2873
rect 23566 2864 23572 2876
rect 23624 2864 23630 2916
rect 23676 2904 23704 3080
rect 23952 3049 23980 3148
rect 24578 3136 24584 3148
rect 24636 3136 24642 3188
rect 25501 3179 25559 3185
rect 25501 3145 25513 3179
rect 25547 3176 25559 3179
rect 25590 3176 25596 3188
rect 25547 3148 25596 3176
rect 25547 3145 25559 3148
rect 25501 3139 25559 3145
rect 25590 3136 25596 3148
rect 25648 3176 25654 3188
rect 26329 3179 26387 3185
rect 26329 3176 26341 3179
rect 25648 3148 26341 3176
rect 25648 3136 25654 3148
rect 26329 3145 26341 3148
rect 26375 3145 26387 3179
rect 26329 3139 26387 3145
rect 24949 3111 25007 3117
rect 24949 3077 24961 3111
rect 24995 3077 25007 3111
rect 24949 3071 25007 3077
rect 23937 3043 23995 3049
rect 23937 3009 23949 3043
rect 23983 3009 23995 3043
rect 24964 3040 24992 3071
rect 24964 3012 26464 3040
rect 23937 3003 23995 3009
rect 24213 2975 24271 2981
rect 24213 2941 24225 2975
rect 24259 2972 24271 2975
rect 24302 2972 24308 2984
rect 24259 2944 24308 2972
rect 24259 2941 24271 2944
rect 24213 2935 24271 2941
rect 24302 2932 24308 2944
rect 24360 2932 24366 2984
rect 25130 2932 25136 2984
rect 25188 2932 25194 2984
rect 25976 2981 26004 3012
rect 26436 2981 26464 3012
rect 25225 2975 25283 2981
rect 25225 2941 25237 2975
rect 25271 2972 25283 2975
rect 25961 2975 26019 2981
rect 25271 2944 25360 2972
rect 25271 2941 25283 2944
rect 25225 2935 25283 2941
rect 25148 2904 25176 2932
rect 23676 2876 25176 2904
rect 20772 2808 22048 2836
rect 22649 2839 22707 2845
rect 20772 2796 20778 2808
rect 22649 2805 22661 2839
rect 22695 2836 22707 2839
rect 23198 2836 23204 2848
rect 22695 2808 23204 2836
rect 22695 2805 22707 2808
rect 22649 2799 22707 2805
rect 23198 2796 23204 2808
rect 23256 2836 23262 2848
rect 24854 2836 24860 2848
rect 23256 2808 24860 2836
rect 23256 2796 23262 2808
rect 24854 2796 24860 2808
rect 24912 2796 24918 2848
rect 25038 2796 25044 2848
rect 25096 2796 25102 2848
rect 25332 2845 25360 2944
rect 25961 2941 25973 2975
rect 26007 2941 26019 2975
rect 25961 2935 26019 2941
rect 26237 2975 26295 2981
rect 26237 2941 26249 2975
rect 26283 2941 26295 2975
rect 26237 2935 26295 2941
rect 26421 2975 26479 2981
rect 26421 2941 26433 2975
rect 26467 2941 26479 2975
rect 26421 2935 26479 2941
rect 25682 2864 25688 2916
rect 25740 2864 25746 2916
rect 26050 2864 26056 2916
rect 26108 2904 26114 2916
rect 26145 2907 26203 2913
rect 26145 2904 26157 2907
rect 26108 2876 26157 2904
rect 26108 2864 26114 2876
rect 26145 2873 26157 2876
rect 26191 2904 26203 2907
rect 26252 2904 26280 2935
rect 26191 2876 26280 2904
rect 26191 2873 26203 2876
rect 26145 2867 26203 2873
rect 25317 2839 25375 2845
rect 25317 2805 25329 2839
rect 25363 2805 25375 2839
rect 25317 2799 25375 2805
rect 25485 2839 25543 2845
rect 25485 2805 25497 2839
rect 25531 2836 25543 2839
rect 25777 2839 25835 2845
rect 25777 2836 25789 2839
rect 25531 2808 25789 2836
rect 25531 2805 25543 2808
rect 25485 2799 25543 2805
rect 25777 2805 25789 2808
rect 25823 2805 25835 2839
rect 25777 2799 25835 2805
rect 552 2746 27576 2768
rect 552 2694 7114 2746
rect 7166 2694 7178 2746
rect 7230 2694 7242 2746
rect 7294 2694 7306 2746
rect 7358 2694 7370 2746
rect 7422 2694 13830 2746
rect 13882 2694 13894 2746
rect 13946 2694 13958 2746
rect 14010 2694 14022 2746
rect 14074 2694 14086 2746
rect 14138 2694 20546 2746
rect 20598 2694 20610 2746
rect 20662 2694 20674 2746
rect 20726 2694 20738 2746
rect 20790 2694 20802 2746
rect 20854 2694 27262 2746
rect 27314 2694 27326 2746
rect 27378 2694 27390 2746
rect 27442 2694 27454 2746
rect 27506 2694 27518 2746
rect 27570 2694 27576 2746
rect 552 2672 27576 2694
rect 4706 2592 4712 2644
rect 4764 2632 4770 2644
rect 5077 2635 5135 2641
rect 5077 2632 5089 2635
rect 4764 2604 5089 2632
rect 4764 2592 4770 2604
rect 5077 2601 5089 2604
rect 5123 2601 5135 2635
rect 5077 2595 5135 2601
rect 6181 2635 6239 2641
rect 6181 2601 6193 2635
rect 6227 2632 6239 2635
rect 6454 2632 6460 2644
rect 6227 2604 6460 2632
rect 6227 2601 6239 2604
rect 6181 2595 6239 2601
rect 6454 2592 6460 2604
rect 6512 2592 6518 2644
rect 6638 2592 6644 2644
rect 6696 2632 6702 2644
rect 6733 2635 6791 2641
rect 6733 2632 6745 2635
rect 6696 2604 6745 2632
rect 6696 2592 6702 2604
rect 6733 2601 6745 2604
rect 6779 2601 6791 2635
rect 6733 2595 6791 2601
rect 8846 2592 8852 2644
rect 8904 2641 8910 2644
rect 8904 2635 8933 2641
rect 8921 2601 8933 2635
rect 8904 2595 8933 2601
rect 9033 2635 9091 2641
rect 9033 2601 9045 2635
rect 9079 2601 9091 2635
rect 9033 2595 9091 2601
rect 9309 2635 9367 2641
rect 9309 2601 9321 2635
rect 9355 2632 9367 2635
rect 9674 2632 9680 2644
rect 9355 2604 9680 2632
rect 9355 2601 9367 2604
rect 9309 2595 9367 2601
rect 8904 2592 8910 2595
rect 5997 2567 6055 2573
rect 3436 2536 4568 2564
rect 2406 2456 2412 2508
rect 2464 2496 2470 2508
rect 2501 2499 2559 2505
rect 2501 2496 2513 2499
rect 2464 2468 2513 2496
rect 2464 2456 2470 2468
rect 2501 2465 2513 2468
rect 2547 2465 2559 2499
rect 2501 2459 2559 2465
rect 2682 2456 2688 2508
rect 2740 2456 2746 2508
rect 3436 2505 3464 2536
rect 4540 2508 4568 2536
rect 5460 2536 5948 2564
rect 3421 2499 3479 2505
rect 3421 2465 3433 2499
rect 3467 2465 3479 2499
rect 3421 2459 3479 2465
rect 3605 2499 3663 2505
rect 3605 2465 3617 2499
rect 3651 2465 3663 2499
rect 3605 2459 3663 2465
rect 3620 2428 3648 2459
rect 4338 2456 4344 2508
rect 4396 2456 4402 2508
rect 4522 2456 4528 2508
rect 4580 2496 4586 2508
rect 4617 2499 4675 2505
rect 4617 2496 4629 2499
rect 4580 2468 4629 2496
rect 4580 2456 4586 2468
rect 4617 2465 4629 2468
rect 4663 2465 4675 2499
rect 4617 2459 4675 2465
rect 4801 2499 4859 2505
rect 4801 2465 4813 2499
rect 4847 2496 4859 2499
rect 4890 2496 4896 2508
rect 4847 2468 4896 2496
rect 4847 2465 4859 2468
rect 4801 2459 4859 2465
rect 4890 2456 4896 2468
rect 4948 2456 4954 2508
rect 4985 2499 5043 2505
rect 4985 2465 4997 2499
rect 5031 2465 5043 2499
rect 4985 2459 5043 2465
rect 3786 2428 3792 2440
rect 3620 2400 3792 2428
rect 3786 2388 3792 2400
rect 3844 2428 3850 2440
rect 5000 2428 5028 2459
rect 5074 2456 5080 2508
rect 5132 2496 5138 2508
rect 5169 2499 5227 2505
rect 5169 2496 5181 2499
rect 5132 2468 5181 2496
rect 5132 2456 5138 2468
rect 5169 2465 5181 2468
rect 5215 2496 5227 2499
rect 5353 2499 5411 2505
rect 5353 2496 5365 2499
rect 5215 2468 5365 2496
rect 5215 2465 5227 2468
rect 5169 2459 5227 2465
rect 5353 2465 5365 2468
rect 5399 2496 5411 2499
rect 5460 2496 5488 2536
rect 5399 2468 5488 2496
rect 5537 2499 5595 2505
rect 5399 2465 5411 2468
rect 5353 2459 5411 2465
rect 5537 2465 5549 2499
rect 5583 2496 5595 2499
rect 5626 2496 5632 2508
rect 5583 2468 5632 2496
rect 5583 2465 5595 2468
rect 5537 2459 5595 2465
rect 5626 2456 5632 2468
rect 5684 2456 5690 2508
rect 5813 2499 5871 2505
rect 5813 2465 5825 2499
rect 5859 2465 5871 2499
rect 5920 2496 5948 2536
rect 5997 2533 6009 2567
rect 6043 2564 6055 2567
rect 8665 2567 8723 2573
rect 6043 2536 6592 2564
rect 6043 2533 6055 2536
rect 5997 2527 6055 2533
rect 6273 2502 6331 2505
rect 6196 2499 6331 2502
rect 6196 2496 6285 2499
rect 5920 2474 6285 2496
rect 5920 2468 6224 2474
rect 5813 2459 5871 2465
rect 6273 2465 6285 2474
rect 6319 2465 6331 2499
rect 6273 2459 6331 2465
rect 5828 2428 5856 2459
rect 6454 2456 6460 2508
rect 6512 2456 6518 2508
rect 3844 2400 5028 2428
rect 5736 2400 5856 2428
rect 3844 2388 3850 2400
rect 2682 2320 2688 2372
rect 2740 2360 2746 2372
rect 5736 2360 5764 2400
rect 2740 2332 5764 2360
rect 6457 2363 6515 2369
rect 2740 2320 2746 2332
rect 6457 2329 6469 2363
rect 6503 2360 6515 2363
rect 6564 2360 6592 2536
rect 8665 2533 8677 2567
rect 8711 2533 8723 2567
rect 8665 2527 8723 2533
rect 6733 2499 6791 2505
rect 6733 2465 6745 2499
rect 6779 2465 6791 2499
rect 6733 2459 6791 2465
rect 6917 2499 6975 2505
rect 6917 2465 6929 2499
rect 6963 2496 6975 2499
rect 7650 2496 7656 2508
rect 6963 2468 7656 2496
rect 6963 2465 6975 2468
rect 6917 2459 6975 2465
rect 6748 2428 6776 2459
rect 7650 2456 7656 2468
rect 7708 2456 7714 2508
rect 6822 2428 6828 2440
rect 6748 2400 6828 2428
rect 6822 2388 6828 2400
rect 6880 2428 6886 2440
rect 8680 2428 8708 2527
rect 9048 2496 9076 2595
rect 9674 2592 9680 2604
rect 9732 2592 9738 2644
rect 10778 2592 10784 2644
rect 10836 2632 10842 2644
rect 11330 2632 11336 2644
rect 10836 2604 11336 2632
rect 10836 2592 10842 2604
rect 11330 2592 11336 2604
rect 11388 2592 11394 2644
rect 12710 2592 12716 2644
rect 12768 2632 12774 2644
rect 12894 2632 12900 2644
rect 12768 2604 12900 2632
rect 12768 2592 12774 2604
rect 12894 2592 12900 2604
rect 12952 2592 12958 2644
rect 13722 2592 13728 2644
rect 13780 2592 13786 2644
rect 15289 2635 15347 2641
rect 15289 2601 15301 2635
rect 15335 2632 15347 2635
rect 15470 2632 15476 2644
rect 15335 2604 15476 2632
rect 15335 2601 15347 2604
rect 15289 2595 15347 2601
rect 15470 2592 15476 2604
rect 15528 2592 15534 2644
rect 18233 2635 18291 2641
rect 18233 2601 18245 2635
rect 18279 2632 18291 2635
rect 22189 2635 22247 2641
rect 18279 2604 18368 2632
rect 18279 2601 18291 2604
rect 18233 2595 18291 2601
rect 18340 2576 18368 2604
rect 22189 2601 22201 2635
rect 22235 2601 22247 2635
rect 22189 2595 22247 2601
rect 22465 2635 22523 2641
rect 22465 2601 22477 2635
rect 22511 2632 22523 2635
rect 22830 2632 22836 2644
rect 22511 2604 22836 2632
rect 22511 2601 22523 2604
rect 22465 2595 22523 2601
rect 14645 2567 14703 2573
rect 12728 2536 13492 2564
rect 12728 2508 12756 2536
rect 9125 2499 9183 2505
rect 9125 2496 9137 2499
rect 9048 2468 9137 2496
rect 9125 2465 9137 2468
rect 9171 2465 9183 2499
rect 9125 2459 9183 2465
rect 11422 2456 11428 2508
rect 11480 2496 11486 2508
rect 11701 2499 11759 2505
rect 11701 2496 11713 2499
rect 11480 2468 11713 2496
rect 11480 2456 11486 2468
rect 11701 2465 11713 2468
rect 11747 2465 11759 2499
rect 11701 2459 11759 2465
rect 9030 2428 9036 2440
rect 6880 2400 7236 2428
rect 8680 2400 9036 2428
rect 6880 2388 6886 2400
rect 7208 2360 7236 2400
rect 9030 2388 9036 2400
rect 9088 2388 9094 2440
rect 9490 2388 9496 2440
rect 9548 2388 9554 2440
rect 11716 2428 11744 2459
rect 11882 2456 11888 2508
rect 11940 2456 11946 2508
rect 12158 2456 12164 2508
rect 12216 2456 12222 2508
rect 12526 2456 12532 2508
rect 12584 2456 12590 2508
rect 12710 2456 12716 2508
rect 12768 2456 12774 2508
rect 12805 2499 12863 2505
rect 12805 2465 12817 2499
rect 12851 2465 12863 2499
rect 12805 2459 12863 2465
rect 12544 2428 12572 2456
rect 12820 2428 12848 2459
rect 12894 2456 12900 2508
rect 12952 2496 12958 2508
rect 12989 2499 13047 2505
rect 12989 2496 13001 2499
rect 12952 2468 13001 2496
rect 12952 2456 12958 2468
rect 12989 2465 13001 2468
rect 13035 2465 13047 2499
rect 12989 2459 13047 2465
rect 11716 2400 12848 2428
rect 9508 2360 9536 2388
rect 6503 2332 7144 2360
rect 7208 2332 9536 2360
rect 6503 2329 6515 2332
rect 6457 2323 6515 2329
rect 7116 2304 7144 2332
rect 10134 2320 10140 2372
rect 10192 2360 10198 2372
rect 10962 2360 10968 2372
rect 10192 2332 10968 2360
rect 10192 2320 10198 2332
rect 10962 2320 10968 2332
rect 11020 2320 11026 2372
rect 12618 2320 12624 2372
rect 12676 2360 12682 2372
rect 12805 2363 12863 2369
rect 12805 2360 12817 2363
rect 12676 2332 12817 2360
rect 12676 2320 12682 2332
rect 12805 2329 12817 2332
rect 12851 2329 12863 2363
rect 13004 2360 13032 2459
rect 13464 2428 13492 2536
rect 13648 2536 14504 2564
rect 13648 2508 13676 2536
rect 13630 2456 13636 2508
rect 13688 2456 13694 2508
rect 13817 2499 13875 2505
rect 13817 2465 13829 2499
rect 13863 2496 13875 2499
rect 14182 2496 14188 2508
rect 13863 2468 14188 2496
rect 13863 2465 13875 2468
rect 13817 2459 13875 2465
rect 14182 2456 14188 2468
rect 14240 2456 14246 2508
rect 14274 2456 14280 2508
rect 14332 2456 14338 2508
rect 14476 2505 14504 2536
rect 14645 2533 14657 2567
rect 14691 2564 14703 2567
rect 15105 2567 15163 2573
rect 15105 2564 15117 2567
rect 14691 2536 15117 2564
rect 14691 2533 14703 2536
rect 14645 2527 14703 2533
rect 15105 2533 15117 2536
rect 15151 2564 15163 2567
rect 15378 2564 15384 2576
rect 15151 2536 15384 2564
rect 15151 2533 15163 2536
rect 15105 2527 15163 2533
rect 15378 2524 15384 2536
rect 15436 2524 15442 2576
rect 17586 2564 17592 2576
rect 16868 2536 17592 2564
rect 14461 2499 14519 2505
rect 14461 2465 14473 2499
rect 14507 2496 14519 2499
rect 14553 2499 14611 2505
rect 14553 2496 14565 2499
rect 14507 2468 14565 2496
rect 14507 2465 14519 2468
rect 14461 2459 14519 2465
rect 14553 2465 14565 2468
rect 14599 2465 14611 2499
rect 14737 2499 14795 2505
rect 14737 2496 14749 2499
rect 14553 2459 14611 2465
rect 14660 2468 14749 2496
rect 14292 2428 14320 2456
rect 13464 2400 14320 2428
rect 14660 2372 14688 2468
rect 14737 2465 14749 2468
rect 14783 2465 14795 2499
rect 14737 2459 14795 2465
rect 14921 2499 14979 2505
rect 14921 2465 14933 2499
rect 14967 2496 14979 2499
rect 15010 2496 15016 2508
rect 14967 2468 15016 2496
rect 14967 2465 14979 2468
rect 14921 2459 14979 2465
rect 15010 2456 15016 2468
rect 15068 2456 15074 2508
rect 16206 2456 16212 2508
rect 16264 2456 16270 2508
rect 16868 2505 16896 2536
rect 17586 2524 17592 2536
rect 17644 2524 17650 2576
rect 18322 2524 18328 2576
rect 18380 2524 18386 2576
rect 18509 2567 18567 2573
rect 18509 2533 18521 2567
rect 18555 2533 18567 2567
rect 20898 2564 20904 2576
rect 18509 2527 18567 2533
rect 20548 2536 20904 2564
rect 16853 2499 16911 2505
rect 16853 2465 16865 2499
rect 16899 2465 16911 2499
rect 16853 2459 16911 2465
rect 16942 2456 16948 2508
rect 17000 2496 17006 2508
rect 17109 2499 17167 2505
rect 17109 2496 17121 2499
rect 17000 2468 17121 2496
rect 17000 2456 17006 2468
rect 17109 2465 17121 2468
rect 17155 2465 17167 2499
rect 17109 2459 17167 2465
rect 18230 2456 18236 2508
rect 18288 2496 18294 2508
rect 18524 2496 18552 2527
rect 18288 2468 18552 2496
rect 18288 2456 18294 2468
rect 20254 2456 20260 2508
rect 20312 2456 20318 2508
rect 20548 2505 20576 2536
rect 20898 2524 20904 2536
rect 20956 2524 20962 2576
rect 22204 2564 22232 2595
rect 22830 2592 22836 2604
rect 22888 2592 22894 2644
rect 23106 2592 23112 2644
rect 23164 2632 23170 2644
rect 23201 2635 23259 2641
rect 23201 2632 23213 2635
rect 23164 2604 23213 2632
rect 23164 2592 23170 2604
rect 23201 2601 23213 2604
rect 23247 2601 23259 2635
rect 23201 2595 23259 2601
rect 25869 2635 25927 2641
rect 25869 2601 25881 2635
rect 25915 2632 25927 2635
rect 26050 2632 26056 2644
rect 25915 2604 26056 2632
rect 25915 2601 25927 2604
rect 25869 2595 25927 2601
rect 26050 2592 26056 2604
rect 26108 2592 26114 2644
rect 23017 2567 23075 2573
rect 23017 2564 23029 2567
rect 21008 2536 21404 2564
rect 22204 2536 23029 2564
rect 21008 2508 21036 2536
rect 20533 2499 20591 2505
rect 20533 2465 20545 2499
rect 20579 2465 20591 2499
rect 20533 2459 20591 2465
rect 20717 2499 20775 2505
rect 20717 2465 20729 2499
rect 20763 2496 20775 2499
rect 20809 2499 20867 2505
rect 20809 2496 20821 2499
rect 20763 2468 20821 2496
rect 20763 2465 20775 2468
rect 20717 2459 20775 2465
rect 20809 2465 20821 2468
rect 20855 2465 20867 2499
rect 20809 2459 20867 2465
rect 18138 2388 18144 2440
rect 18196 2428 18202 2440
rect 18693 2431 18751 2437
rect 18693 2428 18705 2431
rect 18196 2400 18705 2428
rect 18196 2388 18202 2400
rect 18693 2397 18705 2400
rect 18739 2397 18751 2431
rect 20824 2428 20852 2459
rect 20990 2456 20996 2508
rect 21048 2456 21054 2508
rect 21174 2456 21180 2508
rect 21232 2496 21238 2508
rect 21269 2499 21327 2505
rect 21269 2496 21281 2499
rect 21232 2468 21281 2496
rect 21232 2456 21238 2468
rect 21269 2465 21281 2468
rect 21315 2465 21327 2499
rect 21269 2459 21327 2465
rect 21192 2428 21220 2456
rect 18693 2391 18751 2397
rect 19720 2400 20668 2428
rect 20824 2400 21220 2428
rect 21376 2428 21404 2536
rect 23017 2533 23029 2536
rect 23063 2564 23075 2567
rect 24756 2567 24814 2573
rect 23063 2536 23612 2564
rect 23063 2533 23075 2536
rect 23017 2527 23075 2533
rect 21453 2499 21511 2505
rect 21453 2465 21465 2499
rect 21499 2496 21511 2499
rect 21818 2496 21824 2508
rect 21499 2468 21824 2496
rect 21499 2465 21511 2468
rect 21453 2459 21511 2465
rect 21818 2456 21824 2468
rect 21876 2496 21882 2508
rect 22097 2499 22155 2505
rect 22097 2496 22109 2499
rect 21876 2468 22109 2496
rect 21876 2456 21882 2468
rect 22097 2465 22109 2468
rect 22143 2465 22155 2499
rect 22097 2459 22155 2465
rect 22186 2456 22192 2508
rect 22244 2496 22250 2508
rect 22281 2499 22339 2505
rect 22281 2496 22293 2499
rect 22244 2468 22293 2496
rect 22244 2456 22250 2468
rect 22281 2465 22293 2468
rect 22327 2496 22339 2499
rect 22373 2499 22431 2505
rect 22373 2496 22385 2499
rect 22327 2468 22385 2496
rect 22327 2465 22339 2468
rect 22281 2459 22339 2465
rect 22373 2465 22385 2468
rect 22419 2465 22431 2499
rect 22373 2459 22431 2465
rect 22554 2456 22560 2508
rect 22612 2456 22618 2508
rect 23584 2505 23612 2536
rect 24756 2533 24768 2567
rect 24802 2564 24814 2567
rect 25038 2564 25044 2576
rect 24802 2536 25044 2564
rect 24802 2533 24814 2536
rect 24756 2527 24814 2533
rect 25038 2524 25044 2536
rect 25096 2524 25102 2576
rect 22833 2499 22891 2505
rect 22833 2465 22845 2499
rect 22879 2465 22891 2499
rect 22833 2459 22891 2465
rect 23569 2499 23627 2505
rect 23569 2465 23581 2499
rect 23615 2465 23627 2499
rect 23569 2459 23627 2465
rect 22572 2428 22600 2456
rect 21376 2400 22600 2428
rect 19720 2372 19748 2400
rect 14642 2360 14648 2372
rect 13004 2332 14648 2360
rect 12805 2323 12863 2329
rect 14642 2320 14648 2332
rect 14700 2320 14706 2372
rect 19702 2320 19708 2372
rect 19760 2320 19766 2372
rect 20346 2320 20352 2372
rect 20404 2360 20410 2372
rect 20533 2363 20591 2369
rect 20533 2360 20545 2363
rect 20404 2332 20545 2360
rect 20404 2320 20410 2332
rect 20533 2329 20545 2332
rect 20579 2329 20591 2363
rect 20640 2360 20668 2400
rect 22848 2360 22876 2459
rect 24394 2456 24400 2508
rect 24452 2456 24458 2508
rect 24486 2456 24492 2508
rect 24544 2456 24550 2508
rect 23290 2388 23296 2440
rect 23348 2388 23354 2440
rect 20640 2332 22876 2360
rect 20533 2323 20591 2329
rect 3602 2252 3608 2304
rect 3660 2252 3666 2304
rect 4065 2295 4123 2301
rect 4065 2261 4077 2295
rect 4111 2292 4123 2295
rect 4154 2292 4160 2304
rect 4111 2264 4160 2292
rect 4111 2261 4123 2264
rect 4065 2255 4123 2261
rect 4154 2252 4160 2264
rect 4212 2252 4218 2304
rect 4525 2295 4583 2301
rect 4525 2261 4537 2295
rect 4571 2292 4583 2295
rect 4614 2292 4620 2304
rect 4571 2264 4620 2292
rect 4571 2261 4583 2264
rect 4525 2255 4583 2261
rect 4614 2252 4620 2264
rect 4672 2252 4678 2304
rect 4798 2252 4804 2304
rect 4856 2252 4862 2304
rect 5534 2252 5540 2304
rect 5592 2292 5598 2304
rect 6086 2292 6092 2304
rect 5592 2264 6092 2292
rect 5592 2252 5598 2264
rect 6086 2252 6092 2264
rect 6144 2252 6150 2304
rect 7006 2252 7012 2304
rect 7064 2252 7070 2304
rect 7098 2252 7104 2304
rect 7156 2252 7162 2304
rect 8849 2295 8907 2301
rect 8849 2261 8861 2295
rect 8895 2292 8907 2295
rect 9122 2292 9128 2304
rect 8895 2264 9128 2292
rect 8895 2261 8907 2264
rect 8849 2255 8907 2261
rect 9122 2252 9128 2264
rect 9180 2252 9186 2304
rect 10318 2252 10324 2304
rect 10376 2252 10382 2304
rect 11882 2252 11888 2304
rect 11940 2252 11946 2304
rect 11974 2252 11980 2304
rect 12032 2252 12038 2304
rect 12710 2252 12716 2304
rect 12768 2252 12774 2304
rect 14277 2295 14335 2301
rect 14277 2261 14289 2295
rect 14323 2292 14335 2295
rect 14734 2292 14740 2304
rect 14323 2264 14740 2292
rect 14323 2261 14335 2264
rect 14277 2255 14335 2261
rect 14734 2252 14740 2264
rect 14792 2292 14798 2304
rect 14918 2292 14924 2304
rect 14792 2264 14924 2292
rect 14792 2252 14798 2264
rect 14918 2252 14924 2264
rect 14976 2252 14982 2304
rect 20438 2252 20444 2304
rect 20496 2252 20502 2304
rect 20990 2252 20996 2304
rect 21048 2252 21054 2304
rect 21269 2295 21327 2301
rect 21269 2261 21281 2295
rect 21315 2292 21327 2295
rect 21542 2292 21548 2304
rect 21315 2264 21548 2292
rect 21315 2261 21327 2264
rect 21269 2255 21327 2261
rect 21542 2252 21548 2264
rect 21600 2252 21606 2304
rect 552 2202 27416 2224
rect 552 2150 3756 2202
rect 3808 2150 3820 2202
rect 3872 2150 3884 2202
rect 3936 2150 3948 2202
rect 4000 2150 4012 2202
rect 4064 2150 10472 2202
rect 10524 2150 10536 2202
rect 10588 2150 10600 2202
rect 10652 2150 10664 2202
rect 10716 2150 10728 2202
rect 10780 2150 17188 2202
rect 17240 2150 17252 2202
rect 17304 2150 17316 2202
rect 17368 2150 17380 2202
rect 17432 2150 17444 2202
rect 17496 2150 23904 2202
rect 23956 2150 23968 2202
rect 24020 2150 24032 2202
rect 24084 2150 24096 2202
rect 24148 2150 24160 2202
rect 24212 2150 27416 2202
rect 552 2128 27416 2150
rect 4062 2048 4068 2100
rect 4120 2048 4126 2100
rect 4798 2048 4804 2100
rect 4856 2048 4862 2100
rect 4890 2048 4896 2100
rect 4948 2088 4954 2100
rect 5626 2088 5632 2100
rect 4948 2060 5632 2088
rect 4948 2048 4954 2060
rect 5626 2048 5632 2060
rect 5684 2088 5690 2100
rect 6638 2088 6644 2100
rect 5684 2060 6644 2088
rect 5684 2048 5690 2060
rect 6638 2048 6644 2060
rect 6696 2048 6702 2100
rect 7006 2088 7012 2100
rect 6748 2060 7012 2088
rect 4080 1961 4108 2048
rect 4065 1955 4123 1961
rect 4065 1921 4077 1955
rect 4111 1921 4123 1955
rect 4065 1915 4123 1921
rect 934 1844 940 1896
rect 992 1844 998 1896
rect 1118 1844 1124 1896
rect 1176 1884 1182 1896
rect 1305 1887 1363 1893
rect 1305 1884 1317 1887
rect 1176 1856 1317 1884
rect 1176 1844 1182 1856
rect 1305 1853 1317 1856
rect 1351 1853 1363 1887
rect 1305 1847 1363 1853
rect 1765 1887 1823 1893
rect 1765 1853 1777 1887
rect 1811 1884 1823 1887
rect 1857 1887 1915 1893
rect 1857 1884 1869 1887
rect 1811 1856 1869 1884
rect 1811 1853 1823 1856
rect 1765 1847 1823 1853
rect 1857 1853 1869 1856
rect 1903 1853 1915 1887
rect 1857 1847 1915 1853
rect 2133 1887 2191 1893
rect 2133 1853 2145 1887
rect 2179 1884 2191 1887
rect 2682 1884 2688 1896
rect 2179 1856 2688 1884
rect 2179 1853 2191 1856
rect 2133 1847 2191 1853
rect 2682 1844 2688 1856
rect 2740 1844 2746 1896
rect 2958 1844 2964 1896
rect 3016 1844 3022 1896
rect 3237 1887 3295 1893
rect 3237 1853 3249 1887
rect 3283 1884 3295 1887
rect 3326 1884 3332 1896
rect 3283 1856 3332 1884
rect 3283 1853 3295 1856
rect 3237 1847 3295 1853
rect 3326 1844 3332 1856
rect 3384 1844 3390 1896
rect 3510 1844 3516 1896
rect 3568 1884 3574 1896
rect 3697 1887 3755 1893
rect 3697 1884 3709 1887
rect 3568 1856 3709 1884
rect 3568 1844 3574 1856
rect 3697 1853 3709 1856
rect 3743 1853 3755 1887
rect 3697 1847 3755 1853
rect 3973 1887 4031 1893
rect 3973 1853 3985 1887
rect 4019 1853 4031 1887
rect 3973 1847 4031 1853
rect 4341 1887 4399 1893
rect 4341 1853 4353 1887
rect 4387 1884 4399 1887
rect 4816 1884 4844 2048
rect 6748 1961 6776 2060
rect 7006 2048 7012 2060
rect 7064 2048 7070 2100
rect 10318 2048 10324 2100
rect 10376 2048 10382 2100
rect 11054 2048 11060 2100
rect 11112 2088 11118 2100
rect 15010 2088 15016 2100
rect 11112 2060 15016 2088
rect 11112 2048 11118 2060
rect 15010 2048 15016 2060
rect 15068 2048 15074 2100
rect 16942 2048 16948 2100
rect 17000 2088 17006 2100
rect 17497 2091 17555 2097
rect 17497 2088 17509 2091
rect 17000 2060 17509 2088
rect 17000 2048 17006 2060
rect 17497 2057 17509 2060
rect 17543 2057 17555 2091
rect 21361 2091 21419 2097
rect 21361 2088 21373 2091
rect 17497 2051 17555 2057
rect 20180 2060 21373 2088
rect 10336 2020 10364 2048
rect 10336 1992 10456 2020
rect 10428 1961 10456 1992
rect 20180 1961 20208 2060
rect 21361 2057 21373 2060
rect 21407 2057 21419 2091
rect 21361 2051 21419 2057
rect 6733 1955 6791 1961
rect 6733 1921 6745 1955
rect 6779 1921 6791 1955
rect 6733 1915 6791 1921
rect 10413 1955 10471 1961
rect 10413 1921 10425 1955
rect 10459 1921 10471 1955
rect 10413 1915 10471 1921
rect 20165 1955 20223 1961
rect 20165 1921 20177 1955
rect 20211 1921 20223 1955
rect 20165 1915 20223 1921
rect 4387 1856 4844 1884
rect 4387 1853 4399 1856
rect 4341 1847 4399 1853
rect 3988 1816 4016 1847
rect 5166 1844 5172 1896
rect 5224 1844 5230 1896
rect 5258 1844 5264 1896
rect 5316 1844 5322 1896
rect 5537 1887 5595 1893
rect 5537 1853 5549 1887
rect 5583 1884 5595 1887
rect 5718 1884 5724 1896
rect 5583 1856 5724 1884
rect 5583 1853 5595 1856
rect 5537 1847 5595 1853
rect 5718 1844 5724 1856
rect 5776 1844 5782 1896
rect 5810 1844 5816 1896
rect 5868 1844 5874 1896
rect 6638 1844 6644 1896
rect 6696 1844 6702 1896
rect 7009 1887 7067 1893
rect 7009 1853 7021 1887
rect 7055 1884 7067 1887
rect 7098 1884 7104 1896
rect 7055 1856 7104 1884
rect 7055 1853 7067 1856
rect 7009 1847 7067 1853
rect 7098 1844 7104 1856
rect 7156 1844 7162 1896
rect 7834 1844 7840 1896
rect 7892 1844 7898 1896
rect 7926 1844 7932 1896
rect 7984 1844 7990 1896
rect 9214 1844 9220 1896
rect 9272 1844 9278 1896
rect 9309 1887 9367 1893
rect 9309 1853 9321 1887
rect 9355 1853 9367 1887
rect 9309 1847 9367 1853
rect 4062 1816 4068 1828
rect 3988 1788 4068 1816
rect 4062 1776 4068 1788
rect 4120 1776 4126 1828
rect 3510 1708 3516 1760
rect 3568 1708 3574 1760
rect 9324 1748 9352 1847
rect 10134 1844 10140 1896
rect 10192 1844 10198 1896
rect 10505 1887 10563 1893
rect 10505 1853 10517 1887
rect 10551 1853 10563 1887
rect 10505 1847 10563 1853
rect 10318 1776 10324 1828
rect 10376 1816 10382 1828
rect 10520 1816 10548 1847
rect 10778 1844 10784 1896
rect 10836 1844 10842 1896
rect 11606 1844 11612 1896
rect 11664 1844 11670 1896
rect 11698 1844 11704 1896
rect 11756 1844 11762 1896
rect 11974 1844 11980 1896
rect 12032 1844 12038 1896
rect 12802 1844 12808 1896
rect 12860 1844 12866 1896
rect 12894 1844 12900 1896
rect 12952 1844 12958 1896
rect 13170 1844 13176 1896
rect 13228 1844 13234 1896
rect 14182 1844 14188 1896
rect 14240 1844 14246 1896
rect 14642 1844 14648 1896
rect 14700 1844 14706 1896
rect 15105 1887 15163 1893
rect 15105 1853 15117 1887
rect 15151 1884 15163 1887
rect 15197 1887 15255 1893
rect 15197 1884 15209 1887
rect 15151 1856 15209 1884
rect 15151 1853 15163 1856
rect 15105 1847 15163 1853
rect 15197 1853 15209 1856
rect 15243 1853 15255 1887
rect 15197 1847 15255 1853
rect 15378 1844 15384 1896
rect 15436 1884 15442 1896
rect 15473 1887 15531 1893
rect 15473 1884 15485 1887
rect 15436 1856 15485 1884
rect 15436 1844 15442 1856
rect 15473 1853 15485 1856
rect 15519 1853 15531 1887
rect 15473 1847 15531 1853
rect 16298 1844 16304 1896
rect 16356 1844 16362 1896
rect 16390 1844 16396 1896
rect 16448 1844 16454 1896
rect 16853 1887 16911 1893
rect 16853 1853 16865 1887
rect 16899 1884 16911 1887
rect 17310 1884 17316 1896
rect 16899 1856 17316 1884
rect 16899 1853 16911 1856
rect 16853 1847 16911 1853
rect 17310 1844 17316 1856
rect 17368 1844 17374 1896
rect 17678 1844 17684 1896
rect 17736 1844 17742 1896
rect 18877 1887 18935 1893
rect 18877 1853 18889 1887
rect 18923 1884 18935 1887
rect 18969 1887 19027 1893
rect 18969 1884 18981 1887
rect 18923 1856 18981 1884
rect 18923 1853 18935 1856
rect 18877 1847 18935 1853
rect 18969 1853 18981 1856
rect 19015 1853 19027 1887
rect 18969 1847 19027 1853
rect 19245 1887 19303 1893
rect 19245 1853 19257 1887
rect 19291 1884 19303 1887
rect 19794 1884 19800 1896
rect 19291 1856 19800 1884
rect 19291 1853 19303 1856
rect 19245 1847 19303 1853
rect 19794 1844 19800 1856
rect 19852 1844 19858 1896
rect 20070 1844 20076 1896
rect 20128 1844 20134 1896
rect 20438 1844 20444 1896
rect 20496 1844 20502 1896
rect 21266 1844 21272 1896
rect 21324 1844 21330 1896
rect 21450 1844 21456 1896
rect 21508 1884 21514 1896
rect 21637 1887 21695 1893
rect 21637 1884 21649 1887
rect 21508 1856 21649 1884
rect 21508 1844 21514 1856
rect 21637 1853 21649 1856
rect 21683 1853 21695 1887
rect 21637 1847 21695 1853
rect 21910 1844 21916 1896
rect 21968 1844 21974 1896
rect 22373 1887 22431 1893
rect 22373 1853 22385 1887
rect 22419 1884 22431 1887
rect 22554 1884 22560 1896
rect 22419 1856 22560 1884
rect 22419 1853 22431 1856
rect 22373 1847 22431 1853
rect 22554 1844 22560 1856
rect 22612 1844 22618 1896
rect 22646 1844 22652 1896
rect 22704 1844 22710 1896
rect 23290 1844 23296 1896
rect 23348 1884 23354 1896
rect 23477 1887 23535 1893
rect 23477 1884 23489 1887
rect 23348 1856 23489 1884
rect 23348 1844 23354 1856
rect 23477 1853 23489 1856
rect 23523 1853 23535 1887
rect 23477 1847 23535 1853
rect 23750 1844 23756 1896
rect 23808 1884 23814 1896
rect 23845 1887 23903 1893
rect 23845 1884 23857 1887
rect 23808 1856 23857 1884
rect 23808 1844 23814 1856
rect 23845 1853 23857 1856
rect 23891 1853 23903 1887
rect 23845 1847 23903 1853
rect 24581 1887 24639 1893
rect 24581 1853 24593 1887
rect 24627 1853 24639 1887
rect 24581 1847 24639 1853
rect 10376 1788 10548 1816
rect 24596 1816 24624 1847
rect 24854 1844 24860 1896
rect 24912 1844 24918 1896
rect 25685 1887 25743 1893
rect 25685 1853 25697 1887
rect 25731 1884 25743 1887
rect 26050 1884 26056 1896
rect 25731 1856 26056 1884
rect 25731 1853 25743 1856
rect 25685 1847 25743 1853
rect 26050 1844 26056 1856
rect 26108 1844 26114 1896
rect 25314 1816 25320 1828
rect 24596 1788 25320 1816
rect 10376 1776 10382 1788
rect 25314 1776 25320 1788
rect 25372 1776 25378 1828
rect 11146 1748 11152 1760
rect 9324 1720 11152 1748
rect 11146 1708 11152 1720
rect 11204 1708 11210 1760
rect 552 1658 27576 1680
rect 552 1606 7114 1658
rect 7166 1606 7178 1658
rect 7230 1606 7242 1658
rect 7294 1606 7306 1658
rect 7358 1606 7370 1658
rect 7422 1606 13830 1658
rect 13882 1606 13894 1658
rect 13946 1606 13958 1658
rect 14010 1606 14022 1658
rect 14074 1606 14086 1658
rect 14138 1606 20546 1658
rect 20598 1606 20610 1658
rect 20662 1606 20674 1658
rect 20726 1606 20738 1658
rect 20790 1606 20802 1658
rect 20854 1606 27262 1658
rect 27314 1606 27326 1658
rect 27378 1606 27390 1658
rect 27442 1606 27454 1658
rect 27506 1606 27518 1658
rect 27570 1606 27576 1658
rect 552 1584 27576 1606
rect 1302 1504 1308 1556
rect 1360 1504 1366 1556
rect 2038 1504 2044 1556
rect 2096 1504 2102 1556
rect 3510 1504 3516 1556
rect 3568 1504 3574 1556
rect 6270 1504 6276 1556
rect 6328 1544 6334 1556
rect 7374 1544 7380 1556
rect 6328 1516 7380 1544
rect 6328 1504 6334 1516
rect 7374 1504 7380 1516
rect 7432 1504 7438 1556
rect 7926 1504 7932 1556
rect 7984 1504 7990 1556
rect 11882 1504 11888 1556
rect 11940 1504 11946 1556
rect 19702 1504 19708 1556
rect 19760 1504 19766 1556
rect 20990 1504 20996 1556
rect 21048 1504 21054 1556
rect 22830 1504 22836 1556
rect 22888 1504 22894 1556
rect 937 1411 995 1417
rect 937 1377 949 1411
rect 983 1408 995 1411
rect 1118 1408 1124 1420
rect 983 1380 1124 1408
rect 983 1377 995 1380
rect 937 1371 995 1377
rect 1118 1368 1124 1380
rect 1176 1368 1182 1420
rect 1213 1411 1271 1417
rect 1213 1377 1225 1411
rect 1259 1408 1271 1411
rect 1320 1408 1348 1504
rect 2056 1476 2084 1504
rect 2056 1448 2452 1476
rect 1259 1380 1348 1408
rect 2041 1411 2099 1417
rect 1259 1377 1271 1380
rect 1213 1371 1271 1377
rect 2041 1377 2053 1411
rect 2087 1408 2099 1411
rect 2314 1408 2320 1420
rect 2087 1380 2320 1408
rect 2087 1377 2099 1380
rect 2041 1371 2099 1377
rect 2314 1368 2320 1380
rect 2372 1368 2378 1420
rect 2424 1417 2452 1448
rect 2409 1411 2467 1417
rect 2409 1377 2421 1411
rect 2455 1377 2467 1411
rect 2409 1371 2467 1377
rect 3234 1368 3240 1420
rect 3292 1368 3298 1420
rect 3528 1408 3556 1504
rect 6178 1476 6184 1488
rect 4540 1448 5304 1476
rect 3605 1411 3663 1417
rect 3605 1408 3617 1411
rect 3528 1380 3617 1408
rect 3605 1377 3617 1380
rect 3651 1377 3663 1411
rect 3605 1371 3663 1377
rect 4430 1368 4436 1420
rect 4488 1368 4494 1420
rect 4540 1417 4568 1448
rect 5276 1420 5304 1448
rect 5644 1448 6184 1476
rect 4525 1411 4583 1417
rect 4525 1377 4537 1411
rect 4571 1377 4583 1411
rect 4525 1371 4583 1377
rect 4706 1368 4712 1420
rect 4764 1408 4770 1420
rect 4801 1411 4859 1417
rect 4801 1408 4813 1411
rect 4764 1380 4813 1408
rect 4764 1368 4770 1380
rect 4801 1377 4813 1380
rect 4847 1377 4859 1411
rect 4801 1371 4859 1377
rect 5258 1368 5264 1420
rect 5316 1368 5322 1420
rect 5644 1417 5672 1448
rect 6178 1436 6184 1448
rect 6236 1436 6242 1488
rect 7944 1476 7972 1504
rect 8938 1476 8944 1488
rect 7024 1448 7972 1476
rect 8220 1448 8944 1476
rect 5629 1411 5687 1417
rect 5629 1377 5641 1411
rect 5675 1377 5687 1411
rect 5629 1371 5687 1377
rect 5718 1368 5724 1420
rect 5776 1408 5782 1420
rect 5813 1411 5871 1417
rect 5813 1408 5825 1411
rect 5776 1380 5825 1408
rect 5776 1368 5782 1380
rect 5813 1377 5825 1380
rect 5859 1377 5871 1411
rect 7024 1408 7052 1448
rect 5813 1371 5871 1377
rect 6840 1380 7052 1408
rect 2130 1300 2136 1352
rect 2188 1300 2194 1352
rect 3326 1300 3332 1352
rect 3384 1300 3390 1352
rect 6840 1349 6868 1380
rect 7098 1368 7104 1420
rect 7156 1368 7162 1420
rect 7929 1411 7987 1417
rect 7929 1377 7941 1411
rect 7975 1408 7987 1411
rect 8220 1408 8248 1448
rect 8938 1436 8944 1448
rect 8996 1436 9002 1488
rect 7975 1380 8248 1408
rect 7975 1377 7987 1380
rect 7929 1371 7987 1377
rect 8294 1368 8300 1420
rect 8352 1368 8358 1420
rect 9125 1411 9183 1417
rect 9125 1377 9137 1411
rect 9171 1408 9183 1411
rect 9306 1408 9312 1420
rect 9171 1380 9312 1408
rect 9171 1377 9183 1380
rect 9125 1371 9183 1377
rect 9306 1368 9312 1380
rect 9364 1368 9370 1420
rect 9858 1368 9864 1420
rect 9916 1368 9922 1420
rect 10686 1368 10692 1420
rect 10744 1368 10750 1420
rect 11333 1411 11391 1417
rect 11333 1377 11345 1411
rect 11379 1408 11391 1411
rect 11900 1408 11928 1504
rect 12406 1448 12940 1476
rect 11379 1380 11928 1408
rect 11379 1377 11391 1380
rect 11333 1371 11391 1377
rect 12158 1368 12164 1420
rect 12216 1368 12222 1420
rect 12406 1408 12434 1448
rect 12912 1420 12940 1448
rect 17034 1436 17040 1488
rect 17092 1476 17098 1488
rect 17092 1448 17632 1476
rect 17092 1436 17098 1448
rect 12268 1380 12434 1408
rect 12529 1411 12587 1417
rect 6825 1343 6883 1349
rect 6825 1309 6837 1343
rect 6871 1309 6883 1343
rect 6825 1303 6883 1309
rect 8018 1300 8024 1352
rect 8076 1300 8082 1352
rect 9493 1343 9551 1349
rect 9493 1309 9505 1343
rect 9539 1340 9551 1343
rect 9585 1343 9643 1349
rect 9585 1340 9597 1343
rect 9539 1312 9597 1340
rect 9539 1309 9551 1312
rect 9493 1303 9551 1309
rect 9585 1309 9597 1312
rect 9631 1309 9643 1343
rect 9585 1303 9643 1309
rect 11054 1300 11060 1352
rect 11112 1300 11118 1352
rect 12268 1349 12296 1380
rect 12529 1377 12541 1411
rect 12575 1408 12587 1411
rect 12618 1408 12624 1420
rect 12575 1380 12624 1408
rect 12575 1377 12587 1380
rect 12529 1371 12587 1377
rect 12618 1368 12624 1380
rect 12676 1368 12682 1420
rect 12894 1368 12900 1420
rect 12952 1368 12958 1420
rect 13357 1411 13415 1417
rect 13357 1377 13369 1411
rect 13403 1408 13415 1411
rect 13630 1408 13636 1420
rect 13403 1380 13636 1408
rect 13403 1377 13415 1380
rect 13357 1371 13415 1377
rect 13630 1368 13636 1380
rect 13688 1368 13694 1420
rect 13722 1368 13728 1420
rect 13780 1368 13786 1420
rect 14550 1368 14556 1420
rect 14608 1368 14614 1420
rect 14642 1368 14648 1420
rect 14700 1368 14706 1420
rect 14918 1368 14924 1420
rect 14976 1368 14982 1420
rect 15746 1368 15752 1420
rect 15804 1368 15810 1420
rect 15838 1368 15844 1420
rect 15896 1408 15902 1420
rect 16393 1411 16451 1417
rect 16393 1408 16405 1411
rect 15896 1380 16405 1408
rect 15896 1368 15902 1380
rect 16393 1377 16405 1380
rect 16439 1377 16451 1411
rect 16393 1371 16451 1377
rect 16758 1368 16764 1420
rect 16816 1408 16822 1420
rect 17221 1411 17279 1417
rect 17221 1408 17233 1411
rect 16816 1380 17233 1408
rect 16816 1368 16822 1380
rect 17221 1377 17233 1380
rect 17267 1377 17279 1411
rect 17221 1371 17279 1377
rect 17310 1368 17316 1420
rect 17368 1368 17374 1420
rect 17604 1417 17632 1448
rect 17589 1411 17647 1417
rect 17589 1377 17601 1411
rect 17635 1377 17647 1411
rect 17589 1371 17647 1377
rect 17770 1368 17776 1420
rect 17828 1408 17834 1420
rect 18417 1411 18475 1417
rect 18417 1408 18429 1411
rect 17828 1380 18429 1408
rect 17828 1368 17834 1380
rect 18417 1377 18429 1380
rect 18463 1377 18475 1411
rect 18417 1371 18475 1377
rect 18506 1368 18512 1420
rect 18564 1368 18570 1420
rect 19334 1368 19340 1420
rect 19392 1368 19398 1420
rect 19720 1408 19748 1504
rect 19886 1436 19892 1488
rect 19944 1476 19950 1488
rect 21008 1476 21036 1504
rect 19944 1448 20852 1476
rect 21008 1448 21588 1476
rect 19944 1436 19950 1448
rect 20824 1417 20852 1448
rect 19981 1411 20039 1417
rect 19981 1408 19993 1411
rect 19720 1380 19993 1408
rect 19981 1377 19993 1380
rect 20027 1377 20039 1411
rect 19981 1371 20039 1377
rect 20809 1411 20867 1417
rect 20809 1377 20821 1411
rect 20855 1377 20867 1411
rect 20809 1371 20867 1377
rect 21269 1411 21327 1417
rect 21269 1377 21281 1411
rect 21315 1408 21327 1411
rect 21450 1408 21456 1420
rect 21315 1380 21456 1408
rect 21315 1377 21327 1380
rect 21269 1371 21327 1377
rect 21450 1368 21456 1380
rect 21508 1368 21514 1420
rect 21560 1417 21588 1448
rect 22094 1436 22100 1488
rect 22152 1476 22158 1488
rect 22848 1476 22876 1504
rect 22152 1448 22784 1476
rect 22848 1448 23980 1476
rect 22152 1436 22158 1448
rect 21545 1411 21603 1417
rect 21545 1377 21557 1411
rect 21591 1377 21603 1411
rect 21545 1371 21603 1377
rect 22002 1368 22008 1420
rect 22060 1408 22066 1420
rect 22756 1417 22784 1448
rect 22373 1411 22431 1417
rect 22373 1408 22385 1411
rect 22060 1380 22385 1408
rect 22060 1368 22066 1380
rect 22373 1377 22385 1380
rect 22419 1377 22431 1411
rect 22373 1371 22431 1377
rect 22741 1411 22799 1417
rect 22741 1377 22753 1411
rect 22787 1377 22799 1411
rect 22741 1371 22799 1377
rect 22830 1368 22836 1420
rect 22888 1408 22894 1420
rect 23952 1417 23980 1448
rect 23569 1411 23627 1417
rect 23569 1408 23581 1411
rect 22888 1380 23581 1408
rect 22888 1368 22894 1380
rect 23569 1377 23581 1380
rect 23615 1377 23627 1411
rect 23569 1371 23627 1377
rect 23937 1411 23995 1417
rect 23937 1377 23949 1411
rect 23983 1377 23995 1411
rect 23937 1371 23995 1377
rect 24302 1368 24308 1420
rect 24360 1408 24366 1420
rect 24765 1411 24823 1417
rect 24765 1408 24777 1411
rect 24360 1380 24777 1408
rect 24360 1368 24366 1380
rect 24765 1377 24777 1380
rect 24811 1377 24823 1411
rect 24765 1371 24823 1377
rect 25130 1368 25136 1420
rect 25188 1368 25194 1420
rect 25498 1368 25504 1420
rect 25556 1408 25562 1420
rect 25961 1411 26019 1417
rect 25961 1408 25973 1411
rect 25556 1380 25973 1408
rect 25556 1368 25562 1380
rect 25961 1377 25973 1380
rect 26007 1377 26019 1411
rect 25961 1371 26019 1377
rect 12253 1343 12311 1349
rect 12253 1309 12265 1343
rect 12299 1309 12311 1343
rect 12253 1303 12311 1309
rect 13446 1300 13452 1352
rect 13504 1300 13510 1352
rect 16114 1300 16120 1352
rect 16172 1300 16178 1352
rect 19613 1343 19671 1349
rect 19613 1309 19625 1343
rect 19659 1309 19671 1343
rect 19613 1303 19671 1309
rect 6270 1164 6276 1216
rect 6328 1164 6334 1216
rect 6730 1164 6736 1216
rect 6788 1164 6794 1216
rect 17862 1164 17868 1216
rect 17920 1204 17926 1216
rect 19628 1204 19656 1303
rect 19702 1300 19708 1352
rect 19760 1300 19766 1352
rect 22462 1300 22468 1352
rect 22520 1300 22526 1352
rect 23658 1300 23664 1352
rect 23716 1300 23722 1352
rect 24854 1300 24860 1352
rect 24912 1300 24918 1352
rect 17920 1176 19656 1204
rect 17920 1164 17926 1176
rect 21082 1164 21088 1216
rect 21140 1164 21146 1216
rect 552 1114 27416 1136
rect 552 1062 3756 1114
rect 3808 1062 3820 1114
rect 3872 1062 3884 1114
rect 3936 1062 3948 1114
rect 4000 1062 4012 1114
rect 4064 1062 10472 1114
rect 10524 1062 10536 1114
rect 10588 1062 10600 1114
rect 10652 1062 10664 1114
rect 10716 1062 10728 1114
rect 10780 1062 17188 1114
rect 17240 1062 17252 1114
rect 17304 1062 17316 1114
rect 17368 1062 17380 1114
rect 17432 1062 17444 1114
rect 17496 1062 23904 1114
rect 23956 1062 23968 1114
rect 24020 1062 24032 1114
rect 24084 1062 24096 1114
rect 24148 1062 24160 1114
rect 24212 1062 27416 1114
rect 552 1040 27416 1062
rect 2130 960 2136 1012
rect 2188 1000 2194 1012
rect 2225 1003 2283 1009
rect 2225 1000 2237 1003
rect 2188 972 2237 1000
rect 2188 960 2194 972
rect 2225 969 2237 972
rect 2271 969 2283 1003
rect 2225 963 2283 969
rect 4154 960 4160 1012
rect 4212 960 4218 1012
rect 6270 1000 6276 1012
rect 5920 972 6276 1000
rect 934 824 940 876
rect 992 824 998 876
rect 4172 864 4200 960
rect 5920 873 5948 972
rect 6270 960 6276 972
rect 6328 960 6334 1012
rect 6730 960 6736 1012
rect 6788 960 6794 1012
rect 8018 960 8024 1012
rect 8076 1000 8082 1012
rect 8389 1003 8447 1009
rect 8389 1000 8401 1003
rect 8076 972 8401 1000
rect 8076 960 8082 972
rect 8389 969 8401 972
rect 8435 969 8447 1003
rect 8389 963 8447 969
rect 10318 960 10324 1012
rect 10376 1000 10382 1012
rect 10597 1003 10655 1009
rect 10597 1000 10609 1003
rect 10376 972 10609 1000
rect 10376 960 10382 972
rect 10597 969 10609 972
rect 10643 969 10655 1003
rect 10597 963 10655 969
rect 11054 960 11060 1012
rect 11112 1000 11118 1012
rect 11241 1003 11299 1009
rect 11241 1000 11253 1003
rect 11112 972 11253 1000
rect 11112 960 11118 972
rect 11241 969 11253 972
rect 11287 969 11299 1003
rect 11241 963 11299 969
rect 11698 960 11704 1012
rect 11756 960 11762 1012
rect 13170 1000 13176 1012
rect 12268 972 13176 1000
rect 4433 867 4491 873
rect 4433 864 4445 867
rect 4172 836 4445 864
rect 4433 833 4445 836
rect 4479 833 4491 867
rect 4433 827 4491 833
rect 5905 867 5963 873
rect 5905 833 5917 867
rect 5951 833 5963 867
rect 6748 864 6776 960
rect 7101 867 7159 873
rect 7101 864 7113 867
rect 6748 836 7113 864
rect 5905 827 5963 833
rect 7101 833 7113 836
rect 7147 833 7159 867
rect 7101 827 7159 833
rect 9214 824 9220 876
rect 9272 824 9278 876
rect 12268 873 12296 972
rect 13170 960 13176 972
rect 13228 960 13234 1012
rect 13446 960 13452 1012
rect 13504 1000 13510 1012
rect 13541 1003 13599 1009
rect 13541 1000 13553 1003
rect 13504 972 13553 1000
rect 13504 960 13510 972
rect 13541 969 13553 972
rect 13587 969 13599 1003
rect 13541 963 13599 969
rect 14182 960 14188 1012
rect 14240 960 14246 1012
rect 15749 1003 15807 1009
rect 15749 969 15761 1003
rect 15795 1000 15807 1003
rect 16114 1000 16120 1012
rect 15795 972 16120 1000
rect 15795 969 15807 972
rect 15749 963 15807 969
rect 16114 960 16120 972
rect 16172 960 16178 1012
rect 17862 960 17868 1012
rect 17920 960 17926 1012
rect 18509 1003 18567 1009
rect 18509 969 18521 1003
rect 18555 1000 18567 1003
rect 19702 1000 19708 1012
rect 18555 972 19708 1000
rect 18555 969 18567 972
rect 18509 963 18567 969
rect 19702 960 19708 972
rect 19760 960 19766 1012
rect 21082 960 21088 1012
rect 21140 960 21146 1012
rect 21910 1000 21916 1012
rect 21284 972 21916 1000
rect 14200 932 14228 960
rect 14108 904 14228 932
rect 14108 873 14136 904
rect 12253 867 12311 873
rect 12253 833 12265 867
rect 12299 833 12311 867
rect 12253 827 12311 833
rect 14093 867 14151 873
rect 14093 833 14105 867
rect 14139 833 14151 867
rect 14093 827 14151 833
rect 18233 867 18291 873
rect 18233 833 18245 867
rect 18279 864 18291 867
rect 18693 867 18751 873
rect 18693 864 18705 867
rect 18279 836 18705 864
rect 18279 833 18291 836
rect 18233 827 18291 833
rect 18693 833 18705 836
rect 18739 833 18751 867
rect 18693 827 18751 833
rect 20993 867 21051 873
rect 20993 833 21005 867
rect 21039 864 21051 867
rect 21100 864 21128 960
rect 21284 873 21312 972
rect 21910 960 21916 972
rect 21968 960 21974 1012
rect 22462 960 22468 1012
rect 22520 960 22526 1012
rect 22554 960 22560 1012
rect 22612 1000 22618 1012
rect 22741 1003 22799 1009
rect 22741 1000 22753 1003
rect 22612 972 22753 1000
rect 22612 960 22618 972
rect 22741 969 22753 972
rect 22787 969 22799 1003
rect 22741 963 22799 969
rect 23201 1003 23259 1009
rect 23201 969 23213 1003
rect 23247 1000 23259 1003
rect 23658 1000 23664 1012
rect 23247 972 23664 1000
rect 23247 969 23259 972
rect 23201 963 23259 969
rect 23658 960 23664 972
rect 23716 960 23722 1012
rect 24854 960 24860 1012
rect 24912 1000 24918 1012
rect 25041 1003 25099 1009
rect 25041 1000 25053 1003
rect 24912 972 25053 1000
rect 24912 960 24918 972
rect 25041 969 25053 972
rect 25087 969 25099 1003
rect 25041 963 25099 969
rect 25314 960 25320 1012
rect 25372 960 25378 1012
rect 21039 836 21128 864
rect 21269 867 21327 873
rect 21039 833 21051 836
rect 20993 827 21051 833
rect 21269 833 21281 867
rect 21315 833 21327 867
rect 21269 827 21327 833
rect 23750 824 23756 876
rect 23808 864 23814 876
rect 23845 867 23903 873
rect 23845 864 23857 867
rect 23808 836 23857 864
rect 23808 824 23814 836
rect 23845 833 23857 836
rect 23891 833 23903 867
rect 23845 827 23903 833
rect 1213 799 1271 805
rect 1213 765 1225 799
rect 1259 765 1271 799
rect 1213 759 1271 765
rect 1228 728 1256 759
rect 1762 756 1768 808
rect 1820 796 1826 808
rect 2041 799 2099 805
rect 2041 796 2053 799
rect 1820 768 2053 796
rect 1820 756 1826 768
rect 2041 765 2053 768
rect 2087 765 2099 799
rect 2041 759 2099 765
rect 2498 756 2504 808
rect 2556 756 2562 808
rect 3053 799 3111 805
rect 3053 765 3065 799
rect 3099 796 3111 799
rect 3237 799 3295 805
rect 3237 796 3249 799
rect 3099 768 3249 796
rect 3099 765 3111 768
rect 3053 759 3111 765
rect 3237 765 3249 768
rect 3283 765 3295 799
rect 3237 759 3295 765
rect 3513 799 3571 805
rect 3513 765 3525 799
rect 3559 796 3571 799
rect 3602 796 3608 808
rect 3559 768 3608 796
rect 3559 765 3571 768
rect 3513 759 3571 765
rect 3602 756 3608 768
rect 3660 756 3666 808
rect 4062 756 4068 808
rect 4120 796 4126 808
rect 4341 799 4399 805
rect 4341 796 4353 799
rect 4120 768 4353 796
rect 4120 756 4126 768
rect 4341 765 4353 768
rect 4387 765 4399 799
rect 4341 759 4399 765
rect 4614 756 4620 808
rect 4672 796 4678 808
rect 4709 799 4767 805
rect 4709 796 4721 799
rect 4672 768 4721 796
rect 4672 756 4678 768
rect 4709 765 4721 768
rect 4755 765 4767 799
rect 4709 759 4767 765
rect 5534 756 5540 808
rect 5592 756 5598 808
rect 6086 756 6092 808
rect 6144 796 6150 808
rect 6181 799 6239 805
rect 6181 796 6193 799
rect 6144 768 6193 796
rect 6144 756 6150 768
rect 6181 765 6193 768
rect 6227 765 6239 799
rect 6181 759 6239 765
rect 7006 756 7012 808
rect 7064 756 7070 808
rect 7374 756 7380 808
rect 7432 756 7438 808
rect 8205 799 8263 805
rect 8205 765 8217 799
rect 8251 796 8263 799
rect 8294 796 8300 808
rect 8251 768 8300 796
rect 8251 765 8263 768
rect 8205 759 8263 765
rect 8294 756 8300 768
rect 8352 756 8358 808
rect 9493 799 9551 805
rect 9493 765 9505 799
rect 9539 796 9551 799
rect 9674 796 9680 808
rect 9539 768 9680 796
rect 9539 765 9551 768
rect 9493 759 9551 765
rect 9674 756 9680 768
rect 9732 756 9738 808
rect 10042 756 10048 808
rect 10100 796 10106 808
rect 10321 799 10379 805
rect 10321 796 10333 799
rect 10100 768 10333 796
rect 10100 756 10106 768
rect 10321 765 10333 768
rect 10367 765 10379 799
rect 10321 759 10379 765
rect 12529 799 12587 805
rect 12529 765 12541 799
rect 12575 796 12587 799
rect 12710 796 12716 808
rect 12575 768 12716 796
rect 12575 765 12587 768
rect 12529 759 12587 765
rect 12710 756 12716 768
rect 12768 756 12774 808
rect 13354 756 13360 808
rect 13412 756 13418 808
rect 14369 799 14427 805
rect 14369 765 14381 799
rect 14415 796 14427 799
rect 14826 796 14832 808
rect 14415 768 14832 796
rect 14415 765 14427 768
rect 14369 759 14427 765
rect 14826 756 14832 768
rect 14884 756 14890 808
rect 15010 756 15016 808
rect 15068 796 15074 808
rect 15197 799 15255 805
rect 15197 796 15209 799
rect 15068 768 15209 796
rect 15068 756 15074 768
rect 15197 765 15209 768
rect 15243 765 15255 799
rect 15197 759 15255 765
rect 16209 799 16267 805
rect 16209 765 16221 799
rect 16255 796 16267 799
rect 16390 796 16396 808
rect 16255 768 16396 796
rect 16255 765 16267 768
rect 16209 759 16267 765
rect 16390 756 16396 768
rect 16448 756 16454 808
rect 16485 799 16543 805
rect 16485 765 16497 799
rect 16531 765 16543 799
rect 16485 759 16543 765
rect 2516 728 2544 756
rect 1228 700 2544 728
rect 15930 688 15936 740
rect 15988 728 15994 740
rect 16500 728 16528 759
rect 17310 756 17316 808
rect 17368 756 17374 808
rect 18966 756 18972 808
rect 19024 756 19030 808
rect 19334 756 19340 808
rect 19392 796 19398 808
rect 19797 799 19855 805
rect 19797 796 19809 799
rect 19392 768 19809 796
rect 19392 756 19398 768
rect 19797 765 19809 768
rect 19843 765 19855 799
rect 19797 759 19855 765
rect 19889 799 19947 805
rect 19889 765 19901 799
rect 19935 796 19947 799
rect 20254 796 20260 808
rect 19935 768 20260 796
rect 19935 765 19947 768
rect 19889 759 19947 765
rect 20254 756 20260 768
rect 20312 756 20318 808
rect 20346 756 20352 808
rect 20404 796 20410 808
rect 20717 799 20775 805
rect 20717 796 20729 799
rect 20404 768 20729 796
rect 20404 756 20410 768
rect 20717 765 20729 768
rect 20763 765 20775 799
rect 20717 759 20775 765
rect 21542 756 21548 808
rect 21600 756 21606 808
rect 22370 756 22376 808
rect 22428 756 22434 808
rect 23566 756 23572 808
rect 23624 796 23630 808
rect 24121 799 24179 805
rect 24121 796 24133 799
rect 23624 768 24133 796
rect 23624 756 23630 768
rect 24121 765 24133 768
rect 24167 765 24179 799
rect 24121 759 24179 765
rect 24946 756 24952 808
rect 25004 756 25010 808
rect 15988 700 16528 728
rect 15988 688 15994 700
rect 552 570 27576 592
rect 552 518 7114 570
rect 7166 518 7178 570
rect 7230 518 7242 570
rect 7294 518 7306 570
rect 7358 518 7370 570
rect 7422 518 13830 570
rect 13882 518 13894 570
rect 13946 518 13958 570
rect 14010 518 14022 570
rect 14074 518 14086 570
rect 14138 518 20546 570
rect 20598 518 20610 570
rect 20662 518 20674 570
rect 20726 518 20738 570
rect 20790 518 20802 570
rect 20854 518 27262 570
rect 27314 518 27326 570
rect 27378 518 27390 570
rect 27442 518 27454 570
rect 27506 518 27518 570
rect 27570 518 27576 570
rect 552 496 27576 518
<< via1 >>
rect 13452 31152 13504 31204
rect 21088 31152 21140 31204
rect 19432 31084 19484 31136
rect 22744 31084 22796 31136
rect 7114 30982 7166 31034
rect 7178 30982 7230 31034
rect 7242 30982 7294 31034
rect 7306 30982 7358 31034
rect 7370 30982 7422 31034
rect 13830 30982 13882 31034
rect 13894 30982 13946 31034
rect 13958 30982 14010 31034
rect 14022 30982 14074 31034
rect 14086 30982 14138 31034
rect 20546 30982 20598 31034
rect 20610 30982 20662 31034
rect 20674 30982 20726 31034
rect 20738 30982 20790 31034
rect 20802 30982 20854 31034
rect 27262 30982 27314 31034
rect 27326 30982 27378 31034
rect 27390 30982 27442 31034
rect 27454 30982 27506 31034
rect 27518 30982 27570 31034
rect 1400 30880 1452 30932
rect 5816 30880 5868 30932
rect 7472 30880 7524 30932
rect 8760 30880 8812 30932
rect 2044 30787 2096 30796
rect 2044 30753 2073 30787
rect 2073 30753 2096 30787
rect 2044 30744 2096 30753
rect 3516 30744 3568 30796
rect 2320 30719 2372 30728
rect 2320 30685 2329 30719
rect 2329 30685 2363 30719
rect 2363 30685 2372 30719
rect 2320 30676 2372 30685
rect 9680 30787 9732 30796
rect 9680 30753 9689 30787
rect 9689 30753 9723 30787
rect 9723 30753 9732 30787
rect 9680 30744 9732 30753
rect 9864 30787 9916 30796
rect 9864 30753 9873 30787
rect 9873 30753 9907 30787
rect 9907 30753 9916 30787
rect 9864 30744 9916 30753
rect 10324 30744 10376 30796
rect 10232 30676 10284 30728
rect 11060 30608 11112 30660
rect 11704 30744 11756 30796
rect 11244 30719 11296 30728
rect 11244 30685 11253 30719
rect 11253 30685 11287 30719
rect 11287 30685 11296 30719
rect 11244 30676 11296 30685
rect 11796 30719 11848 30728
rect 11796 30685 11805 30719
rect 11805 30685 11839 30719
rect 11839 30685 11848 30719
rect 11796 30676 11848 30685
rect 12716 30744 12768 30796
rect 12440 30676 12492 30728
rect 16120 30880 16172 30932
rect 13176 30744 13228 30796
rect 14648 30744 14700 30796
rect 15292 30787 15344 30796
rect 15292 30753 15301 30787
rect 15301 30753 15335 30787
rect 15335 30753 15344 30787
rect 15292 30744 15344 30753
rect 17592 30812 17644 30864
rect 16764 30744 16816 30796
rect 14096 30719 14148 30728
rect 14096 30685 14105 30719
rect 14105 30685 14139 30719
rect 14139 30685 14148 30719
rect 14096 30676 14148 30685
rect 18052 30787 18104 30796
rect 18052 30753 18061 30787
rect 18061 30753 18095 30787
rect 18095 30753 18104 30787
rect 18052 30744 18104 30753
rect 19432 30787 19484 30796
rect 19432 30753 19441 30787
rect 19441 30753 19475 30787
rect 19475 30753 19484 30787
rect 19432 30744 19484 30753
rect 19616 30855 19668 30864
rect 19616 30821 19625 30855
rect 19625 30821 19659 30855
rect 19659 30821 19668 30855
rect 19616 30812 19668 30821
rect 19708 30812 19760 30864
rect 21088 30880 21140 30932
rect 23480 30880 23532 30932
rect 26424 30880 26476 30932
rect 3608 30540 3660 30592
rect 5908 30583 5960 30592
rect 5908 30549 5917 30583
rect 5917 30549 5951 30583
rect 5951 30549 5960 30583
rect 5908 30540 5960 30549
rect 7380 30583 7432 30592
rect 7380 30549 7389 30583
rect 7389 30549 7423 30583
rect 7423 30549 7432 30583
rect 7380 30540 7432 30549
rect 8484 30583 8536 30592
rect 8484 30549 8493 30583
rect 8493 30549 8527 30583
rect 8527 30549 8536 30583
rect 8484 30540 8536 30549
rect 8760 30540 8812 30592
rect 13636 30608 13688 30660
rect 19064 30676 19116 30728
rect 22008 30744 22060 30796
rect 20812 30719 20864 30728
rect 20812 30685 20821 30719
rect 20821 30685 20855 30719
rect 20855 30685 20864 30719
rect 20812 30676 20864 30685
rect 21732 30719 21784 30728
rect 21732 30685 21741 30719
rect 21741 30685 21775 30719
rect 21775 30685 21784 30719
rect 21732 30676 21784 30685
rect 22468 30719 22520 30728
rect 22468 30685 22477 30719
rect 22477 30685 22511 30719
rect 22511 30685 22520 30719
rect 22468 30676 22520 30685
rect 22744 30744 22796 30796
rect 23204 30676 23256 30728
rect 14556 30608 14608 30660
rect 12164 30583 12216 30592
rect 12164 30549 12173 30583
rect 12173 30549 12207 30583
rect 12207 30549 12216 30583
rect 12164 30540 12216 30549
rect 12624 30540 12676 30592
rect 13544 30583 13596 30592
rect 13544 30549 13553 30583
rect 13553 30549 13587 30583
rect 13587 30549 13596 30583
rect 13544 30540 13596 30549
rect 14648 30540 14700 30592
rect 18144 30608 18196 30660
rect 16396 30583 16448 30592
rect 16396 30549 16405 30583
rect 16405 30549 16439 30583
rect 16439 30549 16448 30583
rect 16396 30540 16448 30549
rect 17776 30583 17828 30592
rect 17776 30549 17785 30583
rect 17785 30549 17819 30583
rect 17819 30549 17828 30583
rect 17776 30540 17828 30549
rect 18236 30583 18288 30592
rect 18236 30549 18245 30583
rect 18245 30549 18279 30583
rect 18279 30549 18288 30583
rect 18236 30540 18288 30549
rect 19524 30540 19576 30592
rect 20076 30583 20128 30592
rect 20076 30549 20085 30583
rect 20085 30549 20119 30583
rect 20119 30549 20128 30583
rect 20076 30540 20128 30549
rect 21364 30583 21416 30592
rect 21364 30549 21373 30583
rect 21373 30549 21407 30583
rect 21407 30549 21416 30583
rect 21364 30540 21416 30549
rect 23020 30583 23072 30592
rect 23020 30549 23029 30583
rect 23029 30549 23063 30583
rect 23063 30549 23072 30583
rect 23020 30540 23072 30549
rect 23112 30583 23164 30592
rect 23112 30549 23121 30583
rect 23121 30549 23155 30583
rect 23155 30549 23164 30583
rect 23112 30540 23164 30549
rect 23572 30540 23624 30592
rect 26516 30583 26568 30592
rect 26516 30549 26525 30583
rect 26525 30549 26559 30583
rect 26559 30549 26568 30583
rect 26516 30540 26568 30549
rect 3756 30438 3808 30490
rect 3820 30438 3872 30490
rect 3884 30438 3936 30490
rect 3948 30438 4000 30490
rect 4012 30438 4064 30490
rect 10472 30438 10524 30490
rect 10536 30438 10588 30490
rect 10600 30438 10652 30490
rect 10664 30438 10716 30490
rect 10728 30438 10780 30490
rect 17188 30438 17240 30490
rect 17252 30438 17304 30490
rect 17316 30438 17368 30490
rect 17380 30438 17432 30490
rect 17444 30438 17496 30490
rect 23904 30438 23956 30490
rect 23968 30438 24020 30490
rect 24032 30438 24084 30490
rect 24096 30438 24148 30490
rect 24160 30438 24212 30490
rect 2872 30268 2924 30320
rect 5908 30336 5960 30388
rect 13268 30336 13320 30388
rect 2320 30132 2372 30184
rect 4528 30132 4580 30184
rect 5908 30175 5960 30184
rect 5908 30141 5917 30175
rect 5917 30141 5951 30175
rect 5951 30141 5960 30175
rect 5908 30132 5960 30141
rect 7380 30268 7432 30320
rect 1860 30107 1912 30116
rect 1860 30073 1894 30107
rect 1894 30073 1912 30107
rect 1860 30064 1912 30073
rect 3608 30107 3660 30116
rect 3608 30073 3642 30107
rect 3642 30073 3660 30107
rect 3608 30064 3660 30073
rect 1768 29996 1820 30048
rect 5448 30064 5500 30116
rect 6828 30132 6880 30184
rect 5172 29996 5224 30048
rect 5540 29996 5592 30048
rect 5816 29996 5868 30048
rect 7472 30064 7524 30116
rect 12992 30311 13044 30320
rect 12992 30277 13001 30311
rect 13001 30277 13035 30311
rect 13035 30277 13044 30311
rect 14096 30336 14148 30388
rect 15660 30336 15712 30388
rect 16396 30336 16448 30388
rect 20812 30336 20864 30388
rect 22468 30336 22520 30388
rect 22652 30379 22704 30388
rect 22652 30345 22661 30379
rect 22661 30345 22695 30379
rect 22695 30345 22704 30379
rect 22652 30336 22704 30345
rect 26516 30336 26568 30388
rect 12992 30268 13044 30277
rect 17040 30311 17092 30320
rect 17040 30277 17049 30311
rect 17049 30277 17083 30311
rect 17083 30277 17092 30311
rect 17040 30268 17092 30277
rect 12624 30200 12676 30252
rect 12808 30200 12860 30252
rect 10968 30132 11020 30184
rect 13084 30175 13136 30184
rect 13084 30141 13093 30175
rect 13093 30141 13127 30175
rect 13127 30141 13136 30175
rect 13084 30132 13136 30141
rect 13544 30132 13596 30184
rect 14556 30132 14608 30184
rect 14648 30132 14700 30184
rect 16948 30200 17000 30252
rect 17316 30200 17368 30252
rect 21272 30243 21324 30252
rect 21272 30209 21281 30243
rect 21281 30209 21315 30243
rect 21315 30209 21324 30243
rect 21272 30200 21324 30209
rect 6736 29996 6788 30048
rect 8024 30064 8076 30116
rect 7656 30039 7708 30048
rect 7656 30005 7665 30039
rect 7665 30005 7699 30039
rect 7699 30005 7708 30039
rect 7656 29996 7708 30005
rect 8668 30064 8720 30116
rect 11060 30064 11112 30116
rect 13728 30064 13780 30116
rect 14280 30064 14332 30116
rect 8760 29996 8812 30048
rect 9588 29996 9640 30048
rect 10232 29996 10284 30048
rect 11152 29996 11204 30048
rect 14648 29996 14700 30048
rect 15108 30064 15160 30116
rect 15568 30064 15620 30116
rect 16120 29996 16172 30048
rect 16396 30175 16448 30184
rect 16396 30141 16405 30175
rect 16405 30141 16439 30175
rect 16439 30141 16448 30175
rect 16396 30132 16448 30141
rect 18144 30175 18196 30184
rect 18144 30141 18162 30175
rect 18162 30141 18196 30175
rect 18144 30132 18196 30141
rect 19432 30132 19484 30184
rect 16580 30064 16632 30116
rect 19524 30064 19576 30116
rect 20444 30132 20496 30184
rect 22744 30200 22796 30252
rect 22652 30132 22704 30184
rect 23020 30200 23072 30252
rect 20996 30039 21048 30048
rect 20996 30005 21005 30039
rect 21005 30005 21039 30039
rect 21039 30005 21048 30039
rect 20996 29996 21048 30005
rect 23020 30107 23072 30116
rect 23020 30073 23029 30107
rect 23029 30073 23063 30107
rect 23063 30073 23072 30107
rect 23020 30064 23072 30073
rect 23204 30064 23256 30116
rect 23480 30107 23532 30116
rect 23480 30073 23489 30107
rect 23489 30073 23523 30107
rect 23523 30073 23532 30107
rect 23480 30064 23532 30073
rect 24400 30107 24452 30116
rect 24400 30073 24409 30107
rect 24409 30073 24443 30107
rect 24443 30073 24452 30107
rect 24400 30064 24452 30073
rect 23664 29996 23716 30048
rect 23940 29996 23992 30048
rect 24216 30039 24268 30048
rect 24216 30005 24225 30039
rect 24225 30005 24259 30039
rect 24259 30005 24268 30039
rect 24216 29996 24268 30005
rect 24492 29996 24544 30048
rect 24860 30039 24912 30048
rect 24860 30005 24869 30039
rect 24869 30005 24903 30039
rect 24903 30005 24912 30039
rect 24860 29996 24912 30005
rect 25228 29996 25280 30048
rect 7114 29894 7166 29946
rect 7178 29894 7230 29946
rect 7242 29894 7294 29946
rect 7306 29894 7358 29946
rect 7370 29894 7422 29946
rect 13830 29894 13882 29946
rect 13894 29894 13946 29946
rect 13958 29894 14010 29946
rect 14022 29894 14074 29946
rect 14086 29894 14138 29946
rect 20546 29894 20598 29946
rect 20610 29894 20662 29946
rect 20674 29894 20726 29946
rect 20738 29894 20790 29946
rect 20802 29894 20854 29946
rect 27262 29894 27314 29946
rect 27326 29894 27378 29946
rect 27390 29894 27442 29946
rect 27454 29894 27506 29946
rect 27518 29894 27570 29946
rect 3516 29792 3568 29844
rect 4160 29724 4212 29776
rect 2044 29656 2096 29708
rect 3608 29656 3660 29708
rect 5816 29792 5868 29844
rect 5908 29792 5960 29844
rect 6736 29724 6788 29776
rect 7472 29792 7524 29844
rect 7932 29792 7984 29844
rect 7840 29724 7892 29776
rect 1860 29588 1912 29640
rect 5080 29631 5132 29640
rect 5080 29597 5089 29631
rect 5089 29597 5123 29631
rect 5123 29597 5132 29631
rect 5080 29588 5132 29597
rect 4252 29452 4304 29504
rect 4344 29452 4396 29504
rect 4804 29452 4856 29504
rect 4896 29495 4948 29504
rect 4896 29461 4905 29495
rect 4905 29461 4939 29495
rect 4939 29461 4948 29495
rect 4896 29452 4948 29461
rect 6368 29588 6420 29640
rect 6920 29699 6972 29708
rect 6920 29665 6929 29699
rect 6929 29665 6963 29699
rect 6963 29665 6972 29699
rect 6920 29656 6972 29665
rect 7104 29656 7156 29708
rect 7748 29699 7800 29708
rect 7748 29665 7782 29699
rect 7782 29665 7800 29699
rect 7748 29656 7800 29665
rect 8300 29699 8352 29708
rect 8300 29665 8309 29699
rect 8309 29665 8343 29699
rect 8343 29665 8352 29699
rect 9588 29724 9640 29776
rect 8300 29656 8352 29665
rect 8760 29699 8812 29708
rect 8760 29665 8769 29699
rect 8769 29665 8803 29699
rect 8803 29665 8812 29699
rect 8760 29656 8812 29665
rect 11796 29792 11848 29844
rect 12716 29835 12768 29844
rect 12716 29801 12725 29835
rect 12725 29801 12759 29835
rect 12759 29801 12768 29835
rect 12716 29792 12768 29801
rect 7012 29588 7064 29640
rect 7196 29631 7248 29640
rect 7196 29597 7205 29631
rect 7205 29597 7239 29631
rect 7239 29597 7248 29631
rect 7196 29588 7248 29597
rect 7656 29588 7708 29640
rect 7104 29452 7156 29504
rect 7748 29520 7800 29572
rect 9864 29724 9916 29776
rect 7564 29452 7616 29504
rect 8760 29452 8812 29504
rect 9404 29495 9456 29504
rect 9404 29461 9413 29495
rect 9413 29461 9447 29495
rect 9447 29461 9456 29495
rect 9404 29452 9456 29461
rect 10232 29699 10284 29708
rect 10232 29665 10241 29699
rect 10241 29665 10275 29699
rect 10275 29665 10284 29699
rect 10232 29656 10284 29665
rect 10324 29699 10376 29708
rect 10324 29665 10333 29699
rect 10333 29665 10367 29699
rect 10367 29665 10376 29699
rect 10324 29656 10376 29665
rect 12440 29767 12492 29776
rect 12440 29733 12449 29767
rect 12449 29733 12483 29767
rect 12483 29733 12492 29767
rect 12440 29724 12492 29733
rect 12992 29792 13044 29844
rect 14280 29792 14332 29844
rect 15016 29792 15068 29844
rect 15292 29835 15344 29844
rect 15292 29801 15301 29835
rect 15301 29801 15335 29835
rect 15335 29801 15344 29835
rect 15292 29792 15344 29801
rect 16120 29792 16172 29844
rect 14464 29767 14516 29776
rect 14464 29733 14491 29767
rect 14491 29733 14516 29767
rect 14464 29724 14516 29733
rect 15384 29724 15436 29776
rect 15568 29724 15620 29776
rect 13084 29656 13136 29708
rect 10968 29631 11020 29640
rect 10968 29597 10977 29631
rect 10977 29597 11011 29631
rect 11011 29597 11020 29631
rect 10968 29588 11020 29597
rect 12164 29588 12216 29640
rect 12440 29588 12492 29640
rect 13544 29588 13596 29640
rect 13360 29563 13412 29572
rect 13360 29529 13369 29563
rect 13369 29529 13403 29563
rect 13403 29529 13412 29563
rect 13360 29520 13412 29529
rect 13452 29520 13504 29572
rect 15568 29588 15620 29640
rect 16212 29724 16264 29776
rect 16488 29767 16540 29776
rect 16488 29733 16497 29767
rect 16497 29733 16531 29767
rect 16531 29733 16540 29767
rect 16488 29724 16540 29733
rect 16764 29835 16816 29844
rect 16764 29801 16773 29835
rect 16773 29801 16807 29835
rect 16807 29801 16816 29835
rect 16764 29792 16816 29801
rect 17040 29792 17092 29844
rect 20628 29792 20680 29844
rect 16948 29767 17000 29776
rect 16948 29733 16957 29767
rect 16957 29733 16991 29767
rect 16991 29733 17000 29767
rect 16948 29724 17000 29733
rect 18236 29724 18288 29776
rect 18972 29724 19024 29776
rect 21548 29724 21600 29776
rect 23848 29792 23900 29844
rect 14464 29520 14516 29572
rect 14648 29520 14700 29572
rect 11244 29452 11296 29504
rect 12992 29452 13044 29504
rect 13084 29495 13136 29504
rect 13084 29461 13093 29495
rect 13093 29461 13127 29495
rect 13127 29461 13136 29495
rect 13084 29452 13136 29461
rect 13636 29452 13688 29504
rect 15660 29452 15712 29504
rect 17316 29656 17368 29708
rect 19524 29656 19576 29708
rect 19708 29699 19760 29708
rect 19708 29665 19742 29699
rect 19742 29665 19760 29699
rect 19708 29656 19760 29665
rect 22928 29699 22980 29708
rect 16120 29563 16172 29572
rect 16120 29529 16129 29563
rect 16129 29529 16163 29563
rect 16163 29529 16172 29563
rect 16120 29520 16172 29529
rect 17040 29520 17092 29572
rect 15936 29495 15988 29504
rect 15936 29461 15945 29495
rect 15945 29461 15979 29495
rect 15979 29461 15988 29495
rect 15936 29452 15988 29461
rect 16672 29495 16724 29504
rect 16672 29461 16681 29495
rect 16681 29461 16715 29495
rect 16715 29461 16724 29495
rect 16672 29452 16724 29461
rect 16764 29452 16816 29504
rect 19248 29588 19300 29640
rect 22652 29631 22704 29640
rect 22652 29597 22661 29631
rect 22661 29597 22695 29631
rect 22695 29597 22704 29631
rect 22652 29588 22704 29597
rect 22928 29665 22934 29699
rect 22934 29665 22968 29699
rect 22968 29665 22980 29699
rect 22928 29656 22980 29665
rect 23388 29699 23440 29708
rect 23388 29665 23397 29699
rect 23397 29665 23431 29699
rect 23431 29665 23440 29699
rect 23388 29656 23440 29665
rect 24400 29792 24452 29844
rect 24860 29792 24912 29844
rect 24676 29724 24728 29776
rect 23112 29588 23164 29640
rect 23756 29631 23808 29640
rect 23756 29597 23765 29631
rect 23765 29597 23799 29631
rect 23799 29597 23808 29631
rect 23756 29588 23808 29597
rect 25964 29656 26016 29708
rect 17592 29452 17644 29504
rect 18144 29452 18196 29504
rect 19156 29452 19208 29504
rect 19616 29452 19668 29504
rect 20076 29452 20128 29504
rect 20628 29452 20680 29504
rect 21732 29452 21784 29504
rect 22836 29452 22888 29504
rect 23296 29495 23348 29504
rect 23296 29461 23305 29495
rect 23305 29461 23339 29495
rect 23339 29461 23348 29495
rect 23296 29452 23348 29461
rect 24584 29520 24636 29572
rect 23756 29452 23808 29504
rect 24216 29495 24268 29504
rect 24216 29461 24225 29495
rect 24225 29461 24259 29495
rect 24259 29461 24268 29495
rect 24216 29452 24268 29461
rect 25228 29495 25280 29504
rect 25228 29461 25237 29495
rect 25237 29461 25271 29495
rect 25271 29461 25280 29495
rect 25228 29452 25280 29461
rect 3756 29350 3808 29402
rect 3820 29350 3872 29402
rect 3884 29350 3936 29402
rect 3948 29350 4000 29402
rect 4012 29350 4064 29402
rect 10472 29350 10524 29402
rect 10536 29350 10588 29402
rect 10600 29350 10652 29402
rect 10664 29350 10716 29402
rect 10728 29350 10780 29402
rect 17188 29350 17240 29402
rect 17252 29350 17304 29402
rect 17316 29350 17368 29402
rect 17380 29350 17432 29402
rect 17444 29350 17496 29402
rect 23904 29350 23956 29402
rect 23968 29350 24020 29402
rect 24032 29350 24084 29402
rect 24096 29350 24148 29402
rect 24160 29350 24212 29402
rect 3608 29248 3660 29300
rect 4160 29248 4212 29300
rect 4896 29248 4948 29300
rect 5080 29248 5132 29300
rect 6460 29291 6512 29300
rect 6460 29257 6469 29291
rect 6469 29257 6503 29291
rect 6503 29257 6512 29291
rect 6460 29248 6512 29257
rect 6920 29291 6972 29300
rect 6920 29257 6929 29291
rect 6929 29257 6963 29291
rect 6963 29257 6972 29291
rect 6920 29248 6972 29257
rect 7196 29248 7248 29300
rect 7656 29248 7708 29300
rect 8484 29248 8536 29300
rect 8668 29291 8720 29300
rect 8668 29257 8677 29291
rect 8677 29257 8711 29291
rect 8711 29257 8720 29291
rect 8668 29248 8720 29257
rect 9404 29248 9456 29300
rect 9496 29248 9548 29300
rect 9680 29248 9732 29300
rect 10232 29248 10284 29300
rect 10324 29248 10376 29300
rect 11152 29248 11204 29300
rect 13268 29248 13320 29300
rect 13544 29248 13596 29300
rect 13728 29248 13780 29300
rect 3056 29044 3108 29096
rect 3976 28976 4028 29028
rect 4620 29087 4672 29096
rect 4620 29053 4629 29087
rect 4629 29053 4663 29087
rect 4663 29053 4672 29087
rect 4620 29044 4672 29053
rect 4804 29019 4856 29028
rect 4804 28985 4813 29019
rect 4813 28985 4847 29019
rect 4847 28985 4856 29019
rect 4804 28976 4856 28985
rect 5908 29180 5960 29232
rect 5448 29044 5500 29096
rect 6368 29087 6420 29096
rect 6368 29053 6377 29087
rect 6377 29053 6411 29087
rect 6411 29053 6420 29087
rect 6368 29044 6420 29053
rect 6644 29087 6696 29096
rect 6644 29053 6653 29087
rect 6653 29053 6687 29087
rect 6687 29053 6696 29087
rect 6644 29044 6696 29053
rect 8300 29180 8352 29232
rect 7012 28951 7064 28960
rect 7012 28917 7021 28951
rect 7021 28917 7055 28951
rect 7055 28917 7064 28951
rect 7012 28908 7064 28917
rect 7472 28976 7524 29028
rect 7932 29087 7984 29096
rect 7932 29053 7941 29087
rect 7941 29053 7975 29087
rect 7975 29053 7984 29087
rect 7932 29044 7984 29053
rect 8024 29044 8076 29096
rect 8760 29044 8812 29096
rect 7656 29019 7708 29028
rect 7656 28985 7665 29019
rect 7665 28985 7699 29019
rect 7699 28985 7708 29019
rect 7656 28976 7708 28985
rect 8392 28976 8444 29028
rect 8944 29019 8996 29028
rect 8944 28985 8953 29019
rect 8953 28985 8987 29019
rect 8987 28985 8996 29019
rect 8944 28976 8996 28985
rect 12440 29180 12492 29232
rect 7748 28908 7800 28960
rect 11612 28976 11664 29028
rect 11980 29019 12032 29028
rect 11980 28985 11989 29019
rect 11989 28985 12023 29019
rect 12023 28985 12032 29019
rect 11980 28976 12032 28985
rect 12072 29019 12124 29028
rect 12072 28985 12081 29019
rect 12081 28985 12115 29019
rect 12115 28985 12124 29019
rect 12072 28976 12124 28985
rect 9496 28908 9548 28960
rect 9680 28908 9732 28960
rect 11704 28951 11756 28960
rect 11704 28917 11713 28951
rect 11713 28917 11747 28951
rect 11747 28917 11756 28951
rect 11704 28908 11756 28917
rect 12624 28908 12676 28960
rect 16580 29248 16632 29300
rect 16948 29248 17000 29300
rect 17132 29291 17184 29300
rect 17132 29257 17141 29291
rect 17141 29257 17175 29291
rect 17175 29257 17184 29291
rect 17132 29248 17184 29257
rect 18052 29248 18104 29300
rect 13360 29112 13412 29164
rect 14464 29044 14516 29096
rect 15016 29112 15068 29164
rect 15108 29087 15160 29096
rect 15108 29053 15117 29087
rect 15117 29053 15151 29087
rect 15151 29053 15160 29087
rect 15108 29044 15160 29053
rect 16120 29180 16172 29232
rect 16672 29180 16724 29232
rect 15752 29087 15804 29096
rect 15752 29053 15761 29087
rect 15761 29053 15795 29087
rect 15795 29053 15804 29087
rect 15752 29044 15804 29053
rect 17040 29044 17092 29096
rect 15936 28976 15988 29028
rect 13452 28908 13504 28960
rect 13544 28908 13596 28960
rect 15568 28951 15620 28960
rect 15568 28917 15577 28951
rect 15577 28917 15611 28951
rect 15611 28917 15620 28951
rect 15568 28908 15620 28917
rect 15844 28951 15896 28960
rect 15844 28917 15853 28951
rect 15853 28917 15887 28951
rect 15887 28917 15896 28951
rect 15844 28908 15896 28917
rect 16396 28908 16448 28960
rect 16764 28908 16816 28960
rect 17592 29019 17644 29028
rect 17592 28985 17601 29019
rect 17601 28985 17635 29019
rect 17635 28985 17644 29019
rect 17592 28976 17644 28985
rect 18144 29087 18196 29096
rect 18144 29053 18153 29087
rect 18153 29053 18187 29087
rect 18187 29053 18196 29087
rect 18144 29044 18196 29053
rect 19340 29248 19392 29300
rect 19708 29248 19760 29300
rect 19616 29180 19668 29232
rect 21548 29180 21600 29232
rect 23020 29248 23072 29300
rect 23756 29248 23808 29300
rect 24308 29248 24360 29300
rect 24400 29248 24452 29300
rect 18696 29087 18748 29096
rect 18696 29053 18705 29087
rect 18705 29053 18739 29087
rect 18739 29053 18748 29087
rect 18696 29044 18748 29053
rect 20628 29155 20680 29164
rect 20628 29121 20637 29155
rect 20637 29121 20671 29155
rect 20671 29121 20680 29155
rect 20628 29112 20680 29121
rect 19156 29087 19208 29096
rect 19156 29053 19165 29087
rect 19165 29053 19199 29087
rect 19199 29053 19208 29087
rect 19156 29044 19208 29053
rect 19248 29087 19300 29096
rect 19248 29053 19257 29087
rect 19257 29053 19291 29087
rect 19291 29053 19300 29087
rect 19248 29044 19300 29053
rect 19340 29087 19392 29096
rect 19340 29053 19349 29087
rect 19349 29053 19383 29087
rect 19383 29053 19392 29087
rect 19340 29044 19392 29053
rect 19800 29044 19852 29096
rect 21180 29044 21232 29096
rect 21640 29087 21692 29096
rect 21640 29053 21649 29087
rect 21649 29053 21683 29087
rect 21683 29053 21692 29087
rect 21640 29044 21692 29053
rect 23296 29044 23348 29096
rect 24308 29112 24360 29164
rect 24584 29223 24636 29232
rect 24584 29189 24593 29223
rect 24593 29189 24627 29223
rect 24627 29189 24636 29223
rect 24584 29180 24636 29189
rect 18236 29019 18288 29028
rect 18236 28985 18245 29019
rect 18245 28985 18279 29019
rect 18279 28985 18288 29019
rect 18236 28976 18288 28985
rect 24492 29044 24544 29096
rect 24768 29044 24820 29096
rect 25320 29044 25372 29096
rect 26424 29019 26476 29028
rect 26424 28985 26442 29019
rect 26442 28985 26476 29019
rect 26424 28976 26476 28985
rect 18880 28951 18932 28960
rect 18880 28917 18889 28951
rect 18889 28917 18923 28951
rect 18923 28917 18932 28951
rect 18880 28908 18932 28917
rect 21732 28908 21784 28960
rect 24400 28951 24452 28960
rect 24400 28917 24409 28951
rect 24409 28917 24443 28951
rect 24443 28917 24452 28951
rect 24400 28908 24452 28917
rect 24492 28951 24544 28960
rect 24492 28917 24501 28951
rect 24501 28917 24535 28951
rect 24535 28917 24544 28951
rect 24492 28908 24544 28917
rect 26240 28908 26292 28960
rect 7114 28806 7166 28858
rect 7178 28806 7230 28858
rect 7242 28806 7294 28858
rect 7306 28806 7358 28858
rect 7370 28806 7422 28858
rect 13830 28806 13882 28858
rect 13894 28806 13946 28858
rect 13958 28806 14010 28858
rect 14022 28806 14074 28858
rect 14086 28806 14138 28858
rect 20546 28806 20598 28858
rect 20610 28806 20662 28858
rect 20674 28806 20726 28858
rect 20738 28806 20790 28858
rect 20802 28806 20854 28858
rect 27262 28806 27314 28858
rect 27326 28806 27378 28858
rect 27390 28806 27442 28858
rect 27454 28806 27506 28858
rect 27518 28806 27570 28858
rect 3240 28747 3292 28756
rect 3240 28713 3249 28747
rect 3249 28713 3283 28747
rect 3283 28713 3292 28747
rect 3240 28704 3292 28713
rect 2136 28611 2188 28620
rect 2136 28577 2170 28611
rect 2170 28577 2188 28611
rect 2136 28568 2188 28577
rect 1860 28543 1912 28552
rect 1860 28509 1869 28543
rect 1869 28509 1903 28543
rect 1903 28509 1912 28543
rect 1860 28500 1912 28509
rect 3608 28611 3660 28620
rect 3608 28577 3617 28611
rect 3617 28577 3651 28611
rect 3651 28577 3660 28611
rect 3608 28568 3660 28577
rect 4252 28679 4304 28688
rect 4252 28645 4263 28679
rect 4263 28645 4304 28679
rect 4252 28636 4304 28645
rect 4436 28679 4488 28688
rect 4436 28645 4445 28679
rect 4445 28645 4479 28679
rect 4479 28645 4488 28679
rect 4436 28636 4488 28645
rect 4804 28636 4856 28688
rect 6644 28704 6696 28756
rect 7288 28704 7340 28756
rect 7472 28704 7524 28756
rect 7564 28704 7616 28756
rect 5908 28568 5960 28620
rect 7196 28568 7248 28620
rect 7564 28611 7616 28620
rect 7564 28577 7573 28611
rect 7573 28577 7607 28611
rect 7607 28577 7616 28611
rect 7564 28568 7616 28577
rect 7748 28611 7800 28620
rect 7748 28577 7757 28611
rect 7757 28577 7791 28611
rect 7791 28577 7800 28611
rect 7748 28568 7800 28577
rect 8944 28611 8996 28620
rect 8944 28577 8978 28611
rect 8978 28577 8996 28611
rect 8944 28568 8996 28577
rect 15384 28704 15436 28756
rect 11704 28636 11756 28688
rect 14556 28636 14608 28688
rect 15936 28704 15988 28756
rect 18696 28704 18748 28756
rect 12716 28568 12768 28620
rect 4252 28500 4304 28552
rect 6828 28500 6880 28552
rect 2228 28364 2280 28416
rect 2780 28364 2832 28416
rect 3424 28364 3476 28416
rect 6920 28432 6972 28484
rect 7932 28432 7984 28484
rect 10968 28543 11020 28552
rect 10968 28509 10977 28543
rect 10977 28509 11011 28543
rect 11011 28509 11020 28543
rect 10968 28500 11020 28509
rect 12808 28543 12860 28552
rect 12808 28509 12817 28543
rect 12817 28509 12851 28543
rect 12851 28509 12860 28543
rect 12808 28500 12860 28509
rect 15660 28568 15712 28620
rect 15936 28568 15988 28620
rect 16396 28568 16448 28620
rect 16672 28636 16724 28688
rect 18880 28636 18932 28688
rect 17592 28568 17644 28620
rect 16580 28500 16632 28552
rect 9680 28364 9732 28416
rect 10140 28407 10192 28416
rect 10140 28373 10149 28407
rect 10149 28373 10183 28407
rect 10183 28373 10192 28407
rect 10140 28364 10192 28373
rect 13544 28364 13596 28416
rect 14280 28407 14332 28416
rect 14280 28373 14289 28407
rect 14289 28373 14323 28407
rect 14323 28373 14332 28407
rect 14280 28364 14332 28373
rect 15292 28364 15344 28416
rect 16672 28475 16724 28484
rect 16672 28441 16681 28475
rect 16681 28441 16715 28475
rect 16715 28441 16724 28475
rect 21732 28636 21784 28688
rect 19616 28568 19668 28620
rect 21272 28611 21324 28620
rect 21272 28577 21281 28611
rect 21281 28577 21315 28611
rect 21315 28577 21324 28611
rect 21272 28568 21324 28577
rect 23112 28611 23164 28620
rect 23112 28577 23121 28611
rect 23121 28577 23155 28611
rect 23155 28577 23164 28611
rect 23112 28568 23164 28577
rect 25320 28704 25372 28756
rect 25688 28747 25740 28756
rect 25688 28713 25697 28747
rect 25697 28713 25731 28747
rect 25731 28713 25740 28747
rect 25688 28704 25740 28713
rect 25044 28679 25096 28688
rect 25044 28645 25071 28679
rect 25071 28645 25096 28679
rect 25044 28636 25096 28645
rect 25228 28679 25280 28688
rect 25228 28645 25237 28679
rect 25237 28645 25271 28679
rect 25271 28645 25280 28679
rect 25228 28636 25280 28645
rect 19524 28543 19576 28552
rect 19524 28509 19533 28543
rect 19533 28509 19567 28543
rect 19567 28509 19576 28543
rect 19524 28500 19576 28509
rect 25596 28611 25648 28620
rect 25596 28577 25605 28611
rect 25605 28577 25639 28611
rect 25639 28577 25648 28611
rect 25596 28568 25648 28577
rect 25872 28611 25924 28620
rect 25872 28577 25881 28611
rect 25881 28577 25915 28611
rect 25915 28577 25924 28611
rect 25872 28568 25924 28577
rect 26424 28568 26476 28620
rect 16672 28432 16724 28441
rect 15660 28407 15712 28416
rect 15660 28373 15669 28407
rect 15669 28373 15703 28407
rect 15703 28373 15712 28407
rect 15660 28364 15712 28373
rect 15752 28364 15804 28416
rect 16120 28364 16172 28416
rect 16764 28364 16816 28416
rect 17132 28364 17184 28416
rect 21180 28364 21232 28416
rect 22008 28364 22060 28416
rect 22836 28364 22888 28416
rect 22928 28407 22980 28416
rect 22928 28373 22937 28407
rect 22937 28373 22971 28407
rect 22971 28373 22980 28407
rect 22928 28364 22980 28373
rect 24584 28364 24636 28416
rect 25044 28407 25096 28416
rect 25044 28373 25053 28407
rect 25053 28373 25087 28407
rect 25087 28373 25096 28407
rect 25044 28364 25096 28373
rect 25136 28364 25188 28416
rect 25780 28364 25832 28416
rect 26056 28407 26108 28416
rect 26056 28373 26065 28407
rect 26065 28373 26099 28407
rect 26099 28373 26108 28407
rect 26056 28364 26108 28373
rect 3756 28262 3808 28314
rect 3820 28262 3872 28314
rect 3884 28262 3936 28314
rect 3948 28262 4000 28314
rect 4012 28262 4064 28314
rect 10472 28262 10524 28314
rect 10536 28262 10588 28314
rect 10600 28262 10652 28314
rect 10664 28262 10716 28314
rect 10728 28262 10780 28314
rect 17188 28262 17240 28314
rect 17252 28262 17304 28314
rect 17316 28262 17368 28314
rect 17380 28262 17432 28314
rect 17444 28262 17496 28314
rect 23904 28262 23956 28314
rect 23968 28262 24020 28314
rect 24032 28262 24084 28314
rect 24096 28262 24148 28314
rect 24160 28262 24212 28314
rect 2136 28160 2188 28212
rect 3424 28160 3476 28212
rect 4528 28203 4580 28212
rect 4528 28169 4537 28203
rect 4537 28169 4571 28203
rect 4571 28169 4580 28203
rect 4528 28160 4580 28169
rect 7012 28160 7064 28212
rect 3056 28135 3108 28144
rect 3056 28101 3065 28135
rect 3065 28101 3099 28135
rect 3099 28101 3108 28135
rect 3056 28092 3108 28101
rect 3240 28092 3292 28144
rect 6552 28092 6604 28144
rect 2872 27956 2924 28008
rect 8760 28024 8812 28076
rect 2780 27931 2832 27940
rect 2780 27897 2789 27931
rect 2789 27897 2823 27931
rect 2823 27897 2832 27931
rect 2780 27888 2832 27897
rect 2504 27863 2556 27872
rect 2504 27829 2513 27863
rect 2513 27829 2547 27863
rect 2547 27829 2556 27863
rect 2504 27820 2556 27829
rect 3240 27931 3292 27940
rect 3240 27897 3249 27931
rect 3249 27897 3283 27931
rect 3283 27897 3292 27931
rect 3240 27888 3292 27897
rect 3608 27888 3660 27940
rect 6736 27999 6788 28008
rect 6736 27965 6745 27999
rect 6745 27965 6779 27999
rect 6779 27965 6788 27999
rect 6736 27956 6788 27965
rect 7564 27888 7616 27940
rect 7840 27888 7892 27940
rect 8024 27999 8076 28008
rect 8024 27965 8033 27999
rect 8033 27965 8067 27999
rect 8067 27965 8076 27999
rect 8024 27956 8076 27965
rect 8852 27956 8904 28008
rect 9220 28024 9272 28076
rect 9680 28160 9732 28212
rect 12716 28203 12768 28212
rect 12716 28169 12725 28203
rect 12725 28169 12759 28203
rect 12759 28169 12768 28203
rect 12716 28160 12768 28169
rect 13452 28160 13504 28212
rect 14280 28160 14332 28212
rect 15844 28160 15896 28212
rect 16580 28160 16632 28212
rect 16672 28160 16724 28212
rect 21640 28203 21692 28212
rect 21640 28169 21649 28203
rect 21649 28169 21683 28203
rect 21683 28169 21692 28203
rect 21640 28160 21692 28169
rect 22192 28160 22244 28212
rect 10876 28135 10928 28144
rect 10876 28101 10885 28135
rect 10885 28101 10919 28135
rect 10919 28101 10928 28135
rect 10876 28092 10928 28101
rect 8392 27888 8444 27940
rect 9404 27999 9456 28008
rect 9404 27965 9413 27999
rect 9413 27965 9447 27999
rect 9447 27965 9456 27999
rect 9404 27956 9456 27965
rect 11704 27956 11756 28008
rect 12532 27999 12584 28008
rect 12532 27965 12541 27999
rect 12541 27965 12575 27999
rect 12575 27965 12584 27999
rect 12532 27956 12584 27965
rect 12624 27956 12676 28008
rect 13544 27999 13596 28008
rect 13544 27965 13553 27999
rect 13553 27965 13587 27999
rect 13587 27965 13596 27999
rect 13544 27956 13596 27965
rect 14556 27956 14608 28008
rect 15292 28092 15344 28144
rect 9772 27931 9824 27940
rect 9772 27897 9806 27931
rect 9806 27897 9824 27931
rect 9772 27888 9824 27897
rect 7748 27863 7800 27872
rect 7748 27829 7757 27863
rect 7757 27829 7791 27863
rect 7791 27829 7800 27863
rect 7748 27820 7800 27829
rect 7932 27820 7984 27872
rect 8576 27863 8628 27872
rect 8576 27829 8585 27863
rect 8585 27829 8619 27863
rect 8619 27829 8628 27863
rect 8576 27820 8628 27829
rect 9864 27820 9916 27872
rect 10968 27863 11020 27872
rect 10968 27829 10977 27863
rect 10977 27829 11011 27863
rect 11011 27829 11020 27863
rect 10968 27820 11020 27829
rect 11520 27820 11572 27872
rect 13084 27931 13136 27940
rect 13084 27897 13093 27931
rect 13093 27897 13127 27931
rect 13127 27897 13136 27931
rect 13084 27888 13136 27897
rect 15016 27999 15068 28008
rect 15016 27965 15025 27999
rect 15025 27965 15059 27999
rect 15059 27965 15068 27999
rect 16948 28024 17000 28076
rect 21272 28024 21324 28076
rect 22652 28160 22704 28212
rect 23296 28160 23348 28212
rect 25044 28160 25096 28212
rect 25228 28092 25280 28144
rect 25872 28160 25924 28212
rect 26056 28160 26108 28212
rect 15016 27956 15068 27965
rect 15108 27888 15160 27940
rect 14832 27820 14884 27872
rect 15384 27863 15436 27872
rect 15384 27829 15393 27863
rect 15393 27829 15427 27863
rect 15427 27829 15436 27863
rect 15384 27820 15436 27829
rect 15476 27863 15528 27872
rect 15476 27829 15485 27863
rect 15485 27829 15519 27863
rect 15519 27829 15528 27863
rect 15476 27820 15528 27829
rect 15568 27820 15620 27872
rect 16396 27820 16448 27872
rect 17132 27999 17184 28008
rect 17132 27965 17141 27999
rect 17141 27965 17175 27999
rect 17175 27965 17184 27999
rect 17132 27956 17184 27965
rect 17776 27956 17828 28008
rect 22376 27956 22428 28008
rect 23664 27956 23716 28008
rect 16672 27820 16724 27872
rect 17224 27820 17276 27872
rect 18328 27820 18380 27872
rect 18512 27863 18564 27872
rect 18512 27829 18521 27863
rect 18521 27829 18555 27863
rect 18555 27829 18564 27863
rect 18512 27820 18564 27829
rect 19524 27820 19576 27872
rect 22928 27888 22980 27940
rect 23572 27888 23624 27940
rect 24216 27956 24268 28008
rect 24400 27999 24452 28008
rect 24400 27965 24409 27999
rect 24409 27965 24443 27999
rect 24443 27965 24452 27999
rect 24400 27956 24452 27965
rect 24492 27956 24544 28008
rect 25228 27956 25280 28008
rect 21824 27863 21876 27872
rect 21824 27829 21833 27863
rect 21833 27829 21867 27863
rect 21867 27829 21876 27863
rect 21824 27820 21876 27829
rect 22192 27820 22244 27872
rect 22652 27820 22704 27872
rect 23296 27820 23348 27872
rect 23388 27820 23440 27872
rect 24584 27931 24636 27940
rect 24584 27897 24593 27931
rect 24593 27897 24627 27931
rect 24627 27897 24636 27931
rect 24584 27888 24636 27897
rect 24768 27931 24820 27940
rect 24768 27897 24777 27931
rect 24777 27897 24811 27931
rect 24811 27897 24820 27931
rect 24768 27888 24820 27897
rect 25320 27888 25372 27940
rect 26240 27956 26292 28008
rect 24492 27820 24544 27872
rect 25504 27820 25556 27872
rect 25596 27820 25648 27872
rect 7114 27718 7166 27770
rect 7178 27718 7230 27770
rect 7242 27718 7294 27770
rect 7306 27718 7358 27770
rect 7370 27718 7422 27770
rect 13830 27718 13882 27770
rect 13894 27718 13946 27770
rect 13958 27718 14010 27770
rect 14022 27718 14074 27770
rect 14086 27718 14138 27770
rect 20546 27718 20598 27770
rect 20610 27718 20662 27770
rect 20674 27718 20726 27770
rect 20738 27718 20790 27770
rect 20802 27718 20854 27770
rect 27262 27718 27314 27770
rect 27326 27718 27378 27770
rect 27390 27718 27442 27770
rect 27454 27718 27506 27770
rect 27518 27718 27570 27770
rect 2872 27616 2924 27668
rect 2504 27591 2556 27600
rect 2504 27557 2538 27591
rect 2538 27557 2556 27591
rect 2504 27548 2556 27557
rect 4436 27616 4488 27668
rect 2228 27455 2280 27464
rect 2228 27421 2237 27455
rect 2237 27421 2271 27455
rect 2271 27421 2280 27455
rect 2228 27412 2280 27421
rect 4252 27548 4304 27600
rect 8944 27616 8996 27668
rect 9404 27616 9456 27668
rect 9772 27616 9824 27668
rect 4620 27523 4672 27532
rect 4620 27489 4629 27523
rect 4629 27489 4663 27523
rect 4663 27489 4672 27523
rect 4620 27480 4672 27489
rect 5264 27523 5316 27532
rect 5264 27489 5273 27523
rect 5273 27489 5307 27523
rect 5307 27489 5316 27523
rect 5264 27480 5316 27489
rect 6828 27480 6880 27532
rect 7840 27480 7892 27532
rect 8024 27523 8076 27532
rect 8024 27489 8033 27523
rect 8033 27489 8067 27523
rect 8067 27489 8076 27523
rect 8024 27480 8076 27489
rect 8392 27480 8444 27532
rect 8760 27480 8812 27532
rect 9588 27480 9640 27532
rect 9956 27523 10008 27532
rect 9956 27489 9965 27523
rect 9965 27489 9999 27523
rect 9999 27489 10008 27523
rect 9956 27480 10008 27489
rect 3608 27387 3660 27396
rect 3608 27353 3617 27387
rect 3617 27353 3651 27387
rect 3651 27353 3660 27387
rect 3608 27344 3660 27353
rect 4620 27276 4672 27328
rect 8024 27344 8076 27396
rect 8576 27344 8628 27396
rect 8852 27412 8904 27464
rect 10140 27480 10192 27532
rect 10968 27616 11020 27668
rect 14832 27616 14884 27668
rect 16396 27616 16448 27668
rect 16672 27616 16724 27668
rect 17224 27616 17276 27668
rect 17776 27616 17828 27668
rect 10876 27548 10928 27600
rect 10968 27523 11020 27532
rect 10968 27489 10977 27523
rect 10977 27489 11011 27523
rect 11011 27489 11020 27523
rect 10968 27480 11020 27489
rect 11060 27480 11112 27532
rect 15568 27591 15620 27600
rect 15568 27557 15577 27591
rect 15577 27557 15611 27591
rect 15611 27557 15620 27591
rect 15568 27548 15620 27557
rect 12808 27523 12860 27532
rect 12808 27489 12817 27523
rect 12817 27489 12851 27523
rect 12851 27489 12860 27523
rect 12808 27480 12860 27489
rect 12900 27480 12952 27532
rect 14556 27480 14608 27532
rect 15108 27480 15160 27532
rect 18512 27548 18564 27600
rect 16948 27480 17000 27532
rect 19340 27523 19392 27532
rect 19340 27489 19358 27523
rect 19358 27489 19392 27523
rect 19340 27480 19392 27489
rect 19524 27480 19576 27532
rect 21548 27616 21600 27668
rect 20076 27591 20128 27600
rect 20076 27557 20085 27591
rect 20085 27557 20119 27591
rect 20119 27557 20128 27591
rect 20076 27548 20128 27557
rect 21824 27548 21876 27600
rect 19800 27480 19852 27532
rect 19984 27523 20036 27532
rect 19984 27489 19993 27523
rect 19993 27489 20027 27523
rect 20027 27489 20036 27523
rect 19984 27480 20036 27489
rect 21732 27480 21784 27532
rect 23112 27616 23164 27668
rect 22744 27591 22796 27600
rect 22744 27557 22753 27591
rect 22753 27557 22787 27591
rect 22787 27557 22796 27591
rect 22744 27548 22796 27557
rect 22836 27548 22888 27600
rect 22284 27480 22336 27532
rect 22928 27480 22980 27532
rect 9312 27344 9364 27396
rect 10048 27344 10100 27396
rect 12532 27344 12584 27396
rect 14188 27387 14240 27396
rect 14188 27353 14197 27387
rect 14197 27353 14231 27387
rect 14231 27353 14240 27387
rect 14188 27344 14240 27353
rect 15016 27344 15068 27396
rect 15200 27387 15252 27396
rect 15200 27353 15209 27387
rect 15209 27353 15243 27387
rect 15243 27353 15252 27387
rect 15200 27344 15252 27353
rect 7288 27276 7340 27328
rect 7932 27319 7984 27328
rect 7932 27285 7941 27319
rect 7941 27285 7975 27319
rect 7975 27285 7984 27319
rect 7932 27276 7984 27285
rect 15936 27344 15988 27396
rect 18420 27344 18472 27396
rect 15384 27276 15436 27328
rect 15844 27276 15896 27328
rect 16488 27276 16540 27328
rect 16580 27276 16632 27328
rect 16948 27319 17000 27328
rect 16948 27285 16957 27319
rect 16957 27285 16991 27319
rect 16991 27285 17000 27319
rect 16948 27276 17000 27285
rect 17776 27276 17828 27328
rect 18052 27276 18104 27328
rect 19800 27276 19852 27328
rect 20904 27276 20956 27328
rect 22284 27344 22336 27396
rect 24584 27616 24636 27668
rect 25504 27616 25556 27668
rect 24676 27548 24728 27600
rect 25596 27591 25648 27600
rect 25596 27557 25605 27591
rect 25605 27557 25639 27591
rect 25639 27557 25648 27591
rect 25596 27548 25648 27557
rect 24584 27523 24636 27532
rect 24584 27489 24593 27523
rect 24593 27489 24627 27523
rect 24627 27489 24636 27523
rect 24584 27480 24636 27489
rect 24860 27523 24912 27532
rect 24860 27489 24869 27523
rect 24869 27489 24903 27523
rect 24903 27489 24912 27523
rect 24860 27480 24912 27489
rect 25688 27523 25740 27532
rect 25688 27489 25697 27523
rect 25697 27489 25731 27523
rect 25731 27489 25740 27523
rect 25688 27480 25740 27489
rect 25780 27480 25832 27532
rect 22192 27276 22244 27328
rect 22652 27276 22704 27328
rect 25136 27319 25188 27328
rect 25136 27285 25145 27319
rect 25145 27285 25179 27319
rect 25179 27285 25188 27319
rect 25136 27276 25188 27285
rect 25228 27319 25280 27328
rect 25228 27285 25237 27319
rect 25237 27285 25271 27319
rect 25271 27285 25280 27319
rect 25228 27276 25280 27285
rect 3756 27174 3808 27226
rect 3820 27174 3872 27226
rect 3884 27174 3936 27226
rect 3948 27174 4000 27226
rect 4012 27174 4064 27226
rect 10472 27174 10524 27226
rect 10536 27174 10588 27226
rect 10600 27174 10652 27226
rect 10664 27174 10716 27226
rect 10728 27174 10780 27226
rect 17188 27174 17240 27226
rect 17252 27174 17304 27226
rect 17316 27174 17368 27226
rect 17380 27174 17432 27226
rect 17444 27174 17496 27226
rect 23904 27174 23956 27226
rect 23968 27174 24020 27226
rect 24032 27174 24084 27226
rect 24096 27174 24148 27226
rect 24160 27174 24212 27226
rect 4252 27072 4304 27124
rect 5264 27115 5316 27124
rect 5264 27081 5273 27115
rect 5273 27081 5307 27115
rect 5307 27081 5316 27115
rect 5264 27072 5316 27081
rect 5356 27115 5408 27124
rect 5356 27081 5365 27115
rect 5365 27081 5399 27115
rect 5399 27081 5408 27115
rect 5356 27072 5408 27081
rect 6092 27072 6144 27124
rect 6736 27115 6788 27124
rect 6736 27081 6745 27115
rect 6745 27081 6779 27115
rect 6779 27081 6788 27115
rect 6736 27072 6788 27081
rect 5264 26936 5316 26988
rect 2504 26868 2556 26920
rect 5080 26868 5132 26920
rect 2320 26800 2372 26852
rect 7472 27047 7524 27056
rect 7472 27013 7481 27047
rect 7481 27013 7515 27047
rect 7515 27013 7524 27047
rect 7472 27004 7524 27013
rect 8852 27072 8904 27124
rect 9036 27072 9088 27124
rect 10048 27072 10100 27124
rect 11060 27072 11112 27124
rect 12808 27072 12860 27124
rect 15200 27072 15252 27124
rect 16948 27072 17000 27124
rect 18052 27072 18104 27124
rect 18328 27115 18380 27124
rect 18328 27081 18337 27115
rect 18337 27081 18371 27115
rect 18371 27081 18380 27115
rect 18328 27072 18380 27081
rect 18420 27072 18472 27124
rect 19340 27072 19392 27124
rect 7288 26936 7340 26988
rect 7748 26979 7800 26988
rect 7748 26945 7757 26979
rect 7757 26945 7791 26979
rect 7791 26945 7800 26979
rect 7748 26936 7800 26945
rect 7840 26936 7892 26988
rect 14188 26979 14240 26988
rect 14188 26945 14197 26979
rect 14197 26945 14231 26979
rect 14231 26945 14240 26979
rect 14188 26936 14240 26945
rect 5816 26843 5868 26852
rect 5816 26809 5825 26843
rect 5825 26809 5859 26843
rect 5859 26809 5868 26843
rect 5816 26800 5868 26809
rect 2596 26775 2648 26784
rect 2596 26741 2605 26775
rect 2605 26741 2639 26775
rect 2639 26741 2648 26775
rect 2596 26732 2648 26741
rect 2688 26732 2740 26784
rect 6920 26732 6972 26784
rect 7012 26732 7064 26784
rect 8576 26911 8628 26920
rect 8576 26877 8585 26911
rect 8585 26877 8619 26911
rect 8619 26877 8628 26911
rect 8576 26868 8628 26877
rect 9680 26868 9732 26920
rect 11428 26868 11480 26920
rect 11520 26911 11572 26920
rect 11520 26877 11529 26911
rect 11529 26877 11563 26911
rect 11563 26877 11572 26911
rect 11520 26868 11572 26877
rect 11612 26911 11664 26920
rect 11612 26877 11621 26911
rect 11621 26877 11655 26911
rect 11655 26877 11664 26911
rect 11612 26868 11664 26877
rect 12808 26868 12860 26920
rect 13636 26868 13688 26920
rect 15292 27004 15344 27056
rect 15660 26868 15712 26920
rect 17868 27004 17920 27056
rect 20904 27115 20956 27124
rect 20904 27081 20913 27115
rect 20913 27081 20947 27115
rect 20947 27081 20956 27115
rect 20904 27072 20956 27081
rect 21456 27072 21508 27124
rect 21916 27115 21968 27124
rect 21916 27081 21925 27115
rect 21925 27081 21959 27115
rect 21959 27081 21968 27115
rect 21916 27072 21968 27081
rect 22468 27072 22520 27124
rect 21272 27004 21324 27056
rect 22744 27115 22796 27124
rect 22744 27081 22753 27115
rect 22753 27081 22787 27115
rect 22787 27081 22796 27115
rect 22744 27072 22796 27081
rect 22836 27072 22888 27124
rect 23388 27115 23440 27124
rect 23388 27081 23397 27115
rect 23397 27081 23431 27115
rect 23431 27081 23440 27115
rect 23388 27072 23440 27081
rect 17500 26911 17552 26920
rect 9864 26800 9916 26852
rect 11060 26800 11112 26852
rect 11336 26843 11388 26852
rect 11336 26809 11345 26843
rect 11345 26809 11379 26843
rect 11379 26809 11388 26843
rect 11336 26800 11388 26809
rect 15568 26800 15620 26852
rect 17500 26877 17509 26911
rect 17509 26877 17543 26911
rect 17543 26877 17552 26911
rect 17500 26868 17552 26877
rect 7656 26732 7708 26784
rect 13544 26775 13596 26784
rect 13544 26741 13553 26775
rect 13553 26741 13587 26775
rect 13587 26741 13596 26775
rect 13544 26732 13596 26741
rect 15384 26732 15436 26784
rect 15660 26775 15712 26784
rect 15660 26741 15669 26775
rect 15669 26741 15703 26775
rect 15703 26741 15712 26775
rect 15660 26732 15712 26741
rect 15752 26775 15804 26784
rect 15752 26741 15761 26775
rect 15761 26741 15795 26775
rect 15795 26741 15804 26775
rect 15752 26732 15804 26741
rect 17408 26800 17460 26852
rect 18512 26868 18564 26920
rect 19524 26979 19576 26988
rect 19524 26945 19533 26979
rect 19533 26945 19567 26979
rect 19567 26945 19576 26979
rect 19524 26936 19576 26945
rect 19800 26911 19852 26920
rect 19800 26877 19834 26911
rect 19834 26877 19852 26911
rect 19800 26868 19852 26877
rect 21548 26936 21600 26988
rect 22192 26936 22244 26988
rect 21272 26868 21324 26920
rect 22376 26911 22428 26920
rect 17960 26775 18012 26784
rect 17960 26741 17985 26775
rect 17985 26741 18012 26775
rect 21548 26800 21600 26852
rect 21824 26800 21876 26852
rect 22376 26877 22385 26911
rect 22385 26877 22419 26911
rect 22419 26877 22428 26911
rect 22376 26868 22428 26877
rect 22928 26868 22980 26920
rect 23480 26868 23532 26920
rect 24676 26868 24728 26920
rect 17960 26732 18012 26741
rect 18696 26775 18748 26784
rect 18696 26741 18705 26775
rect 18705 26741 18739 26775
rect 18739 26741 18748 26775
rect 18696 26732 18748 26741
rect 22100 26775 22152 26784
rect 22100 26741 22127 26775
rect 22127 26741 22152 26775
rect 22100 26732 22152 26741
rect 25320 26843 25372 26852
rect 25320 26809 25329 26843
rect 25329 26809 25363 26843
rect 25363 26809 25372 26843
rect 25320 26800 25372 26809
rect 23020 26732 23072 26784
rect 23388 26732 23440 26784
rect 23480 26732 23532 26784
rect 26240 26732 26292 26784
rect 7114 26630 7166 26682
rect 7178 26630 7230 26682
rect 7242 26630 7294 26682
rect 7306 26630 7358 26682
rect 7370 26630 7422 26682
rect 13830 26630 13882 26682
rect 13894 26630 13946 26682
rect 13958 26630 14010 26682
rect 14022 26630 14074 26682
rect 14086 26630 14138 26682
rect 20546 26630 20598 26682
rect 20610 26630 20662 26682
rect 20674 26630 20726 26682
rect 20738 26630 20790 26682
rect 20802 26630 20854 26682
rect 27262 26630 27314 26682
rect 27326 26630 27378 26682
rect 27390 26630 27442 26682
rect 27454 26630 27506 26682
rect 27518 26630 27570 26682
rect 2228 26528 2280 26580
rect 5816 26528 5868 26580
rect 7012 26528 7064 26580
rect 7472 26528 7524 26580
rect 1216 26435 1268 26444
rect 1216 26401 1250 26435
rect 1250 26401 1268 26435
rect 1216 26392 1268 26401
rect 2688 26392 2740 26444
rect 2320 26299 2372 26308
rect 2320 26265 2329 26299
rect 2329 26265 2363 26299
rect 2363 26265 2372 26299
rect 2320 26256 2372 26265
rect 2412 26231 2464 26240
rect 2412 26197 2421 26231
rect 2421 26197 2455 26231
rect 2455 26197 2464 26231
rect 2412 26188 2464 26197
rect 2596 26231 2648 26240
rect 2596 26197 2605 26231
rect 2605 26197 2639 26231
rect 2639 26197 2648 26231
rect 2596 26188 2648 26197
rect 3332 26392 3384 26444
rect 3516 26392 3568 26444
rect 4988 26435 5040 26444
rect 4988 26401 4997 26435
rect 4997 26401 5031 26435
rect 5031 26401 5040 26435
rect 4988 26392 5040 26401
rect 7104 26392 7156 26444
rect 9588 26528 9640 26580
rect 9680 26528 9732 26580
rect 12072 26528 12124 26580
rect 12900 26528 12952 26580
rect 13544 26528 13596 26580
rect 15752 26528 15804 26580
rect 15844 26528 15896 26580
rect 7564 26435 7616 26444
rect 7564 26401 7573 26435
rect 7573 26401 7607 26435
rect 7607 26401 7616 26435
rect 7564 26392 7616 26401
rect 6184 26324 6236 26376
rect 2964 26299 3016 26308
rect 2964 26265 2973 26299
rect 2973 26265 3007 26299
rect 3007 26265 3016 26299
rect 2964 26256 3016 26265
rect 5080 26256 5132 26308
rect 3148 26188 3200 26240
rect 3424 26231 3476 26240
rect 3424 26197 3433 26231
rect 3433 26197 3467 26231
rect 3467 26197 3476 26231
rect 3424 26188 3476 26197
rect 3608 26231 3660 26240
rect 3608 26197 3617 26231
rect 3617 26197 3651 26231
rect 3651 26197 3660 26231
rect 3608 26188 3660 26197
rect 5448 26231 5500 26240
rect 5448 26197 5457 26231
rect 5457 26197 5491 26231
rect 5491 26197 5500 26231
rect 5448 26188 5500 26197
rect 5632 26188 5684 26240
rect 7012 26367 7064 26376
rect 7012 26333 7021 26367
rect 7021 26333 7055 26367
rect 7055 26333 7064 26367
rect 7012 26324 7064 26333
rect 8392 26435 8444 26444
rect 8392 26401 8401 26435
rect 8401 26401 8435 26435
rect 8435 26401 8444 26435
rect 8392 26392 8444 26401
rect 11152 26460 11204 26512
rect 11336 26460 11388 26512
rect 12256 26460 12308 26512
rect 13084 26460 13136 26512
rect 8484 26324 8536 26376
rect 9036 26435 9088 26444
rect 9036 26401 9045 26435
rect 9045 26401 9079 26435
rect 9079 26401 9088 26435
rect 9036 26392 9088 26401
rect 10140 26392 10192 26444
rect 11428 26435 11480 26444
rect 11428 26401 11437 26435
rect 11437 26401 11471 26435
rect 11471 26401 11480 26435
rect 11428 26392 11480 26401
rect 11704 26392 11756 26444
rect 12072 26392 12124 26444
rect 12624 26392 12676 26444
rect 12900 26435 12952 26444
rect 12900 26401 12909 26435
rect 12909 26401 12943 26435
rect 12943 26401 12952 26435
rect 12900 26392 12952 26401
rect 13452 26392 13504 26444
rect 14280 26392 14332 26444
rect 15660 26460 15712 26512
rect 15568 26435 15620 26444
rect 15568 26401 15577 26435
rect 15577 26401 15611 26435
rect 15611 26401 15620 26435
rect 15568 26392 15620 26401
rect 17500 26528 17552 26580
rect 18696 26528 18748 26580
rect 19524 26528 19576 26580
rect 21272 26528 21324 26580
rect 16764 26392 16816 26444
rect 9864 26367 9916 26376
rect 9864 26333 9873 26367
rect 9873 26333 9907 26367
rect 9907 26333 9916 26367
rect 9864 26324 9916 26333
rect 12532 26367 12584 26376
rect 12532 26333 12541 26367
rect 12541 26333 12575 26367
rect 12575 26333 12584 26367
rect 12532 26324 12584 26333
rect 15936 26324 15988 26376
rect 6920 26188 6972 26240
rect 7748 26299 7800 26308
rect 7748 26265 7757 26299
rect 7757 26265 7791 26299
rect 7791 26265 7800 26299
rect 7748 26256 7800 26265
rect 8392 26256 8444 26308
rect 9036 26256 9088 26308
rect 14188 26256 14240 26308
rect 15292 26299 15344 26308
rect 15292 26265 15301 26299
rect 15301 26265 15335 26299
rect 15335 26265 15344 26299
rect 15292 26256 15344 26265
rect 16580 26299 16632 26308
rect 16580 26265 16589 26299
rect 16589 26265 16623 26299
rect 16623 26265 16632 26299
rect 16580 26256 16632 26265
rect 16672 26256 16724 26308
rect 17408 26324 17460 26376
rect 19524 26435 19576 26444
rect 19524 26401 19542 26435
rect 19542 26401 19576 26435
rect 19524 26392 19576 26401
rect 19800 26435 19852 26444
rect 19800 26401 19809 26435
rect 19809 26401 19843 26435
rect 19843 26401 19852 26435
rect 19800 26392 19852 26401
rect 17592 26256 17644 26308
rect 8024 26231 8076 26240
rect 8024 26197 8033 26231
rect 8033 26197 8067 26231
rect 8067 26197 8076 26231
rect 8024 26188 8076 26197
rect 8760 26188 8812 26240
rect 11244 26231 11296 26240
rect 11244 26197 11253 26231
rect 11253 26197 11287 26231
rect 11287 26197 11296 26231
rect 11244 26188 11296 26197
rect 13728 26188 13780 26240
rect 13820 26231 13872 26240
rect 13820 26197 13829 26231
rect 13829 26197 13863 26231
rect 13863 26197 13872 26231
rect 13820 26188 13872 26197
rect 14556 26188 14608 26240
rect 16856 26188 16908 26240
rect 17960 26231 18012 26240
rect 17960 26197 17969 26231
rect 17969 26197 18003 26231
rect 18003 26197 18012 26231
rect 17960 26188 18012 26197
rect 18144 26231 18196 26240
rect 18144 26197 18153 26231
rect 18153 26197 18187 26231
rect 18187 26197 18196 26231
rect 18144 26188 18196 26197
rect 18420 26231 18472 26240
rect 18420 26197 18429 26231
rect 18429 26197 18463 26231
rect 18463 26197 18472 26231
rect 18420 26188 18472 26197
rect 20720 26231 20772 26240
rect 20720 26197 20729 26231
rect 20729 26197 20763 26231
rect 20763 26197 20772 26231
rect 20720 26188 20772 26197
rect 21732 26528 21784 26580
rect 22468 26528 22520 26580
rect 24308 26571 24360 26580
rect 24308 26537 24317 26571
rect 24317 26537 24351 26571
rect 24351 26537 24360 26571
rect 24308 26528 24360 26537
rect 21548 26460 21600 26512
rect 21916 26503 21968 26512
rect 21916 26469 21925 26503
rect 21925 26469 21959 26503
rect 21959 26469 21968 26503
rect 21916 26460 21968 26469
rect 21456 26324 21508 26376
rect 22008 26435 22060 26444
rect 22008 26401 22017 26435
rect 22017 26401 22051 26435
rect 22051 26401 22060 26435
rect 22008 26392 22060 26401
rect 24400 26460 24452 26512
rect 24952 26460 25004 26512
rect 22836 26392 22888 26444
rect 23480 26435 23532 26444
rect 23480 26401 23489 26435
rect 23489 26401 23523 26435
rect 23523 26401 23532 26435
rect 23480 26392 23532 26401
rect 22652 26324 22704 26376
rect 24308 26392 24360 26444
rect 25136 26392 25188 26444
rect 25228 26392 25280 26444
rect 25964 26503 26016 26512
rect 25964 26469 25973 26503
rect 25973 26469 26007 26503
rect 26007 26469 26016 26503
rect 25964 26460 26016 26469
rect 23112 26299 23164 26308
rect 23112 26265 23121 26299
rect 23121 26265 23155 26299
rect 23155 26265 23164 26299
rect 23112 26256 23164 26265
rect 23572 26256 23624 26308
rect 24860 26324 24912 26376
rect 26148 26324 26200 26376
rect 21916 26188 21968 26240
rect 22284 26188 22336 26240
rect 24584 26188 24636 26240
rect 25412 26188 25464 26240
rect 25504 26188 25556 26240
rect 26056 26231 26108 26240
rect 26056 26197 26065 26231
rect 26065 26197 26099 26231
rect 26099 26197 26108 26231
rect 26056 26188 26108 26197
rect 3756 26086 3808 26138
rect 3820 26086 3872 26138
rect 3884 26086 3936 26138
rect 3948 26086 4000 26138
rect 4012 26086 4064 26138
rect 10472 26086 10524 26138
rect 10536 26086 10588 26138
rect 10600 26086 10652 26138
rect 10664 26086 10716 26138
rect 10728 26086 10780 26138
rect 17188 26086 17240 26138
rect 17252 26086 17304 26138
rect 17316 26086 17368 26138
rect 17380 26086 17432 26138
rect 17444 26086 17496 26138
rect 23904 26086 23956 26138
rect 23968 26086 24020 26138
rect 24032 26086 24084 26138
rect 24096 26086 24148 26138
rect 24160 26086 24212 26138
rect 1216 25984 1268 26036
rect 2412 25984 2464 26036
rect 2320 25823 2372 25832
rect 2320 25789 2329 25823
rect 2329 25789 2363 25823
rect 2363 25789 2372 25823
rect 2320 25780 2372 25789
rect 2412 25823 2464 25832
rect 2412 25789 2421 25823
rect 2421 25789 2455 25823
rect 2455 25789 2464 25823
rect 2412 25780 2464 25789
rect 4528 25984 4580 26036
rect 7104 25984 7156 26036
rect 2964 25916 3016 25968
rect 7012 25916 7064 25968
rect 3148 25780 3200 25832
rect 7656 25848 7708 25900
rect 9864 25984 9916 26036
rect 12532 25984 12584 26036
rect 15568 25984 15620 26036
rect 17960 25984 18012 26036
rect 13176 25916 13228 25968
rect 13728 25916 13780 25968
rect 18512 25984 18564 26036
rect 19524 25984 19576 26036
rect 21548 25984 21600 26036
rect 22284 25984 22336 26036
rect 22468 26027 22520 26036
rect 22468 25993 22477 26027
rect 22477 25993 22511 26027
rect 22511 25993 22520 26027
rect 22468 25984 22520 25993
rect 22836 26027 22888 26036
rect 22836 25993 22845 26027
rect 22845 25993 22879 26027
rect 22879 25993 22888 26027
rect 22836 25984 22888 25993
rect 22928 25984 22980 26036
rect 23572 25984 23624 26036
rect 24308 25984 24360 26036
rect 24952 25984 25004 26036
rect 25412 26027 25464 26036
rect 3332 25712 3384 25764
rect 3608 25712 3660 25764
rect 5264 25755 5316 25764
rect 5264 25721 5298 25755
rect 5298 25721 5316 25755
rect 5264 25712 5316 25721
rect 2504 25644 2556 25696
rect 2872 25687 2924 25696
rect 2872 25653 2897 25687
rect 2897 25653 2924 25687
rect 2872 25644 2924 25653
rect 3056 25687 3108 25696
rect 3056 25653 3065 25687
rect 3065 25653 3099 25687
rect 3099 25653 3108 25687
rect 3056 25644 3108 25653
rect 5632 25644 5684 25696
rect 5724 25644 5776 25696
rect 6184 25644 6236 25696
rect 10968 25780 11020 25832
rect 6460 25687 6512 25696
rect 6460 25653 6469 25687
rect 6469 25653 6503 25687
rect 6503 25653 6512 25687
rect 6460 25644 6512 25653
rect 8760 25712 8812 25764
rect 11244 25712 11296 25764
rect 11888 25755 11940 25764
rect 11888 25721 11922 25755
rect 11922 25721 11940 25755
rect 11888 25712 11940 25721
rect 13636 25780 13688 25832
rect 13728 25780 13780 25832
rect 14188 25780 14240 25832
rect 14372 25823 14424 25832
rect 14372 25789 14381 25823
rect 14381 25789 14415 25823
rect 14415 25789 14424 25823
rect 14372 25780 14424 25789
rect 17040 25848 17092 25900
rect 10140 25644 10192 25696
rect 13544 25687 13596 25696
rect 13544 25653 13553 25687
rect 13553 25653 13587 25687
rect 13587 25653 13596 25687
rect 13544 25644 13596 25653
rect 13820 25644 13872 25696
rect 17868 25823 17920 25832
rect 17868 25789 17877 25823
rect 17877 25789 17911 25823
rect 17911 25789 17920 25823
rect 17868 25780 17920 25789
rect 18420 25848 18472 25900
rect 18144 25780 18196 25832
rect 19800 25848 19852 25900
rect 24492 25916 24544 25968
rect 24768 25916 24820 25968
rect 25412 25993 25421 26027
rect 25421 25993 25455 26027
rect 25455 25993 25464 26027
rect 25412 25984 25464 25993
rect 25964 25984 26016 26036
rect 15844 25712 15896 25764
rect 16304 25755 16356 25764
rect 16304 25721 16322 25755
rect 16322 25721 16356 25755
rect 16304 25712 16356 25721
rect 21824 25780 21876 25832
rect 20720 25712 20772 25764
rect 22008 25780 22060 25832
rect 22284 25780 22336 25832
rect 23020 25823 23072 25832
rect 23020 25789 23029 25823
rect 23029 25789 23063 25823
rect 23063 25789 23072 25823
rect 23020 25780 23072 25789
rect 23480 25848 23532 25900
rect 24584 25780 24636 25832
rect 25228 25780 25280 25832
rect 25412 25780 25464 25832
rect 26240 25780 26292 25832
rect 26792 25755 26844 25764
rect 26792 25721 26810 25755
rect 26810 25721 26844 25755
rect 26792 25712 26844 25721
rect 15200 25687 15252 25696
rect 15200 25653 15209 25687
rect 15209 25653 15243 25687
rect 15243 25653 15252 25687
rect 15200 25644 15252 25653
rect 21640 25687 21692 25696
rect 21640 25653 21649 25687
rect 21649 25653 21683 25687
rect 21683 25653 21692 25687
rect 21640 25644 21692 25653
rect 24308 25687 24360 25696
rect 24308 25653 24317 25687
rect 24317 25653 24351 25687
rect 24351 25653 24360 25687
rect 24308 25644 24360 25653
rect 24492 25644 24544 25696
rect 25504 25644 25556 25696
rect 25596 25687 25648 25696
rect 25596 25653 25605 25687
rect 25605 25653 25639 25687
rect 25639 25653 25648 25687
rect 25596 25644 25648 25653
rect 7114 25542 7166 25594
rect 7178 25542 7230 25594
rect 7242 25542 7294 25594
rect 7306 25542 7358 25594
rect 7370 25542 7422 25594
rect 13830 25542 13882 25594
rect 13894 25542 13946 25594
rect 13958 25542 14010 25594
rect 14022 25542 14074 25594
rect 14086 25542 14138 25594
rect 20546 25542 20598 25594
rect 20610 25542 20662 25594
rect 20674 25542 20726 25594
rect 20738 25542 20790 25594
rect 20802 25542 20854 25594
rect 27262 25542 27314 25594
rect 27326 25542 27378 25594
rect 27390 25542 27442 25594
rect 27454 25542 27506 25594
rect 27518 25542 27570 25594
rect 3056 25440 3108 25492
rect 3424 25440 3476 25492
rect 3516 25440 3568 25492
rect 5264 25440 5316 25492
rect 5448 25440 5500 25492
rect 6460 25440 6512 25492
rect 9864 25440 9916 25492
rect 11888 25440 11940 25492
rect 1216 25347 1268 25356
rect 1216 25313 1225 25347
rect 1225 25313 1259 25347
rect 1259 25313 1268 25347
rect 1216 25304 1268 25313
rect 2228 25347 2280 25356
rect 2228 25313 2237 25347
rect 2237 25313 2271 25347
rect 2271 25313 2280 25347
rect 2228 25304 2280 25313
rect 2412 25347 2464 25356
rect 2412 25313 2421 25347
rect 2421 25313 2455 25347
rect 2455 25313 2464 25347
rect 2412 25304 2464 25313
rect 4436 25304 4488 25356
rect 8024 25372 8076 25424
rect 9956 25372 10008 25424
rect 6828 25236 6880 25288
rect 9036 25236 9088 25288
rect 12256 25304 12308 25356
rect 13544 25440 13596 25492
rect 13636 25483 13688 25492
rect 13636 25449 13645 25483
rect 13645 25449 13679 25483
rect 13679 25449 13688 25483
rect 13636 25440 13688 25449
rect 14188 25440 14240 25492
rect 14832 25440 14884 25492
rect 16856 25440 16908 25492
rect 17960 25440 18012 25492
rect 19708 25440 19760 25492
rect 20076 25440 20128 25492
rect 20536 25440 20588 25492
rect 13728 25415 13780 25424
rect 13728 25381 13737 25415
rect 13737 25381 13771 25415
rect 13771 25381 13780 25415
rect 13728 25372 13780 25381
rect 14924 25415 14976 25424
rect 14924 25381 14933 25415
rect 14933 25381 14967 25415
rect 14967 25381 14976 25415
rect 14924 25372 14976 25381
rect 13176 25347 13228 25356
rect 13176 25313 13185 25347
rect 13185 25313 13219 25347
rect 13219 25313 13228 25347
rect 13176 25304 13228 25313
rect 14096 25347 14148 25356
rect 14096 25313 14105 25347
rect 14105 25313 14139 25347
rect 14139 25313 14148 25347
rect 14096 25304 14148 25313
rect 15476 25372 15528 25424
rect 16396 25304 16448 25356
rect 14372 25236 14424 25288
rect 17040 25304 17092 25356
rect 17776 25304 17828 25356
rect 13820 25168 13872 25220
rect 1124 25100 1176 25152
rect 2596 25143 2648 25152
rect 2596 25109 2605 25143
rect 2605 25109 2639 25143
rect 2639 25109 2648 25143
rect 2596 25100 2648 25109
rect 4436 25100 4488 25152
rect 6920 25143 6972 25152
rect 6920 25109 6929 25143
rect 6929 25109 6963 25143
rect 6963 25109 6972 25143
rect 6920 25100 6972 25109
rect 9404 25143 9456 25152
rect 9404 25109 9413 25143
rect 9413 25109 9447 25143
rect 9447 25109 9456 25143
rect 9404 25100 9456 25109
rect 10140 25100 10192 25152
rect 11060 25100 11112 25152
rect 12072 25100 12124 25152
rect 13452 25143 13504 25152
rect 13452 25109 13461 25143
rect 13461 25109 13495 25143
rect 13495 25109 13504 25143
rect 13452 25100 13504 25109
rect 13728 25100 13780 25152
rect 14004 25100 14056 25152
rect 14648 25168 14700 25220
rect 15016 25168 15068 25220
rect 16948 25236 17000 25288
rect 18328 25415 18380 25424
rect 18328 25381 18337 25415
rect 18337 25381 18371 25415
rect 18371 25381 18380 25415
rect 18328 25372 18380 25381
rect 20352 25372 20404 25424
rect 24492 25440 24544 25492
rect 24584 25440 24636 25492
rect 25596 25440 25648 25492
rect 20076 25304 20128 25356
rect 20904 25304 20956 25356
rect 26056 25372 26108 25424
rect 26148 25372 26200 25424
rect 26240 25347 26292 25356
rect 26240 25313 26249 25347
rect 26249 25313 26283 25347
rect 26283 25313 26292 25347
rect 26240 25304 26292 25313
rect 26332 25304 26384 25356
rect 26792 25440 26844 25492
rect 22008 25236 22060 25288
rect 22560 25279 22612 25288
rect 22560 25245 22569 25279
rect 22569 25245 22603 25279
rect 22603 25245 22612 25279
rect 22560 25236 22612 25245
rect 23756 25236 23808 25288
rect 22928 25211 22980 25220
rect 22928 25177 22937 25211
rect 22937 25177 22971 25211
rect 22971 25177 22980 25211
rect 22928 25168 22980 25177
rect 24676 25168 24728 25220
rect 14832 25100 14884 25152
rect 15200 25100 15252 25152
rect 15384 25100 15436 25152
rect 15660 25100 15712 25152
rect 15752 25143 15804 25152
rect 15752 25109 15761 25143
rect 15761 25109 15795 25143
rect 15795 25109 15804 25143
rect 15752 25100 15804 25109
rect 16672 25143 16724 25152
rect 16672 25109 16681 25143
rect 16681 25109 16715 25143
rect 16715 25109 16724 25143
rect 16672 25100 16724 25109
rect 18144 25143 18196 25152
rect 18144 25109 18153 25143
rect 18153 25109 18187 25143
rect 18187 25109 18196 25143
rect 18144 25100 18196 25109
rect 20444 25143 20496 25152
rect 20444 25109 20453 25143
rect 20453 25109 20487 25143
rect 20487 25109 20496 25143
rect 20444 25100 20496 25109
rect 23020 25143 23072 25152
rect 23020 25109 23029 25143
rect 23029 25109 23063 25143
rect 23063 25109 23072 25143
rect 23020 25100 23072 25109
rect 25504 25100 25556 25152
rect 3756 24998 3808 25050
rect 3820 24998 3872 25050
rect 3884 24998 3936 25050
rect 3948 24998 4000 25050
rect 4012 24998 4064 25050
rect 10472 24998 10524 25050
rect 10536 24998 10588 25050
rect 10600 24998 10652 25050
rect 10664 24998 10716 25050
rect 10728 24998 10780 25050
rect 17188 24998 17240 25050
rect 17252 24998 17304 25050
rect 17316 24998 17368 25050
rect 17380 24998 17432 25050
rect 17444 24998 17496 25050
rect 23904 24998 23956 25050
rect 23968 24998 24020 25050
rect 24032 24998 24084 25050
rect 24096 24998 24148 25050
rect 24160 24998 24212 25050
rect 2412 24896 2464 24948
rect 2596 24896 2648 24948
rect 3056 24896 3108 24948
rect 4804 24896 4856 24948
rect 6920 24896 6972 24948
rect 9036 24896 9088 24948
rect 10968 24896 11020 24948
rect 2872 24871 2924 24880
rect 2872 24837 2881 24871
rect 2881 24837 2915 24871
rect 2915 24837 2924 24871
rect 2872 24828 2924 24837
rect 4528 24871 4580 24880
rect 4528 24837 4537 24871
rect 4537 24837 4571 24871
rect 4571 24837 4580 24871
rect 4528 24828 4580 24837
rect 1124 24667 1176 24676
rect 1124 24633 1158 24667
rect 1158 24633 1176 24667
rect 1124 24624 1176 24633
rect 1216 24624 1268 24676
rect 1860 24624 1912 24676
rect 3148 24624 3200 24676
rect 3424 24692 3476 24744
rect 5080 24760 5132 24812
rect 5724 24871 5776 24880
rect 5724 24837 5733 24871
rect 5733 24837 5767 24871
rect 5767 24837 5776 24871
rect 5724 24828 5776 24837
rect 6460 24828 6512 24880
rect 14096 24896 14148 24948
rect 14924 24939 14976 24948
rect 14924 24905 14933 24939
rect 14933 24905 14967 24939
rect 14967 24905 14976 24939
rect 14924 24896 14976 24905
rect 15016 24939 15068 24948
rect 15016 24905 15025 24939
rect 15025 24905 15059 24939
rect 15059 24905 15068 24939
rect 15016 24896 15068 24905
rect 15568 24896 15620 24948
rect 15752 24896 15804 24948
rect 16304 24896 16356 24948
rect 16396 24939 16448 24948
rect 16396 24905 16405 24939
rect 16405 24905 16439 24939
rect 16439 24905 16448 24939
rect 16396 24896 16448 24905
rect 6920 24692 6972 24744
rect 14280 24828 14332 24880
rect 14464 24828 14516 24880
rect 14832 24828 14884 24880
rect 13452 24760 13504 24812
rect 13820 24760 13872 24812
rect 7564 24735 7616 24744
rect 5632 24624 5684 24676
rect 2688 24556 2740 24608
rect 4804 24599 4856 24608
rect 4804 24565 4813 24599
rect 4813 24565 4847 24599
rect 4847 24565 4856 24599
rect 4804 24556 4856 24565
rect 4896 24599 4948 24608
rect 4896 24565 4905 24599
rect 4905 24565 4939 24599
rect 4939 24565 4948 24599
rect 4896 24556 4948 24565
rect 5448 24599 5500 24608
rect 5448 24565 5457 24599
rect 5457 24565 5491 24599
rect 5491 24565 5500 24599
rect 5448 24556 5500 24565
rect 6828 24556 6880 24608
rect 7564 24701 7573 24735
rect 7573 24701 7607 24735
rect 7607 24701 7616 24735
rect 7564 24692 7616 24701
rect 7840 24692 7892 24744
rect 10048 24735 10100 24744
rect 7656 24667 7708 24676
rect 7656 24633 7665 24667
rect 7665 24633 7699 24667
rect 7699 24633 7708 24667
rect 7656 24624 7708 24633
rect 8668 24624 8720 24676
rect 7472 24599 7524 24608
rect 7472 24565 7481 24599
rect 7481 24565 7515 24599
rect 7515 24565 7524 24599
rect 7472 24556 7524 24565
rect 8852 24556 8904 24608
rect 10048 24701 10057 24735
rect 10057 24701 10091 24735
rect 10091 24701 10100 24735
rect 10048 24692 10100 24701
rect 10140 24735 10192 24744
rect 10140 24701 10149 24735
rect 10149 24701 10183 24735
rect 10183 24701 10192 24735
rect 10140 24692 10192 24701
rect 10416 24735 10468 24744
rect 10416 24701 10425 24735
rect 10425 24701 10459 24735
rect 10459 24701 10468 24735
rect 10416 24692 10468 24701
rect 10232 24667 10284 24676
rect 10232 24633 10241 24667
rect 10241 24633 10275 24667
rect 10275 24633 10284 24667
rect 10232 24624 10284 24633
rect 10324 24624 10376 24676
rect 11060 24692 11112 24744
rect 14188 24760 14240 24812
rect 14556 24760 14608 24812
rect 12900 24624 12952 24676
rect 9864 24599 9916 24608
rect 9864 24565 9873 24599
rect 9873 24565 9907 24599
rect 9907 24565 9916 24599
rect 9864 24556 9916 24565
rect 11796 24556 11848 24608
rect 13084 24599 13136 24608
rect 13084 24565 13093 24599
rect 13093 24565 13127 24599
rect 13127 24565 13136 24599
rect 14004 24692 14056 24744
rect 15108 24760 15160 24812
rect 15200 24760 15252 24812
rect 21456 24896 21508 24948
rect 24124 24896 24176 24948
rect 24768 24896 24820 24948
rect 16580 24803 16632 24812
rect 16580 24769 16589 24803
rect 16589 24769 16623 24803
rect 16623 24769 16632 24803
rect 16580 24760 16632 24769
rect 16672 24803 16724 24812
rect 16672 24769 16681 24803
rect 16681 24769 16715 24803
rect 16715 24769 16724 24803
rect 16672 24760 16724 24769
rect 22008 24871 22060 24880
rect 22008 24837 22017 24871
rect 22017 24837 22051 24871
rect 22051 24837 22060 24871
rect 22008 24828 22060 24837
rect 24308 24828 24360 24880
rect 25872 24896 25924 24948
rect 19800 24760 19852 24812
rect 21824 24760 21876 24812
rect 22560 24760 22612 24812
rect 23296 24760 23348 24812
rect 16304 24735 16356 24744
rect 16304 24701 16313 24735
rect 16313 24701 16347 24735
rect 16347 24701 16356 24735
rect 16304 24692 16356 24701
rect 14464 24624 14516 24676
rect 17408 24735 17460 24744
rect 17408 24701 17417 24735
rect 17417 24701 17451 24735
rect 17451 24701 17460 24735
rect 17408 24692 17460 24701
rect 18144 24692 18196 24744
rect 20444 24735 20496 24744
rect 20444 24701 20478 24735
rect 20478 24701 20496 24735
rect 20444 24692 20496 24701
rect 22652 24735 22704 24744
rect 22652 24701 22661 24735
rect 22661 24701 22695 24735
rect 22695 24701 22704 24735
rect 22652 24692 22704 24701
rect 23020 24735 23072 24744
rect 23020 24701 23029 24735
rect 23029 24701 23063 24735
rect 23063 24701 23072 24735
rect 23020 24692 23072 24701
rect 23112 24735 23164 24744
rect 23112 24701 23121 24735
rect 23121 24701 23155 24735
rect 23155 24701 23164 24735
rect 23112 24692 23164 24701
rect 23480 24735 23532 24744
rect 23480 24701 23489 24735
rect 23489 24701 23523 24735
rect 23523 24701 23532 24735
rect 23480 24692 23532 24701
rect 24124 24692 24176 24744
rect 13084 24556 13136 24565
rect 14740 24556 14792 24608
rect 15200 24599 15252 24608
rect 15200 24565 15227 24599
rect 15227 24565 15252 24599
rect 15200 24556 15252 24565
rect 15660 24556 15712 24608
rect 15936 24556 15988 24608
rect 17224 24556 17276 24608
rect 17316 24556 17368 24608
rect 21640 24667 21692 24676
rect 21640 24633 21649 24667
rect 21649 24633 21683 24667
rect 21683 24633 21692 24667
rect 21640 24624 21692 24633
rect 18512 24556 18564 24608
rect 19708 24556 19760 24608
rect 20076 24599 20128 24608
rect 20076 24565 20085 24599
rect 20085 24565 20119 24599
rect 20119 24565 20128 24599
rect 20076 24556 20128 24565
rect 22836 24556 22888 24608
rect 23756 24556 23808 24608
rect 24308 24735 24360 24744
rect 24308 24701 24317 24735
rect 24317 24701 24351 24735
rect 24351 24701 24360 24735
rect 24308 24692 24360 24701
rect 25412 24828 25464 24880
rect 24768 24667 24820 24676
rect 24768 24633 24777 24667
rect 24777 24633 24811 24667
rect 24811 24633 24820 24667
rect 24768 24624 24820 24633
rect 25504 24692 25556 24744
rect 25412 24624 25464 24676
rect 26424 24556 26476 24608
rect 26976 24599 27028 24608
rect 26976 24565 26985 24599
rect 26985 24565 27019 24599
rect 27019 24565 27028 24599
rect 26976 24556 27028 24565
rect 7114 24454 7166 24506
rect 7178 24454 7230 24506
rect 7242 24454 7294 24506
rect 7306 24454 7358 24506
rect 7370 24454 7422 24506
rect 13830 24454 13882 24506
rect 13894 24454 13946 24506
rect 13958 24454 14010 24506
rect 14022 24454 14074 24506
rect 14086 24454 14138 24506
rect 20546 24454 20598 24506
rect 20610 24454 20662 24506
rect 20674 24454 20726 24506
rect 20738 24454 20790 24506
rect 20802 24454 20854 24506
rect 27262 24454 27314 24506
rect 27326 24454 27378 24506
rect 27390 24454 27442 24506
rect 27454 24454 27506 24506
rect 27518 24454 27570 24506
rect 1860 24259 1912 24268
rect 1860 24225 1869 24259
rect 1869 24225 1903 24259
rect 1903 24225 1912 24259
rect 1860 24216 1912 24225
rect 2228 24284 2280 24336
rect 2780 24284 2832 24336
rect 3056 24352 3108 24404
rect 3148 24352 3200 24404
rect 4804 24284 4856 24336
rect 1124 24012 1176 24064
rect 3516 24259 3568 24268
rect 3516 24225 3550 24259
rect 3550 24225 3568 24259
rect 3516 24216 3568 24225
rect 6092 24284 6144 24336
rect 7012 24352 7064 24404
rect 7656 24395 7708 24404
rect 7656 24361 7665 24395
rect 7665 24361 7699 24395
rect 7699 24361 7708 24395
rect 7656 24352 7708 24361
rect 8668 24395 8720 24404
rect 8668 24361 8677 24395
rect 8677 24361 8711 24395
rect 8711 24361 8720 24395
rect 8668 24352 8720 24361
rect 10324 24352 10376 24404
rect 10416 24352 10468 24404
rect 5264 24259 5316 24268
rect 5264 24225 5273 24259
rect 5273 24225 5307 24259
rect 5307 24225 5316 24259
rect 5264 24216 5316 24225
rect 6184 24259 6236 24268
rect 6184 24225 6193 24259
rect 6193 24225 6227 24259
rect 6227 24225 6236 24259
rect 6184 24216 6236 24225
rect 6460 24216 6512 24268
rect 6828 24259 6880 24268
rect 6828 24225 6837 24259
rect 6837 24225 6871 24259
rect 6871 24225 6880 24259
rect 6828 24216 6880 24225
rect 7012 24259 7064 24268
rect 7012 24225 7021 24259
rect 7021 24225 7055 24259
rect 7055 24225 7064 24259
rect 7012 24216 7064 24225
rect 3424 24012 3476 24064
rect 3608 24012 3660 24064
rect 4896 24080 4948 24132
rect 6552 24080 6604 24132
rect 6368 24012 6420 24064
rect 6460 24055 6512 24064
rect 6460 24021 6469 24055
rect 6469 24021 6503 24055
rect 6503 24021 6512 24055
rect 6460 24012 6512 24021
rect 6920 24012 6972 24064
rect 7932 24216 7984 24268
rect 7472 24148 7524 24200
rect 8116 24191 8168 24200
rect 8116 24157 8125 24191
rect 8125 24157 8159 24191
rect 8159 24157 8168 24191
rect 8852 24259 8904 24268
rect 8852 24225 8861 24259
rect 8861 24225 8895 24259
rect 8895 24225 8904 24259
rect 8852 24216 8904 24225
rect 8944 24259 8996 24268
rect 8944 24225 8953 24259
rect 8953 24225 8987 24259
rect 8987 24225 8996 24259
rect 8944 24216 8996 24225
rect 8116 24148 8168 24157
rect 8576 24148 8628 24200
rect 9404 24216 9456 24268
rect 10232 24284 10284 24336
rect 11796 24352 11848 24404
rect 10048 24216 10100 24268
rect 10968 24216 11020 24268
rect 7932 24080 7984 24132
rect 12164 24216 12216 24268
rect 13084 24352 13136 24404
rect 13728 24327 13780 24336
rect 13728 24293 13737 24327
rect 13737 24293 13771 24327
rect 13771 24293 13780 24327
rect 13728 24284 13780 24293
rect 15200 24352 15252 24404
rect 15292 24352 15344 24404
rect 15476 24395 15528 24404
rect 15476 24361 15485 24395
rect 15485 24361 15519 24395
rect 15519 24361 15528 24395
rect 15476 24352 15528 24361
rect 16304 24395 16356 24404
rect 16304 24361 16306 24395
rect 16306 24361 16340 24395
rect 16340 24361 16356 24395
rect 16304 24352 16356 24361
rect 16580 24395 16632 24404
rect 16580 24361 16589 24395
rect 16589 24361 16623 24395
rect 16623 24361 16632 24395
rect 16580 24352 16632 24361
rect 17224 24395 17276 24404
rect 17224 24361 17233 24395
rect 17233 24361 17267 24395
rect 17267 24361 17276 24395
rect 17224 24352 17276 24361
rect 17316 24352 17368 24404
rect 17408 24352 17460 24404
rect 13820 24216 13872 24268
rect 12808 24080 12860 24132
rect 14280 24148 14332 24200
rect 14740 24191 14792 24200
rect 14740 24157 14749 24191
rect 14749 24157 14783 24191
rect 14783 24157 14792 24191
rect 14740 24148 14792 24157
rect 15016 24259 15068 24268
rect 15016 24225 15025 24259
rect 15025 24225 15059 24259
rect 15059 24225 15068 24259
rect 15016 24216 15068 24225
rect 15384 24216 15436 24268
rect 15568 24259 15620 24268
rect 15568 24225 15577 24259
rect 15577 24225 15611 24259
rect 15611 24225 15620 24259
rect 15568 24216 15620 24225
rect 18512 24352 18564 24404
rect 22652 24352 22704 24404
rect 22928 24352 22980 24404
rect 19340 24327 19392 24336
rect 16764 24259 16816 24268
rect 16764 24225 16773 24259
rect 16773 24225 16807 24259
rect 16807 24225 16816 24259
rect 16764 24216 16816 24225
rect 15476 24148 15528 24200
rect 16396 24148 16448 24200
rect 14464 24080 14516 24132
rect 16948 24259 17000 24268
rect 16948 24225 16957 24259
rect 16957 24225 16991 24259
rect 16991 24225 17000 24259
rect 16948 24216 17000 24225
rect 17040 24216 17092 24268
rect 17500 24259 17552 24268
rect 17500 24225 17509 24259
rect 17509 24225 17543 24259
rect 17543 24225 17552 24259
rect 17500 24216 17552 24225
rect 19340 24293 19349 24327
rect 19349 24293 19383 24327
rect 19383 24293 19392 24327
rect 19340 24284 19392 24293
rect 18328 24216 18380 24268
rect 18420 24216 18472 24268
rect 18788 24216 18840 24268
rect 19800 24216 19852 24268
rect 19984 24259 20036 24268
rect 19984 24225 20018 24259
rect 20018 24225 20036 24259
rect 19984 24216 20036 24225
rect 21640 24216 21692 24268
rect 23480 24352 23532 24404
rect 23664 24352 23716 24404
rect 24308 24352 24360 24404
rect 24860 24352 24912 24404
rect 7380 24012 7432 24064
rect 7656 24012 7708 24064
rect 11336 24012 11388 24064
rect 13084 24055 13136 24064
rect 13084 24021 13093 24055
rect 13093 24021 13127 24055
rect 13127 24021 13136 24055
rect 13084 24012 13136 24021
rect 13176 24012 13228 24064
rect 13452 24012 13504 24064
rect 14188 24012 14240 24064
rect 18696 24191 18748 24200
rect 18696 24157 18705 24191
rect 18705 24157 18739 24191
rect 18739 24157 18748 24191
rect 18696 24148 18748 24157
rect 19708 24080 19760 24132
rect 22836 24148 22888 24200
rect 23296 24216 23348 24268
rect 15200 24012 15252 24064
rect 18420 24012 18472 24064
rect 21272 24055 21324 24064
rect 21272 24021 21281 24055
rect 21281 24021 21315 24055
rect 21315 24021 21324 24055
rect 21272 24012 21324 24021
rect 22008 24012 22060 24064
rect 24768 24284 24820 24336
rect 25412 24352 25464 24404
rect 26424 24395 26476 24404
rect 26424 24361 26433 24395
rect 26433 24361 26467 24395
rect 26467 24361 26476 24395
rect 26424 24352 26476 24361
rect 26976 24352 27028 24404
rect 24400 24148 24452 24200
rect 25044 24148 25096 24200
rect 26240 24216 26292 24268
rect 24584 24055 24636 24064
rect 24584 24021 24593 24055
rect 24593 24021 24627 24055
rect 24627 24021 24636 24055
rect 24584 24012 24636 24021
rect 25964 24012 26016 24064
rect 26056 24055 26108 24064
rect 26056 24021 26065 24055
rect 26065 24021 26099 24055
rect 26099 24021 26108 24055
rect 26056 24012 26108 24021
rect 26424 24012 26476 24064
rect 3756 23910 3808 23962
rect 3820 23910 3872 23962
rect 3884 23910 3936 23962
rect 3948 23910 4000 23962
rect 4012 23910 4064 23962
rect 10472 23910 10524 23962
rect 10536 23910 10588 23962
rect 10600 23910 10652 23962
rect 10664 23910 10716 23962
rect 10728 23910 10780 23962
rect 17188 23910 17240 23962
rect 17252 23910 17304 23962
rect 17316 23910 17368 23962
rect 17380 23910 17432 23962
rect 17444 23910 17496 23962
rect 23904 23910 23956 23962
rect 23968 23910 24020 23962
rect 24032 23910 24084 23962
rect 24096 23910 24148 23962
rect 24160 23910 24212 23962
rect 3056 23808 3108 23860
rect 3516 23851 3568 23860
rect 3516 23817 3525 23851
rect 3525 23817 3559 23851
rect 3559 23817 3568 23851
rect 3516 23808 3568 23817
rect 4712 23740 4764 23792
rect 848 23647 900 23656
rect 848 23613 857 23647
rect 857 23613 891 23647
rect 891 23613 900 23647
rect 848 23604 900 23613
rect 1124 23647 1176 23656
rect 1124 23613 1158 23647
rect 1158 23613 1176 23647
rect 1124 23604 1176 23613
rect 3332 23647 3384 23656
rect 3332 23613 3341 23647
rect 3341 23613 3375 23647
rect 3375 23613 3384 23647
rect 3332 23604 3384 23613
rect 3608 23604 3660 23656
rect 5264 23808 5316 23860
rect 6460 23808 6512 23860
rect 6552 23808 6604 23860
rect 6920 23808 6972 23860
rect 8116 23851 8168 23860
rect 8116 23817 8125 23851
rect 8125 23817 8159 23851
rect 8159 23817 8168 23851
rect 8116 23808 8168 23817
rect 9864 23808 9916 23860
rect 10232 23808 10284 23860
rect 5540 23647 5592 23656
rect 5540 23613 5554 23647
rect 5554 23613 5588 23647
rect 5588 23613 5592 23647
rect 5540 23604 5592 23613
rect 2688 23579 2740 23588
rect 2688 23545 2697 23579
rect 2697 23545 2731 23579
rect 2731 23545 2740 23579
rect 2688 23536 2740 23545
rect 5172 23579 5224 23588
rect 5172 23545 5181 23579
rect 5181 23545 5215 23579
rect 5215 23545 5224 23579
rect 5172 23536 5224 23545
rect 5356 23579 5408 23588
rect 5356 23545 5365 23579
rect 5365 23545 5399 23579
rect 5399 23545 5408 23579
rect 5356 23536 5408 23545
rect 7564 23740 7616 23792
rect 7380 23647 7432 23656
rect 7380 23613 7389 23647
rect 7389 23613 7423 23647
rect 7423 23613 7432 23647
rect 7380 23604 7432 23613
rect 7564 23604 7616 23656
rect 7840 23604 7892 23656
rect 7932 23604 7984 23656
rect 8208 23647 8260 23656
rect 8208 23613 8217 23647
rect 8217 23613 8251 23647
rect 8251 23613 8260 23647
rect 8208 23604 8260 23613
rect 8576 23604 8628 23656
rect 8852 23647 8904 23656
rect 8852 23613 8861 23647
rect 8861 23613 8895 23647
rect 8895 23613 8904 23647
rect 8852 23604 8904 23613
rect 3056 23511 3108 23520
rect 3056 23477 3065 23511
rect 3065 23477 3099 23511
rect 3099 23477 3108 23511
rect 3056 23468 3108 23477
rect 3516 23468 3568 23520
rect 4896 23511 4948 23520
rect 4896 23477 4905 23511
rect 4905 23477 4939 23511
rect 4939 23477 4948 23511
rect 4896 23468 4948 23477
rect 4988 23468 5040 23520
rect 5264 23468 5316 23520
rect 7012 23468 7064 23520
rect 9312 23536 9364 23588
rect 11336 23851 11388 23860
rect 11336 23817 11345 23851
rect 11345 23817 11379 23851
rect 11379 23817 11388 23851
rect 11336 23808 11388 23817
rect 12164 23808 12216 23860
rect 12900 23851 12952 23860
rect 12900 23817 12909 23851
rect 12909 23817 12943 23851
rect 12943 23817 12952 23851
rect 12900 23808 12952 23817
rect 13084 23808 13136 23860
rect 14464 23851 14516 23860
rect 14464 23817 14473 23851
rect 14473 23817 14507 23851
rect 14507 23817 14516 23851
rect 14464 23808 14516 23817
rect 11060 23604 11112 23656
rect 13820 23740 13872 23792
rect 13176 23672 13228 23724
rect 14740 23740 14792 23792
rect 11888 23536 11940 23588
rect 15568 23808 15620 23860
rect 15844 23808 15896 23860
rect 18420 23808 18472 23860
rect 19984 23851 20036 23860
rect 19984 23817 19993 23851
rect 19993 23817 20027 23851
rect 20027 23817 20036 23851
rect 19984 23808 20036 23817
rect 20352 23808 20404 23860
rect 21272 23808 21324 23860
rect 24768 23808 24820 23860
rect 15200 23783 15252 23792
rect 15200 23749 15209 23783
rect 15209 23749 15243 23783
rect 15243 23749 15252 23783
rect 15200 23740 15252 23749
rect 18512 23740 18564 23792
rect 15476 23604 15528 23656
rect 9036 23511 9088 23520
rect 9036 23477 9045 23511
rect 9045 23477 9079 23511
rect 9079 23477 9088 23511
rect 9036 23468 9088 23477
rect 18788 23647 18840 23656
rect 18788 23613 18797 23647
rect 18797 23613 18831 23647
rect 18831 23613 18840 23647
rect 18788 23604 18840 23613
rect 19616 23604 19668 23656
rect 20444 23604 20496 23656
rect 22652 23672 22704 23724
rect 21824 23647 21876 23656
rect 21824 23613 21833 23647
rect 21833 23613 21867 23647
rect 21867 23613 21876 23647
rect 21824 23604 21876 23613
rect 21916 23604 21968 23656
rect 24492 23604 24544 23656
rect 19432 23536 19484 23588
rect 22100 23536 22152 23588
rect 24400 23536 24452 23588
rect 24952 23647 25004 23656
rect 24952 23613 24961 23647
rect 24961 23613 24995 23647
rect 24995 23613 25004 23647
rect 24952 23604 25004 23613
rect 13544 23511 13596 23520
rect 13544 23477 13553 23511
rect 13553 23477 13587 23511
rect 13587 23477 13596 23511
rect 13544 23468 13596 23477
rect 14740 23468 14792 23520
rect 15016 23468 15068 23520
rect 18696 23468 18748 23520
rect 19524 23468 19576 23520
rect 19800 23468 19852 23520
rect 22192 23468 22244 23520
rect 23480 23468 23532 23520
rect 25504 23604 25556 23656
rect 25780 23604 25832 23656
rect 25596 23536 25648 23588
rect 26240 23468 26292 23520
rect 7114 23366 7166 23418
rect 7178 23366 7230 23418
rect 7242 23366 7294 23418
rect 7306 23366 7358 23418
rect 7370 23366 7422 23418
rect 13830 23366 13882 23418
rect 13894 23366 13946 23418
rect 13958 23366 14010 23418
rect 14022 23366 14074 23418
rect 14086 23366 14138 23418
rect 20546 23366 20598 23418
rect 20610 23366 20662 23418
rect 20674 23366 20726 23418
rect 20738 23366 20790 23418
rect 20802 23366 20854 23418
rect 27262 23366 27314 23418
rect 27326 23366 27378 23418
rect 27390 23366 27442 23418
rect 27454 23366 27506 23418
rect 27518 23366 27570 23418
rect 2688 23264 2740 23316
rect 2780 23264 2832 23316
rect 3332 23264 3384 23316
rect 3516 23307 3568 23316
rect 2872 23128 2924 23180
rect 3516 23273 3543 23307
rect 3543 23273 3568 23307
rect 3516 23264 3568 23273
rect 4896 23264 4948 23316
rect 5448 23264 5500 23316
rect 6920 23264 6972 23316
rect 3608 23196 3660 23248
rect 4068 23128 4120 23180
rect 4712 23171 4764 23180
rect 4712 23137 4721 23171
rect 4721 23137 4755 23171
rect 4755 23137 4764 23171
rect 4712 23128 4764 23137
rect 4988 23128 5040 23180
rect 5172 23128 5224 23180
rect 6092 23128 6144 23180
rect 6828 23171 6880 23180
rect 6828 23137 6837 23171
rect 6837 23137 6871 23171
rect 6871 23137 6880 23171
rect 6828 23128 6880 23137
rect 7012 23128 7064 23180
rect 2228 23103 2280 23112
rect 2228 23069 2237 23103
rect 2237 23069 2271 23103
rect 2271 23069 2280 23103
rect 2228 23060 2280 23069
rect 3424 23060 3476 23112
rect 8208 23264 8260 23316
rect 9956 23264 10008 23316
rect 10416 23264 10468 23316
rect 7748 23196 7800 23248
rect 9036 23196 9088 23248
rect 9680 23239 9732 23248
rect 9680 23205 9689 23239
rect 9689 23205 9723 23239
rect 9723 23205 9732 23239
rect 9680 23196 9732 23205
rect 9864 23171 9916 23180
rect 9864 23137 9873 23171
rect 9873 23137 9907 23171
rect 9907 23137 9916 23171
rect 9864 23128 9916 23137
rect 9956 23171 10008 23180
rect 9956 23137 9965 23171
rect 9965 23137 9999 23171
rect 9999 23137 10008 23171
rect 9956 23128 10008 23137
rect 10048 23128 10100 23180
rect 10140 23171 10192 23180
rect 10140 23137 10149 23171
rect 10149 23137 10183 23171
rect 10183 23137 10192 23171
rect 10140 23128 10192 23137
rect 10232 23128 10284 23180
rect 10416 23171 10468 23180
rect 10416 23137 10425 23171
rect 10425 23137 10459 23171
rect 10459 23137 10468 23171
rect 10416 23128 10468 23137
rect 11152 23196 11204 23248
rect 11520 23239 11572 23248
rect 11520 23205 11529 23239
rect 11529 23205 11563 23239
rect 11563 23205 11572 23239
rect 11520 23196 11572 23205
rect 14740 23307 14792 23316
rect 14740 23273 14749 23307
rect 14749 23273 14783 23307
rect 14783 23273 14792 23307
rect 14740 23264 14792 23273
rect 15476 23264 15528 23316
rect 16580 23264 16632 23316
rect 16948 23264 17000 23316
rect 19340 23307 19392 23316
rect 19340 23273 19349 23307
rect 19349 23273 19383 23307
rect 19383 23273 19392 23307
rect 19340 23264 19392 23273
rect 21824 23307 21876 23316
rect 21824 23273 21833 23307
rect 21833 23273 21867 23307
rect 21867 23273 21876 23307
rect 21824 23264 21876 23273
rect 17040 23196 17092 23248
rect 11060 23128 11112 23180
rect 11980 23128 12032 23180
rect 12072 23171 12124 23180
rect 12072 23137 12081 23171
rect 12081 23137 12115 23171
rect 12115 23137 12124 23171
rect 12072 23128 12124 23137
rect 12256 23171 12308 23180
rect 12256 23137 12265 23171
rect 12265 23137 12299 23171
rect 12299 23137 12308 23171
rect 12256 23128 12308 23137
rect 13544 23128 13596 23180
rect 14280 23171 14332 23180
rect 4528 23035 4580 23044
rect 3056 22967 3108 22976
rect 3056 22933 3065 22967
rect 3065 22933 3099 22967
rect 3099 22933 3108 22967
rect 3056 22924 3108 22933
rect 4528 23001 4537 23035
rect 4537 23001 4571 23035
rect 4571 23001 4580 23035
rect 4528 22992 4580 23001
rect 7656 22992 7708 23044
rect 12808 23060 12860 23112
rect 12072 22992 12124 23044
rect 3608 22924 3660 22976
rect 5540 22924 5592 22976
rect 6276 22967 6328 22976
rect 6276 22933 6285 22967
rect 6285 22933 6319 22967
rect 6319 22933 6328 22967
rect 6276 22924 6328 22933
rect 7472 22967 7524 22976
rect 7472 22933 7481 22967
rect 7481 22933 7515 22967
rect 7515 22933 7524 22967
rect 7472 22924 7524 22933
rect 11152 22924 11204 22976
rect 11244 22967 11296 22976
rect 11244 22933 11253 22967
rect 11253 22933 11287 22967
rect 11287 22933 11296 22967
rect 11244 22924 11296 22933
rect 11888 22967 11940 22976
rect 11888 22933 11897 22967
rect 11897 22933 11931 22967
rect 11931 22933 11940 22967
rect 11888 22924 11940 22933
rect 14280 23137 14289 23171
rect 14289 23137 14323 23171
rect 14323 23137 14332 23171
rect 14280 23128 14332 23137
rect 17868 23128 17920 23180
rect 22284 23264 22336 23316
rect 22652 23264 22704 23316
rect 24400 23264 24452 23316
rect 24492 23307 24544 23316
rect 24492 23273 24501 23307
rect 24501 23273 24535 23307
rect 24535 23273 24544 23307
rect 24492 23264 24544 23273
rect 22192 23239 22244 23248
rect 22192 23205 22204 23239
rect 22204 23205 22244 23239
rect 22192 23196 22244 23205
rect 17960 23103 18012 23112
rect 17960 23069 17969 23103
rect 17969 23069 18003 23103
rect 18003 23069 18012 23103
rect 17960 23060 18012 23069
rect 13820 22992 13872 23044
rect 22008 23128 22060 23180
rect 24584 23196 24636 23248
rect 24952 23196 25004 23248
rect 20352 23103 20404 23112
rect 20352 23069 20361 23103
rect 20361 23069 20395 23103
rect 20395 23069 20404 23103
rect 20352 23060 20404 23069
rect 21916 23103 21968 23112
rect 21916 23069 21925 23103
rect 21925 23069 21959 23103
rect 21959 23069 21968 23103
rect 21916 23060 21968 23069
rect 24400 23128 24452 23180
rect 25136 23171 25188 23180
rect 25136 23137 25145 23171
rect 25145 23137 25179 23171
rect 25179 23137 25188 23171
rect 25136 23128 25188 23137
rect 26056 23264 26108 23316
rect 26240 23264 26292 23316
rect 25872 23196 25924 23248
rect 26424 23171 26476 23180
rect 26424 23137 26433 23171
rect 26433 23137 26467 23171
rect 26467 23137 26476 23171
rect 26424 23128 26476 23137
rect 15016 22924 15068 22976
rect 18972 22924 19024 22976
rect 24492 23060 24544 23112
rect 24676 23060 24728 23112
rect 25688 23060 25740 23112
rect 23480 22924 23532 22976
rect 23572 22924 23624 22976
rect 25044 22924 25096 22976
rect 25412 22924 25464 22976
rect 26148 22967 26200 22976
rect 26148 22933 26157 22967
rect 26157 22933 26191 22967
rect 26191 22933 26200 22967
rect 26148 22924 26200 22933
rect 26976 22967 27028 22976
rect 26976 22933 26985 22967
rect 26985 22933 27019 22967
rect 27019 22933 27028 22967
rect 26976 22924 27028 22933
rect 3756 22822 3808 22874
rect 3820 22822 3872 22874
rect 3884 22822 3936 22874
rect 3948 22822 4000 22874
rect 4012 22822 4064 22874
rect 10472 22822 10524 22874
rect 10536 22822 10588 22874
rect 10600 22822 10652 22874
rect 10664 22822 10716 22874
rect 10728 22822 10780 22874
rect 17188 22822 17240 22874
rect 17252 22822 17304 22874
rect 17316 22822 17368 22874
rect 17380 22822 17432 22874
rect 17444 22822 17496 22874
rect 23904 22822 23956 22874
rect 23968 22822 24020 22874
rect 24032 22822 24084 22874
rect 24096 22822 24148 22874
rect 24160 22822 24212 22874
rect 2228 22763 2280 22772
rect 2228 22729 2237 22763
rect 2237 22729 2271 22763
rect 2271 22729 2280 22763
rect 2228 22720 2280 22729
rect 2504 22763 2556 22772
rect 2504 22729 2513 22763
rect 2513 22729 2547 22763
rect 2547 22729 2556 22763
rect 2504 22720 2556 22729
rect 2964 22720 3016 22772
rect 4528 22720 4580 22772
rect 5448 22720 5500 22772
rect 8392 22720 8444 22772
rect 11980 22720 12032 22772
rect 2688 22652 2740 22704
rect 4712 22652 4764 22704
rect 848 22627 900 22636
rect 848 22593 857 22627
rect 857 22593 891 22627
rect 891 22593 900 22627
rect 848 22584 900 22593
rect 3424 22559 3476 22568
rect 3424 22525 3433 22559
rect 3433 22525 3467 22559
rect 3467 22525 3476 22559
rect 3424 22516 3476 22525
rect 4988 22516 5040 22568
rect 5080 22559 5132 22568
rect 5080 22525 5089 22559
rect 5089 22525 5123 22559
rect 5123 22525 5132 22559
rect 5080 22516 5132 22525
rect 6276 22584 6328 22636
rect 6644 22652 6696 22704
rect 1216 22448 1268 22500
rect 2320 22423 2372 22432
rect 2320 22389 2329 22423
rect 2329 22389 2363 22423
rect 2363 22389 2372 22423
rect 2320 22380 2372 22389
rect 2780 22380 2832 22432
rect 3148 22380 3200 22432
rect 3608 22380 3660 22432
rect 4896 22423 4948 22432
rect 4896 22389 4905 22423
rect 4905 22389 4939 22423
rect 4939 22389 4948 22423
rect 4896 22380 4948 22389
rect 5540 22516 5592 22568
rect 5816 22559 5868 22568
rect 5816 22525 5825 22559
rect 5825 22525 5859 22559
rect 5859 22525 5868 22559
rect 5816 22516 5868 22525
rect 5172 22448 5224 22500
rect 6276 22491 6328 22500
rect 6276 22457 6310 22491
rect 6310 22457 6328 22491
rect 6276 22448 6328 22457
rect 7012 22559 7064 22568
rect 7012 22525 7021 22559
rect 7021 22525 7055 22559
rect 7055 22525 7064 22559
rect 7012 22516 7064 22525
rect 7104 22516 7156 22568
rect 7932 22584 7984 22636
rect 7748 22516 7800 22568
rect 12072 22652 12124 22704
rect 9864 22584 9916 22636
rect 12440 22584 12492 22636
rect 13728 22763 13780 22772
rect 13728 22729 13737 22763
rect 13737 22729 13771 22763
rect 13771 22729 13780 22763
rect 13728 22720 13780 22729
rect 17040 22720 17092 22772
rect 17868 22763 17920 22772
rect 17868 22729 17877 22763
rect 17877 22729 17911 22763
rect 17911 22729 17920 22763
rect 17868 22720 17920 22729
rect 18696 22720 18748 22772
rect 20444 22720 20496 22772
rect 14280 22652 14332 22704
rect 7840 22448 7892 22500
rect 10048 22516 10100 22568
rect 10876 22516 10928 22568
rect 11612 22516 11664 22568
rect 9956 22448 10008 22500
rect 5632 22380 5684 22432
rect 6552 22423 6604 22432
rect 6552 22389 6561 22423
rect 6561 22389 6595 22423
rect 6595 22389 6604 22423
rect 6552 22380 6604 22389
rect 7472 22380 7524 22432
rect 9680 22423 9732 22432
rect 9680 22389 9689 22423
rect 9689 22389 9723 22423
rect 9723 22389 9732 22423
rect 9680 22380 9732 22389
rect 10324 22380 10376 22432
rect 11060 22423 11112 22432
rect 11060 22389 11069 22423
rect 11069 22389 11103 22423
rect 11103 22389 11112 22423
rect 11060 22380 11112 22389
rect 12440 22448 12492 22500
rect 12900 22559 12952 22568
rect 12900 22525 12909 22559
rect 12909 22525 12943 22559
rect 12943 22525 12952 22559
rect 12900 22516 12952 22525
rect 13820 22516 13872 22568
rect 14648 22516 14700 22568
rect 15016 22516 15068 22568
rect 13452 22448 13504 22500
rect 14556 22448 14608 22500
rect 16580 22584 16632 22636
rect 19340 22652 19392 22704
rect 17408 22559 17460 22568
rect 17408 22525 17417 22559
rect 17417 22525 17451 22559
rect 17451 22525 17460 22559
rect 17408 22516 17460 22525
rect 17868 22516 17920 22568
rect 18236 22584 18288 22636
rect 18972 22584 19024 22636
rect 19064 22559 19116 22568
rect 19064 22525 19073 22559
rect 19073 22525 19107 22559
rect 19107 22525 19116 22559
rect 19064 22516 19116 22525
rect 19156 22559 19208 22568
rect 19156 22525 19165 22559
rect 19165 22525 19199 22559
rect 19199 22525 19208 22559
rect 19156 22516 19208 22525
rect 19340 22559 19392 22568
rect 19340 22525 19349 22559
rect 19349 22525 19383 22559
rect 19383 22525 19392 22559
rect 19340 22516 19392 22525
rect 19432 22516 19484 22568
rect 24952 22720 25004 22772
rect 25596 22763 25648 22772
rect 25596 22729 25605 22763
rect 25605 22729 25639 22763
rect 25639 22729 25648 22763
rect 25596 22720 25648 22729
rect 25688 22763 25740 22772
rect 25688 22729 25697 22763
rect 25697 22729 25731 22763
rect 25731 22729 25740 22763
rect 25688 22720 25740 22729
rect 23572 22652 23624 22704
rect 24400 22652 24452 22704
rect 24860 22652 24912 22704
rect 21916 22627 21968 22636
rect 21916 22593 21925 22627
rect 21925 22593 21959 22627
rect 21959 22593 21968 22627
rect 21916 22584 21968 22593
rect 25504 22584 25556 22636
rect 13176 22380 13228 22432
rect 13636 22380 13688 22432
rect 16672 22380 16724 22432
rect 17040 22380 17092 22432
rect 17684 22380 17736 22432
rect 19248 22448 19300 22500
rect 19892 22448 19944 22500
rect 21640 22559 21692 22568
rect 21640 22525 21649 22559
rect 21649 22525 21683 22559
rect 21683 22525 21692 22559
rect 21640 22516 21692 22525
rect 21364 22448 21416 22500
rect 21456 22491 21508 22500
rect 21456 22457 21465 22491
rect 21465 22457 21499 22491
rect 21499 22457 21508 22491
rect 21456 22448 21508 22457
rect 21732 22380 21784 22432
rect 23572 22448 23624 22500
rect 24584 22559 24636 22568
rect 24584 22525 24593 22559
rect 24593 22525 24627 22559
rect 24627 22525 24636 22559
rect 24584 22516 24636 22525
rect 24860 22559 24912 22568
rect 24860 22525 24869 22559
rect 24869 22525 24903 22559
rect 24903 22525 24912 22559
rect 24860 22516 24912 22525
rect 24676 22448 24728 22500
rect 25412 22559 25464 22568
rect 25412 22525 25421 22559
rect 25421 22525 25455 22559
rect 25455 22525 25464 22559
rect 25412 22516 25464 22525
rect 26516 22516 26568 22568
rect 24492 22380 24544 22432
rect 26148 22448 26200 22500
rect 26792 22491 26844 22500
rect 26792 22457 26810 22491
rect 26810 22457 26844 22491
rect 26792 22448 26844 22457
rect 7114 22278 7166 22330
rect 7178 22278 7230 22330
rect 7242 22278 7294 22330
rect 7306 22278 7358 22330
rect 7370 22278 7422 22330
rect 13830 22278 13882 22330
rect 13894 22278 13946 22330
rect 13958 22278 14010 22330
rect 14022 22278 14074 22330
rect 14086 22278 14138 22330
rect 20546 22278 20598 22330
rect 20610 22278 20662 22330
rect 20674 22278 20726 22330
rect 20738 22278 20790 22330
rect 20802 22278 20854 22330
rect 27262 22278 27314 22330
rect 27326 22278 27378 22330
rect 27390 22278 27442 22330
rect 27454 22278 27506 22330
rect 27518 22278 27570 22330
rect 1216 22219 1268 22228
rect 1216 22185 1225 22219
rect 1225 22185 1259 22219
rect 1259 22185 1268 22219
rect 1216 22176 1268 22185
rect 2320 22176 2372 22228
rect 2504 22176 2556 22228
rect 2964 22176 3016 22228
rect 3148 22176 3200 22228
rect 4068 22219 4120 22228
rect 4068 22185 4077 22219
rect 4077 22185 4111 22219
rect 4111 22185 4120 22219
rect 4068 22176 4120 22185
rect 5816 22176 5868 22228
rect 2872 22108 2924 22160
rect 5540 22040 5592 22092
rect 6000 21972 6052 22024
rect 6276 22219 6328 22228
rect 6276 22185 6285 22219
rect 6285 22185 6319 22219
rect 6319 22185 6328 22219
rect 6276 22176 6328 22185
rect 6368 22176 6420 22228
rect 6552 22176 6604 22228
rect 7472 22176 7524 22228
rect 7656 22176 7708 22228
rect 10140 22219 10192 22228
rect 10140 22185 10149 22219
rect 10149 22185 10183 22219
rect 10183 22185 10192 22219
rect 10140 22176 10192 22185
rect 12808 22219 12860 22228
rect 12808 22185 12817 22219
rect 12817 22185 12851 22219
rect 12851 22185 12860 22219
rect 12808 22176 12860 22185
rect 14648 22176 14700 22228
rect 16580 22176 16632 22228
rect 17684 22176 17736 22228
rect 6736 22040 6788 22092
rect 11244 22108 11296 22160
rect 19156 22176 19208 22228
rect 7564 22040 7616 22092
rect 7748 22083 7800 22092
rect 7748 22049 7757 22083
rect 7757 22049 7791 22083
rect 7791 22049 7800 22083
rect 7748 22040 7800 22049
rect 7932 22083 7984 22092
rect 7932 22049 7941 22083
rect 7941 22049 7975 22083
rect 7975 22049 7984 22083
rect 7932 22040 7984 22049
rect 8760 22040 8812 22092
rect 11060 22040 11112 22092
rect 11428 22083 11480 22092
rect 11428 22049 11437 22083
rect 11437 22049 11471 22083
rect 11471 22049 11480 22083
rect 11428 22040 11480 22049
rect 14188 22083 14240 22092
rect 14188 22049 14206 22083
rect 14206 22049 14240 22083
rect 14188 22040 14240 22049
rect 7012 21972 7064 22024
rect 5448 21947 5500 21956
rect 5448 21913 5457 21947
rect 5457 21913 5491 21947
rect 5491 21913 5500 21947
rect 5448 21904 5500 21913
rect 6644 21947 6696 21956
rect 6644 21913 6653 21947
rect 6653 21913 6687 21947
rect 6687 21913 6696 21947
rect 6644 21904 6696 21913
rect 6920 21904 6972 21956
rect 8024 21972 8076 22024
rect 8208 21904 8260 21956
rect 10048 21947 10100 21956
rect 10048 21913 10057 21947
rect 10057 21913 10091 21947
rect 10091 21913 10100 21947
rect 10048 21904 10100 21913
rect 4896 21836 4948 21888
rect 6092 21879 6144 21888
rect 6092 21845 6101 21879
rect 6101 21845 6135 21879
rect 6135 21845 6144 21879
rect 6092 21836 6144 21845
rect 10140 21836 10192 21888
rect 13820 21836 13872 21888
rect 16120 22015 16172 22024
rect 16120 21981 16129 22015
rect 16129 21981 16163 22015
rect 16163 21981 16172 22015
rect 16120 21972 16172 21981
rect 16304 21972 16356 22024
rect 16580 22083 16632 22092
rect 16580 22049 16589 22083
rect 16589 22049 16623 22083
rect 16623 22049 16632 22083
rect 16580 22040 16632 22049
rect 16672 22083 16724 22092
rect 16672 22049 16681 22083
rect 16681 22049 16715 22083
rect 16715 22049 16724 22083
rect 16672 22040 16724 22049
rect 16856 22083 16908 22092
rect 16856 22049 16865 22083
rect 16865 22049 16899 22083
rect 16899 22049 16908 22083
rect 16856 22040 16908 22049
rect 15752 21836 15804 21888
rect 16212 21879 16264 21888
rect 16212 21845 16221 21879
rect 16221 21845 16255 21879
rect 16255 21845 16264 21879
rect 17408 21904 17460 21956
rect 17776 22040 17828 22092
rect 19064 22040 19116 22092
rect 19616 22219 19668 22228
rect 19616 22185 19625 22219
rect 19625 22185 19659 22219
rect 19659 22185 19668 22219
rect 19616 22176 19668 22185
rect 19892 22219 19944 22228
rect 19892 22185 19901 22219
rect 19901 22185 19935 22219
rect 19935 22185 19944 22219
rect 19892 22176 19944 22185
rect 20352 22176 20404 22228
rect 24492 22176 24544 22228
rect 26792 22176 26844 22228
rect 18052 21972 18104 22024
rect 18512 21972 18564 22024
rect 18696 21972 18748 22024
rect 19248 22015 19300 22024
rect 19248 21981 19257 22015
rect 19257 21981 19291 22015
rect 19291 21981 19300 22015
rect 19248 21972 19300 21981
rect 19892 22040 19944 22092
rect 19156 21904 19208 21956
rect 19984 21904 20036 21956
rect 21364 22040 21416 22092
rect 21456 22040 21508 22092
rect 21640 22040 21692 22092
rect 21732 22040 21784 22092
rect 24400 22040 24452 22092
rect 25872 22108 25924 22160
rect 26976 22108 27028 22160
rect 20904 21904 20956 21956
rect 16212 21836 16264 21845
rect 17868 21836 17920 21888
rect 21088 21836 21140 21888
rect 22928 22015 22980 22024
rect 22928 21981 22937 22015
rect 22937 21981 22971 22015
rect 22971 21981 22980 22015
rect 22928 21972 22980 21981
rect 23572 22015 23624 22024
rect 23572 21981 23581 22015
rect 23581 21981 23615 22015
rect 23615 21981 23624 22015
rect 23572 21972 23624 21981
rect 25504 22015 25556 22024
rect 25504 21981 25513 22015
rect 25513 21981 25547 22015
rect 25547 21981 25556 22015
rect 25504 21972 25556 21981
rect 21824 21904 21876 21956
rect 24400 21904 24452 21956
rect 21548 21836 21600 21888
rect 25872 21879 25924 21888
rect 25872 21845 25881 21879
rect 25881 21845 25915 21879
rect 25915 21845 25924 21879
rect 25872 21836 25924 21845
rect 26424 21836 26476 21888
rect 3756 21734 3808 21786
rect 3820 21734 3872 21786
rect 3884 21734 3936 21786
rect 3948 21734 4000 21786
rect 4012 21734 4064 21786
rect 10472 21734 10524 21786
rect 10536 21734 10588 21786
rect 10600 21734 10652 21786
rect 10664 21734 10716 21786
rect 10728 21734 10780 21786
rect 17188 21734 17240 21786
rect 17252 21734 17304 21786
rect 17316 21734 17368 21786
rect 17380 21734 17432 21786
rect 17444 21734 17496 21786
rect 23904 21734 23956 21786
rect 23968 21734 24020 21786
rect 24032 21734 24084 21786
rect 24096 21734 24148 21786
rect 24160 21734 24212 21786
rect 3792 21632 3844 21684
rect 5264 21632 5316 21684
rect 6000 21632 6052 21684
rect 7012 21632 7064 21684
rect 7748 21632 7800 21684
rect 3516 21564 3568 21616
rect 1032 21292 1084 21344
rect 1584 21428 1636 21480
rect 2228 21428 2280 21480
rect 2412 21428 2464 21480
rect 2780 21428 2832 21480
rect 3424 21428 3476 21480
rect 3792 21471 3844 21480
rect 3792 21437 3801 21471
rect 3801 21437 3835 21471
rect 3835 21437 3844 21471
rect 3792 21428 3844 21437
rect 5172 21496 5224 21548
rect 5540 21496 5592 21548
rect 7748 21496 7800 21548
rect 8208 21632 8260 21684
rect 8760 21675 8812 21684
rect 8760 21641 8769 21675
rect 8769 21641 8803 21675
rect 8803 21641 8812 21675
rect 8760 21632 8812 21641
rect 12256 21632 12308 21684
rect 13636 21675 13688 21684
rect 13636 21641 13645 21675
rect 13645 21641 13679 21675
rect 13679 21641 13688 21675
rect 13636 21632 13688 21641
rect 14188 21675 14240 21684
rect 14188 21641 14197 21675
rect 14197 21641 14231 21675
rect 14231 21641 14240 21675
rect 14188 21632 14240 21641
rect 16672 21632 16724 21684
rect 10140 21564 10192 21616
rect 16212 21564 16264 21616
rect 16304 21564 16356 21616
rect 19340 21632 19392 21684
rect 19892 21675 19944 21684
rect 19892 21641 19901 21675
rect 19901 21641 19935 21675
rect 19935 21641 19944 21675
rect 19892 21632 19944 21641
rect 21548 21632 21600 21684
rect 23572 21632 23624 21684
rect 24676 21632 24728 21684
rect 25136 21632 25188 21684
rect 25504 21632 25556 21684
rect 25688 21632 25740 21684
rect 26516 21632 26568 21684
rect 18328 21564 18380 21616
rect 19064 21564 19116 21616
rect 4988 21471 5040 21480
rect 4988 21437 4997 21471
rect 4997 21437 5031 21471
rect 5031 21437 5040 21471
rect 4988 21428 5040 21437
rect 7012 21428 7064 21480
rect 5448 21360 5500 21412
rect 7564 21360 7616 21412
rect 8852 21428 8904 21480
rect 9588 21496 9640 21548
rect 10232 21496 10284 21548
rect 10416 21496 10468 21548
rect 12900 21496 12952 21548
rect 9680 21428 9732 21480
rect 11152 21471 11204 21480
rect 11152 21437 11170 21471
rect 11170 21437 11204 21471
rect 11152 21428 11204 21437
rect 11428 21471 11480 21480
rect 11428 21437 11437 21471
rect 11437 21437 11471 21471
rect 11471 21437 11480 21471
rect 11428 21428 11480 21437
rect 11796 21428 11848 21480
rect 9220 21360 9272 21412
rect 9864 21360 9916 21412
rect 10968 21360 11020 21412
rect 12440 21471 12492 21480
rect 12440 21437 12449 21471
rect 12449 21437 12483 21471
rect 12483 21437 12492 21471
rect 12440 21428 12492 21437
rect 13820 21471 13872 21480
rect 13820 21437 13829 21471
rect 13829 21437 13863 21471
rect 13863 21437 13872 21471
rect 13820 21428 13872 21437
rect 14648 21496 14700 21548
rect 12808 21360 12860 21412
rect 14372 21471 14424 21480
rect 14372 21437 14381 21471
rect 14381 21437 14415 21471
rect 14415 21437 14424 21471
rect 14372 21428 14424 21437
rect 14188 21360 14240 21412
rect 2688 21335 2740 21344
rect 2688 21301 2697 21335
rect 2697 21301 2731 21335
rect 2731 21301 2740 21335
rect 2688 21292 2740 21301
rect 3332 21335 3384 21344
rect 3332 21301 3341 21335
rect 3341 21301 3375 21335
rect 3375 21301 3384 21335
rect 3332 21292 3384 21301
rect 4896 21335 4948 21344
rect 4896 21301 4905 21335
rect 4905 21301 4939 21335
rect 4939 21301 4948 21335
rect 4896 21292 4948 21301
rect 7472 21335 7524 21344
rect 7472 21301 7481 21335
rect 7481 21301 7515 21335
rect 7515 21301 7524 21335
rect 7472 21292 7524 21301
rect 7656 21292 7708 21344
rect 7932 21292 7984 21344
rect 14280 21292 14332 21344
rect 14372 21292 14424 21344
rect 16120 21292 16172 21344
rect 16856 21292 16908 21344
rect 19156 21539 19208 21548
rect 19156 21505 19165 21539
rect 19165 21505 19199 21539
rect 19199 21505 19208 21539
rect 19156 21496 19208 21505
rect 17960 21428 18012 21480
rect 19340 21428 19392 21480
rect 21364 21471 21416 21480
rect 21364 21437 21373 21471
rect 21373 21437 21407 21471
rect 21407 21437 21416 21471
rect 21364 21428 21416 21437
rect 21640 21428 21692 21480
rect 24032 21496 24084 21548
rect 23848 21471 23900 21480
rect 18144 21360 18196 21412
rect 20352 21292 20404 21344
rect 20444 21292 20496 21344
rect 21732 21335 21784 21344
rect 21732 21301 21741 21335
rect 21741 21301 21775 21335
rect 21775 21301 21784 21335
rect 21732 21292 21784 21301
rect 23848 21437 23857 21471
rect 23857 21437 23891 21471
rect 23891 21437 23900 21471
rect 23848 21428 23900 21437
rect 24400 21471 24452 21480
rect 24400 21437 24410 21471
rect 24410 21437 24452 21471
rect 24400 21428 24452 21437
rect 25320 21471 25372 21480
rect 25320 21437 25329 21471
rect 25329 21437 25363 21471
rect 25363 21437 25372 21471
rect 25320 21428 25372 21437
rect 21916 21360 21968 21412
rect 22928 21360 22980 21412
rect 22284 21292 22336 21344
rect 7114 21190 7166 21242
rect 7178 21190 7230 21242
rect 7242 21190 7294 21242
rect 7306 21190 7358 21242
rect 7370 21190 7422 21242
rect 13830 21190 13882 21242
rect 13894 21190 13946 21242
rect 13958 21190 14010 21242
rect 14022 21190 14074 21242
rect 14086 21190 14138 21242
rect 20546 21190 20598 21242
rect 20610 21190 20662 21242
rect 20674 21190 20726 21242
rect 20738 21190 20790 21242
rect 20802 21190 20854 21242
rect 27262 21190 27314 21242
rect 27326 21190 27378 21242
rect 27390 21190 27442 21242
rect 27454 21190 27506 21242
rect 27518 21190 27570 21242
rect 2688 21088 2740 21140
rect 3424 21088 3476 21140
rect 5080 21088 5132 21140
rect 7012 21088 7064 21140
rect 848 20952 900 21004
rect 3240 21020 3292 21072
rect 1584 20927 1636 20936
rect 1584 20893 1593 20927
rect 1593 20893 1627 20927
rect 1627 20893 1636 20927
rect 1584 20884 1636 20893
rect 3608 20927 3660 20936
rect 3608 20893 3617 20927
rect 3617 20893 3651 20927
rect 3651 20893 3660 20927
rect 3608 20884 3660 20893
rect 5816 20952 5868 21004
rect 5908 20952 5960 21004
rect 7472 21088 7524 21140
rect 7840 21131 7892 21140
rect 7840 21097 7849 21131
rect 7849 21097 7883 21131
rect 7883 21097 7892 21131
rect 7840 21088 7892 21097
rect 10416 21088 10468 21140
rect 12440 21088 12492 21140
rect 13268 21020 13320 21072
rect 7472 20995 7524 21004
rect 7472 20961 7481 20995
rect 7481 20961 7515 20995
rect 7515 20961 7524 20995
rect 7472 20952 7524 20961
rect 9220 20952 9272 21004
rect 9956 20952 10008 21004
rect 10968 20995 11020 21004
rect 10968 20961 10977 20995
rect 10977 20961 11011 20995
rect 11011 20961 11020 20995
rect 10968 20952 11020 20961
rect 11796 20952 11848 21004
rect 14280 21088 14332 21140
rect 16304 21088 16356 21140
rect 17868 21088 17920 21140
rect 19248 21088 19300 21140
rect 21732 21088 21784 21140
rect 18420 21020 18472 21072
rect 20444 21020 20496 21072
rect 1124 20748 1176 20800
rect 5080 20791 5132 20800
rect 5080 20757 5089 20791
rect 5089 20757 5123 20791
rect 5123 20757 5132 20791
rect 5080 20748 5132 20757
rect 5540 20748 5592 20800
rect 7656 20884 7708 20936
rect 9772 20884 9824 20936
rect 7012 20859 7064 20868
rect 7012 20825 7021 20859
rect 7021 20825 7055 20859
rect 7055 20825 7064 20859
rect 15200 20952 15252 21004
rect 16672 20952 16724 21004
rect 18052 20952 18104 21004
rect 18512 20952 18564 21004
rect 19156 20952 19208 21004
rect 19616 20995 19668 21004
rect 19616 20961 19625 20995
rect 19625 20961 19659 20995
rect 19659 20961 19668 20995
rect 19616 20952 19668 20961
rect 20996 20952 21048 21004
rect 21364 20952 21416 21004
rect 12624 20884 12676 20936
rect 13636 20884 13688 20936
rect 17960 20927 18012 20936
rect 7012 20816 7064 20825
rect 7840 20748 7892 20800
rect 7932 20791 7984 20800
rect 7932 20757 7941 20791
rect 7941 20757 7975 20791
rect 7975 20757 7984 20791
rect 7932 20748 7984 20757
rect 15936 20816 15988 20868
rect 9404 20791 9456 20800
rect 9404 20757 9413 20791
rect 9413 20757 9447 20791
rect 9447 20757 9456 20791
rect 9404 20748 9456 20757
rect 12348 20748 12400 20800
rect 14096 20748 14148 20800
rect 15108 20748 15160 20800
rect 15844 20748 15896 20800
rect 17960 20893 17969 20927
rect 17969 20893 18003 20927
rect 18003 20893 18012 20927
rect 17960 20884 18012 20893
rect 20260 20884 20312 20936
rect 21640 20995 21692 21004
rect 21640 20961 21649 20995
rect 21649 20961 21683 20995
rect 21683 20961 21692 20995
rect 21640 20952 21692 20961
rect 21732 20952 21784 21004
rect 16672 20816 16724 20868
rect 21916 21020 21968 21072
rect 22928 21088 22980 21140
rect 23848 21088 23900 21140
rect 24032 21131 24084 21140
rect 24032 21097 24041 21131
rect 24041 21097 24075 21131
rect 24075 21097 24084 21131
rect 24032 21088 24084 21097
rect 25504 21088 25556 21140
rect 25872 21088 25924 21140
rect 26424 21131 26476 21140
rect 26424 21097 26433 21131
rect 26433 21097 26467 21131
rect 26467 21097 26476 21131
rect 26424 21088 26476 21097
rect 26976 21131 27028 21140
rect 26976 21097 26985 21131
rect 26985 21097 27019 21131
rect 27019 21097 27028 21131
rect 26976 21088 27028 21097
rect 25136 21020 25188 21072
rect 26148 21020 26200 21072
rect 26516 20952 26568 21004
rect 26700 20952 26752 21004
rect 26976 20952 27028 21004
rect 18696 20748 18748 20800
rect 19340 20748 19392 20800
rect 20904 20791 20956 20800
rect 20904 20757 20913 20791
rect 20913 20757 20947 20791
rect 20947 20757 20956 20791
rect 20904 20748 20956 20757
rect 24584 20816 24636 20868
rect 22284 20748 22336 20800
rect 3756 20646 3808 20698
rect 3820 20646 3872 20698
rect 3884 20646 3936 20698
rect 3948 20646 4000 20698
rect 4012 20646 4064 20698
rect 10472 20646 10524 20698
rect 10536 20646 10588 20698
rect 10600 20646 10652 20698
rect 10664 20646 10716 20698
rect 10728 20646 10780 20698
rect 17188 20646 17240 20698
rect 17252 20646 17304 20698
rect 17316 20646 17368 20698
rect 17380 20646 17432 20698
rect 17444 20646 17496 20698
rect 23904 20646 23956 20698
rect 23968 20646 24020 20698
rect 24032 20646 24084 20698
rect 24096 20646 24148 20698
rect 24160 20646 24212 20698
rect 2228 20587 2280 20596
rect 2228 20553 2237 20587
rect 2237 20553 2271 20587
rect 2271 20553 2280 20587
rect 2228 20544 2280 20553
rect 2780 20544 2832 20596
rect 3332 20544 3384 20596
rect 848 20383 900 20392
rect 848 20349 857 20383
rect 857 20349 891 20383
rect 891 20349 900 20383
rect 848 20340 900 20349
rect 1124 20383 1176 20392
rect 1124 20349 1158 20383
rect 1158 20349 1176 20383
rect 1124 20340 1176 20349
rect 3516 20544 3568 20596
rect 3608 20544 3660 20596
rect 4988 20544 5040 20596
rect 3332 20408 3384 20460
rect 5540 20476 5592 20528
rect 2320 20340 2372 20392
rect 3424 20315 3476 20324
rect 3424 20281 3449 20315
rect 3449 20281 3476 20315
rect 3424 20272 3476 20281
rect 2872 20247 2924 20256
rect 2872 20213 2881 20247
rect 2881 20213 2915 20247
rect 2915 20213 2924 20247
rect 2872 20204 2924 20213
rect 4436 20340 4488 20392
rect 3976 20315 4028 20324
rect 3976 20281 4010 20315
rect 4010 20281 4028 20315
rect 3976 20272 4028 20281
rect 6276 20340 6328 20392
rect 7472 20544 7524 20596
rect 7932 20544 7984 20596
rect 8576 20544 8628 20596
rect 14188 20544 14240 20596
rect 14832 20544 14884 20596
rect 9404 20451 9456 20460
rect 9404 20417 9413 20451
rect 9413 20417 9447 20451
rect 9447 20417 9456 20451
rect 9404 20408 9456 20417
rect 9772 20408 9824 20460
rect 10232 20408 10284 20460
rect 11796 20451 11848 20460
rect 11796 20417 11805 20451
rect 11805 20417 11839 20451
rect 11839 20417 11848 20451
rect 11796 20408 11848 20417
rect 7748 20340 7800 20392
rect 12348 20340 12400 20392
rect 9404 20272 9456 20324
rect 5264 20204 5316 20256
rect 9036 20247 9088 20256
rect 9036 20213 9045 20247
rect 9045 20213 9079 20247
rect 9079 20213 9088 20247
rect 9036 20204 9088 20213
rect 10048 20247 10100 20256
rect 10048 20213 10057 20247
rect 10057 20213 10091 20247
rect 10091 20213 10100 20247
rect 10048 20204 10100 20213
rect 11060 20272 11112 20324
rect 11336 20272 11388 20324
rect 14464 20476 14516 20528
rect 13268 20408 13320 20460
rect 13636 20383 13688 20392
rect 11152 20204 11204 20256
rect 12532 20204 12584 20256
rect 13084 20204 13136 20256
rect 13636 20349 13645 20383
rect 13645 20349 13679 20383
rect 13679 20349 13688 20383
rect 13636 20340 13688 20349
rect 14188 20408 14240 20460
rect 14372 20408 14424 20460
rect 14096 20383 14148 20392
rect 14096 20349 14105 20383
rect 14105 20349 14139 20383
rect 14139 20349 14148 20383
rect 14096 20340 14148 20349
rect 16856 20451 16908 20460
rect 16856 20417 16865 20451
rect 16865 20417 16899 20451
rect 16899 20417 16908 20451
rect 16856 20408 16908 20417
rect 18144 20587 18196 20596
rect 18144 20553 18153 20587
rect 18153 20553 18187 20587
rect 18187 20553 18196 20587
rect 18144 20544 18196 20553
rect 19984 20544 20036 20596
rect 17684 20340 17736 20392
rect 17960 20383 18012 20392
rect 17960 20349 17969 20383
rect 17969 20349 18003 20383
rect 18003 20349 18012 20383
rect 17960 20340 18012 20349
rect 18512 20340 18564 20392
rect 18972 20340 19024 20392
rect 20812 20476 20864 20528
rect 15844 20272 15896 20324
rect 15936 20315 15988 20324
rect 15936 20281 15954 20315
rect 15954 20281 15988 20315
rect 15936 20272 15988 20281
rect 19340 20272 19392 20324
rect 14648 20204 14700 20256
rect 14740 20247 14792 20256
rect 14740 20213 14749 20247
rect 14749 20213 14783 20247
rect 14783 20213 14792 20247
rect 14740 20204 14792 20213
rect 14832 20247 14884 20256
rect 14832 20213 14841 20247
rect 14841 20213 14875 20247
rect 14875 20213 14884 20247
rect 14832 20204 14884 20213
rect 15292 20204 15344 20256
rect 19524 20204 19576 20256
rect 20812 20340 20864 20392
rect 20904 20340 20956 20392
rect 22284 20383 22336 20392
rect 22284 20349 22293 20383
rect 22293 20349 22327 20383
rect 22327 20349 22336 20383
rect 22284 20340 22336 20349
rect 23020 20340 23072 20392
rect 23664 20383 23716 20392
rect 23664 20349 23673 20383
rect 23673 20349 23707 20383
rect 23707 20349 23716 20383
rect 23664 20340 23716 20349
rect 26240 20340 26292 20392
rect 26516 20340 26568 20392
rect 25596 20272 25648 20324
rect 22100 20204 22152 20256
rect 22192 20204 22244 20256
rect 23480 20247 23532 20256
rect 23480 20213 23489 20247
rect 23489 20213 23523 20247
rect 23523 20213 23532 20247
rect 23480 20204 23532 20213
rect 27068 20247 27120 20256
rect 27068 20213 27077 20247
rect 27077 20213 27111 20247
rect 27111 20213 27120 20247
rect 27068 20204 27120 20213
rect 7114 20102 7166 20154
rect 7178 20102 7230 20154
rect 7242 20102 7294 20154
rect 7306 20102 7358 20154
rect 7370 20102 7422 20154
rect 13830 20102 13882 20154
rect 13894 20102 13946 20154
rect 13958 20102 14010 20154
rect 14022 20102 14074 20154
rect 14086 20102 14138 20154
rect 20546 20102 20598 20154
rect 20610 20102 20662 20154
rect 20674 20102 20726 20154
rect 20738 20102 20790 20154
rect 20802 20102 20854 20154
rect 27262 20102 27314 20154
rect 27326 20102 27378 20154
rect 27390 20102 27442 20154
rect 27454 20102 27506 20154
rect 27518 20102 27570 20154
rect 3976 20000 4028 20052
rect 5080 20000 5132 20052
rect 5264 20000 5316 20052
rect 7656 20043 7708 20052
rect 7656 20009 7665 20043
rect 7665 20009 7699 20043
rect 7699 20009 7708 20043
rect 7656 20000 7708 20009
rect 8484 20000 8536 20052
rect 8944 20000 8996 20052
rect 9036 20000 9088 20052
rect 9220 20043 9272 20052
rect 9220 20009 9229 20043
rect 9229 20009 9263 20043
rect 9263 20009 9272 20043
rect 9220 20000 9272 20009
rect 9956 20000 10008 20052
rect 10968 20000 11020 20052
rect 11060 20043 11112 20052
rect 11060 20009 11069 20043
rect 11069 20009 11103 20043
rect 11103 20009 11112 20043
rect 11060 20000 11112 20009
rect 12624 20043 12676 20052
rect 12624 20009 12633 20043
rect 12633 20009 12667 20043
rect 12667 20009 12676 20043
rect 12624 20000 12676 20009
rect 12992 20000 13044 20052
rect 13084 20043 13136 20052
rect 13084 20009 13093 20043
rect 13093 20009 13127 20043
rect 13127 20009 13136 20043
rect 13084 20000 13136 20009
rect 14188 20000 14240 20052
rect 14648 20000 14700 20052
rect 15200 20043 15252 20052
rect 15200 20009 15209 20043
rect 15209 20009 15243 20043
rect 15243 20009 15252 20043
rect 15200 20000 15252 20009
rect 15568 20043 15620 20052
rect 15568 20009 15577 20043
rect 15577 20009 15611 20043
rect 15611 20009 15620 20043
rect 15568 20000 15620 20009
rect 2872 19932 2924 19984
rect 1400 19907 1452 19916
rect 1400 19873 1409 19907
rect 1409 19873 1443 19907
rect 1443 19873 1452 19907
rect 1400 19864 1452 19873
rect 4436 19932 4488 19984
rect 6552 19932 6604 19984
rect 4988 19907 5040 19916
rect 4988 19873 4997 19907
rect 4997 19873 5031 19907
rect 5031 19873 5040 19907
rect 4988 19864 5040 19873
rect 7840 19864 7892 19916
rect 11336 19975 11388 19984
rect 11336 19941 11345 19975
rect 11345 19941 11379 19975
rect 11379 19941 11388 19975
rect 11336 19932 11388 19941
rect 5448 19796 5500 19848
rect 7564 19839 7616 19848
rect 7564 19805 7573 19839
rect 7573 19805 7607 19839
rect 7607 19805 7616 19839
rect 7564 19796 7616 19805
rect 8576 19796 8628 19848
rect 1124 19660 1176 19712
rect 4896 19660 4948 19712
rect 6368 19703 6420 19712
rect 6368 19669 6377 19703
rect 6377 19669 6411 19703
rect 6411 19669 6420 19703
rect 6368 19660 6420 19669
rect 7012 19660 7064 19712
rect 8944 19907 8996 19916
rect 8944 19873 8953 19907
rect 8953 19873 8987 19907
rect 8987 19873 8996 19907
rect 8944 19864 8996 19873
rect 9680 19907 9732 19916
rect 9680 19873 9689 19907
rect 9689 19873 9723 19907
rect 9723 19873 9732 19907
rect 9680 19864 9732 19873
rect 10048 19864 10100 19916
rect 8852 19728 8904 19780
rect 9588 19728 9640 19780
rect 11244 19907 11296 19916
rect 11244 19873 11253 19907
rect 11253 19873 11287 19907
rect 11287 19873 11296 19907
rect 11244 19864 11296 19873
rect 11428 19907 11480 19916
rect 11428 19873 11437 19907
rect 11437 19873 11471 19907
rect 11471 19873 11480 19907
rect 11428 19864 11480 19873
rect 12532 19864 12584 19916
rect 15292 19932 15344 19984
rect 12992 19907 13044 19916
rect 12992 19873 13001 19907
rect 13001 19873 13035 19907
rect 13035 19873 13044 19907
rect 12992 19864 13044 19873
rect 13636 19864 13688 19916
rect 14188 19907 14240 19916
rect 14188 19873 14197 19907
rect 14197 19873 14231 19907
rect 14231 19873 14240 19907
rect 14188 19864 14240 19873
rect 16028 19864 16080 19916
rect 16948 19907 17000 19916
rect 16948 19873 16957 19907
rect 16957 19873 16991 19907
rect 16991 19873 17000 19907
rect 16948 19864 17000 19873
rect 18972 20000 19024 20052
rect 19340 20000 19392 20052
rect 19524 20000 19576 20052
rect 19616 20000 19668 20052
rect 20996 20000 21048 20052
rect 18052 19932 18104 19984
rect 25320 19932 25372 19984
rect 14648 19796 14700 19848
rect 14096 19728 14148 19780
rect 10968 19660 11020 19712
rect 11152 19660 11204 19712
rect 14556 19660 14608 19712
rect 15016 19660 15068 19712
rect 16120 19703 16172 19712
rect 16120 19669 16129 19703
rect 16129 19669 16163 19703
rect 16163 19669 16172 19703
rect 16120 19660 16172 19669
rect 19800 19864 19852 19916
rect 20076 19907 20128 19916
rect 20076 19873 20085 19907
rect 20085 19873 20119 19907
rect 20119 19873 20128 19907
rect 20076 19864 20128 19873
rect 20168 19864 20220 19916
rect 19616 19796 19668 19848
rect 20260 19839 20312 19848
rect 20260 19805 20269 19839
rect 20269 19805 20303 19839
rect 20303 19805 20312 19839
rect 20260 19796 20312 19805
rect 20904 19907 20956 19916
rect 20904 19873 20913 19907
rect 20913 19873 20947 19907
rect 20947 19873 20956 19907
rect 20904 19864 20956 19873
rect 22192 19907 22244 19916
rect 22192 19873 22201 19907
rect 22201 19873 22235 19907
rect 22235 19873 22244 19907
rect 22192 19864 22244 19873
rect 27068 19907 27120 19916
rect 27068 19873 27077 19907
rect 27077 19873 27111 19907
rect 27111 19873 27120 19907
rect 27068 19864 27120 19873
rect 21180 19796 21232 19848
rect 21824 19839 21876 19848
rect 21824 19805 21833 19839
rect 21833 19805 21867 19839
rect 21867 19805 21876 19839
rect 21824 19796 21876 19805
rect 17960 19660 18012 19712
rect 18604 19703 18656 19712
rect 18604 19669 18613 19703
rect 18613 19669 18647 19703
rect 18647 19669 18656 19703
rect 18604 19660 18656 19669
rect 19892 19703 19944 19712
rect 19892 19669 19901 19703
rect 19901 19669 19935 19703
rect 19935 19669 19944 19703
rect 19892 19660 19944 19669
rect 20352 19703 20404 19712
rect 20352 19669 20361 19703
rect 20361 19669 20395 19703
rect 20395 19669 20404 19703
rect 20352 19660 20404 19669
rect 22100 19728 22152 19780
rect 22376 19728 22428 19780
rect 21088 19660 21140 19712
rect 22652 19660 22704 19712
rect 23020 19660 23072 19712
rect 25504 19660 25556 19712
rect 26424 19703 26476 19712
rect 26424 19669 26433 19703
rect 26433 19669 26467 19703
rect 26467 19669 26476 19703
rect 26424 19660 26476 19669
rect 3756 19558 3808 19610
rect 3820 19558 3872 19610
rect 3884 19558 3936 19610
rect 3948 19558 4000 19610
rect 4012 19558 4064 19610
rect 10472 19558 10524 19610
rect 10536 19558 10588 19610
rect 10600 19558 10652 19610
rect 10664 19558 10716 19610
rect 10728 19558 10780 19610
rect 17188 19558 17240 19610
rect 17252 19558 17304 19610
rect 17316 19558 17368 19610
rect 17380 19558 17432 19610
rect 17444 19558 17496 19610
rect 23904 19558 23956 19610
rect 23968 19558 24020 19610
rect 24032 19558 24084 19610
rect 24096 19558 24148 19610
rect 24160 19558 24212 19610
rect 4436 19456 4488 19508
rect 9220 19499 9272 19508
rect 9220 19465 9229 19499
rect 9229 19465 9263 19499
rect 9263 19465 9272 19499
rect 9220 19456 9272 19465
rect 8944 19388 8996 19440
rect 11060 19456 11112 19508
rect 11428 19456 11480 19508
rect 12072 19456 12124 19508
rect 13452 19456 13504 19508
rect 14096 19499 14148 19508
rect 14096 19465 14105 19499
rect 14105 19465 14139 19499
rect 14139 19465 14148 19499
rect 14096 19456 14148 19465
rect 14740 19456 14792 19508
rect 15292 19456 15344 19508
rect 16028 19456 16080 19508
rect 16948 19456 17000 19508
rect 19340 19456 19392 19508
rect 23572 19456 23624 19508
rect 23664 19499 23716 19508
rect 23664 19465 23673 19499
rect 23673 19465 23707 19499
rect 23707 19465 23716 19499
rect 23664 19456 23716 19465
rect 25596 19456 25648 19508
rect 848 19295 900 19304
rect 848 19261 857 19295
rect 857 19261 891 19295
rect 891 19261 900 19295
rect 848 19252 900 19261
rect 1124 19295 1176 19304
rect 1124 19261 1158 19295
rect 1158 19261 1176 19295
rect 1124 19252 1176 19261
rect 2596 19295 2648 19304
rect 2596 19261 2605 19295
rect 2605 19261 2639 19295
rect 2639 19261 2648 19295
rect 2596 19252 2648 19261
rect 2872 19252 2924 19304
rect 3148 19252 3200 19304
rect 4160 19252 4212 19304
rect 1032 19116 1084 19168
rect 3332 19184 3384 19236
rect 4620 19295 4672 19304
rect 4620 19261 4629 19295
rect 4629 19261 4663 19295
rect 4663 19261 4672 19295
rect 4620 19252 4672 19261
rect 2780 19116 2832 19168
rect 4988 19227 5040 19236
rect 4988 19193 4997 19227
rect 4997 19193 5031 19227
rect 5031 19193 5040 19227
rect 4988 19184 5040 19193
rect 5080 19227 5132 19236
rect 5080 19193 5089 19227
rect 5089 19193 5123 19227
rect 5123 19193 5132 19227
rect 5080 19184 5132 19193
rect 4252 19116 4304 19168
rect 6092 19252 6144 19304
rect 6276 19252 6328 19304
rect 8024 19252 8076 19304
rect 8484 19252 8536 19304
rect 9404 19320 9456 19372
rect 8668 19295 8720 19304
rect 8668 19261 8677 19295
rect 8677 19261 8711 19295
rect 8711 19261 8720 19295
rect 8668 19252 8720 19261
rect 8760 19295 8812 19304
rect 8760 19261 8769 19295
rect 8769 19261 8803 19295
rect 8803 19261 8812 19295
rect 8760 19252 8812 19261
rect 8944 19252 8996 19304
rect 12256 19388 12308 19440
rect 11244 19320 11296 19372
rect 15016 19388 15068 19440
rect 15200 19388 15252 19440
rect 5908 19227 5960 19236
rect 5908 19193 5917 19227
rect 5917 19193 5951 19227
rect 5951 19193 5960 19227
rect 5908 19184 5960 19193
rect 8208 19116 8260 19168
rect 8392 19159 8444 19168
rect 8392 19125 8401 19159
rect 8401 19125 8435 19159
rect 8435 19125 8444 19159
rect 8392 19116 8444 19125
rect 8852 19116 8904 19168
rect 8944 19116 8996 19168
rect 9128 19116 9180 19168
rect 9404 19159 9456 19168
rect 9404 19125 9413 19159
rect 9413 19125 9447 19159
rect 9447 19125 9456 19159
rect 9404 19116 9456 19125
rect 10416 19295 10468 19304
rect 10416 19261 10425 19295
rect 10425 19261 10459 19295
rect 10459 19261 10468 19295
rect 10416 19252 10468 19261
rect 10508 19295 10560 19304
rect 10508 19261 10517 19295
rect 10517 19261 10551 19295
rect 10551 19261 10560 19295
rect 10508 19252 10560 19261
rect 11060 19252 11112 19304
rect 9864 19227 9916 19236
rect 9864 19193 9873 19227
rect 9873 19193 9907 19227
rect 9907 19193 9916 19227
rect 9864 19184 9916 19193
rect 12256 19295 12308 19304
rect 12256 19261 12265 19295
rect 12265 19261 12299 19295
rect 12299 19261 12308 19295
rect 12256 19252 12308 19261
rect 12624 19252 12676 19304
rect 12808 19252 12860 19304
rect 9956 19116 10008 19168
rect 12072 19227 12124 19236
rect 12072 19193 12081 19227
rect 12081 19193 12115 19227
rect 12115 19193 12124 19227
rect 12072 19184 12124 19193
rect 10324 19116 10376 19168
rect 11152 19116 11204 19168
rect 11980 19116 12032 19168
rect 12256 19116 12308 19168
rect 13544 19252 13596 19304
rect 14924 19184 14976 19236
rect 13544 19116 13596 19168
rect 13728 19116 13780 19168
rect 14280 19159 14332 19168
rect 14280 19125 14289 19159
rect 14289 19125 14323 19159
rect 14323 19125 14332 19159
rect 14280 19116 14332 19125
rect 15108 19116 15160 19168
rect 15384 19363 15436 19372
rect 15384 19329 15393 19363
rect 15393 19329 15427 19363
rect 15427 19329 15436 19363
rect 15384 19320 15436 19329
rect 15844 19363 15896 19372
rect 15844 19329 15853 19363
rect 15853 19329 15887 19363
rect 15887 19329 15896 19363
rect 15844 19320 15896 19329
rect 17868 19363 17920 19372
rect 17868 19329 17877 19363
rect 17877 19329 17911 19363
rect 17911 19329 17920 19363
rect 17868 19320 17920 19329
rect 18604 19388 18656 19440
rect 22744 19388 22796 19440
rect 19616 19320 19668 19372
rect 21824 19320 21876 19372
rect 22100 19363 22152 19372
rect 22100 19329 22109 19363
rect 22109 19329 22143 19363
rect 22143 19329 22152 19363
rect 22100 19320 22152 19329
rect 15476 19252 15528 19304
rect 15568 19295 15620 19304
rect 15568 19261 15577 19295
rect 15577 19261 15611 19295
rect 15611 19261 15620 19295
rect 15568 19252 15620 19261
rect 16120 19295 16172 19304
rect 16120 19261 16154 19295
rect 16154 19261 16172 19295
rect 16120 19252 16172 19261
rect 17592 19252 17644 19304
rect 18052 19252 18104 19304
rect 18328 19295 18380 19304
rect 18328 19261 18337 19295
rect 18337 19261 18371 19295
rect 18371 19261 18380 19295
rect 18328 19252 18380 19261
rect 19708 19252 19760 19304
rect 22284 19295 22336 19304
rect 22284 19261 22293 19295
rect 22293 19261 22327 19295
rect 22327 19261 22336 19295
rect 22284 19252 22336 19261
rect 22468 19295 22520 19304
rect 22468 19261 22477 19295
rect 22477 19261 22511 19295
rect 22511 19261 22520 19295
rect 22468 19252 22520 19261
rect 22560 19295 22612 19304
rect 22560 19261 22569 19295
rect 22569 19261 22603 19295
rect 22603 19261 22612 19295
rect 22560 19252 22612 19261
rect 24032 19295 24084 19304
rect 16488 19116 16540 19168
rect 19984 19184 20036 19236
rect 24032 19261 24041 19295
rect 24041 19261 24075 19295
rect 24075 19261 24084 19295
rect 24032 19252 24084 19261
rect 24492 19252 24544 19304
rect 20444 19116 20496 19168
rect 20996 19159 21048 19168
rect 20996 19125 21005 19159
rect 21005 19125 21039 19159
rect 21039 19125 21048 19159
rect 20996 19116 21048 19125
rect 22836 19159 22888 19168
rect 22836 19125 22845 19159
rect 22845 19125 22879 19159
rect 22879 19125 22888 19159
rect 22836 19116 22888 19125
rect 23112 19159 23164 19168
rect 23112 19125 23121 19159
rect 23121 19125 23155 19159
rect 23155 19125 23164 19159
rect 23112 19116 23164 19125
rect 23388 19184 23440 19236
rect 25228 19252 25280 19304
rect 25780 19252 25832 19304
rect 26240 19252 26292 19304
rect 24676 19116 24728 19168
rect 24860 19116 24912 19168
rect 25872 19184 25924 19236
rect 26424 19116 26476 19168
rect 7114 19014 7166 19066
rect 7178 19014 7230 19066
rect 7242 19014 7294 19066
rect 7306 19014 7358 19066
rect 7370 19014 7422 19066
rect 13830 19014 13882 19066
rect 13894 19014 13946 19066
rect 13958 19014 14010 19066
rect 14022 19014 14074 19066
rect 14086 19014 14138 19066
rect 20546 19014 20598 19066
rect 20610 19014 20662 19066
rect 20674 19014 20726 19066
rect 20738 19014 20790 19066
rect 20802 19014 20854 19066
rect 27262 19014 27314 19066
rect 27326 19014 27378 19066
rect 27390 19014 27442 19066
rect 27454 19014 27506 19066
rect 27518 19014 27570 19066
rect 1400 18912 1452 18964
rect 1952 18955 2004 18964
rect 1952 18921 1961 18955
rect 1961 18921 1995 18955
rect 1995 18921 2004 18955
rect 1952 18912 2004 18921
rect 2596 18912 2648 18964
rect 5080 18912 5132 18964
rect 7564 18955 7616 18964
rect 7564 18921 7573 18955
rect 7573 18921 7607 18955
rect 7607 18921 7616 18955
rect 7564 18912 7616 18921
rect 848 18776 900 18828
rect 1032 18819 1084 18828
rect 1032 18785 1041 18819
rect 1041 18785 1075 18819
rect 1075 18785 1084 18819
rect 1032 18776 1084 18785
rect 2228 18776 2280 18828
rect 2780 18844 2832 18896
rect 9220 18912 9272 18964
rect 9404 18912 9456 18964
rect 8668 18887 8720 18896
rect 4252 18819 4304 18828
rect 4252 18785 4286 18819
rect 4286 18785 4304 18819
rect 4252 18776 4304 18785
rect 5448 18819 5500 18828
rect 5448 18785 5457 18819
rect 5457 18785 5491 18819
rect 5491 18785 5500 18819
rect 5448 18776 5500 18785
rect 8668 18853 8677 18887
rect 8677 18853 8711 18887
rect 8711 18853 8720 18887
rect 8668 18844 8720 18853
rect 6276 18776 6328 18828
rect 6460 18819 6512 18828
rect 6460 18785 6494 18819
rect 6494 18785 6512 18819
rect 6460 18776 6512 18785
rect 1400 18683 1452 18692
rect 1400 18649 1409 18683
rect 1409 18649 1443 18683
rect 1443 18649 1452 18683
rect 1400 18640 1452 18649
rect 3608 18572 3660 18624
rect 4160 18572 4212 18624
rect 5816 18640 5868 18692
rect 6092 18572 6144 18624
rect 8576 18776 8628 18828
rect 8760 18819 8812 18828
rect 8760 18785 8769 18819
rect 8769 18785 8803 18819
rect 8803 18785 8812 18819
rect 11060 18955 11112 18964
rect 11060 18921 11069 18955
rect 11069 18921 11103 18955
rect 11103 18921 11112 18955
rect 11060 18912 11112 18921
rect 12348 18912 12400 18964
rect 13728 18912 13780 18964
rect 14280 18912 14332 18964
rect 15568 18912 15620 18964
rect 16488 18912 16540 18964
rect 8760 18776 8812 18785
rect 8208 18640 8260 18692
rect 8300 18640 8352 18692
rect 9036 18640 9088 18692
rect 6920 18572 6972 18624
rect 7840 18615 7892 18624
rect 7840 18581 7849 18615
rect 7849 18581 7883 18615
rect 7883 18581 7892 18615
rect 7840 18572 7892 18581
rect 10232 18819 10284 18828
rect 10232 18785 10241 18819
rect 10241 18785 10275 18819
rect 10275 18785 10284 18819
rect 10232 18776 10284 18785
rect 12164 18819 12216 18828
rect 12164 18785 12193 18819
rect 12193 18785 12216 18819
rect 12164 18776 12216 18785
rect 12440 18819 12492 18828
rect 12440 18785 12449 18819
rect 12449 18785 12483 18819
rect 12483 18785 12492 18819
rect 12440 18776 12492 18785
rect 12532 18819 12584 18828
rect 12532 18785 12541 18819
rect 12541 18785 12575 18819
rect 12575 18785 12584 18819
rect 12532 18776 12584 18785
rect 14924 18844 14976 18896
rect 17592 18912 17644 18964
rect 20444 18912 20496 18964
rect 20996 18912 21048 18964
rect 21916 18912 21968 18964
rect 10232 18640 10284 18692
rect 10416 18640 10468 18692
rect 15384 18776 15436 18828
rect 14556 18708 14608 18760
rect 14648 18708 14700 18760
rect 9312 18572 9364 18624
rect 10508 18572 10560 18624
rect 14280 18572 14332 18624
rect 17040 18819 17092 18828
rect 17040 18785 17049 18819
rect 17049 18785 17083 18819
rect 17083 18785 17092 18819
rect 17040 18776 17092 18785
rect 17960 18844 18012 18896
rect 19340 18844 19392 18896
rect 20352 18844 20404 18896
rect 22560 18955 22612 18964
rect 22560 18921 22569 18955
rect 22569 18921 22603 18955
rect 22603 18921 22612 18955
rect 22560 18912 22612 18921
rect 23112 18912 23164 18964
rect 24032 18912 24084 18964
rect 24676 18955 24728 18964
rect 24676 18921 24685 18955
rect 24685 18921 24719 18955
rect 24719 18921 24728 18955
rect 24676 18912 24728 18921
rect 20260 18708 20312 18760
rect 20904 18819 20956 18828
rect 20904 18785 20913 18819
rect 20913 18785 20947 18819
rect 20947 18785 20956 18819
rect 20904 18776 20956 18785
rect 21088 18751 21140 18760
rect 21088 18717 21097 18751
rect 21097 18717 21131 18751
rect 21131 18717 21140 18751
rect 21088 18708 21140 18717
rect 18236 18572 18288 18624
rect 18696 18615 18748 18624
rect 18696 18581 18705 18615
rect 18705 18581 18739 18615
rect 18739 18581 18748 18615
rect 18696 18572 18748 18581
rect 22192 18819 22244 18828
rect 22192 18785 22201 18819
rect 22201 18785 22235 18819
rect 22235 18785 22244 18819
rect 22192 18776 22244 18785
rect 23480 18844 23532 18896
rect 24860 18844 24912 18896
rect 23020 18776 23072 18828
rect 24308 18776 24360 18828
rect 24492 18708 24544 18760
rect 22836 18640 22888 18692
rect 24860 18640 24912 18692
rect 25872 18955 25924 18964
rect 25872 18921 25881 18955
rect 25881 18921 25915 18955
rect 25915 18921 25924 18955
rect 25872 18912 25924 18921
rect 27068 18708 27120 18760
rect 19708 18572 19760 18624
rect 20444 18615 20496 18624
rect 20444 18581 20453 18615
rect 20453 18581 20487 18615
rect 20487 18581 20496 18615
rect 20444 18572 20496 18581
rect 21180 18572 21232 18624
rect 22192 18572 22244 18624
rect 24768 18572 24820 18624
rect 25412 18615 25464 18624
rect 25412 18581 25421 18615
rect 25421 18581 25455 18615
rect 25455 18581 25464 18615
rect 25412 18572 25464 18581
rect 3756 18470 3808 18522
rect 3820 18470 3872 18522
rect 3884 18470 3936 18522
rect 3948 18470 4000 18522
rect 4012 18470 4064 18522
rect 10472 18470 10524 18522
rect 10536 18470 10588 18522
rect 10600 18470 10652 18522
rect 10664 18470 10716 18522
rect 10728 18470 10780 18522
rect 17188 18470 17240 18522
rect 17252 18470 17304 18522
rect 17316 18470 17368 18522
rect 17380 18470 17432 18522
rect 17444 18470 17496 18522
rect 23904 18470 23956 18522
rect 23968 18470 24020 18522
rect 24032 18470 24084 18522
rect 24096 18470 24148 18522
rect 24160 18470 24212 18522
rect 2872 18368 2924 18420
rect 2412 18300 2464 18352
rect 1952 18232 2004 18284
rect 3056 18300 3108 18352
rect 3148 18300 3200 18352
rect 3424 18300 3476 18352
rect 3608 18300 3660 18352
rect 6460 18368 6512 18420
rect 8392 18368 8444 18420
rect 9956 18368 10008 18420
rect 12440 18411 12492 18420
rect 12440 18377 12449 18411
rect 12449 18377 12483 18411
rect 12483 18377 12492 18411
rect 12440 18368 12492 18377
rect 15108 18411 15160 18420
rect 15108 18377 15117 18411
rect 15117 18377 15151 18411
rect 15151 18377 15160 18411
rect 15108 18368 15160 18377
rect 16212 18368 16264 18420
rect 17040 18368 17092 18420
rect 1400 18207 1452 18216
rect 1400 18173 1409 18207
rect 1409 18173 1443 18207
rect 1443 18173 1452 18207
rect 1400 18164 1452 18173
rect 2228 18164 2280 18216
rect 3608 18164 3660 18216
rect 5080 18164 5132 18216
rect 5816 18207 5868 18216
rect 5816 18173 5825 18207
rect 5825 18173 5859 18207
rect 5859 18173 5868 18207
rect 6920 18232 6972 18284
rect 7840 18300 7892 18352
rect 5816 18164 5868 18173
rect 6368 18164 6420 18216
rect 6736 18164 6788 18216
rect 8484 18164 8536 18216
rect 8944 18300 8996 18352
rect 9036 18300 9088 18352
rect 9588 18300 9640 18352
rect 9680 18232 9732 18284
rect 11060 18275 11112 18284
rect 8944 18207 8996 18216
rect 8944 18173 8953 18207
rect 8953 18173 8987 18207
rect 8987 18173 8996 18207
rect 8944 18164 8996 18173
rect 9036 18207 9088 18216
rect 9036 18173 9045 18207
rect 9045 18173 9079 18207
rect 9079 18173 9088 18207
rect 9036 18164 9088 18173
rect 11060 18241 11069 18275
rect 11069 18241 11103 18275
rect 11103 18241 11112 18275
rect 11060 18232 11112 18241
rect 15016 18232 15068 18284
rect 10048 18207 10100 18216
rect 10048 18173 10057 18207
rect 10057 18173 10091 18207
rect 10091 18173 10100 18207
rect 10048 18164 10100 18173
rect 8852 18096 8904 18148
rect 11612 18164 11664 18216
rect 13268 18164 13320 18216
rect 15476 18164 15528 18216
rect 14188 18096 14240 18148
rect 15108 18096 15160 18148
rect 15200 18139 15252 18148
rect 15200 18105 15209 18139
rect 15209 18105 15243 18139
rect 15243 18105 15252 18139
rect 15200 18096 15252 18105
rect 17868 18232 17920 18284
rect 19708 18368 19760 18420
rect 20168 18368 20220 18420
rect 20996 18368 21048 18420
rect 21088 18368 21140 18420
rect 16856 18164 16908 18216
rect 18512 18164 18564 18216
rect 19432 18232 19484 18284
rect 19892 18164 19944 18216
rect 20444 18164 20496 18216
rect 1676 18071 1728 18080
rect 1676 18037 1685 18071
rect 1685 18037 1719 18071
rect 1719 18037 1728 18071
rect 1676 18028 1728 18037
rect 1768 18071 1820 18080
rect 1768 18037 1777 18071
rect 1777 18037 1811 18071
rect 1811 18037 1820 18071
rect 1768 18028 1820 18037
rect 2320 18028 2372 18080
rect 6920 18028 6972 18080
rect 7012 18028 7064 18080
rect 8668 18028 8720 18080
rect 9220 18028 9272 18080
rect 9496 18071 9548 18080
rect 9496 18037 9505 18071
rect 9505 18037 9539 18071
rect 9539 18037 9548 18071
rect 9496 18028 9548 18037
rect 22284 18368 22336 18420
rect 22468 18368 22520 18420
rect 22744 18368 22796 18420
rect 22836 18368 22888 18420
rect 23572 18368 23624 18420
rect 24124 18368 24176 18420
rect 25412 18368 25464 18420
rect 24308 18300 24360 18352
rect 24492 18300 24544 18352
rect 21916 18164 21968 18216
rect 16764 18028 16816 18080
rect 18144 18071 18196 18080
rect 18144 18037 18153 18071
rect 18153 18037 18187 18071
rect 18187 18037 18196 18071
rect 18144 18028 18196 18037
rect 18696 18028 18748 18080
rect 21180 18028 21232 18080
rect 22192 18139 22244 18148
rect 22192 18105 22201 18139
rect 22201 18105 22235 18139
rect 22235 18105 22244 18139
rect 22192 18096 22244 18105
rect 23112 18164 23164 18216
rect 23204 18207 23256 18216
rect 23204 18173 23213 18207
rect 23213 18173 23247 18207
rect 23247 18173 23256 18207
rect 23204 18164 23256 18173
rect 23296 18207 23348 18216
rect 23296 18173 23305 18207
rect 23305 18173 23339 18207
rect 23339 18173 23348 18207
rect 23296 18164 23348 18173
rect 24124 18207 24176 18216
rect 24124 18173 24133 18207
rect 24133 18173 24167 18207
rect 24167 18173 24176 18207
rect 24124 18164 24176 18173
rect 25780 18164 25832 18216
rect 25964 18139 26016 18148
rect 25964 18105 25998 18139
rect 25998 18105 26016 18139
rect 25964 18096 26016 18105
rect 25044 18028 25096 18080
rect 7114 17926 7166 17978
rect 7178 17926 7230 17978
rect 7242 17926 7294 17978
rect 7306 17926 7358 17978
rect 7370 17926 7422 17978
rect 13830 17926 13882 17978
rect 13894 17926 13946 17978
rect 13958 17926 14010 17978
rect 14022 17926 14074 17978
rect 14086 17926 14138 17978
rect 20546 17926 20598 17978
rect 20610 17926 20662 17978
rect 20674 17926 20726 17978
rect 20738 17926 20790 17978
rect 20802 17926 20854 17978
rect 27262 17926 27314 17978
rect 27326 17926 27378 17978
rect 27390 17926 27442 17978
rect 27454 17926 27506 17978
rect 27518 17926 27570 17978
rect 1768 17824 1820 17876
rect 3424 17756 3476 17808
rect 3516 17756 3568 17808
rect 848 17731 900 17740
rect 848 17697 857 17731
rect 857 17697 891 17731
rect 891 17697 900 17731
rect 848 17688 900 17697
rect 1400 17688 1452 17740
rect 2780 17552 2832 17604
rect 3424 17663 3476 17672
rect 3424 17629 3433 17663
rect 3433 17629 3467 17663
rect 3467 17629 3476 17663
rect 3424 17620 3476 17629
rect 3608 17731 3660 17740
rect 3608 17697 3617 17731
rect 3617 17697 3651 17731
rect 3651 17697 3660 17731
rect 3608 17688 3660 17697
rect 4620 17824 4672 17876
rect 4896 17824 4948 17876
rect 8300 17824 8352 17876
rect 8668 17824 8720 17876
rect 9128 17824 9180 17876
rect 9496 17824 9548 17876
rect 9680 17824 9732 17876
rect 11060 17824 11112 17876
rect 13176 17824 13228 17876
rect 5080 17756 5132 17808
rect 4620 17731 4672 17740
rect 4620 17697 4629 17731
rect 4629 17697 4663 17731
rect 4663 17697 4672 17731
rect 4620 17688 4672 17697
rect 4988 17731 5040 17740
rect 4988 17697 4997 17731
rect 4997 17697 5031 17731
rect 5031 17697 5040 17731
rect 4988 17688 5040 17697
rect 6276 17688 6328 17740
rect 6644 17731 6696 17740
rect 6644 17697 6678 17731
rect 6678 17697 6696 17731
rect 6644 17688 6696 17697
rect 4160 17552 4212 17604
rect 5356 17552 5408 17604
rect 8484 17688 8536 17740
rect 8760 17688 8812 17740
rect 8944 17731 8996 17740
rect 8944 17697 8953 17731
rect 8953 17697 8987 17731
rect 8987 17697 8996 17731
rect 8944 17688 8996 17697
rect 9128 17731 9180 17740
rect 9128 17697 9137 17731
rect 9137 17697 9171 17731
rect 9171 17697 9180 17731
rect 9128 17688 9180 17697
rect 9220 17731 9272 17740
rect 9220 17697 9229 17731
rect 9229 17697 9263 17731
rect 9263 17697 9272 17731
rect 9220 17688 9272 17697
rect 9312 17688 9364 17740
rect 9772 17688 9824 17740
rect 10324 17688 10376 17740
rect 10140 17620 10192 17672
rect 9220 17552 9272 17604
rect 10876 17688 10928 17740
rect 10876 17552 10928 17604
rect 3332 17484 3384 17536
rect 4436 17527 4488 17536
rect 4436 17493 4445 17527
rect 4445 17493 4479 17527
rect 4479 17493 4488 17527
rect 4436 17484 4488 17493
rect 7932 17484 7984 17536
rect 9128 17484 9180 17536
rect 10232 17484 10284 17536
rect 10324 17484 10376 17536
rect 11152 17484 11204 17536
rect 12624 17688 12676 17740
rect 13268 17731 13320 17740
rect 13268 17697 13277 17731
rect 13277 17697 13311 17731
rect 13311 17697 13320 17731
rect 13268 17688 13320 17697
rect 14004 17756 14056 17808
rect 13452 17688 13504 17740
rect 13728 17731 13780 17740
rect 13728 17697 13737 17731
rect 13737 17697 13771 17731
rect 13771 17697 13780 17731
rect 13728 17688 13780 17697
rect 13820 17688 13872 17740
rect 14372 17824 14424 17876
rect 15108 17824 15160 17876
rect 15292 17824 15344 17876
rect 13636 17620 13688 17672
rect 15200 17688 15252 17740
rect 17684 17824 17736 17876
rect 18144 17824 18196 17876
rect 23204 17824 23256 17876
rect 18052 17756 18104 17808
rect 16856 17731 16908 17740
rect 16856 17697 16865 17731
rect 16865 17697 16899 17731
rect 16899 17697 16908 17731
rect 16856 17688 16908 17697
rect 13912 17527 13964 17536
rect 13912 17493 13921 17527
rect 13921 17493 13955 17527
rect 13955 17493 13964 17527
rect 13912 17484 13964 17493
rect 14740 17484 14792 17536
rect 16580 17620 16632 17672
rect 17592 17688 17644 17740
rect 17776 17731 17828 17740
rect 17776 17697 17785 17731
rect 17785 17697 17819 17731
rect 17819 17697 17828 17731
rect 17776 17688 17828 17697
rect 20076 17756 20128 17808
rect 23572 17756 23624 17808
rect 24308 17756 24360 17808
rect 15292 17552 15344 17604
rect 18696 17731 18748 17740
rect 18696 17697 18705 17731
rect 18705 17697 18739 17731
rect 18739 17697 18748 17731
rect 18696 17688 18748 17697
rect 19064 17731 19116 17740
rect 19064 17697 19073 17731
rect 19073 17697 19107 17731
rect 19107 17697 19116 17731
rect 19064 17688 19116 17697
rect 17960 17620 18012 17672
rect 18328 17620 18380 17672
rect 20444 17688 20496 17740
rect 20904 17688 20956 17740
rect 18052 17552 18104 17604
rect 19892 17552 19944 17604
rect 21824 17620 21876 17672
rect 22468 17731 22520 17740
rect 22468 17697 22477 17731
rect 22477 17697 22511 17731
rect 22511 17697 22520 17731
rect 22468 17688 22520 17697
rect 22744 17731 22796 17740
rect 22744 17697 22753 17731
rect 22753 17697 22787 17731
rect 22787 17697 22796 17731
rect 22744 17688 22796 17697
rect 24676 17688 24728 17740
rect 24860 17756 24912 17808
rect 24492 17620 24544 17672
rect 25044 17756 25096 17808
rect 25228 17799 25280 17808
rect 25228 17765 25237 17799
rect 25237 17765 25271 17799
rect 25271 17765 25280 17799
rect 25228 17756 25280 17765
rect 25964 17824 26016 17876
rect 20260 17552 20312 17604
rect 15936 17527 15988 17536
rect 15936 17493 15945 17527
rect 15945 17493 15979 17527
rect 15979 17493 15988 17527
rect 15936 17484 15988 17493
rect 16304 17484 16356 17536
rect 18420 17484 18472 17536
rect 19248 17527 19300 17536
rect 19248 17493 19257 17527
rect 19257 17493 19291 17527
rect 19291 17493 19300 17527
rect 19248 17484 19300 17493
rect 19616 17527 19668 17536
rect 19616 17493 19625 17527
rect 19625 17493 19659 17527
rect 19659 17493 19668 17527
rect 19616 17484 19668 17493
rect 21640 17527 21692 17536
rect 21640 17493 21649 17527
rect 21649 17493 21683 17527
rect 21683 17493 21692 17527
rect 21640 17484 21692 17493
rect 22560 17484 22612 17536
rect 23296 17484 23348 17536
rect 23756 17484 23808 17536
rect 24860 17552 24912 17604
rect 24400 17527 24452 17536
rect 24400 17493 24409 17527
rect 24409 17493 24443 17527
rect 24443 17493 24452 17527
rect 24400 17484 24452 17493
rect 25136 17484 25188 17536
rect 3756 17382 3808 17434
rect 3820 17382 3872 17434
rect 3884 17382 3936 17434
rect 3948 17382 4000 17434
rect 4012 17382 4064 17434
rect 10472 17382 10524 17434
rect 10536 17382 10588 17434
rect 10600 17382 10652 17434
rect 10664 17382 10716 17434
rect 10728 17382 10780 17434
rect 17188 17382 17240 17434
rect 17252 17382 17304 17434
rect 17316 17382 17368 17434
rect 17380 17382 17432 17434
rect 17444 17382 17496 17434
rect 23904 17382 23956 17434
rect 23968 17382 24020 17434
rect 24032 17382 24084 17434
rect 24096 17382 24148 17434
rect 24160 17382 24212 17434
rect 1400 17323 1452 17332
rect 1400 17289 1409 17323
rect 1409 17289 1443 17323
rect 1443 17289 1452 17323
rect 1400 17280 1452 17289
rect 1768 17280 1820 17332
rect 2780 17323 2832 17332
rect 2780 17289 2789 17323
rect 2789 17289 2823 17323
rect 2823 17289 2832 17323
rect 2780 17280 2832 17289
rect 4160 17280 4212 17332
rect 4252 17280 4304 17332
rect 4620 17280 4672 17332
rect 6644 17280 6696 17332
rect 2964 17212 3016 17264
rect 1952 17144 2004 17196
rect 2504 17144 2556 17196
rect 1676 17076 1728 17128
rect 3516 17076 3568 17128
rect 3332 17008 3384 17060
rect 9036 17280 9088 17332
rect 9128 17280 9180 17332
rect 9680 17280 9732 17332
rect 10600 17280 10652 17332
rect 10968 17280 11020 17332
rect 6276 17144 6328 17196
rect 7932 17144 7984 17196
rect 6092 17119 6144 17128
rect 6092 17085 6101 17119
rect 6101 17085 6135 17119
rect 6135 17085 6144 17119
rect 6092 17076 6144 17085
rect 7012 17119 7064 17128
rect 7012 17085 7021 17119
rect 7021 17085 7055 17119
rect 7055 17085 7064 17119
rect 7012 17076 7064 17085
rect 4896 17051 4948 17060
rect 4896 17017 4930 17051
rect 4930 17017 4948 17051
rect 4896 17008 4948 17017
rect 6920 17008 6972 17060
rect 8024 17076 8076 17128
rect 14188 17280 14240 17332
rect 15016 17280 15068 17332
rect 16304 17280 16356 17332
rect 10232 17187 10284 17196
rect 10232 17153 10241 17187
rect 10241 17153 10275 17187
rect 10275 17153 10284 17187
rect 10232 17144 10284 17153
rect 10324 17187 10376 17196
rect 10324 17153 10333 17187
rect 10333 17153 10367 17187
rect 10367 17153 10376 17187
rect 10324 17144 10376 17153
rect 9956 17076 10008 17128
rect 10048 17119 10100 17128
rect 10048 17085 10057 17119
rect 10057 17085 10091 17119
rect 10091 17085 10100 17119
rect 10048 17076 10100 17085
rect 10416 17119 10468 17128
rect 10416 17085 10421 17119
rect 10421 17085 10455 17119
rect 10455 17085 10468 17119
rect 10416 17076 10468 17085
rect 10508 17076 10560 17128
rect 10968 17076 11020 17128
rect 11152 17119 11204 17128
rect 11152 17085 11161 17119
rect 11161 17085 11195 17119
rect 11195 17085 11204 17119
rect 16488 17212 16540 17264
rect 17776 17280 17828 17332
rect 13912 17144 13964 17196
rect 14004 17144 14056 17196
rect 15016 17144 15068 17196
rect 17960 17212 18012 17264
rect 18052 17187 18104 17196
rect 11152 17076 11204 17085
rect 7564 17008 7616 17060
rect 2412 16940 2464 16992
rect 2504 16940 2556 16992
rect 3240 16983 3292 16992
rect 3240 16949 3249 16983
rect 3249 16949 3283 16983
rect 3283 16949 3292 16983
rect 3240 16940 3292 16949
rect 8024 16983 8076 16992
rect 8024 16949 8033 16983
rect 8033 16949 8067 16983
rect 8067 16949 8076 16983
rect 8024 16940 8076 16949
rect 8300 17008 8352 17060
rect 9036 17008 9088 17060
rect 12440 17008 12492 17060
rect 14280 17076 14332 17128
rect 16672 17076 16724 17128
rect 16764 17119 16816 17128
rect 16764 17085 16773 17119
rect 16773 17085 16807 17119
rect 16807 17085 16816 17119
rect 16764 17076 16816 17085
rect 18052 17153 18061 17187
rect 18061 17153 18095 17187
rect 18095 17153 18104 17187
rect 18052 17144 18104 17153
rect 16948 17076 17000 17128
rect 17132 17119 17184 17128
rect 17132 17085 17141 17119
rect 17141 17085 17175 17119
rect 17175 17085 17184 17119
rect 20260 17323 20312 17332
rect 20260 17289 20269 17323
rect 20269 17289 20303 17323
rect 20303 17289 20312 17323
rect 20260 17280 20312 17289
rect 21824 17323 21876 17332
rect 21824 17289 21833 17323
rect 21833 17289 21867 17323
rect 21867 17289 21876 17323
rect 21824 17280 21876 17289
rect 24400 17280 24452 17332
rect 17132 17076 17184 17085
rect 18880 17119 18932 17128
rect 18880 17085 18889 17119
rect 18889 17085 18923 17119
rect 18923 17085 18932 17119
rect 18880 17076 18932 17085
rect 19432 17076 19484 17128
rect 22468 17212 22520 17264
rect 22744 17212 22796 17264
rect 23940 17255 23992 17264
rect 23940 17221 23949 17255
rect 23949 17221 23983 17255
rect 23983 17221 23992 17255
rect 23940 17212 23992 17221
rect 13544 17051 13596 17060
rect 13544 17017 13553 17051
rect 13553 17017 13587 17051
rect 13587 17017 13596 17051
rect 13544 17008 13596 17017
rect 13820 17008 13872 17060
rect 14740 17008 14792 17060
rect 16120 17051 16172 17060
rect 16120 17017 16129 17051
rect 16129 17017 16163 17051
rect 16163 17017 16172 17051
rect 16120 17008 16172 17017
rect 18972 17008 19024 17060
rect 19248 17008 19300 17060
rect 20352 17008 20404 17060
rect 10140 16940 10192 16992
rect 11888 16983 11940 16992
rect 11888 16949 11897 16983
rect 11897 16949 11931 16983
rect 11931 16949 11940 16983
rect 11888 16940 11940 16949
rect 14832 16983 14884 16992
rect 14832 16949 14841 16983
rect 14841 16949 14875 16983
rect 14875 16949 14884 16983
rect 14832 16940 14884 16949
rect 16304 16983 16356 16992
rect 16304 16949 16313 16983
rect 16313 16949 16347 16983
rect 16347 16949 16356 16983
rect 16304 16940 16356 16949
rect 16948 16983 17000 16992
rect 16948 16949 16957 16983
rect 16957 16949 16991 16983
rect 16991 16949 17000 16983
rect 16948 16940 17000 16949
rect 17868 16983 17920 16992
rect 17868 16949 17877 16983
rect 17877 16949 17911 16983
rect 17911 16949 17920 16983
rect 17868 16940 17920 16949
rect 21364 16940 21416 16992
rect 22376 16983 22428 16992
rect 22376 16949 22385 16983
rect 22385 16949 22419 16983
rect 22419 16949 22428 16983
rect 22376 16940 22428 16949
rect 22836 17076 22888 17128
rect 23204 17076 23256 17128
rect 23296 17119 23348 17128
rect 23296 17085 23305 17119
rect 23305 17085 23339 17119
rect 23339 17085 23348 17119
rect 23296 17076 23348 17085
rect 24860 17144 24912 17196
rect 25044 17076 25096 17128
rect 25320 17076 25372 17128
rect 25504 17187 25556 17196
rect 25504 17153 25513 17187
rect 25513 17153 25547 17187
rect 25547 17153 25556 17187
rect 25504 17144 25556 17153
rect 24952 17051 25004 17060
rect 24952 17017 24961 17051
rect 24961 17017 24995 17051
rect 24995 17017 25004 17051
rect 24952 17008 25004 17017
rect 23020 16940 23072 16992
rect 23112 16983 23164 16992
rect 23112 16949 23121 16983
rect 23121 16949 23155 16983
rect 23155 16949 23164 16983
rect 23112 16940 23164 16949
rect 24124 16983 24176 16992
rect 24124 16949 24133 16983
rect 24133 16949 24167 16983
rect 24167 16949 24176 16983
rect 24124 16940 24176 16949
rect 24216 16940 24268 16992
rect 24400 16983 24452 16992
rect 24400 16949 24409 16983
rect 24409 16949 24443 16983
rect 24443 16949 24452 16983
rect 24400 16940 24452 16949
rect 25044 16940 25096 16992
rect 25228 16983 25280 16992
rect 25228 16949 25237 16983
rect 25237 16949 25271 16983
rect 25271 16949 25280 16983
rect 25228 16940 25280 16949
rect 25780 17051 25832 17060
rect 25780 17017 25814 17051
rect 25814 17017 25832 17051
rect 25780 17008 25832 17017
rect 7114 16838 7166 16890
rect 7178 16838 7230 16890
rect 7242 16838 7294 16890
rect 7306 16838 7358 16890
rect 7370 16838 7422 16890
rect 13830 16838 13882 16890
rect 13894 16838 13946 16890
rect 13958 16838 14010 16890
rect 14022 16838 14074 16890
rect 14086 16838 14138 16890
rect 20546 16838 20598 16890
rect 20610 16838 20662 16890
rect 20674 16838 20726 16890
rect 20738 16838 20790 16890
rect 20802 16838 20854 16890
rect 27262 16838 27314 16890
rect 27326 16838 27378 16890
rect 27390 16838 27442 16890
rect 27454 16838 27506 16890
rect 27518 16838 27570 16890
rect 2412 16779 2464 16788
rect 2412 16745 2421 16779
rect 2421 16745 2455 16779
rect 2455 16745 2464 16779
rect 2412 16736 2464 16745
rect 3332 16736 3384 16788
rect 4436 16736 4488 16788
rect 1032 16643 1084 16652
rect 1032 16609 1041 16643
rect 1041 16609 1075 16643
rect 1075 16609 1084 16643
rect 1032 16600 1084 16609
rect 2688 16643 2740 16652
rect 2688 16609 2697 16643
rect 2697 16609 2731 16643
rect 2731 16609 2740 16643
rect 2688 16600 2740 16609
rect 2872 16600 2924 16652
rect 3240 16600 3292 16652
rect 7840 16736 7892 16788
rect 8024 16736 8076 16788
rect 8484 16736 8536 16788
rect 6828 16643 6880 16652
rect 6828 16609 6837 16643
rect 6837 16609 6871 16643
rect 6871 16609 6880 16643
rect 6828 16600 6880 16609
rect 6920 16600 6972 16652
rect 7012 16643 7064 16652
rect 7012 16609 7021 16643
rect 7021 16609 7055 16643
rect 7055 16609 7064 16643
rect 7012 16600 7064 16609
rect 7564 16600 7616 16652
rect 9036 16779 9088 16788
rect 9036 16745 9045 16779
rect 9045 16745 9079 16779
rect 9079 16745 9088 16779
rect 9036 16736 9088 16745
rect 10232 16736 10284 16788
rect 10324 16736 10376 16788
rect 10876 16736 10928 16788
rect 10968 16779 11020 16788
rect 10968 16745 10977 16779
rect 10977 16745 11011 16779
rect 11011 16745 11020 16779
rect 10968 16736 11020 16745
rect 13084 16736 13136 16788
rect 15108 16736 15160 16788
rect 8208 16600 8260 16652
rect 8392 16600 8444 16652
rect 8576 16600 8628 16652
rect 10048 16600 10100 16652
rect 2964 16464 3016 16516
rect 4436 16396 4488 16448
rect 6552 16532 6604 16584
rect 6644 16532 6696 16584
rect 9036 16532 9088 16584
rect 10324 16643 10376 16652
rect 10324 16609 10333 16643
rect 10333 16609 10367 16643
rect 10367 16609 10376 16643
rect 10324 16600 10376 16609
rect 11060 16600 11112 16652
rect 12440 16600 12492 16652
rect 12624 16600 12676 16652
rect 14096 16643 14148 16652
rect 14096 16609 14130 16643
rect 14130 16609 14148 16643
rect 14096 16600 14148 16609
rect 6460 16396 6512 16448
rect 10600 16464 10652 16516
rect 15936 16736 15988 16788
rect 16488 16736 16540 16788
rect 15384 16600 15436 16652
rect 17684 16736 17736 16788
rect 17868 16736 17920 16788
rect 18880 16736 18932 16788
rect 18972 16736 19024 16788
rect 19064 16779 19116 16788
rect 19064 16745 19073 16779
rect 19073 16745 19107 16779
rect 19107 16745 19116 16779
rect 19064 16736 19116 16745
rect 19616 16736 19668 16788
rect 20352 16736 20404 16788
rect 16856 16600 16908 16652
rect 17132 16600 17184 16652
rect 17592 16600 17644 16652
rect 17684 16600 17736 16652
rect 19432 16600 19484 16652
rect 21640 16779 21692 16788
rect 21640 16745 21649 16779
rect 21649 16745 21683 16779
rect 21683 16745 21692 16779
rect 21640 16736 21692 16745
rect 22008 16736 22060 16788
rect 22100 16736 22152 16788
rect 22376 16736 22428 16788
rect 22560 16736 22612 16788
rect 23020 16736 23072 16788
rect 21364 16600 21416 16652
rect 19708 16575 19760 16584
rect 19708 16541 19717 16575
rect 19717 16541 19751 16575
rect 19751 16541 19760 16575
rect 19708 16532 19760 16541
rect 23020 16643 23072 16652
rect 23020 16609 23029 16643
rect 23029 16609 23063 16643
rect 23063 16609 23072 16643
rect 23020 16600 23072 16609
rect 23756 16668 23808 16720
rect 24308 16736 24360 16788
rect 24768 16736 24820 16788
rect 24952 16736 25004 16788
rect 25136 16736 25188 16788
rect 24124 16600 24176 16652
rect 24952 16600 25004 16652
rect 25044 16600 25096 16652
rect 25780 16779 25832 16788
rect 25780 16745 25789 16779
rect 25789 16745 25823 16779
rect 25823 16745 25832 16779
rect 25780 16736 25832 16745
rect 26240 16668 26292 16720
rect 24308 16575 24360 16584
rect 7564 16396 7616 16448
rect 8300 16396 8352 16448
rect 10876 16396 10928 16448
rect 11244 16396 11296 16448
rect 13728 16396 13780 16448
rect 15292 16439 15344 16448
rect 15292 16405 15301 16439
rect 15301 16405 15335 16439
rect 15335 16405 15344 16439
rect 15292 16396 15344 16405
rect 22376 16396 22428 16448
rect 23020 16464 23072 16516
rect 24308 16541 24317 16575
rect 24317 16541 24351 16575
rect 24351 16541 24360 16575
rect 24308 16532 24360 16541
rect 24584 16532 24636 16584
rect 23112 16439 23164 16448
rect 23112 16405 23121 16439
rect 23121 16405 23155 16439
rect 23155 16405 23164 16439
rect 23112 16396 23164 16405
rect 23296 16396 23348 16448
rect 23388 16439 23440 16448
rect 23388 16405 23397 16439
rect 23397 16405 23431 16439
rect 23431 16405 23440 16439
rect 23388 16396 23440 16405
rect 25228 16396 25280 16448
rect 3756 16294 3808 16346
rect 3820 16294 3872 16346
rect 3884 16294 3936 16346
rect 3948 16294 4000 16346
rect 4012 16294 4064 16346
rect 10472 16294 10524 16346
rect 10536 16294 10588 16346
rect 10600 16294 10652 16346
rect 10664 16294 10716 16346
rect 10728 16294 10780 16346
rect 17188 16294 17240 16346
rect 17252 16294 17304 16346
rect 17316 16294 17368 16346
rect 17380 16294 17432 16346
rect 17444 16294 17496 16346
rect 23904 16294 23956 16346
rect 23968 16294 24020 16346
rect 24032 16294 24084 16346
rect 24096 16294 24148 16346
rect 24160 16294 24212 16346
rect 2688 16235 2740 16244
rect 2688 16201 2697 16235
rect 2697 16201 2731 16235
rect 2731 16201 2740 16235
rect 2688 16192 2740 16201
rect 6184 16192 6236 16244
rect 8852 16235 8904 16244
rect 8852 16201 8861 16235
rect 8861 16201 8895 16235
rect 8895 16201 8904 16235
rect 8852 16192 8904 16201
rect 9404 16192 9456 16244
rect 11060 16235 11112 16244
rect 11060 16201 11069 16235
rect 11069 16201 11103 16235
rect 11103 16201 11112 16235
rect 11060 16192 11112 16201
rect 11152 16192 11204 16244
rect 11428 16192 11480 16244
rect 14096 16192 14148 16244
rect 2596 16056 2648 16108
rect 11336 16124 11388 16176
rect 12900 16124 12952 16176
rect 2136 16031 2188 16040
rect 2136 15997 2145 16031
rect 2145 15997 2179 16031
rect 2179 15997 2188 16031
rect 2136 15988 2188 15997
rect 1676 15920 1728 15972
rect 1768 15895 1820 15904
rect 1768 15861 1777 15895
rect 1777 15861 1811 15895
rect 1811 15861 1820 15895
rect 1768 15852 1820 15861
rect 1952 15920 2004 15972
rect 2412 16031 2464 16040
rect 2412 15997 2421 16031
rect 2421 15997 2455 16031
rect 2455 15997 2464 16031
rect 2412 15988 2464 15997
rect 2320 15920 2372 15972
rect 2872 16031 2924 16040
rect 2872 15997 2881 16031
rect 2881 15997 2915 16031
rect 2915 15997 2924 16031
rect 2872 15988 2924 15997
rect 2964 16031 3016 16040
rect 2964 15997 2973 16031
rect 2973 15997 3007 16031
rect 3007 15997 3016 16031
rect 2964 15988 3016 15997
rect 8208 16056 8260 16108
rect 9036 16056 9088 16108
rect 4436 15988 4488 16040
rect 6092 15988 6144 16040
rect 3332 15920 3384 15972
rect 6552 15920 6604 15972
rect 6460 15852 6512 15904
rect 7472 15895 7524 15904
rect 7472 15861 7481 15895
rect 7481 15861 7515 15895
rect 7515 15861 7524 15895
rect 7472 15852 7524 15861
rect 7656 15920 7708 15972
rect 9956 15920 10008 15972
rect 10692 15963 10744 15972
rect 10692 15929 10701 15963
rect 10701 15929 10735 15963
rect 10735 15929 10744 15963
rect 10692 15920 10744 15929
rect 11060 15920 11112 15972
rect 11244 16031 11296 16040
rect 11244 15997 11253 16031
rect 11253 15997 11287 16031
rect 11287 15997 11296 16031
rect 11244 15988 11296 15997
rect 11336 16031 11388 16040
rect 11336 15997 11345 16031
rect 11345 15997 11379 16031
rect 11379 15997 11388 16031
rect 11336 15988 11388 15997
rect 11888 15988 11940 16040
rect 13452 15988 13504 16040
rect 11704 15852 11756 15904
rect 14924 16056 14976 16108
rect 15568 16192 15620 16244
rect 16488 16192 16540 16244
rect 19708 16192 19760 16244
rect 19984 16235 20036 16244
rect 19984 16201 19993 16235
rect 19993 16201 20027 16235
rect 20027 16201 20036 16235
rect 19984 16192 20036 16201
rect 25320 16192 25372 16244
rect 15752 16099 15804 16108
rect 15752 16065 15761 16099
rect 15761 16065 15795 16099
rect 15795 16065 15804 16099
rect 15752 16056 15804 16065
rect 15292 15988 15344 16040
rect 15476 15988 15528 16040
rect 16212 15988 16264 16040
rect 17776 15988 17828 16040
rect 18328 16031 18380 16040
rect 18328 15997 18337 16031
rect 18337 15997 18371 16031
rect 18371 15997 18380 16031
rect 18328 15988 18380 15997
rect 18420 16031 18472 16040
rect 18420 15997 18429 16031
rect 18429 15997 18463 16031
rect 18463 15997 18472 16031
rect 18420 15988 18472 15997
rect 20444 15988 20496 16040
rect 14832 15920 14884 15972
rect 18788 15920 18840 15972
rect 21088 16031 21140 16040
rect 21088 15997 21097 16031
rect 21097 15997 21131 16031
rect 21131 15997 21140 16031
rect 21088 15988 21140 15997
rect 22652 15988 22704 16040
rect 23756 15988 23808 16040
rect 24124 16031 24176 16040
rect 24124 15997 24133 16031
rect 24133 15997 24167 16031
rect 24167 15997 24176 16031
rect 24124 15988 24176 15997
rect 24768 15988 24820 16040
rect 26240 15988 26292 16040
rect 26884 15988 26936 16040
rect 15476 15895 15528 15904
rect 15476 15861 15485 15895
rect 15485 15861 15519 15895
rect 15519 15861 15528 15895
rect 15476 15852 15528 15861
rect 17684 15895 17736 15904
rect 17684 15861 17693 15895
rect 17693 15861 17727 15895
rect 17727 15861 17736 15895
rect 17684 15852 17736 15861
rect 17960 15852 18012 15904
rect 20904 15895 20956 15904
rect 20904 15861 20913 15895
rect 20913 15861 20947 15895
rect 20947 15861 20956 15895
rect 20904 15852 20956 15861
rect 21456 15852 21508 15904
rect 23572 15852 23624 15904
rect 24676 15852 24728 15904
rect 7114 15750 7166 15802
rect 7178 15750 7230 15802
rect 7242 15750 7294 15802
rect 7306 15750 7358 15802
rect 7370 15750 7422 15802
rect 13830 15750 13882 15802
rect 13894 15750 13946 15802
rect 13958 15750 14010 15802
rect 14022 15750 14074 15802
rect 14086 15750 14138 15802
rect 20546 15750 20598 15802
rect 20610 15750 20662 15802
rect 20674 15750 20726 15802
rect 20738 15750 20790 15802
rect 20802 15750 20854 15802
rect 27262 15750 27314 15802
rect 27326 15750 27378 15802
rect 27390 15750 27442 15802
rect 27454 15750 27506 15802
rect 27518 15750 27570 15802
rect 1676 15648 1728 15700
rect 1768 15648 1820 15700
rect 2596 15648 2648 15700
rect 6828 15648 6880 15700
rect 7472 15648 7524 15700
rect 7564 15648 7616 15700
rect 940 15512 992 15564
rect 2412 15512 2464 15564
rect 3148 15487 3200 15496
rect 3148 15453 3157 15487
rect 3157 15453 3191 15487
rect 3191 15453 3200 15487
rect 3148 15444 3200 15453
rect 4436 15580 4488 15632
rect 8484 15648 8536 15700
rect 9036 15691 9088 15700
rect 9036 15657 9045 15691
rect 9045 15657 9079 15691
rect 9079 15657 9088 15691
rect 9036 15648 9088 15657
rect 3516 15555 3568 15564
rect 3516 15521 3550 15555
rect 3550 15521 3568 15555
rect 3516 15512 3568 15521
rect 4252 15512 4304 15564
rect 6092 15512 6144 15564
rect 6184 15512 6236 15564
rect 8024 15623 8076 15632
rect 8024 15589 8049 15623
rect 8049 15589 8076 15623
rect 8024 15580 8076 15589
rect 10876 15648 10928 15700
rect 15660 15648 15712 15700
rect 15936 15648 15988 15700
rect 16212 15648 16264 15700
rect 17684 15648 17736 15700
rect 18328 15648 18380 15700
rect 6644 15512 6696 15564
rect 6736 15512 6788 15564
rect 2136 15376 2188 15428
rect 1124 15308 1176 15360
rect 1584 15308 1636 15360
rect 2320 15308 2372 15360
rect 2412 15351 2464 15360
rect 2412 15317 2421 15351
rect 2421 15317 2455 15351
rect 2455 15317 2464 15351
rect 2412 15308 2464 15317
rect 2780 15308 2832 15360
rect 4160 15308 4212 15360
rect 5724 15376 5776 15428
rect 7472 15487 7524 15496
rect 7472 15453 7481 15487
rect 7481 15453 7515 15487
rect 7515 15453 7524 15487
rect 7472 15444 7524 15453
rect 8392 15444 8444 15496
rect 4712 15351 4764 15360
rect 4712 15317 4721 15351
rect 4721 15317 4755 15351
rect 4755 15317 4764 15351
rect 4712 15308 4764 15317
rect 5540 15351 5592 15360
rect 5540 15317 5549 15351
rect 5549 15317 5583 15351
rect 5583 15317 5592 15351
rect 5540 15308 5592 15317
rect 8668 15308 8720 15360
rect 10324 15512 10376 15564
rect 13544 15580 13596 15632
rect 11244 15555 11296 15564
rect 11244 15521 11278 15555
rect 11278 15521 11296 15555
rect 11244 15512 11296 15521
rect 12440 15555 12492 15564
rect 12440 15521 12449 15555
rect 12449 15521 12483 15555
rect 12483 15521 12492 15555
rect 12440 15512 12492 15521
rect 12716 15555 12768 15564
rect 12716 15521 12750 15555
rect 12750 15521 12768 15555
rect 12716 15512 12768 15521
rect 12992 15512 13044 15564
rect 14280 15555 14332 15564
rect 14280 15521 14289 15555
rect 14289 15521 14323 15555
rect 14323 15521 14332 15555
rect 14280 15512 14332 15521
rect 13820 15444 13872 15496
rect 15476 15580 15528 15632
rect 18788 15580 18840 15632
rect 21272 15648 21324 15700
rect 15200 15555 15252 15564
rect 15200 15521 15209 15555
rect 15209 15521 15243 15555
rect 15243 15521 15252 15555
rect 15200 15512 15252 15521
rect 15568 15444 15620 15496
rect 19616 15512 19668 15564
rect 23296 15648 23348 15700
rect 20996 15512 21048 15564
rect 17592 15487 17644 15496
rect 17592 15453 17601 15487
rect 17601 15453 17635 15487
rect 17635 15453 17644 15487
rect 17592 15444 17644 15453
rect 19432 15487 19484 15496
rect 19432 15453 19441 15487
rect 19441 15453 19475 15487
rect 19475 15453 19484 15487
rect 19432 15444 19484 15453
rect 20260 15487 20312 15496
rect 20260 15453 20269 15487
rect 20269 15453 20303 15487
rect 20303 15453 20312 15487
rect 20260 15444 20312 15453
rect 12348 15351 12400 15360
rect 12348 15317 12357 15351
rect 12357 15317 12391 15351
rect 12391 15317 12400 15351
rect 12348 15308 12400 15317
rect 19340 15419 19392 15428
rect 19340 15385 19349 15419
rect 19349 15385 19383 15419
rect 19383 15385 19392 15419
rect 19340 15376 19392 15385
rect 22652 15512 22704 15564
rect 23480 15512 23532 15564
rect 23756 15512 23808 15564
rect 24124 15580 24176 15632
rect 24308 15580 24360 15632
rect 24584 15623 24636 15632
rect 24584 15589 24593 15623
rect 24593 15589 24627 15623
rect 24627 15589 24636 15623
rect 24584 15580 24636 15589
rect 22928 15444 22980 15496
rect 23296 15487 23348 15496
rect 22284 15376 22336 15428
rect 13452 15308 13504 15360
rect 13912 15351 13964 15360
rect 13912 15317 13921 15351
rect 13921 15317 13955 15351
rect 13955 15317 13964 15351
rect 13912 15308 13964 15317
rect 14832 15351 14884 15360
rect 14832 15317 14841 15351
rect 14841 15317 14875 15351
rect 14875 15317 14884 15351
rect 14832 15308 14884 15317
rect 21916 15351 21968 15360
rect 21916 15317 21925 15351
rect 21925 15317 21959 15351
rect 21959 15317 21968 15351
rect 21916 15308 21968 15317
rect 23296 15453 23305 15487
rect 23305 15453 23339 15487
rect 23339 15453 23348 15487
rect 23296 15444 23348 15453
rect 23572 15308 23624 15360
rect 24492 15512 24544 15564
rect 25412 15555 25464 15564
rect 25412 15521 25421 15555
rect 25421 15521 25455 15555
rect 25455 15521 25464 15555
rect 25412 15512 25464 15521
rect 24768 15351 24820 15360
rect 24768 15317 24777 15351
rect 24777 15317 24811 15351
rect 24811 15317 24820 15351
rect 24768 15308 24820 15317
rect 26240 15308 26292 15360
rect 3756 15206 3808 15258
rect 3820 15206 3872 15258
rect 3884 15206 3936 15258
rect 3948 15206 4000 15258
rect 4012 15206 4064 15258
rect 10472 15206 10524 15258
rect 10536 15206 10588 15258
rect 10600 15206 10652 15258
rect 10664 15206 10716 15258
rect 10728 15206 10780 15258
rect 17188 15206 17240 15258
rect 17252 15206 17304 15258
rect 17316 15206 17368 15258
rect 17380 15206 17432 15258
rect 17444 15206 17496 15258
rect 23904 15206 23956 15258
rect 23968 15206 24020 15258
rect 24032 15206 24084 15258
rect 24096 15206 24148 15258
rect 24160 15206 24212 15258
rect 940 15147 992 15156
rect 940 15113 949 15147
rect 949 15113 983 15147
rect 983 15113 992 15147
rect 940 15104 992 15113
rect 1032 14968 1084 15020
rect 2044 15104 2096 15156
rect 2688 15104 2740 15156
rect 3516 15104 3568 15156
rect 4436 15104 4488 15156
rect 2412 14900 2464 14952
rect 2504 14900 2556 14952
rect 4528 15036 4580 15088
rect 4712 15036 4764 15088
rect 6552 15147 6604 15156
rect 6552 15113 6561 15147
rect 6561 15113 6595 15147
rect 6595 15113 6604 15147
rect 6552 15104 6604 15113
rect 7012 15104 7064 15156
rect 8392 15104 8444 15156
rect 10232 15104 10284 15156
rect 12992 15104 13044 15156
rect 13820 15104 13872 15156
rect 14740 15104 14792 15156
rect 15200 15104 15252 15156
rect 17776 15104 17828 15156
rect 20260 15104 20312 15156
rect 21088 15104 21140 15156
rect 23296 15147 23348 15156
rect 23296 15113 23305 15147
rect 23305 15113 23339 15147
rect 23339 15113 23348 15147
rect 23296 15104 23348 15113
rect 24768 15104 24820 15156
rect 25412 15104 25464 15156
rect 6276 14968 6328 15020
rect 6460 14968 6512 15020
rect 6828 15011 6880 15020
rect 6828 14977 6837 15011
rect 6837 14977 6871 15011
rect 6871 14977 6880 15011
rect 6828 14968 6880 14977
rect 12624 15036 12676 15088
rect 12716 15079 12768 15088
rect 12716 15045 12725 15079
rect 12725 15045 12759 15079
rect 12759 15045 12768 15079
rect 12716 15036 12768 15045
rect 14096 15036 14148 15088
rect 14556 15036 14608 15088
rect 15568 15079 15620 15088
rect 15568 15045 15577 15079
rect 15577 15045 15611 15079
rect 15611 15045 15620 15079
rect 15568 15036 15620 15045
rect 22928 15036 22980 15088
rect 3700 14900 3752 14952
rect 5080 14832 5132 14884
rect 5540 14832 5592 14884
rect 2320 14764 2372 14816
rect 3148 14764 3200 14816
rect 3424 14764 3476 14816
rect 6184 14832 6236 14884
rect 6368 14875 6420 14884
rect 6368 14841 6377 14875
rect 6377 14841 6411 14875
rect 6411 14841 6420 14875
rect 6368 14832 6420 14841
rect 6736 14943 6788 14952
rect 6736 14909 6745 14943
rect 6745 14909 6779 14943
rect 6779 14909 6788 14943
rect 6736 14900 6788 14909
rect 8668 14943 8720 14952
rect 8668 14909 8677 14943
rect 8677 14909 8711 14943
rect 8711 14909 8720 14943
rect 8668 14900 8720 14909
rect 8852 14900 8904 14952
rect 9680 14900 9732 14952
rect 9128 14832 9180 14884
rect 9404 14832 9456 14884
rect 10876 14900 10928 14952
rect 12348 14900 12400 14952
rect 13912 14968 13964 15020
rect 15384 14968 15436 15020
rect 16212 14968 16264 15020
rect 18052 14968 18104 15020
rect 23664 14968 23716 15020
rect 13084 14943 13136 14952
rect 13084 14909 13093 14943
rect 13093 14909 13127 14943
rect 13127 14909 13136 14943
rect 13084 14900 13136 14909
rect 13176 14943 13228 14952
rect 13176 14909 13185 14943
rect 13185 14909 13219 14943
rect 13219 14909 13228 14943
rect 13176 14900 13228 14909
rect 13452 14900 13504 14952
rect 6736 14764 6788 14816
rect 8300 14764 8352 14816
rect 10232 14764 10284 14816
rect 10508 14807 10560 14816
rect 10508 14773 10517 14807
rect 10517 14773 10551 14807
rect 10551 14773 10560 14807
rect 10508 14764 10560 14773
rect 11704 14832 11756 14884
rect 14096 14832 14148 14884
rect 12072 14764 12124 14816
rect 13544 14764 13596 14816
rect 14372 14900 14424 14952
rect 14740 14900 14792 14952
rect 14924 14943 14976 14952
rect 14924 14909 14933 14943
rect 14933 14909 14967 14943
rect 14967 14909 14976 14943
rect 14924 14900 14976 14909
rect 15292 14832 15344 14884
rect 17960 14943 18012 14952
rect 17960 14909 17969 14943
rect 17969 14909 18003 14943
rect 18003 14909 18012 14943
rect 17960 14900 18012 14909
rect 18420 14832 18472 14884
rect 19248 14832 19300 14884
rect 20904 14900 20956 14952
rect 21916 14900 21968 14952
rect 22836 14943 22888 14952
rect 22836 14909 22845 14943
rect 22845 14909 22879 14943
rect 22879 14909 22888 14943
rect 22836 14900 22888 14909
rect 23480 14943 23532 14952
rect 23480 14909 23489 14943
rect 23489 14909 23523 14943
rect 23523 14909 23532 14943
rect 23480 14900 23532 14909
rect 24400 14943 24452 14952
rect 24400 14909 24409 14943
rect 24409 14909 24443 14943
rect 24443 14909 24452 14943
rect 24400 14900 24452 14909
rect 24584 14943 24636 14952
rect 24584 14909 24593 14943
rect 24593 14909 24627 14943
rect 24627 14909 24636 14943
rect 24584 14900 24636 14909
rect 18236 14764 18288 14816
rect 18328 14764 18380 14816
rect 20812 14764 20864 14816
rect 22284 14807 22336 14816
rect 22284 14773 22293 14807
rect 22293 14773 22327 14807
rect 22327 14773 22336 14807
rect 22284 14764 22336 14773
rect 23020 14807 23072 14816
rect 23020 14773 23029 14807
rect 23029 14773 23063 14807
rect 23063 14773 23072 14807
rect 23020 14764 23072 14773
rect 24124 14807 24176 14816
rect 24124 14773 24133 14807
rect 24133 14773 24167 14807
rect 24167 14773 24176 14807
rect 24124 14764 24176 14773
rect 24400 14764 24452 14816
rect 24676 14875 24728 14884
rect 24676 14841 24685 14875
rect 24685 14841 24719 14875
rect 24719 14841 24728 14875
rect 24676 14832 24728 14841
rect 26240 14900 26292 14952
rect 26884 14900 26936 14952
rect 25228 14764 25280 14816
rect 7114 14662 7166 14714
rect 7178 14662 7230 14714
rect 7242 14662 7294 14714
rect 7306 14662 7358 14714
rect 7370 14662 7422 14714
rect 13830 14662 13882 14714
rect 13894 14662 13946 14714
rect 13958 14662 14010 14714
rect 14022 14662 14074 14714
rect 14086 14662 14138 14714
rect 20546 14662 20598 14714
rect 20610 14662 20662 14714
rect 20674 14662 20726 14714
rect 20738 14662 20790 14714
rect 20802 14662 20854 14714
rect 27262 14662 27314 14714
rect 27326 14662 27378 14714
rect 27390 14662 27442 14714
rect 27454 14662 27506 14714
rect 27518 14662 27570 14714
rect 1032 14560 1084 14612
rect 4528 14560 4580 14612
rect 6368 14560 6420 14612
rect 6920 14560 6972 14612
rect 7472 14560 7524 14612
rect 8024 14560 8076 14612
rect 8116 14603 8168 14612
rect 8116 14569 8125 14603
rect 8125 14569 8159 14603
rect 8159 14569 8168 14603
rect 8116 14560 8168 14569
rect 1124 14535 1176 14544
rect 1124 14501 1158 14535
rect 1158 14501 1176 14535
rect 1124 14492 1176 14501
rect 1768 14492 1820 14544
rect 2136 14492 2188 14544
rect 2688 14492 2740 14544
rect 2504 14424 2556 14476
rect 2780 14467 2832 14476
rect 2780 14433 2789 14467
rect 2789 14433 2823 14467
rect 2823 14433 2832 14467
rect 2780 14424 2832 14433
rect 3332 14492 3384 14544
rect 6276 14492 6328 14544
rect 9036 14535 9088 14544
rect 4528 14424 4580 14476
rect 9036 14501 9047 14535
rect 9047 14501 9088 14535
rect 9036 14492 9088 14501
rect 9404 14603 9456 14612
rect 9404 14569 9413 14603
rect 9413 14569 9447 14603
rect 9447 14569 9456 14603
rect 9404 14560 9456 14569
rect 9496 14560 9548 14612
rect 6828 14424 6880 14476
rect 3516 14356 3568 14408
rect 4804 14356 4856 14408
rect 8668 14467 8720 14476
rect 8668 14433 8677 14467
rect 8677 14433 8711 14467
rect 8711 14433 8720 14467
rect 8668 14424 8720 14433
rect 4344 14288 4396 14340
rect 6368 14288 6420 14340
rect 2320 14220 2372 14272
rect 5908 14263 5960 14272
rect 5908 14229 5917 14263
rect 5917 14229 5951 14263
rect 5951 14229 5960 14263
rect 5908 14220 5960 14229
rect 9128 14356 9180 14408
rect 9588 14467 9640 14476
rect 9588 14433 9597 14467
rect 9597 14433 9631 14467
rect 9631 14433 9640 14467
rect 9588 14424 9640 14433
rect 9772 14467 9824 14476
rect 9772 14433 9781 14467
rect 9781 14433 9815 14467
rect 9815 14433 9824 14467
rect 9772 14424 9824 14433
rect 10232 14492 10284 14544
rect 11888 14560 11940 14612
rect 13636 14560 13688 14612
rect 11060 14492 11112 14544
rect 11980 14492 12032 14544
rect 14832 14560 14884 14612
rect 15292 14603 15344 14612
rect 15292 14569 15301 14603
rect 15301 14569 15335 14603
rect 15335 14569 15344 14603
rect 15292 14560 15344 14569
rect 19248 14560 19300 14612
rect 14924 14424 14976 14476
rect 19616 14492 19668 14544
rect 19892 14492 19944 14544
rect 21272 14492 21324 14544
rect 9588 14288 9640 14340
rect 7012 14220 7064 14272
rect 8484 14220 8536 14272
rect 9864 14220 9916 14272
rect 10416 14288 10468 14340
rect 10968 14399 11020 14408
rect 10968 14365 10977 14399
rect 10977 14365 11011 14399
rect 11011 14365 11020 14399
rect 10968 14356 11020 14365
rect 12072 14399 12124 14408
rect 12072 14365 12081 14399
rect 12081 14365 12115 14399
rect 12115 14365 12124 14399
rect 12072 14356 12124 14365
rect 12164 14399 12216 14408
rect 12164 14365 12173 14399
rect 12173 14365 12207 14399
rect 12207 14365 12216 14399
rect 12164 14356 12216 14365
rect 11244 14288 11296 14340
rect 11612 14263 11664 14272
rect 11612 14229 11621 14263
rect 11621 14229 11655 14263
rect 11655 14229 11664 14263
rect 11612 14220 11664 14229
rect 11796 14220 11848 14272
rect 12624 14263 12676 14272
rect 12624 14229 12633 14263
rect 12633 14229 12667 14263
rect 12667 14229 12676 14263
rect 12624 14220 12676 14229
rect 16856 14399 16908 14408
rect 16856 14365 16865 14399
rect 16865 14365 16899 14399
rect 16899 14365 16908 14399
rect 16856 14356 16908 14365
rect 18420 14467 18472 14476
rect 18420 14433 18429 14467
rect 18429 14433 18463 14467
rect 18463 14433 18472 14467
rect 18420 14424 18472 14433
rect 18604 14424 18656 14476
rect 17040 14356 17092 14408
rect 18144 14399 18196 14408
rect 18144 14365 18153 14399
rect 18153 14365 18187 14399
rect 18187 14365 18196 14399
rect 18144 14356 18196 14365
rect 18696 14356 18748 14408
rect 18880 14467 18932 14476
rect 18880 14433 18889 14467
rect 18889 14433 18923 14467
rect 18923 14433 18932 14467
rect 18880 14424 18932 14433
rect 20352 14424 20404 14476
rect 19708 14356 19760 14408
rect 19892 14356 19944 14408
rect 22284 14560 22336 14612
rect 22376 14560 22428 14612
rect 23020 14560 23072 14612
rect 24124 14560 24176 14612
rect 24308 14560 24360 14612
rect 24584 14603 24636 14612
rect 24584 14569 24593 14603
rect 24593 14569 24627 14603
rect 24627 14569 24636 14603
rect 24584 14560 24636 14569
rect 24676 14560 24728 14612
rect 23388 14492 23440 14544
rect 23020 14467 23072 14476
rect 23020 14433 23029 14467
rect 23029 14433 23063 14467
rect 23063 14433 23072 14467
rect 23020 14424 23072 14433
rect 23204 14467 23256 14476
rect 23204 14433 23237 14467
rect 23237 14433 23256 14467
rect 23204 14424 23256 14433
rect 24400 14492 24452 14544
rect 25044 14424 25096 14476
rect 25228 14560 25280 14612
rect 25504 14492 25556 14544
rect 25412 14424 25464 14476
rect 24768 14288 24820 14340
rect 24860 14331 24912 14340
rect 24860 14297 24869 14331
rect 24869 14297 24903 14331
rect 24903 14297 24912 14331
rect 24860 14288 24912 14297
rect 14648 14220 14700 14272
rect 16488 14263 16540 14272
rect 16488 14229 16497 14263
rect 16497 14229 16531 14263
rect 16531 14229 16540 14263
rect 16488 14220 16540 14229
rect 19524 14220 19576 14272
rect 19708 14263 19760 14272
rect 19708 14229 19717 14263
rect 19717 14229 19751 14263
rect 19751 14229 19760 14263
rect 19708 14220 19760 14229
rect 19800 14220 19852 14272
rect 20260 14220 20312 14272
rect 20996 14220 21048 14272
rect 21548 14220 21600 14272
rect 22284 14263 22336 14272
rect 22284 14229 22293 14263
rect 22293 14229 22327 14263
rect 22327 14229 22336 14263
rect 22284 14220 22336 14229
rect 22468 14263 22520 14272
rect 22468 14229 22477 14263
rect 22477 14229 22511 14263
rect 22511 14229 22520 14263
rect 22468 14220 22520 14229
rect 23756 14220 23808 14272
rect 25136 14288 25188 14340
rect 25320 14263 25372 14272
rect 25320 14229 25329 14263
rect 25329 14229 25363 14263
rect 25363 14229 25372 14263
rect 25320 14220 25372 14229
rect 26148 14288 26200 14340
rect 26240 14263 26292 14272
rect 26240 14229 26249 14263
rect 26249 14229 26283 14263
rect 26283 14229 26292 14263
rect 26240 14220 26292 14229
rect 3756 14118 3808 14170
rect 3820 14118 3872 14170
rect 3884 14118 3936 14170
rect 3948 14118 4000 14170
rect 4012 14118 4064 14170
rect 10472 14118 10524 14170
rect 10536 14118 10588 14170
rect 10600 14118 10652 14170
rect 10664 14118 10716 14170
rect 10728 14118 10780 14170
rect 17188 14118 17240 14170
rect 17252 14118 17304 14170
rect 17316 14118 17368 14170
rect 17380 14118 17432 14170
rect 17444 14118 17496 14170
rect 23904 14118 23956 14170
rect 23968 14118 24020 14170
rect 24032 14118 24084 14170
rect 24096 14118 24148 14170
rect 24160 14118 24212 14170
rect 2780 14016 2832 14068
rect 3516 14016 3568 14068
rect 4436 14016 4488 14068
rect 5080 14016 5132 14068
rect 6828 14016 6880 14068
rect 7012 14059 7064 14068
rect 7012 14025 7021 14059
rect 7021 14025 7055 14059
rect 7055 14025 7064 14059
rect 7012 14016 7064 14025
rect 1308 13744 1360 13796
rect 2872 13855 2924 13864
rect 2872 13821 2881 13855
rect 2881 13821 2915 13855
rect 2915 13821 2924 13855
rect 2872 13812 2924 13821
rect 6184 13923 6236 13932
rect 6184 13889 6193 13923
rect 6193 13889 6227 13923
rect 6227 13889 6236 13923
rect 7472 14016 7524 14068
rect 8668 14016 8720 14068
rect 11060 14016 11112 14068
rect 12164 14016 12216 14068
rect 17040 14016 17092 14068
rect 19892 14016 19944 14068
rect 22744 14016 22796 14068
rect 24216 14016 24268 14068
rect 6184 13880 6236 13889
rect 4068 13812 4120 13864
rect 4344 13855 4396 13864
rect 4344 13821 4362 13855
rect 4362 13821 4396 13855
rect 4344 13812 4396 13821
rect 5908 13855 5960 13864
rect 5908 13821 5926 13855
rect 5926 13821 5960 13855
rect 5908 13812 5960 13821
rect 6092 13812 6144 13864
rect 7656 13880 7708 13932
rect 1124 13676 1176 13728
rect 3332 13744 3384 13796
rect 2136 13719 2188 13728
rect 2136 13685 2145 13719
rect 2145 13685 2179 13719
rect 2179 13685 2188 13719
rect 2136 13676 2188 13685
rect 2228 13719 2280 13728
rect 2228 13685 2237 13719
rect 2237 13685 2271 13719
rect 2271 13685 2280 13719
rect 2228 13676 2280 13685
rect 3056 13676 3108 13728
rect 4804 13719 4856 13728
rect 4804 13685 4813 13719
rect 4813 13685 4847 13719
rect 4847 13685 4856 13719
rect 4804 13676 4856 13685
rect 6276 13787 6328 13796
rect 6276 13753 6285 13787
rect 6285 13753 6319 13787
rect 6319 13753 6328 13787
rect 6276 13744 6328 13753
rect 6368 13744 6420 13796
rect 8852 13812 8904 13864
rect 13084 13923 13136 13932
rect 13084 13889 13093 13923
rect 13093 13889 13127 13923
rect 13127 13889 13136 13923
rect 13084 13880 13136 13889
rect 8208 13744 8260 13796
rect 11336 13812 11388 13864
rect 12716 13812 12768 13864
rect 12256 13744 12308 13796
rect 14372 13880 14424 13932
rect 14832 13948 14884 14000
rect 14740 13880 14792 13932
rect 10324 13719 10376 13728
rect 10324 13685 10333 13719
rect 10333 13685 10367 13719
rect 10367 13685 10376 13719
rect 10324 13676 10376 13685
rect 10784 13676 10836 13728
rect 11060 13676 11112 13728
rect 12716 13676 12768 13728
rect 13084 13676 13136 13728
rect 14556 13855 14608 13864
rect 14556 13821 14565 13855
rect 14565 13821 14599 13855
rect 14599 13821 14608 13855
rect 14556 13812 14608 13821
rect 15476 13855 15528 13864
rect 15476 13821 15485 13855
rect 15485 13821 15519 13855
rect 15519 13821 15528 13855
rect 15476 13812 15528 13821
rect 13636 13676 13688 13728
rect 14188 13676 14240 13728
rect 14280 13676 14332 13728
rect 14464 13676 14516 13728
rect 15016 13719 15068 13728
rect 15016 13685 15025 13719
rect 15025 13685 15059 13719
rect 15059 13685 15068 13719
rect 15016 13676 15068 13685
rect 23204 13948 23256 14000
rect 18052 13923 18104 13932
rect 16672 13744 16724 13796
rect 18052 13889 18061 13923
rect 18061 13889 18095 13923
rect 18095 13889 18104 13923
rect 18052 13880 18104 13889
rect 18604 13880 18656 13932
rect 23848 13991 23900 14000
rect 23848 13957 23857 13991
rect 23857 13957 23891 13991
rect 23891 13957 23900 13991
rect 24952 14059 25004 14068
rect 24952 14025 24961 14059
rect 24961 14025 24995 14059
rect 24995 14025 25004 14059
rect 24952 14016 25004 14025
rect 25044 14016 25096 14068
rect 23848 13948 23900 13957
rect 23756 13880 23808 13932
rect 17776 13812 17828 13864
rect 19984 13812 20036 13864
rect 20444 13812 20496 13864
rect 22836 13812 22888 13864
rect 21088 13744 21140 13796
rect 23664 13744 23716 13796
rect 24216 13812 24268 13864
rect 24400 13744 24452 13796
rect 24768 13880 24820 13932
rect 26240 13812 26292 13864
rect 26884 13812 26936 13864
rect 17316 13676 17368 13728
rect 17868 13719 17920 13728
rect 17868 13685 17877 13719
rect 17877 13685 17911 13719
rect 17911 13685 17920 13719
rect 17868 13676 17920 13685
rect 20904 13719 20956 13728
rect 20904 13685 20913 13719
rect 20913 13685 20947 13719
rect 20947 13685 20956 13719
rect 20904 13676 20956 13685
rect 22928 13719 22980 13728
rect 22928 13685 22937 13719
rect 22937 13685 22971 13719
rect 22971 13685 22980 13719
rect 22928 13676 22980 13685
rect 23480 13676 23532 13728
rect 24860 13676 24912 13728
rect 7114 13574 7166 13626
rect 7178 13574 7230 13626
rect 7242 13574 7294 13626
rect 7306 13574 7358 13626
rect 7370 13574 7422 13626
rect 13830 13574 13882 13626
rect 13894 13574 13946 13626
rect 13958 13574 14010 13626
rect 14022 13574 14074 13626
rect 14086 13574 14138 13626
rect 20546 13574 20598 13626
rect 20610 13574 20662 13626
rect 20674 13574 20726 13626
rect 20738 13574 20790 13626
rect 20802 13574 20854 13626
rect 27262 13574 27314 13626
rect 27326 13574 27378 13626
rect 27390 13574 27442 13626
rect 27454 13574 27506 13626
rect 27518 13574 27570 13626
rect 2228 13472 2280 13524
rect 2504 13472 2556 13524
rect 2688 13472 2740 13524
rect 2872 13472 2924 13524
rect 2136 13336 2188 13388
rect 2228 13379 2280 13388
rect 2228 13345 2237 13379
rect 2237 13345 2271 13379
rect 2271 13345 2280 13379
rect 2228 13336 2280 13345
rect 2412 13336 2464 13388
rect 3332 13404 3384 13456
rect 3424 13447 3476 13456
rect 3424 13413 3433 13447
rect 3433 13413 3467 13447
rect 3467 13413 3476 13447
rect 3424 13404 3476 13413
rect 3516 13336 3568 13388
rect 4804 13472 4856 13524
rect 6092 13472 6144 13524
rect 9772 13472 9824 13524
rect 10968 13472 11020 13524
rect 12256 13515 12308 13524
rect 12256 13481 12265 13515
rect 12265 13481 12299 13515
rect 12299 13481 12308 13515
rect 12256 13472 12308 13481
rect 4160 13379 4212 13388
rect 4160 13345 4169 13379
rect 4169 13345 4203 13379
rect 4203 13345 4212 13379
rect 4160 13336 4212 13345
rect 6000 13404 6052 13456
rect 6276 13404 6328 13456
rect 11796 13404 11848 13456
rect 4804 13311 4856 13320
rect 4804 13277 4813 13311
rect 4813 13277 4847 13311
rect 4847 13277 4856 13311
rect 4804 13268 4856 13277
rect 8116 13336 8168 13388
rect 1216 13132 1268 13184
rect 3148 13175 3200 13184
rect 3148 13141 3157 13175
rect 3157 13141 3191 13175
rect 3191 13141 3200 13175
rect 3148 13132 3200 13141
rect 4068 13132 4120 13184
rect 5908 13200 5960 13252
rect 7656 13268 7708 13320
rect 8392 13311 8444 13320
rect 8392 13277 8401 13311
rect 8401 13277 8435 13311
rect 8435 13277 8444 13311
rect 8392 13268 8444 13277
rect 7748 13200 7800 13252
rect 11060 13336 11112 13388
rect 11888 13379 11940 13388
rect 11888 13345 11897 13379
rect 11897 13345 11931 13379
rect 11931 13345 11940 13379
rect 11888 13336 11940 13345
rect 12624 13472 12676 13524
rect 14464 13472 14516 13524
rect 15476 13472 15528 13524
rect 16488 13515 16540 13524
rect 16488 13481 16497 13515
rect 16497 13481 16531 13515
rect 16531 13481 16540 13515
rect 16488 13472 16540 13481
rect 18420 13515 18472 13524
rect 18420 13481 18429 13515
rect 18429 13481 18463 13515
rect 18463 13481 18472 13515
rect 18420 13472 18472 13481
rect 18880 13472 18932 13524
rect 21088 13472 21140 13524
rect 22836 13472 22888 13524
rect 23020 13472 23072 13524
rect 12808 13379 12860 13388
rect 12808 13345 12842 13379
rect 12842 13345 12860 13379
rect 10784 13311 10836 13320
rect 10784 13277 10793 13311
rect 10793 13277 10827 13311
rect 10827 13277 10836 13311
rect 10784 13268 10836 13277
rect 10876 13268 10928 13320
rect 12808 13336 12860 13345
rect 14280 13379 14332 13388
rect 14280 13345 14314 13379
rect 14314 13345 14332 13379
rect 14280 13336 14332 13345
rect 14740 13336 14792 13388
rect 13912 13268 13964 13320
rect 15200 13268 15252 13320
rect 16672 13311 16724 13320
rect 16672 13277 16681 13311
rect 16681 13277 16715 13311
rect 16715 13277 16724 13311
rect 16672 13268 16724 13277
rect 6920 13132 6972 13184
rect 7380 13175 7432 13184
rect 7380 13141 7389 13175
rect 7389 13141 7423 13175
rect 7423 13141 7432 13175
rect 7380 13132 7432 13141
rect 8576 13175 8628 13184
rect 8576 13141 8585 13175
rect 8585 13141 8619 13175
rect 8619 13141 8628 13175
rect 8576 13132 8628 13141
rect 10968 13175 11020 13184
rect 10968 13141 10977 13175
rect 10977 13141 11011 13175
rect 11011 13141 11020 13175
rect 10968 13132 11020 13141
rect 13636 13132 13688 13184
rect 17316 13379 17368 13388
rect 17316 13345 17350 13379
rect 17350 13345 17368 13379
rect 17316 13336 17368 13345
rect 17592 13336 17644 13388
rect 19892 13379 19944 13388
rect 20904 13404 20956 13456
rect 19892 13345 19910 13379
rect 19910 13345 19944 13379
rect 19892 13336 19944 13345
rect 20260 13336 20312 13388
rect 20352 13336 20404 13388
rect 20536 13336 20588 13388
rect 21272 13379 21324 13388
rect 21272 13345 21281 13379
rect 21281 13345 21315 13379
rect 21315 13345 21324 13379
rect 21272 13336 21324 13345
rect 22928 13404 22980 13456
rect 21548 13379 21600 13388
rect 21548 13345 21582 13379
rect 21582 13345 21600 13379
rect 21548 13336 21600 13345
rect 22468 13336 22520 13388
rect 23296 13336 23348 13388
rect 23480 13336 23532 13388
rect 23112 13311 23164 13320
rect 23112 13277 23121 13311
rect 23121 13277 23155 13311
rect 23155 13277 23164 13311
rect 23112 13268 23164 13277
rect 21088 13200 21140 13252
rect 22836 13200 22888 13252
rect 23664 13379 23716 13388
rect 23664 13345 23673 13379
rect 23673 13345 23707 13379
rect 23707 13345 23716 13379
rect 23664 13336 23716 13345
rect 23756 13336 23808 13388
rect 23848 13379 23900 13388
rect 23848 13345 23857 13379
rect 23857 13345 23891 13379
rect 23891 13345 23900 13379
rect 23848 13336 23900 13345
rect 24860 13515 24912 13524
rect 24860 13481 24869 13515
rect 24869 13481 24903 13515
rect 24903 13481 24912 13515
rect 24860 13472 24912 13481
rect 24952 13472 25004 13524
rect 26148 13404 26200 13456
rect 26884 13336 26936 13388
rect 24400 13200 24452 13252
rect 25044 13268 25096 13320
rect 25136 13268 25188 13320
rect 20260 13132 20312 13184
rect 20628 13132 20680 13184
rect 23572 13132 23624 13184
rect 24308 13175 24360 13184
rect 24308 13141 24317 13175
rect 24317 13141 24351 13175
rect 24351 13141 24360 13175
rect 24308 13132 24360 13141
rect 3756 13030 3808 13082
rect 3820 13030 3872 13082
rect 3884 13030 3936 13082
rect 3948 13030 4000 13082
rect 4012 13030 4064 13082
rect 10472 13030 10524 13082
rect 10536 13030 10588 13082
rect 10600 13030 10652 13082
rect 10664 13030 10716 13082
rect 10728 13030 10780 13082
rect 17188 13030 17240 13082
rect 17252 13030 17304 13082
rect 17316 13030 17368 13082
rect 17380 13030 17432 13082
rect 17444 13030 17496 13082
rect 23904 13030 23956 13082
rect 23968 13030 24020 13082
rect 24032 13030 24084 13082
rect 24096 13030 24148 13082
rect 24160 13030 24212 13082
rect 2412 12928 2464 12980
rect 6276 12971 6328 12980
rect 6276 12937 6285 12971
rect 6285 12937 6319 12971
rect 6319 12937 6328 12971
rect 6276 12928 6328 12937
rect 7380 12928 7432 12980
rect 8116 12928 8168 12980
rect 8576 12928 8628 12980
rect 10968 12928 11020 12980
rect 11704 12971 11756 12980
rect 11704 12937 11713 12971
rect 11713 12937 11747 12971
rect 11747 12937 11756 12971
rect 11704 12928 11756 12937
rect 11888 12971 11940 12980
rect 11888 12937 11897 12971
rect 11897 12937 11931 12971
rect 11931 12937 11940 12971
rect 11888 12928 11940 12937
rect 12808 12971 12860 12980
rect 12808 12937 12817 12971
rect 12817 12937 12851 12971
rect 12851 12937 12860 12971
rect 12808 12928 12860 12937
rect 1124 12724 1176 12776
rect 2228 12724 2280 12776
rect 5080 12860 5132 12912
rect 2320 12656 2372 12708
rect 2688 12656 2740 12708
rect 2780 12699 2832 12708
rect 2780 12665 2798 12699
rect 2798 12665 2832 12699
rect 2780 12656 2832 12665
rect 4436 12767 4488 12776
rect 4436 12733 4445 12767
rect 4445 12733 4479 12767
rect 4479 12733 4488 12767
rect 4436 12724 4488 12733
rect 4804 12724 4856 12776
rect 4988 12656 5040 12708
rect 5724 12724 5776 12776
rect 7748 12792 7800 12844
rect 9772 12835 9824 12844
rect 9772 12801 9781 12835
rect 9781 12801 9815 12835
rect 9815 12801 9824 12835
rect 9772 12792 9824 12801
rect 6460 12767 6512 12776
rect 6460 12733 6469 12767
rect 6469 12733 6503 12767
rect 6503 12733 6512 12767
rect 6460 12724 6512 12733
rect 1308 12588 1360 12640
rect 3148 12588 3200 12640
rect 3240 12631 3292 12640
rect 3240 12597 3249 12631
rect 3249 12597 3283 12631
rect 3283 12597 3292 12631
rect 3240 12588 3292 12597
rect 3976 12631 4028 12640
rect 3976 12597 3985 12631
rect 3985 12597 4019 12631
rect 4019 12597 4028 12631
rect 3976 12588 4028 12597
rect 5080 12588 5132 12640
rect 5908 12588 5960 12640
rect 12072 12860 12124 12912
rect 14556 12971 14608 12980
rect 14556 12937 14565 12971
rect 14565 12937 14599 12971
rect 14599 12937 14608 12971
rect 14556 12928 14608 12937
rect 17868 12928 17920 12980
rect 19892 12928 19944 12980
rect 13084 12792 13136 12844
rect 7012 12699 7064 12708
rect 7012 12665 7021 12699
rect 7021 12665 7055 12699
rect 7055 12665 7064 12699
rect 7012 12656 7064 12665
rect 7472 12699 7524 12708
rect 7472 12665 7481 12699
rect 7481 12665 7515 12699
rect 7515 12665 7524 12699
rect 7472 12656 7524 12665
rect 10876 12656 10928 12708
rect 11612 12656 11664 12708
rect 11980 12724 12032 12776
rect 12440 12724 12492 12776
rect 18788 12860 18840 12912
rect 19156 12860 19208 12912
rect 20352 12860 20404 12912
rect 13820 12792 13872 12844
rect 14188 12792 14240 12844
rect 15752 12792 15804 12844
rect 16304 12792 16356 12844
rect 18512 12835 18564 12844
rect 18512 12801 18521 12835
rect 18521 12801 18555 12835
rect 18555 12801 18564 12835
rect 18512 12792 18564 12801
rect 18880 12792 18932 12844
rect 19524 12792 19576 12844
rect 15016 12724 15068 12776
rect 16212 12767 16264 12776
rect 16212 12733 16221 12767
rect 16221 12733 16255 12767
rect 16255 12733 16264 12767
rect 16212 12724 16264 12733
rect 18236 12724 18288 12776
rect 18420 12724 18472 12776
rect 13912 12699 13964 12708
rect 13912 12665 13921 12699
rect 13921 12665 13955 12699
rect 13955 12665 13964 12699
rect 13912 12656 13964 12665
rect 15108 12656 15160 12708
rect 8300 12588 8352 12640
rect 9220 12631 9272 12640
rect 9220 12597 9229 12631
rect 9229 12597 9263 12631
rect 9263 12597 9272 12631
rect 9220 12588 9272 12597
rect 10140 12631 10192 12640
rect 10140 12597 10149 12631
rect 10149 12597 10183 12631
rect 10183 12597 10192 12631
rect 10140 12588 10192 12597
rect 11980 12631 12032 12640
rect 11980 12597 11989 12631
rect 11989 12597 12023 12631
rect 12023 12597 12032 12631
rect 11980 12588 12032 12597
rect 12348 12631 12400 12640
rect 12348 12597 12357 12631
rect 12357 12597 12391 12631
rect 12391 12597 12400 12631
rect 12348 12588 12400 12597
rect 12532 12588 12584 12640
rect 12900 12588 12952 12640
rect 15200 12588 15252 12640
rect 15844 12631 15896 12640
rect 15844 12597 15853 12631
rect 15853 12597 15887 12631
rect 15887 12597 15896 12631
rect 15844 12588 15896 12597
rect 19616 12724 19668 12776
rect 19708 12724 19760 12776
rect 20628 12792 20680 12844
rect 20536 12724 20588 12776
rect 20720 12767 20772 12776
rect 20720 12733 20729 12767
rect 20729 12733 20763 12767
rect 20763 12733 20772 12767
rect 20720 12724 20772 12733
rect 18788 12656 18840 12708
rect 22468 12767 22520 12776
rect 22468 12733 22477 12767
rect 22477 12733 22511 12767
rect 22511 12733 22520 12767
rect 22468 12724 22520 12733
rect 23112 12928 23164 12980
rect 23848 12928 23900 12980
rect 24308 12860 24360 12912
rect 24676 12928 24728 12980
rect 26240 12928 26292 12980
rect 25320 12860 25372 12912
rect 25504 12792 25556 12844
rect 26884 12835 26936 12844
rect 26884 12801 26893 12835
rect 26893 12801 26927 12835
rect 26927 12801 26936 12835
rect 26884 12792 26936 12801
rect 23112 12767 23164 12776
rect 23112 12733 23121 12767
rect 23121 12733 23155 12767
rect 23155 12733 23164 12767
rect 23112 12724 23164 12733
rect 23664 12724 23716 12776
rect 25228 12724 25280 12776
rect 25320 12767 25372 12776
rect 25320 12733 25329 12767
rect 25329 12733 25363 12767
rect 25363 12733 25372 12767
rect 25320 12724 25372 12733
rect 21088 12699 21140 12708
rect 21088 12665 21097 12699
rect 21097 12665 21131 12699
rect 21131 12665 21140 12699
rect 21088 12656 21140 12665
rect 21180 12699 21232 12708
rect 21180 12665 21189 12699
rect 21189 12665 21223 12699
rect 21223 12665 21232 12699
rect 21180 12656 21232 12665
rect 20996 12588 21048 12640
rect 21456 12631 21508 12640
rect 21456 12597 21465 12631
rect 21465 12597 21499 12631
rect 21499 12597 21508 12631
rect 21456 12588 21508 12597
rect 22560 12631 22612 12640
rect 22560 12597 22569 12631
rect 22569 12597 22603 12631
rect 22603 12597 22612 12631
rect 22560 12588 22612 12597
rect 23388 12699 23440 12708
rect 23388 12665 23397 12699
rect 23397 12665 23431 12699
rect 23431 12665 23440 12699
rect 23388 12656 23440 12665
rect 23572 12699 23624 12708
rect 23572 12665 23581 12699
rect 23581 12665 23615 12699
rect 23615 12665 23624 12699
rect 23572 12656 23624 12665
rect 24952 12656 25004 12708
rect 26608 12699 26660 12708
rect 26608 12665 26626 12699
rect 26626 12665 26660 12699
rect 26608 12656 26660 12665
rect 24676 12631 24728 12640
rect 24676 12597 24685 12631
rect 24685 12597 24719 12631
rect 24719 12597 24728 12631
rect 24676 12588 24728 12597
rect 24768 12631 24820 12640
rect 24768 12597 24777 12631
rect 24777 12597 24811 12631
rect 24811 12597 24820 12631
rect 24768 12588 24820 12597
rect 25044 12588 25096 12640
rect 7114 12486 7166 12538
rect 7178 12486 7230 12538
rect 7242 12486 7294 12538
rect 7306 12486 7358 12538
rect 7370 12486 7422 12538
rect 13830 12486 13882 12538
rect 13894 12486 13946 12538
rect 13958 12486 14010 12538
rect 14022 12486 14074 12538
rect 14086 12486 14138 12538
rect 20546 12486 20598 12538
rect 20610 12486 20662 12538
rect 20674 12486 20726 12538
rect 20738 12486 20790 12538
rect 20802 12486 20854 12538
rect 27262 12486 27314 12538
rect 27326 12486 27378 12538
rect 27390 12486 27442 12538
rect 27454 12486 27506 12538
rect 27518 12486 27570 12538
rect 1952 12384 2004 12436
rect 2780 12384 2832 12436
rect 3240 12384 3292 12436
rect 4160 12384 4212 12436
rect 7748 12427 7800 12436
rect 7748 12393 7757 12427
rect 7757 12393 7791 12427
rect 7791 12393 7800 12427
rect 7748 12384 7800 12393
rect 10140 12427 10192 12436
rect 10140 12393 10149 12427
rect 10149 12393 10183 12427
rect 10183 12393 10192 12427
rect 10140 12384 10192 12393
rect 1032 12291 1084 12300
rect 1032 12257 1041 12291
rect 1041 12257 1075 12291
rect 1075 12257 1084 12291
rect 1032 12248 1084 12257
rect 1676 12291 1728 12300
rect 1676 12257 1685 12291
rect 1685 12257 1719 12291
rect 1719 12257 1728 12291
rect 1676 12248 1728 12257
rect 1768 12291 1820 12300
rect 1768 12257 1777 12291
rect 1777 12257 1811 12291
rect 1811 12257 1820 12291
rect 1768 12248 1820 12257
rect 3516 12316 3568 12368
rect 3976 12316 4028 12368
rect 2504 12248 2556 12300
rect 2964 12291 3016 12300
rect 2964 12257 2973 12291
rect 2973 12257 3007 12291
rect 3007 12257 3016 12291
rect 2964 12248 3016 12257
rect 3148 12291 3200 12300
rect 3148 12257 3157 12291
rect 3157 12257 3191 12291
rect 3191 12257 3200 12291
rect 3148 12248 3200 12257
rect 2780 12180 2832 12232
rect 4988 12291 5040 12300
rect 4988 12257 4997 12291
rect 4997 12257 5031 12291
rect 5031 12257 5040 12291
rect 4988 12248 5040 12257
rect 5080 12248 5132 12300
rect 8944 12316 8996 12368
rect 9680 12316 9732 12368
rect 11980 12384 12032 12436
rect 14740 12384 14792 12436
rect 11520 12316 11572 12368
rect 15660 12384 15712 12436
rect 15844 12384 15896 12436
rect 16212 12384 16264 12436
rect 19616 12427 19668 12436
rect 19616 12393 19625 12427
rect 19625 12393 19659 12427
rect 19659 12393 19668 12427
rect 19616 12384 19668 12393
rect 20904 12384 20956 12436
rect 1124 12044 1176 12096
rect 7012 12248 7064 12300
rect 7656 12291 7708 12300
rect 7656 12257 7665 12291
rect 7665 12257 7699 12291
rect 7699 12257 7708 12291
rect 7656 12248 7708 12257
rect 8208 12248 8260 12300
rect 8300 12291 8352 12300
rect 8300 12257 8309 12291
rect 8309 12257 8343 12291
rect 8343 12257 8352 12291
rect 8300 12248 8352 12257
rect 8484 12291 8536 12300
rect 8484 12257 8493 12291
rect 8493 12257 8527 12291
rect 8527 12257 8536 12291
rect 8484 12248 8536 12257
rect 8668 12248 8720 12300
rect 6552 12180 6604 12232
rect 7564 12223 7616 12232
rect 7564 12189 7573 12223
rect 7573 12189 7607 12223
rect 7607 12189 7616 12223
rect 7564 12180 7616 12189
rect 4436 12044 4488 12096
rect 4804 12044 4856 12096
rect 5448 12044 5500 12096
rect 6460 12044 6512 12096
rect 6828 12044 6880 12096
rect 9128 12248 9180 12300
rect 9312 12291 9364 12300
rect 9312 12257 9321 12291
rect 9321 12257 9355 12291
rect 9355 12257 9364 12291
rect 9312 12248 9364 12257
rect 10048 12223 10100 12232
rect 10048 12189 10057 12223
rect 10057 12189 10091 12223
rect 10091 12189 10100 12223
rect 10048 12180 10100 12189
rect 11060 12291 11112 12300
rect 11060 12257 11069 12291
rect 11069 12257 11103 12291
rect 11103 12257 11112 12291
rect 11060 12248 11112 12257
rect 11888 12248 11940 12300
rect 20260 12359 20312 12368
rect 20260 12325 20269 12359
rect 20269 12325 20303 12359
rect 20303 12325 20312 12359
rect 22008 12384 22060 12436
rect 22468 12384 22520 12436
rect 22928 12384 22980 12436
rect 23112 12384 23164 12436
rect 21548 12359 21600 12368
rect 20260 12316 20312 12325
rect 21548 12325 21560 12359
rect 21560 12325 21600 12359
rect 21548 12316 21600 12325
rect 25320 12384 25372 12436
rect 26608 12427 26660 12436
rect 26608 12393 26617 12427
rect 26617 12393 26651 12427
rect 26651 12393 26660 12427
rect 26608 12384 26660 12393
rect 14556 12291 14608 12300
rect 14556 12257 14565 12291
rect 14565 12257 14599 12291
rect 14599 12257 14608 12291
rect 14556 12248 14608 12257
rect 14832 12248 14884 12300
rect 15660 12248 15712 12300
rect 16672 12248 16724 12300
rect 17960 12291 18012 12300
rect 17960 12257 17994 12291
rect 17994 12257 18012 12291
rect 17960 12248 18012 12257
rect 19524 12291 19576 12300
rect 19524 12257 19533 12291
rect 19533 12257 19567 12291
rect 19567 12257 19576 12291
rect 19524 12248 19576 12257
rect 19800 12248 19852 12300
rect 21272 12291 21324 12300
rect 21272 12257 21281 12291
rect 21281 12257 21315 12291
rect 21315 12257 21324 12291
rect 21272 12248 21324 12257
rect 9312 12044 9364 12096
rect 9588 12087 9640 12096
rect 9588 12053 9597 12087
rect 9597 12053 9631 12087
rect 9631 12053 9640 12087
rect 9588 12044 9640 12053
rect 10324 12044 10376 12096
rect 12532 12044 12584 12096
rect 13360 12044 13412 12096
rect 14372 12044 14424 12096
rect 17684 12044 17736 12096
rect 19984 12180 20036 12232
rect 22836 12223 22888 12232
rect 22836 12189 22845 12223
rect 22845 12189 22879 12223
rect 22879 12189 22888 12223
rect 22836 12180 22888 12189
rect 23664 12316 23716 12368
rect 23848 12248 23900 12300
rect 25964 12316 26016 12368
rect 26884 12316 26936 12368
rect 23572 12180 23624 12232
rect 24768 12180 24820 12232
rect 26424 12291 26476 12300
rect 26424 12257 26433 12291
rect 26433 12257 26467 12291
rect 26467 12257 26476 12291
rect 26424 12248 26476 12257
rect 19064 12087 19116 12096
rect 19064 12053 19073 12087
rect 19073 12053 19107 12087
rect 19107 12053 19116 12087
rect 19064 12044 19116 12053
rect 19156 12087 19208 12096
rect 19156 12053 19165 12087
rect 19165 12053 19199 12087
rect 19199 12053 19208 12087
rect 19156 12044 19208 12053
rect 23388 12044 23440 12096
rect 23756 12044 23808 12096
rect 24860 12044 24912 12096
rect 3756 11942 3808 11994
rect 3820 11942 3872 11994
rect 3884 11942 3936 11994
rect 3948 11942 4000 11994
rect 4012 11942 4064 11994
rect 10472 11942 10524 11994
rect 10536 11942 10588 11994
rect 10600 11942 10652 11994
rect 10664 11942 10716 11994
rect 10728 11942 10780 11994
rect 17188 11942 17240 11994
rect 17252 11942 17304 11994
rect 17316 11942 17368 11994
rect 17380 11942 17432 11994
rect 17444 11942 17496 11994
rect 23904 11942 23956 11994
rect 23968 11942 24020 11994
rect 24032 11942 24084 11994
rect 24096 11942 24148 11994
rect 24160 11942 24212 11994
rect 1216 11679 1268 11688
rect 1216 11645 1225 11679
rect 1225 11645 1259 11679
rect 1259 11645 1268 11679
rect 1216 11636 1268 11645
rect 3332 11840 3384 11892
rect 4068 11840 4120 11892
rect 7472 11840 7524 11892
rect 8484 11840 8536 11892
rect 12440 11883 12492 11892
rect 12440 11849 12449 11883
rect 12449 11849 12483 11883
rect 12483 11849 12492 11883
rect 12440 11840 12492 11849
rect 13728 11840 13780 11892
rect 17960 11883 18012 11892
rect 17960 11849 17969 11883
rect 17969 11849 18003 11883
rect 18003 11849 18012 11883
rect 17960 11840 18012 11849
rect 19524 11840 19576 11892
rect 1768 11679 1820 11688
rect 1768 11645 1777 11679
rect 1777 11645 1811 11679
rect 1811 11645 1820 11679
rect 1768 11636 1820 11645
rect 2688 11772 2740 11824
rect 2964 11772 3016 11824
rect 1492 11543 1544 11552
rect 1492 11509 1501 11543
rect 1501 11509 1535 11543
rect 1535 11509 1544 11543
rect 1492 11500 1544 11509
rect 2504 11636 2556 11688
rect 2688 11636 2740 11688
rect 4988 11772 5040 11824
rect 4436 11704 4488 11756
rect 4896 11704 4948 11756
rect 11060 11704 11112 11756
rect 12348 11704 12400 11756
rect 14740 11704 14792 11756
rect 4528 11679 4580 11688
rect 4528 11645 4537 11679
rect 4537 11645 4571 11679
rect 4571 11645 4580 11679
rect 4528 11636 4580 11645
rect 4620 11679 4672 11688
rect 4620 11645 4629 11679
rect 4629 11645 4663 11679
rect 4663 11645 4672 11679
rect 4620 11636 4672 11645
rect 7564 11636 7616 11688
rect 7748 11568 7800 11620
rect 8760 11679 8812 11688
rect 8760 11645 8769 11679
rect 8769 11645 8803 11679
rect 8803 11645 8812 11679
rect 8760 11636 8812 11645
rect 8852 11679 8904 11688
rect 8852 11645 8861 11679
rect 8861 11645 8895 11679
rect 8895 11645 8904 11679
rect 8852 11636 8904 11645
rect 9128 11636 9180 11688
rect 9312 11636 9364 11688
rect 10324 11568 10376 11620
rect 12072 11679 12124 11688
rect 12072 11645 12081 11679
rect 12081 11645 12115 11679
rect 12115 11645 12124 11679
rect 12072 11636 12124 11645
rect 12900 11679 12952 11688
rect 12900 11645 12909 11679
rect 12909 11645 12943 11679
rect 12943 11645 12952 11679
rect 12900 11636 12952 11645
rect 14464 11636 14516 11688
rect 15752 11747 15804 11756
rect 15752 11713 15761 11747
rect 15761 11713 15795 11747
rect 15795 11713 15804 11747
rect 15752 11704 15804 11713
rect 16948 11704 17000 11756
rect 17684 11704 17736 11756
rect 2136 11500 2188 11552
rect 2780 11500 2832 11552
rect 3240 11500 3292 11552
rect 4160 11500 4212 11552
rect 6552 11500 6604 11552
rect 8392 11543 8444 11552
rect 8392 11509 8401 11543
rect 8401 11509 8435 11543
rect 8435 11509 8444 11543
rect 8392 11500 8444 11509
rect 11244 11500 11296 11552
rect 11612 11543 11664 11552
rect 11612 11509 11621 11543
rect 11621 11509 11655 11543
rect 11655 11509 11664 11543
rect 11612 11500 11664 11509
rect 14188 11568 14240 11620
rect 14280 11568 14332 11620
rect 16580 11636 16632 11688
rect 19156 11772 19208 11824
rect 19064 11704 19116 11756
rect 21272 11840 21324 11892
rect 22836 11840 22888 11892
rect 22928 11840 22980 11892
rect 18236 11636 18288 11688
rect 18696 11679 18748 11688
rect 18696 11645 18705 11679
rect 18705 11645 18739 11679
rect 18739 11645 18748 11679
rect 18696 11636 18748 11645
rect 20352 11679 20404 11688
rect 20352 11645 20370 11679
rect 20370 11645 20404 11679
rect 20352 11636 20404 11645
rect 22560 11636 22612 11688
rect 15016 11568 15068 11620
rect 23020 11568 23072 11620
rect 23480 11840 23532 11892
rect 24584 11840 24636 11892
rect 24768 11883 24820 11892
rect 24768 11849 24777 11883
rect 24777 11849 24811 11883
rect 24811 11849 24820 11883
rect 24768 11840 24820 11849
rect 24952 11840 25004 11892
rect 26884 11840 26936 11892
rect 23572 11772 23624 11824
rect 23388 11704 23440 11756
rect 23572 11679 23624 11688
rect 23572 11645 23581 11679
rect 23581 11645 23615 11679
rect 23615 11645 23624 11679
rect 23572 11636 23624 11645
rect 24952 11704 25004 11756
rect 23388 11568 23440 11620
rect 12992 11543 13044 11552
rect 12992 11509 13001 11543
rect 13001 11509 13035 11543
rect 13035 11509 13044 11543
rect 12992 11500 13044 11509
rect 15108 11543 15160 11552
rect 15108 11509 15117 11543
rect 15117 11509 15151 11543
rect 15151 11509 15160 11543
rect 15108 11500 15160 11509
rect 16580 11500 16632 11552
rect 17408 11543 17460 11552
rect 17408 11509 17417 11543
rect 17417 11509 17451 11543
rect 17451 11509 17460 11543
rect 17408 11500 17460 11509
rect 19248 11543 19300 11552
rect 19248 11509 19257 11543
rect 19257 11509 19291 11543
rect 19291 11509 19300 11543
rect 19248 11500 19300 11509
rect 23296 11500 23348 11552
rect 25136 11636 25188 11688
rect 25044 11611 25096 11620
rect 25044 11577 25053 11611
rect 25053 11577 25087 11611
rect 25087 11577 25096 11611
rect 25044 11568 25096 11577
rect 24492 11500 24544 11552
rect 24676 11500 24728 11552
rect 24768 11500 24820 11552
rect 7114 11398 7166 11450
rect 7178 11398 7230 11450
rect 7242 11398 7294 11450
rect 7306 11398 7358 11450
rect 7370 11398 7422 11450
rect 13830 11398 13882 11450
rect 13894 11398 13946 11450
rect 13958 11398 14010 11450
rect 14022 11398 14074 11450
rect 14086 11398 14138 11450
rect 20546 11398 20598 11450
rect 20610 11398 20662 11450
rect 20674 11398 20726 11450
rect 20738 11398 20790 11450
rect 20802 11398 20854 11450
rect 27262 11398 27314 11450
rect 27326 11398 27378 11450
rect 27390 11398 27442 11450
rect 27454 11398 27506 11450
rect 27518 11398 27570 11450
rect 1768 11296 1820 11348
rect 2136 11296 2188 11348
rect 2964 11296 3016 11348
rect 4620 11339 4672 11348
rect 4620 11305 4629 11339
rect 4629 11305 4663 11339
rect 4663 11305 4672 11339
rect 4620 11296 4672 11305
rect 6920 11296 6972 11348
rect 7748 11339 7800 11348
rect 7748 11305 7757 11339
rect 7757 11305 7791 11339
rect 7791 11305 7800 11339
rect 7748 11296 7800 11305
rect 8392 11296 8444 11348
rect 8760 11296 8812 11348
rect 8852 11296 8904 11348
rect 9588 11296 9640 11348
rect 10048 11296 10100 11348
rect 12992 11296 13044 11348
rect 14188 11296 14240 11348
rect 1124 11203 1176 11212
rect 1124 11169 1158 11203
rect 1158 11169 1176 11203
rect 1124 11160 1176 11169
rect 4804 11228 4856 11280
rect 2964 11203 3016 11212
rect 2964 11169 2998 11203
rect 2998 11169 3016 11203
rect 2964 11160 3016 11169
rect 4068 11160 4120 11212
rect 4252 11160 4304 11212
rect 7472 11228 7524 11280
rect 4988 11203 5040 11212
rect 4988 11169 4997 11203
rect 4997 11169 5031 11203
rect 5031 11169 5040 11203
rect 4988 11160 5040 11169
rect 5448 11160 5500 11212
rect 6552 11203 6604 11212
rect 6552 11169 6561 11203
rect 6561 11169 6595 11203
rect 6595 11169 6604 11203
rect 6552 11160 6604 11169
rect 6644 11203 6696 11212
rect 6644 11169 6653 11203
rect 6653 11169 6687 11203
rect 6687 11169 6696 11203
rect 6644 11160 6696 11169
rect 6736 11160 6788 11212
rect 6828 11203 6880 11212
rect 6828 11169 6837 11203
rect 6837 11169 6871 11203
rect 6871 11169 6880 11203
rect 6828 11160 6880 11169
rect 6920 11203 6972 11212
rect 6920 11169 6929 11203
rect 6929 11169 6963 11203
rect 6963 11169 6972 11203
rect 6920 11160 6972 11169
rect 8668 11160 8720 11212
rect 8944 11160 8996 11212
rect 2504 11024 2556 11076
rect 4160 11024 4212 11076
rect 2136 10956 2188 11008
rect 6092 10956 6144 11008
rect 9680 11228 9732 11280
rect 11612 11228 11664 11280
rect 14556 11296 14608 11348
rect 15016 11339 15068 11348
rect 15016 11305 15025 11339
rect 15025 11305 15059 11339
rect 15059 11305 15068 11339
rect 15016 11296 15068 11305
rect 15108 11296 15160 11348
rect 16580 11296 16632 11348
rect 9772 11160 9824 11212
rect 10048 11203 10100 11212
rect 10048 11169 10057 11203
rect 10057 11169 10091 11203
rect 10091 11169 10100 11203
rect 10048 11160 10100 11169
rect 11244 11160 11296 11212
rect 11888 11203 11940 11212
rect 11888 11169 11904 11203
rect 11904 11169 11938 11203
rect 11938 11169 11940 11203
rect 11888 11160 11940 11169
rect 11060 11024 11112 11076
rect 8484 10956 8536 11008
rect 9404 10956 9456 11008
rect 9772 10956 9824 11008
rect 10232 10999 10284 11008
rect 10232 10965 10241 10999
rect 10241 10965 10275 10999
rect 10275 10965 10284 10999
rect 10232 10956 10284 10965
rect 12992 10956 13044 11008
rect 14188 11160 14240 11212
rect 14280 11203 14332 11212
rect 14280 11169 14289 11203
rect 14289 11169 14323 11203
rect 14323 11169 14332 11203
rect 14280 11160 14332 11169
rect 17408 11296 17460 11348
rect 19800 11339 19852 11348
rect 19800 11305 19809 11339
rect 19809 11305 19843 11339
rect 19843 11305 19852 11339
rect 19800 11296 19852 11305
rect 22836 11296 22888 11348
rect 23572 11296 23624 11348
rect 19248 11228 19300 11280
rect 18420 11203 18472 11212
rect 16672 11092 16724 11144
rect 14832 11024 14884 11076
rect 18420 11169 18429 11203
rect 18429 11169 18463 11203
rect 18463 11169 18472 11203
rect 18420 11160 18472 11169
rect 23480 11228 23532 11280
rect 23756 11228 23808 11280
rect 23020 11160 23072 11212
rect 18236 11092 18288 11144
rect 19432 11135 19484 11144
rect 19432 11101 19441 11135
rect 19441 11101 19475 11135
rect 19475 11101 19484 11135
rect 19432 11092 19484 11101
rect 25320 11160 25372 11212
rect 23664 11135 23716 11144
rect 23664 11101 23673 11135
rect 23673 11101 23707 11135
rect 23707 11101 23716 11135
rect 23664 11092 23716 11101
rect 23388 11024 23440 11076
rect 14280 10956 14332 11008
rect 3756 10854 3808 10906
rect 3820 10854 3872 10906
rect 3884 10854 3936 10906
rect 3948 10854 4000 10906
rect 4012 10854 4064 10906
rect 10472 10854 10524 10906
rect 10536 10854 10588 10906
rect 10600 10854 10652 10906
rect 10664 10854 10716 10906
rect 10728 10854 10780 10906
rect 17188 10854 17240 10906
rect 17252 10854 17304 10906
rect 17316 10854 17368 10906
rect 17380 10854 17432 10906
rect 17444 10854 17496 10906
rect 23904 10854 23956 10906
rect 23968 10854 24020 10906
rect 24032 10854 24084 10906
rect 24096 10854 24148 10906
rect 24160 10854 24212 10906
rect 1124 10752 1176 10804
rect 1676 10752 1728 10804
rect 4988 10752 5040 10804
rect 6736 10752 6788 10804
rect 6828 10752 6880 10804
rect 1492 10616 1544 10668
rect 1032 10591 1084 10600
rect 1032 10557 1041 10591
rect 1041 10557 1075 10591
rect 1075 10557 1084 10591
rect 1032 10548 1084 10557
rect 1216 10591 1268 10600
rect 1216 10557 1225 10591
rect 1225 10557 1259 10591
rect 1259 10557 1268 10591
rect 1216 10548 1268 10557
rect 5540 10684 5592 10736
rect 3332 10616 3384 10668
rect 5816 10684 5868 10736
rect 6276 10727 6328 10736
rect 6276 10693 6285 10727
rect 6285 10693 6319 10727
rect 6319 10693 6328 10727
rect 6276 10684 6328 10693
rect 3700 10591 3752 10600
rect 3700 10557 3709 10591
rect 3709 10557 3743 10591
rect 3743 10557 3752 10591
rect 3700 10548 3752 10557
rect 3516 10480 3568 10532
rect 4988 10548 5040 10600
rect 5172 10591 5224 10600
rect 5172 10557 5181 10591
rect 5181 10557 5215 10591
rect 5215 10557 5224 10591
rect 5172 10548 5224 10557
rect 5540 10591 5592 10600
rect 5540 10557 5549 10591
rect 5549 10557 5583 10591
rect 5583 10557 5592 10591
rect 5540 10548 5592 10557
rect 6552 10548 6604 10600
rect 6736 10591 6788 10600
rect 6736 10557 6745 10591
rect 6745 10557 6779 10591
rect 6779 10557 6788 10591
rect 6736 10548 6788 10557
rect 6828 10591 6880 10600
rect 6828 10557 6837 10591
rect 6837 10557 6871 10591
rect 6871 10557 6880 10591
rect 6828 10548 6880 10557
rect 7472 10591 7524 10600
rect 7472 10557 7481 10591
rect 7481 10557 7515 10591
rect 7515 10557 7524 10591
rect 7472 10548 7524 10557
rect 8208 10591 8260 10600
rect 8208 10557 8217 10591
rect 8217 10557 8251 10591
rect 8251 10557 8260 10591
rect 8208 10548 8260 10557
rect 9128 10548 9180 10600
rect 9404 10591 9456 10600
rect 9404 10557 9413 10591
rect 9413 10557 9447 10591
rect 9447 10557 9456 10591
rect 9404 10548 9456 10557
rect 10048 10752 10100 10804
rect 24952 10795 25004 10804
rect 24952 10761 24961 10795
rect 24961 10761 24995 10795
rect 24995 10761 25004 10795
rect 24952 10752 25004 10761
rect 13084 10684 13136 10736
rect 18144 10684 18196 10736
rect 10232 10616 10284 10668
rect 10140 10591 10192 10600
rect 10140 10557 10149 10591
rect 10149 10557 10183 10591
rect 10183 10557 10192 10591
rect 10140 10548 10192 10557
rect 10876 10548 10928 10600
rect 12164 10591 12216 10600
rect 12164 10557 12173 10591
rect 12173 10557 12207 10591
rect 12207 10557 12216 10591
rect 12164 10548 12216 10557
rect 19432 10616 19484 10668
rect 2320 10412 2372 10464
rect 3056 10412 3108 10464
rect 4160 10412 4212 10464
rect 4804 10455 4856 10464
rect 4804 10421 4813 10455
rect 4813 10421 4847 10455
rect 4847 10421 4856 10455
rect 4804 10412 4856 10421
rect 5172 10412 5224 10464
rect 6276 10412 6328 10464
rect 6368 10455 6420 10464
rect 6368 10421 6377 10455
rect 6377 10421 6411 10455
rect 6411 10421 6420 10455
rect 6368 10412 6420 10421
rect 6460 10412 6512 10464
rect 9680 10480 9732 10532
rect 8024 10455 8076 10464
rect 8024 10421 8033 10455
rect 8033 10421 8067 10455
rect 8067 10421 8076 10455
rect 8024 10412 8076 10421
rect 10784 10412 10836 10464
rect 11980 10455 12032 10464
rect 11980 10421 11989 10455
rect 11989 10421 12023 10455
rect 12023 10421 12032 10455
rect 11980 10412 12032 10421
rect 12992 10548 13044 10600
rect 13636 10548 13688 10600
rect 14924 10591 14976 10600
rect 14924 10557 14933 10591
rect 14933 10557 14967 10591
rect 14967 10557 14976 10591
rect 14924 10548 14976 10557
rect 13452 10480 13504 10532
rect 15660 10548 15712 10600
rect 16028 10591 16080 10600
rect 16028 10557 16037 10591
rect 16037 10557 16071 10591
rect 16071 10557 16080 10591
rect 16028 10548 16080 10557
rect 18420 10548 18472 10600
rect 18604 10480 18656 10532
rect 19064 10548 19116 10600
rect 19248 10548 19300 10600
rect 19708 10591 19760 10600
rect 19708 10557 19717 10591
rect 19717 10557 19751 10591
rect 19751 10557 19760 10591
rect 19708 10548 19760 10557
rect 21272 10616 21324 10668
rect 22284 10659 22336 10668
rect 22284 10625 22293 10659
rect 22293 10625 22327 10659
rect 22327 10625 22336 10659
rect 22284 10616 22336 10625
rect 24492 10616 24544 10668
rect 20352 10523 20404 10532
rect 20352 10489 20361 10523
rect 20361 10489 20395 10523
rect 20395 10489 20404 10523
rect 20352 10480 20404 10489
rect 20904 10548 20956 10600
rect 21548 10548 21600 10600
rect 21916 10548 21968 10600
rect 22192 10548 22244 10600
rect 24676 10548 24728 10600
rect 12900 10412 12952 10464
rect 13084 10412 13136 10464
rect 13268 10455 13320 10464
rect 13268 10421 13277 10455
rect 13277 10421 13311 10455
rect 13311 10421 13320 10455
rect 13268 10412 13320 10421
rect 14740 10455 14792 10464
rect 14740 10421 14749 10455
rect 14749 10421 14783 10455
rect 14783 10421 14792 10455
rect 14740 10412 14792 10421
rect 15200 10455 15252 10464
rect 15200 10421 15209 10455
rect 15209 10421 15243 10455
rect 15243 10421 15252 10455
rect 15200 10412 15252 10421
rect 15476 10412 15528 10464
rect 16764 10412 16816 10464
rect 18788 10455 18840 10464
rect 18788 10421 18797 10455
rect 18797 10421 18831 10455
rect 18831 10421 18840 10455
rect 18788 10412 18840 10421
rect 18880 10412 18932 10464
rect 19892 10455 19944 10464
rect 19892 10421 19901 10455
rect 19901 10421 19935 10455
rect 19935 10421 19944 10455
rect 19892 10412 19944 10421
rect 20996 10412 21048 10464
rect 21088 10412 21140 10464
rect 7114 10310 7166 10362
rect 7178 10310 7230 10362
rect 7242 10310 7294 10362
rect 7306 10310 7358 10362
rect 7370 10310 7422 10362
rect 13830 10310 13882 10362
rect 13894 10310 13946 10362
rect 13958 10310 14010 10362
rect 14022 10310 14074 10362
rect 14086 10310 14138 10362
rect 20546 10310 20598 10362
rect 20610 10310 20662 10362
rect 20674 10310 20726 10362
rect 20738 10310 20790 10362
rect 20802 10310 20854 10362
rect 27262 10310 27314 10362
rect 27326 10310 27378 10362
rect 27390 10310 27442 10362
rect 27454 10310 27506 10362
rect 27518 10310 27570 10362
rect 1860 10251 1912 10260
rect 1860 10217 1869 10251
rect 1869 10217 1903 10251
rect 1903 10217 1912 10251
rect 1860 10208 1912 10217
rect 2688 10208 2740 10260
rect 3700 10208 3752 10260
rect 4896 10251 4948 10260
rect 4896 10217 4905 10251
rect 4905 10217 4939 10251
rect 4939 10217 4948 10251
rect 4896 10208 4948 10217
rect 6644 10208 6696 10260
rect 7564 10208 7616 10260
rect 8024 10208 8076 10260
rect 8944 10208 8996 10260
rect 10140 10208 10192 10260
rect 10784 10208 10836 10260
rect 13452 10251 13504 10260
rect 13452 10217 13461 10251
rect 13461 10217 13495 10251
rect 13495 10217 13504 10251
rect 13452 10208 13504 10217
rect 14556 10208 14608 10260
rect 15936 10208 15988 10260
rect 16028 10208 16080 10260
rect 3148 10140 3200 10192
rect 3608 10183 3660 10192
rect 3608 10149 3617 10183
rect 3617 10149 3651 10183
rect 3651 10149 3660 10183
rect 3608 10140 3660 10149
rect 5816 10183 5868 10192
rect 5816 10149 5825 10183
rect 5825 10149 5859 10183
rect 5859 10149 5868 10183
rect 5816 10140 5868 10149
rect 1308 10004 1360 10056
rect 1860 10072 1912 10124
rect 2412 10115 2464 10124
rect 2412 10081 2446 10115
rect 2446 10081 2464 10115
rect 2412 10072 2464 10081
rect 6092 10115 6144 10124
rect 6092 10081 6101 10115
rect 6101 10081 6135 10115
rect 6135 10081 6144 10115
rect 6092 10072 6144 10081
rect 6460 10072 6512 10124
rect 6920 10072 6972 10124
rect 10876 10140 10928 10192
rect 14740 10183 14792 10192
rect 2136 10047 2188 10056
rect 2136 10013 2145 10047
rect 2145 10013 2179 10047
rect 2179 10013 2188 10047
rect 2136 10004 2188 10013
rect 6000 10047 6052 10056
rect 6000 10013 6009 10047
rect 6009 10013 6043 10047
rect 6043 10013 6052 10047
rect 6000 10004 6052 10013
rect 9496 10072 9548 10124
rect 10968 10072 11020 10124
rect 11060 10115 11112 10124
rect 11060 10081 11069 10115
rect 11069 10081 11103 10115
rect 11103 10081 11112 10115
rect 11060 10072 11112 10081
rect 12992 10115 13044 10124
rect 12992 10081 13001 10115
rect 13001 10081 13035 10115
rect 13035 10081 13044 10115
rect 12992 10072 13044 10081
rect 13084 10072 13136 10124
rect 13268 10115 13320 10124
rect 13268 10081 13277 10115
rect 13277 10081 13311 10115
rect 13311 10081 13320 10115
rect 13268 10072 13320 10081
rect 13360 10115 13412 10124
rect 13360 10081 13369 10115
rect 13369 10081 13403 10115
rect 13403 10081 13412 10115
rect 13360 10072 13412 10081
rect 14188 10072 14240 10124
rect 14280 10115 14332 10124
rect 14280 10081 14289 10115
rect 14289 10081 14323 10115
rect 14323 10081 14332 10115
rect 14280 10072 14332 10081
rect 14740 10149 14763 10183
rect 14763 10149 14792 10183
rect 14740 10140 14792 10149
rect 18788 10208 18840 10260
rect 16580 10140 16632 10192
rect 2044 9868 2096 9920
rect 2504 9868 2556 9920
rect 3056 9868 3108 9920
rect 6460 9911 6512 9920
rect 6460 9877 6469 9911
rect 6469 9877 6503 9911
rect 6503 9877 6512 9911
rect 6460 9868 6512 9877
rect 8668 9868 8720 9920
rect 13084 9868 13136 9920
rect 17776 10115 17828 10124
rect 17776 10081 17785 10115
rect 17785 10081 17819 10115
rect 17819 10081 17828 10115
rect 17776 10072 17828 10081
rect 18604 10115 18656 10124
rect 18604 10081 18613 10115
rect 18613 10081 18647 10115
rect 18647 10081 18656 10115
rect 18604 10072 18656 10081
rect 19892 10208 19944 10260
rect 21272 10251 21324 10260
rect 21272 10217 21281 10251
rect 21281 10217 21315 10251
rect 21315 10217 21324 10251
rect 21272 10208 21324 10217
rect 14464 10047 14516 10056
rect 14464 10013 14473 10047
rect 14473 10013 14507 10047
rect 14507 10013 14516 10047
rect 14464 10004 14516 10013
rect 15568 10004 15620 10056
rect 15752 10004 15804 10056
rect 15936 10004 15988 10056
rect 14464 9868 14516 9920
rect 17684 9936 17736 9988
rect 18696 10004 18748 10056
rect 19156 10004 19208 10056
rect 19340 10004 19392 10056
rect 19984 10047 20036 10056
rect 19984 10013 19993 10047
rect 19993 10013 20027 10047
rect 20027 10013 20036 10047
rect 19984 10004 20036 10013
rect 21180 10140 21232 10192
rect 22100 10072 22152 10124
rect 23664 10072 23716 10124
rect 24676 10115 24728 10124
rect 24676 10081 24685 10115
rect 24685 10081 24719 10115
rect 24719 10081 24728 10115
rect 24676 10072 24728 10081
rect 21088 10047 21140 10056
rect 21088 10013 21097 10047
rect 21097 10013 21131 10047
rect 21131 10013 21140 10047
rect 21088 10004 21140 10013
rect 15476 9868 15528 9920
rect 17592 9868 17644 9920
rect 19064 9911 19116 9920
rect 19064 9877 19073 9911
rect 19073 9877 19107 9911
rect 19107 9877 19116 9911
rect 19064 9868 19116 9877
rect 20996 9868 21048 9920
rect 24860 9911 24912 9920
rect 24860 9877 24869 9911
rect 24869 9877 24903 9911
rect 24903 9877 24912 9911
rect 24860 9868 24912 9877
rect 3756 9766 3808 9818
rect 3820 9766 3872 9818
rect 3884 9766 3936 9818
rect 3948 9766 4000 9818
rect 4012 9766 4064 9818
rect 10472 9766 10524 9818
rect 10536 9766 10588 9818
rect 10600 9766 10652 9818
rect 10664 9766 10716 9818
rect 10728 9766 10780 9818
rect 17188 9766 17240 9818
rect 17252 9766 17304 9818
rect 17316 9766 17368 9818
rect 17380 9766 17432 9818
rect 17444 9766 17496 9818
rect 23904 9766 23956 9818
rect 23968 9766 24020 9818
rect 24032 9766 24084 9818
rect 24096 9766 24148 9818
rect 24160 9766 24212 9818
rect 2228 9664 2280 9716
rect 2688 9664 2740 9716
rect 3516 9664 3568 9716
rect 2964 9596 3016 9648
rect 4344 9596 4396 9648
rect 4896 9664 4948 9716
rect 5816 9664 5868 9716
rect 6920 9664 6972 9716
rect 7472 9664 7524 9716
rect 8208 9707 8260 9716
rect 8208 9673 8217 9707
rect 8217 9673 8251 9707
rect 8251 9673 8260 9707
rect 8208 9664 8260 9673
rect 8852 9571 8904 9580
rect 8852 9537 8861 9571
rect 8861 9537 8895 9571
rect 8895 9537 8904 9571
rect 8852 9528 8904 9537
rect 9036 9571 9088 9580
rect 9036 9537 9045 9571
rect 9045 9537 9079 9571
rect 9079 9537 9088 9571
rect 9036 9528 9088 9537
rect 9312 9639 9364 9648
rect 9312 9605 9321 9639
rect 9321 9605 9355 9639
rect 9355 9605 9364 9639
rect 9312 9596 9364 9605
rect 10968 9664 11020 9716
rect 11060 9664 11112 9716
rect 14924 9707 14976 9716
rect 14924 9673 14933 9707
rect 14933 9673 14967 9707
rect 14967 9673 14976 9707
rect 14924 9664 14976 9673
rect 2136 9460 2188 9512
rect 1952 9435 2004 9444
rect 1952 9401 1970 9435
rect 1970 9401 2004 9435
rect 1952 9392 2004 9401
rect 2504 9460 2556 9512
rect 2596 9503 2648 9512
rect 2596 9469 2605 9503
rect 2605 9469 2639 9503
rect 2639 9469 2648 9503
rect 2596 9460 2648 9469
rect 2688 9503 2740 9512
rect 2688 9469 2697 9503
rect 2697 9469 2731 9503
rect 2731 9469 2740 9503
rect 2688 9460 2740 9469
rect 3240 9460 3292 9512
rect 3424 9460 3476 9512
rect 3884 9460 3936 9512
rect 4804 9503 4856 9512
rect 4804 9469 4838 9503
rect 4838 9469 4856 9503
rect 4804 9460 4856 9469
rect 7932 9460 7984 9512
rect 848 9367 900 9376
rect 848 9333 857 9367
rect 857 9333 891 9367
rect 891 9333 900 9367
rect 848 9324 900 9333
rect 2320 9324 2372 9376
rect 2504 9324 2556 9376
rect 2964 9324 3016 9376
rect 6000 9392 6052 9444
rect 6368 9392 6420 9444
rect 8668 9392 8720 9444
rect 9496 9460 9548 9512
rect 10140 9528 10192 9580
rect 12808 9596 12860 9648
rect 17776 9664 17828 9716
rect 12164 9528 12216 9580
rect 17684 9596 17736 9648
rect 19340 9664 19392 9716
rect 19708 9664 19760 9716
rect 20260 9664 20312 9716
rect 20904 9664 20956 9716
rect 21088 9664 21140 9716
rect 10324 9435 10376 9444
rect 10324 9401 10333 9435
rect 10333 9401 10367 9435
rect 10367 9401 10376 9435
rect 12348 9460 12400 9512
rect 12624 9503 12676 9512
rect 12624 9469 12633 9503
rect 12633 9469 12667 9503
rect 12667 9469 12676 9503
rect 12624 9460 12676 9469
rect 13176 9503 13228 9512
rect 13176 9469 13185 9503
rect 13185 9469 13219 9503
rect 13219 9469 13228 9503
rect 13176 9460 13228 9469
rect 15752 9528 15804 9580
rect 10324 9392 10376 9401
rect 12992 9392 13044 9444
rect 14188 9503 14240 9512
rect 14188 9469 14197 9503
rect 14197 9469 14231 9503
rect 14231 9469 14240 9503
rect 14188 9460 14240 9469
rect 14372 9503 14424 9512
rect 14372 9469 14381 9503
rect 14381 9469 14415 9503
rect 14415 9469 14424 9503
rect 14372 9460 14424 9469
rect 14464 9503 14516 9512
rect 14464 9469 14473 9503
rect 14473 9469 14507 9503
rect 14507 9469 14516 9503
rect 14464 9460 14516 9469
rect 15200 9460 15252 9512
rect 16672 9460 16724 9512
rect 17132 9460 17184 9512
rect 22100 9596 22152 9648
rect 23480 9596 23532 9648
rect 24308 9528 24360 9580
rect 25964 9571 26016 9580
rect 25964 9537 25973 9571
rect 25973 9537 26007 9571
rect 26007 9537 26016 9571
rect 25964 9528 26016 9537
rect 17592 9503 17644 9512
rect 17592 9469 17601 9503
rect 17601 9469 17635 9503
rect 17635 9469 17644 9503
rect 17592 9460 17644 9469
rect 18052 9503 18104 9512
rect 18052 9469 18061 9503
rect 18061 9469 18095 9503
rect 18095 9469 18104 9503
rect 18052 9460 18104 9469
rect 18144 9503 18196 9512
rect 18144 9469 18153 9503
rect 18153 9469 18187 9503
rect 18187 9469 18196 9503
rect 18144 9460 18196 9469
rect 19064 9460 19116 9512
rect 6460 9324 6512 9376
rect 9220 9367 9272 9376
rect 9220 9333 9229 9367
rect 9229 9333 9263 9367
rect 9263 9333 9272 9367
rect 9220 9324 9272 9333
rect 9496 9367 9548 9376
rect 9496 9333 9505 9367
rect 9505 9333 9539 9367
rect 9539 9333 9548 9367
rect 9496 9324 9548 9333
rect 9956 9367 10008 9376
rect 9956 9333 9965 9367
rect 9965 9333 9999 9367
rect 9999 9333 10008 9367
rect 9956 9324 10008 9333
rect 10140 9367 10192 9376
rect 10140 9333 10167 9367
rect 10167 9333 10192 9367
rect 10140 9324 10192 9333
rect 12532 9367 12584 9376
rect 12532 9333 12541 9367
rect 12541 9333 12575 9367
rect 12575 9333 12584 9367
rect 12532 9324 12584 9333
rect 14648 9324 14700 9376
rect 15384 9324 15436 9376
rect 15844 9367 15896 9376
rect 15844 9333 15853 9367
rect 15853 9333 15887 9367
rect 15887 9333 15896 9367
rect 15844 9324 15896 9333
rect 16764 9392 16816 9444
rect 17408 9367 17460 9376
rect 17408 9333 17417 9367
rect 17417 9333 17451 9367
rect 17451 9333 17460 9367
rect 17408 9324 17460 9333
rect 18972 9324 19024 9376
rect 20996 9367 21048 9376
rect 20996 9333 21005 9367
rect 21005 9333 21039 9367
rect 21039 9333 21048 9367
rect 20996 9324 21048 9333
rect 21272 9392 21324 9444
rect 22192 9460 22244 9512
rect 23020 9460 23072 9512
rect 21916 9392 21968 9444
rect 23112 9367 23164 9376
rect 23112 9333 23121 9367
rect 23121 9333 23155 9367
rect 23155 9333 23164 9367
rect 24860 9460 24912 9512
rect 23112 9324 23164 9333
rect 24400 9367 24452 9376
rect 24400 9333 24409 9367
rect 24409 9333 24443 9367
rect 24443 9333 24452 9367
rect 24400 9324 24452 9333
rect 7114 9222 7166 9274
rect 7178 9222 7230 9274
rect 7242 9222 7294 9274
rect 7306 9222 7358 9274
rect 7370 9222 7422 9274
rect 13830 9222 13882 9274
rect 13894 9222 13946 9274
rect 13958 9222 14010 9274
rect 14022 9222 14074 9274
rect 14086 9222 14138 9274
rect 20546 9222 20598 9274
rect 20610 9222 20662 9274
rect 20674 9222 20726 9274
rect 20738 9222 20790 9274
rect 20802 9222 20854 9274
rect 27262 9222 27314 9274
rect 27326 9222 27378 9274
rect 27390 9222 27442 9274
rect 27454 9222 27506 9274
rect 27518 9222 27570 9274
rect 1308 9120 1360 9172
rect 3148 9163 3200 9172
rect 3148 9129 3157 9163
rect 3157 9129 3191 9163
rect 3191 9129 3200 9163
rect 3148 9120 3200 9129
rect 3332 9120 3384 9172
rect 6000 9120 6052 9172
rect 848 8984 900 9036
rect 1676 8984 1728 9036
rect 1860 8984 1912 9036
rect 2044 8984 2096 9036
rect 2136 9030 2188 9036
rect 2136 8996 2145 9030
rect 2145 8996 2179 9030
rect 2179 8996 2188 9030
rect 2136 8984 2188 8996
rect 2228 9027 2280 9036
rect 2228 8993 2237 9027
rect 2237 8993 2271 9027
rect 2271 8993 2280 9027
rect 2228 8984 2280 8993
rect 2504 9052 2556 9104
rect 8852 9120 8904 9172
rect 9036 9120 9088 9172
rect 9220 9120 9272 9172
rect 12808 9120 12860 9172
rect 12900 9120 12952 9172
rect 2412 8916 2464 8968
rect 2872 8916 2924 8968
rect 3056 8984 3108 9036
rect 3424 8984 3476 9036
rect 4160 9027 4212 9036
rect 4160 8993 4194 9027
rect 4194 8993 4212 9027
rect 4160 8984 4212 8993
rect 7472 9027 7524 9036
rect 7472 8993 7481 9027
rect 7481 8993 7515 9027
rect 7515 8993 7524 9027
rect 7472 8984 7524 8993
rect 7932 9027 7984 9036
rect 7932 8993 7946 9027
rect 7946 8993 7980 9027
rect 7980 8993 7984 9027
rect 7932 8984 7984 8993
rect 3884 8959 3936 8968
rect 3884 8925 3893 8959
rect 3893 8925 3927 8959
rect 3927 8925 3936 8959
rect 3884 8916 3936 8925
rect 2964 8848 3016 8900
rect 9496 9052 9548 9104
rect 9404 8984 9456 9036
rect 9956 8984 10008 9036
rect 10140 8984 10192 9036
rect 11060 9027 11112 9036
rect 11060 8993 11069 9027
rect 11069 8993 11103 9027
rect 11103 8993 11112 9027
rect 11060 8984 11112 8993
rect 14096 9120 14148 9172
rect 13176 8984 13228 9036
rect 13360 9027 13412 9036
rect 13360 8993 13369 9027
rect 13369 8993 13403 9027
rect 13403 8993 13412 9027
rect 13360 8984 13412 8993
rect 13728 8984 13780 9036
rect 14188 8984 14240 9036
rect 9496 8916 9548 8968
rect 8024 8823 8076 8832
rect 8024 8789 8033 8823
rect 8033 8789 8067 8823
rect 8067 8789 8076 8823
rect 8024 8780 8076 8789
rect 12440 8916 12492 8968
rect 14464 8984 14516 9036
rect 14924 9027 14976 9036
rect 14924 8993 14933 9027
rect 14933 8993 14967 9027
rect 14967 8993 14976 9027
rect 14924 8984 14976 8993
rect 15476 8984 15528 9036
rect 15384 8916 15436 8968
rect 9128 8780 9180 8832
rect 9680 8780 9732 8832
rect 13544 8823 13596 8832
rect 13544 8789 13553 8823
rect 13553 8789 13587 8823
rect 13587 8789 13596 8823
rect 13544 8780 13596 8789
rect 14280 8780 14332 8832
rect 14740 8780 14792 8832
rect 15108 8823 15160 8832
rect 15108 8789 15117 8823
rect 15117 8789 15151 8823
rect 15151 8789 15160 8823
rect 15108 8780 15160 8789
rect 15844 9120 15896 9172
rect 16580 9163 16632 9172
rect 16580 9129 16589 9163
rect 16589 9129 16623 9163
rect 16623 9129 16632 9163
rect 16580 9120 16632 9129
rect 18052 9120 18104 9172
rect 18880 9120 18932 9172
rect 17408 9095 17460 9104
rect 15660 8984 15712 9036
rect 17408 9061 17431 9095
rect 17431 9061 17460 9095
rect 17408 9052 17460 9061
rect 18144 8984 18196 9036
rect 18788 8984 18840 9036
rect 17040 8916 17092 8968
rect 18972 9027 19024 9036
rect 18972 8993 18981 9027
rect 18981 8993 19015 9027
rect 19015 8993 19024 9027
rect 18972 8984 19024 8993
rect 19340 9120 19392 9172
rect 19524 9052 19576 9104
rect 23112 9120 23164 9172
rect 23480 9120 23532 9172
rect 24400 9120 24452 9172
rect 24676 9120 24728 9172
rect 18604 8848 18656 8900
rect 19248 8848 19300 8900
rect 20260 9027 20312 9036
rect 20260 8993 20269 9027
rect 20269 8993 20303 9027
rect 20303 8993 20312 9027
rect 20260 8984 20312 8993
rect 22652 9027 22704 9036
rect 22652 8993 22661 9027
rect 22661 8993 22695 9027
rect 22695 8993 22704 9027
rect 22652 8984 22704 8993
rect 20628 8916 20680 8968
rect 22284 8916 22336 8968
rect 22836 8848 22888 8900
rect 23112 8984 23164 9036
rect 23572 9027 23624 9036
rect 23572 8993 23581 9027
rect 23581 8993 23615 9027
rect 23615 8993 23624 9027
rect 23572 8984 23624 8993
rect 23480 8848 23532 8900
rect 24400 8959 24452 8968
rect 24400 8925 24409 8959
rect 24409 8925 24443 8959
rect 24443 8925 24452 8959
rect 24400 8916 24452 8925
rect 21088 8780 21140 8832
rect 22008 8780 22060 8832
rect 22928 8780 22980 8832
rect 23020 8780 23072 8832
rect 3756 8678 3808 8730
rect 3820 8678 3872 8730
rect 3884 8678 3936 8730
rect 3948 8678 4000 8730
rect 4012 8678 4064 8730
rect 10472 8678 10524 8730
rect 10536 8678 10588 8730
rect 10600 8678 10652 8730
rect 10664 8678 10716 8730
rect 10728 8678 10780 8730
rect 17188 8678 17240 8730
rect 17252 8678 17304 8730
rect 17316 8678 17368 8730
rect 17380 8678 17432 8730
rect 17444 8678 17496 8730
rect 23904 8678 23956 8730
rect 23968 8678 24020 8730
rect 24032 8678 24084 8730
rect 24096 8678 24148 8730
rect 24160 8678 24212 8730
rect 1584 8440 1636 8492
rect 1676 8483 1728 8492
rect 1676 8449 1685 8483
rect 1685 8449 1719 8483
rect 1719 8449 1728 8483
rect 1676 8440 1728 8449
rect 1952 8440 2004 8492
rect 1860 8372 1912 8424
rect 2596 8619 2648 8628
rect 2596 8585 2605 8619
rect 2605 8585 2639 8619
rect 2639 8585 2648 8619
rect 2596 8576 2648 8585
rect 8852 8576 8904 8628
rect 10324 8576 10376 8628
rect 18052 8576 18104 8628
rect 2412 8508 2464 8560
rect 2872 8508 2924 8560
rect 12900 8508 12952 8560
rect 14372 8508 14424 8560
rect 16856 8508 16908 8560
rect 18144 8508 18196 8560
rect 11060 8483 11112 8492
rect 11060 8449 11069 8483
rect 11069 8449 11103 8483
rect 11103 8449 11112 8483
rect 11060 8440 11112 8449
rect 12532 8440 12584 8492
rect 12624 8483 12676 8492
rect 12624 8449 12633 8483
rect 12633 8449 12667 8483
rect 12667 8449 12676 8483
rect 12624 8440 12676 8449
rect 14740 8440 14792 8492
rect 2412 8415 2464 8424
rect 2412 8381 2421 8415
rect 2421 8381 2455 8415
rect 2455 8381 2464 8415
rect 2412 8372 2464 8381
rect 2872 8372 2924 8424
rect 6092 8372 6144 8424
rect 9220 8415 9272 8424
rect 9220 8381 9229 8415
rect 9229 8381 9263 8415
rect 9263 8381 9272 8415
rect 9220 8372 9272 8381
rect 10968 8415 11020 8424
rect 10968 8381 10977 8415
rect 10977 8381 11011 8415
rect 11011 8381 11020 8415
rect 10968 8372 11020 8381
rect 12348 8372 12400 8424
rect 13176 8372 13228 8424
rect 2780 8347 2832 8356
rect 2780 8313 2789 8347
rect 2789 8313 2823 8347
rect 2823 8313 2832 8347
rect 2780 8304 2832 8313
rect 3056 8304 3108 8356
rect 3148 8304 3200 8356
rect 6368 8304 6420 8356
rect 8024 8304 8076 8356
rect 9496 8347 9548 8356
rect 9496 8313 9530 8347
rect 9530 8313 9548 8347
rect 9496 8304 9548 8313
rect 12808 8347 12860 8356
rect 12808 8313 12817 8347
rect 12817 8313 12851 8347
rect 12851 8313 12860 8347
rect 12808 8304 12860 8313
rect 14464 8415 14516 8424
rect 14464 8381 14473 8415
rect 14473 8381 14507 8415
rect 14507 8381 14516 8415
rect 14464 8372 14516 8381
rect 14924 8415 14976 8424
rect 14924 8381 14933 8415
rect 14933 8381 14967 8415
rect 14967 8381 14976 8415
rect 14924 8372 14976 8381
rect 13728 8304 13780 8356
rect 16212 8415 16264 8424
rect 16212 8381 16221 8415
rect 16221 8381 16255 8415
rect 16255 8381 16264 8415
rect 16212 8372 16264 8381
rect 17592 8372 17644 8424
rect 21824 8576 21876 8628
rect 22928 8619 22980 8628
rect 22928 8585 22937 8619
rect 22937 8585 22971 8619
rect 22971 8585 22980 8619
rect 22928 8576 22980 8585
rect 19616 8440 19668 8492
rect 20628 8483 20680 8492
rect 20628 8449 20637 8483
rect 20637 8449 20671 8483
rect 20671 8449 20680 8483
rect 20628 8440 20680 8449
rect 22008 8508 22060 8560
rect 24216 8576 24268 8628
rect 24400 8576 24452 8628
rect 18604 8372 18656 8424
rect 19156 8372 19208 8424
rect 20444 8415 20496 8424
rect 20444 8381 20453 8415
rect 20453 8381 20487 8415
rect 20487 8381 20496 8415
rect 20444 8372 20496 8381
rect 21640 8372 21692 8424
rect 22100 8440 22152 8492
rect 22836 8440 22888 8492
rect 22008 8372 22060 8424
rect 22928 8347 22980 8356
rect 22928 8313 22937 8347
rect 22937 8313 22971 8347
rect 22971 8313 22980 8347
rect 22928 8304 22980 8313
rect 23112 8415 23164 8424
rect 23112 8381 23121 8415
rect 23121 8381 23155 8415
rect 23155 8381 23164 8415
rect 23112 8372 23164 8381
rect 23388 8440 23440 8492
rect 25136 8551 25188 8560
rect 25136 8517 25145 8551
rect 25145 8517 25179 8551
rect 25179 8517 25188 8551
rect 25136 8508 25188 8517
rect 23480 8415 23532 8424
rect 23480 8381 23489 8415
rect 23489 8381 23523 8415
rect 23523 8381 23532 8415
rect 23480 8372 23532 8381
rect 23572 8372 23624 8424
rect 23756 8372 23808 8424
rect 24216 8415 24268 8424
rect 24216 8381 24225 8415
rect 24225 8381 24259 8415
rect 24259 8381 24268 8415
rect 24216 8372 24268 8381
rect 24768 8440 24820 8492
rect 25596 8415 25648 8424
rect 25596 8381 25605 8415
rect 25605 8381 25639 8415
rect 25639 8381 25648 8415
rect 25596 8372 25648 8381
rect 24584 8304 24636 8356
rect 24768 8347 24820 8356
rect 24768 8313 24777 8347
rect 24777 8313 24811 8347
rect 24811 8313 24820 8347
rect 24768 8304 24820 8313
rect 26240 8304 26292 8356
rect 2412 8236 2464 8288
rect 4160 8236 4212 8288
rect 4620 8279 4672 8288
rect 4620 8245 4629 8279
rect 4629 8245 4663 8279
rect 4663 8245 4672 8279
rect 4620 8236 4672 8245
rect 6644 8279 6696 8288
rect 6644 8245 6653 8279
rect 6653 8245 6687 8279
rect 6687 8245 6696 8279
rect 6644 8236 6696 8245
rect 13360 8236 13412 8288
rect 13636 8236 13688 8288
rect 15016 8236 15068 8288
rect 18052 8236 18104 8288
rect 18420 8279 18472 8288
rect 18420 8245 18429 8279
rect 18429 8245 18463 8279
rect 18463 8245 18472 8279
rect 18420 8236 18472 8245
rect 19432 8236 19484 8288
rect 20904 8279 20956 8288
rect 20904 8245 20913 8279
rect 20913 8245 20947 8279
rect 20947 8245 20956 8279
rect 20904 8236 20956 8245
rect 21640 8236 21692 8288
rect 21916 8279 21968 8288
rect 21916 8245 21925 8279
rect 21925 8245 21959 8279
rect 21959 8245 21968 8279
rect 21916 8236 21968 8245
rect 25228 8279 25280 8288
rect 25228 8245 25237 8279
rect 25237 8245 25271 8279
rect 25271 8245 25280 8279
rect 25228 8236 25280 8245
rect 7114 8134 7166 8186
rect 7178 8134 7230 8186
rect 7242 8134 7294 8186
rect 7306 8134 7358 8186
rect 7370 8134 7422 8186
rect 13830 8134 13882 8186
rect 13894 8134 13946 8186
rect 13958 8134 14010 8186
rect 14022 8134 14074 8186
rect 14086 8134 14138 8186
rect 20546 8134 20598 8186
rect 20610 8134 20662 8186
rect 20674 8134 20726 8186
rect 20738 8134 20790 8186
rect 20802 8134 20854 8186
rect 27262 8134 27314 8186
rect 27326 8134 27378 8186
rect 27390 8134 27442 8186
rect 27454 8134 27506 8186
rect 27518 8134 27570 8186
rect 2136 8032 2188 8084
rect 3056 8007 3108 8016
rect 3056 7973 3065 8007
rect 3065 7973 3099 8007
rect 3099 7973 3108 8007
rect 3056 7964 3108 7973
rect 3332 7964 3384 8016
rect 3516 7964 3568 8016
rect 3240 7896 3292 7948
rect 2964 7828 3016 7880
rect 3148 7760 3200 7812
rect 3608 7828 3660 7880
rect 4160 7939 4212 7948
rect 4160 7905 4169 7939
rect 4169 7905 4203 7939
rect 4203 7905 4212 7939
rect 4160 7896 4212 7905
rect 6368 8075 6420 8084
rect 6368 8041 6377 8075
rect 6377 8041 6411 8075
rect 6411 8041 6420 8075
rect 6368 8032 6420 8041
rect 9496 8075 9548 8084
rect 9496 8041 9505 8075
rect 9505 8041 9539 8075
rect 9539 8041 9548 8075
rect 9496 8032 9548 8041
rect 9680 8032 9732 8084
rect 12532 8032 12584 8084
rect 14188 8032 14240 8084
rect 5080 7939 5132 7948
rect 5080 7905 5089 7939
rect 5089 7905 5123 7939
rect 5123 7905 5132 7939
rect 5080 7896 5132 7905
rect 6828 7939 6880 7948
rect 6828 7905 6837 7939
rect 6837 7905 6871 7939
rect 6871 7905 6880 7939
rect 6828 7896 6880 7905
rect 11888 7939 11940 7948
rect 11888 7905 11897 7939
rect 11897 7905 11931 7939
rect 11931 7905 11940 7939
rect 11888 7896 11940 7905
rect 12440 7964 12492 8016
rect 4344 7871 4396 7880
rect 4344 7837 4353 7871
rect 4353 7837 4387 7871
rect 4387 7837 4396 7871
rect 4344 7828 4396 7837
rect 8852 7828 8904 7880
rect 12348 7939 12400 7948
rect 12348 7905 12357 7939
rect 12357 7905 12391 7939
rect 12391 7905 12400 7939
rect 12348 7896 12400 7905
rect 12532 7939 12584 7948
rect 12532 7905 12541 7939
rect 12541 7905 12575 7939
rect 12575 7905 12584 7939
rect 12532 7896 12584 7905
rect 14924 8032 14976 8084
rect 18420 8032 18472 8084
rect 16856 7964 16908 8016
rect 17040 7964 17092 8016
rect 14556 7939 14608 7948
rect 14556 7905 14565 7939
rect 14565 7905 14599 7939
rect 14599 7905 14608 7939
rect 14556 7896 14608 7905
rect 14832 7939 14884 7948
rect 14832 7905 14841 7939
rect 14841 7905 14875 7939
rect 14875 7905 14884 7939
rect 14832 7896 14884 7905
rect 15108 7896 15160 7948
rect 15200 7896 15252 7948
rect 18144 7896 18196 7948
rect 4436 7760 4488 7812
rect 12164 7828 12216 7880
rect 12900 7828 12952 7880
rect 4252 7692 4304 7744
rect 14556 7760 14608 7812
rect 15384 7871 15436 7880
rect 15384 7837 15393 7871
rect 15393 7837 15427 7871
rect 15427 7837 15436 7871
rect 15384 7828 15436 7837
rect 19156 8032 19208 8084
rect 20904 8032 20956 8084
rect 21824 8032 21876 8084
rect 22100 8032 22152 8084
rect 22652 8032 22704 8084
rect 19064 7939 19116 7948
rect 19064 7905 19073 7939
rect 19073 7905 19107 7939
rect 19107 7905 19116 7939
rect 19064 7896 19116 7905
rect 19248 7896 19300 7948
rect 19340 7939 19392 7948
rect 19340 7905 19349 7939
rect 19349 7905 19383 7939
rect 19383 7905 19392 7939
rect 19340 7896 19392 7905
rect 21640 7939 21692 7948
rect 21640 7905 21649 7939
rect 21649 7905 21683 7939
rect 21683 7905 21692 7939
rect 21640 7896 21692 7905
rect 21916 7896 21968 7948
rect 23756 8032 23808 8084
rect 24216 8032 24268 8084
rect 25964 8032 26016 8084
rect 26240 8032 26292 8084
rect 22468 7896 22520 7948
rect 22744 7896 22796 7948
rect 22836 7939 22888 7948
rect 22836 7905 22845 7939
rect 22845 7905 22879 7939
rect 22879 7905 22888 7939
rect 23480 8007 23532 8016
rect 23480 7973 23489 8007
rect 23489 7973 23523 8007
rect 23523 7973 23532 8007
rect 23480 7964 23532 7973
rect 22836 7896 22888 7905
rect 23572 7896 23624 7948
rect 15016 7760 15068 7812
rect 19432 7760 19484 7812
rect 4988 7735 5040 7744
rect 4988 7701 4997 7735
rect 4997 7701 5031 7735
rect 5031 7701 5040 7735
rect 4988 7692 5040 7701
rect 5172 7735 5224 7744
rect 5172 7701 5181 7735
rect 5181 7701 5215 7735
rect 5215 7701 5224 7735
rect 5172 7692 5224 7701
rect 11704 7735 11756 7744
rect 11704 7701 11713 7735
rect 11713 7701 11747 7735
rect 11747 7701 11756 7735
rect 11704 7692 11756 7701
rect 12348 7692 12400 7744
rect 14188 7692 14240 7744
rect 15200 7692 15252 7744
rect 15752 7735 15804 7744
rect 15752 7701 15761 7735
rect 15761 7701 15795 7735
rect 15795 7701 15804 7735
rect 15752 7692 15804 7701
rect 16856 7692 16908 7744
rect 20444 7692 20496 7744
rect 22560 7735 22612 7744
rect 22560 7701 22569 7735
rect 22569 7701 22603 7735
rect 22603 7701 22612 7735
rect 22560 7692 22612 7701
rect 24768 7964 24820 8016
rect 24308 7828 24360 7880
rect 25136 7896 25188 7948
rect 25504 7896 25556 7948
rect 25044 7828 25096 7880
rect 24768 7692 24820 7744
rect 25320 7692 25372 7744
rect 3756 7590 3808 7642
rect 3820 7590 3872 7642
rect 3884 7590 3936 7642
rect 3948 7590 4000 7642
rect 4012 7590 4064 7642
rect 10472 7590 10524 7642
rect 10536 7590 10588 7642
rect 10600 7590 10652 7642
rect 10664 7590 10716 7642
rect 10728 7590 10780 7642
rect 17188 7590 17240 7642
rect 17252 7590 17304 7642
rect 17316 7590 17368 7642
rect 17380 7590 17432 7642
rect 17444 7590 17496 7642
rect 23904 7590 23956 7642
rect 23968 7590 24020 7642
rect 24032 7590 24084 7642
rect 24096 7590 24148 7642
rect 24160 7590 24212 7642
rect 2412 7531 2464 7540
rect 2412 7497 2421 7531
rect 2421 7497 2455 7531
rect 2455 7497 2464 7531
rect 2412 7488 2464 7497
rect 3240 7488 3292 7540
rect 4344 7488 4396 7540
rect 3608 7463 3660 7472
rect 3608 7429 3617 7463
rect 3617 7429 3651 7463
rect 3651 7429 3660 7463
rect 3608 7420 3660 7429
rect 4160 7420 4212 7472
rect 1584 7352 1636 7404
rect 4252 7352 4304 7404
rect 5080 7488 5132 7540
rect 5172 7488 5224 7540
rect 6828 7488 6880 7540
rect 11704 7488 11756 7540
rect 4620 7420 4672 7472
rect 1860 7327 1912 7336
rect 1860 7293 1869 7327
rect 1869 7293 1903 7327
rect 1903 7293 1912 7327
rect 1860 7284 1912 7293
rect 2136 7327 2188 7336
rect 2136 7293 2145 7327
rect 2145 7293 2179 7327
rect 2179 7293 2188 7327
rect 2136 7284 2188 7293
rect 1768 7259 1820 7268
rect 1768 7225 1777 7259
rect 1777 7225 1811 7259
rect 1811 7225 1820 7259
rect 1768 7216 1820 7225
rect 2504 7259 2556 7268
rect 2504 7225 2513 7259
rect 2513 7225 2547 7259
rect 2547 7225 2556 7259
rect 2504 7216 2556 7225
rect 3056 7216 3108 7268
rect 3700 7327 3752 7336
rect 3700 7293 3709 7327
rect 3709 7293 3743 7327
rect 3743 7293 3752 7327
rect 3700 7284 3752 7293
rect 4160 7327 4212 7336
rect 4160 7293 4169 7327
rect 4169 7293 4203 7327
rect 4203 7293 4212 7327
rect 4160 7284 4212 7293
rect 4528 7284 4580 7336
rect 7012 7395 7064 7404
rect 7012 7361 7021 7395
rect 7021 7361 7055 7395
rect 7055 7361 7064 7395
rect 7012 7352 7064 7361
rect 8852 7395 8904 7404
rect 8852 7361 8861 7395
rect 8861 7361 8895 7395
rect 8895 7361 8904 7395
rect 8852 7352 8904 7361
rect 6920 7327 6972 7336
rect 6920 7293 6929 7327
rect 6929 7293 6963 7327
rect 6963 7293 6972 7327
rect 6920 7284 6972 7293
rect 8668 7327 8720 7336
rect 8668 7293 8677 7327
rect 8677 7293 8711 7327
rect 8711 7293 8720 7327
rect 8668 7284 8720 7293
rect 10140 7327 10192 7336
rect 10140 7293 10149 7327
rect 10149 7293 10183 7327
rect 10183 7293 10192 7327
rect 10140 7284 10192 7293
rect 7472 7216 7524 7268
rect 9864 7259 9916 7268
rect 9864 7225 9873 7259
rect 9873 7225 9907 7259
rect 9907 7225 9916 7259
rect 9864 7216 9916 7225
rect 1676 7191 1728 7200
rect 1676 7157 1685 7191
rect 1685 7157 1719 7191
rect 1719 7157 1728 7191
rect 1676 7148 1728 7157
rect 4160 7148 4212 7200
rect 4988 7148 5040 7200
rect 5356 7148 5408 7200
rect 8484 7191 8536 7200
rect 8484 7157 8493 7191
rect 8493 7157 8527 7191
rect 8527 7157 8536 7191
rect 8484 7148 8536 7157
rect 9680 7148 9732 7200
rect 10324 7327 10376 7336
rect 10324 7293 10333 7327
rect 10333 7293 10367 7327
rect 10367 7293 10376 7327
rect 10324 7284 10376 7293
rect 10508 7327 10560 7336
rect 10508 7293 10517 7327
rect 10517 7293 10551 7327
rect 10551 7293 10560 7327
rect 12624 7352 12676 7404
rect 10508 7284 10560 7293
rect 12440 7327 12492 7336
rect 12440 7293 12449 7327
rect 12449 7293 12483 7327
rect 12483 7293 12492 7327
rect 12440 7284 12492 7293
rect 12900 7531 12952 7540
rect 12900 7497 12909 7531
rect 12909 7497 12943 7531
rect 12943 7497 12952 7531
rect 12900 7488 12952 7497
rect 13636 7488 13688 7540
rect 14556 7488 14608 7540
rect 15752 7488 15804 7540
rect 16212 7488 16264 7540
rect 17592 7531 17644 7540
rect 17592 7497 17601 7531
rect 17601 7497 17635 7531
rect 17635 7497 17644 7531
rect 17592 7488 17644 7497
rect 18052 7488 18104 7540
rect 11060 7191 11112 7200
rect 11060 7157 11069 7191
rect 11069 7157 11103 7191
rect 11103 7157 11112 7191
rect 11060 7148 11112 7157
rect 12992 7327 13044 7336
rect 12992 7293 13001 7327
rect 13001 7293 13035 7327
rect 13035 7293 13044 7327
rect 12992 7284 13044 7293
rect 14464 7284 14516 7336
rect 19616 7420 19668 7472
rect 23480 7488 23532 7540
rect 25596 7488 25648 7540
rect 24400 7420 24452 7472
rect 19064 7352 19116 7404
rect 24308 7352 24360 7404
rect 25228 7352 25280 7404
rect 25320 7352 25372 7404
rect 17040 7216 17092 7268
rect 19156 7284 19208 7336
rect 19340 7327 19392 7336
rect 19340 7293 19349 7327
rect 19349 7293 19383 7327
rect 19383 7293 19392 7327
rect 19340 7284 19392 7293
rect 19248 7216 19300 7268
rect 21640 7327 21692 7336
rect 21640 7293 21649 7327
rect 21649 7293 21683 7327
rect 21683 7293 21692 7327
rect 21640 7284 21692 7293
rect 23756 7284 23808 7336
rect 22560 7259 22612 7268
rect 22560 7225 22594 7259
rect 22594 7225 22612 7259
rect 22560 7216 22612 7225
rect 25044 7327 25096 7336
rect 25044 7293 25053 7327
rect 25053 7293 25087 7327
rect 25087 7293 25096 7327
rect 25044 7284 25096 7293
rect 25412 7284 25464 7336
rect 20352 7148 20404 7200
rect 25504 7191 25556 7200
rect 25504 7157 25513 7191
rect 25513 7157 25547 7191
rect 25547 7157 25556 7191
rect 25504 7148 25556 7157
rect 7114 7046 7166 7098
rect 7178 7046 7230 7098
rect 7242 7046 7294 7098
rect 7306 7046 7358 7098
rect 7370 7046 7422 7098
rect 13830 7046 13882 7098
rect 13894 7046 13946 7098
rect 13958 7046 14010 7098
rect 14022 7046 14074 7098
rect 14086 7046 14138 7098
rect 20546 7046 20598 7098
rect 20610 7046 20662 7098
rect 20674 7046 20726 7098
rect 20738 7046 20790 7098
rect 20802 7046 20854 7098
rect 27262 7046 27314 7098
rect 27326 7046 27378 7098
rect 27390 7046 27442 7098
rect 27454 7046 27506 7098
rect 27518 7046 27570 7098
rect 1860 6944 1912 6996
rect 2964 6944 3016 6996
rect 2872 6876 2924 6928
rect 1124 6851 1176 6860
rect 1124 6817 1158 6851
rect 1158 6817 1176 6851
rect 1124 6808 1176 6817
rect 2504 6808 2556 6860
rect 3608 6808 3660 6860
rect 4528 6876 4580 6928
rect 5356 6919 5408 6928
rect 5356 6885 5374 6919
rect 5374 6885 5408 6919
rect 5356 6876 5408 6885
rect 7012 6944 7064 6996
rect 7472 6987 7524 6996
rect 7472 6953 7481 6987
rect 7481 6953 7515 6987
rect 7515 6953 7524 6987
rect 7472 6944 7524 6953
rect 10048 6944 10100 6996
rect 10324 6944 10376 6996
rect 11888 6944 11940 6996
rect 12164 6944 12216 6996
rect 10508 6876 10560 6928
rect 11060 6876 11112 6928
rect 2136 6604 2188 6656
rect 2228 6647 2280 6656
rect 2228 6613 2237 6647
rect 2237 6613 2271 6647
rect 2271 6613 2280 6647
rect 2228 6604 2280 6613
rect 3700 6740 3752 6792
rect 4620 6808 4672 6860
rect 6092 6808 6144 6860
rect 6184 6851 6236 6860
rect 6184 6817 6193 6851
rect 6193 6817 6227 6851
rect 6227 6817 6236 6851
rect 6184 6808 6236 6817
rect 6644 6808 6696 6860
rect 6920 6808 6972 6860
rect 4252 6715 4304 6724
rect 4252 6681 4261 6715
rect 4261 6681 4295 6715
rect 4295 6681 4304 6715
rect 4252 6672 4304 6681
rect 8484 6808 8536 6860
rect 8576 6808 8628 6860
rect 9220 6808 9272 6860
rect 10140 6808 10192 6860
rect 10232 6851 10284 6860
rect 10232 6817 10241 6851
rect 10241 6817 10275 6851
rect 10275 6817 10284 6851
rect 10232 6808 10284 6817
rect 9680 6740 9732 6792
rect 6644 6604 6696 6656
rect 7932 6647 7984 6656
rect 7932 6613 7941 6647
rect 7941 6613 7975 6647
rect 7975 6613 7984 6647
rect 7932 6604 7984 6613
rect 8576 6604 8628 6656
rect 11244 6740 11296 6792
rect 11796 6808 11848 6860
rect 12900 6919 12952 6928
rect 12900 6885 12909 6919
rect 12909 6885 12943 6919
rect 12943 6885 12952 6919
rect 12900 6876 12952 6885
rect 12532 6808 12584 6860
rect 12716 6851 12768 6860
rect 12716 6817 12725 6851
rect 12725 6817 12759 6851
rect 12759 6817 12768 6851
rect 12716 6808 12768 6817
rect 14464 6987 14516 6996
rect 14464 6953 14473 6987
rect 14473 6953 14507 6987
rect 14507 6953 14516 6987
rect 14464 6944 14516 6953
rect 15384 6944 15436 6996
rect 22744 6944 22796 6996
rect 16856 6876 16908 6928
rect 19892 6876 19944 6928
rect 20444 6876 20496 6928
rect 15384 6851 15436 6860
rect 15384 6817 15393 6851
rect 15393 6817 15427 6851
rect 15427 6817 15436 6851
rect 15384 6808 15436 6817
rect 16580 6851 16632 6860
rect 16580 6817 16589 6851
rect 16589 6817 16623 6851
rect 16623 6817 16632 6851
rect 16580 6808 16632 6817
rect 18052 6808 18104 6860
rect 19064 6851 19116 6860
rect 19064 6817 19073 6851
rect 19073 6817 19107 6851
rect 19107 6817 19116 6851
rect 19064 6808 19116 6817
rect 19524 6808 19576 6860
rect 19800 6808 19852 6860
rect 10324 6672 10376 6724
rect 12440 6672 12492 6724
rect 12716 6672 12768 6724
rect 11704 6647 11756 6656
rect 11704 6613 11713 6647
rect 11713 6613 11747 6647
rect 11747 6613 11756 6647
rect 11704 6604 11756 6613
rect 12072 6647 12124 6656
rect 12072 6613 12081 6647
rect 12081 6613 12115 6647
rect 12115 6613 12124 6647
rect 12072 6604 12124 6613
rect 15108 6783 15160 6792
rect 15108 6749 15117 6783
rect 15117 6749 15151 6783
rect 15151 6749 15160 6783
rect 15108 6740 15160 6749
rect 17960 6783 18012 6792
rect 17960 6749 17969 6783
rect 17969 6749 18003 6783
rect 18003 6749 18012 6783
rect 17960 6740 18012 6749
rect 21180 6740 21232 6792
rect 21640 6851 21692 6860
rect 21640 6817 21649 6851
rect 21649 6817 21683 6851
rect 21683 6817 21692 6851
rect 21640 6808 21692 6817
rect 21548 6740 21600 6792
rect 25044 6808 25096 6860
rect 24952 6740 25004 6792
rect 14372 6647 14424 6656
rect 14372 6613 14381 6647
rect 14381 6613 14415 6647
rect 14415 6613 14424 6647
rect 14372 6604 14424 6613
rect 14648 6604 14700 6656
rect 15200 6672 15252 6724
rect 18328 6715 18380 6724
rect 18328 6681 18337 6715
rect 18337 6681 18371 6715
rect 18371 6681 18380 6715
rect 18328 6672 18380 6681
rect 21088 6672 21140 6724
rect 23112 6672 23164 6724
rect 15292 6647 15344 6656
rect 15292 6613 15301 6647
rect 15301 6613 15335 6647
rect 15335 6613 15344 6647
rect 15292 6604 15344 6613
rect 16672 6647 16724 6656
rect 16672 6613 16681 6647
rect 16681 6613 16715 6647
rect 16715 6613 16724 6647
rect 16672 6604 16724 6613
rect 18420 6647 18472 6656
rect 18420 6613 18429 6647
rect 18429 6613 18463 6647
rect 18463 6613 18472 6647
rect 18420 6604 18472 6613
rect 19524 6647 19576 6656
rect 19524 6613 19533 6647
rect 19533 6613 19567 6647
rect 19567 6613 19576 6647
rect 19524 6604 19576 6613
rect 19984 6647 20036 6656
rect 19984 6613 19993 6647
rect 19993 6613 20027 6647
rect 20027 6613 20036 6647
rect 19984 6604 20036 6613
rect 24492 6604 24544 6656
rect 25596 6604 25648 6656
rect 25688 6647 25740 6656
rect 25688 6613 25697 6647
rect 25697 6613 25731 6647
rect 25731 6613 25740 6647
rect 25688 6604 25740 6613
rect 25780 6604 25832 6656
rect 3756 6502 3808 6554
rect 3820 6502 3872 6554
rect 3884 6502 3936 6554
rect 3948 6502 4000 6554
rect 4012 6502 4064 6554
rect 10472 6502 10524 6554
rect 10536 6502 10588 6554
rect 10600 6502 10652 6554
rect 10664 6502 10716 6554
rect 10728 6502 10780 6554
rect 17188 6502 17240 6554
rect 17252 6502 17304 6554
rect 17316 6502 17368 6554
rect 17380 6502 17432 6554
rect 17444 6502 17496 6554
rect 23904 6502 23956 6554
rect 23968 6502 24020 6554
rect 24032 6502 24084 6554
rect 24096 6502 24148 6554
rect 24160 6502 24212 6554
rect 1124 6400 1176 6452
rect 1860 6400 1912 6452
rect 2136 6443 2188 6452
rect 2136 6409 2145 6443
rect 2145 6409 2179 6443
rect 2179 6409 2188 6443
rect 2136 6400 2188 6409
rect 2228 6400 2280 6452
rect 2504 6400 2556 6452
rect 3608 6400 3660 6452
rect 4252 6400 4304 6452
rect 6184 6400 6236 6452
rect 6644 6443 6696 6452
rect 6644 6409 6653 6443
rect 6653 6409 6687 6443
rect 6687 6409 6696 6443
rect 6644 6400 6696 6409
rect 6920 6400 6972 6452
rect 8668 6400 8720 6452
rect 9220 6400 9272 6452
rect 10324 6400 10376 6452
rect 11704 6443 11756 6452
rect 11704 6409 11713 6443
rect 11713 6409 11747 6443
rect 11747 6409 11756 6443
rect 11704 6400 11756 6409
rect 12072 6400 12124 6452
rect 12900 6400 12952 6452
rect 14096 6400 14148 6452
rect 14372 6400 14424 6452
rect 14648 6443 14700 6452
rect 14648 6409 14657 6443
rect 14657 6409 14691 6443
rect 14691 6409 14700 6443
rect 14648 6400 14700 6409
rect 15016 6400 15068 6452
rect 15384 6400 15436 6452
rect 17040 6443 17092 6452
rect 17040 6409 17049 6443
rect 17049 6409 17083 6443
rect 17083 6409 17092 6443
rect 17040 6400 17092 6409
rect 18420 6400 18472 6452
rect 19064 6400 19116 6452
rect 19984 6400 20036 6452
rect 1768 6264 1820 6316
rect 1676 6196 1728 6248
rect 2688 6239 2740 6248
rect 2688 6205 2697 6239
rect 2697 6205 2731 6239
rect 2731 6205 2740 6239
rect 2688 6196 2740 6205
rect 3516 6196 3568 6248
rect 8116 6375 8168 6384
rect 4804 6239 4856 6248
rect 4804 6205 4813 6239
rect 4813 6205 4847 6239
rect 4847 6205 4856 6239
rect 4804 6196 4856 6205
rect 5816 6239 5868 6248
rect 5816 6205 5825 6239
rect 5825 6205 5859 6239
rect 5859 6205 5868 6239
rect 5816 6196 5868 6205
rect 6552 6239 6604 6248
rect 6552 6205 6561 6239
rect 6561 6205 6595 6239
rect 6595 6205 6604 6239
rect 6552 6196 6604 6205
rect 6736 6239 6788 6248
rect 6736 6205 6745 6239
rect 6745 6205 6779 6239
rect 6779 6205 6788 6239
rect 6736 6196 6788 6205
rect 8116 6341 8125 6375
rect 8125 6341 8159 6375
rect 8159 6341 8168 6375
rect 8116 6332 8168 6341
rect 8300 6332 8352 6384
rect 7748 6307 7800 6316
rect 7748 6273 7757 6307
rect 7757 6273 7791 6307
rect 7791 6273 7800 6307
rect 7748 6264 7800 6273
rect 2228 6060 2280 6112
rect 11244 6196 11296 6248
rect 11520 6239 11572 6248
rect 11520 6205 11529 6239
rect 11529 6205 11563 6239
rect 11563 6205 11572 6239
rect 11520 6196 11572 6205
rect 11796 6196 11848 6248
rect 11888 6239 11940 6248
rect 11888 6205 11897 6239
rect 11897 6205 11931 6239
rect 11931 6205 11940 6239
rect 11888 6196 11940 6205
rect 8208 6060 8260 6112
rect 10324 6060 10376 6112
rect 11520 6060 11572 6112
rect 11612 6060 11664 6112
rect 12532 6264 12584 6316
rect 12624 6264 12676 6316
rect 13728 6239 13780 6248
rect 13728 6205 13737 6239
rect 13737 6205 13771 6239
rect 13771 6205 13780 6239
rect 13728 6196 13780 6205
rect 15200 6332 15252 6384
rect 12716 6128 12768 6180
rect 15016 6239 15068 6248
rect 15016 6205 15025 6239
rect 15025 6205 15059 6239
rect 15059 6205 15068 6239
rect 15016 6196 15068 6205
rect 16672 6332 16724 6384
rect 20996 6400 21048 6452
rect 22468 6443 22520 6452
rect 22468 6409 22477 6443
rect 22477 6409 22511 6443
rect 22511 6409 22520 6443
rect 22468 6400 22520 6409
rect 23572 6443 23624 6452
rect 23572 6409 23581 6443
rect 23581 6409 23615 6443
rect 23615 6409 23624 6443
rect 23572 6400 23624 6409
rect 24952 6400 25004 6452
rect 25596 6443 25648 6452
rect 25596 6409 25605 6443
rect 25605 6409 25639 6443
rect 25639 6409 25648 6443
rect 25596 6400 25648 6409
rect 25780 6332 25832 6384
rect 23756 6264 23808 6316
rect 14280 6060 14332 6112
rect 14464 6103 14516 6112
rect 14464 6069 14473 6103
rect 14473 6069 14507 6103
rect 14507 6069 14516 6103
rect 14464 6060 14516 6069
rect 17592 6196 17644 6248
rect 18052 6196 18104 6248
rect 19432 6196 19484 6248
rect 17684 6171 17736 6180
rect 17684 6137 17693 6171
rect 17693 6137 17727 6171
rect 17727 6137 17736 6171
rect 17684 6128 17736 6137
rect 19524 6128 19576 6180
rect 21456 6239 21508 6248
rect 21456 6205 21465 6239
rect 21465 6205 21499 6239
rect 21499 6205 21508 6239
rect 21456 6196 21508 6205
rect 22560 6239 22612 6248
rect 22560 6205 22569 6239
rect 22569 6205 22603 6239
rect 22603 6205 22612 6239
rect 22560 6196 22612 6205
rect 22836 6239 22888 6248
rect 22836 6205 22845 6239
rect 22845 6205 22879 6239
rect 22879 6205 22888 6239
rect 22836 6196 22888 6205
rect 23480 6196 23532 6248
rect 24492 6239 24544 6248
rect 24492 6205 24526 6239
rect 24526 6205 24544 6239
rect 24492 6196 24544 6205
rect 26148 6196 26200 6248
rect 25688 6128 25740 6180
rect 15200 6060 15252 6112
rect 15844 6103 15896 6112
rect 15844 6069 15853 6103
rect 15853 6069 15887 6103
rect 15887 6069 15896 6103
rect 15844 6060 15896 6069
rect 18880 6103 18932 6112
rect 18880 6069 18889 6103
rect 18889 6069 18923 6103
rect 18923 6069 18932 6103
rect 18880 6060 18932 6069
rect 20444 6060 20496 6112
rect 21732 6060 21784 6112
rect 7114 5958 7166 6010
rect 7178 5958 7230 6010
rect 7242 5958 7294 6010
rect 7306 5958 7358 6010
rect 7370 5958 7422 6010
rect 13830 5958 13882 6010
rect 13894 5958 13946 6010
rect 13958 5958 14010 6010
rect 14022 5958 14074 6010
rect 14086 5958 14138 6010
rect 20546 5958 20598 6010
rect 20610 5958 20662 6010
rect 20674 5958 20726 6010
rect 20738 5958 20790 6010
rect 20802 5958 20854 6010
rect 27262 5958 27314 6010
rect 27326 5958 27378 6010
rect 27390 5958 27442 6010
rect 27454 5958 27506 6010
rect 27518 5958 27570 6010
rect 2688 5856 2740 5908
rect 3608 5856 3660 5908
rect 4528 5899 4580 5908
rect 4528 5865 4537 5899
rect 4537 5865 4571 5899
rect 4571 5865 4580 5899
rect 4528 5856 4580 5865
rect 4804 5856 4856 5908
rect 5816 5856 5868 5908
rect 6736 5856 6788 5908
rect 7748 5856 7800 5908
rect 8116 5899 8168 5908
rect 8116 5865 8125 5899
rect 8125 5865 8159 5899
rect 8159 5865 8168 5899
rect 8116 5856 8168 5865
rect 9680 5856 9732 5908
rect 2320 5763 2372 5772
rect 2320 5729 2329 5763
rect 2329 5729 2363 5763
rect 2363 5729 2372 5763
rect 2320 5720 2372 5729
rect 2964 5763 3016 5772
rect 2964 5729 2973 5763
rect 2973 5729 3007 5763
rect 3007 5729 3016 5763
rect 2964 5720 3016 5729
rect 5264 5763 5316 5772
rect 5264 5729 5273 5763
rect 5273 5729 5307 5763
rect 5307 5729 5316 5763
rect 5264 5720 5316 5729
rect 6092 5763 6144 5772
rect 6092 5729 6101 5763
rect 6101 5729 6135 5763
rect 6135 5729 6144 5763
rect 6092 5720 6144 5729
rect 7656 5720 7708 5772
rect 7932 5763 7984 5772
rect 7932 5729 7941 5763
rect 7941 5729 7975 5763
rect 7975 5729 7984 5763
rect 7932 5720 7984 5729
rect 9496 5788 9548 5840
rect 14188 5856 14240 5908
rect 11612 5788 11664 5840
rect 13544 5788 13596 5840
rect 13728 5788 13780 5840
rect 15108 5856 15160 5908
rect 15844 5856 15896 5908
rect 17592 5899 17644 5908
rect 17592 5865 17601 5899
rect 17601 5865 17635 5899
rect 17635 5865 17644 5899
rect 17592 5856 17644 5865
rect 17684 5856 17736 5908
rect 2596 5695 2648 5704
rect 2596 5661 2605 5695
rect 2605 5661 2639 5695
rect 2639 5661 2648 5695
rect 2596 5652 2648 5661
rect 8300 5720 8352 5772
rect 9680 5720 9732 5772
rect 10508 5695 10560 5704
rect 10508 5661 10517 5695
rect 10517 5661 10551 5695
rect 10551 5661 10560 5695
rect 10508 5652 10560 5661
rect 1216 5516 1268 5568
rect 2136 5559 2188 5568
rect 2136 5525 2145 5559
rect 2145 5525 2179 5559
rect 2179 5525 2188 5559
rect 2136 5516 2188 5525
rect 3240 5516 3292 5568
rect 6920 5559 6972 5568
rect 6920 5525 6929 5559
rect 6929 5525 6963 5559
rect 6963 5525 6972 5559
rect 6920 5516 6972 5525
rect 9772 5516 9824 5568
rect 10140 5516 10192 5568
rect 11796 5720 11848 5772
rect 11980 5720 12032 5772
rect 12256 5763 12308 5772
rect 12256 5729 12265 5763
rect 12265 5729 12299 5763
rect 12299 5729 12308 5763
rect 12256 5720 12308 5729
rect 12348 5763 12400 5772
rect 12348 5729 12357 5763
rect 12357 5729 12391 5763
rect 12391 5729 12400 5763
rect 12348 5720 12400 5729
rect 12532 5763 12584 5772
rect 12532 5729 12541 5763
rect 12541 5729 12575 5763
rect 12575 5729 12584 5763
rect 12532 5720 12584 5729
rect 12900 5720 12952 5772
rect 12992 5695 13044 5704
rect 12992 5661 13001 5695
rect 13001 5661 13035 5695
rect 13035 5661 13044 5695
rect 12992 5652 13044 5661
rect 16580 5763 16632 5772
rect 16580 5729 16589 5763
rect 16589 5729 16623 5763
rect 16623 5729 16632 5763
rect 16580 5720 16632 5729
rect 16856 5720 16908 5772
rect 18328 5856 18380 5908
rect 18880 5856 18932 5908
rect 21456 5856 21508 5908
rect 22560 5856 22612 5908
rect 22836 5899 22888 5908
rect 22836 5865 22845 5899
rect 22845 5865 22879 5899
rect 22879 5865 22888 5899
rect 22836 5856 22888 5865
rect 17960 5763 18012 5772
rect 17960 5729 17969 5763
rect 17969 5729 18003 5763
rect 18003 5729 18012 5763
rect 17960 5720 18012 5729
rect 18052 5763 18104 5772
rect 18052 5729 18061 5763
rect 18061 5729 18095 5763
rect 18095 5729 18104 5763
rect 18052 5720 18104 5729
rect 18144 5763 18196 5772
rect 18144 5729 18153 5763
rect 18153 5729 18187 5763
rect 18187 5729 18196 5763
rect 18144 5720 18196 5729
rect 15292 5652 15344 5704
rect 14464 5584 14516 5636
rect 15016 5584 15068 5636
rect 18144 5584 18196 5636
rect 23020 5763 23072 5772
rect 23020 5729 23029 5763
rect 23029 5729 23063 5763
rect 23063 5729 23072 5763
rect 23020 5720 23072 5729
rect 23204 5763 23256 5772
rect 23204 5729 23213 5763
rect 23213 5729 23247 5763
rect 23247 5729 23256 5763
rect 23204 5720 23256 5729
rect 24308 5856 24360 5908
rect 25412 5899 25464 5908
rect 25412 5865 25421 5899
rect 25421 5865 25455 5899
rect 25455 5865 25464 5899
rect 25412 5856 25464 5865
rect 25780 5720 25832 5772
rect 23480 5695 23532 5704
rect 23480 5661 23489 5695
rect 23489 5661 23523 5695
rect 23523 5661 23532 5695
rect 23480 5652 23532 5661
rect 25688 5652 25740 5704
rect 26148 5652 26200 5704
rect 24308 5584 24360 5636
rect 11520 5559 11572 5568
rect 11520 5525 11529 5559
rect 11529 5525 11563 5559
rect 11563 5525 11572 5559
rect 11520 5516 11572 5525
rect 12072 5516 12124 5568
rect 12716 5559 12768 5568
rect 12716 5525 12725 5559
rect 12725 5525 12759 5559
rect 12759 5525 12768 5559
rect 12716 5516 12768 5525
rect 14188 5559 14240 5568
rect 14188 5525 14197 5559
rect 14197 5525 14231 5559
rect 14231 5525 14240 5559
rect 14188 5516 14240 5525
rect 15568 5516 15620 5568
rect 20720 5516 20772 5568
rect 21548 5516 21600 5568
rect 3756 5414 3808 5466
rect 3820 5414 3872 5466
rect 3884 5414 3936 5466
rect 3948 5414 4000 5466
rect 4012 5414 4064 5466
rect 10472 5414 10524 5466
rect 10536 5414 10588 5466
rect 10600 5414 10652 5466
rect 10664 5414 10716 5466
rect 10728 5414 10780 5466
rect 17188 5414 17240 5466
rect 17252 5414 17304 5466
rect 17316 5414 17368 5466
rect 17380 5414 17432 5466
rect 17444 5414 17496 5466
rect 23904 5414 23956 5466
rect 23968 5414 24020 5466
rect 24032 5414 24084 5466
rect 24096 5414 24148 5466
rect 24160 5414 24212 5466
rect 2228 5355 2280 5364
rect 2228 5321 2237 5355
rect 2237 5321 2271 5355
rect 2271 5321 2280 5355
rect 2228 5312 2280 5321
rect 2964 5312 3016 5364
rect 5264 5312 5316 5364
rect 6092 5312 6144 5364
rect 6920 5312 6972 5364
rect 7656 5355 7708 5364
rect 7656 5321 7665 5355
rect 7665 5321 7699 5355
rect 7699 5321 7708 5355
rect 7656 5312 7708 5321
rect 11888 5312 11940 5364
rect 11980 5312 12032 5364
rect 11244 5287 11296 5296
rect 11244 5253 11253 5287
rect 11253 5253 11287 5287
rect 11287 5253 11296 5287
rect 11244 5244 11296 5253
rect 12900 5312 12952 5364
rect 12992 5355 13044 5364
rect 12992 5321 13001 5355
rect 13001 5321 13035 5355
rect 13035 5321 13044 5355
rect 12992 5312 13044 5321
rect 15200 5355 15252 5364
rect 15200 5321 15209 5355
rect 15209 5321 15243 5355
rect 15243 5321 15252 5355
rect 15200 5312 15252 5321
rect 16580 5355 16632 5364
rect 16580 5321 16589 5355
rect 16589 5321 16623 5355
rect 16623 5321 16632 5355
rect 16580 5312 16632 5321
rect 18696 5244 18748 5296
rect 8852 5176 8904 5228
rect 14188 5219 14240 5228
rect 14188 5185 14197 5219
rect 14197 5185 14231 5219
rect 14231 5185 14240 5219
rect 14188 5176 14240 5185
rect 1124 5151 1176 5160
rect 1124 5117 1133 5151
rect 1133 5117 1167 5151
rect 1167 5117 1176 5151
rect 1124 5108 1176 5117
rect 1216 5151 1268 5160
rect 1216 5117 1225 5151
rect 1225 5117 1259 5151
rect 1259 5117 1268 5151
rect 1216 5108 1268 5117
rect 2136 5108 2188 5160
rect 3332 5108 3384 5160
rect 5080 5108 5132 5160
rect 5724 5151 5776 5160
rect 5724 5117 5733 5151
rect 5733 5117 5767 5151
rect 5767 5117 5776 5151
rect 5724 5108 5776 5117
rect 6368 5151 6420 5160
rect 6368 5117 6377 5151
rect 6377 5117 6411 5151
rect 6411 5117 6420 5151
rect 6368 5108 6420 5117
rect 3424 4972 3476 5024
rect 8576 5151 8628 5160
rect 8576 5117 8585 5151
rect 8585 5117 8619 5151
rect 8619 5117 8628 5151
rect 8576 5108 8628 5117
rect 8484 4972 8536 5024
rect 8760 5015 8812 5024
rect 8760 4981 8769 5015
rect 8769 4981 8803 5015
rect 8803 4981 8812 5015
rect 8760 4972 8812 4981
rect 9588 4972 9640 5024
rect 10232 5108 10284 5160
rect 10784 5151 10836 5160
rect 10784 5117 10793 5151
rect 10793 5117 10827 5151
rect 10827 5117 10836 5151
rect 10784 5108 10836 5117
rect 11520 5040 11572 5092
rect 12072 5108 12124 5160
rect 12164 5040 12216 5092
rect 12716 5151 12768 5160
rect 12716 5117 12725 5151
rect 12725 5117 12759 5151
rect 12759 5117 12768 5151
rect 12716 5108 12768 5117
rect 13084 5108 13136 5160
rect 14464 5151 14516 5160
rect 14464 5117 14473 5151
rect 14473 5117 14507 5151
rect 14507 5117 14516 5151
rect 14464 5108 14516 5117
rect 15292 5151 15344 5160
rect 15292 5117 15301 5151
rect 15301 5117 15335 5151
rect 15335 5117 15344 5151
rect 15292 5108 15344 5117
rect 15568 5151 15620 5160
rect 15568 5117 15577 5151
rect 15577 5117 15611 5151
rect 15611 5117 15620 5151
rect 15568 5108 15620 5117
rect 19984 5312 20036 5364
rect 20720 5312 20772 5364
rect 21732 5312 21784 5364
rect 23204 5312 23256 5364
rect 23756 5312 23808 5364
rect 24492 5312 24544 5364
rect 26332 5312 26384 5364
rect 21548 5287 21600 5296
rect 21548 5253 21557 5287
rect 21557 5253 21591 5287
rect 21591 5253 21600 5287
rect 21548 5244 21600 5253
rect 25780 5244 25832 5296
rect 19800 5151 19852 5160
rect 19800 5117 19809 5151
rect 19809 5117 19843 5151
rect 19843 5117 19852 5151
rect 19800 5108 19852 5117
rect 20352 5108 20404 5160
rect 20720 5151 20772 5160
rect 20720 5117 20729 5151
rect 20729 5117 20763 5151
rect 20763 5117 20772 5151
rect 20720 5108 20772 5117
rect 21180 5219 21232 5228
rect 21180 5185 21189 5219
rect 21189 5185 21223 5219
rect 21223 5185 21232 5219
rect 21180 5176 21232 5185
rect 21456 5108 21508 5160
rect 22744 5151 22796 5160
rect 22744 5117 22753 5151
rect 22753 5117 22787 5151
rect 22787 5117 22796 5151
rect 22744 5108 22796 5117
rect 22928 5151 22980 5160
rect 22928 5117 22937 5151
rect 22937 5117 22971 5151
rect 22971 5117 22980 5151
rect 22928 5108 22980 5117
rect 23756 5108 23808 5160
rect 24584 5151 24636 5160
rect 24584 5117 24593 5151
rect 24593 5117 24627 5151
rect 24627 5117 24636 5151
rect 24584 5108 24636 5117
rect 25596 5108 25648 5160
rect 26056 5108 26108 5160
rect 11336 4972 11388 5024
rect 11888 4972 11940 5024
rect 12072 4972 12124 5024
rect 20076 5015 20128 5024
rect 20076 4981 20085 5015
rect 20085 4981 20119 5015
rect 20119 4981 20128 5015
rect 20076 4972 20128 4981
rect 20168 4972 20220 5024
rect 20904 5040 20956 5092
rect 21088 5040 21140 5092
rect 20720 4972 20772 5024
rect 22100 5015 22152 5024
rect 22100 4981 22109 5015
rect 22109 4981 22143 5015
rect 22143 4981 22152 5015
rect 22100 4972 22152 4981
rect 22192 4972 22244 5024
rect 26792 5015 26844 5024
rect 26792 4981 26801 5015
rect 26801 4981 26835 5015
rect 26835 4981 26844 5015
rect 26792 4972 26844 4981
rect 7114 4870 7166 4922
rect 7178 4870 7230 4922
rect 7242 4870 7294 4922
rect 7306 4870 7358 4922
rect 7370 4870 7422 4922
rect 13830 4870 13882 4922
rect 13894 4870 13946 4922
rect 13958 4870 14010 4922
rect 14022 4870 14074 4922
rect 14086 4870 14138 4922
rect 20546 4870 20598 4922
rect 20610 4870 20662 4922
rect 20674 4870 20726 4922
rect 20738 4870 20790 4922
rect 20802 4870 20854 4922
rect 27262 4870 27314 4922
rect 27326 4870 27378 4922
rect 27390 4870 27442 4922
rect 27454 4870 27506 4922
rect 27518 4870 27570 4922
rect 1124 4768 1176 4820
rect 1952 4768 2004 4820
rect 5724 4768 5776 4820
rect 8208 4811 8260 4820
rect 8208 4777 8217 4811
rect 8217 4777 8251 4811
rect 8251 4777 8260 4811
rect 8208 4768 8260 4777
rect 8760 4768 8812 4820
rect 9772 4811 9824 4820
rect 9772 4777 9781 4811
rect 9781 4777 9815 4811
rect 9815 4777 9824 4811
rect 9772 4768 9824 4777
rect 10784 4768 10836 4820
rect 12256 4768 12308 4820
rect 2596 4700 2648 4752
rect 2136 4632 2188 4684
rect 3056 4632 3108 4684
rect 2596 4564 2648 4616
rect 3332 4632 3384 4684
rect 4160 4700 4212 4752
rect 3516 4675 3568 4684
rect 3516 4641 3525 4675
rect 3525 4641 3559 4675
rect 3559 4641 3568 4675
rect 3516 4632 3568 4641
rect 4344 4632 4396 4684
rect 4252 4564 4304 4616
rect 4804 4632 4856 4684
rect 5540 4632 5592 4684
rect 8300 4700 8352 4752
rect 8576 4700 8628 4752
rect 9036 4700 9088 4752
rect 9588 4700 9640 4752
rect 10692 4700 10744 4752
rect 6000 4564 6052 4616
rect 8024 4564 8076 4616
rect 8852 4675 8904 4684
rect 8852 4641 8861 4675
rect 8861 4641 8895 4675
rect 8895 4641 8904 4675
rect 8852 4632 8904 4641
rect 3424 4539 3476 4548
rect 3424 4505 3433 4539
rect 3433 4505 3467 4539
rect 3467 4505 3476 4539
rect 3424 4496 3476 4505
rect 4436 4539 4488 4548
rect 4436 4505 4445 4539
rect 4445 4505 4479 4539
rect 4479 4505 4488 4539
rect 4436 4496 4488 4505
rect 5448 4428 5500 4480
rect 8484 4496 8536 4548
rect 11244 4632 11296 4684
rect 11796 4632 11848 4684
rect 12072 4743 12124 4752
rect 12072 4709 12081 4743
rect 12081 4709 12115 4743
rect 12115 4709 12124 4743
rect 14464 4768 14516 4820
rect 15292 4768 15344 4820
rect 18052 4768 18104 4820
rect 21456 4811 21508 4820
rect 21456 4777 21481 4811
rect 21481 4777 21508 4811
rect 21456 4768 21508 4777
rect 22100 4768 22152 4820
rect 12072 4700 12124 4709
rect 12072 4564 12124 4616
rect 12532 4632 12584 4684
rect 13452 4675 13504 4684
rect 12808 4564 12860 4616
rect 13452 4641 13461 4675
rect 13461 4641 13495 4675
rect 13495 4641 13504 4675
rect 13452 4632 13504 4641
rect 14188 4675 14240 4684
rect 14188 4641 14197 4675
rect 14197 4641 14231 4675
rect 14231 4641 14240 4675
rect 14188 4632 14240 4641
rect 14740 4675 14792 4684
rect 14740 4641 14749 4675
rect 14749 4641 14783 4675
rect 14783 4641 14792 4675
rect 14740 4632 14792 4641
rect 14924 4675 14976 4684
rect 14924 4641 14933 4675
rect 14933 4641 14967 4675
rect 14967 4641 14976 4675
rect 14924 4632 14976 4641
rect 16580 4675 16632 4684
rect 16580 4641 16589 4675
rect 16589 4641 16623 4675
rect 16623 4641 16632 4675
rect 16580 4632 16632 4641
rect 17592 4632 17644 4684
rect 17684 4675 17736 4684
rect 17684 4641 17693 4675
rect 17693 4641 17727 4675
rect 17727 4641 17736 4675
rect 17684 4632 17736 4641
rect 19340 4675 19392 4684
rect 19340 4641 19358 4675
rect 19358 4641 19392 4675
rect 19340 4632 19392 4641
rect 19708 4632 19760 4684
rect 20076 4700 20128 4752
rect 21180 4700 21232 4752
rect 7012 4428 7064 4480
rect 9128 4471 9180 4480
rect 9128 4437 9137 4471
rect 9137 4437 9171 4471
rect 9171 4437 9180 4471
rect 9128 4428 9180 4437
rect 9680 4428 9732 4480
rect 10968 4471 11020 4480
rect 10968 4437 10977 4471
rect 10977 4437 11011 4471
rect 11011 4437 11020 4471
rect 10968 4428 11020 4437
rect 13084 4539 13136 4548
rect 13084 4505 13093 4539
rect 13093 4505 13127 4539
rect 13127 4505 13136 4539
rect 13084 4496 13136 4505
rect 12808 4428 12860 4480
rect 13176 4428 13228 4480
rect 14280 4428 14332 4480
rect 17868 4564 17920 4616
rect 18144 4496 18196 4548
rect 18236 4471 18288 4480
rect 18236 4437 18245 4471
rect 18245 4437 18279 4471
rect 18279 4437 18288 4471
rect 18236 4428 18288 4437
rect 19432 4428 19484 4480
rect 20444 4496 20496 4548
rect 22560 4564 22612 4616
rect 21364 4428 21416 4480
rect 23388 4632 23440 4684
rect 25044 4811 25096 4820
rect 25044 4777 25053 4811
rect 25053 4777 25087 4811
rect 25087 4777 25096 4811
rect 25044 4768 25096 4777
rect 25780 4768 25832 4820
rect 26148 4811 26200 4820
rect 26148 4777 26157 4811
rect 26157 4777 26191 4811
rect 26191 4777 26200 4811
rect 26148 4768 26200 4777
rect 26424 4743 26476 4752
rect 26424 4709 26433 4743
rect 26433 4709 26467 4743
rect 26467 4709 26476 4743
rect 26424 4700 26476 4709
rect 25596 4632 25648 4684
rect 25780 4632 25832 4684
rect 22284 4428 22336 4480
rect 22468 4471 22520 4480
rect 22468 4437 22477 4471
rect 22477 4437 22511 4471
rect 22511 4437 22520 4471
rect 22468 4428 22520 4437
rect 23112 4471 23164 4480
rect 23112 4437 23121 4471
rect 23121 4437 23155 4471
rect 23155 4437 23164 4471
rect 23112 4428 23164 4437
rect 25504 4496 25556 4548
rect 26056 4632 26108 4684
rect 26792 4564 26844 4616
rect 24308 4428 24360 4480
rect 26884 4471 26936 4480
rect 26884 4437 26893 4471
rect 26893 4437 26927 4471
rect 26927 4437 26936 4471
rect 26884 4428 26936 4437
rect 3756 4326 3808 4378
rect 3820 4326 3872 4378
rect 3884 4326 3936 4378
rect 3948 4326 4000 4378
rect 4012 4326 4064 4378
rect 10472 4326 10524 4378
rect 10536 4326 10588 4378
rect 10600 4326 10652 4378
rect 10664 4326 10716 4378
rect 10728 4326 10780 4378
rect 17188 4326 17240 4378
rect 17252 4326 17304 4378
rect 17316 4326 17368 4378
rect 17380 4326 17432 4378
rect 17444 4326 17496 4378
rect 23904 4326 23956 4378
rect 23968 4326 24020 4378
rect 24032 4326 24084 4378
rect 24096 4326 24148 4378
rect 24160 4326 24212 4378
rect 3056 4156 3108 4208
rect 3424 4156 3476 4208
rect 4252 4224 4304 4276
rect 4436 4267 4488 4276
rect 4436 4233 4445 4267
rect 4445 4233 4479 4267
rect 4479 4233 4488 4267
rect 4436 4224 4488 4233
rect 4896 4224 4948 4276
rect 3332 4088 3384 4140
rect 4988 4156 5040 4208
rect 6368 4224 6420 4276
rect 8024 4267 8076 4276
rect 8024 4233 8033 4267
rect 8033 4233 8067 4267
rect 8067 4233 8076 4267
rect 8024 4224 8076 4233
rect 8484 4224 8536 4276
rect 9128 4224 9180 4276
rect 13084 4267 13136 4276
rect 13084 4233 13093 4267
rect 13093 4233 13127 4267
rect 13127 4233 13136 4267
rect 13084 4224 13136 4233
rect 17684 4224 17736 4276
rect 19340 4267 19392 4276
rect 19340 4233 19349 4267
rect 19349 4233 19383 4267
rect 19383 4233 19392 4267
rect 19340 4224 19392 4233
rect 6460 4156 6512 4208
rect 10876 4156 10928 4208
rect 15016 4156 15068 4208
rect 18236 4156 18288 4208
rect 2228 4020 2280 4072
rect 2596 4063 2648 4072
rect 2596 4029 2605 4063
rect 2605 4029 2639 4063
rect 2639 4029 2648 4063
rect 2596 4020 2648 4029
rect 3516 4020 3568 4072
rect 4160 4063 4212 4072
rect 4160 4029 4169 4063
rect 4169 4029 4203 4063
rect 4203 4029 4212 4063
rect 4160 4020 4212 4029
rect 4804 4063 4856 4072
rect 4804 4029 4813 4063
rect 4813 4029 4847 4063
rect 4847 4029 4856 4063
rect 4804 4020 4856 4029
rect 4896 4020 4948 4072
rect 10968 4088 11020 4140
rect 5448 4020 5500 4072
rect 5816 4020 5868 4072
rect 2320 3952 2372 4004
rect 2780 3995 2832 4004
rect 2780 3961 2789 3995
rect 2789 3961 2823 3995
rect 2823 3961 2832 3995
rect 2780 3952 2832 3961
rect 4068 3952 4120 4004
rect 4252 3995 4304 4004
rect 4252 3961 4261 3995
rect 4261 3961 4295 3995
rect 4295 3961 4304 3995
rect 4252 3952 4304 3961
rect 4344 3952 4396 4004
rect 6736 4063 6788 4072
rect 6736 4029 6745 4063
rect 6745 4029 6779 4063
rect 6779 4029 6788 4063
rect 6736 4020 6788 4029
rect 7012 4063 7064 4072
rect 7012 4029 7021 4063
rect 7021 4029 7055 4063
rect 7055 4029 7064 4063
rect 7012 4020 7064 4029
rect 2136 3927 2188 3936
rect 2136 3893 2145 3927
rect 2145 3893 2179 3927
rect 2179 3893 2188 3927
rect 6184 3952 6236 4004
rect 8576 4063 8628 4072
rect 8576 4029 8585 4063
rect 8585 4029 8619 4063
rect 8619 4029 8628 4063
rect 8576 4020 8628 4029
rect 8852 4020 8904 4072
rect 9128 4020 9180 4072
rect 9680 4020 9732 4072
rect 2136 3884 2188 3893
rect 4896 3927 4948 3936
rect 4896 3893 4905 3927
rect 4905 3893 4939 3927
rect 4939 3893 4948 3927
rect 4896 3884 4948 3893
rect 5264 3927 5316 3936
rect 5264 3893 5273 3927
rect 5273 3893 5307 3927
rect 5307 3893 5316 3927
rect 5264 3884 5316 3893
rect 5448 3927 5500 3936
rect 5448 3893 5457 3927
rect 5457 3893 5491 3927
rect 5491 3893 5500 3927
rect 5448 3884 5500 3893
rect 6000 3884 6052 3936
rect 6644 3884 6696 3936
rect 9956 3952 10008 4004
rect 10324 3952 10376 4004
rect 10600 4063 10652 4072
rect 10600 4029 10609 4063
rect 10609 4029 10643 4063
rect 10643 4029 10652 4063
rect 10600 4020 10652 4029
rect 11796 4020 11848 4072
rect 12072 4020 12124 4072
rect 13360 4020 13412 4072
rect 13452 4020 13504 4072
rect 13176 3952 13228 4004
rect 15292 4063 15344 4072
rect 15292 4029 15301 4063
rect 15301 4029 15335 4063
rect 15335 4029 15344 4063
rect 15292 4020 15344 4029
rect 15568 4063 15620 4072
rect 15568 4029 15577 4063
rect 15577 4029 15611 4063
rect 15611 4029 15620 4063
rect 15568 4020 15620 4029
rect 16580 4020 16632 4072
rect 21180 4156 21232 4208
rect 8300 3884 8352 3936
rect 11060 3884 11112 3936
rect 12992 3884 13044 3936
rect 13636 3927 13688 3936
rect 13636 3893 13645 3927
rect 13645 3893 13679 3927
rect 13679 3893 13688 3927
rect 13636 3884 13688 3893
rect 15384 3884 15436 3936
rect 17868 4020 17920 4072
rect 22560 4224 22612 4276
rect 22928 4267 22980 4276
rect 22928 4233 22937 4267
rect 22937 4233 22971 4267
rect 22971 4233 22980 4267
rect 22928 4224 22980 4233
rect 23204 4267 23256 4276
rect 23204 4233 23213 4267
rect 23213 4233 23247 4267
rect 23247 4233 23256 4267
rect 23204 4224 23256 4233
rect 25504 4224 25556 4276
rect 26332 4224 26384 4276
rect 21364 4156 21416 4208
rect 17592 3952 17644 4004
rect 18696 3995 18748 4004
rect 18696 3961 18705 3995
rect 18705 3961 18739 3995
rect 18739 3961 18748 3995
rect 18696 3952 18748 3961
rect 17868 3884 17920 3936
rect 18052 3884 18104 3936
rect 19984 4020 20036 4072
rect 20260 4020 20312 4072
rect 20904 4063 20956 4072
rect 20904 4029 20913 4063
rect 20913 4029 20947 4063
rect 20947 4029 20956 4063
rect 20904 4020 20956 4029
rect 21180 4020 21232 4072
rect 19800 3927 19852 3936
rect 19800 3893 19809 3927
rect 19809 3893 19843 3927
rect 19843 3893 19852 3927
rect 19800 3884 19852 3893
rect 21180 3884 21232 3936
rect 21456 3884 21508 3936
rect 21824 4063 21876 4072
rect 21824 4029 21833 4063
rect 21833 4029 21867 4063
rect 21867 4029 21876 4063
rect 21824 4020 21876 4029
rect 22284 4156 22336 4208
rect 22652 4156 22704 4208
rect 23756 4088 23808 4140
rect 22008 3952 22060 4004
rect 22560 4020 22612 4072
rect 22652 4020 22704 4072
rect 23296 4063 23348 4072
rect 23296 4029 23305 4063
rect 23305 4029 23339 4063
rect 23339 4029 23348 4063
rect 23296 4020 23348 4029
rect 24216 4063 24268 4072
rect 24216 4029 24225 4063
rect 24225 4029 24259 4063
rect 24259 4029 24268 4063
rect 24216 4020 24268 4029
rect 26884 3952 26936 4004
rect 21824 3884 21876 3936
rect 22560 3927 22612 3936
rect 22560 3893 22569 3927
rect 22569 3893 22603 3927
rect 22603 3893 22612 3927
rect 22560 3884 22612 3893
rect 23480 3927 23532 3936
rect 23480 3893 23489 3927
rect 23489 3893 23523 3927
rect 23523 3893 23532 3927
rect 23480 3884 23532 3893
rect 24952 3927 25004 3936
rect 24952 3893 24961 3927
rect 24961 3893 24995 3927
rect 24995 3893 25004 3927
rect 24952 3884 25004 3893
rect 25688 3927 25740 3936
rect 25688 3893 25697 3927
rect 25697 3893 25731 3927
rect 25731 3893 25740 3927
rect 25688 3884 25740 3893
rect 7114 3782 7166 3834
rect 7178 3782 7230 3834
rect 7242 3782 7294 3834
rect 7306 3782 7358 3834
rect 7370 3782 7422 3834
rect 13830 3782 13882 3834
rect 13894 3782 13946 3834
rect 13958 3782 14010 3834
rect 14022 3782 14074 3834
rect 14086 3782 14138 3834
rect 20546 3782 20598 3834
rect 20610 3782 20662 3834
rect 20674 3782 20726 3834
rect 20738 3782 20790 3834
rect 20802 3782 20854 3834
rect 27262 3782 27314 3834
rect 27326 3782 27378 3834
rect 27390 3782 27442 3834
rect 27454 3782 27506 3834
rect 27518 3782 27570 3834
rect 2044 3408 2096 3460
rect 2964 3680 3016 3732
rect 3056 3723 3108 3732
rect 3056 3689 3065 3723
rect 3065 3689 3099 3723
rect 3099 3689 3108 3723
rect 3056 3680 3108 3689
rect 5080 3723 5132 3732
rect 5080 3689 5089 3723
rect 5089 3689 5123 3723
rect 5123 3689 5132 3723
rect 5080 3680 5132 3689
rect 6736 3680 6788 3732
rect 9772 3680 9824 3732
rect 10784 3680 10836 3732
rect 12072 3680 12124 3732
rect 12808 3680 12860 3732
rect 12992 3680 13044 3732
rect 13728 3680 13780 3732
rect 14924 3723 14976 3732
rect 14924 3689 14933 3723
rect 14933 3689 14967 3723
rect 14967 3689 14976 3723
rect 14924 3680 14976 3689
rect 3332 3587 3384 3596
rect 3332 3553 3341 3587
rect 3341 3553 3375 3587
rect 3375 3553 3384 3587
rect 3332 3544 3384 3553
rect 3424 3587 3476 3596
rect 3424 3553 3434 3587
rect 3434 3553 3468 3587
rect 3468 3553 3476 3587
rect 3424 3544 3476 3553
rect 3240 3408 3292 3460
rect 4160 3544 4212 3596
rect 4344 3587 4396 3596
rect 4344 3553 4353 3587
rect 4353 3553 4387 3587
rect 4387 3553 4396 3587
rect 4344 3544 4396 3553
rect 4528 3587 4580 3596
rect 4528 3553 4537 3587
rect 4537 3553 4571 3587
rect 4571 3553 4580 3587
rect 4528 3544 4580 3553
rect 4712 3587 4764 3596
rect 4712 3553 4721 3587
rect 4721 3553 4755 3587
rect 4755 3553 4764 3587
rect 4712 3544 4764 3553
rect 4436 3476 4488 3528
rect 5816 3476 5868 3528
rect 6276 3476 6328 3528
rect 6644 3587 6696 3596
rect 6644 3553 6653 3587
rect 6653 3553 6687 3587
rect 6687 3553 6696 3587
rect 6644 3544 6696 3553
rect 6828 3544 6880 3596
rect 8576 3544 8628 3596
rect 8208 3476 8260 3528
rect 10232 3544 10284 3596
rect 10600 3587 10652 3596
rect 10600 3553 10609 3587
rect 10609 3553 10643 3587
rect 10643 3553 10652 3587
rect 10600 3544 10652 3553
rect 11336 3476 11388 3528
rect 12532 3544 12584 3596
rect 13268 3655 13320 3664
rect 13268 3621 13277 3655
rect 13277 3621 13311 3655
rect 13311 3621 13320 3655
rect 13268 3612 13320 3621
rect 13544 3612 13596 3664
rect 15292 3680 15344 3732
rect 17684 3680 17736 3732
rect 18052 3723 18104 3732
rect 18052 3689 18061 3723
rect 18061 3689 18095 3723
rect 18095 3689 18104 3723
rect 18052 3680 18104 3689
rect 19340 3680 19392 3732
rect 19708 3680 19760 3732
rect 19800 3680 19852 3732
rect 21824 3680 21876 3732
rect 21916 3680 21968 3732
rect 22560 3680 22612 3732
rect 22928 3680 22980 3732
rect 23296 3680 23348 3732
rect 23480 3680 23532 3732
rect 24216 3680 24268 3732
rect 24952 3680 25004 3732
rect 25688 3680 25740 3732
rect 13176 3587 13228 3596
rect 13176 3553 13185 3587
rect 13185 3553 13219 3587
rect 13219 3553 13228 3587
rect 13176 3544 13228 3553
rect 13360 3587 13412 3596
rect 13360 3553 13369 3587
rect 13369 3553 13403 3587
rect 13403 3553 13412 3587
rect 13360 3544 13412 3553
rect 4436 3340 4488 3392
rect 6368 3383 6420 3392
rect 6368 3349 6377 3383
rect 6377 3349 6411 3383
rect 6411 3349 6420 3383
rect 6368 3340 6420 3349
rect 6460 3340 6512 3392
rect 6920 3340 6972 3392
rect 7380 3340 7432 3392
rect 7472 3383 7524 3392
rect 7472 3349 7481 3383
rect 7481 3349 7515 3383
rect 7515 3349 7524 3383
rect 7472 3340 7524 3349
rect 8852 3340 8904 3392
rect 9128 3340 9180 3392
rect 11428 3383 11480 3392
rect 11428 3349 11437 3383
rect 11437 3349 11471 3383
rect 11471 3349 11480 3383
rect 11428 3340 11480 3349
rect 11796 3408 11848 3460
rect 12808 3476 12860 3528
rect 13912 3476 13964 3528
rect 14372 3544 14424 3596
rect 14556 3587 14608 3596
rect 14556 3553 14565 3587
rect 14565 3553 14599 3587
rect 14599 3553 14608 3587
rect 14556 3544 14608 3553
rect 14280 3476 14332 3528
rect 14832 3544 14884 3596
rect 14924 3476 14976 3528
rect 15384 3544 15436 3596
rect 15660 3544 15712 3596
rect 15752 3587 15804 3596
rect 15752 3553 15761 3587
rect 15761 3553 15795 3587
rect 15795 3553 15804 3587
rect 15752 3544 15804 3553
rect 17868 3587 17920 3596
rect 17868 3553 17877 3587
rect 17877 3553 17911 3587
rect 17911 3553 17920 3587
rect 17868 3544 17920 3553
rect 17592 3476 17644 3528
rect 20168 3544 20220 3596
rect 21272 3544 21324 3596
rect 21456 3544 21508 3596
rect 21088 3476 21140 3528
rect 22100 3587 22152 3596
rect 22100 3553 22109 3587
rect 22109 3553 22143 3587
rect 22143 3553 22152 3587
rect 22100 3544 22152 3553
rect 22468 3544 22520 3596
rect 22744 3544 22796 3596
rect 21732 3476 21784 3528
rect 12256 3383 12308 3392
rect 12256 3349 12265 3383
rect 12265 3349 12299 3383
rect 12299 3349 12308 3383
rect 12256 3340 12308 3349
rect 14372 3408 14424 3460
rect 19524 3408 19576 3460
rect 23020 3476 23072 3528
rect 14464 3340 14516 3392
rect 15108 3383 15160 3392
rect 15108 3349 15117 3383
rect 15117 3349 15151 3383
rect 15151 3349 15160 3383
rect 15108 3340 15160 3349
rect 15476 3340 15528 3392
rect 16488 3383 16540 3392
rect 16488 3349 16497 3383
rect 16497 3349 16531 3383
rect 16531 3349 16540 3383
rect 16488 3340 16540 3349
rect 17040 3340 17092 3392
rect 17684 3340 17736 3392
rect 19432 3340 19484 3392
rect 19708 3340 19760 3392
rect 21456 3383 21508 3392
rect 21456 3349 21465 3383
rect 21465 3349 21499 3383
rect 21499 3349 21508 3383
rect 21456 3340 21508 3349
rect 21824 3340 21876 3392
rect 22008 3340 22060 3392
rect 24308 3408 24360 3460
rect 25780 3476 25832 3528
rect 25688 3408 25740 3460
rect 26424 3408 26476 3460
rect 23112 3383 23164 3392
rect 23112 3349 23121 3383
rect 23121 3349 23155 3383
rect 23155 3349 23164 3383
rect 23112 3340 23164 3349
rect 23756 3340 23808 3392
rect 24584 3340 24636 3392
rect 3756 3238 3808 3290
rect 3820 3238 3872 3290
rect 3884 3238 3936 3290
rect 3948 3238 4000 3290
rect 4012 3238 4064 3290
rect 10472 3238 10524 3290
rect 10536 3238 10588 3290
rect 10600 3238 10652 3290
rect 10664 3238 10716 3290
rect 10728 3238 10780 3290
rect 17188 3238 17240 3290
rect 17252 3238 17304 3290
rect 17316 3238 17368 3290
rect 17380 3238 17432 3290
rect 17444 3238 17496 3290
rect 23904 3238 23956 3290
rect 23968 3238 24020 3290
rect 24032 3238 24084 3290
rect 24096 3238 24148 3290
rect 24160 3238 24212 3290
rect 2228 3136 2280 3188
rect 6276 3136 6328 3188
rect 2044 2932 2096 2984
rect 2780 3000 2832 3052
rect 1308 2796 1360 2848
rect 2044 2839 2096 2848
rect 2044 2805 2053 2839
rect 2053 2805 2087 2839
rect 2087 2805 2096 2839
rect 2044 2796 2096 2805
rect 2412 2975 2464 2984
rect 2412 2941 2421 2975
rect 2421 2941 2455 2975
rect 2455 2941 2464 2975
rect 2412 2932 2464 2941
rect 3056 3000 3108 3052
rect 5264 3068 5316 3120
rect 7012 3136 7064 3188
rect 6920 3068 6972 3120
rect 3792 3043 3844 3052
rect 3792 3009 3801 3043
rect 3801 3009 3835 3043
rect 3835 3009 3844 3043
rect 7472 3136 7524 3188
rect 8208 3179 8260 3188
rect 8208 3145 8217 3179
rect 8217 3145 8251 3179
rect 8251 3145 8260 3179
rect 8208 3136 8260 3145
rect 8576 3179 8628 3188
rect 8576 3145 8585 3179
rect 8585 3145 8619 3179
rect 8619 3145 8628 3179
rect 8576 3136 8628 3145
rect 10232 3136 10284 3188
rect 3792 3000 3844 3009
rect 3240 2932 3292 2984
rect 2504 2864 2556 2916
rect 4344 2864 4396 2916
rect 5264 2864 5316 2916
rect 6644 2975 6696 2984
rect 6644 2941 6653 2975
rect 6653 2941 6687 2975
rect 6687 2941 6696 2975
rect 6644 2932 6696 2941
rect 9956 3043 10008 3052
rect 9956 3009 9965 3043
rect 9965 3009 9999 3043
rect 9999 3009 10008 3043
rect 9956 3000 10008 3009
rect 2688 2796 2740 2848
rect 4252 2796 4304 2848
rect 7380 2932 7432 2984
rect 10692 3111 10744 3120
rect 10692 3077 10701 3111
rect 10701 3077 10735 3111
rect 10735 3077 10744 3111
rect 10692 3068 10744 3077
rect 11888 3179 11940 3188
rect 11888 3145 11897 3179
rect 11897 3145 11931 3179
rect 11931 3145 11940 3179
rect 11888 3136 11940 3145
rect 12900 3068 12952 3120
rect 13820 3179 13872 3188
rect 13820 3145 13829 3179
rect 13829 3145 13863 3179
rect 13863 3145 13872 3179
rect 13820 3136 13872 3145
rect 14188 3179 14240 3188
rect 14188 3145 14197 3179
rect 14197 3145 14231 3179
rect 14231 3145 14240 3179
rect 14188 3136 14240 3145
rect 15108 3136 15160 3188
rect 15476 3179 15528 3188
rect 15476 3145 15485 3179
rect 15485 3145 15519 3179
rect 15519 3145 15528 3179
rect 15476 3136 15528 3145
rect 15568 3136 15620 3188
rect 14096 3068 14148 3120
rect 14372 3068 14424 3120
rect 7196 2864 7248 2916
rect 9680 2907 9732 2916
rect 9680 2873 9698 2907
rect 9698 2873 9732 2907
rect 9680 2864 9732 2873
rect 10784 2975 10836 2984
rect 10784 2941 10793 2975
rect 10793 2941 10827 2975
rect 10827 2941 10836 2975
rect 10784 2932 10836 2941
rect 11060 2975 11112 2984
rect 11060 2941 11069 2975
rect 11069 2941 11103 2975
rect 11103 2941 11112 2975
rect 11060 2932 11112 2941
rect 11244 2975 11296 2984
rect 11244 2941 11253 2975
rect 11253 2941 11287 2975
rect 11287 2941 11296 2975
rect 11244 2932 11296 2941
rect 12348 2932 12400 2984
rect 12900 2932 12952 2984
rect 13268 3000 13320 3052
rect 13544 2932 13596 2984
rect 13728 2932 13780 2984
rect 13820 2975 13872 2984
rect 13820 2941 13829 2975
rect 13829 2941 13863 2975
rect 13863 2941 13872 2975
rect 13820 2932 13872 2941
rect 11336 2864 11388 2916
rect 14280 2975 14332 2984
rect 14280 2941 14289 2975
rect 14289 2941 14323 2975
rect 14323 2941 14332 2975
rect 14280 2932 14332 2941
rect 14188 2864 14240 2916
rect 15016 2932 15068 2984
rect 16488 3136 16540 3188
rect 17592 3136 17644 3188
rect 18696 3136 18748 3188
rect 23756 3136 23808 3188
rect 16212 2975 16264 2984
rect 16212 2941 16221 2975
rect 16221 2941 16255 2975
rect 16255 2941 16264 2975
rect 16212 2932 16264 2941
rect 19248 3068 19300 3120
rect 19340 3068 19392 3120
rect 18144 2975 18196 2984
rect 6276 2839 6328 2848
rect 6276 2805 6285 2839
rect 6285 2805 6319 2839
rect 6319 2805 6328 2839
rect 6276 2796 6328 2805
rect 6368 2796 6420 2848
rect 8300 2796 8352 2848
rect 10048 2796 10100 2848
rect 10968 2796 11020 2848
rect 12716 2839 12768 2848
rect 12716 2805 12725 2839
rect 12725 2805 12759 2839
rect 12759 2805 12768 2839
rect 12716 2796 12768 2805
rect 12900 2839 12952 2848
rect 12900 2805 12909 2839
rect 12909 2805 12943 2839
rect 12943 2805 12952 2839
rect 12900 2796 12952 2805
rect 15844 2864 15896 2916
rect 18144 2941 18153 2975
rect 18153 2941 18187 2975
rect 18187 2941 18196 2975
rect 18144 2932 18196 2941
rect 18328 2975 18380 2984
rect 18328 2941 18337 2975
rect 18337 2941 18371 2975
rect 18371 2941 18380 2975
rect 18328 2932 18380 2941
rect 19892 3068 19944 3120
rect 21088 3068 21140 3120
rect 21456 3068 21508 3120
rect 20996 3000 21048 3052
rect 18696 2864 18748 2916
rect 19708 2932 19760 2984
rect 20352 2975 20404 2984
rect 22100 3043 22152 3052
rect 22100 3009 22109 3043
rect 22109 3009 22143 3043
rect 22143 3009 22152 3043
rect 22100 3000 22152 3009
rect 20352 2941 20367 2975
rect 20367 2941 20401 2975
rect 20401 2941 20404 2975
rect 20352 2932 20404 2941
rect 20168 2864 20220 2916
rect 21732 2864 21784 2916
rect 22192 2975 22244 2984
rect 22192 2941 22201 2975
rect 22201 2941 22235 2975
rect 22235 2941 22244 2975
rect 22192 2932 22244 2941
rect 22560 3068 22612 3120
rect 22744 3068 22796 3120
rect 23388 2975 23440 2984
rect 23388 2941 23397 2975
rect 23397 2941 23431 2975
rect 23431 2941 23440 2975
rect 23388 2932 23440 2941
rect 17684 2839 17736 2848
rect 17684 2805 17693 2839
rect 17693 2805 17727 2839
rect 17727 2805 17736 2839
rect 17684 2796 17736 2805
rect 18144 2796 18196 2848
rect 19156 2839 19208 2848
rect 19156 2805 19165 2839
rect 19165 2805 19199 2839
rect 19199 2805 19208 2839
rect 19156 2796 19208 2805
rect 19708 2839 19760 2848
rect 19708 2805 19717 2839
rect 19717 2805 19751 2839
rect 19751 2805 19760 2839
rect 19708 2796 19760 2805
rect 19984 2839 20036 2848
rect 19984 2805 19993 2839
rect 19993 2805 20027 2839
rect 20027 2805 20036 2839
rect 19984 2796 20036 2805
rect 20720 2839 20772 2848
rect 20720 2805 20729 2839
rect 20729 2805 20763 2839
rect 20763 2805 20772 2839
rect 23572 2864 23624 2916
rect 24584 3136 24636 3188
rect 25596 3136 25648 3188
rect 24308 2932 24360 2984
rect 25136 2932 25188 2984
rect 20720 2796 20772 2805
rect 23204 2796 23256 2848
rect 24860 2796 24912 2848
rect 25044 2839 25096 2848
rect 25044 2805 25053 2839
rect 25053 2805 25087 2839
rect 25087 2805 25096 2839
rect 25044 2796 25096 2805
rect 25688 2907 25740 2916
rect 25688 2873 25697 2907
rect 25697 2873 25731 2907
rect 25731 2873 25740 2907
rect 25688 2864 25740 2873
rect 26056 2864 26108 2916
rect 7114 2694 7166 2746
rect 7178 2694 7230 2746
rect 7242 2694 7294 2746
rect 7306 2694 7358 2746
rect 7370 2694 7422 2746
rect 13830 2694 13882 2746
rect 13894 2694 13946 2746
rect 13958 2694 14010 2746
rect 14022 2694 14074 2746
rect 14086 2694 14138 2746
rect 20546 2694 20598 2746
rect 20610 2694 20662 2746
rect 20674 2694 20726 2746
rect 20738 2694 20790 2746
rect 20802 2694 20854 2746
rect 27262 2694 27314 2746
rect 27326 2694 27378 2746
rect 27390 2694 27442 2746
rect 27454 2694 27506 2746
rect 27518 2694 27570 2746
rect 4712 2592 4764 2644
rect 6460 2592 6512 2644
rect 6644 2592 6696 2644
rect 8852 2635 8904 2644
rect 8852 2601 8887 2635
rect 8887 2601 8904 2635
rect 8852 2592 8904 2601
rect 2412 2456 2464 2508
rect 2688 2499 2740 2508
rect 2688 2465 2697 2499
rect 2697 2465 2731 2499
rect 2731 2465 2740 2499
rect 2688 2456 2740 2465
rect 4344 2499 4396 2508
rect 4344 2465 4353 2499
rect 4353 2465 4387 2499
rect 4387 2465 4396 2499
rect 4344 2456 4396 2465
rect 4528 2499 4580 2508
rect 4528 2465 4537 2499
rect 4537 2465 4571 2499
rect 4571 2465 4580 2499
rect 4528 2456 4580 2465
rect 4896 2456 4948 2508
rect 3792 2388 3844 2440
rect 5080 2456 5132 2508
rect 5632 2456 5684 2508
rect 6460 2499 6512 2508
rect 6460 2465 6469 2499
rect 6469 2465 6503 2499
rect 6503 2465 6512 2499
rect 6460 2456 6512 2465
rect 2688 2363 2740 2372
rect 2688 2329 2697 2363
rect 2697 2329 2731 2363
rect 2731 2329 2740 2363
rect 2688 2320 2740 2329
rect 7656 2456 7708 2508
rect 6828 2388 6880 2440
rect 9680 2592 9732 2644
rect 10784 2592 10836 2644
rect 11336 2592 11388 2644
rect 12716 2592 12768 2644
rect 12900 2592 12952 2644
rect 13728 2635 13780 2644
rect 13728 2601 13737 2635
rect 13737 2601 13771 2635
rect 13771 2601 13780 2635
rect 13728 2592 13780 2601
rect 15476 2592 15528 2644
rect 11428 2456 11480 2508
rect 9036 2388 9088 2440
rect 9496 2388 9548 2440
rect 11888 2499 11940 2508
rect 11888 2465 11897 2499
rect 11897 2465 11931 2499
rect 11931 2465 11940 2499
rect 11888 2456 11940 2465
rect 12164 2499 12216 2508
rect 12164 2465 12173 2499
rect 12173 2465 12207 2499
rect 12207 2465 12216 2499
rect 12164 2456 12216 2465
rect 12532 2499 12584 2508
rect 12532 2465 12541 2499
rect 12541 2465 12575 2499
rect 12575 2465 12584 2499
rect 12532 2456 12584 2465
rect 12716 2499 12768 2508
rect 12716 2465 12725 2499
rect 12725 2465 12759 2499
rect 12759 2465 12768 2499
rect 12716 2456 12768 2465
rect 12900 2456 12952 2508
rect 10140 2320 10192 2372
rect 10968 2320 11020 2372
rect 12624 2320 12676 2372
rect 13636 2499 13688 2508
rect 13636 2465 13645 2499
rect 13645 2465 13679 2499
rect 13679 2465 13688 2499
rect 13636 2456 13688 2465
rect 14188 2456 14240 2508
rect 14280 2499 14332 2508
rect 14280 2465 14289 2499
rect 14289 2465 14323 2499
rect 14323 2465 14332 2499
rect 14280 2456 14332 2465
rect 15384 2524 15436 2576
rect 15016 2456 15068 2508
rect 16212 2499 16264 2508
rect 16212 2465 16221 2499
rect 16221 2465 16255 2499
rect 16255 2465 16264 2499
rect 16212 2456 16264 2465
rect 17592 2524 17644 2576
rect 18328 2567 18380 2576
rect 18328 2533 18337 2567
rect 18337 2533 18371 2567
rect 18371 2533 18380 2567
rect 18328 2524 18380 2533
rect 16948 2456 17000 2508
rect 18236 2456 18288 2508
rect 20260 2499 20312 2508
rect 20260 2465 20269 2499
rect 20269 2465 20303 2499
rect 20303 2465 20312 2499
rect 20260 2456 20312 2465
rect 20904 2524 20956 2576
rect 22836 2592 22888 2644
rect 23112 2592 23164 2644
rect 26056 2592 26108 2644
rect 18144 2388 18196 2440
rect 20996 2499 21048 2508
rect 20996 2465 21005 2499
rect 21005 2465 21039 2499
rect 21039 2465 21048 2499
rect 20996 2456 21048 2465
rect 21180 2456 21232 2508
rect 21824 2456 21876 2508
rect 22192 2456 22244 2508
rect 22560 2499 22612 2508
rect 22560 2465 22569 2499
rect 22569 2465 22603 2499
rect 22603 2465 22612 2499
rect 22560 2456 22612 2465
rect 25044 2524 25096 2576
rect 14648 2320 14700 2372
rect 19708 2320 19760 2372
rect 20352 2320 20404 2372
rect 24400 2499 24452 2508
rect 24400 2465 24409 2499
rect 24409 2465 24443 2499
rect 24443 2465 24452 2499
rect 24400 2456 24452 2465
rect 24492 2499 24544 2508
rect 24492 2465 24501 2499
rect 24501 2465 24535 2499
rect 24535 2465 24544 2499
rect 24492 2456 24544 2465
rect 23296 2431 23348 2440
rect 23296 2397 23305 2431
rect 23305 2397 23339 2431
rect 23339 2397 23348 2431
rect 23296 2388 23348 2397
rect 3608 2295 3660 2304
rect 3608 2261 3617 2295
rect 3617 2261 3651 2295
rect 3651 2261 3660 2295
rect 3608 2252 3660 2261
rect 4160 2252 4212 2304
rect 4620 2252 4672 2304
rect 4804 2295 4856 2304
rect 4804 2261 4813 2295
rect 4813 2261 4847 2295
rect 4847 2261 4856 2295
rect 4804 2252 4856 2261
rect 5540 2295 5592 2304
rect 5540 2261 5549 2295
rect 5549 2261 5583 2295
rect 5583 2261 5592 2295
rect 5540 2252 5592 2261
rect 6092 2252 6144 2304
rect 7012 2295 7064 2304
rect 7012 2261 7021 2295
rect 7021 2261 7055 2295
rect 7055 2261 7064 2295
rect 7012 2252 7064 2261
rect 7104 2252 7156 2304
rect 9128 2252 9180 2304
rect 10324 2295 10376 2304
rect 10324 2261 10333 2295
rect 10333 2261 10367 2295
rect 10367 2261 10376 2295
rect 10324 2252 10376 2261
rect 11888 2295 11940 2304
rect 11888 2261 11897 2295
rect 11897 2261 11931 2295
rect 11931 2261 11940 2295
rect 11888 2252 11940 2261
rect 11980 2295 12032 2304
rect 11980 2261 11989 2295
rect 11989 2261 12023 2295
rect 12023 2261 12032 2295
rect 11980 2252 12032 2261
rect 12716 2295 12768 2304
rect 12716 2261 12725 2295
rect 12725 2261 12759 2295
rect 12759 2261 12768 2295
rect 12716 2252 12768 2261
rect 14740 2252 14792 2304
rect 14924 2252 14976 2304
rect 20444 2295 20496 2304
rect 20444 2261 20453 2295
rect 20453 2261 20487 2295
rect 20487 2261 20496 2295
rect 20444 2252 20496 2261
rect 20996 2295 21048 2304
rect 20996 2261 21005 2295
rect 21005 2261 21039 2295
rect 21039 2261 21048 2295
rect 20996 2252 21048 2261
rect 21548 2252 21600 2304
rect 3756 2150 3808 2202
rect 3820 2150 3872 2202
rect 3884 2150 3936 2202
rect 3948 2150 4000 2202
rect 4012 2150 4064 2202
rect 10472 2150 10524 2202
rect 10536 2150 10588 2202
rect 10600 2150 10652 2202
rect 10664 2150 10716 2202
rect 10728 2150 10780 2202
rect 17188 2150 17240 2202
rect 17252 2150 17304 2202
rect 17316 2150 17368 2202
rect 17380 2150 17432 2202
rect 17444 2150 17496 2202
rect 23904 2150 23956 2202
rect 23968 2150 24020 2202
rect 24032 2150 24084 2202
rect 24096 2150 24148 2202
rect 24160 2150 24212 2202
rect 4068 2048 4120 2100
rect 4804 2048 4856 2100
rect 4896 2048 4948 2100
rect 5632 2048 5684 2100
rect 6644 2048 6696 2100
rect 940 1887 992 1896
rect 940 1853 949 1887
rect 949 1853 983 1887
rect 983 1853 992 1887
rect 940 1844 992 1853
rect 1124 1844 1176 1896
rect 2688 1844 2740 1896
rect 2964 1887 3016 1896
rect 2964 1853 2973 1887
rect 2973 1853 3007 1887
rect 3007 1853 3016 1887
rect 2964 1844 3016 1853
rect 3332 1844 3384 1896
rect 3516 1844 3568 1896
rect 7012 2048 7064 2100
rect 10324 2048 10376 2100
rect 11060 2048 11112 2100
rect 15016 2048 15068 2100
rect 16948 2048 17000 2100
rect 5172 1887 5224 1896
rect 5172 1853 5181 1887
rect 5181 1853 5215 1887
rect 5215 1853 5224 1887
rect 5172 1844 5224 1853
rect 5264 1887 5316 1896
rect 5264 1853 5273 1887
rect 5273 1853 5307 1887
rect 5307 1853 5316 1887
rect 5264 1844 5316 1853
rect 5724 1844 5776 1896
rect 5816 1887 5868 1896
rect 5816 1853 5825 1887
rect 5825 1853 5859 1887
rect 5859 1853 5868 1887
rect 5816 1844 5868 1853
rect 6644 1887 6696 1896
rect 6644 1853 6653 1887
rect 6653 1853 6687 1887
rect 6687 1853 6696 1887
rect 6644 1844 6696 1853
rect 7104 1844 7156 1896
rect 7840 1887 7892 1896
rect 7840 1853 7849 1887
rect 7849 1853 7883 1887
rect 7883 1853 7892 1887
rect 7840 1844 7892 1853
rect 7932 1887 7984 1896
rect 7932 1853 7941 1887
rect 7941 1853 7975 1887
rect 7975 1853 7984 1887
rect 7932 1844 7984 1853
rect 9220 1887 9272 1896
rect 9220 1853 9229 1887
rect 9229 1853 9263 1887
rect 9263 1853 9272 1887
rect 9220 1844 9272 1853
rect 4068 1776 4120 1828
rect 3516 1751 3568 1760
rect 3516 1717 3525 1751
rect 3525 1717 3559 1751
rect 3559 1717 3568 1751
rect 3516 1708 3568 1717
rect 10140 1887 10192 1896
rect 10140 1853 10149 1887
rect 10149 1853 10183 1887
rect 10183 1853 10192 1887
rect 10140 1844 10192 1853
rect 10324 1776 10376 1828
rect 10784 1887 10836 1896
rect 10784 1853 10793 1887
rect 10793 1853 10827 1887
rect 10827 1853 10836 1887
rect 10784 1844 10836 1853
rect 11612 1887 11664 1896
rect 11612 1853 11621 1887
rect 11621 1853 11655 1887
rect 11655 1853 11664 1887
rect 11612 1844 11664 1853
rect 11704 1887 11756 1896
rect 11704 1853 11713 1887
rect 11713 1853 11747 1887
rect 11747 1853 11756 1887
rect 11704 1844 11756 1853
rect 11980 1887 12032 1896
rect 11980 1853 11989 1887
rect 11989 1853 12023 1887
rect 12023 1853 12032 1887
rect 11980 1844 12032 1853
rect 12808 1887 12860 1896
rect 12808 1853 12817 1887
rect 12817 1853 12851 1887
rect 12851 1853 12860 1887
rect 12808 1844 12860 1853
rect 12900 1887 12952 1896
rect 12900 1853 12909 1887
rect 12909 1853 12943 1887
rect 12943 1853 12952 1887
rect 12900 1844 12952 1853
rect 13176 1887 13228 1896
rect 13176 1853 13185 1887
rect 13185 1853 13219 1887
rect 13219 1853 13228 1887
rect 13176 1844 13228 1853
rect 14188 1887 14240 1896
rect 14188 1853 14197 1887
rect 14197 1853 14231 1887
rect 14231 1853 14240 1887
rect 14188 1844 14240 1853
rect 14648 1887 14700 1896
rect 14648 1853 14657 1887
rect 14657 1853 14691 1887
rect 14691 1853 14700 1887
rect 14648 1844 14700 1853
rect 15384 1844 15436 1896
rect 16304 1887 16356 1896
rect 16304 1853 16313 1887
rect 16313 1853 16347 1887
rect 16347 1853 16356 1887
rect 16304 1844 16356 1853
rect 16396 1887 16448 1896
rect 16396 1853 16405 1887
rect 16405 1853 16439 1887
rect 16439 1853 16448 1887
rect 16396 1844 16448 1853
rect 17316 1844 17368 1896
rect 17684 1887 17736 1896
rect 17684 1853 17693 1887
rect 17693 1853 17727 1887
rect 17727 1853 17736 1887
rect 17684 1844 17736 1853
rect 19800 1844 19852 1896
rect 20076 1887 20128 1896
rect 20076 1853 20085 1887
rect 20085 1853 20119 1887
rect 20119 1853 20128 1887
rect 20076 1844 20128 1853
rect 20444 1887 20496 1896
rect 20444 1853 20453 1887
rect 20453 1853 20487 1887
rect 20487 1853 20496 1887
rect 20444 1844 20496 1853
rect 21272 1887 21324 1896
rect 21272 1853 21281 1887
rect 21281 1853 21315 1887
rect 21315 1853 21324 1887
rect 21272 1844 21324 1853
rect 21456 1844 21508 1896
rect 21916 1887 21968 1896
rect 21916 1853 21925 1887
rect 21925 1853 21959 1887
rect 21959 1853 21968 1887
rect 21916 1844 21968 1853
rect 22560 1844 22612 1896
rect 22652 1887 22704 1896
rect 22652 1853 22661 1887
rect 22661 1853 22695 1887
rect 22695 1853 22704 1887
rect 22652 1844 22704 1853
rect 23296 1844 23348 1896
rect 23756 1844 23808 1896
rect 24860 1887 24912 1896
rect 24860 1853 24869 1887
rect 24869 1853 24903 1887
rect 24903 1853 24912 1887
rect 24860 1844 24912 1853
rect 26056 1844 26108 1896
rect 25320 1776 25372 1828
rect 11152 1708 11204 1760
rect 7114 1606 7166 1658
rect 7178 1606 7230 1658
rect 7242 1606 7294 1658
rect 7306 1606 7358 1658
rect 7370 1606 7422 1658
rect 13830 1606 13882 1658
rect 13894 1606 13946 1658
rect 13958 1606 14010 1658
rect 14022 1606 14074 1658
rect 14086 1606 14138 1658
rect 20546 1606 20598 1658
rect 20610 1606 20662 1658
rect 20674 1606 20726 1658
rect 20738 1606 20790 1658
rect 20802 1606 20854 1658
rect 27262 1606 27314 1658
rect 27326 1606 27378 1658
rect 27390 1606 27442 1658
rect 27454 1606 27506 1658
rect 27518 1606 27570 1658
rect 1308 1504 1360 1556
rect 2044 1504 2096 1556
rect 3516 1504 3568 1556
rect 6276 1504 6328 1556
rect 7380 1504 7432 1556
rect 7932 1504 7984 1556
rect 11888 1504 11940 1556
rect 19708 1504 19760 1556
rect 20996 1504 21048 1556
rect 22836 1504 22888 1556
rect 1124 1368 1176 1420
rect 2320 1368 2372 1420
rect 3240 1411 3292 1420
rect 3240 1377 3249 1411
rect 3249 1377 3283 1411
rect 3283 1377 3292 1411
rect 3240 1368 3292 1377
rect 4436 1411 4488 1420
rect 4436 1377 4445 1411
rect 4445 1377 4479 1411
rect 4479 1377 4488 1411
rect 4436 1368 4488 1377
rect 4712 1368 4764 1420
rect 5264 1368 5316 1420
rect 6184 1436 6236 1488
rect 5724 1368 5776 1420
rect 2136 1343 2188 1352
rect 2136 1309 2145 1343
rect 2145 1309 2179 1343
rect 2179 1309 2188 1343
rect 2136 1300 2188 1309
rect 3332 1343 3384 1352
rect 3332 1309 3341 1343
rect 3341 1309 3375 1343
rect 3375 1309 3384 1343
rect 3332 1300 3384 1309
rect 7104 1411 7156 1420
rect 7104 1377 7113 1411
rect 7113 1377 7147 1411
rect 7147 1377 7156 1411
rect 7104 1368 7156 1377
rect 8944 1436 8996 1488
rect 8300 1411 8352 1420
rect 8300 1377 8309 1411
rect 8309 1377 8343 1411
rect 8343 1377 8352 1411
rect 8300 1368 8352 1377
rect 9312 1368 9364 1420
rect 9864 1411 9916 1420
rect 9864 1377 9873 1411
rect 9873 1377 9907 1411
rect 9907 1377 9916 1411
rect 9864 1368 9916 1377
rect 10692 1411 10744 1420
rect 10692 1377 10701 1411
rect 10701 1377 10735 1411
rect 10735 1377 10744 1411
rect 10692 1368 10744 1377
rect 12164 1411 12216 1420
rect 12164 1377 12173 1411
rect 12173 1377 12207 1411
rect 12207 1377 12216 1411
rect 12164 1368 12216 1377
rect 17040 1436 17092 1488
rect 8024 1343 8076 1352
rect 8024 1309 8033 1343
rect 8033 1309 8067 1343
rect 8067 1309 8076 1343
rect 8024 1300 8076 1309
rect 11060 1343 11112 1352
rect 11060 1309 11069 1343
rect 11069 1309 11103 1343
rect 11103 1309 11112 1343
rect 11060 1300 11112 1309
rect 12624 1368 12676 1420
rect 12900 1368 12952 1420
rect 13636 1368 13688 1420
rect 13728 1411 13780 1420
rect 13728 1377 13737 1411
rect 13737 1377 13771 1411
rect 13771 1377 13780 1411
rect 13728 1368 13780 1377
rect 14556 1411 14608 1420
rect 14556 1377 14565 1411
rect 14565 1377 14599 1411
rect 14599 1377 14608 1411
rect 14556 1368 14608 1377
rect 14648 1411 14700 1420
rect 14648 1377 14657 1411
rect 14657 1377 14691 1411
rect 14691 1377 14700 1411
rect 14648 1368 14700 1377
rect 14924 1411 14976 1420
rect 14924 1377 14933 1411
rect 14933 1377 14967 1411
rect 14967 1377 14976 1411
rect 14924 1368 14976 1377
rect 15752 1411 15804 1420
rect 15752 1377 15761 1411
rect 15761 1377 15795 1411
rect 15795 1377 15804 1411
rect 15752 1368 15804 1377
rect 15844 1368 15896 1420
rect 16764 1368 16816 1420
rect 17316 1411 17368 1420
rect 17316 1377 17325 1411
rect 17325 1377 17359 1411
rect 17359 1377 17368 1411
rect 17316 1368 17368 1377
rect 17776 1368 17828 1420
rect 18512 1411 18564 1420
rect 18512 1377 18521 1411
rect 18521 1377 18555 1411
rect 18555 1377 18564 1411
rect 18512 1368 18564 1377
rect 19340 1411 19392 1420
rect 19340 1377 19349 1411
rect 19349 1377 19383 1411
rect 19383 1377 19392 1411
rect 19340 1368 19392 1377
rect 19892 1436 19944 1488
rect 21456 1368 21508 1420
rect 22100 1436 22152 1488
rect 22008 1368 22060 1420
rect 22836 1368 22888 1420
rect 24308 1368 24360 1420
rect 25136 1411 25188 1420
rect 25136 1377 25145 1411
rect 25145 1377 25179 1411
rect 25179 1377 25188 1411
rect 25136 1368 25188 1377
rect 25504 1368 25556 1420
rect 13452 1343 13504 1352
rect 13452 1309 13461 1343
rect 13461 1309 13495 1343
rect 13495 1309 13504 1343
rect 13452 1300 13504 1309
rect 16120 1343 16172 1352
rect 16120 1309 16129 1343
rect 16129 1309 16163 1343
rect 16163 1309 16172 1343
rect 16120 1300 16172 1309
rect 6276 1207 6328 1216
rect 6276 1173 6285 1207
rect 6285 1173 6319 1207
rect 6319 1173 6328 1207
rect 6276 1164 6328 1173
rect 6736 1207 6788 1216
rect 6736 1173 6745 1207
rect 6745 1173 6779 1207
rect 6779 1173 6788 1207
rect 6736 1164 6788 1173
rect 17868 1164 17920 1216
rect 19708 1343 19760 1352
rect 19708 1309 19717 1343
rect 19717 1309 19751 1343
rect 19751 1309 19760 1343
rect 19708 1300 19760 1309
rect 22468 1343 22520 1352
rect 22468 1309 22477 1343
rect 22477 1309 22511 1343
rect 22511 1309 22520 1343
rect 22468 1300 22520 1309
rect 23664 1343 23716 1352
rect 23664 1309 23673 1343
rect 23673 1309 23707 1343
rect 23707 1309 23716 1343
rect 23664 1300 23716 1309
rect 24860 1343 24912 1352
rect 24860 1309 24869 1343
rect 24869 1309 24903 1343
rect 24903 1309 24912 1343
rect 24860 1300 24912 1309
rect 21088 1207 21140 1216
rect 21088 1173 21097 1207
rect 21097 1173 21131 1207
rect 21131 1173 21140 1207
rect 21088 1164 21140 1173
rect 3756 1062 3808 1114
rect 3820 1062 3872 1114
rect 3884 1062 3936 1114
rect 3948 1062 4000 1114
rect 4012 1062 4064 1114
rect 10472 1062 10524 1114
rect 10536 1062 10588 1114
rect 10600 1062 10652 1114
rect 10664 1062 10716 1114
rect 10728 1062 10780 1114
rect 17188 1062 17240 1114
rect 17252 1062 17304 1114
rect 17316 1062 17368 1114
rect 17380 1062 17432 1114
rect 17444 1062 17496 1114
rect 23904 1062 23956 1114
rect 23968 1062 24020 1114
rect 24032 1062 24084 1114
rect 24096 1062 24148 1114
rect 24160 1062 24212 1114
rect 2136 960 2188 1012
rect 4160 960 4212 1012
rect 940 867 992 876
rect 940 833 949 867
rect 949 833 983 867
rect 983 833 992 867
rect 940 824 992 833
rect 6276 960 6328 1012
rect 6736 960 6788 1012
rect 8024 960 8076 1012
rect 10324 960 10376 1012
rect 11060 960 11112 1012
rect 11704 1003 11756 1012
rect 11704 969 11713 1003
rect 11713 969 11747 1003
rect 11747 969 11756 1003
rect 11704 960 11756 969
rect 9220 867 9272 876
rect 9220 833 9229 867
rect 9229 833 9263 867
rect 9263 833 9272 867
rect 9220 824 9272 833
rect 13176 960 13228 1012
rect 13452 960 13504 1012
rect 14188 960 14240 1012
rect 16120 960 16172 1012
rect 17868 1003 17920 1012
rect 17868 969 17877 1003
rect 17877 969 17911 1003
rect 17911 969 17920 1003
rect 17868 960 17920 969
rect 19708 960 19760 1012
rect 21088 960 21140 1012
rect 21916 960 21968 1012
rect 22468 1003 22520 1012
rect 22468 969 22477 1003
rect 22477 969 22511 1003
rect 22511 969 22520 1003
rect 22468 960 22520 969
rect 22560 960 22612 1012
rect 23664 960 23716 1012
rect 24860 960 24912 1012
rect 25320 1003 25372 1012
rect 25320 969 25329 1003
rect 25329 969 25363 1003
rect 25363 969 25372 1003
rect 25320 960 25372 969
rect 23756 824 23808 876
rect 1768 756 1820 808
rect 2504 756 2556 808
rect 3608 756 3660 808
rect 4068 756 4120 808
rect 4620 756 4672 808
rect 5540 799 5592 808
rect 5540 765 5549 799
rect 5549 765 5583 799
rect 5583 765 5592 799
rect 5540 756 5592 765
rect 6092 756 6144 808
rect 7012 799 7064 808
rect 7012 765 7021 799
rect 7021 765 7055 799
rect 7055 765 7064 799
rect 7012 756 7064 765
rect 7380 799 7432 808
rect 7380 765 7389 799
rect 7389 765 7423 799
rect 7423 765 7432 799
rect 7380 756 7432 765
rect 8300 756 8352 808
rect 9680 756 9732 808
rect 10048 756 10100 808
rect 12716 756 12768 808
rect 13360 799 13412 808
rect 13360 765 13369 799
rect 13369 765 13403 799
rect 13403 765 13412 799
rect 13360 756 13412 765
rect 14832 756 14884 808
rect 15016 756 15068 808
rect 16396 756 16448 808
rect 15936 688 15988 740
rect 17316 799 17368 808
rect 17316 765 17325 799
rect 17325 765 17359 799
rect 17359 765 17368 799
rect 17316 756 17368 765
rect 18972 799 19024 808
rect 18972 765 18981 799
rect 18981 765 19015 799
rect 19015 765 19024 799
rect 18972 756 19024 765
rect 19340 756 19392 808
rect 20260 756 20312 808
rect 20352 756 20404 808
rect 21548 799 21600 808
rect 21548 765 21557 799
rect 21557 765 21591 799
rect 21591 765 21600 799
rect 21548 756 21600 765
rect 22376 799 22428 808
rect 22376 765 22385 799
rect 22385 765 22419 799
rect 22419 765 22428 799
rect 22376 756 22428 765
rect 23572 756 23624 808
rect 24952 799 25004 808
rect 24952 765 24961 799
rect 24961 765 24995 799
rect 24995 765 25004 799
rect 24952 756 25004 765
rect 7114 518 7166 570
rect 7178 518 7230 570
rect 7242 518 7294 570
rect 7306 518 7358 570
rect 7370 518 7422 570
rect 13830 518 13882 570
rect 13894 518 13946 570
rect 13958 518 14010 570
rect 14022 518 14074 570
rect 14086 518 14138 570
rect 20546 518 20598 570
rect 20610 518 20662 570
rect 20674 518 20726 570
rect 20738 518 20790 570
rect 20802 518 20854 570
rect 27262 518 27314 570
rect 27326 518 27378 570
rect 27390 518 27442 570
rect 27454 518 27506 570
rect 27518 518 27570 570
<< metal2 >>
rect 1398 31600 1454 32000
rect 2870 31600 2926 32000
rect 4342 31600 4398 32000
rect 5814 31600 5870 32000
rect 7286 31600 7342 32000
rect 8758 31600 8814 32000
rect 10230 31600 10286 32000
rect 11702 31600 11758 32000
rect 13174 31600 13230 32000
rect 14646 31600 14702 32000
rect 16118 31600 16174 32000
rect 17590 31600 17646 32000
rect 19062 31600 19118 32000
rect 20534 31600 20590 32000
rect 22006 31600 22062 32000
rect 23478 31600 23534 32000
rect 24950 31600 25006 32000
rect 26422 31600 26478 32000
rect 1412 30938 1440 31600
rect 1400 30932 1452 30938
rect 1400 30874 1452 30880
rect 2044 30796 2096 30802
rect 2044 30738 2096 30744
rect 2056 30433 2084 30738
rect 2320 30728 2372 30734
rect 2320 30670 2372 30676
rect 2042 30424 2098 30433
rect 2042 30359 2098 30368
rect 2332 30190 2360 30670
rect 2884 30326 2912 31600
rect 3516 30796 3568 30802
rect 3516 30738 3568 30744
rect 2872 30320 2924 30326
rect 2872 30262 2924 30268
rect 2320 30184 2372 30190
rect 2320 30126 2372 30132
rect 1860 30116 1912 30122
rect 1860 30058 1912 30064
rect 1768 30048 1820 30054
rect 1768 29990 1820 29996
rect 1780 29594 1808 29990
rect 1872 29753 1900 30058
rect 3528 29850 3556 30738
rect 3608 30592 3660 30598
rect 3608 30534 3660 30540
rect 3620 30122 3648 30534
rect 3756 30492 4064 30501
rect 3756 30490 3762 30492
rect 3818 30490 3842 30492
rect 3898 30490 3922 30492
rect 3978 30490 4002 30492
rect 4058 30490 4064 30492
rect 3818 30438 3820 30490
rect 4000 30438 4002 30490
rect 3756 30436 3762 30438
rect 3818 30436 3842 30438
rect 3898 30436 3922 30438
rect 3978 30436 4002 30438
rect 4058 30436 4064 30438
rect 3756 30427 4064 30436
rect 3608 30116 3660 30122
rect 3608 30058 3660 30064
rect 3516 29844 3568 29850
rect 3516 29786 3568 29792
rect 4160 29776 4212 29782
rect 1858 29744 1914 29753
rect 4160 29718 4212 29724
rect 1858 29679 1914 29688
rect 2044 29708 2096 29714
rect 2044 29650 2096 29656
rect 3608 29708 3660 29714
rect 3608 29650 3660 29656
rect 1860 29640 1912 29646
rect 1780 29588 1860 29594
rect 1780 29582 1912 29588
rect 1780 29566 1900 29582
rect 1872 28558 1900 29566
rect 1860 28552 1912 28558
rect 1860 28494 1912 28500
rect 1216 26444 1268 26450
rect 1216 26386 1268 26392
rect 1228 26042 1256 26386
rect 1216 26036 1268 26042
rect 1216 25978 1268 25984
rect 1216 25356 1268 25362
rect 1216 25298 1268 25304
rect 1124 25152 1176 25158
rect 1124 25094 1176 25100
rect 1136 24682 1164 25094
rect 1228 24682 1256 25298
rect 1124 24676 1176 24682
rect 1124 24618 1176 24624
rect 1216 24676 1268 24682
rect 1216 24618 1268 24624
rect 1860 24676 1912 24682
rect 1860 24618 1912 24624
rect 1872 24274 1900 24618
rect 1860 24268 1912 24274
rect 1860 24210 1912 24216
rect 1124 24064 1176 24070
rect 1124 24006 1176 24012
rect 1136 23662 1164 24006
rect 848 23656 900 23662
rect 848 23598 900 23604
rect 1124 23656 1176 23662
rect 1124 23598 1176 23604
rect 860 22642 888 23598
rect 848 22636 900 22642
rect 848 22578 900 22584
rect 860 21010 888 22578
rect 1216 22500 1268 22506
rect 1216 22442 1268 22448
rect 1228 22234 1256 22442
rect 1216 22228 1268 22234
rect 1216 22170 1268 22176
rect 2056 22094 2084 29650
rect 3620 29306 3648 29650
rect 3756 29404 4064 29413
rect 3756 29402 3762 29404
rect 3818 29402 3842 29404
rect 3898 29402 3922 29404
rect 3978 29402 4002 29404
rect 4058 29402 4064 29404
rect 3818 29350 3820 29402
rect 4000 29350 4002 29402
rect 3756 29348 3762 29350
rect 3818 29348 3842 29350
rect 3898 29348 3922 29350
rect 3978 29348 4002 29350
rect 4058 29348 4064 29350
rect 3756 29339 4064 29348
rect 4172 29306 4200 29718
rect 4356 29510 4384 31600
rect 5828 30938 5856 31600
rect 7300 31226 7328 31600
rect 7300 31198 7512 31226
rect 7114 31036 7422 31045
rect 7114 31034 7120 31036
rect 7176 31034 7200 31036
rect 7256 31034 7280 31036
rect 7336 31034 7360 31036
rect 7416 31034 7422 31036
rect 7176 30982 7178 31034
rect 7358 30982 7360 31034
rect 7114 30980 7120 30982
rect 7176 30980 7200 30982
rect 7256 30980 7280 30982
rect 7336 30980 7360 30982
rect 7416 30980 7422 30982
rect 7114 30971 7422 30980
rect 7484 30938 7512 31198
rect 8772 30938 8800 31600
rect 5816 30932 5868 30938
rect 5816 30874 5868 30880
rect 7472 30932 7524 30938
rect 7472 30874 7524 30880
rect 8760 30932 8812 30938
rect 8760 30874 8812 30880
rect 10244 30818 10272 31600
rect 10244 30802 10364 30818
rect 11716 30802 11744 31600
rect 13188 30802 13216 31600
rect 13452 31204 13504 31210
rect 13452 31146 13504 31152
rect 9680 30796 9732 30802
rect 9680 30738 9732 30744
rect 9864 30796 9916 30802
rect 10244 30796 10376 30802
rect 10244 30790 10324 30796
rect 9864 30738 9916 30744
rect 10324 30738 10376 30744
rect 11704 30796 11756 30802
rect 11704 30738 11756 30744
rect 12716 30796 12768 30802
rect 12716 30738 12768 30744
rect 13176 30796 13228 30802
rect 13176 30738 13228 30744
rect 5908 30592 5960 30598
rect 5908 30534 5960 30540
rect 7380 30592 7432 30598
rect 7380 30534 7432 30540
rect 8484 30592 8536 30598
rect 8484 30534 8536 30540
rect 8760 30592 8812 30598
rect 8760 30534 8812 30540
rect 5920 30394 5948 30534
rect 5908 30388 5960 30394
rect 5908 30330 5960 30336
rect 7392 30326 7420 30534
rect 7380 30320 7432 30326
rect 7380 30262 7432 30268
rect 4528 30184 4580 30190
rect 4528 30126 4580 30132
rect 5908 30184 5960 30190
rect 5908 30126 5960 30132
rect 6828 30184 6880 30190
rect 6828 30126 6880 30132
rect 4252 29504 4304 29510
rect 4252 29446 4304 29452
rect 4344 29504 4396 29510
rect 4344 29446 4396 29452
rect 4264 29322 4292 29446
rect 3608 29300 3660 29306
rect 3608 29242 3660 29248
rect 4160 29300 4212 29306
rect 4264 29294 4476 29322
rect 4160 29242 4212 29248
rect 3056 29096 3108 29102
rect 3056 29038 3108 29044
rect 4158 29064 4214 29073
rect 2136 28620 2188 28626
rect 2136 28562 2188 28568
rect 2148 28218 2176 28562
rect 2228 28416 2280 28422
rect 2228 28358 2280 28364
rect 2780 28416 2832 28422
rect 2780 28358 2832 28364
rect 2136 28212 2188 28218
rect 2136 28154 2188 28160
rect 2240 27470 2268 28358
rect 2792 27946 2820 28358
rect 3068 28150 3096 29038
rect 3976 29028 4028 29034
rect 4028 29008 4158 29016
rect 4214 29008 4292 29016
rect 4028 28988 4292 29008
rect 3976 28970 4028 28976
rect 3240 28756 3292 28762
rect 3240 28698 3292 28704
rect 3252 28150 3280 28698
rect 4264 28694 4292 28988
rect 4448 28694 4476 29294
rect 4252 28688 4304 28694
rect 4252 28630 4304 28636
rect 4436 28688 4488 28694
rect 4436 28630 4488 28636
rect 3608 28620 3660 28626
rect 3608 28562 3660 28568
rect 3424 28416 3476 28422
rect 3424 28358 3476 28364
rect 3436 28218 3464 28358
rect 3424 28212 3476 28218
rect 3424 28154 3476 28160
rect 3056 28144 3108 28150
rect 3056 28086 3108 28092
rect 3240 28144 3292 28150
rect 3240 28086 3292 28092
rect 2872 28008 2924 28014
rect 2872 27950 2924 27956
rect 2780 27940 2832 27946
rect 2780 27882 2832 27888
rect 2504 27872 2556 27878
rect 2504 27814 2556 27820
rect 2516 27606 2544 27814
rect 2884 27674 2912 27950
rect 3620 27946 3648 28562
rect 4252 28552 4304 28558
rect 4252 28494 4304 28500
rect 3756 28316 4064 28325
rect 3756 28314 3762 28316
rect 3818 28314 3842 28316
rect 3898 28314 3922 28316
rect 3978 28314 4002 28316
rect 4058 28314 4064 28316
rect 3818 28262 3820 28314
rect 4000 28262 4002 28314
rect 3756 28260 3762 28262
rect 3818 28260 3842 28262
rect 3898 28260 3922 28262
rect 3978 28260 4002 28262
rect 4058 28260 4064 28262
rect 3756 28251 4064 28260
rect 3240 27940 3292 27946
rect 3240 27882 3292 27888
rect 3608 27940 3660 27946
rect 3608 27882 3660 27888
rect 2872 27668 2924 27674
rect 2872 27610 2924 27616
rect 2504 27600 2556 27606
rect 2504 27542 2556 27548
rect 2228 27464 2280 27470
rect 2228 27406 2280 27412
rect 2240 26586 2268 27406
rect 2504 26920 2556 26926
rect 2504 26862 2556 26868
rect 2320 26852 2372 26858
rect 2320 26794 2372 26800
rect 2228 26580 2280 26586
rect 2228 26522 2280 26528
rect 2332 26314 2360 26794
rect 2320 26308 2372 26314
rect 2320 26250 2372 26256
rect 2332 25838 2360 26250
rect 2412 26240 2464 26246
rect 2412 26182 2464 26188
rect 2424 26042 2452 26182
rect 2412 26036 2464 26042
rect 2412 25978 2464 25984
rect 2320 25832 2372 25838
rect 2320 25774 2372 25780
rect 2412 25832 2464 25838
rect 2516 25820 2544 26862
rect 2596 26784 2648 26790
rect 2596 26726 2648 26732
rect 2688 26784 2740 26790
rect 2688 26726 2740 26732
rect 2608 26246 2636 26726
rect 2700 26450 2728 26726
rect 2688 26444 2740 26450
rect 2688 26386 2740 26392
rect 2596 26240 2648 26246
rect 2596 26182 2648 26188
rect 2464 25792 2544 25820
rect 2412 25774 2464 25780
rect 2516 25702 2544 25792
rect 2504 25696 2556 25702
rect 2504 25638 2556 25644
rect 2228 25356 2280 25362
rect 2228 25298 2280 25304
rect 2412 25356 2464 25362
rect 2412 25298 2464 25304
rect 2240 24342 2268 25298
rect 2424 24954 2452 25298
rect 2596 25152 2648 25158
rect 2596 25094 2648 25100
rect 2608 24954 2636 25094
rect 2412 24948 2464 24954
rect 2412 24890 2464 24896
rect 2596 24948 2648 24954
rect 2596 24890 2648 24896
rect 2700 24614 2728 26386
rect 2964 26308 3016 26314
rect 2964 26250 3016 26256
rect 2976 25974 3004 26250
rect 3148 26240 3200 26246
rect 3148 26182 3200 26188
rect 2964 25968 3016 25974
rect 2964 25910 3016 25916
rect 3160 25838 3188 26182
rect 3148 25832 3200 25838
rect 3148 25774 3200 25780
rect 2872 25696 2924 25702
rect 2872 25638 2924 25644
rect 3056 25696 3108 25702
rect 3056 25638 3108 25644
rect 2884 24886 2912 25638
rect 3068 25498 3096 25638
rect 3056 25492 3108 25498
rect 3056 25434 3108 25440
rect 3056 24948 3108 24954
rect 3056 24890 3108 24896
rect 2872 24880 2924 24886
rect 2872 24822 2924 24828
rect 2688 24608 2740 24614
rect 2688 24550 2740 24556
rect 2228 24336 2280 24342
rect 2228 24278 2280 24284
rect 2700 24324 2728 24550
rect 3068 24410 3096 24890
rect 3160 24682 3188 25774
rect 3148 24676 3200 24682
rect 3148 24618 3200 24624
rect 3160 24410 3188 24618
rect 3056 24404 3108 24410
rect 3056 24346 3108 24352
rect 3148 24404 3200 24410
rect 3148 24346 3200 24352
rect 2780 24336 2832 24342
rect 2700 24296 2780 24324
rect 2700 23746 2728 24296
rect 2780 24278 2832 24284
rect 3068 23866 3096 24346
rect 3056 23860 3108 23866
rect 3056 23802 3108 23808
rect 2700 23718 2820 23746
rect 2688 23588 2740 23594
rect 2688 23530 2740 23536
rect 2700 23322 2728 23530
rect 2792 23322 2820 23718
rect 3056 23520 3108 23526
rect 3056 23462 3108 23468
rect 2688 23316 2740 23322
rect 2688 23258 2740 23264
rect 2780 23316 2832 23322
rect 2780 23258 2832 23264
rect 2228 23112 2280 23118
rect 2228 23054 2280 23060
rect 2240 22778 2268 23054
rect 2228 22772 2280 22778
rect 2228 22714 2280 22720
rect 2504 22772 2556 22778
rect 2504 22714 2556 22720
rect 2320 22432 2372 22438
rect 2320 22374 2372 22380
rect 2332 22234 2360 22374
rect 2516 22234 2544 22714
rect 2700 22710 2728 23258
rect 2688 22704 2740 22710
rect 2688 22646 2740 22652
rect 2792 22438 2820 23258
rect 2872 23180 2924 23186
rect 2872 23122 2924 23128
rect 2780 22432 2832 22438
rect 2780 22374 2832 22380
rect 2320 22228 2372 22234
rect 2320 22170 2372 22176
rect 2504 22228 2556 22234
rect 2504 22170 2556 22176
rect 2884 22166 2912 23122
rect 3068 22982 3096 23462
rect 3056 22976 3108 22982
rect 3056 22918 3108 22924
rect 2964 22772 3016 22778
rect 2964 22714 3016 22720
rect 2976 22234 3004 22714
rect 3148 22432 3200 22438
rect 3148 22374 3200 22380
rect 3160 22234 3188 22374
rect 2964 22228 3016 22234
rect 2964 22170 3016 22176
rect 3148 22228 3200 22234
rect 3148 22170 3200 22176
rect 2872 22160 2924 22166
rect 2872 22102 2924 22108
rect 1872 22066 2084 22094
rect 1584 21480 1636 21486
rect 1584 21422 1636 21428
rect 1032 21344 1084 21350
rect 1032 21286 1084 21292
rect 848 21004 900 21010
rect 848 20946 900 20952
rect 860 20398 888 20946
rect 848 20392 900 20398
rect 848 20334 900 20340
rect 860 19310 888 20334
rect 848 19304 900 19310
rect 848 19246 900 19252
rect 860 18834 888 19246
rect 1044 19174 1072 21286
rect 1596 20942 1624 21422
rect 1584 20936 1636 20942
rect 1584 20878 1636 20884
rect 1124 20800 1176 20806
rect 1124 20742 1176 20748
rect 1136 20398 1164 20742
rect 1124 20392 1176 20398
rect 1124 20334 1176 20340
rect 1400 19916 1452 19922
rect 1400 19858 1452 19864
rect 1124 19712 1176 19718
rect 1124 19654 1176 19660
rect 1136 19310 1164 19654
rect 1124 19304 1176 19310
rect 1124 19246 1176 19252
rect 1032 19168 1084 19174
rect 1032 19110 1084 19116
rect 1044 18834 1072 19110
rect 1412 18970 1440 19858
rect 1400 18964 1452 18970
rect 1400 18906 1452 18912
rect 848 18828 900 18834
rect 848 18770 900 18776
rect 1032 18828 1084 18834
rect 1032 18770 1084 18776
rect 860 17746 888 18770
rect 1400 18692 1452 18698
rect 1400 18634 1452 18640
rect 1412 18222 1440 18634
rect 1400 18216 1452 18222
rect 1400 18158 1452 18164
rect 1676 18080 1728 18086
rect 1676 18022 1728 18028
rect 1768 18080 1820 18086
rect 1768 18022 1820 18028
rect 848 17740 900 17746
rect 848 17682 900 17688
rect 1400 17740 1452 17746
rect 1400 17682 1452 17688
rect 1412 17338 1440 17682
rect 1400 17332 1452 17338
rect 1400 17274 1452 17280
rect 1688 17134 1716 18022
rect 1780 17882 1808 18022
rect 1768 17876 1820 17882
rect 1768 17818 1820 17824
rect 1780 17338 1808 17818
rect 1768 17332 1820 17338
rect 1768 17274 1820 17280
rect 1676 17128 1728 17134
rect 1676 17070 1728 17076
rect 1032 16652 1084 16658
rect 1032 16594 1084 16600
rect 940 15564 992 15570
rect 940 15506 992 15512
rect 952 15162 980 15506
rect 940 15156 992 15162
rect 940 15098 992 15104
rect 1044 15026 1072 16594
rect 1676 15972 1728 15978
rect 1676 15914 1728 15920
rect 1688 15706 1716 15914
rect 1768 15904 1820 15910
rect 1768 15846 1820 15852
rect 1780 15706 1808 15846
rect 1676 15700 1728 15706
rect 1676 15642 1728 15648
rect 1768 15700 1820 15706
rect 1768 15642 1820 15648
rect 1124 15360 1176 15366
rect 1124 15302 1176 15308
rect 1584 15360 1636 15366
rect 1584 15302 1636 15308
rect 1032 15020 1084 15026
rect 1032 14962 1084 14968
rect 1044 14618 1072 14962
rect 1032 14612 1084 14618
rect 1032 14554 1084 14560
rect 1136 14550 1164 15302
rect 1124 14544 1176 14550
rect 1124 14486 1176 14492
rect 1308 13796 1360 13802
rect 1308 13738 1360 13744
rect 1124 13728 1176 13734
rect 1320 13682 1348 13738
rect 1124 13670 1176 13676
rect 1136 12782 1164 13670
rect 1228 13654 1348 13682
rect 1228 13190 1256 13654
rect 1216 13184 1268 13190
rect 1216 13126 1268 13132
rect 1124 12776 1176 12782
rect 1124 12718 1176 12724
rect 1136 12434 1164 12718
rect 1044 12406 1164 12434
rect 1044 12306 1072 12406
rect 1032 12300 1084 12306
rect 1032 12242 1084 12248
rect 1044 10606 1072 12242
rect 1228 12186 1256 13126
rect 1308 12640 1360 12646
rect 1308 12582 1360 12588
rect 1136 12158 1256 12186
rect 1136 12102 1164 12158
rect 1124 12096 1176 12102
rect 1320 12050 1348 12582
rect 1124 12038 1176 12044
rect 1136 11540 1164 12038
rect 1228 12022 1348 12050
rect 1228 11694 1256 12022
rect 1216 11688 1268 11694
rect 1216 11630 1268 11636
rect 1492 11552 1544 11558
rect 1136 11512 1256 11540
rect 1124 11212 1176 11218
rect 1124 11154 1176 11160
rect 1136 10810 1164 11154
rect 1124 10804 1176 10810
rect 1124 10746 1176 10752
rect 1228 10606 1256 11512
rect 1492 11494 1544 11500
rect 1504 10674 1532 11494
rect 1492 10668 1544 10674
rect 1492 10610 1544 10616
rect 1032 10600 1084 10606
rect 1032 10542 1084 10548
rect 1216 10600 1268 10606
rect 1216 10542 1268 10548
rect 1308 10056 1360 10062
rect 1308 9998 1360 10004
rect 848 9376 900 9382
rect 848 9318 900 9324
rect 860 9042 888 9318
rect 1320 9178 1348 9998
rect 1308 9172 1360 9178
rect 1308 9114 1360 9120
rect 848 9036 900 9042
rect 848 8978 900 8984
rect 1596 8498 1624 15302
rect 1768 14544 1820 14550
rect 1768 14486 1820 14492
rect 1780 12306 1808 14486
rect 1676 12300 1728 12306
rect 1676 12242 1728 12248
rect 1768 12300 1820 12306
rect 1768 12242 1820 12248
rect 1688 10810 1716 12242
rect 1768 11688 1820 11694
rect 1768 11630 1820 11636
rect 1780 11354 1808 11630
rect 1768 11348 1820 11354
rect 1768 11290 1820 11296
rect 1676 10804 1728 10810
rect 1676 10746 1728 10752
rect 1872 10266 1900 22066
rect 2228 21480 2280 21486
rect 2228 21422 2280 21428
rect 2412 21480 2464 21486
rect 2412 21422 2464 21428
rect 2780 21480 2832 21486
rect 2780 21422 2832 21428
rect 2240 20602 2268 21422
rect 2228 20596 2280 20602
rect 2228 20538 2280 20544
rect 2320 20392 2372 20398
rect 2320 20334 2372 20340
rect 2332 19334 2360 20334
rect 2240 19306 2360 19334
rect 1952 18964 2004 18970
rect 1952 18906 2004 18912
rect 1964 18290 1992 18906
rect 2240 18834 2268 19306
rect 2228 18828 2280 18834
rect 2228 18770 2280 18776
rect 1952 18284 2004 18290
rect 1952 18226 2004 18232
rect 1964 17202 1992 18226
rect 2240 18222 2268 18770
rect 2424 18358 2452 21422
rect 2688 21344 2740 21350
rect 2688 21286 2740 21292
rect 2700 21146 2728 21286
rect 2688 21140 2740 21146
rect 2688 21082 2740 21088
rect 2792 20602 2820 21422
rect 2780 20596 2832 20602
rect 2780 20538 2832 20544
rect 2872 20256 2924 20262
rect 2872 20198 2924 20204
rect 2884 19990 2912 20198
rect 2872 19984 2924 19990
rect 2872 19926 2924 19932
rect 3160 19310 3188 22170
rect 3252 21078 3280 27882
rect 3620 27402 3648 27882
rect 4264 27606 4292 28494
rect 4448 27674 4476 28630
rect 4540 28218 4568 30126
rect 5448 30116 5500 30122
rect 5448 30058 5500 30064
rect 5172 30048 5224 30054
rect 5172 29990 5224 29996
rect 5080 29640 5132 29646
rect 5080 29582 5132 29588
rect 4804 29504 4856 29510
rect 4804 29446 4856 29452
rect 4896 29504 4948 29510
rect 4896 29446 4948 29452
rect 4620 29096 4672 29102
rect 4618 29064 4620 29073
rect 4672 29064 4674 29073
rect 4816 29034 4844 29446
rect 4908 29306 4936 29446
rect 5092 29306 5120 29582
rect 4896 29300 4948 29306
rect 4896 29242 4948 29248
rect 5080 29300 5132 29306
rect 5080 29242 5132 29248
rect 4618 28999 4674 29008
rect 4804 29028 4856 29034
rect 4804 28970 4856 28976
rect 4816 28694 4844 28970
rect 4804 28688 4856 28694
rect 4804 28630 4856 28636
rect 4528 28212 4580 28218
rect 4528 28154 4580 28160
rect 4436 27668 4488 27674
rect 4436 27610 4488 27616
rect 4252 27600 4304 27606
rect 4252 27542 4304 27548
rect 3608 27396 3660 27402
rect 3608 27338 3660 27344
rect 3756 27228 4064 27237
rect 3756 27226 3762 27228
rect 3818 27226 3842 27228
rect 3898 27226 3922 27228
rect 3978 27226 4002 27228
rect 4058 27226 4064 27228
rect 3818 27174 3820 27226
rect 4000 27174 4002 27226
rect 3756 27172 3762 27174
rect 3818 27172 3842 27174
rect 3898 27172 3922 27174
rect 3978 27172 4002 27174
rect 4058 27172 4064 27174
rect 3756 27163 4064 27172
rect 4264 27130 4292 27542
rect 4252 27124 4304 27130
rect 4252 27066 4304 27072
rect 3332 26444 3384 26450
rect 3332 26386 3384 26392
rect 3516 26444 3568 26450
rect 3516 26386 3568 26392
rect 3344 25770 3372 26386
rect 3424 26240 3476 26246
rect 3424 26182 3476 26188
rect 3332 25764 3384 25770
rect 3332 25706 3384 25712
rect 3436 25498 3464 26182
rect 3528 25498 3556 26386
rect 3608 26240 3660 26246
rect 3608 26182 3660 26188
rect 3620 25770 3648 26182
rect 3756 26140 4064 26149
rect 3756 26138 3762 26140
rect 3818 26138 3842 26140
rect 3898 26138 3922 26140
rect 3978 26138 4002 26140
rect 4058 26138 4064 26140
rect 3818 26086 3820 26138
rect 4000 26086 4002 26138
rect 3756 26084 3762 26086
rect 3818 26084 3842 26086
rect 3898 26084 3922 26086
rect 3978 26084 4002 26086
rect 4058 26084 4064 26086
rect 3756 26075 4064 26084
rect 3608 25764 3660 25770
rect 3608 25706 3660 25712
rect 3424 25492 3476 25498
rect 3424 25434 3476 25440
rect 3516 25492 3568 25498
rect 3516 25434 3568 25440
rect 4448 25362 4476 27610
rect 4620 27532 4672 27538
rect 4620 27474 4672 27480
rect 4632 27334 4660 27474
rect 4620 27328 4672 27334
rect 4620 27270 4672 27276
rect 5080 26920 5132 26926
rect 5080 26862 5132 26868
rect 4988 26444 5040 26450
rect 4988 26386 5040 26392
rect 4528 26036 4580 26042
rect 4528 25978 4580 25984
rect 4436 25356 4488 25362
rect 4436 25298 4488 25304
rect 4448 25158 4476 25298
rect 4436 25152 4488 25158
rect 4436 25094 4488 25100
rect 3756 25052 4064 25061
rect 3756 25050 3762 25052
rect 3818 25050 3842 25052
rect 3898 25050 3922 25052
rect 3978 25050 4002 25052
rect 4058 25050 4064 25052
rect 3818 24998 3820 25050
rect 4000 24998 4002 25050
rect 3756 24996 3762 24998
rect 3818 24996 3842 24998
rect 3898 24996 3922 24998
rect 3978 24996 4002 24998
rect 4058 24996 4064 24998
rect 3756 24987 4064 24996
rect 3424 24744 3476 24750
rect 3424 24686 3476 24692
rect 3436 24070 3464 24686
rect 3516 24268 3568 24274
rect 3516 24210 3568 24216
rect 3424 24064 3476 24070
rect 3424 24006 3476 24012
rect 3332 23656 3384 23662
rect 3332 23598 3384 23604
rect 3344 23322 3372 23598
rect 3332 23316 3384 23322
rect 3332 23258 3384 23264
rect 3436 23118 3464 24006
rect 3528 23866 3556 24210
rect 3608 24064 3660 24070
rect 3608 24006 3660 24012
rect 3516 23860 3568 23866
rect 3516 23802 3568 23808
rect 3620 23662 3648 24006
rect 3756 23964 4064 23973
rect 3756 23962 3762 23964
rect 3818 23962 3842 23964
rect 3898 23962 3922 23964
rect 3978 23962 4002 23964
rect 4058 23962 4064 23964
rect 3818 23910 3820 23962
rect 4000 23910 4002 23962
rect 3756 23908 3762 23910
rect 3818 23908 3842 23910
rect 3898 23908 3922 23910
rect 3978 23908 4002 23910
rect 4058 23908 4064 23910
rect 3756 23899 4064 23908
rect 3608 23656 3660 23662
rect 3608 23598 3660 23604
rect 3516 23520 3568 23526
rect 3516 23462 3568 23468
rect 3528 23322 3556 23462
rect 3516 23316 3568 23322
rect 3516 23258 3568 23264
rect 3620 23254 3648 23598
rect 3608 23248 3660 23254
rect 3608 23190 3660 23196
rect 4068 23180 4120 23186
rect 4068 23122 4120 23128
rect 3424 23112 3476 23118
rect 3424 23054 3476 23060
rect 4080 23066 4108 23122
rect 4080 23038 4200 23066
rect 3608 22976 3660 22982
rect 3608 22918 3660 22924
rect 3424 22568 3476 22574
rect 3424 22510 3476 22516
rect 3436 22094 3464 22510
rect 3620 22438 3648 22918
rect 3756 22876 4064 22885
rect 3756 22874 3762 22876
rect 3818 22874 3842 22876
rect 3898 22874 3922 22876
rect 3978 22874 4002 22876
rect 4058 22874 4064 22876
rect 3818 22822 3820 22874
rect 4000 22822 4002 22874
rect 3756 22820 3762 22822
rect 3818 22820 3842 22822
rect 3898 22820 3922 22822
rect 3978 22820 4002 22822
rect 4058 22820 4064 22822
rect 3756 22811 4064 22820
rect 4172 22760 4200 23038
rect 4080 22732 4200 22760
rect 3608 22432 3660 22438
rect 3608 22374 3660 22380
rect 4080 22234 4108 22732
rect 4068 22228 4120 22234
rect 4068 22170 4120 22176
rect 3436 22066 3648 22094
rect 3516 21616 3568 21622
rect 3516 21558 3568 21564
rect 3424 21480 3476 21486
rect 3424 21422 3476 21428
rect 3332 21344 3384 21350
rect 3332 21286 3384 21292
rect 3240 21072 3292 21078
rect 3240 21014 3292 21020
rect 3344 20602 3372 21286
rect 3436 21146 3464 21422
rect 3424 21140 3476 21146
rect 3424 21082 3476 21088
rect 3332 20596 3384 20602
rect 3332 20538 3384 20544
rect 3332 20460 3384 20466
rect 3332 20402 3384 20408
rect 2596 19304 2648 19310
rect 2596 19246 2648 19252
rect 2872 19304 2924 19310
rect 2872 19246 2924 19252
rect 3148 19304 3200 19310
rect 3148 19246 3200 19252
rect 2608 18970 2636 19246
rect 2780 19168 2832 19174
rect 2780 19110 2832 19116
rect 2596 18964 2648 18970
rect 2596 18906 2648 18912
rect 2792 18902 2820 19110
rect 2780 18896 2832 18902
rect 2780 18838 2832 18844
rect 2884 18426 2912 19246
rect 2872 18420 2924 18426
rect 2872 18362 2924 18368
rect 3160 18358 3188 19246
rect 3344 19242 3372 20402
rect 3436 20330 3464 21082
rect 3528 20602 3556 21558
rect 3620 20942 3648 22066
rect 3756 21788 4064 21797
rect 3756 21786 3762 21788
rect 3818 21786 3842 21788
rect 3898 21786 3922 21788
rect 3978 21786 4002 21788
rect 4058 21786 4064 21788
rect 3818 21734 3820 21786
rect 4000 21734 4002 21786
rect 3756 21732 3762 21734
rect 3818 21732 3842 21734
rect 3898 21732 3922 21734
rect 3978 21732 4002 21734
rect 4058 21732 4064 21734
rect 3756 21723 4064 21732
rect 3792 21684 3844 21690
rect 3792 21626 3844 21632
rect 3804 21486 3832 21626
rect 3792 21480 3844 21486
rect 3792 21422 3844 21428
rect 3608 20936 3660 20942
rect 3608 20878 3660 20884
rect 3620 20602 3648 20878
rect 3756 20700 4064 20709
rect 3756 20698 3762 20700
rect 3818 20698 3842 20700
rect 3898 20698 3922 20700
rect 3978 20698 4002 20700
rect 4058 20698 4064 20700
rect 3818 20646 3820 20698
rect 4000 20646 4002 20698
rect 3756 20644 3762 20646
rect 3818 20644 3842 20646
rect 3898 20644 3922 20646
rect 3978 20644 4002 20646
rect 4058 20644 4064 20646
rect 3756 20635 4064 20644
rect 3516 20596 3568 20602
rect 3516 20538 3568 20544
rect 3608 20596 3660 20602
rect 3608 20538 3660 20544
rect 4448 20398 4476 25094
rect 4540 24886 4568 25978
rect 4804 24948 4856 24954
rect 4804 24890 4856 24896
rect 4528 24880 4580 24886
rect 4528 24822 4580 24828
rect 4816 24614 4844 24890
rect 4804 24608 4856 24614
rect 4804 24550 4856 24556
rect 4896 24608 4948 24614
rect 4896 24550 4948 24556
rect 4816 24342 4844 24550
rect 4804 24336 4856 24342
rect 4804 24278 4856 24284
rect 4908 24138 4936 24550
rect 4896 24132 4948 24138
rect 4896 24074 4948 24080
rect 4712 23792 4764 23798
rect 4712 23734 4764 23740
rect 4724 23186 4752 23734
rect 5000 23610 5028 26386
rect 5092 26314 5120 26862
rect 5080 26308 5132 26314
rect 5080 26250 5132 26256
rect 5092 24818 5120 26250
rect 5080 24812 5132 24818
rect 5080 24754 5132 24760
rect 5000 23582 5120 23610
rect 5184 23594 5212 29990
rect 5460 29102 5488 30058
rect 5540 30048 5592 30054
rect 5540 29990 5592 29996
rect 5816 30048 5868 30054
rect 5816 29990 5868 29996
rect 5448 29096 5500 29102
rect 5448 29038 5500 29044
rect 5264 27532 5316 27538
rect 5264 27474 5316 27480
rect 5276 27130 5304 27474
rect 5264 27124 5316 27130
rect 5264 27066 5316 27072
rect 5356 27124 5408 27130
rect 5356 27066 5408 27072
rect 5264 26988 5316 26994
rect 5368 26976 5396 27066
rect 5316 26948 5396 26976
rect 5264 26930 5316 26936
rect 5448 26240 5500 26246
rect 5448 26182 5500 26188
rect 5264 25764 5316 25770
rect 5264 25706 5316 25712
rect 5276 25498 5304 25706
rect 5460 25498 5488 26182
rect 5264 25492 5316 25498
rect 5264 25434 5316 25440
rect 5448 25492 5500 25498
rect 5448 25434 5500 25440
rect 5448 24608 5500 24614
rect 5448 24550 5500 24556
rect 5264 24268 5316 24274
rect 5264 24210 5316 24216
rect 5276 23866 5304 24210
rect 5264 23860 5316 23866
rect 5264 23802 5316 23808
rect 4896 23520 4948 23526
rect 4896 23462 4948 23468
rect 4988 23520 5040 23526
rect 4988 23462 5040 23468
rect 4908 23322 4936 23462
rect 4896 23316 4948 23322
rect 4896 23258 4948 23264
rect 5000 23186 5028 23462
rect 4712 23180 4764 23186
rect 4712 23122 4764 23128
rect 4988 23180 5040 23186
rect 4988 23122 5040 23128
rect 4528 23044 4580 23050
rect 4528 22986 4580 22992
rect 4540 22778 4568 22986
rect 4528 22772 4580 22778
rect 4528 22714 4580 22720
rect 4724 22710 4752 23122
rect 4712 22704 4764 22710
rect 4712 22646 4764 22652
rect 5000 22574 5028 23122
rect 5092 22574 5120 23582
rect 5172 23588 5224 23594
rect 5172 23530 5224 23536
rect 5356 23588 5408 23594
rect 5356 23530 5408 23536
rect 5264 23520 5316 23526
rect 5264 23462 5316 23468
rect 5172 23180 5224 23186
rect 5172 23122 5224 23128
rect 4988 22568 5040 22574
rect 4988 22510 5040 22516
rect 5080 22568 5132 22574
rect 5080 22510 5132 22516
rect 4896 22432 4948 22438
rect 4896 22374 4948 22380
rect 4908 21894 4936 22374
rect 4896 21888 4948 21894
rect 4896 21830 4948 21836
rect 5000 21486 5028 22510
rect 5184 22506 5212 23122
rect 5172 22500 5224 22506
rect 5172 22442 5224 22448
rect 5184 21554 5212 22442
rect 5276 21690 5304 23462
rect 5264 21684 5316 21690
rect 5264 21626 5316 21632
rect 5172 21548 5224 21554
rect 5172 21490 5224 21496
rect 4988 21480 5040 21486
rect 5040 21440 5120 21468
rect 4988 21422 5040 21428
rect 4896 21344 4948 21350
rect 4896 21286 4948 21292
rect 4436 20392 4488 20398
rect 4436 20334 4488 20340
rect 3424 20324 3476 20330
rect 3424 20266 3476 20272
rect 3976 20324 4028 20330
rect 3976 20266 4028 20272
rect 3988 20058 4016 20266
rect 3976 20052 4028 20058
rect 3976 19994 4028 20000
rect 4448 19990 4476 20334
rect 4436 19984 4488 19990
rect 4436 19926 4488 19932
rect 3756 19612 4064 19621
rect 3756 19610 3762 19612
rect 3818 19610 3842 19612
rect 3898 19610 3922 19612
rect 3978 19610 4002 19612
rect 4058 19610 4064 19612
rect 3818 19558 3820 19610
rect 4000 19558 4002 19610
rect 3756 19556 3762 19558
rect 3818 19556 3842 19558
rect 3898 19556 3922 19558
rect 3978 19556 4002 19558
rect 4058 19556 4064 19558
rect 3756 19547 4064 19556
rect 4448 19514 4476 19926
rect 4908 19718 4936 21286
rect 5092 21146 5120 21440
rect 5080 21140 5132 21146
rect 5000 21100 5080 21128
rect 5000 20602 5028 21100
rect 5080 21082 5132 21088
rect 5080 20800 5132 20806
rect 5080 20742 5132 20748
rect 4988 20596 5040 20602
rect 4988 20538 5040 20544
rect 5000 19922 5028 20538
rect 5092 20058 5120 20742
rect 5264 20256 5316 20262
rect 5264 20198 5316 20204
rect 5276 20058 5304 20198
rect 5080 20052 5132 20058
rect 5080 19994 5132 20000
rect 5264 20052 5316 20058
rect 5264 19994 5316 20000
rect 4988 19916 5040 19922
rect 4988 19858 5040 19864
rect 4896 19712 4948 19718
rect 4896 19654 4948 19660
rect 4436 19508 4488 19514
rect 4436 19450 4488 19456
rect 4160 19304 4212 19310
rect 4160 19246 4212 19252
rect 4620 19304 4672 19310
rect 4620 19246 4672 19252
rect 3332 19236 3384 19242
rect 3332 19178 3384 19184
rect 4172 18630 4200 19246
rect 4252 19168 4304 19174
rect 4252 19110 4304 19116
rect 4264 18834 4292 19110
rect 4252 18828 4304 18834
rect 4252 18770 4304 18776
rect 3608 18624 3660 18630
rect 3608 18566 3660 18572
rect 4160 18624 4212 18630
rect 4160 18566 4212 18572
rect 3620 18358 3648 18566
rect 3756 18524 4064 18533
rect 3756 18522 3762 18524
rect 3818 18522 3842 18524
rect 3898 18522 3922 18524
rect 3978 18522 4002 18524
rect 4058 18522 4064 18524
rect 3818 18470 3820 18522
rect 4000 18470 4002 18522
rect 3756 18468 3762 18470
rect 3818 18468 3842 18470
rect 3898 18468 3922 18470
rect 3978 18468 4002 18470
rect 4058 18468 4064 18470
rect 3756 18459 4064 18468
rect 2412 18352 2464 18358
rect 2412 18294 2464 18300
rect 3056 18352 3108 18358
rect 3056 18294 3108 18300
rect 3148 18352 3200 18358
rect 3148 18294 3200 18300
rect 3424 18352 3476 18358
rect 3424 18294 3476 18300
rect 3608 18352 3660 18358
rect 3608 18294 3660 18300
rect 2228 18216 2280 18222
rect 2228 18158 2280 18164
rect 2320 18080 2372 18086
rect 2320 18022 2372 18028
rect 1952 17196 2004 17202
rect 1952 17138 2004 17144
rect 2136 16040 2188 16046
rect 2136 15982 2188 15988
rect 1952 15972 2004 15978
rect 1952 15914 2004 15920
rect 1964 12442 1992 15914
rect 2148 15434 2176 15982
rect 2332 15978 2360 18022
rect 2780 17604 2832 17610
rect 2780 17546 2832 17552
rect 2792 17338 2820 17546
rect 2780 17332 2832 17338
rect 2780 17274 2832 17280
rect 2964 17264 3016 17270
rect 2964 17206 3016 17212
rect 2504 17196 2556 17202
rect 2504 17138 2556 17144
rect 2516 16998 2544 17138
rect 2412 16992 2464 16998
rect 2412 16934 2464 16940
rect 2504 16992 2556 16998
rect 2504 16934 2556 16940
rect 2424 16794 2452 16934
rect 2412 16788 2464 16794
rect 2412 16730 2464 16736
rect 2688 16652 2740 16658
rect 2688 16594 2740 16600
rect 2872 16652 2924 16658
rect 2872 16594 2924 16600
rect 2700 16250 2728 16594
rect 2688 16244 2740 16250
rect 2688 16186 2740 16192
rect 2596 16108 2648 16114
rect 2596 16050 2648 16056
rect 2412 16040 2464 16046
rect 2412 15982 2464 15988
rect 2320 15972 2372 15978
rect 2320 15914 2372 15920
rect 2136 15428 2188 15434
rect 2136 15370 2188 15376
rect 2044 15156 2096 15162
rect 2044 15098 2096 15104
rect 2056 13274 2084 15098
rect 2148 14550 2176 15370
rect 2332 15366 2360 15914
rect 2424 15570 2452 15982
rect 2608 15706 2636 16050
rect 2884 16046 2912 16594
rect 2976 16522 3004 17206
rect 2964 16516 3016 16522
rect 2964 16458 3016 16464
rect 2976 16046 3004 16458
rect 2872 16040 2924 16046
rect 2872 15982 2924 15988
rect 2964 16040 3016 16046
rect 2964 15982 3016 15988
rect 2596 15700 2648 15706
rect 2596 15642 2648 15648
rect 2412 15564 2464 15570
rect 2412 15506 2464 15512
rect 2424 15450 2452 15506
rect 2424 15422 2544 15450
rect 2320 15360 2372 15366
rect 2320 15302 2372 15308
rect 2412 15360 2464 15366
rect 2412 15302 2464 15308
rect 2424 14958 2452 15302
rect 2516 14958 2544 15422
rect 2780 15360 2832 15366
rect 2780 15302 2832 15308
rect 2792 15178 2820 15302
rect 2700 15162 2820 15178
rect 2688 15156 2820 15162
rect 2740 15150 2820 15156
rect 2688 15098 2740 15104
rect 2412 14952 2464 14958
rect 2412 14894 2464 14900
rect 2504 14952 2556 14958
rect 2504 14894 2556 14900
rect 2320 14816 2372 14822
rect 2320 14758 2372 14764
rect 2136 14544 2188 14550
rect 2136 14486 2188 14492
rect 2332 14278 2360 14758
rect 2516 14482 2544 14894
rect 2688 14544 2740 14550
rect 2688 14486 2740 14492
rect 2504 14476 2556 14482
rect 2504 14418 2556 14424
rect 2320 14272 2372 14278
rect 2320 14214 2372 14220
rect 2136 13728 2188 13734
rect 2136 13670 2188 13676
rect 2228 13728 2280 13734
rect 2228 13670 2280 13676
rect 2148 13394 2176 13670
rect 2240 13530 2268 13670
rect 2228 13524 2280 13530
rect 2228 13466 2280 13472
rect 2136 13388 2188 13394
rect 2136 13330 2188 13336
rect 2228 13388 2280 13394
rect 2228 13330 2280 13336
rect 2240 13274 2268 13330
rect 2056 13246 2268 13274
rect 2240 12782 2268 13246
rect 2228 12776 2280 12782
rect 2228 12718 2280 12724
rect 2332 12714 2360 14214
rect 2516 13530 2544 14418
rect 2700 13530 2728 14486
rect 2780 14476 2832 14482
rect 2780 14418 2832 14424
rect 2792 14074 2820 14418
rect 2780 14068 2832 14074
rect 2780 14010 2832 14016
rect 2872 13864 2924 13870
rect 2872 13806 2924 13812
rect 2884 13530 2912 13806
rect 3068 13734 3096 18294
rect 3436 17814 3464 18294
rect 3608 18216 3660 18222
rect 3608 18158 3660 18164
rect 3424 17808 3476 17814
rect 3424 17750 3476 17756
rect 3516 17808 3568 17814
rect 3516 17750 3568 17756
rect 3436 17678 3464 17750
rect 3424 17672 3476 17678
rect 3424 17614 3476 17620
rect 3332 17536 3384 17542
rect 3332 17478 3384 17484
rect 3344 17066 3372 17478
rect 3528 17134 3556 17750
rect 3620 17746 3648 18158
rect 4632 17882 4660 19246
rect 4988 19236 5040 19242
rect 4988 19178 5040 19184
rect 5080 19236 5132 19242
rect 5080 19178 5132 19184
rect 4620 17876 4672 17882
rect 4620 17818 4672 17824
rect 4896 17876 4948 17882
rect 4896 17818 4948 17824
rect 3608 17740 3660 17746
rect 3608 17682 3660 17688
rect 4620 17740 4672 17746
rect 4620 17682 4672 17688
rect 4160 17604 4212 17610
rect 4160 17546 4212 17552
rect 3756 17436 4064 17445
rect 3756 17434 3762 17436
rect 3818 17434 3842 17436
rect 3898 17434 3922 17436
rect 3978 17434 4002 17436
rect 4058 17434 4064 17436
rect 3818 17382 3820 17434
rect 4000 17382 4002 17434
rect 3756 17380 3762 17382
rect 3818 17380 3842 17382
rect 3898 17380 3922 17382
rect 3978 17380 4002 17382
rect 4058 17380 4064 17382
rect 3756 17371 4064 17380
rect 4172 17338 4200 17546
rect 4436 17536 4488 17542
rect 4436 17478 4488 17484
rect 4160 17332 4212 17338
rect 4160 17274 4212 17280
rect 4252 17332 4304 17338
rect 4252 17274 4304 17280
rect 3516 17128 3568 17134
rect 3516 17070 3568 17076
rect 3332 17060 3384 17066
rect 3332 17002 3384 17008
rect 3240 16992 3292 16998
rect 3240 16934 3292 16940
rect 3252 16658 3280 16934
rect 3344 16794 3372 17002
rect 3332 16788 3384 16794
rect 3332 16730 3384 16736
rect 3240 16652 3292 16658
rect 3240 16594 3292 16600
rect 3756 16348 4064 16357
rect 3756 16346 3762 16348
rect 3818 16346 3842 16348
rect 3898 16346 3922 16348
rect 3978 16346 4002 16348
rect 4058 16346 4064 16348
rect 3818 16294 3820 16346
rect 4000 16294 4002 16346
rect 3756 16292 3762 16294
rect 3818 16292 3842 16294
rect 3898 16292 3922 16294
rect 3978 16292 4002 16294
rect 4058 16292 4064 16294
rect 3756 16283 4064 16292
rect 3332 15972 3384 15978
rect 3332 15914 3384 15920
rect 3148 15496 3200 15502
rect 3148 15438 3200 15444
rect 3160 14822 3188 15438
rect 3148 14816 3200 14822
rect 3148 14758 3200 14764
rect 3344 14550 3372 15914
rect 4264 15570 4292 17274
rect 4448 16794 4476 17478
rect 4632 17338 4660 17682
rect 4620 17332 4672 17338
rect 4620 17274 4672 17280
rect 4908 17066 4936 17818
rect 5000 17746 5028 19178
rect 5092 18970 5120 19178
rect 5080 18964 5132 18970
rect 5080 18906 5132 18912
rect 5080 18216 5132 18222
rect 5080 18158 5132 18164
rect 5092 17814 5120 18158
rect 5080 17808 5132 17814
rect 5080 17750 5132 17756
rect 4988 17740 5040 17746
rect 4988 17682 5040 17688
rect 5368 17610 5396 23530
rect 5460 23322 5488 24550
rect 5552 23662 5580 29990
rect 5828 29850 5856 29990
rect 5920 29850 5948 30126
rect 6736 30048 6788 30054
rect 6736 29990 6788 29996
rect 5816 29844 5868 29850
rect 5816 29786 5868 29792
rect 5908 29844 5960 29850
rect 5908 29786 5960 29792
rect 6748 29782 6776 29990
rect 6736 29776 6788 29782
rect 6736 29718 6788 29724
rect 6368 29640 6420 29646
rect 6368 29582 6420 29588
rect 5908 29232 5960 29238
rect 5908 29174 5960 29180
rect 5920 28626 5948 29174
rect 6380 29102 6408 29582
rect 6458 29472 6514 29481
rect 6458 29407 6514 29416
rect 6472 29306 6500 29407
rect 6460 29300 6512 29306
rect 6460 29242 6512 29248
rect 6368 29096 6420 29102
rect 6368 29038 6420 29044
rect 6644 29096 6696 29102
rect 6644 29038 6696 29044
rect 6656 28762 6684 29038
rect 6644 28756 6696 28762
rect 6644 28698 6696 28704
rect 5908 28620 5960 28626
rect 5908 28562 5960 28568
rect 6840 28558 6868 30126
rect 7472 30116 7524 30122
rect 7472 30058 7524 30064
rect 8024 30116 8076 30122
rect 8024 30058 8076 30064
rect 7114 29948 7422 29957
rect 7114 29946 7120 29948
rect 7176 29946 7200 29948
rect 7256 29946 7280 29948
rect 7336 29946 7360 29948
rect 7416 29946 7422 29948
rect 7176 29894 7178 29946
rect 7358 29894 7360 29946
rect 7114 29892 7120 29894
rect 7176 29892 7200 29894
rect 7256 29892 7280 29894
rect 7336 29892 7360 29894
rect 7416 29892 7422 29894
rect 7114 29883 7422 29892
rect 7484 29850 7512 30058
rect 7656 30048 7708 30054
rect 7656 29990 7708 29996
rect 7472 29844 7524 29850
rect 7472 29786 7524 29792
rect 6920 29708 6972 29714
rect 6920 29650 6972 29656
rect 7104 29708 7156 29714
rect 7104 29650 7156 29656
rect 6932 29306 6960 29650
rect 7012 29640 7064 29646
rect 7012 29582 7064 29588
rect 6920 29300 6972 29306
rect 6920 29242 6972 29248
rect 7024 29050 7052 29582
rect 7116 29510 7144 29650
rect 7668 29646 7696 29990
rect 7932 29844 7984 29850
rect 7932 29786 7984 29792
rect 7840 29776 7892 29782
rect 7840 29718 7892 29724
rect 7748 29708 7800 29714
rect 7748 29650 7800 29656
rect 7196 29640 7248 29646
rect 7196 29582 7248 29588
rect 7656 29640 7708 29646
rect 7656 29582 7708 29588
rect 7104 29504 7156 29510
rect 7104 29446 7156 29452
rect 7208 29306 7236 29582
rect 7564 29504 7616 29510
rect 7564 29446 7616 29452
rect 7196 29300 7248 29306
rect 7196 29242 7248 29248
rect 6932 29022 7052 29050
rect 7472 29028 7524 29034
rect 6828 28552 6880 28558
rect 6828 28494 6880 28500
rect 6552 28144 6604 28150
rect 6552 28086 6604 28092
rect 6092 27124 6144 27130
rect 6092 27066 6144 27072
rect 5816 26852 5868 26858
rect 5816 26794 5868 26800
rect 5828 26586 5856 26794
rect 5816 26580 5868 26586
rect 5816 26522 5868 26528
rect 5632 26240 5684 26246
rect 5632 26182 5684 26188
rect 5644 25702 5672 26182
rect 5632 25696 5684 25702
rect 5632 25638 5684 25644
rect 5724 25696 5776 25702
rect 5724 25638 5776 25644
rect 5644 24682 5672 25638
rect 5736 24886 5764 25638
rect 5724 24880 5776 24886
rect 5724 24822 5776 24828
rect 6104 24834 6132 27066
rect 6184 26376 6236 26382
rect 6184 26318 6236 26324
rect 6196 25702 6224 26318
rect 6184 25696 6236 25702
rect 6184 25638 6236 25644
rect 6460 25696 6512 25702
rect 6460 25638 6512 25644
rect 6472 25498 6500 25638
rect 6460 25492 6512 25498
rect 6460 25434 6512 25440
rect 6460 24880 6512 24886
rect 6366 24848 6422 24857
rect 6104 24806 6366 24834
rect 5632 24676 5684 24682
rect 5632 24618 5684 24624
rect 6104 24342 6132 24806
rect 6460 24822 6512 24828
rect 6366 24783 6422 24792
rect 6366 24712 6422 24721
rect 6196 24670 6366 24698
rect 6092 24336 6144 24342
rect 6092 24278 6144 24284
rect 6196 24274 6224 24670
rect 6366 24647 6422 24656
rect 6366 24304 6422 24313
rect 6184 24268 6236 24274
rect 6472 24274 6500 24822
rect 6564 24290 6592 28086
rect 6736 28008 6788 28014
rect 6736 27950 6788 27956
rect 6748 27130 6776 27950
rect 6840 27538 6868 28494
rect 6932 28490 6960 29022
rect 7472 28970 7524 28976
rect 7012 28960 7064 28966
rect 7012 28902 7064 28908
rect 6920 28484 6972 28490
rect 6920 28426 6972 28432
rect 7024 28218 7052 28902
rect 7114 28860 7422 28869
rect 7114 28858 7120 28860
rect 7176 28858 7200 28860
rect 7256 28858 7280 28860
rect 7336 28858 7360 28860
rect 7416 28858 7422 28860
rect 7176 28806 7178 28858
rect 7358 28806 7360 28858
rect 7114 28804 7120 28806
rect 7176 28804 7200 28806
rect 7256 28804 7280 28806
rect 7336 28804 7360 28806
rect 7416 28804 7422 28806
rect 7114 28795 7422 28804
rect 7484 28762 7512 28970
rect 7576 28762 7604 29446
rect 7668 29306 7696 29582
rect 7760 29578 7788 29650
rect 7748 29572 7800 29578
rect 7748 29514 7800 29520
rect 7760 29481 7788 29514
rect 7746 29472 7802 29481
rect 7746 29407 7802 29416
rect 7656 29300 7708 29306
rect 7656 29242 7708 29248
rect 7656 29028 7708 29034
rect 7656 28970 7708 28976
rect 7288 28756 7340 28762
rect 7288 28698 7340 28704
rect 7472 28756 7524 28762
rect 7472 28698 7524 28704
rect 7564 28756 7616 28762
rect 7564 28698 7616 28704
rect 7300 28642 7328 28698
rect 7300 28626 7604 28642
rect 7196 28620 7248 28626
rect 7300 28620 7616 28626
rect 7300 28614 7564 28620
rect 7196 28562 7248 28568
rect 7564 28562 7616 28568
rect 7208 28506 7236 28562
rect 7668 28506 7696 28970
rect 7748 28960 7800 28966
rect 7748 28902 7800 28908
rect 7760 28626 7788 28902
rect 7748 28620 7800 28626
rect 7748 28562 7800 28568
rect 7208 28478 7696 28506
rect 7012 28212 7064 28218
rect 7012 28154 7064 28160
rect 7852 27946 7880 29718
rect 7944 29102 7972 29786
rect 8036 29102 8064 30058
rect 8300 29708 8352 29714
rect 8300 29650 8352 29656
rect 8312 29238 8340 29650
rect 8496 29306 8524 30534
rect 8668 30116 8720 30122
rect 8668 30058 8720 30064
rect 8680 29306 8708 30058
rect 8772 30054 8800 30534
rect 8760 30048 8812 30054
rect 8760 29990 8812 29996
rect 9588 30048 9640 30054
rect 9588 29990 9640 29996
rect 8772 29714 8800 29990
rect 9600 29782 9628 29990
rect 9588 29776 9640 29782
rect 9588 29718 9640 29724
rect 8760 29708 8812 29714
rect 8760 29650 8812 29656
rect 8760 29504 8812 29510
rect 8760 29446 8812 29452
rect 9404 29504 9456 29510
rect 9404 29446 9456 29452
rect 8484 29300 8536 29306
rect 8484 29242 8536 29248
rect 8668 29300 8720 29306
rect 8668 29242 8720 29248
rect 8300 29232 8352 29238
rect 8300 29174 8352 29180
rect 8772 29102 8800 29446
rect 9416 29306 9444 29446
rect 9692 29306 9720 30738
rect 9876 29782 9904 30738
rect 10232 30728 10284 30734
rect 10232 30670 10284 30676
rect 11244 30728 11296 30734
rect 11244 30670 11296 30676
rect 11796 30728 11848 30734
rect 11796 30670 11848 30676
rect 12440 30728 12492 30734
rect 12440 30670 12492 30676
rect 10244 30054 10272 30670
rect 11060 30660 11112 30666
rect 11060 30602 11112 30608
rect 10472 30492 10780 30501
rect 10472 30490 10478 30492
rect 10534 30490 10558 30492
rect 10614 30490 10638 30492
rect 10694 30490 10718 30492
rect 10774 30490 10780 30492
rect 10534 30438 10536 30490
rect 10716 30438 10718 30490
rect 10472 30436 10478 30438
rect 10534 30436 10558 30438
rect 10614 30436 10638 30438
rect 10694 30436 10718 30438
rect 10774 30436 10780 30438
rect 10472 30427 10780 30436
rect 10968 30184 11020 30190
rect 10968 30126 11020 30132
rect 10232 30048 10284 30054
rect 10232 29990 10284 29996
rect 9864 29776 9916 29782
rect 9864 29718 9916 29724
rect 10232 29708 10284 29714
rect 10232 29650 10284 29656
rect 10324 29708 10376 29714
rect 10324 29650 10376 29656
rect 10244 29306 10272 29650
rect 10336 29306 10364 29650
rect 10980 29646 11008 30126
rect 11072 30122 11100 30602
rect 11060 30116 11112 30122
rect 11060 30058 11112 30064
rect 11152 30048 11204 30054
rect 11152 29990 11204 29996
rect 10968 29640 11020 29646
rect 10968 29582 11020 29588
rect 10472 29404 10780 29413
rect 10472 29402 10478 29404
rect 10534 29402 10558 29404
rect 10614 29402 10638 29404
rect 10694 29402 10718 29404
rect 10774 29402 10780 29404
rect 10534 29350 10536 29402
rect 10716 29350 10718 29402
rect 10472 29348 10478 29350
rect 10534 29348 10558 29350
rect 10614 29348 10638 29350
rect 10694 29348 10718 29350
rect 10774 29348 10780 29350
rect 10472 29339 10780 29348
rect 9404 29300 9456 29306
rect 9404 29242 9456 29248
rect 9496 29300 9548 29306
rect 9496 29242 9548 29248
rect 9680 29300 9732 29306
rect 9680 29242 9732 29248
rect 10232 29300 10284 29306
rect 10232 29242 10284 29248
rect 10324 29300 10376 29306
rect 10324 29242 10376 29248
rect 7932 29096 7984 29102
rect 7932 29038 7984 29044
rect 8024 29096 8076 29102
rect 8024 29038 8076 29044
rect 8760 29096 8812 29102
rect 8760 29038 8812 29044
rect 7944 28490 7972 29038
rect 8392 29028 8444 29034
rect 8392 28970 8444 28976
rect 7932 28484 7984 28490
rect 7932 28426 7984 28432
rect 8024 28008 8076 28014
rect 8024 27950 8076 27956
rect 7564 27940 7616 27946
rect 7564 27882 7616 27888
rect 7840 27940 7892 27946
rect 7840 27882 7892 27888
rect 7114 27772 7422 27781
rect 7114 27770 7120 27772
rect 7176 27770 7200 27772
rect 7256 27770 7280 27772
rect 7336 27770 7360 27772
rect 7416 27770 7422 27772
rect 7176 27718 7178 27770
rect 7358 27718 7360 27770
rect 7114 27716 7120 27718
rect 7176 27716 7200 27718
rect 7256 27716 7280 27718
rect 7336 27716 7360 27718
rect 7416 27716 7422 27718
rect 7114 27707 7422 27716
rect 6828 27532 6880 27538
rect 6828 27474 6880 27480
rect 6736 27124 6788 27130
rect 6736 27066 6788 27072
rect 6840 25294 6868 27474
rect 7288 27328 7340 27334
rect 7288 27270 7340 27276
rect 7300 26994 7328 27270
rect 7472 27056 7524 27062
rect 7472 26998 7524 27004
rect 7288 26988 7340 26994
rect 7288 26930 7340 26936
rect 6920 26784 6972 26790
rect 6920 26726 6972 26732
rect 7012 26784 7064 26790
rect 7012 26726 7064 26732
rect 6932 26246 6960 26726
rect 7024 26586 7052 26726
rect 7114 26684 7422 26693
rect 7114 26682 7120 26684
rect 7176 26682 7200 26684
rect 7256 26682 7280 26684
rect 7336 26682 7360 26684
rect 7416 26682 7422 26684
rect 7176 26630 7178 26682
rect 7358 26630 7360 26682
rect 7114 26628 7120 26630
rect 7176 26628 7200 26630
rect 7256 26628 7280 26630
rect 7336 26628 7360 26630
rect 7416 26628 7422 26630
rect 7114 26619 7422 26628
rect 7484 26586 7512 26998
rect 7012 26580 7064 26586
rect 7012 26522 7064 26528
rect 7472 26580 7524 26586
rect 7472 26522 7524 26528
rect 7576 26450 7604 27882
rect 7748 27872 7800 27878
rect 7748 27814 7800 27820
rect 7932 27872 7984 27878
rect 7932 27814 7984 27820
rect 7760 26994 7788 27814
rect 7840 27532 7892 27538
rect 7840 27474 7892 27480
rect 7852 26994 7880 27474
rect 7944 27334 7972 27814
rect 8036 27538 8064 27950
rect 8404 27946 8432 28970
rect 8772 28082 8800 29038
rect 8944 29028 8996 29034
rect 8944 28970 8996 28976
rect 8956 28778 8984 28970
rect 9508 28966 9536 29242
rect 9496 28960 9548 28966
rect 9496 28902 9548 28908
rect 9680 28960 9732 28966
rect 9680 28902 9732 28908
rect 8956 28750 9076 28778
rect 8944 28620 8996 28626
rect 8944 28562 8996 28568
rect 8760 28076 8812 28082
rect 8760 28018 8812 28024
rect 8392 27940 8444 27946
rect 8392 27882 8444 27888
rect 8404 27538 8432 27882
rect 8576 27872 8628 27878
rect 8576 27814 8628 27820
rect 8024 27532 8076 27538
rect 8024 27474 8076 27480
rect 8392 27532 8444 27538
rect 8392 27474 8444 27480
rect 8036 27402 8064 27474
rect 8024 27396 8076 27402
rect 8024 27338 8076 27344
rect 7932 27328 7984 27334
rect 7932 27270 7984 27276
rect 7748 26988 7800 26994
rect 7748 26930 7800 26936
rect 7840 26988 7892 26994
rect 7840 26930 7892 26936
rect 7656 26784 7708 26790
rect 7656 26726 7708 26732
rect 7104 26444 7156 26450
rect 7104 26386 7156 26392
rect 7564 26444 7616 26450
rect 7564 26386 7616 26392
rect 7012 26376 7064 26382
rect 7012 26318 7064 26324
rect 6920 26240 6972 26246
rect 6920 26182 6972 26188
rect 7024 25974 7052 26318
rect 7116 26042 7144 26386
rect 7104 26036 7156 26042
rect 7104 25978 7156 25984
rect 7012 25968 7064 25974
rect 7012 25910 7064 25916
rect 7668 25906 7696 26726
rect 8404 26450 8432 27474
rect 8588 27402 8616 27814
rect 8772 27538 8800 28018
rect 8852 28008 8904 28014
rect 8852 27950 8904 27956
rect 8760 27532 8812 27538
rect 8760 27474 8812 27480
rect 8864 27470 8892 27950
rect 8956 27674 8984 28562
rect 8944 27668 8996 27674
rect 8944 27610 8996 27616
rect 9048 27554 9076 28750
rect 9692 28422 9720 28902
rect 10980 28558 11008 29582
rect 11164 29306 11192 29990
rect 11256 29510 11284 30670
rect 11808 29850 11836 30670
rect 12164 30592 12216 30598
rect 12164 30534 12216 30540
rect 11796 29844 11848 29850
rect 11796 29786 11848 29792
rect 12176 29646 12204 30534
rect 12452 29782 12480 30670
rect 12624 30592 12676 30598
rect 12624 30534 12676 30540
rect 12636 30258 12664 30534
rect 12624 30252 12676 30258
rect 12624 30194 12676 30200
rect 12728 29850 12756 30738
rect 13268 30388 13320 30394
rect 13268 30330 13320 30336
rect 12992 30320 13044 30326
rect 12992 30262 13044 30268
rect 12808 30252 12860 30258
rect 12808 30194 12860 30200
rect 12716 29844 12768 29850
rect 12716 29786 12768 29792
rect 12440 29776 12492 29782
rect 12440 29718 12492 29724
rect 12164 29640 12216 29646
rect 11978 29608 12034 29617
rect 12164 29582 12216 29588
rect 12440 29640 12492 29646
rect 12440 29582 12492 29588
rect 11978 29543 12034 29552
rect 11244 29504 11296 29510
rect 11244 29446 11296 29452
rect 11152 29300 11204 29306
rect 11152 29242 11204 29248
rect 10968 28552 11020 28558
rect 10968 28494 11020 28500
rect 9680 28416 9732 28422
rect 9680 28358 9732 28364
rect 10140 28416 10192 28422
rect 10140 28358 10192 28364
rect 9692 28218 9720 28358
rect 9680 28212 9732 28218
rect 9680 28154 9732 28160
rect 9220 28076 9272 28082
rect 9220 28018 9272 28024
rect 8956 27526 9076 27554
rect 8852 27464 8904 27470
rect 8852 27406 8904 27412
rect 8576 27396 8628 27402
rect 8576 27338 8628 27344
rect 8588 26926 8616 27338
rect 8864 27130 8892 27406
rect 8852 27124 8904 27130
rect 8852 27066 8904 27072
rect 8576 26920 8628 26926
rect 8576 26862 8628 26868
rect 8392 26444 8444 26450
rect 8392 26386 8444 26392
rect 8404 26314 8432 26386
rect 8484 26376 8536 26382
rect 8484 26318 8536 26324
rect 7748 26308 7800 26314
rect 7748 26250 7800 26256
rect 8392 26308 8444 26314
rect 8392 26250 8444 26256
rect 7656 25900 7708 25906
rect 7656 25842 7708 25848
rect 7114 25596 7422 25605
rect 7114 25594 7120 25596
rect 7176 25594 7200 25596
rect 7256 25594 7280 25596
rect 7336 25594 7360 25596
rect 7416 25594 7422 25596
rect 7176 25542 7178 25594
rect 7358 25542 7360 25594
rect 7114 25540 7120 25542
rect 7176 25540 7200 25542
rect 7256 25540 7280 25542
rect 7336 25540 7360 25542
rect 7416 25540 7422 25542
rect 7114 25531 7422 25540
rect 6828 25288 6880 25294
rect 6828 25230 6880 25236
rect 6920 25152 6972 25158
rect 6920 25094 6972 25100
rect 6932 24954 6960 25094
rect 6920 24948 6972 24954
rect 6920 24890 6972 24896
rect 6920 24744 6972 24750
rect 7564 24744 7616 24750
rect 6972 24692 7052 24698
rect 6920 24686 7052 24692
rect 7564 24686 7616 24692
rect 7654 24712 7710 24721
rect 6932 24670 7052 24686
rect 6828 24608 6880 24614
rect 6828 24550 6880 24556
rect 6366 24239 6422 24248
rect 6460 24268 6512 24274
rect 6184 24210 6236 24216
rect 6380 24070 6408 24239
rect 6564 24262 6776 24290
rect 6840 24274 6868 24550
rect 7024 24410 7052 24670
rect 7472 24608 7524 24614
rect 7472 24550 7524 24556
rect 7114 24508 7422 24517
rect 7114 24506 7120 24508
rect 7176 24506 7200 24508
rect 7256 24506 7280 24508
rect 7336 24506 7360 24508
rect 7416 24506 7422 24508
rect 7176 24454 7178 24506
rect 7358 24454 7360 24506
rect 7114 24452 7120 24454
rect 7176 24452 7200 24454
rect 7256 24452 7280 24454
rect 7336 24452 7360 24454
rect 7416 24452 7422 24454
rect 7114 24443 7422 24452
rect 7012 24404 7064 24410
rect 7012 24346 7064 24352
rect 7024 24274 7052 24346
rect 6460 24210 6512 24216
rect 6552 24132 6604 24138
rect 6552 24074 6604 24080
rect 6368 24064 6420 24070
rect 6368 24006 6420 24012
rect 6460 24064 6512 24070
rect 6460 24006 6512 24012
rect 6472 23866 6500 24006
rect 6564 23866 6592 24074
rect 6460 23860 6512 23866
rect 6460 23802 6512 23808
rect 6552 23860 6604 23866
rect 6552 23802 6604 23808
rect 5540 23656 5592 23662
rect 5540 23598 5592 23604
rect 5448 23316 5500 23322
rect 5448 23258 5500 23264
rect 6092 23180 6144 23186
rect 6092 23122 6144 23128
rect 5540 22976 5592 22982
rect 5540 22918 5592 22924
rect 5448 22772 5500 22778
rect 5448 22714 5500 22720
rect 5460 21962 5488 22714
rect 5552 22574 5580 22918
rect 5540 22568 5592 22574
rect 5540 22510 5592 22516
rect 5816 22568 5868 22574
rect 5816 22510 5868 22516
rect 5552 22098 5580 22510
rect 5632 22432 5684 22438
rect 5632 22374 5684 22380
rect 5540 22092 5592 22098
rect 5644 22094 5672 22374
rect 5828 22234 5856 22510
rect 5816 22228 5868 22234
rect 5816 22170 5868 22176
rect 5644 22066 5856 22094
rect 5540 22034 5592 22040
rect 5448 21956 5500 21962
rect 5448 21898 5500 21904
rect 5540 21548 5592 21554
rect 5540 21490 5592 21496
rect 5448 21412 5500 21418
rect 5448 21354 5500 21360
rect 5460 19854 5488 21354
rect 5552 20806 5580 21490
rect 5828 21010 5856 22066
rect 6000 22024 6052 22030
rect 6000 21966 6052 21972
rect 6012 21690 6040 21966
rect 6104 21894 6132 23122
rect 6276 22976 6328 22982
rect 6276 22918 6328 22924
rect 6288 22642 6316 22918
rect 6644 22704 6696 22710
rect 6644 22646 6696 22652
rect 6276 22636 6328 22642
rect 6328 22596 6408 22624
rect 6276 22578 6328 22584
rect 6276 22500 6328 22506
rect 6276 22442 6328 22448
rect 6288 22234 6316 22442
rect 6380 22234 6408 22596
rect 6552 22432 6604 22438
rect 6552 22374 6604 22380
rect 6564 22234 6592 22374
rect 6276 22228 6328 22234
rect 6276 22170 6328 22176
rect 6368 22228 6420 22234
rect 6368 22170 6420 22176
rect 6552 22228 6604 22234
rect 6552 22170 6604 22176
rect 6656 22094 6684 22646
rect 6748 22098 6776 24262
rect 6828 24268 6880 24274
rect 6828 24210 6880 24216
rect 7012 24268 7064 24274
rect 7012 24210 7064 24216
rect 7484 24206 7512 24550
rect 7472 24200 7524 24206
rect 7472 24142 7524 24148
rect 6920 24064 6972 24070
rect 6918 24032 6920 24041
rect 7380 24064 7432 24070
rect 6972 24032 6974 24041
rect 7380 24006 7432 24012
rect 6918 23967 6974 23976
rect 6920 23860 6972 23866
rect 6920 23802 6972 23808
rect 6932 23322 6960 23802
rect 7392 23662 7420 24006
rect 7380 23656 7432 23662
rect 7484 23644 7512 24142
rect 7576 23798 7604 24686
rect 7654 24647 7656 24656
rect 7708 24647 7710 24656
rect 7656 24618 7708 24624
rect 7656 24404 7708 24410
rect 7656 24346 7708 24352
rect 7668 24070 7696 24346
rect 7656 24064 7708 24070
rect 7656 24006 7708 24012
rect 7564 23792 7616 23798
rect 7564 23734 7616 23740
rect 7564 23656 7616 23662
rect 7484 23616 7564 23644
rect 7380 23598 7432 23604
rect 7564 23598 7616 23604
rect 7012 23520 7064 23526
rect 7012 23462 7064 23468
rect 6920 23316 6972 23322
rect 6920 23258 6972 23264
rect 7024 23186 7052 23462
rect 7114 23420 7422 23429
rect 7114 23418 7120 23420
rect 7176 23418 7200 23420
rect 7256 23418 7280 23420
rect 7336 23418 7360 23420
rect 7416 23418 7422 23420
rect 7176 23366 7178 23418
rect 7358 23366 7360 23418
rect 7114 23364 7120 23366
rect 7176 23364 7200 23366
rect 7256 23364 7280 23366
rect 7336 23364 7360 23366
rect 7416 23364 7422 23366
rect 7114 23355 7422 23364
rect 7760 23254 7788 26250
rect 8024 26240 8076 26246
rect 8024 26182 8076 26188
rect 8036 25430 8064 26182
rect 8024 25424 8076 25430
rect 8024 25366 8076 25372
rect 8114 24848 8170 24857
rect 8036 24806 8114 24834
rect 7840 24744 7892 24750
rect 7840 24686 7892 24692
rect 7852 24041 7880 24686
rect 7930 24304 7986 24313
rect 7930 24239 7932 24248
rect 7984 24239 7986 24248
rect 7932 24210 7984 24216
rect 7932 24132 7984 24138
rect 7932 24074 7984 24080
rect 7838 24032 7894 24041
rect 7838 23967 7894 23976
rect 7852 23662 7880 23967
rect 7944 23662 7972 24074
rect 7840 23656 7892 23662
rect 7840 23598 7892 23604
rect 7932 23656 7984 23662
rect 7932 23598 7984 23604
rect 7748 23248 7800 23254
rect 7748 23190 7800 23196
rect 6828 23180 6880 23186
rect 6828 23122 6880 23128
rect 7012 23180 7064 23186
rect 7012 23122 7064 23128
rect 6564 22066 6684 22094
rect 6736 22092 6788 22098
rect 6092 21888 6144 21894
rect 6092 21830 6144 21836
rect 6000 21684 6052 21690
rect 6000 21626 6052 21632
rect 5816 21004 5868 21010
rect 5816 20946 5868 20952
rect 5908 21004 5960 21010
rect 5908 20946 5960 20952
rect 5540 20800 5592 20806
rect 5540 20742 5592 20748
rect 5552 20534 5580 20742
rect 5540 20528 5592 20534
rect 5540 20470 5592 20476
rect 5448 19848 5500 19854
rect 5448 19790 5500 19796
rect 5460 18834 5488 19790
rect 5448 18828 5500 18834
rect 5448 18770 5500 18776
rect 5828 18698 5856 20946
rect 5920 19242 5948 20946
rect 6276 20392 6328 20398
rect 6276 20334 6328 20340
rect 6288 19310 6316 20334
rect 6564 19990 6592 22066
rect 6736 22034 6788 22040
rect 6840 21978 6868 23122
rect 7024 22658 7052 23122
rect 7656 23044 7708 23050
rect 7656 22986 7708 22992
rect 7472 22976 7524 22982
rect 7472 22918 7524 22924
rect 7024 22630 7144 22658
rect 7116 22574 7144 22630
rect 7012 22568 7064 22574
rect 7012 22510 7064 22516
rect 7104 22568 7156 22574
rect 7104 22510 7156 22516
rect 7484 22522 7512 22918
rect 7024 22030 7052 22510
rect 7484 22494 7604 22522
rect 7472 22432 7524 22438
rect 7472 22374 7524 22380
rect 7114 22332 7422 22341
rect 7114 22330 7120 22332
rect 7176 22330 7200 22332
rect 7256 22330 7280 22332
rect 7336 22330 7360 22332
rect 7416 22330 7422 22332
rect 7176 22278 7178 22330
rect 7358 22278 7360 22330
rect 7114 22276 7120 22278
rect 7176 22276 7200 22278
rect 7256 22276 7280 22278
rect 7336 22276 7360 22278
rect 7416 22276 7422 22278
rect 7114 22267 7422 22276
rect 7484 22234 7512 22374
rect 7472 22228 7524 22234
rect 7472 22170 7524 22176
rect 7576 22098 7604 22494
rect 7668 22234 7696 22986
rect 7760 22574 7788 23190
rect 7932 22636 7984 22642
rect 7932 22578 7984 22584
rect 7748 22568 7800 22574
rect 7748 22510 7800 22516
rect 7840 22500 7892 22506
rect 7840 22442 7892 22448
rect 7656 22228 7708 22234
rect 7656 22170 7708 22176
rect 7564 22092 7616 22098
rect 7564 22034 7616 22040
rect 7748 22092 7800 22098
rect 7748 22034 7800 22040
rect 6656 21962 6868 21978
rect 7012 22024 7064 22030
rect 7012 21966 7064 21972
rect 6644 21956 6868 21962
rect 6696 21950 6868 21956
rect 6920 21956 6972 21962
rect 6644 21898 6696 21904
rect 6920 21898 6972 21904
rect 6552 19984 6604 19990
rect 6552 19926 6604 19932
rect 6368 19712 6420 19718
rect 6368 19654 6420 19660
rect 6092 19304 6144 19310
rect 6092 19246 6144 19252
rect 6276 19304 6328 19310
rect 6276 19246 6328 19252
rect 5908 19236 5960 19242
rect 5908 19178 5960 19184
rect 5816 18692 5868 18698
rect 5816 18634 5868 18640
rect 5828 18222 5856 18634
rect 6104 18630 6132 19246
rect 6288 18834 6316 19246
rect 6276 18828 6328 18834
rect 6276 18770 6328 18776
rect 6092 18624 6144 18630
rect 6092 18566 6144 18572
rect 5816 18216 5868 18222
rect 5816 18158 5868 18164
rect 5356 17604 5408 17610
rect 5356 17546 5408 17552
rect 6104 17134 6132 18566
rect 6288 17746 6316 18770
rect 6380 18222 6408 19654
rect 6460 18828 6512 18834
rect 6460 18770 6512 18776
rect 6472 18426 6500 18770
rect 6460 18420 6512 18426
rect 6460 18362 6512 18368
rect 6368 18216 6420 18222
rect 6368 18158 6420 18164
rect 6276 17740 6328 17746
rect 6276 17682 6328 17688
rect 6288 17202 6316 17682
rect 6276 17196 6328 17202
rect 6276 17138 6328 17144
rect 6092 17128 6144 17134
rect 6092 17070 6144 17076
rect 4896 17060 4948 17066
rect 4896 17002 4948 17008
rect 4436 16788 4488 16794
rect 4436 16730 4488 16736
rect 6564 16590 6592 19926
rect 6932 18630 6960 21898
rect 7024 21690 7052 21966
rect 7760 21690 7788 22034
rect 7012 21684 7064 21690
rect 7012 21626 7064 21632
rect 7748 21684 7800 21690
rect 7748 21626 7800 21632
rect 7748 21548 7800 21554
rect 7748 21490 7800 21496
rect 7012 21480 7064 21486
rect 7012 21422 7064 21428
rect 7024 21146 7052 21422
rect 7564 21412 7616 21418
rect 7564 21354 7616 21360
rect 7472 21344 7524 21350
rect 7472 21286 7524 21292
rect 7114 21244 7422 21253
rect 7114 21242 7120 21244
rect 7176 21242 7200 21244
rect 7256 21242 7280 21244
rect 7336 21242 7360 21244
rect 7416 21242 7422 21244
rect 7176 21190 7178 21242
rect 7358 21190 7360 21242
rect 7114 21188 7120 21190
rect 7176 21188 7200 21190
rect 7256 21188 7280 21190
rect 7336 21188 7360 21190
rect 7416 21188 7422 21190
rect 7114 21179 7422 21188
rect 7484 21146 7512 21286
rect 7012 21140 7064 21146
rect 7012 21082 7064 21088
rect 7472 21140 7524 21146
rect 7472 21082 7524 21088
rect 7576 21026 7604 21354
rect 7656 21344 7708 21350
rect 7656 21286 7708 21292
rect 7484 21010 7604 21026
rect 7472 21004 7604 21010
rect 7524 20998 7604 21004
rect 7472 20946 7524 20952
rect 7012 20868 7064 20874
rect 7012 20810 7064 20816
rect 7024 19718 7052 20810
rect 7484 20602 7512 20946
rect 7668 20942 7696 21286
rect 7656 20936 7708 20942
rect 7656 20878 7708 20884
rect 7472 20596 7524 20602
rect 7472 20538 7524 20544
rect 7114 20156 7422 20165
rect 7114 20154 7120 20156
rect 7176 20154 7200 20156
rect 7256 20154 7280 20156
rect 7336 20154 7360 20156
rect 7416 20154 7422 20156
rect 7176 20102 7178 20154
rect 7358 20102 7360 20154
rect 7114 20100 7120 20102
rect 7176 20100 7200 20102
rect 7256 20100 7280 20102
rect 7336 20100 7360 20102
rect 7416 20100 7422 20102
rect 7114 20091 7422 20100
rect 7668 20058 7696 20878
rect 7760 20398 7788 21490
rect 7852 21146 7880 22442
rect 7944 22098 7972 22578
rect 7932 22092 7984 22098
rect 8036 22094 8064 24806
rect 8114 24783 8170 24792
rect 8116 24200 8168 24206
rect 8116 24142 8168 24148
rect 8128 23866 8156 24142
rect 8116 23860 8168 23866
rect 8116 23802 8168 23808
rect 8208 23656 8260 23662
rect 8208 23598 8260 23604
rect 8220 23322 8248 23598
rect 8208 23316 8260 23322
rect 8208 23258 8260 23264
rect 8404 22778 8432 26250
rect 8392 22772 8444 22778
rect 8392 22714 8444 22720
rect 8036 22066 8156 22094
rect 7932 22034 7984 22040
rect 8024 22024 8076 22030
rect 8024 21966 8076 21972
rect 7932 21344 7984 21350
rect 7932 21286 7984 21292
rect 7840 21140 7892 21146
rect 7840 21082 7892 21088
rect 7944 20806 7972 21286
rect 7840 20800 7892 20806
rect 7840 20742 7892 20748
rect 7932 20800 7984 20806
rect 7932 20742 7984 20748
rect 7748 20392 7800 20398
rect 7748 20334 7800 20340
rect 7656 20052 7708 20058
rect 7656 19994 7708 20000
rect 7852 19922 7880 20742
rect 7944 20602 7972 20742
rect 7932 20596 7984 20602
rect 7932 20538 7984 20544
rect 7840 19916 7892 19922
rect 7840 19858 7892 19864
rect 7564 19848 7616 19854
rect 7564 19790 7616 19796
rect 7012 19712 7064 19718
rect 7012 19654 7064 19660
rect 7114 19068 7422 19077
rect 7114 19066 7120 19068
rect 7176 19066 7200 19068
rect 7256 19066 7280 19068
rect 7336 19066 7360 19068
rect 7416 19066 7422 19068
rect 7176 19014 7178 19066
rect 7358 19014 7360 19066
rect 7114 19012 7120 19014
rect 7176 19012 7200 19014
rect 7256 19012 7280 19014
rect 7336 19012 7360 19014
rect 7416 19012 7422 19014
rect 7114 19003 7422 19012
rect 7576 18970 7604 19790
rect 8036 19310 8064 21966
rect 8128 19394 8156 22066
rect 8208 21956 8260 21962
rect 8208 21898 8260 21904
rect 8220 21690 8248 21898
rect 8208 21684 8260 21690
rect 8208 21626 8260 21632
rect 8496 20058 8524 26318
rect 8760 26240 8812 26246
rect 8760 26182 8812 26188
rect 8772 25770 8800 26182
rect 8760 25764 8812 25770
rect 8760 25706 8812 25712
rect 8668 24676 8720 24682
rect 8668 24618 8720 24624
rect 8680 24410 8708 24618
rect 8852 24608 8904 24614
rect 8852 24550 8904 24556
rect 8668 24404 8720 24410
rect 8668 24346 8720 24352
rect 8864 24274 8892 24550
rect 8956 24274 8984 27526
rect 9036 27124 9088 27130
rect 9036 27066 9088 27072
rect 9048 26450 9076 27066
rect 9036 26444 9088 26450
rect 9036 26386 9088 26392
rect 9048 26314 9076 26386
rect 9036 26308 9088 26314
rect 9036 26250 9088 26256
rect 9036 25288 9088 25294
rect 9036 25230 9088 25236
rect 9048 24954 9076 25230
rect 9036 24948 9088 24954
rect 9036 24890 9088 24896
rect 8852 24268 8904 24274
rect 8852 24210 8904 24216
rect 8944 24268 8996 24274
rect 8944 24210 8996 24216
rect 8576 24200 8628 24206
rect 8576 24142 8628 24148
rect 8588 23662 8616 24142
rect 8864 23662 8892 24210
rect 8576 23656 8628 23662
rect 8576 23598 8628 23604
rect 8852 23656 8904 23662
rect 8852 23598 8904 23604
rect 8760 22092 8812 22098
rect 8760 22034 8812 22040
rect 8772 21690 8800 22034
rect 8760 21684 8812 21690
rect 8760 21626 8812 21632
rect 8864 21486 8892 23598
rect 9036 23520 9088 23526
rect 9036 23462 9088 23468
rect 9048 23254 9076 23462
rect 9036 23248 9088 23254
rect 9036 23190 9088 23196
rect 8852 21480 8904 21486
rect 8852 21422 8904 21428
rect 8576 20596 8628 20602
rect 8576 20538 8628 20544
rect 8484 20052 8536 20058
rect 8484 19994 8536 20000
rect 8588 19854 8616 20538
rect 8576 19848 8628 19854
rect 8576 19790 8628 19796
rect 8128 19366 8248 19394
rect 8024 19304 8076 19310
rect 8024 19246 8076 19252
rect 8220 19174 8248 19366
rect 8484 19304 8536 19310
rect 8484 19246 8536 19252
rect 8208 19168 8260 19174
rect 8208 19110 8260 19116
rect 8392 19168 8444 19174
rect 8392 19110 8444 19116
rect 7564 18964 7616 18970
rect 7564 18906 7616 18912
rect 8220 18698 8248 19110
rect 8208 18692 8260 18698
rect 8208 18634 8260 18640
rect 8300 18692 8352 18698
rect 8300 18634 8352 18640
rect 6920 18624 6972 18630
rect 6920 18566 6972 18572
rect 7840 18624 7892 18630
rect 7840 18566 7892 18572
rect 6932 18290 6960 18566
rect 7852 18358 7880 18566
rect 7840 18352 7892 18358
rect 7840 18294 7892 18300
rect 6920 18284 6972 18290
rect 6920 18226 6972 18232
rect 6736 18216 6788 18222
rect 6788 18164 6960 18170
rect 6736 18158 6960 18164
rect 6748 18142 6960 18158
rect 6932 18086 6960 18142
rect 6920 18080 6972 18086
rect 6920 18022 6972 18028
rect 7012 18080 7064 18086
rect 7012 18022 7064 18028
rect 6644 17740 6696 17746
rect 6644 17682 6696 17688
rect 6656 17338 6684 17682
rect 6644 17332 6696 17338
rect 6644 17274 6696 17280
rect 6932 17066 6960 18022
rect 7024 17134 7052 18022
rect 7114 17980 7422 17989
rect 7114 17978 7120 17980
rect 7176 17978 7200 17980
rect 7256 17978 7280 17980
rect 7336 17978 7360 17980
rect 7416 17978 7422 17980
rect 7176 17926 7178 17978
rect 7358 17926 7360 17978
rect 7114 17924 7120 17926
rect 7176 17924 7200 17926
rect 7256 17924 7280 17926
rect 7336 17924 7360 17926
rect 7416 17924 7422 17926
rect 7114 17915 7422 17924
rect 7012 17128 7064 17134
rect 7012 17070 7064 17076
rect 6920 17060 6972 17066
rect 6920 17002 6972 17008
rect 7564 17060 7616 17066
rect 7564 17002 7616 17008
rect 6932 16658 6960 17002
rect 7114 16892 7422 16901
rect 7114 16890 7120 16892
rect 7176 16890 7200 16892
rect 7256 16890 7280 16892
rect 7336 16890 7360 16892
rect 7416 16890 7422 16892
rect 7176 16838 7178 16890
rect 7358 16838 7360 16890
rect 7114 16836 7120 16838
rect 7176 16836 7200 16838
rect 7256 16836 7280 16838
rect 7336 16836 7360 16838
rect 7416 16836 7422 16838
rect 7114 16827 7422 16836
rect 7576 16658 7604 17002
rect 7852 16794 7880 18294
rect 8312 17882 8340 18634
rect 8404 18426 8432 19110
rect 8392 18420 8444 18426
rect 8392 18362 8444 18368
rect 8496 18222 8524 19246
rect 8588 18834 8616 19790
rect 8864 19786 8892 21422
rect 9232 21418 9260 28018
rect 9404 28008 9456 28014
rect 9404 27950 9456 27956
rect 9416 27674 9444 27950
rect 9404 27668 9456 27674
rect 9404 27610 9456 27616
rect 9588 27532 9640 27538
rect 9588 27474 9640 27480
rect 9312 27396 9364 27402
rect 9312 27338 9364 27344
rect 9324 23594 9352 27338
rect 9600 26586 9628 27474
rect 9692 26926 9720 28154
rect 9772 27940 9824 27946
rect 9772 27882 9824 27888
rect 9784 27674 9812 27882
rect 9864 27872 9916 27878
rect 9864 27814 9916 27820
rect 9772 27668 9824 27674
rect 9772 27610 9824 27616
rect 9680 26920 9732 26926
rect 9680 26862 9732 26868
rect 9876 26858 9904 27814
rect 10152 27538 10180 28358
rect 10472 28316 10780 28325
rect 10472 28314 10478 28316
rect 10534 28314 10558 28316
rect 10614 28314 10638 28316
rect 10694 28314 10718 28316
rect 10774 28314 10780 28316
rect 10534 28262 10536 28314
rect 10716 28262 10718 28314
rect 10472 28260 10478 28262
rect 10534 28260 10558 28262
rect 10614 28260 10638 28262
rect 10694 28260 10718 28262
rect 10774 28260 10780 28262
rect 10472 28251 10780 28260
rect 10876 28144 10928 28150
rect 10876 28086 10928 28092
rect 10888 27606 10916 28086
rect 10968 27872 11020 27878
rect 10968 27814 11020 27820
rect 10980 27674 11008 27814
rect 10968 27668 11020 27674
rect 10968 27610 11020 27616
rect 10876 27600 10928 27606
rect 10876 27542 10928 27548
rect 9956 27532 10008 27538
rect 9956 27474 10008 27480
rect 10140 27532 10192 27538
rect 10140 27474 10192 27480
rect 10968 27532 11020 27538
rect 10968 27474 11020 27480
rect 11060 27532 11112 27538
rect 11060 27474 11112 27480
rect 9864 26852 9916 26858
rect 9864 26794 9916 26800
rect 9588 26580 9640 26586
rect 9588 26522 9640 26528
rect 9680 26580 9732 26586
rect 9680 26522 9732 26528
rect 9404 25152 9456 25158
rect 9404 25094 9456 25100
rect 9416 24274 9444 25094
rect 9404 24268 9456 24274
rect 9404 24210 9456 24216
rect 9312 23588 9364 23594
rect 9312 23530 9364 23536
rect 9220 21412 9272 21418
rect 9220 21354 9272 21360
rect 9220 21004 9272 21010
rect 9220 20946 9272 20952
rect 9036 20256 9088 20262
rect 9036 20198 9088 20204
rect 9048 20058 9076 20198
rect 9232 20058 9260 20946
rect 8944 20052 8996 20058
rect 8944 19994 8996 20000
rect 9036 20052 9088 20058
rect 9036 19994 9088 20000
rect 9220 20052 9272 20058
rect 9220 19994 9272 20000
rect 8956 19922 8984 19994
rect 8944 19916 8996 19922
rect 8944 19858 8996 19864
rect 8852 19780 8904 19786
rect 8852 19722 8904 19728
rect 8956 19446 8984 19858
rect 9220 19508 9272 19514
rect 9220 19450 9272 19456
rect 8944 19440 8996 19446
rect 8944 19382 8996 19388
rect 8668 19304 8720 19310
rect 8668 19246 8720 19252
rect 8760 19304 8812 19310
rect 8760 19246 8812 19252
rect 8944 19304 8996 19310
rect 8996 19264 9076 19292
rect 8944 19246 8996 19252
rect 8680 18902 8708 19246
rect 8668 18896 8720 18902
rect 8668 18838 8720 18844
rect 8576 18828 8628 18834
rect 8576 18770 8628 18776
rect 8484 18216 8536 18222
rect 8484 18158 8536 18164
rect 8300 17876 8352 17882
rect 8300 17818 8352 17824
rect 8496 17746 8524 18158
rect 8680 18086 8708 18838
rect 8772 18834 8800 19246
rect 8852 19168 8904 19174
rect 8852 19110 8904 19116
rect 8944 19168 8996 19174
rect 8944 19110 8996 19116
rect 8760 18828 8812 18834
rect 8760 18770 8812 18776
rect 8668 18080 8720 18086
rect 8668 18022 8720 18028
rect 8680 17882 8708 18022
rect 8668 17876 8720 17882
rect 8668 17818 8720 17824
rect 8772 17746 8800 18770
rect 8864 18154 8892 19110
rect 8956 18358 8984 19110
rect 9048 18698 9076 19264
rect 9128 19168 9180 19174
rect 9128 19110 9180 19116
rect 9036 18692 9088 18698
rect 9036 18634 9088 18640
rect 9048 18358 9076 18634
rect 8944 18352 8996 18358
rect 8944 18294 8996 18300
rect 9036 18352 9088 18358
rect 9036 18294 9088 18300
rect 9048 18222 9076 18294
rect 8944 18216 8996 18222
rect 8944 18158 8996 18164
rect 9036 18216 9088 18222
rect 9036 18158 9088 18164
rect 8852 18148 8904 18154
rect 8852 18090 8904 18096
rect 8484 17740 8536 17746
rect 8484 17682 8536 17688
rect 8760 17740 8812 17746
rect 8760 17682 8812 17688
rect 7932 17536 7984 17542
rect 7932 17478 7984 17484
rect 7944 17202 7972 17478
rect 8496 17241 8524 17682
rect 8482 17232 8538 17241
rect 7932 17196 7984 17202
rect 7932 17138 7984 17144
rect 8036 17190 8248 17218
rect 8036 17134 8064 17190
rect 8220 17184 8248 17190
rect 8220 17156 8432 17184
rect 8482 17167 8538 17176
rect 8024 17128 8076 17134
rect 8024 17070 8076 17076
rect 8300 17060 8352 17066
rect 8300 17002 8352 17008
rect 8024 16992 8076 16998
rect 8024 16934 8076 16940
rect 8036 16794 8064 16934
rect 7840 16788 7892 16794
rect 7840 16730 7892 16736
rect 8024 16788 8076 16794
rect 8024 16730 8076 16736
rect 6828 16652 6880 16658
rect 6828 16594 6880 16600
rect 6920 16652 6972 16658
rect 6920 16594 6972 16600
rect 7012 16652 7064 16658
rect 7012 16594 7064 16600
rect 7564 16652 7616 16658
rect 7564 16594 7616 16600
rect 8208 16652 8260 16658
rect 8208 16594 8260 16600
rect 6552 16584 6604 16590
rect 6552 16526 6604 16532
rect 6644 16584 6696 16590
rect 6644 16526 6696 16532
rect 4436 16448 4488 16454
rect 4436 16390 4488 16396
rect 6460 16448 6512 16454
rect 6460 16390 6512 16396
rect 4448 16046 4476 16390
rect 6184 16244 6236 16250
rect 6184 16186 6236 16192
rect 4436 16040 4488 16046
rect 4436 15982 4488 15988
rect 6092 16040 6144 16046
rect 6092 15982 6144 15988
rect 4448 15638 4476 15982
rect 4436 15632 4488 15638
rect 4436 15574 4488 15580
rect 3516 15564 3568 15570
rect 3516 15506 3568 15512
rect 4252 15564 4304 15570
rect 4252 15506 4304 15512
rect 3528 15162 3556 15506
rect 4160 15360 4212 15366
rect 4160 15302 4212 15308
rect 3756 15260 4064 15269
rect 3756 15258 3762 15260
rect 3818 15258 3842 15260
rect 3898 15258 3922 15260
rect 3978 15258 4002 15260
rect 4058 15258 4064 15260
rect 3818 15206 3820 15258
rect 4000 15206 4002 15258
rect 3756 15204 3762 15206
rect 3818 15204 3842 15206
rect 3898 15204 3922 15206
rect 3978 15204 4002 15206
rect 4058 15204 4064 15206
rect 3756 15195 4064 15204
rect 3516 15156 3568 15162
rect 3516 15098 3568 15104
rect 3700 14952 3752 14958
rect 3620 14912 3700 14940
rect 3424 14816 3476 14822
rect 3424 14758 3476 14764
rect 3332 14544 3384 14550
rect 3332 14486 3384 14492
rect 3344 13802 3372 14486
rect 3332 13796 3384 13802
rect 3332 13738 3384 13744
rect 3056 13728 3108 13734
rect 3056 13670 3108 13676
rect 2504 13524 2556 13530
rect 2504 13466 2556 13472
rect 2688 13524 2740 13530
rect 2688 13466 2740 13472
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 2412 13388 2464 13394
rect 2412 13330 2464 13336
rect 2424 12986 2452 13330
rect 2412 12980 2464 12986
rect 2412 12922 2464 12928
rect 2320 12708 2372 12714
rect 2320 12650 2372 12656
rect 1952 12436 2004 12442
rect 1952 12378 2004 12384
rect 2516 12306 2544 13466
rect 3344 13462 3372 13738
rect 3436 13462 3464 14758
rect 3516 14408 3568 14414
rect 3516 14350 3568 14356
rect 3528 14074 3556 14350
rect 3516 14068 3568 14074
rect 3516 14010 3568 14016
rect 3332 13456 3384 13462
rect 3332 13398 3384 13404
rect 3424 13456 3476 13462
rect 3424 13398 3476 13404
rect 3528 13394 3556 14010
rect 3516 13388 3568 13394
rect 3516 13330 3568 13336
rect 3148 13184 3200 13190
rect 3148 13126 3200 13132
rect 3160 12764 3188 13126
rect 3160 12736 3372 12764
rect 2688 12708 2740 12714
rect 2688 12650 2740 12656
rect 2780 12708 2832 12714
rect 2780 12650 2832 12656
rect 2700 12322 2728 12650
rect 2792 12442 2820 12650
rect 3148 12640 3200 12646
rect 3148 12582 3200 12588
rect 3240 12640 3292 12646
rect 3240 12582 3292 12588
rect 2780 12436 2832 12442
rect 2780 12378 2832 12384
rect 2504 12300 2556 12306
rect 2700 12294 2820 12322
rect 3160 12306 3188 12582
rect 3252 12442 3280 12582
rect 3240 12436 3292 12442
rect 3240 12378 3292 12384
rect 2504 12242 2556 12248
rect 2516 11694 2544 12242
rect 2792 12238 2820 12294
rect 2964 12300 3016 12306
rect 2964 12242 3016 12248
rect 3148 12300 3200 12306
rect 3148 12242 3200 12248
rect 2780 12232 2832 12238
rect 2780 12174 2832 12180
rect 2976 11830 3004 12242
rect 3344 11898 3372 12736
rect 3528 12374 3556 13330
rect 3516 12368 3568 12374
rect 3516 12310 3568 12316
rect 3332 11892 3384 11898
rect 3384 11852 3464 11880
rect 3332 11834 3384 11840
rect 2688 11824 2740 11830
rect 2688 11766 2740 11772
rect 2964 11824 3016 11830
rect 2964 11766 3016 11772
rect 2700 11694 2728 11766
rect 2504 11688 2556 11694
rect 2504 11630 2556 11636
rect 2688 11688 2740 11694
rect 2688 11630 2740 11636
rect 2136 11552 2188 11558
rect 2136 11494 2188 11500
rect 2148 11354 2176 11494
rect 2136 11348 2188 11354
rect 2136 11290 2188 11296
rect 2516 11082 2544 11630
rect 2504 11076 2556 11082
rect 2504 11018 2556 11024
rect 2136 11008 2188 11014
rect 2136 10950 2188 10956
rect 1860 10260 1912 10266
rect 1860 10202 1912 10208
rect 1860 10124 1912 10130
rect 1860 10066 1912 10072
rect 1872 9042 1900 10066
rect 2148 10062 2176 10950
rect 2320 10464 2372 10470
rect 2320 10406 2372 10412
rect 2136 10056 2188 10062
rect 2136 9998 2188 10004
rect 2044 9920 2096 9926
rect 2044 9862 2096 9868
rect 1952 9444 2004 9450
rect 1952 9386 2004 9392
rect 1676 9036 1728 9042
rect 1676 8978 1728 8984
rect 1860 9036 1912 9042
rect 1860 8978 1912 8984
rect 1688 8498 1716 8978
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 1596 7410 1624 8434
rect 1872 8430 1900 8978
rect 1964 8498 1992 9386
rect 2056 9042 2084 9862
rect 2148 9518 2176 9998
rect 2228 9716 2280 9722
rect 2228 9658 2280 9664
rect 2136 9512 2188 9518
rect 2136 9454 2188 9460
rect 2240 9042 2268 9658
rect 2332 9382 2360 10406
rect 2412 10124 2464 10130
rect 2412 10066 2464 10072
rect 2320 9376 2372 9382
rect 2320 9318 2372 9324
rect 2044 9036 2096 9042
rect 2044 8978 2096 8984
rect 2136 9036 2188 9042
rect 2136 8978 2188 8984
rect 2228 9036 2280 9042
rect 2228 8978 2280 8984
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 1860 8424 1912 8430
rect 1912 8372 1992 8378
rect 1860 8366 1992 8372
rect 1872 8350 1992 8366
rect 1584 7404 1636 7410
rect 1584 7346 1636 7352
rect 1860 7336 1912 7342
rect 1860 7278 1912 7284
rect 1768 7268 1820 7274
rect 1768 7210 1820 7216
rect 1676 7200 1728 7206
rect 1676 7142 1728 7148
rect 1124 6860 1176 6866
rect 1124 6802 1176 6808
rect 1136 6458 1164 6802
rect 1124 6452 1176 6458
rect 1124 6394 1176 6400
rect 1688 6254 1716 7142
rect 1780 6322 1808 7210
rect 1872 7002 1900 7278
rect 1860 6996 1912 7002
rect 1860 6938 1912 6944
rect 1872 6458 1900 6938
rect 1860 6452 1912 6458
rect 1860 6394 1912 6400
rect 1768 6316 1820 6322
rect 1768 6258 1820 6264
rect 1676 6248 1728 6254
rect 1676 6190 1728 6196
rect 1216 5568 1268 5574
rect 1216 5510 1268 5516
rect 1228 5166 1256 5510
rect 1124 5160 1176 5166
rect 1124 5102 1176 5108
rect 1216 5160 1268 5166
rect 1216 5102 1268 5108
rect 1136 4826 1164 5102
rect 1964 4826 1992 8350
rect 2148 8090 2176 8978
rect 2424 8974 2452 10066
rect 2516 9926 2544 11018
rect 2700 10266 2728 11630
rect 2780 11552 2832 11558
rect 2780 11494 2832 11500
rect 2688 10260 2740 10266
rect 2688 10202 2740 10208
rect 2504 9920 2556 9926
rect 2504 9862 2556 9868
rect 2516 9518 2544 9862
rect 2700 9722 2728 10202
rect 2688 9716 2740 9722
rect 2688 9658 2740 9664
rect 2700 9518 2728 9658
rect 2504 9512 2556 9518
rect 2504 9454 2556 9460
rect 2596 9512 2648 9518
rect 2596 9454 2648 9460
rect 2688 9512 2740 9518
rect 2688 9454 2740 9460
rect 2504 9376 2556 9382
rect 2504 9318 2556 9324
rect 2516 9110 2544 9318
rect 2504 9104 2556 9110
rect 2504 9046 2556 9052
rect 2412 8968 2464 8974
rect 2412 8910 2464 8916
rect 2608 8634 2636 9454
rect 2596 8628 2648 8634
rect 2596 8570 2648 8576
rect 2412 8560 2464 8566
rect 2412 8502 2464 8508
rect 2424 8430 2452 8502
rect 2412 8424 2464 8430
rect 2412 8366 2464 8372
rect 2424 8294 2452 8366
rect 2792 8362 2820 11494
rect 2976 11354 3004 11766
rect 3240 11552 3292 11558
rect 3240 11494 3292 11500
rect 2964 11348 3016 11354
rect 2964 11290 3016 11296
rect 2964 11212 3016 11218
rect 2964 11154 3016 11160
rect 2976 9654 3004 11154
rect 3056 10464 3108 10470
rect 3056 10406 3108 10412
rect 3068 9926 3096 10406
rect 3148 10192 3200 10198
rect 3148 10134 3200 10140
rect 3056 9920 3108 9926
rect 3056 9862 3108 9868
rect 2964 9648 3016 9654
rect 2964 9590 3016 9596
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 2884 8566 2912 8910
rect 2976 8906 3004 9318
rect 3160 9178 3188 10134
rect 3252 9518 3280 11494
rect 3332 10668 3384 10674
rect 3332 10610 3384 10616
rect 3240 9512 3292 9518
rect 3240 9454 3292 9460
rect 3148 9172 3200 9178
rect 3148 9114 3200 9120
rect 3056 9036 3108 9042
rect 3056 8978 3108 8984
rect 2964 8900 3016 8906
rect 2964 8842 3016 8848
rect 2872 8560 2924 8566
rect 2872 8502 2924 8508
rect 2872 8424 2924 8430
rect 2976 8412 3004 8842
rect 2924 8384 3004 8412
rect 2872 8366 2924 8372
rect 2780 8356 2832 8362
rect 2780 8298 2832 8304
rect 2412 8288 2464 8294
rect 2412 8230 2464 8236
rect 2136 8084 2188 8090
rect 2136 8026 2188 8032
rect 2424 7546 2452 8230
rect 2412 7540 2464 7546
rect 2412 7482 2464 7488
rect 2136 7336 2188 7342
rect 2136 7278 2188 7284
rect 2148 6662 2176 7278
rect 2504 7268 2556 7274
rect 2504 7210 2556 7216
rect 2516 6866 2544 7210
rect 2884 6934 2912 8366
rect 3068 8362 3096 8978
rect 3252 8922 3280 9454
rect 3344 9178 3372 10610
rect 3436 9518 3464 11852
rect 3516 10532 3568 10538
rect 3516 10474 3568 10480
rect 3528 9722 3556 10474
rect 3620 10198 3648 14912
rect 3700 14894 3752 14900
rect 3756 14172 4064 14181
rect 3756 14170 3762 14172
rect 3818 14170 3842 14172
rect 3898 14170 3922 14172
rect 3978 14170 4002 14172
rect 4058 14170 4064 14172
rect 3818 14118 3820 14170
rect 4000 14118 4002 14170
rect 3756 14116 3762 14118
rect 3818 14116 3842 14118
rect 3898 14116 3922 14118
rect 3978 14116 4002 14118
rect 4058 14116 4064 14118
rect 3756 14107 4064 14116
rect 4068 13864 4120 13870
rect 4172 13818 4200 15302
rect 4120 13812 4200 13818
rect 4068 13806 4200 13812
rect 4080 13790 4200 13806
rect 4080 13190 4108 13790
rect 4160 13388 4212 13394
rect 4160 13330 4212 13336
rect 4068 13184 4120 13190
rect 4068 13126 4120 13132
rect 3756 13084 4064 13093
rect 3756 13082 3762 13084
rect 3818 13082 3842 13084
rect 3898 13082 3922 13084
rect 3978 13082 4002 13084
rect 4058 13082 4064 13084
rect 3818 13030 3820 13082
rect 4000 13030 4002 13082
rect 3756 13028 3762 13030
rect 3818 13028 3842 13030
rect 3898 13028 3922 13030
rect 3978 13028 4002 13030
rect 4058 13028 4064 13030
rect 3756 13019 4064 13028
rect 3976 12640 4028 12646
rect 3976 12582 4028 12588
rect 3988 12374 4016 12582
rect 4172 12442 4200 13330
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 3976 12368 4028 12374
rect 3976 12310 4028 12316
rect 3756 11996 4064 12005
rect 3756 11994 3762 11996
rect 3818 11994 3842 11996
rect 3898 11994 3922 11996
rect 3978 11994 4002 11996
rect 4058 11994 4064 11996
rect 3818 11942 3820 11994
rect 4000 11942 4002 11994
rect 3756 11940 3762 11942
rect 3818 11940 3842 11942
rect 3898 11940 3922 11942
rect 3978 11940 4002 11942
rect 4058 11940 4064 11942
rect 3756 11931 4064 11940
rect 4068 11892 4120 11898
rect 4068 11834 4120 11840
rect 4080 11218 4108 11834
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 4068 11212 4120 11218
rect 4068 11154 4120 11160
rect 4172 11082 4200 11494
rect 4264 11218 4292 15506
rect 4448 15162 4476 15574
rect 6104 15570 6132 15982
rect 6196 15570 6224 16186
rect 6472 15910 6500 16390
rect 6552 15972 6604 15978
rect 6552 15914 6604 15920
rect 6460 15904 6512 15910
rect 6460 15846 6512 15852
rect 6092 15564 6144 15570
rect 6092 15506 6144 15512
rect 6184 15564 6236 15570
rect 6184 15506 6236 15512
rect 5724 15428 5776 15434
rect 5724 15370 5776 15376
rect 4712 15360 4764 15366
rect 4712 15302 4764 15308
rect 5540 15360 5592 15366
rect 5540 15302 5592 15308
rect 4436 15156 4488 15162
rect 4436 15098 4488 15104
rect 4344 14340 4396 14346
rect 4344 14282 4396 14288
rect 4356 13870 4384 14282
rect 4448 14074 4476 15098
rect 4724 15094 4752 15302
rect 4528 15088 4580 15094
rect 4528 15030 4580 15036
rect 4712 15088 4764 15094
rect 4712 15030 4764 15036
rect 4540 14618 4568 15030
rect 5552 14890 5580 15302
rect 5080 14884 5132 14890
rect 5080 14826 5132 14832
rect 5540 14884 5592 14890
rect 5540 14826 5592 14832
rect 4528 14612 4580 14618
rect 4528 14554 4580 14560
rect 4540 14482 4568 14554
rect 4528 14476 4580 14482
rect 4528 14418 4580 14424
rect 4436 14068 4488 14074
rect 4436 14010 4488 14016
rect 4344 13864 4396 13870
rect 4344 13806 4396 13812
rect 4436 12776 4488 12782
rect 4436 12718 4488 12724
rect 4448 12186 4476 12718
rect 4356 12158 4476 12186
rect 4252 11212 4304 11218
rect 4252 11154 4304 11160
rect 4160 11076 4212 11082
rect 4160 11018 4212 11024
rect 3756 10908 4064 10917
rect 3756 10906 3762 10908
rect 3818 10906 3842 10908
rect 3898 10906 3922 10908
rect 3978 10906 4002 10908
rect 4058 10906 4064 10908
rect 3818 10854 3820 10906
rect 4000 10854 4002 10906
rect 3756 10852 3762 10854
rect 3818 10852 3842 10854
rect 3898 10852 3922 10854
rect 3978 10852 4002 10854
rect 4058 10852 4064 10854
rect 3756 10843 4064 10852
rect 3700 10600 3752 10606
rect 3700 10542 3752 10548
rect 3712 10266 3740 10542
rect 4160 10464 4212 10470
rect 4160 10406 4212 10412
rect 3700 10260 3752 10266
rect 3700 10202 3752 10208
rect 3608 10192 3660 10198
rect 3608 10134 3660 10140
rect 3756 9820 4064 9829
rect 3756 9818 3762 9820
rect 3818 9818 3842 9820
rect 3898 9818 3922 9820
rect 3978 9818 4002 9820
rect 4058 9818 4064 9820
rect 3818 9766 3820 9818
rect 4000 9766 4002 9818
rect 3756 9764 3762 9766
rect 3818 9764 3842 9766
rect 3898 9764 3922 9766
rect 3978 9764 4002 9766
rect 4058 9764 4064 9766
rect 3756 9755 4064 9764
rect 3516 9716 3568 9722
rect 3516 9658 3568 9664
rect 3424 9512 3476 9518
rect 3424 9454 3476 9460
rect 3884 9512 3936 9518
rect 3884 9454 3936 9460
rect 3332 9172 3384 9178
rect 3332 9114 3384 9120
rect 3436 9042 3464 9454
rect 3424 9036 3476 9042
rect 3424 8978 3476 8984
rect 3252 8894 3372 8922
rect 3056 8356 3108 8362
rect 3056 8298 3108 8304
rect 3148 8356 3200 8362
rect 3148 8298 3200 8304
rect 3056 8016 3108 8022
rect 3056 7958 3108 7964
rect 2964 7880 3016 7886
rect 2964 7822 3016 7828
rect 2976 7002 3004 7822
rect 3068 7274 3096 7958
rect 3160 7818 3188 8298
rect 3344 8022 3372 8894
rect 3332 8016 3384 8022
rect 3436 8004 3464 8978
rect 3896 8974 3924 9454
rect 4172 9042 4200 10406
rect 4356 9654 4384 12158
rect 4436 12096 4488 12102
rect 4436 12038 4488 12044
rect 4448 11762 4476 12038
rect 4436 11756 4488 11762
rect 4436 11698 4488 11704
rect 4540 11694 4568 14418
rect 4804 14408 4856 14414
rect 4804 14350 4856 14356
rect 4816 13734 4844 14350
rect 5092 14074 5120 14826
rect 5080 14068 5132 14074
rect 5080 14010 5132 14016
rect 4804 13728 4856 13734
rect 4804 13670 4856 13676
rect 4816 13530 4844 13670
rect 4804 13524 4856 13530
rect 4804 13466 4856 13472
rect 4804 13320 4856 13326
rect 4804 13262 4856 13268
rect 4816 12782 4844 13262
rect 5080 12912 5132 12918
rect 5080 12854 5132 12860
rect 4804 12776 4856 12782
rect 4804 12718 4856 12724
rect 4816 12102 4844 12718
rect 4988 12708 5040 12714
rect 4988 12650 5040 12656
rect 5000 12306 5028 12650
rect 5092 12646 5120 12854
rect 5736 12782 5764 15370
rect 6196 14890 6224 15506
rect 6472 15026 6500 15846
rect 6564 15162 6592 15914
rect 6656 15570 6684 16526
rect 6840 15706 6868 16594
rect 6828 15700 6880 15706
rect 6828 15642 6880 15648
rect 6644 15564 6696 15570
rect 6644 15506 6696 15512
rect 6736 15564 6788 15570
rect 6736 15506 6788 15512
rect 6552 15156 6604 15162
rect 6552 15098 6604 15104
rect 6276 15020 6328 15026
rect 6276 14962 6328 14968
rect 6460 15020 6512 15026
rect 6460 14962 6512 14968
rect 6184 14884 6236 14890
rect 6184 14826 6236 14832
rect 6288 14550 6316 14962
rect 6748 14958 6776 15506
rect 6828 15020 6880 15026
rect 6828 14962 6880 14968
rect 6736 14952 6788 14958
rect 6736 14894 6788 14900
rect 6368 14884 6420 14890
rect 6368 14826 6420 14832
rect 6380 14618 6408 14826
rect 6748 14822 6776 14894
rect 6736 14816 6788 14822
rect 6736 14758 6788 14764
rect 6368 14612 6420 14618
rect 6368 14554 6420 14560
rect 6276 14544 6328 14550
rect 6276 14486 6328 14492
rect 5908 14272 5960 14278
rect 5908 14214 5960 14220
rect 5920 13870 5948 14214
rect 6012 13938 6224 13954
rect 6012 13932 6236 13938
rect 6012 13926 6184 13932
rect 5908 13864 5960 13870
rect 5908 13806 5960 13812
rect 6012 13462 6040 13926
rect 6184 13874 6236 13880
rect 6092 13864 6144 13870
rect 6092 13806 6144 13812
rect 6104 13530 6132 13806
rect 6288 13802 6316 14486
rect 6840 14482 6868 14962
rect 6932 14618 6960 16594
rect 7024 15162 7052 16594
rect 7564 16448 7616 16454
rect 7564 16390 7616 16396
rect 7472 15904 7524 15910
rect 7472 15846 7524 15852
rect 7114 15804 7422 15813
rect 7114 15802 7120 15804
rect 7176 15802 7200 15804
rect 7256 15802 7280 15804
rect 7336 15802 7360 15804
rect 7416 15802 7422 15804
rect 7176 15750 7178 15802
rect 7358 15750 7360 15802
rect 7114 15748 7120 15750
rect 7176 15748 7200 15750
rect 7256 15748 7280 15750
rect 7336 15748 7360 15750
rect 7416 15748 7422 15750
rect 7114 15739 7422 15748
rect 7484 15706 7512 15846
rect 7576 15706 7604 16390
rect 8220 16114 8248 16594
rect 8312 16454 8340 17002
rect 8404 16776 8432 17156
rect 8484 16788 8536 16794
rect 8404 16748 8484 16776
rect 8484 16730 8536 16736
rect 8392 16652 8444 16658
rect 8576 16652 8628 16658
rect 8444 16612 8576 16640
rect 8392 16594 8444 16600
rect 8576 16594 8628 16600
rect 8300 16448 8352 16454
rect 8300 16390 8352 16396
rect 8864 16250 8892 18090
rect 8956 17746 8984 18158
rect 9140 17882 9168 19110
rect 9232 18970 9260 19450
rect 9220 18964 9272 18970
rect 9220 18906 9272 18912
rect 9324 18714 9352 23530
rect 9692 23254 9720 26522
rect 9864 26376 9916 26382
rect 9864 26318 9916 26324
rect 9876 26042 9904 26318
rect 9864 26036 9916 26042
rect 9864 25978 9916 25984
rect 9876 25498 9904 25978
rect 9864 25492 9916 25498
rect 9864 25434 9916 25440
rect 9968 25430 9996 27474
rect 10048 27396 10100 27402
rect 10048 27338 10100 27344
rect 10060 27130 10088 27338
rect 10472 27228 10780 27237
rect 10472 27226 10478 27228
rect 10534 27226 10558 27228
rect 10614 27226 10638 27228
rect 10694 27226 10718 27228
rect 10774 27226 10780 27228
rect 10534 27174 10536 27226
rect 10716 27174 10718 27226
rect 10472 27172 10478 27174
rect 10534 27172 10558 27174
rect 10614 27172 10638 27174
rect 10694 27172 10718 27174
rect 10774 27172 10780 27174
rect 10472 27163 10780 27172
rect 10048 27124 10100 27130
rect 10048 27066 10100 27072
rect 10140 26444 10192 26450
rect 10140 26386 10192 26392
rect 10152 25702 10180 26386
rect 10472 26140 10780 26149
rect 10472 26138 10478 26140
rect 10534 26138 10558 26140
rect 10614 26138 10638 26140
rect 10694 26138 10718 26140
rect 10774 26138 10780 26140
rect 10534 26086 10536 26138
rect 10716 26086 10718 26138
rect 10472 26084 10478 26086
rect 10534 26084 10558 26086
rect 10614 26084 10638 26086
rect 10694 26084 10718 26086
rect 10774 26084 10780 26086
rect 10472 26075 10780 26084
rect 10980 25838 11008 27474
rect 11072 27130 11100 27474
rect 11060 27124 11112 27130
rect 11060 27066 11112 27072
rect 11060 26852 11112 26858
rect 11164 26840 11192 29242
rect 11992 29034 12020 29543
rect 12452 29238 12480 29582
rect 12440 29232 12492 29238
rect 12440 29174 12492 29180
rect 11612 29028 11664 29034
rect 11612 28970 11664 28976
rect 11980 29028 12032 29034
rect 11980 28970 12032 28976
rect 12072 29028 12124 29034
rect 12072 28970 12124 28976
rect 11520 27872 11572 27878
rect 11520 27814 11572 27820
rect 11532 26926 11560 27814
rect 11624 26926 11652 28970
rect 11704 28960 11756 28966
rect 11704 28902 11756 28908
rect 11716 28694 11744 28902
rect 11704 28688 11756 28694
rect 11704 28630 11756 28636
rect 11704 28008 11756 28014
rect 11704 27950 11756 27956
rect 11428 26920 11480 26926
rect 11428 26862 11480 26868
rect 11520 26920 11572 26926
rect 11520 26862 11572 26868
rect 11612 26920 11664 26926
rect 11612 26862 11664 26868
rect 11112 26812 11192 26840
rect 11336 26852 11388 26858
rect 11060 26794 11112 26800
rect 11336 26794 11388 26800
rect 10968 25832 11020 25838
rect 10968 25774 11020 25780
rect 10140 25696 10192 25702
rect 10140 25638 10192 25644
rect 9956 25424 10008 25430
rect 9956 25366 10008 25372
rect 9864 24608 9916 24614
rect 9864 24550 9916 24556
rect 9876 23866 9904 24550
rect 9864 23860 9916 23866
rect 9864 23802 9916 23808
rect 9968 23322 9996 25366
rect 10140 25152 10192 25158
rect 10140 25094 10192 25100
rect 10152 24750 10180 25094
rect 10472 25052 10780 25061
rect 10472 25050 10478 25052
rect 10534 25050 10558 25052
rect 10614 25050 10638 25052
rect 10694 25050 10718 25052
rect 10774 25050 10780 25052
rect 10534 24998 10536 25050
rect 10716 24998 10718 25050
rect 10472 24996 10478 24998
rect 10534 24996 10558 24998
rect 10614 24996 10638 24998
rect 10694 24996 10718 24998
rect 10774 24996 10780 24998
rect 10472 24987 10780 24996
rect 10980 24954 11008 25774
rect 11072 25158 11100 26794
rect 11348 26518 11376 26794
rect 11152 26512 11204 26518
rect 11152 26454 11204 26460
rect 11336 26512 11388 26518
rect 11336 26454 11388 26460
rect 11060 25152 11112 25158
rect 11060 25094 11112 25100
rect 10968 24948 11020 24954
rect 10968 24890 11020 24896
rect 10048 24744 10100 24750
rect 10048 24686 10100 24692
rect 10140 24744 10192 24750
rect 10140 24686 10192 24692
rect 10416 24744 10468 24750
rect 10416 24686 10468 24692
rect 10060 24274 10088 24686
rect 10232 24676 10284 24682
rect 10232 24618 10284 24624
rect 10324 24676 10376 24682
rect 10324 24618 10376 24624
rect 10244 24342 10272 24618
rect 10336 24410 10364 24618
rect 10428 24410 10456 24686
rect 10324 24404 10376 24410
rect 10324 24346 10376 24352
rect 10416 24404 10468 24410
rect 10416 24346 10468 24352
rect 10232 24336 10284 24342
rect 10232 24278 10284 24284
rect 10048 24268 10100 24274
rect 10048 24210 10100 24216
rect 9956 23316 10008 23322
rect 9956 23258 10008 23264
rect 9680 23248 9732 23254
rect 9680 23190 9732 23196
rect 10060 23186 10088 24210
rect 10244 23866 10272 24278
rect 10980 24274 11008 24890
rect 11060 24744 11112 24750
rect 11060 24686 11112 24692
rect 10968 24268 11020 24274
rect 10968 24210 11020 24216
rect 10472 23964 10780 23973
rect 10472 23962 10478 23964
rect 10534 23962 10558 23964
rect 10614 23962 10638 23964
rect 10694 23962 10718 23964
rect 10774 23962 10780 23964
rect 10534 23910 10536 23962
rect 10716 23910 10718 23962
rect 10472 23908 10478 23910
rect 10534 23908 10558 23910
rect 10614 23908 10638 23910
rect 10694 23908 10718 23910
rect 10774 23908 10780 23910
rect 10472 23899 10780 23908
rect 10232 23860 10284 23866
rect 10232 23802 10284 23808
rect 10244 23186 10272 23802
rect 11072 23662 11100 24686
rect 11060 23656 11112 23662
rect 11060 23598 11112 23604
rect 10416 23316 10468 23322
rect 10416 23258 10468 23264
rect 10428 23186 10456 23258
rect 11072 23186 11100 23598
rect 11164 23254 11192 26454
rect 11440 26450 11468 26862
rect 11428 26444 11480 26450
rect 11428 26386 11480 26392
rect 11244 26240 11296 26246
rect 11244 26182 11296 26188
rect 11256 25770 11284 26182
rect 11244 25764 11296 25770
rect 11244 25706 11296 25712
rect 11336 24064 11388 24070
rect 11336 24006 11388 24012
rect 11348 23866 11376 24006
rect 11336 23860 11388 23866
rect 11336 23802 11388 23808
rect 11152 23248 11204 23254
rect 11152 23190 11204 23196
rect 11520 23248 11572 23254
rect 11520 23190 11572 23196
rect 9864 23180 9916 23186
rect 9864 23122 9916 23128
rect 9956 23180 10008 23186
rect 9956 23122 10008 23128
rect 10048 23180 10100 23186
rect 10048 23122 10100 23128
rect 10140 23180 10192 23186
rect 10140 23122 10192 23128
rect 10232 23180 10284 23186
rect 10232 23122 10284 23128
rect 10416 23180 10468 23186
rect 10416 23122 10468 23128
rect 11060 23180 11112 23186
rect 11060 23122 11112 23128
rect 9876 22642 9904 23122
rect 9864 22636 9916 22642
rect 9864 22578 9916 22584
rect 9968 22506 9996 23122
rect 10048 22568 10100 22574
rect 10048 22510 10100 22516
rect 9956 22500 10008 22506
rect 9956 22442 10008 22448
rect 9680 22432 9732 22438
rect 9680 22374 9732 22380
rect 9588 21548 9640 21554
rect 9588 21490 9640 21496
rect 9404 20800 9456 20806
rect 9404 20742 9456 20748
rect 9416 20466 9444 20742
rect 9404 20460 9456 20466
rect 9404 20402 9456 20408
rect 9404 20324 9456 20330
rect 9404 20266 9456 20272
rect 9416 19378 9444 20266
rect 9600 19904 9628 21490
rect 9692 21486 9720 22374
rect 10060 21962 10088 22510
rect 10152 22234 10180 23122
rect 10140 22228 10192 22234
rect 10140 22170 10192 22176
rect 10048 21956 10100 21962
rect 10048 21898 10100 21904
rect 10140 21888 10192 21894
rect 10140 21830 10192 21836
rect 10152 21622 10180 21830
rect 10140 21616 10192 21622
rect 10140 21558 10192 21564
rect 10244 21554 10272 23122
rect 10428 23066 10456 23122
rect 10336 23038 10456 23066
rect 10336 22438 10364 23038
rect 10472 22876 10780 22885
rect 10472 22874 10478 22876
rect 10534 22874 10558 22876
rect 10614 22874 10638 22876
rect 10694 22874 10718 22876
rect 10774 22874 10780 22876
rect 10534 22822 10536 22874
rect 10716 22822 10718 22874
rect 10472 22820 10478 22822
rect 10534 22820 10558 22822
rect 10614 22820 10638 22822
rect 10694 22820 10718 22822
rect 10774 22820 10780 22822
rect 10472 22811 10780 22820
rect 10876 22568 10928 22574
rect 10876 22510 10928 22516
rect 10324 22432 10376 22438
rect 10324 22374 10376 22380
rect 10472 21788 10780 21797
rect 10472 21786 10478 21788
rect 10534 21786 10558 21788
rect 10614 21786 10638 21788
rect 10694 21786 10718 21788
rect 10774 21786 10780 21788
rect 10534 21734 10536 21786
rect 10716 21734 10718 21786
rect 10472 21732 10478 21734
rect 10534 21732 10558 21734
rect 10614 21732 10638 21734
rect 10694 21732 10718 21734
rect 10774 21732 10780 21734
rect 10472 21723 10780 21732
rect 10232 21548 10284 21554
rect 10232 21490 10284 21496
rect 10416 21548 10468 21554
rect 10416 21490 10468 21496
rect 9680 21480 9732 21486
rect 9680 21422 9732 21428
rect 9864 21412 9916 21418
rect 9864 21354 9916 21360
rect 9772 20936 9824 20942
rect 9772 20878 9824 20884
rect 9784 20466 9812 20878
rect 9772 20460 9824 20466
rect 9772 20402 9824 20408
rect 9680 19916 9732 19922
rect 9600 19876 9680 19904
rect 9600 19786 9628 19876
rect 9680 19858 9732 19864
rect 9588 19780 9640 19786
rect 9588 19722 9640 19728
rect 9404 19372 9456 19378
rect 9404 19314 9456 19320
rect 9876 19242 9904 21354
rect 10428 21146 10456 21490
rect 10416 21140 10468 21146
rect 10416 21082 10468 21088
rect 9956 21004 10008 21010
rect 9956 20946 10008 20952
rect 9968 20058 9996 20946
rect 10472 20700 10780 20709
rect 10472 20698 10478 20700
rect 10534 20698 10558 20700
rect 10614 20698 10638 20700
rect 10694 20698 10718 20700
rect 10774 20698 10780 20700
rect 10534 20646 10536 20698
rect 10716 20646 10718 20698
rect 10472 20644 10478 20646
rect 10534 20644 10558 20646
rect 10614 20644 10638 20646
rect 10694 20644 10718 20646
rect 10774 20644 10780 20646
rect 10472 20635 10780 20644
rect 10232 20460 10284 20466
rect 10232 20402 10284 20408
rect 10048 20256 10100 20262
rect 10048 20198 10100 20204
rect 9956 20052 10008 20058
rect 9956 19994 10008 20000
rect 10060 19922 10088 20198
rect 10048 19916 10100 19922
rect 10048 19858 10100 19864
rect 9864 19236 9916 19242
rect 9864 19178 9916 19184
rect 9404 19168 9456 19174
rect 9404 19110 9456 19116
rect 9416 18970 9444 19110
rect 9404 18964 9456 18970
rect 9404 18906 9456 18912
rect 9324 18686 9444 18714
rect 9312 18624 9364 18630
rect 9312 18566 9364 18572
rect 9220 18080 9272 18086
rect 9220 18022 9272 18028
rect 9128 17876 9180 17882
rect 9128 17818 9180 17824
rect 9232 17746 9260 18022
rect 9324 17746 9352 18566
rect 8944 17740 8996 17746
rect 8944 17682 8996 17688
rect 9128 17740 9180 17746
rect 9128 17682 9180 17688
rect 9220 17740 9272 17746
rect 9220 17682 9272 17688
rect 9312 17740 9364 17746
rect 9312 17682 9364 17688
rect 9140 17626 9168 17682
rect 9140 17610 9260 17626
rect 9140 17604 9272 17610
rect 9140 17598 9220 17604
rect 9220 17546 9272 17552
rect 9128 17536 9180 17542
rect 9128 17478 9180 17484
rect 9140 17338 9168 17478
rect 9036 17332 9088 17338
rect 9036 17274 9088 17280
rect 9128 17332 9180 17338
rect 9128 17274 9180 17280
rect 9048 17184 9076 17274
rect 8956 17156 9076 17184
rect 8852 16244 8904 16250
rect 8852 16186 8904 16192
rect 8208 16108 8260 16114
rect 8208 16050 8260 16056
rect 7656 15972 7708 15978
rect 7656 15914 7708 15920
rect 7472 15700 7524 15706
rect 7472 15642 7524 15648
rect 7564 15700 7616 15706
rect 7564 15642 7616 15648
rect 7472 15496 7524 15502
rect 7472 15438 7524 15444
rect 7012 15156 7064 15162
rect 7012 15098 7064 15104
rect 7114 14716 7422 14725
rect 7114 14714 7120 14716
rect 7176 14714 7200 14716
rect 7256 14714 7280 14716
rect 7336 14714 7360 14716
rect 7416 14714 7422 14716
rect 7176 14662 7178 14714
rect 7358 14662 7360 14714
rect 7114 14660 7120 14662
rect 7176 14660 7200 14662
rect 7256 14660 7280 14662
rect 7336 14660 7360 14662
rect 7416 14660 7422 14662
rect 7114 14651 7422 14660
rect 7484 14618 7512 15438
rect 6920 14612 6972 14618
rect 6920 14554 6972 14560
rect 7472 14612 7524 14618
rect 7472 14554 7524 14560
rect 6828 14476 6880 14482
rect 6828 14418 6880 14424
rect 6368 14340 6420 14346
rect 6368 14282 6420 14288
rect 6380 13802 6408 14282
rect 6840 14074 6868 14418
rect 7012 14272 7064 14278
rect 7012 14214 7064 14220
rect 7024 14074 7052 14214
rect 7484 14074 7512 14554
rect 6828 14068 6880 14074
rect 6828 14010 6880 14016
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 7472 14068 7524 14074
rect 7472 14010 7524 14016
rect 7668 13938 7696 15914
rect 8484 15700 8536 15706
rect 8484 15642 8536 15648
rect 8024 15632 8076 15638
rect 8024 15574 8076 15580
rect 8036 14618 8064 15574
rect 8392 15496 8444 15502
rect 8392 15438 8444 15444
rect 8404 15162 8432 15438
rect 8392 15156 8444 15162
rect 8392 15098 8444 15104
rect 8300 14816 8352 14822
rect 8220 14776 8300 14804
rect 8024 14612 8076 14618
rect 8024 14554 8076 14560
rect 8116 14612 8168 14618
rect 8116 14554 8168 14560
rect 7656 13932 7708 13938
rect 7656 13874 7708 13880
rect 6276 13796 6328 13802
rect 6276 13738 6328 13744
rect 6368 13796 6420 13802
rect 6368 13738 6420 13744
rect 7114 13628 7422 13637
rect 7114 13626 7120 13628
rect 7176 13626 7200 13628
rect 7256 13626 7280 13628
rect 7336 13626 7360 13628
rect 7416 13626 7422 13628
rect 7176 13574 7178 13626
rect 7358 13574 7360 13626
rect 7114 13572 7120 13574
rect 7176 13572 7200 13574
rect 7256 13572 7280 13574
rect 7336 13572 7360 13574
rect 7416 13572 7422 13574
rect 7114 13563 7422 13572
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 6000 13456 6052 13462
rect 6000 13398 6052 13404
rect 6276 13456 6328 13462
rect 6276 13398 6328 13404
rect 5908 13252 5960 13258
rect 5908 13194 5960 13200
rect 5724 12776 5776 12782
rect 5724 12718 5776 12724
rect 5920 12646 5948 13194
rect 6288 12986 6316 13398
rect 8128 13394 8156 14554
rect 8220 13802 8248 14776
rect 8300 14758 8352 14764
rect 8208 13796 8260 13802
rect 8208 13738 8260 13744
rect 8116 13388 8168 13394
rect 8116 13330 8168 13336
rect 7656 13320 7708 13326
rect 7656 13262 7708 13268
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 6276 12980 6328 12986
rect 6276 12922 6328 12928
rect 6460 12776 6512 12782
rect 6460 12718 6512 12724
rect 5080 12640 5132 12646
rect 5080 12582 5132 12588
rect 5908 12640 5960 12646
rect 5908 12582 5960 12588
rect 5092 12306 5120 12582
rect 4988 12300 5040 12306
rect 4988 12242 5040 12248
rect 5080 12300 5132 12306
rect 5080 12242 5132 12248
rect 4804 12096 4856 12102
rect 4804 12038 4856 12044
rect 4528 11688 4580 11694
rect 4528 11630 4580 11636
rect 4620 11688 4672 11694
rect 4620 11630 4672 11636
rect 4632 11354 4660 11630
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 4816 11286 4844 12038
rect 4988 11824 5040 11830
rect 5092 11812 5120 12242
rect 6472 12102 6500 12718
rect 6552 12232 6604 12238
rect 6552 12174 6604 12180
rect 5448 12096 5500 12102
rect 5448 12038 5500 12044
rect 6460 12096 6512 12102
rect 6460 12038 6512 12044
rect 5040 11784 5120 11812
rect 4988 11766 5040 11772
rect 4896 11756 4948 11762
rect 4896 11698 4948 11704
rect 4804 11280 4856 11286
rect 4804 11222 4856 11228
rect 4804 10464 4856 10470
rect 4804 10406 4856 10412
rect 4344 9648 4396 9654
rect 4344 9590 4396 9596
rect 4816 9518 4844 10406
rect 4908 10266 4936 11698
rect 5000 11218 5028 11766
rect 5460 11218 5488 12038
rect 6564 11642 6592 12174
rect 6828 12096 6880 12102
rect 6828 12038 6880 12044
rect 6564 11614 6684 11642
rect 6552 11552 6604 11558
rect 6552 11494 6604 11500
rect 6564 11218 6592 11494
rect 6656 11370 6684 11614
rect 6656 11342 6776 11370
rect 6748 11218 6776 11342
rect 6840 11218 6868 12038
rect 6932 11354 6960 13126
rect 7392 12986 7420 13126
rect 7380 12980 7432 12986
rect 7380 12922 7432 12928
rect 7012 12708 7064 12714
rect 7012 12650 7064 12656
rect 7472 12708 7524 12714
rect 7472 12650 7524 12656
rect 7024 12306 7052 12650
rect 7114 12540 7422 12549
rect 7114 12538 7120 12540
rect 7176 12538 7200 12540
rect 7256 12538 7280 12540
rect 7336 12538 7360 12540
rect 7416 12538 7422 12540
rect 7176 12486 7178 12538
rect 7358 12486 7360 12538
rect 7114 12484 7120 12486
rect 7176 12484 7200 12486
rect 7256 12484 7280 12486
rect 7336 12484 7360 12486
rect 7416 12484 7422 12486
rect 7114 12475 7422 12484
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 7484 11898 7512 12650
rect 7668 12306 7696 13262
rect 7748 13252 7800 13258
rect 7748 13194 7800 13200
rect 7760 12850 7788 13194
rect 8128 12986 8156 13330
rect 8116 12980 8168 12986
rect 8116 12922 8168 12928
rect 7748 12844 7800 12850
rect 7748 12786 7800 12792
rect 7760 12442 7788 12786
rect 7748 12436 7800 12442
rect 7748 12378 7800 12384
rect 8220 12306 8248 13738
rect 8404 13326 8432 15098
rect 8496 14278 8524 15642
rect 8668 15360 8720 15366
rect 8668 15302 8720 15308
rect 8680 14958 8708 15302
rect 8864 14958 8892 16186
rect 8668 14952 8720 14958
rect 8668 14894 8720 14900
rect 8852 14952 8904 14958
rect 8852 14894 8904 14900
rect 8668 14476 8720 14482
rect 8668 14418 8720 14424
rect 8484 14272 8536 14278
rect 8484 14214 8536 14220
rect 8680 14074 8708 14418
rect 8668 14068 8720 14074
rect 8668 14010 8720 14016
rect 8864 13870 8892 14894
rect 8852 13864 8904 13870
rect 8852 13806 8904 13812
rect 8392 13320 8444 13326
rect 8392 13262 8444 13268
rect 8576 13184 8628 13190
rect 8576 13126 8628 13132
rect 8588 12986 8616 13126
rect 8576 12980 8628 12986
rect 8576 12922 8628 12928
rect 8300 12640 8352 12646
rect 8300 12582 8352 12588
rect 8312 12306 8340 12582
rect 8956 12434 8984 17156
rect 9036 17060 9088 17066
rect 9036 17002 9088 17008
rect 9048 16794 9076 17002
rect 9036 16788 9088 16794
rect 9036 16730 9088 16736
rect 9036 16584 9088 16590
rect 9036 16526 9088 16532
rect 9048 16114 9076 16526
rect 9416 16250 9444 18686
rect 9588 18352 9640 18358
rect 9588 18294 9640 18300
rect 9496 18080 9548 18086
rect 9496 18022 9548 18028
rect 9508 17882 9536 18022
rect 9496 17876 9548 17882
rect 9496 17818 9548 17824
rect 9600 17728 9628 18294
rect 9680 18284 9732 18290
rect 9680 18226 9732 18232
rect 9692 17882 9720 18226
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9772 17740 9824 17746
rect 9600 17700 9772 17728
rect 9772 17682 9824 17688
rect 9680 17332 9732 17338
rect 9680 17274 9732 17280
rect 9404 16244 9456 16250
rect 9404 16186 9456 16192
rect 9036 16108 9088 16114
rect 9036 16050 9088 16056
rect 9048 15706 9076 16050
rect 9036 15700 9088 15706
rect 9036 15642 9088 15648
rect 9692 14958 9720 17274
rect 9680 14952 9732 14958
rect 9680 14894 9732 14900
rect 9128 14884 9180 14890
rect 9128 14826 9180 14832
rect 9404 14884 9456 14890
rect 9404 14826 9456 14832
rect 9036 14544 9088 14550
rect 9036 14486 9088 14492
rect 9048 14260 9076 14486
rect 9140 14414 9168 14826
rect 9416 14618 9444 14826
rect 9404 14612 9456 14618
rect 9404 14554 9456 14560
rect 9496 14612 9548 14618
rect 9496 14554 9548 14560
rect 9128 14408 9180 14414
rect 9128 14350 9180 14356
rect 9508 14260 9536 14554
rect 9588 14476 9640 14482
rect 9588 14418 9640 14424
rect 9600 14346 9628 14418
rect 9588 14340 9640 14346
rect 9588 14282 9640 14288
rect 9048 14232 9536 14260
rect 9220 12640 9272 12646
rect 9220 12582 9272 12588
rect 8680 12406 8984 12434
rect 9232 12434 9260 12582
rect 9232 12406 9352 12434
rect 8680 12306 8708 12406
rect 8944 12368 8996 12374
rect 8944 12310 8996 12316
rect 7656 12300 7708 12306
rect 7656 12242 7708 12248
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 8300 12300 8352 12306
rect 8300 12242 8352 12248
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 8668 12300 8720 12306
rect 8668 12242 8720 12248
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7472 11892 7524 11898
rect 7472 11834 7524 11840
rect 7114 11452 7422 11461
rect 7114 11450 7120 11452
rect 7176 11450 7200 11452
rect 7256 11450 7280 11452
rect 7336 11450 7360 11452
rect 7416 11450 7422 11452
rect 7176 11398 7178 11450
rect 7358 11398 7360 11450
rect 7114 11396 7120 11398
rect 7176 11396 7200 11398
rect 7256 11396 7280 11398
rect 7336 11396 7360 11398
rect 7416 11396 7422 11398
rect 7114 11387 7422 11396
rect 6920 11348 6972 11354
rect 6920 11290 6972 11296
rect 7484 11286 7512 11834
rect 7576 11694 7604 12174
rect 8496 11898 8524 12242
rect 8484 11892 8536 11898
rect 8484 11834 8536 11840
rect 7564 11688 7616 11694
rect 7564 11630 7616 11636
rect 7472 11280 7524 11286
rect 7472 11222 7524 11228
rect 4988 11212 5040 11218
rect 4988 11154 5040 11160
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 6552 11212 6604 11218
rect 6552 11154 6604 11160
rect 6644 11212 6696 11218
rect 6644 11154 6696 11160
rect 6736 11212 6788 11218
rect 6736 11154 6788 11160
rect 6828 11212 6880 11218
rect 6828 11154 6880 11160
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 5000 10810 5028 11154
rect 5460 11098 5488 11154
rect 5460 11070 5580 11098
rect 4988 10804 5040 10810
rect 4988 10746 5040 10752
rect 5000 10606 5028 10746
rect 5552 10742 5580 11070
rect 6092 11008 6144 11014
rect 6092 10950 6144 10956
rect 5540 10736 5592 10742
rect 5540 10678 5592 10684
rect 5816 10736 5868 10742
rect 5816 10678 5868 10684
rect 5552 10606 5580 10678
rect 4988 10600 5040 10606
rect 4988 10542 5040 10548
rect 5172 10600 5224 10606
rect 5172 10542 5224 10548
rect 5540 10600 5592 10606
rect 5540 10542 5592 10548
rect 5184 10470 5212 10542
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 4896 10260 4948 10266
rect 4896 10202 4948 10208
rect 4908 9722 4936 10202
rect 5828 10198 5856 10678
rect 5816 10192 5868 10198
rect 5816 10134 5868 10140
rect 5828 9722 5856 10134
rect 6104 10130 6132 10950
rect 6276 10736 6328 10742
rect 6276 10678 6328 10684
rect 6288 10470 6316 10678
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 6276 10464 6328 10470
rect 6276 10406 6328 10412
rect 6368 10464 6420 10470
rect 6368 10406 6420 10412
rect 6460 10464 6512 10470
rect 6460 10406 6512 10412
rect 6092 10124 6144 10130
rect 6092 10066 6144 10072
rect 6000 10056 6052 10062
rect 6000 9998 6052 10004
rect 4896 9716 4948 9722
rect 4896 9658 4948 9664
rect 5816 9716 5868 9722
rect 5816 9658 5868 9664
rect 4804 9512 4856 9518
rect 4804 9454 4856 9460
rect 6012 9450 6040 9998
rect 6380 9450 6408 10406
rect 6472 10130 6500 10406
rect 6460 10124 6512 10130
rect 6460 10066 6512 10072
rect 6460 9920 6512 9926
rect 6564 9908 6592 10542
rect 6656 10266 6684 11154
rect 6736 10804 6788 10810
rect 6736 10746 6788 10752
rect 6828 10804 6880 10810
rect 6828 10746 6880 10752
rect 6748 10606 6776 10746
rect 6840 10606 6868 10746
rect 6736 10600 6788 10606
rect 6736 10542 6788 10548
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 6644 10260 6696 10266
rect 6644 10202 6696 10208
rect 6932 10130 6960 11154
rect 7484 10606 7512 11222
rect 7472 10600 7524 10606
rect 7472 10542 7524 10548
rect 7114 10364 7422 10373
rect 7114 10362 7120 10364
rect 7176 10362 7200 10364
rect 7256 10362 7280 10364
rect 7336 10362 7360 10364
rect 7416 10362 7422 10364
rect 7176 10310 7178 10362
rect 7358 10310 7360 10362
rect 7114 10308 7120 10310
rect 7176 10308 7200 10310
rect 7256 10308 7280 10310
rect 7336 10308 7360 10310
rect 7416 10308 7422 10310
rect 7114 10299 7422 10308
rect 7576 10266 7604 11630
rect 7748 11620 7800 11626
rect 7748 11562 7800 11568
rect 7760 11354 7788 11562
rect 8392 11552 8444 11558
rect 8392 11494 8444 11500
rect 8404 11354 8432 11494
rect 7748 11348 7800 11354
rect 7748 11290 7800 11296
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 8496 11014 8524 11834
rect 8680 11218 8708 12242
rect 8760 11688 8812 11694
rect 8760 11630 8812 11636
rect 8852 11688 8904 11694
rect 8852 11630 8904 11636
rect 8772 11354 8800 11630
rect 8864 11354 8892 11630
rect 8760 11348 8812 11354
rect 8760 11290 8812 11296
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 8956 11218 8984 12310
rect 9324 12306 9352 12406
rect 9692 12374 9720 14894
rect 9772 14476 9824 14482
rect 9876 14464 9904 19178
rect 9956 19168 10008 19174
rect 9956 19110 10008 19116
rect 9968 18426 9996 19110
rect 10244 18834 10272 20402
rect 10472 19612 10780 19621
rect 10472 19610 10478 19612
rect 10534 19610 10558 19612
rect 10614 19610 10638 19612
rect 10694 19610 10718 19612
rect 10774 19610 10780 19612
rect 10534 19558 10536 19610
rect 10716 19558 10718 19610
rect 10472 19556 10478 19558
rect 10534 19556 10558 19558
rect 10614 19556 10638 19558
rect 10694 19556 10718 19558
rect 10774 19556 10780 19558
rect 10472 19547 10780 19556
rect 10416 19304 10468 19310
rect 10416 19246 10468 19252
rect 10508 19304 10560 19310
rect 10508 19246 10560 19252
rect 10324 19168 10376 19174
rect 10324 19110 10376 19116
rect 10232 18828 10284 18834
rect 10152 18788 10232 18816
rect 9956 18420 10008 18426
rect 9956 18362 10008 18368
rect 10152 18306 10180 18788
rect 10232 18770 10284 18776
rect 10232 18692 10284 18698
rect 10232 18634 10284 18640
rect 9968 18278 10180 18306
rect 9968 17134 9996 18278
rect 10048 18216 10100 18222
rect 10048 18158 10100 18164
rect 10060 17134 10088 18158
rect 10140 17672 10192 17678
rect 10140 17614 10192 17620
rect 9956 17128 10008 17134
rect 9956 17070 10008 17076
rect 10048 17128 10100 17134
rect 10048 17070 10100 17076
rect 10060 16658 10088 17070
rect 10152 16998 10180 17614
rect 10244 17542 10272 18634
rect 10336 17746 10364 19110
rect 10428 18698 10456 19246
rect 10416 18692 10468 18698
rect 10416 18634 10468 18640
rect 10520 18630 10548 19246
rect 10508 18624 10560 18630
rect 10508 18566 10560 18572
rect 10472 18524 10780 18533
rect 10472 18522 10478 18524
rect 10534 18522 10558 18524
rect 10614 18522 10638 18524
rect 10694 18522 10718 18524
rect 10774 18522 10780 18524
rect 10534 18470 10536 18522
rect 10716 18470 10718 18522
rect 10472 18468 10478 18470
rect 10534 18468 10558 18470
rect 10614 18468 10638 18470
rect 10694 18468 10718 18470
rect 10774 18468 10780 18470
rect 10472 18459 10780 18468
rect 10888 17746 10916 22510
rect 11072 22438 11100 23122
rect 11152 22976 11204 22982
rect 11152 22918 11204 22924
rect 11244 22976 11296 22982
rect 11244 22918 11296 22924
rect 11060 22432 11112 22438
rect 11060 22374 11112 22380
rect 11072 22098 11100 22374
rect 11060 22092 11112 22098
rect 11060 22034 11112 22040
rect 10966 21992 11022 22001
rect 10966 21927 11022 21936
rect 10980 21418 11008 21927
rect 11164 21486 11192 22918
rect 11256 22166 11284 22918
rect 11244 22160 11296 22166
rect 11244 22102 11296 22108
rect 11428 22092 11480 22098
rect 11428 22034 11480 22040
rect 11440 21486 11468 22034
rect 11152 21480 11204 21486
rect 11152 21422 11204 21428
rect 11428 21480 11480 21486
rect 11428 21422 11480 21428
rect 10968 21412 11020 21418
rect 10968 21354 11020 21360
rect 10968 21004 11020 21010
rect 10968 20946 11020 20952
rect 10980 20058 11008 20946
rect 11532 20618 11560 23190
rect 11624 22574 11652 26862
rect 11716 26450 11744 27950
rect 12084 26586 12112 28970
rect 12624 28960 12676 28966
rect 12624 28902 12676 28908
rect 12636 28014 12664 28902
rect 12716 28620 12768 28626
rect 12716 28562 12768 28568
rect 12728 28218 12756 28562
rect 12820 28558 12848 30194
rect 13004 29850 13032 30262
rect 13084 30184 13136 30190
rect 13084 30126 13136 30132
rect 12992 29844 13044 29850
rect 12992 29786 13044 29792
rect 13096 29714 13124 30126
rect 13084 29708 13136 29714
rect 13084 29650 13136 29656
rect 12992 29504 13044 29510
rect 12992 29446 13044 29452
rect 13084 29504 13136 29510
rect 13136 29464 13216 29492
rect 13084 29446 13136 29452
rect 12808 28552 12860 28558
rect 12808 28494 12860 28500
rect 12716 28212 12768 28218
rect 12716 28154 12768 28160
rect 12532 28008 12584 28014
rect 12532 27950 12584 27956
rect 12624 28008 12676 28014
rect 12624 27950 12676 27956
rect 12544 27402 12572 27950
rect 12532 27396 12584 27402
rect 12532 27338 12584 27344
rect 12072 26580 12124 26586
rect 12072 26522 12124 26528
rect 12256 26512 12308 26518
rect 12256 26454 12308 26460
rect 11704 26444 11756 26450
rect 11704 26386 11756 26392
rect 12072 26444 12124 26450
rect 12072 26386 12124 26392
rect 11888 25764 11940 25770
rect 11888 25706 11940 25712
rect 11900 25498 11928 25706
rect 11888 25492 11940 25498
rect 11888 25434 11940 25440
rect 12084 25158 12112 26386
rect 12268 25362 12296 26454
rect 12636 26450 12664 27950
rect 12820 27538 12848 28494
rect 12808 27532 12860 27538
rect 12808 27474 12860 27480
rect 12900 27532 12952 27538
rect 12900 27474 12952 27480
rect 12820 27130 12848 27474
rect 12808 27124 12860 27130
rect 12808 27066 12860 27072
rect 12808 26920 12860 26926
rect 12808 26862 12860 26868
rect 12624 26444 12676 26450
rect 12624 26386 12676 26392
rect 12820 26432 12848 26862
rect 12912 26586 12940 27474
rect 12900 26580 12952 26586
rect 12900 26522 12952 26528
rect 12900 26444 12952 26450
rect 12820 26404 12900 26432
rect 12532 26376 12584 26382
rect 12532 26318 12584 26324
rect 12544 26042 12572 26318
rect 12532 26036 12584 26042
rect 12532 25978 12584 25984
rect 12256 25356 12308 25362
rect 12256 25298 12308 25304
rect 12072 25152 12124 25158
rect 12072 25094 12124 25100
rect 11796 24608 11848 24614
rect 11796 24550 11848 24556
rect 11808 24410 11836 24550
rect 11796 24404 11848 24410
rect 11796 24346 11848 24352
rect 11888 23588 11940 23594
rect 11888 23530 11940 23536
rect 11900 22982 11928 23530
rect 12084 23186 12112 25094
rect 12164 24268 12216 24274
rect 12164 24210 12216 24216
rect 12176 23866 12204 24210
rect 12164 23860 12216 23866
rect 12164 23802 12216 23808
rect 12268 23186 12296 25298
rect 12820 24138 12848 26404
rect 12900 26386 12952 26392
rect 12900 24676 12952 24682
rect 12900 24618 12952 24624
rect 12808 24132 12860 24138
rect 12808 24074 12860 24080
rect 12912 23866 12940 24618
rect 12900 23860 12952 23866
rect 12900 23802 12952 23808
rect 11980 23180 12032 23186
rect 11980 23122 12032 23128
rect 12072 23180 12124 23186
rect 12072 23122 12124 23128
rect 12256 23180 12308 23186
rect 12256 23122 12308 23128
rect 11888 22976 11940 22982
rect 11888 22918 11940 22924
rect 11992 22778 12020 23122
rect 12084 23050 12112 23122
rect 12072 23044 12124 23050
rect 12072 22986 12124 22992
rect 11980 22772 12032 22778
rect 11980 22714 12032 22720
rect 11612 22568 11664 22574
rect 11612 22510 11664 22516
rect 11348 20590 11560 20618
rect 11348 20330 11376 20590
rect 11060 20324 11112 20330
rect 11060 20266 11112 20272
rect 11336 20324 11388 20330
rect 11336 20266 11388 20272
rect 11072 20058 11100 20266
rect 11152 20256 11204 20262
rect 11152 20198 11204 20204
rect 10968 20052 11020 20058
rect 10968 19994 11020 20000
rect 11060 20052 11112 20058
rect 11060 19994 11112 20000
rect 11164 19718 11192 20198
rect 11348 19990 11376 20266
rect 11336 19984 11388 19990
rect 11336 19926 11388 19932
rect 11244 19916 11296 19922
rect 11244 19858 11296 19864
rect 11428 19916 11480 19922
rect 11428 19858 11480 19864
rect 10968 19712 11020 19718
rect 10968 19654 11020 19660
rect 11152 19712 11204 19718
rect 11152 19654 11204 19660
rect 10324 17740 10376 17746
rect 10324 17682 10376 17688
rect 10876 17740 10928 17746
rect 10876 17682 10928 17688
rect 10876 17604 10928 17610
rect 10876 17546 10928 17552
rect 10232 17536 10284 17542
rect 10232 17478 10284 17484
rect 10324 17536 10376 17542
rect 10324 17478 10376 17484
rect 10336 17320 10364 17478
rect 10472 17436 10780 17445
rect 10472 17434 10478 17436
rect 10534 17434 10558 17436
rect 10614 17434 10638 17436
rect 10694 17434 10718 17436
rect 10774 17434 10780 17436
rect 10534 17382 10536 17434
rect 10716 17382 10718 17434
rect 10472 17380 10478 17382
rect 10534 17380 10558 17382
rect 10614 17380 10638 17382
rect 10694 17380 10718 17382
rect 10774 17380 10780 17382
rect 10472 17371 10780 17380
rect 10600 17332 10652 17338
rect 10336 17292 10456 17320
rect 10232 17196 10284 17202
rect 10232 17138 10284 17144
rect 10324 17196 10376 17202
rect 10324 17138 10376 17144
rect 10140 16992 10192 16998
rect 10140 16934 10192 16940
rect 10048 16652 10100 16658
rect 10152 16640 10180 16934
rect 10244 16794 10272 17138
rect 10336 16794 10364 17138
rect 10428 17134 10456 17292
rect 10600 17274 10652 17280
rect 10506 17232 10562 17241
rect 10506 17167 10562 17176
rect 10520 17134 10548 17167
rect 10416 17128 10468 17134
rect 10416 17070 10468 17076
rect 10508 17128 10560 17134
rect 10508 17070 10560 17076
rect 10232 16788 10284 16794
rect 10232 16730 10284 16736
rect 10324 16788 10376 16794
rect 10324 16730 10376 16736
rect 10324 16652 10376 16658
rect 10152 16612 10324 16640
rect 10048 16594 10100 16600
rect 10324 16594 10376 16600
rect 10612 16522 10640 17274
rect 10888 16794 10916 17546
rect 10980 17338 11008 19654
rect 11060 19508 11112 19514
rect 11060 19450 11112 19456
rect 11072 19394 11100 19450
rect 11072 19366 11192 19394
rect 11256 19378 11284 19858
rect 11440 19514 11468 19858
rect 11428 19508 11480 19514
rect 11428 19450 11480 19456
rect 11060 19304 11112 19310
rect 11060 19246 11112 19252
rect 11072 18970 11100 19246
rect 11164 19174 11192 19366
rect 11244 19372 11296 19378
rect 11244 19314 11296 19320
rect 11152 19168 11204 19174
rect 11152 19110 11204 19116
rect 11060 18964 11112 18970
rect 11060 18906 11112 18912
rect 11060 18284 11112 18290
rect 11060 18226 11112 18232
rect 11072 17882 11100 18226
rect 11624 18222 11652 22510
rect 11796 21480 11848 21486
rect 11796 21422 11848 21428
rect 11808 21010 11836 21422
rect 11796 21004 11848 21010
rect 11796 20946 11848 20952
rect 11808 20466 11836 20946
rect 11796 20460 11848 20466
rect 11796 20402 11848 20408
rect 11992 19174 12020 22714
rect 12084 22710 12112 22986
rect 12072 22704 12124 22710
rect 12072 22646 12124 22652
rect 12268 21690 12296 23122
rect 12808 23112 12860 23118
rect 12808 23054 12860 23060
rect 12440 22636 12492 22642
rect 12440 22578 12492 22584
rect 12452 22506 12480 22578
rect 12440 22500 12492 22506
rect 12440 22442 12492 22448
rect 12256 21684 12308 21690
rect 12256 21626 12308 21632
rect 12452 21486 12480 22442
rect 12820 22234 12848 23054
rect 12900 22568 12952 22574
rect 12900 22510 12952 22516
rect 12808 22228 12860 22234
rect 12808 22170 12860 22176
rect 12912 21554 12940 22510
rect 12900 21548 12952 21554
rect 12900 21490 12952 21496
rect 12440 21480 12492 21486
rect 12440 21422 12492 21428
rect 12452 21146 12480 21422
rect 12808 21412 12860 21418
rect 12808 21354 12860 21360
rect 12440 21140 12492 21146
rect 12440 21082 12492 21088
rect 12624 20936 12676 20942
rect 12624 20878 12676 20884
rect 12348 20800 12400 20806
rect 12348 20742 12400 20748
rect 12360 20398 12388 20742
rect 12348 20392 12400 20398
rect 12348 20334 12400 20340
rect 12532 20256 12584 20262
rect 12532 20198 12584 20204
rect 12544 19922 12572 20198
rect 12636 20058 12664 20878
rect 12624 20052 12676 20058
rect 12624 19994 12676 20000
rect 12532 19916 12584 19922
rect 12532 19858 12584 19864
rect 12072 19508 12124 19514
rect 12072 19450 12124 19456
rect 12084 19242 12112 19450
rect 12256 19440 12308 19446
rect 12256 19382 12308 19388
rect 12268 19310 12296 19382
rect 12256 19304 12308 19310
rect 12308 19264 12388 19292
rect 12256 19246 12308 19252
rect 12072 19236 12124 19242
rect 12072 19178 12124 19184
rect 11980 19168 12032 19174
rect 12256 19168 12308 19174
rect 11980 19110 12032 19116
rect 12176 19116 12256 19122
rect 12176 19110 12308 19116
rect 11612 18216 11664 18222
rect 11612 18158 11664 18164
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 11152 17536 11204 17542
rect 11152 17478 11204 17484
rect 10968 17332 11020 17338
rect 10968 17274 11020 17280
rect 11164 17134 11192 17478
rect 10968 17128 11020 17134
rect 10968 17070 11020 17076
rect 11152 17128 11204 17134
rect 11152 17070 11204 17076
rect 10980 16794 11008 17070
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 10876 16788 10928 16794
rect 10876 16730 10928 16736
rect 10968 16788 11020 16794
rect 10968 16730 11020 16736
rect 11060 16652 11112 16658
rect 11060 16594 11112 16600
rect 10600 16516 10652 16522
rect 10600 16458 10652 16464
rect 10876 16448 10928 16454
rect 10876 16390 10928 16396
rect 10472 16348 10780 16357
rect 10472 16346 10478 16348
rect 10534 16346 10558 16348
rect 10614 16346 10638 16348
rect 10694 16346 10718 16348
rect 10774 16346 10780 16348
rect 10534 16294 10536 16346
rect 10716 16294 10718 16346
rect 10472 16292 10478 16294
rect 10534 16292 10558 16294
rect 10614 16292 10638 16294
rect 10694 16292 10718 16294
rect 10774 16292 10780 16294
rect 10472 16283 10780 16292
rect 10690 16008 10746 16017
rect 9956 15972 10008 15978
rect 10690 15943 10692 15952
rect 9956 15914 10008 15920
rect 10744 15943 10746 15952
rect 10692 15914 10744 15920
rect 9824 14436 9904 14464
rect 9772 14418 9824 14424
rect 9862 14376 9918 14385
rect 9862 14311 9918 14320
rect 9876 14278 9904 14311
rect 9864 14272 9916 14278
rect 9864 14214 9916 14220
rect 9772 13524 9824 13530
rect 9772 13466 9824 13472
rect 9784 12850 9812 13466
rect 9772 12844 9824 12850
rect 9772 12786 9824 12792
rect 9680 12368 9732 12374
rect 9680 12310 9732 12316
rect 9128 12300 9180 12306
rect 9128 12242 9180 12248
rect 9312 12300 9364 12306
rect 9312 12242 9364 12248
rect 9140 11694 9168 12242
rect 9312 12096 9364 12102
rect 9312 12038 9364 12044
rect 9588 12096 9640 12102
rect 9588 12038 9640 12044
rect 9324 11694 9352 12038
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 9312 11688 9364 11694
rect 9312 11630 9364 11636
rect 8668 11212 8720 11218
rect 8668 11154 8720 11160
rect 8944 11212 8996 11218
rect 8944 11154 8996 11160
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 8208 10600 8260 10606
rect 8208 10542 8260 10548
rect 8024 10464 8076 10470
rect 8024 10406 8076 10412
rect 8036 10266 8064 10406
rect 7564 10260 7616 10266
rect 7564 10202 7616 10208
rect 8024 10260 8076 10266
rect 8024 10202 8076 10208
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6512 9880 6592 9908
rect 6460 9862 6512 9868
rect 6000 9444 6052 9450
rect 6000 9386 6052 9392
rect 6368 9444 6420 9450
rect 6368 9386 6420 9392
rect 6012 9178 6040 9386
rect 6472 9382 6500 9862
rect 6932 9722 6960 10066
rect 8220 9722 8248 10542
rect 8956 10266 8984 11154
rect 9140 10606 9168 11630
rect 9128 10600 9180 10606
rect 9128 10542 9180 10548
rect 8944 10260 8996 10266
rect 8996 10220 9076 10248
rect 8944 10202 8996 10208
rect 8668 9920 8720 9926
rect 8668 9862 8720 9868
rect 6920 9716 6972 9722
rect 6920 9658 6972 9664
rect 7472 9716 7524 9722
rect 7472 9658 7524 9664
rect 8208 9716 8260 9722
rect 8208 9658 8260 9664
rect 6460 9376 6512 9382
rect 6460 9318 6512 9324
rect 7114 9276 7422 9285
rect 7114 9274 7120 9276
rect 7176 9274 7200 9276
rect 7256 9274 7280 9276
rect 7336 9274 7360 9276
rect 7416 9274 7422 9276
rect 7176 9222 7178 9274
rect 7358 9222 7360 9274
rect 7114 9220 7120 9222
rect 7176 9220 7200 9222
rect 7256 9220 7280 9222
rect 7336 9220 7360 9222
rect 7416 9220 7422 9222
rect 7114 9211 7422 9220
rect 6000 9172 6052 9178
rect 6000 9114 6052 9120
rect 7484 9042 7512 9658
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 7944 9042 7972 9454
rect 8680 9450 8708 9862
rect 9048 9586 9076 10220
rect 8852 9580 8904 9586
rect 8852 9522 8904 9528
rect 9036 9580 9088 9586
rect 9036 9522 9088 9528
rect 8668 9444 8720 9450
rect 8668 9386 8720 9392
rect 8864 9178 8892 9522
rect 9048 9178 9076 9522
rect 8852 9172 8904 9178
rect 8852 9114 8904 9120
rect 9036 9172 9088 9178
rect 9036 9114 9088 9120
rect 4160 9036 4212 9042
rect 4160 8978 4212 8984
rect 7472 9036 7524 9042
rect 7472 8978 7524 8984
rect 7932 9036 7984 9042
rect 7932 8978 7984 8984
rect 3884 8968 3936 8974
rect 3884 8910 3936 8916
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 3756 8732 4064 8741
rect 3756 8730 3762 8732
rect 3818 8730 3842 8732
rect 3898 8730 3922 8732
rect 3978 8730 4002 8732
rect 4058 8730 4064 8732
rect 3818 8678 3820 8730
rect 4000 8678 4002 8730
rect 3756 8676 3762 8678
rect 3818 8676 3842 8678
rect 3898 8676 3922 8678
rect 3978 8676 4002 8678
rect 4058 8676 4064 8678
rect 3756 8667 4064 8676
rect 6092 8424 6144 8430
rect 6092 8366 6144 8372
rect 4160 8288 4212 8294
rect 4160 8230 4212 8236
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 3516 8016 3568 8022
rect 3436 7976 3516 8004
rect 3332 7958 3384 7964
rect 3516 7958 3568 7964
rect 4172 7954 4200 8230
rect 3240 7948 3292 7954
rect 3240 7890 3292 7896
rect 4160 7948 4212 7954
rect 4160 7890 4212 7896
rect 3148 7812 3200 7818
rect 3148 7754 3200 7760
rect 3252 7546 3280 7890
rect 3608 7880 3660 7886
rect 3608 7822 3660 7828
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 3240 7540 3292 7546
rect 3240 7482 3292 7488
rect 3620 7478 3648 7822
rect 4252 7744 4304 7750
rect 4252 7686 4304 7692
rect 3756 7644 4064 7653
rect 3756 7642 3762 7644
rect 3818 7642 3842 7644
rect 3898 7642 3922 7644
rect 3978 7642 4002 7644
rect 4058 7642 4064 7644
rect 3818 7590 3820 7642
rect 4000 7590 4002 7642
rect 3756 7588 3762 7590
rect 3818 7588 3842 7590
rect 3898 7588 3922 7590
rect 3978 7588 4002 7590
rect 4058 7588 4064 7590
rect 3756 7579 4064 7588
rect 3608 7472 3660 7478
rect 3528 7432 3608 7460
rect 3056 7268 3108 7274
rect 3056 7210 3108 7216
rect 2964 6996 3016 7002
rect 2964 6938 3016 6944
rect 2872 6928 2924 6934
rect 2872 6870 2924 6876
rect 2504 6860 2556 6866
rect 2504 6802 2556 6808
rect 2136 6656 2188 6662
rect 2136 6598 2188 6604
rect 2228 6656 2280 6662
rect 2228 6598 2280 6604
rect 2148 6458 2176 6598
rect 2240 6458 2268 6598
rect 2516 6458 2544 6802
rect 2136 6452 2188 6458
rect 2136 6394 2188 6400
rect 2228 6452 2280 6458
rect 2228 6394 2280 6400
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 3528 6254 3556 7432
rect 3608 7414 3660 7420
rect 4160 7472 4212 7478
rect 4160 7414 4212 7420
rect 4172 7342 4200 7414
rect 4264 7410 4292 7686
rect 4356 7546 4384 7822
rect 4436 7812 4488 7818
rect 4436 7754 4488 7760
rect 4344 7540 4396 7546
rect 4344 7482 4396 7488
rect 4252 7404 4304 7410
rect 4252 7346 4304 7352
rect 3700 7336 3752 7342
rect 3700 7278 3752 7284
rect 4160 7336 4212 7342
rect 4448 7324 4476 7754
rect 4632 7478 4660 8230
rect 5080 7948 5132 7954
rect 5080 7890 5132 7896
rect 4988 7744 5040 7750
rect 4988 7686 5040 7692
rect 4620 7472 4672 7478
rect 4620 7414 4672 7420
rect 4528 7336 4580 7342
rect 4448 7296 4528 7324
rect 4160 7278 4212 7284
rect 4528 7278 4580 7284
rect 3608 6860 3660 6866
rect 3608 6802 3660 6808
rect 3620 6458 3648 6802
rect 3712 6798 3740 7278
rect 4172 7206 4200 7278
rect 4160 7200 4212 7206
rect 4160 7142 4212 7148
rect 4540 6934 4568 7278
rect 4528 6928 4580 6934
rect 4528 6870 4580 6876
rect 3700 6792 3752 6798
rect 3700 6734 3752 6740
rect 4252 6724 4304 6730
rect 4252 6666 4304 6672
rect 3756 6556 4064 6565
rect 3756 6554 3762 6556
rect 3818 6554 3842 6556
rect 3898 6554 3922 6556
rect 3978 6554 4002 6556
rect 4058 6554 4064 6556
rect 3818 6502 3820 6554
rect 4000 6502 4002 6554
rect 3756 6500 3762 6502
rect 3818 6500 3842 6502
rect 3898 6500 3922 6502
rect 3978 6500 4002 6502
rect 4058 6500 4064 6502
rect 3756 6491 4064 6500
rect 4264 6458 4292 6666
rect 3608 6452 3660 6458
rect 3608 6394 3660 6400
rect 4252 6452 4304 6458
rect 4252 6394 4304 6400
rect 2688 6248 2740 6254
rect 2688 6190 2740 6196
rect 3516 6248 3568 6254
rect 3516 6190 3568 6196
rect 2228 6112 2280 6118
rect 2228 6054 2280 6060
rect 2136 5568 2188 5574
rect 2136 5510 2188 5516
rect 2148 5166 2176 5510
rect 2240 5370 2268 6054
rect 2700 5914 2728 6190
rect 3620 5914 3648 6394
rect 4540 5914 4568 6870
rect 4632 6866 4660 7414
rect 5000 7206 5028 7686
rect 5092 7546 5120 7890
rect 5172 7744 5224 7750
rect 5172 7686 5224 7692
rect 5184 7546 5212 7686
rect 5080 7540 5132 7546
rect 5080 7482 5132 7488
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 5356 7200 5408 7206
rect 5356 7142 5408 7148
rect 5368 6934 5396 7142
rect 5356 6928 5408 6934
rect 5356 6870 5408 6876
rect 6104 6866 6132 8366
rect 8036 8362 8064 8774
rect 8864 8634 8892 9114
rect 9140 8838 9168 10542
rect 9324 9654 9352 11630
rect 9600 11354 9628 12038
rect 9588 11348 9640 11354
rect 9588 11290 9640 11296
rect 9680 11280 9732 11286
rect 9680 11222 9732 11228
rect 9404 11008 9456 11014
rect 9404 10950 9456 10956
rect 9416 10606 9444 10950
rect 9404 10600 9456 10606
rect 9404 10542 9456 10548
rect 9312 9648 9364 9654
rect 9312 9590 9364 9596
rect 9220 9376 9272 9382
rect 9220 9318 9272 9324
rect 9232 9178 9260 9318
rect 9220 9172 9272 9178
rect 9220 9114 9272 9120
rect 9416 9042 9444 10542
rect 9692 10538 9720 11222
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 9784 11014 9812 11154
rect 9772 11008 9824 11014
rect 9772 10950 9824 10956
rect 9680 10532 9732 10538
rect 9680 10474 9732 10480
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9508 9518 9536 10066
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 9968 9466 9996 15914
rect 10888 15706 10916 16390
rect 11072 16250 11100 16594
rect 11244 16448 11296 16454
rect 11244 16390 11296 16396
rect 11060 16244 11112 16250
rect 11060 16186 11112 16192
rect 11152 16244 11204 16250
rect 11152 16186 11204 16192
rect 11060 15972 11112 15978
rect 11164 15960 11192 16186
rect 11256 16046 11284 16390
rect 11428 16244 11480 16250
rect 11428 16186 11480 16192
rect 11336 16176 11388 16182
rect 11336 16118 11388 16124
rect 11348 16046 11376 16118
rect 11244 16040 11296 16046
rect 11244 15982 11296 15988
rect 11336 16040 11388 16046
rect 11336 15982 11388 15988
rect 11112 15932 11192 15960
rect 11060 15914 11112 15920
rect 10876 15700 10928 15706
rect 10876 15642 10928 15648
rect 10324 15564 10376 15570
rect 10324 15506 10376 15512
rect 11244 15564 11296 15570
rect 11244 15506 11296 15512
rect 10232 15156 10284 15162
rect 10232 15098 10284 15104
rect 10244 14822 10272 15098
rect 10232 14816 10284 14822
rect 10232 14758 10284 14764
rect 10232 14544 10284 14550
rect 10232 14486 10284 14492
rect 10244 14385 10272 14486
rect 10230 14376 10286 14385
rect 10230 14311 10286 14320
rect 10336 13734 10364 15506
rect 10472 15260 10780 15269
rect 10472 15258 10478 15260
rect 10534 15258 10558 15260
rect 10614 15258 10638 15260
rect 10694 15258 10718 15260
rect 10774 15258 10780 15260
rect 10534 15206 10536 15258
rect 10716 15206 10718 15258
rect 10472 15204 10478 15206
rect 10534 15204 10558 15206
rect 10614 15204 10638 15206
rect 10694 15204 10718 15206
rect 10774 15204 10780 15206
rect 10472 15195 10780 15204
rect 10876 14952 10928 14958
rect 10876 14894 10928 14900
rect 10508 14816 10560 14822
rect 10508 14758 10560 14764
rect 10520 14362 10548 14758
rect 10428 14346 10548 14362
rect 10416 14340 10548 14346
rect 10468 14334 10548 14340
rect 10416 14282 10468 14288
rect 10472 14172 10780 14181
rect 10472 14170 10478 14172
rect 10534 14170 10558 14172
rect 10614 14170 10638 14172
rect 10694 14170 10718 14172
rect 10774 14170 10780 14172
rect 10534 14118 10536 14170
rect 10716 14118 10718 14170
rect 10472 14116 10478 14118
rect 10534 14116 10558 14118
rect 10614 14116 10638 14118
rect 10694 14116 10718 14118
rect 10774 14116 10780 14118
rect 10472 14107 10780 14116
rect 10324 13728 10376 13734
rect 10324 13670 10376 13676
rect 10784 13728 10836 13734
rect 10784 13670 10836 13676
rect 10796 13326 10824 13670
rect 10888 13326 10916 14894
rect 11060 14544 11112 14550
rect 11060 14486 11112 14492
rect 10968 14408 11020 14414
rect 10968 14350 11020 14356
rect 10980 13530 11008 14350
rect 11072 14074 11100 14486
rect 11256 14346 11284 15506
rect 11440 14770 11468 16186
rect 11900 16046 11928 16934
rect 11888 16040 11940 16046
rect 11888 15982 11940 15988
rect 11704 15904 11756 15910
rect 11704 15846 11756 15852
rect 11716 14890 11744 15846
rect 11704 14884 11756 14890
rect 11704 14826 11756 14832
rect 11348 14742 11468 14770
rect 11244 14340 11296 14346
rect 11244 14282 11296 14288
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 11348 13954 11376 14742
rect 11612 14272 11664 14278
rect 11612 14214 11664 14220
rect 11256 13926 11376 13954
rect 11060 13728 11112 13734
rect 11060 13670 11112 13676
rect 10968 13524 11020 13530
rect 10968 13466 11020 13472
rect 11072 13394 11100 13670
rect 11060 13388 11112 13394
rect 11060 13330 11112 13336
rect 10784 13320 10836 13326
rect 10784 13262 10836 13268
rect 10876 13320 10928 13326
rect 10876 13262 10928 13268
rect 10472 13084 10780 13093
rect 10472 13082 10478 13084
rect 10534 13082 10558 13084
rect 10614 13082 10638 13084
rect 10694 13082 10718 13084
rect 10774 13082 10780 13084
rect 10534 13030 10536 13082
rect 10716 13030 10718 13082
rect 10472 13028 10478 13030
rect 10534 13028 10558 13030
rect 10614 13028 10638 13030
rect 10694 13028 10718 13030
rect 10774 13028 10780 13030
rect 10472 13019 10780 13028
rect 10888 12714 10916 13262
rect 10968 13184 11020 13190
rect 10968 13126 11020 13132
rect 10980 12986 11008 13126
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 10876 12708 10928 12714
rect 10876 12650 10928 12656
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 10152 12442 10180 12582
rect 10140 12436 10192 12442
rect 11256 12434 11284 13926
rect 11336 13864 11388 13870
rect 11388 13824 11560 13852
rect 11336 13806 11388 13812
rect 11256 12406 11376 12434
rect 10140 12378 10192 12384
rect 11060 12300 11112 12306
rect 11060 12242 11112 12248
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 10060 11354 10088 12174
rect 10324 12096 10376 12102
rect 10324 12038 10376 12044
rect 10336 11626 10364 12038
rect 10472 11996 10780 12005
rect 10472 11994 10478 11996
rect 10534 11994 10558 11996
rect 10614 11994 10638 11996
rect 10694 11994 10718 11996
rect 10774 11994 10780 11996
rect 10534 11942 10536 11994
rect 10716 11942 10718 11994
rect 10472 11940 10478 11942
rect 10534 11940 10558 11942
rect 10614 11940 10638 11942
rect 10694 11940 10718 11942
rect 10774 11940 10780 11942
rect 10472 11931 10780 11940
rect 11072 11762 11100 12242
rect 11060 11756 11112 11762
rect 10980 11716 11060 11744
rect 10324 11620 10376 11626
rect 10324 11562 10376 11568
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 10060 10810 10088 11154
rect 10232 11008 10284 11014
rect 10232 10950 10284 10956
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 10244 10674 10272 10950
rect 10472 10908 10780 10917
rect 10472 10906 10478 10908
rect 10534 10906 10558 10908
rect 10614 10906 10638 10908
rect 10694 10906 10718 10908
rect 10774 10906 10780 10908
rect 10534 10854 10536 10906
rect 10716 10854 10718 10906
rect 10472 10852 10478 10854
rect 10534 10852 10558 10854
rect 10614 10852 10638 10854
rect 10694 10852 10718 10854
rect 10774 10852 10780 10854
rect 10472 10843 10780 10852
rect 10232 10668 10284 10674
rect 10232 10610 10284 10616
rect 10140 10600 10192 10606
rect 10140 10542 10192 10548
rect 10876 10600 10928 10606
rect 10876 10542 10928 10548
rect 10152 10266 10180 10542
rect 10784 10464 10836 10470
rect 10784 10406 10836 10412
rect 10796 10266 10824 10406
rect 10140 10260 10192 10266
rect 10140 10202 10192 10208
rect 10784 10260 10836 10266
rect 10784 10202 10836 10208
rect 10152 9586 10180 10202
rect 10888 10198 10916 10542
rect 10876 10192 10928 10198
rect 10876 10134 10928 10140
rect 10980 10130 11008 11716
rect 11060 11698 11112 11704
rect 11244 11552 11296 11558
rect 11244 11494 11296 11500
rect 11256 11218 11284 11494
rect 11244 11212 11296 11218
rect 11244 11154 11296 11160
rect 11060 11076 11112 11082
rect 11060 11018 11112 11024
rect 11072 10130 11100 11018
rect 10968 10124 11020 10130
rect 10968 10066 11020 10072
rect 11060 10124 11112 10130
rect 11060 10066 11112 10072
rect 10472 9820 10780 9829
rect 10472 9818 10478 9820
rect 10534 9818 10558 9820
rect 10614 9818 10638 9820
rect 10694 9818 10718 9820
rect 10774 9818 10780 9820
rect 10534 9766 10536 9818
rect 10716 9766 10718 9818
rect 10472 9764 10478 9766
rect 10534 9764 10558 9766
rect 10614 9764 10638 9766
rect 10694 9764 10718 9766
rect 10774 9764 10780 9766
rect 10472 9755 10780 9764
rect 11072 9722 11100 10066
rect 10968 9716 11020 9722
rect 10968 9658 11020 9664
rect 11060 9716 11112 9722
rect 11060 9658 11112 9664
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 9508 9382 9536 9454
rect 9968 9438 10088 9466
rect 9496 9376 9548 9382
rect 9496 9318 9548 9324
rect 9956 9376 10008 9382
rect 9956 9318 10008 9324
rect 9508 9110 9536 9318
rect 9496 9104 9548 9110
rect 9496 9046 9548 9052
rect 9404 9036 9456 9042
rect 9404 8978 9456 8984
rect 9508 8974 9536 9046
rect 9968 9042 9996 9318
rect 9956 9036 10008 9042
rect 9956 8978 10008 8984
rect 9496 8968 9548 8974
rect 9496 8910 9548 8916
rect 9128 8832 9180 8838
rect 9128 8774 9180 8780
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 8852 8628 8904 8634
rect 8852 8570 8904 8576
rect 9220 8424 9272 8430
rect 9220 8366 9272 8372
rect 6368 8356 6420 8362
rect 6368 8298 6420 8304
rect 8024 8356 8076 8362
rect 8024 8298 8076 8304
rect 6380 8090 6408 8298
rect 6644 8288 6696 8294
rect 6644 8230 6696 8236
rect 6368 8084 6420 8090
rect 6368 8026 6420 8032
rect 6656 6866 6684 8230
rect 7114 8188 7422 8197
rect 7114 8186 7120 8188
rect 7176 8186 7200 8188
rect 7256 8186 7280 8188
rect 7336 8186 7360 8188
rect 7416 8186 7422 8188
rect 7176 8134 7178 8186
rect 7358 8134 7360 8186
rect 7114 8132 7120 8134
rect 7176 8132 7200 8134
rect 7256 8132 7280 8134
rect 7336 8132 7360 8134
rect 7416 8132 7422 8134
rect 7114 8123 7422 8132
rect 6828 7948 6880 7954
rect 6828 7890 6880 7896
rect 6840 7546 6868 7890
rect 8852 7880 8904 7886
rect 8852 7822 8904 7828
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 8864 7410 8892 7822
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 8852 7404 8904 7410
rect 8852 7346 8904 7352
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 6932 6866 6960 7278
rect 7024 7002 7052 7346
rect 8668 7336 8720 7342
rect 8668 7278 8720 7284
rect 7472 7268 7524 7274
rect 7472 7210 7524 7216
rect 7114 7100 7422 7109
rect 7114 7098 7120 7100
rect 7176 7098 7200 7100
rect 7256 7098 7280 7100
rect 7336 7098 7360 7100
rect 7416 7098 7422 7100
rect 7176 7046 7178 7098
rect 7358 7046 7360 7098
rect 7114 7044 7120 7046
rect 7176 7044 7200 7046
rect 7256 7044 7280 7046
rect 7336 7044 7360 7046
rect 7416 7044 7422 7046
rect 7114 7035 7422 7044
rect 7484 7002 7512 7210
rect 8484 7200 8536 7206
rect 8484 7142 8536 7148
rect 7012 6996 7064 7002
rect 7012 6938 7064 6944
rect 7472 6996 7524 7002
rect 7472 6938 7524 6944
rect 8496 6866 8524 7142
rect 4620 6860 4672 6866
rect 4620 6802 4672 6808
rect 6092 6860 6144 6866
rect 6092 6802 6144 6808
rect 6184 6860 6236 6866
rect 6644 6860 6696 6866
rect 6184 6802 6236 6808
rect 6564 6820 6644 6848
rect 6196 6458 6224 6802
rect 6184 6452 6236 6458
rect 6184 6394 6236 6400
rect 6564 6254 6592 6820
rect 6644 6802 6696 6808
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 8484 6860 8536 6866
rect 8484 6802 8536 6808
rect 8576 6860 8628 6866
rect 8576 6802 8628 6808
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 6656 6458 6684 6598
rect 6932 6458 6960 6802
rect 8588 6662 8616 6802
rect 7932 6656 7984 6662
rect 7932 6598 7984 6604
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6920 6452 6972 6458
rect 6920 6394 6972 6400
rect 7748 6316 7800 6322
rect 7748 6258 7800 6264
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 5816 6248 5868 6254
rect 5816 6190 5868 6196
rect 6552 6248 6604 6254
rect 6552 6190 6604 6196
rect 6736 6248 6788 6254
rect 6736 6190 6788 6196
rect 4816 5914 4844 6190
rect 5828 5914 5856 6190
rect 6748 5914 6776 6190
rect 7114 6012 7422 6021
rect 7114 6010 7120 6012
rect 7176 6010 7200 6012
rect 7256 6010 7280 6012
rect 7336 6010 7360 6012
rect 7416 6010 7422 6012
rect 7176 5958 7178 6010
rect 7358 5958 7360 6010
rect 7114 5956 7120 5958
rect 7176 5956 7200 5958
rect 7256 5956 7280 5958
rect 7336 5956 7360 5958
rect 7416 5956 7422 5958
rect 7114 5947 7422 5956
rect 7760 5914 7788 6258
rect 2688 5908 2740 5914
rect 2688 5850 2740 5856
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 4528 5908 4580 5914
rect 4528 5850 4580 5856
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 5816 5908 5868 5914
rect 5816 5850 5868 5856
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 7944 5778 7972 6598
rect 8680 6458 8708 7278
rect 9232 6866 9260 8366
rect 9496 8356 9548 8362
rect 9496 8298 9548 8304
rect 9508 8090 9536 8298
rect 9692 8090 9720 8774
rect 9496 8084 9548 8090
rect 9496 8026 9548 8032
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 9862 7304 9918 7313
rect 9862 7239 9864 7248
rect 9916 7239 9918 7248
rect 9864 7210 9916 7216
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9220 6860 9272 6866
rect 9220 6802 9272 6808
rect 9232 6458 9260 6802
rect 9692 6798 9720 7142
rect 10060 7002 10088 9438
rect 10324 9444 10376 9450
rect 10324 9386 10376 9392
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 10152 9042 10180 9318
rect 10140 9036 10192 9042
rect 10140 8978 10192 8984
rect 10336 8634 10364 9386
rect 10472 8732 10780 8741
rect 10472 8730 10478 8732
rect 10534 8730 10558 8732
rect 10614 8730 10638 8732
rect 10694 8730 10718 8732
rect 10774 8730 10780 8732
rect 10534 8678 10536 8730
rect 10716 8678 10718 8730
rect 10472 8676 10478 8678
rect 10534 8676 10558 8678
rect 10614 8676 10638 8678
rect 10694 8676 10718 8678
rect 10774 8676 10780 8678
rect 10472 8667 10780 8676
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 10980 8430 11008 9658
rect 11072 9042 11100 9658
rect 11060 9036 11112 9042
rect 11060 8978 11112 8984
rect 11072 8498 11100 8978
rect 11060 8492 11112 8498
rect 11060 8434 11112 8440
rect 10968 8424 11020 8430
rect 10968 8366 11020 8372
rect 10472 7644 10780 7653
rect 10472 7642 10478 7644
rect 10534 7642 10558 7644
rect 10614 7642 10638 7644
rect 10694 7642 10718 7644
rect 10774 7642 10780 7644
rect 10534 7590 10536 7642
rect 10716 7590 10718 7642
rect 10472 7588 10478 7590
rect 10534 7588 10558 7590
rect 10614 7588 10638 7590
rect 10694 7588 10718 7590
rect 10774 7588 10780 7590
rect 10472 7579 10780 7588
rect 10140 7336 10192 7342
rect 10140 7278 10192 7284
rect 10324 7336 10376 7342
rect 10324 7278 10376 7284
rect 10508 7336 10560 7342
rect 10508 7278 10560 7284
rect 10048 6996 10100 7002
rect 10048 6938 10100 6944
rect 10152 6866 10180 7278
rect 10336 7002 10364 7278
rect 10324 6996 10376 7002
rect 10324 6938 10376 6944
rect 10520 6934 10548 7278
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 11072 6934 11100 7142
rect 10508 6928 10560 6934
rect 10508 6870 10560 6876
rect 11060 6928 11112 6934
rect 11060 6870 11112 6876
rect 10140 6860 10192 6866
rect 10140 6802 10192 6808
rect 10232 6860 10284 6866
rect 10232 6802 10284 6808
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 9220 6452 9272 6458
rect 9220 6394 9272 6400
rect 8116 6384 8168 6390
rect 8116 6326 8168 6332
rect 8300 6384 8352 6390
rect 8300 6326 8352 6332
rect 8128 5914 8156 6326
rect 8208 6112 8260 6118
rect 8208 6054 8260 6060
rect 8116 5908 8168 5914
rect 8116 5850 8168 5856
rect 2320 5772 2372 5778
rect 2320 5714 2372 5720
rect 2964 5772 3016 5778
rect 2964 5714 3016 5720
rect 5264 5772 5316 5778
rect 5264 5714 5316 5720
rect 6092 5772 6144 5778
rect 6092 5714 6144 5720
rect 7656 5772 7708 5778
rect 7656 5714 7708 5720
rect 7932 5772 7984 5778
rect 7932 5714 7984 5720
rect 2228 5364 2280 5370
rect 2228 5306 2280 5312
rect 2136 5160 2188 5166
rect 2136 5102 2188 5108
rect 1124 4820 1176 4826
rect 1124 4762 1176 4768
rect 1952 4820 2004 4826
rect 1952 4762 2004 4768
rect 2136 4684 2188 4690
rect 2136 4626 2188 4632
rect 2148 3942 2176 4626
rect 2228 4072 2280 4078
rect 2228 4014 2280 4020
rect 2136 3936 2188 3942
rect 2136 3878 2188 3884
rect 2044 3460 2096 3466
rect 2044 3402 2096 3408
rect 2056 2990 2084 3402
rect 2240 3194 2268 4014
rect 2332 4010 2360 5714
rect 2596 5704 2648 5710
rect 2596 5646 2648 5652
rect 2608 4758 2636 5646
rect 2976 5370 3004 5714
rect 3240 5568 3292 5574
rect 3240 5510 3292 5516
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 2596 4752 2648 4758
rect 2596 4694 2648 4700
rect 3056 4684 3108 4690
rect 3056 4626 3108 4632
rect 2596 4616 2648 4622
rect 2596 4558 2648 4564
rect 2608 4078 2636 4558
rect 3068 4214 3096 4626
rect 3056 4208 3108 4214
rect 3056 4150 3108 4156
rect 2596 4072 2648 4078
rect 2596 4014 2648 4020
rect 2962 4040 3018 4049
rect 2320 4004 2372 4010
rect 2320 3946 2372 3952
rect 2780 4004 2832 4010
rect 2962 3975 3018 3984
rect 2780 3946 2832 3952
rect 2228 3188 2280 3194
rect 2228 3130 2280 3136
rect 2792 3058 2820 3946
rect 2976 3738 3004 3975
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 3056 3732 3108 3738
rect 3056 3674 3108 3680
rect 3068 3058 3096 3674
rect 3252 3466 3280 5510
rect 3756 5468 4064 5477
rect 3756 5466 3762 5468
rect 3818 5466 3842 5468
rect 3898 5466 3922 5468
rect 3978 5466 4002 5468
rect 4058 5466 4064 5468
rect 3818 5414 3820 5466
rect 4000 5414 4002 5466
rect 3756 5412 3762 5414
rect 3818 5412 3842 5414
rect 3898 5412 3922 5414
rect 3978 5412 4002 5414
rect 4058 5412 4064 5414
rect 3756 5403 4064 5412
rect 5276 5370 5304 5714
rect 6104 5370 6132 5714
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 6932 5370 6960 5510
rect 7668 5370 7696 5714
rect 5264 5364 5316 5370
rect 5264 5306 5316 5312
rect 6092 5364 6144 5370
rect 6092 5306 6144 5312
rect 6920 5364 6972 5370
rect 6920 5306 6972 5312
rect 7656 5364 7708 5370
rect 7656 5306 7708 5312
rect 3332 5160 3384 5166
rect 3332 5102 3384 5108
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 5724 5160 5776 5166
rect 5724 5102 5776 5108
rect 6368 5160 6420 5166
rect 6368 5102 6420 5108
rect 3344 4690 3372 5102
rect 3424 5024 3476 5030
rect 3424 4966 3476 4972
rect 3332 4684 3384 4690
rect 3332 4626 3384 4632
rect 3344 4146 3372 4626
rect 3436 4554 3464 4966
rect 4160 4752 4212 4758
rect 4160 4694 4212 4700
rect 3516 4684 3568 4690
rect 3568 4644 3648 4672
rect 3516 4626 3568 4632
rect 3424 4548 3476 4554
rect 3424 4490 3476 4496
rect 3424 4208 3476 4214
rect 3424 4150 3476 4156
rect 3332 4140 3384 4146
rect 3332 4082 3384 4088
rect 3344 3602 3372 4082
rect 3436 3602 3464 4150
rect 3516 4072 3568 4078
rect 3620 4049 3648 4644
rect 3756 4380 4064 4389
rect 3756 4378 3762 4380
rect 3818 4378 3842 4380
rect 3898 4378 3922 4380
rect 3978 4378 4002 4380
rect 4058 4378 4064 4380
rect 3818 4326 3820 4378
rect 4000 4326 4002 4378
rect 3756 4324 3762 4326
rect 3818 4324 3842 4326
rect 3898 4324 3922 4326
rect 3978 4324 4002 4326
rect 4058 4324 4064 4326
rect 3756 4315 4064 4324
rect 4172 4078 4200 4694
rect 4344 4684 4396 4690
rect 4344 4626 4396 4632
rect 4804 4684 4856 4690
rect 4804 4626 4856 4632
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 4264 4282 4292 4558
rect 4252 4276 4304 4282
rect 4252 4218 4304 4224
rect 4160 4072 4212 4078
rect 3516 4014 3568 4020
rect 3606 4040 3662 4049
rect 3332 3596 3384 3602
rect 3332 3538 3384 3544
rect 3424 3596 3476 3602
rect 3424 3538 3476 3544
rect 3240 3460 3292 3466
rect 3240 3402 3292 3408
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 3056 3052 3108 3058
rect 3056 2994 3108 3000
rect 3252 2990 3280 3402
rect 2044 2984 2096 2990
rect 2044 2926 2096 2932
rect 2412 2984 2464 2990
rect 2412 2926 2464 2932
rect 3240 2984 3292 2990
rect 3240 2926 3292 2932
rect 1308 2848 1360 2854
rect 1308 2790 1360 2796
rect 2044 2848 2096 2854
rect 2044 2790 2096 2796
rect 940 1896 992 1902
rect 940 1838 992 1844
rect 1124 1896 1176 1902
rect 1124 1838 1176 1844
rect 952 882 980 1838
rect 1136 1426 1164 1838
rect 1320 1562 1348 2790
rect 2056 1562 2084 2790
rect 2424 2514 2452 2926
rect 2504 2916 2556 2922
rect 2504 2858 2556 2864
rect 2412 2508 2464 2514
rect 2412 2450 2464 2456
rect 1308 1556 1360 1562
rect 1308 1498 1360 1504
rect 2044 1556 2096 1562
rect 2044 1498 2096 1504
rect 1124 1420 1176 1426
rect 1124 1362 1176 1368
rect 2320 1420 2372 1426
rect 2320 1362 2372 1368
rect 2136 1352 2188 1358
rect 2136 1294 2188 1300
rect 2148 1018 2176 1294
rect 2136 1012 2188 1018
rect 2136 954 2188 960
rect 940 876 992 882
rect 940 818 992 824
rect 1768 808 1820 814
rect 1768 750 1820 756
rect 1780 400 1808 750
rect 2332 400 2360 1362
rect 2516 814 2544 2858
rect 2688 2848 2740 2854
rect 2688 2790 2740 2796
rect 2700 2514 2728 2790
rect 2688 2508 2740 2514
rect 2688 2450 2740 2456
rect 2688 2372 2740 2378
rect 2688 2314 2740 2320
rect 2700 1902 2728 2314
rect 3528 1902 3556 4014
rect 4160 4014 4212 4020
rect 4264 4010 4292 4218
rect 4356 4162 4384 4626
rect 4436 4548 4488 4554
rect 4436 4490 4488 4496
rect 4448 4282 4476 4490
rect 4436 4276 4488 4282
rect 4436 4218 4488 4224
rect 4356 4134 4476 4162
rect 3606 3975 3662 3984
rect 4068 4004 4120 4010
rect 4068 3946 4120 3952
rect 4252 4004 4304 4010
rect 4252 3946 4304 3952
rect 4344 4004 4396 4010
rect 4344 3946 4396 3952
rect 4080 3584 4108 3946
rect 4160 3596 4212 3602
rect 4080 3556 4160 3584
rect 4160 3538 4212 3544
rect 3756 3292 4064 3301
rect 3756 3290 3762 3292
rect 3818 3290 3842 3292
rect 3898 3290 3922 3292
rect 3978 3290 4002 3292
rect 4058 3290 4064 3292
rect 3818 3238 3820 3290
rect 4000 3238 4002 3290
rect 3756 3236 3762 3238
rect 3818 3236 3842 3238
rect 3898 3236 3922 3238
rect 3978 3236 4002 3238
rect 4058 3236 4064 3238
rect 3756 3227 4064 3236
rect 3792 3052 3844 3058
rect 3792 2994 3844 3000
rect 3804 2446 3832 2994
rect 4264 2854 4292 3946
rect 4356 3602 4384 3946
rect 4344 3596 4396 3602
rect 4344 3538 4396 3544
rect 4448 3534 4476 4134
rect 4816 4078 4844 4626
rect 4896 4276 4948 4282
rect 4896 4218 4948 4224
rect 4908 4078 4936 4218
rect 4988 4208 5040 4214
rect 4988 4150 5040 4156
rect 4804 4072 4856 4078
rect 4804 4014 4856 4020
rect 4896 4072 4948 4078
rect 4896 4014 4948 4020
rect 4896 3936 4948 3942
rect 4896 3878 4948 3884
rect 4528 3596 4580 3602
rect 4528 3538 4580 3544
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 4436 3528 4488 3534
rect 4356 3476 4436 3482
rect 4356 3470 4488 3476
rect 4356 3454 4476 3470
rect 4356 2922 4384 3454
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 4344 2916 4396 2922
rect 4344 2858 4396 2864
rect 4252 2848 4304 2854
rect 4252 2790 4304 2796
rect 4448 2553 4476 3334
rect 4434 2544 4490 2553
rect 4356 2514 4434 2530
rect 4344 2508 4434 2514
rect 4396 2502 4434 2508
rect 4540 2514 4568 3538
rect 4724 2650 4752 3538
rect 4908 2836 4936 3878
rect 5000 3505 5028 4150
rect 5092 3738 5120 5102
rect 5736 4826 5764 5102
rect 5724 4820 5776 4826
rect 5724 4762 5776 4768
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 5448 4480 5500 4486
rect 5448 4422 5500 4428
rect 5460 4078 5488 4422
rect 5448 4072 5500 4078
rect 5448 4014 5500 4020
rect 5264 3936 5316 3942
rect 5264 3878 5316 3884
rect 5448 3936 5500 3942
rect 5448 3878 5500 3884
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 4986 3496 5042 3505
rect 4986 3431 5042 3440
rect 5276 3126 5304 3878
rect 5264 3120 5316 3126
rect 5264 3062 5316 3068
rect 5276 2922 5304 3062
rect 5264 2916 5316 2922
rect 5264 2858 5316 2864
rect 4908 2808 5120 2836
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 4434 2479 4490 2488
rect 4528 2508 4580 2514
rect 4344 2450 4396 2456
rect 4528 2450 4580 2456
rect 3792 2440 3844 2446
rect 3792 2382 3844 2388
rect 3608 2304 3660 2310
rect 3608 2246 3660 2252
rect 4160 2304 4212 2310
rect 4160 2246 4212 2252
rect 4620 2304 4672 2310
rect 4620 2246 4672 2252
rect 2688 1896 2740 1902
rect 2964 1896 3016 1902
rect 2688 1838 2740 1844
rect 2884 1856 2964 1884
rect 2504 808 2556 814
rect 2504 750 2556 756
rect 2884 400 2912 1856
rect 2964 1838 3016 1844
rect 3332 1896 3384 1902
rect 3332 1838 3384 1844
rect 3516 1896 3568 1902
rect 3516 1838 3568 1844
rect 3240 1420 3292 1426
rect 3240 1362 3292 1368
rect 3252 762 3280 1362
rect 3344 1358 3372 1838
rect 3516 1760 3568 1766
rect 3516 1702 3568 1708
rect 3528 1562 3556 1702
rect 3516 1556 3568 1562
rect 3516 1498 3568 1504
rect 3332 1352 3384 1358
rect 3332 1294 3384 1300
rect 3620 814 3648 2246
rect 3756 2204 4064 2213
rect 3756 2202 3762 2204
rect 3818 2202 3842 2204
rect 3898 2202 3922 2204
rect 3978 2202 4002 2204
rect 4058 2202 4064 2204
rect 3818 2150 3820 2202
rect 4000 2150 4002 2202
rect 3756 2148 3762 2150
rect 3818 2148 3842 2150
rect 3898 2148 3922 2150
rect 3978 2148 4002 2150
rect 4058 2148 4064 2150
rect 3756 2139 4064 2148
rect 4068 2100 4120 2106
rect 4172 2088 4200 2246
rect 4120 2060 4200 2088
rect 4068 2042 4120 2048
rect 4068 1828 4120 1834
rect 4068 1770 4120 1776
rect 4080 1306 4108 1770
rect 4436 1420 4488 1426
rect 4488 1380 4568 1408
rect 4436 1362 4488 1368
rect 4080 1278 4200 1306
rect 3756 1116 4064 1125
rect 3756 1114 3762 1116
rect 3818 1114 3842 1116
rect 3898 1114 3922 1116
rect 3978 1114 4002 1116
rect 4058 1114 4064 1116
rect 3818 1062 3820 1114
rect 4000 1062 4002 1114
rect 3756 1060 3762 1062
rect 3818 1060 3842 1062
rect 3898 1060 3922 1062
rect 3978 1060 4002 1062
rect 4058 1060 4064 1062
rect 3756 1051 4064 1060
rect 4172 1018 4200 1278
rect 4160 1012 4212 1018
rect 4160 954 4212 960
rect 3608 808 3660 814
rect 3252 734 3464 762
rect 4068 808 4120 814
rect 3608 750 3660 756
rect 3988 768 4068 796
rect 3436 400 3464 734
rect 3988 400 4016 768
rect 4068 750 4120 756
rect 4540 400 4568 1380
rect 4632 814 4660 2246
rect 4724 1426 4752 2586
rect 5092 2514 5120 2808
rect 5460 2553 5488 3878
rect 5446 2544 5502 2553
rect 4896 2508 4948 2514
rect 4896 2450 4948 2456
rect 5080 2508 5132 2514
rect 5446 2479 5502 2488
rect 5080 2450 5132 2456
rect 4804 2304 4856 2310
rect 4804 2246 4856 2252
rect 4816 2106 4844 2246
rect 4908 2106 4936 2450
rect 5552 2310 5580 4626
rect 6000 4616 6052 4622
rect 6000 4558 6052 4564
rect 5816 4072 5868 4078
rect 5816 4014 5868 4020
rect 5828 3534 5856 4014
rect 6012 3942 6040 4558
rect 6380 4282 6408 5102
rect 7114 4924 7422 4933
rect 7114 4922 7120 4924
rect 7176 4922 7200 4924
rect 7256 4922 7280 4924
rect 7336 4922 7360 4924
rect 7416 4922 7422 4924
rect 7176 4870 7178 4922
rect 7358 4870 7360 4922
rect 7114 4868 7120 4870
rect 7176 4868 7200 4870
rect 7256 4868 7280 4870
rect 7336 4868 7360 4870
rect 7416 4868 7422 4870
rect 7114 4859 7422 4868
rect 8220 4826 8248 6054
rect 8312 5778 8340 6326
rect 9692 5914 9720 6734
rect 9680 5908 9732 5914
rect 9680 5850 9732 5856
rect 9496 5840 9548 5846
rect 9496 5782 9548 5788
rect 8300 5772 8352 5778
rect 8300 5714 8352 5720
rect 8852 5228 8904 5234
rect 8852 5170 8904 5176
rect 8576 5160 8628 5166
rect 8576 5102 8628 5108
rect 8484 5024 8536 5030
rect 8484 4966 8536 4972
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 8300 4752 8352 4758
rect 8300 4694 8352 4700
rect 8024 4616 8076 4622
rect 8024 4558 8076 4564
rect 7012 4480 7064 4486
rect 7012 4422 7064 4428
rect 6368 4276 6420 4282
rect 6368 4218 6420 4224
rect 6460 4208 6512 4214
rect 6460 4150 6512 4156
rect 6184 4004 6236 4010
rect 6184 3946 6236 3952
rect 6000 3936 6052 3942
rect 6000 3878 6052 3884
rect 5816 3528 5868 3534
rect 5816 3470 5868 3476
rect 5632 2508 5684 2514
rect 5632 2450 5684 2456
rect 5540 2304 5592 2310
rect 5540 2246 5592 2252
rect 5644 2106 5672 2450
rect 4804 2100 4856 2106
rect 4804 2042 4856 2048
rect 4896 2100 4948 2106
rect 4896 2042 4948 2048
rect 5632 2100 5684 2106
rect 5632 2042 5684 2048
rect 5828 1902 5856 3470
rect 6196 2836 6224 3946
rect 6276 3528 6328 3534
rect 6276 3470 6328 3476
rect 6288 3194 6316 3470
rect 6472 3398 6500 4150
rect 7024 4078 7052 4422
rect 8036 4282 8064 4558
rect 8024 4276 8076 4282
rect 8024 4218 8076 4224
rect 6736 4072 6788 4078
rect 6736 4014 6788 4020
rect 7012 4072 7064 4078
rect 7012 4014 7064 4020
rect 7654 4040 7710 4049
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 6656 3602 6684 3878
rect 6748 3738 6776 4014
rect 7654 3975 7710 3984
rect 7114 3836 7422 3845
rect 7114 3834 7120 3836
rect 7176 3834 7200 3836
rect 7256 3834 7280 3836
rect 7336 3834 7360 3836
rect 7416 3834 7422 3836
rect 7176 3782 7178 3834
rect 7358 3782 7360 3834
rect 7114 3780 7120 3782
rect 7176 3780 7200 3782
rect 7256 3780 7280 3782
rect 7336 3780 7360 3782
rect 7416 3780 7422 3782
rect 7114 3771 7422 3780
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 6644 3596 6696 3602
rect 6644 3538 6696 3544
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 6368 3392 6420 3398
rect 6368 3334 6420 3340
rect 6460 3392 6512 3398
rect 6460 3334 6512 3340
rect 6276 3188 6328 3194
rect 6276 3130 6328 3136
rect 6380 2854 6408 3334
rect 6276 2848 6328 2854
rect 6196 2808 6276 2836
rect 6276 2790 6328 2796
rect 6368 2848 6420 2854
rect 6368 2790 6420 2796
rect 6092 2304 6144 2310
rect 6092 2246 6144 2252
rect 5172 1896 5224 1902
rect 5092 1856 5172 1884
rect 4712 1420 4764 1426
rect 4712 1362 4764 1368
rect 4620 808 4672 814
rect 4620 750 4672 756
rect 5092 400 5120 1856
rect 5172 1838 5224 1844
rect 5264 1896 5316 1902
rect 5264 1838 5316 1844
rect 5724 1896 5776 1902
rect 5724 1838 5776 1844
rect 5816 1896 5868 1902
rect 5816 1838 5868 1844
rect 5276 1426 5304 1838
rect 5736 1426 5764 1838
rect 5264 1420 5316 1426
rect 5264 1362 5316 1368
rect 5724 1420 5776 1426
rect 5724 1362 5776 1368
rect 6104 814 6132 2246
rect 6288 1562 6316 2790
rect 6472 2650 6500 3334
rect 6644 2984 6696 2990
rect 6644 2926 6696 2932
rect 6656 2650 6684 2926
rect 6460 2644 6512 2650
rect 6460 2586 6512 2592
rect 6644 2644 6696 2650
rect 6644 2586 6696 2592
rect 6458 2544 6514 2553
rect 6458 2479 6460 2488
rect 6512 2479 6514 2488
rect 6460 2450 6512 2456
rect 6656 2106 6684 2586
rect 6840 2446 6868 3538
rect 7194 3496 7250 3505
rect 7194 3431 7250 3440
rect 6920 3392 6972 3398
rect 6920 3334 6972 3340
rect 6932 3126 6960 3334
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 6920 3120 6972 3126
rect 6920 3062 6972 3068
rect 7024 2774 7052 3130
rect 7208 2922 7236 3431
rect 7380 3392 7432 3398
rect 7380 3334 7432 3340
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 7392 2990 7420 3334
rect 7484 3194 7512 3334
rect 7472 3188 7524 3194
rect 7472 3130 7524 3136
rect 7380 2984 7432 2990
rect 7380 2926 7432 2932
rect 7196 2916 7248 2922
rect 7196 2858 7248 2864
rect 6932 2746 7052 2774
rect 7114 2748 7422 2757
rect 7114 2746 7120 2748
rect 7176 2746 7200 2748
rect 7256 2746 7280 2748
rect 7336 2746 7360 2748
rect 7416 2746 7422 2748
rect 6828 2440 6880 2446
rect 6828 2382 6880 2388
rect 6644 2100 6696 2106
rect 6644 2042 6696 2048
rect 6644 1896 6696 1902
rect 6644 1838 6696 1844
rect 6276 1556 6328 1562
rect 6276 1498 6328 1504
rect 6184 1488 6236 1494
rect 6184 1430 6236 1436
rect 5540 808 5592 814
rect 6092 808 6144 814
rect 5592 768 5672 796
rect 5540 750 5592 756
rect 5644 400 5672 768
rect 6092 750 6144 756
rect 6196 400 6224 1430
rect 6276 1216 6328 1222
rect 6276 1158 6328 1164
rect 6288 1018 6316 1158
rect 6276 1012 6328 1018
rect 6276 954 6328 960
rect 6656 490 6684 1838
rect 6932 1408 6960 2746
rect 7176 2694 7178 2746
rect 7358 2694 7360 2746
rect 7114 2692 7120 2694
rect 7176 2692 7200 2694
rect 7256 2692 7280 2694
rect 7336 2692 7360 2694
rect 7416 2692 7422 2694
rect 7114 2683 7422 2692
rect 7668 2514 7696 3975
rect 8312 3942 8340 4694
rect 8496 4554 8524 4966
rect 8588 4758 8616 5102
rect 8760 5024 8812 5030
rect 8760 4966 8812 4972
rect 8772 4826 8800 4966
rect 8760 4820 8812 4826
rect 8760 4762 8812 4768
rect 8576 4752 8628 4758
rect 8576 4694 8628 4700
rect 8484 4548 8536 4554
rect 8484 4490 8536 4496
rect 8496 4282 8524 4490
rect 8484 4276 8536 4282
rect 8484 4218 8536 4224
rect 8588 4078 8616 4694
rect 8864 4690 8892 5170
rect 9036 4752 9088 4758
rect 9036 4694 9088 4700
rect 8852 4684 8904 4690
rect 8852 4626 8904 4632
rect 8864 4078 8892 4626
rect 8576 4072 8628 4078
rect 8576 4014 8628 4020
rect 8852 4072 8904 4078
rect 8852 4014 8904 4020
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 8576 3596 8628 3602
rect 8576 3538 8628 3544
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8220 3194 8248 3470
rect 8588 3194 8616 3538
rect 8852 3392 8904 3398
rect 8852 3334 8904 3340
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 8576 3188 8628 3194
rect 8576 3130 8628 3136
rect 8300 2848 8352 2854
rect 8300 2790 8352 2796
rect 7656 2508 7708 2514
rect 7656 2450 7708 2456
rect 7012 2304 7064 2310
rect 7012 2246 7064 2252
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7024 2106 7052 2246
rect 7012 2100 7064 2106
rect 7012 2042 7064 2048
rect 7116 1902 7144 2246
rect 7104 1896 7156 1902
rect 7104 1838 7156 1844
rect 7840 1896 7892 1902
rect 7840 1838 7892 1844
rect 7932 1896 7984 1902
rect 7932 1838 7984 1844
rect 7114 1660 7422 1669
rect 7114 1658 7120 1660
rect 7176 1658 7200 1660
rect 7256 1658 7280 1660
rect 7336 1658 7360 1660
rect 7416 1658 7422 1660
rect 7176 1606 7178 1658
rect 7358 1606 7360 1658
rect 7114 1604 7120 1606
rect 7176 1604 7200 1606
rect 7256 1604 7280 1606
rect 7336 1604 7360 1606
rect 7416 1604 7422 1606
rect 7114 1595 7422 1604
rect 7380 1556 7432 1562
rect 7380 1498 7432 1504
rect 7104 1420 7156 1426
rect 6932 1380 7104 1408
rect 7104 1362 7156 1368
rect 6736 1216 6788 1222
rect 6736 1158 6788 1164
rect 6748 1018 6776 1158
rect 6736 1012 6788 1018
rect 6736 954 6788 960
rect 7392 814 7420 1498
rect 7012 808 7064 814
rect 7012 750 7064 756
rect 7380 808 7432 814
rect 7380 750 7432 756
rect 6656 462 6776 490
rect 6748 400 6776 462
rect 1766 0 1822 400
rect 2318 0 2374 400
rect 2870 0 2926 400
rect 3422 0 3478 400
rect 3974 0 4030 400
rect 4526 0 4582 400
rect 5078 0 5134 400
rect 5630 0 5686 400
rect 6182 0 6238 400
rect 6734 0 6790 400
rect 7024 354 7052 750
rect 7114 572 7422 581
rect 7114 570 7120 572
rect 7176 570 7200 572
rect 7256 570 7280 572
rect 7336 570 7360 572
rect 7416 570 7422 572
rect 7176 518 7178 570
rect 7358 518 7360 570
rect 7114 516 7120 518
rect 7176 516 7200 518
rect 7256 516 7280 518
rect 7336 516 7360 518
rect 7416 516 7422 518
rect 7114 507 7422 516
rect 7208 428 7328 456
rect 7208 354 7236 428
rect 7300 400 7328 428
rect 7852 400 7880 1838
rect 7944 1562 7972 1838
rect 7932 1556 7984 1562
rect 7932 1498 7984 1504
rect 8312 1426 8340 2790
rect 8864 2650 8892 3334
rect 8852 2644 8904 2650
rect 8852 2586 8904 2592
rect 9048 2446 9076 4694
rect 9128 4480 9180 4486
rect 9128 4422 9180 4428
rect 9140 4282 9168 4422
rect 9128 4276 9180 4282
rect 9128 4218 9180 4224
rect 9128 4072 9180 4078
rect 9128 4014 9180 4020
rect 9140 3398 9168 4014
rect 9128 3392 9180 3398
rect 9128 3334 9180 3340
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 9140 2310 9168 3334
rect 9508 2446 9536 5782
rect 9692 5778 9720 5850
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 10152 5574 10180 6802
rect 9772 5568 9824 5574
rect 9772 5510 9824 5516
rect 10140 5568 10192 5574
rect 10140 5510 10192 5516
rect 9588 5024 9640 5030
rect 9588 4966 9640 4972
rect 9600 4758 9628 4966
rect 9784 4826 9812 5510
rect 10244 5166 10272 6802
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 10324 6724 10376 6730
rect 10324 6666 10376 6672
rect 10336 6458 10364 6666
rect 10472 6556 10780 6565
rect 10472 6554 10478 6556
rect 10534 6554 10558 6556
rect 10614 6554 10638 6556
rect 10694 6554 10718 6556
rect 10774 6554 10780 6556
rect 10534 6502 10536 6554
rect 10716 6502 10718 6554
rect 10472 6500 10478 6502
rect 10534 6500 10558 6502
rect 10614 6500 10638 6502
rect 10694 6500 10718 6502
rect 10774 6500 10780 6502
rect 10472 6491 10780 6500
rect 10324 6452 10376 6458
rect 10324 6394 10376 6400
rect 10336 6118 10364 6394
rect 11256 6254 11284 6734
rect 11244 6248 11296 6254
rect 11244 6190 11296 6196
rect 10324 6112 10376 6118
rect 10324 6054 10376 6060
rect 10336 5692 10364 6054
rect 10508 5704 10560 5710
rect 10336 5664 10508 5692
rect 10232 5160 10284 5166
rect 10232 5102 10284 5108
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 9588 4752 9640 4758
rect 9588 4694 9640 4700
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9692 4078 9720 4422
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 10336 4010 10364 5664
rect 10508 5646 10560 5652
rect 10472 5468 10780 5477
rect 10472 5466 10478 5468
rect 10534 5466 10558 5468
rect 10614 5466 10638 5468
rect 10694 5466 10718 5468
rect 10774 5466 10780 5468
rect 10534 5414 10536 5466
rect 10716 5414 10718 5466
rect 10472 5412 10478 5414
rect 10534 5412 10558 5414
rect 10614 5412 10638 5414
rect 10694 5412 10718 5414
rect 10774 5412 10780 5414
rect 10472 5403 10780 5412
rect 11256 5302 11284 6190
rect 11244 5296 11296 5302
rect 11244 5238 11296 5244
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 10796 4826 10824 5102
rect 11348 5030 11376 12406
rect 11532 12374 11560 13824
rect 11624 12714 11652 14214
rect 11716 12986 11744 14826
rect 11888 14612 11940 14618
rect 11888 14554 11940 14560
rect 11796 14272 11848 14278
rect 11796 14214 11848 14220
rect 11808 13462 11836 14214
rect 11900 13512 11928 14554
rect 11992 14550 12020 19110
rect 12176 19094 12296 19110
rect 12176 18834 12204 19094
rect 12360 18970 12388 19264
rect 12348 18964 12400 18970
rect 12348 18906 12400 18912
rect 12544 18834 12572 19858
rect 12820 19310 12848 21354
rect 13004 20058 13032 29446
rect 13188 28994 13216 29464
rect 13280 29306 13308 30330
rect 13464 29578 13492 31146
rect 13830 31036 14138 31045
rect 13830 31034 13836 31036
rect 13892 31034 13916 31036
rect 13972 31034 13996 31036
rect 14052 31034 14076 31036
rect 14132 31034 14138 31036
rect 13892 30982 13894 31034
rect 14074 30982 14076 31034
rect 13830 30980 13836 30982
rect 13892 30980 13916 30982
rect 13972 30980 13996 30982
rect 14052 30980 14076 30982
rect 14132 30980 14138 30982
rect 13830 30971 14138 30980
rect 14660 30802 14688 31600
rect 16132 30938 16160 31600
rect 16120 30932 16172 30938
rect 16120 30874 16172 30880
rect 17604 30870 17632 31600
rect 17592 30864 17644 30870
rect 17592 30806 17644 30812
rect 14648 30796 14700 30802
rect 14648 30738 14700 30744
rect 15292 30796 15344 30802
rect 15292 30738 15344 30744
rect 16764 30796 16816 30802
rect 16764 30738 16816 30744
rect 18052 30796 18104 30802
rect 18052 30738 18104 30744
rect 14096 30728 14148 30734
rect 14096 30670 14148 30676
rect 13636 30660 13688 30666
rect 13636 30602 13688 30608
rect 13544 30592 13596 30598
rect 13544 30534 13596 30540
rect 13556 30190 13584 30534
rect 13544 30184 13596 30190
rect 13544 30126 13596 30132
rect 13544 29640 13596 29646
rect 13544 29582 13596 29588
rect 13360 29572 13412 29578
rect 13360 29514 13412 29520
rect 13452 29572 13504 29578
rect 13452 29514 13504 29520
rect 13268 29300 13320 29306
rect 13268 29242 13320 29248
rect 13372 29170 13400 29514
rect 13360 29164 13412 29170
rect 13360 29106 13412 29112
rect 13188 28966 13308 28994
rect 13464 28966 13492 29514
rect 13556 29306 13584 29582
rect 13648 29510 13676 30602
rect 14108 30394 14136 30670
rect 14556 30660 14608 30666
rect 14556 30602 14608 30608
rect 14096 30388 14148 30394
rect 14096 30330 14148 30336
rect 14568 30190 14596 30602
rect 14648 30592 14700 30598
rect 14648 30534 14700 30540
rect 14660 30190 14688 30534
rect 14556 30184 14608 30190
rect 14556 30126 14608 30132
rect 14648 30184 14700 30190
rect 14648 30126 14700 30132
rect 13728 30116 13780 30122
rect 13728 30058 13780 30064
rect 14280 30116 14332 30122
rect 14280 30058 14332 30064
rect 13636 29504 13688 29510
rect 13636 29446 13688 29452
rect 13544 29300 13596 29306
rect 13544 29242 13596 29248
rect 13084 27940 13136 27946
rect 13084 27882 13136 27888
rect 13096 26518 13124 27882
rect 13084 26512 13136 26518
rect 13084 26454 13136 26460
rect 13176 25968 13228 25974
rect 13176 25910 13228 25916
rect 13188 25362 13216 25910
rect 13176 25356 13228 25362
rect 13176 25298 13228 25304
rect 13084 24608 13136 24614
rect 13084 24550 13136 24556
rect 13096 24410 13124 24550
rect 13084 24404 13136 24410
rect 13084 24346 13136 24352
rect 13084 24064 13136 24070
rect 13084 24006 13136 24012
rect 13176 24064 13228 24070
rect 13176 24006 13228 24012
rect 13096 23866 13124 24006
rect 13084 23860 13136 23866
rect 13084 23802 13136 23808
rect 13188 23730 13216 24006
rect 13176 23724 13228 23730
rect 13176 23666 13228 23672
rect 13176 22432 13228 22438
rect 13176 22374 13228 22380
rect 13084 20256 13136 20262
rect 13084 20198 13136 20204
rect 13096 20058 13124 20198
rect 12992 20052 13044 20058
rect 12992 19994 13044 20000
rect 13084 20052 13136 20058
rect 13084 19994 13136 20000
rect 12992 19916 13044 19922
rect 12992 19858 13044 19864
rect 13004 19825 13032 19858
rect 12990 19816 13046 19825
rect 12990 19751 13046 19760
rect 12624 19304 12676 19310
rect 12624 19246 12676 19252
rect 12808 19304 12860 19310
rect 12808 19246 12860 19252
rect 12164 18828 12216 18834
rect 12164 18770 12216 18776
rect 12440 18828 12492 18834
rect 12440 18770 12492 18776
rect 12532 18828 12584 18834
rect 12532 18770 12584 18776
rect 12452 18426 12480 18770
rect 12440 18420 12492 18426
rect 12440 18362 12492 18368
rect 12452 17066 12480 18362
rect 12636 17746 12664 19246
rect 12624 17740 12676 17746
rect 12624 17682 12676 17688
rect 12440 17060 12492 17066
rect 12440 17002 12492 17008
rect 12452 16658 12480 17002
rect 12440 16652 12492 16658
rect 12440 16594 12492 16600
rect 12624 16652 12676 16658
rect 12624 16594 12676 16600
rect 12452 15570 12480 16594
rect 12440 15564 12492 15570
rect 12440 15506 12492 15512
rect 12348 15360 12400 15366
rect 12348 15302 12400 15308
rect 12360 14958 12388 15302
rect 12636 15094 12664 16594
rect 12716 15564 12768 15570
rect 12716 15506 12768 15512
rect 12728 15094 12756 15506
rect 12624 15088 12676 15094
rect 12624 15030 12676 15036
rect 12716 15088 12768 15094
rect 12716 15030 12768 15036
rect 12348 14952 12400 14958
rect 12348 14894 12400 14900
rect 12072 14816 12124 14822
rect 12072 14758 12124 14764
rect 11980 14544 12032 14550
rect 11980 14486 12032 14492
rect 12084 14414 12112 14758
rect 12072 14408 12124 14414
rect 12072 14350 12124 14356
rect 12164 14408 12216 14414
rect 12164 14350 12216 14356
rect 12714 14376 12770 14385
rect 12176 14074 12204 14350
rect 12820 14362 12848 19246
rect 13188 17882 13216 22374
rect 13280 21078 13308 28966
rect 13452 28960 13504 28966
rect 13452 28902 13504 28908
rect 13544 28960 13596 28966
rect 13544 28902 13596 28908
rect 13464 28218 13492 28902
rect 13556 28422 13584 28902
rect 13544 28416 13596 28422
rect 13544 28358 13596 28364
rect 13452 28212 13504 28218
rect 13452 28154 13504 28160
rect 13556 28014 13584 28358
rect 13544 28008 13596 28014
rect 13544 27950 13596 27956
rect 13648 26926 13676 29446
rect 13740 29306 13768 30058
rect 13830 29948 14138 29957
rect 13830 29946 13836 29948
rect 13892 29946 13916 29948
rect 13972 29946 13996 29948
rect 14052 29946 14076 29948
rect 14132 29946 14138 29948
rect 13892 29894 13894 29946
rect 14074 29894 14076 29946
rect 13830 29892 13836 29894
rect 13892 29892 13916 29894
rect 13972 29892 13996 29894
rect 14052 29892 14076 29894
rect 14132 29892 14138 29894
rect 13830 29883 14138 29892
rect 14292 29850 14320 30058
rect 14660 30054 14688 30126
rect 15108 30116 15160 30122
rect 15108 30058 15160 30064
rect 14648 30048 14700 30054
rect 14648 29990 14700 29996
rect 14280 29844 14332 29850
rect 14280 29786 14332 29792
rect 15016 29844 15068 29850
rect 15016 29786 15068 29792
rect 14464 29776 14516 29782
rect 14464 29718 14516 29724
rect 14476 29578 14504 29718
rect 14464 29572 14516 29578
rect 14464 29514 14516 29520
rect 14648 29572 14700 29578
rect 14648 29514 14700 29520
rect 13728 29300 13780 29306
rect 13728 29242 13780 29248
rect 14464 29096 14516 29102
rect 14464 29038 14516 29044
rect 13830 28860 14138 28869
rect 13830 28858 13836 28860
rect 13892 28858 13916 28860
rect 13972 28858 13996 28860
rect 14052 28858 14076 28860
rect 14132 28858 14138 28860
rect 13892 28806 13894 28858
rect 14074 28806 14076 28858
rect 13830 28804 13836 28806
rect 13892 28804 13916 28806
rect 13972 28804 13996 28806
rect 14052 28804 14076 28806
rect 14132 28804 14138 28806
rect 13830 28795 14138 28804
rect 14280 28416 14332 28422
rect 14280 28358 14332 28364
rect 14292 28218 14320 28358
rect 14280 28212 14332 28218
rect 14280 28154 14332 28160
rect 13830 27772 14138 27781
rect 13830 27770 13836 27772
rect 13892 27770 13916 27772
rect 13972 27770 13996 27772
rect 14052 27770 14076 27772
rect 14132 27770 14138 27772
rect 13892 27718 13894 27770
rect 14074 27718 14076 27770
rect 13830 27716 13836 27718
rect 13892 27716 13916 27718
rect 13972 27716 13996 27718
rect 14052 27716 14076 27718
rect 14132 27716 14138 27718
rect 13830 27707 14138 27716
rect 14188 27396 14240 27402
rect 14188 27338 14240 27344
rect 14200 26994 14228 27338
rect 14188 26988 14240 26994
rect 14188 26930 14240 26936
rect 13636 26920 13688 26926
rect 13636 26862 13688 26868
rect 13544 26784 13596 26790
rect 13544 26726 13596 26732
rect 13556 26586 13584 26726
rect 13830 26684 14138 26693
rect 13830 26682 13836 26684
rect 13892 26682 13916 26684
rect 13972 26682 13996 26684
rect 14052 26682 14076 26684
rect 14132 26682 14138 26684
rect 13892 26630 13894 26682
rect 14074 26630 14076 26682
rect 13830 26628 13836 26630
rect 13892 26628 13916 26630
rect 13972 26628 13996 26630
rect 14052 26628 14076 26630
rect 14132 26628 14138 26630
rect 13830 26619 14138 26628
rect 13544 26580 13596 26586
rect 13544 26522 13596 26528
rect 13452 26444 13504 26450
rect 13452 26386 13504 26392
rect 14280 26444 14332 26450
rect 14280 26386 14332 26392
rect 13464 25158 13492 26386
rect 14188 26308 14240 26314
rect 14188 26250 14240 26256
rect 13728 26240 13780 26246
rect 13728 26182 13780 26188
rect 13820 26240 13872 26246
rect 13820 26182 13872 26188
rect 13740 25974 13768 26182
rect 13728 25968 13780 25974
rect 13728 25910 13780 25916
rect 13740 25838 13768 25910
rect 13636 25832 13688 25838
rect 13636 25774 13688 25780
rect 13728 25832 13780 25838
rect 13728 25774 13780 25780
rect 13544 25696 13596 25702
rect 13544 25638 13596 25644
rect 13556 25498 13584 25638
rect 13648 25498 13676 25774
rect 13832 25702 13860 26182
rect 14200 25838 14228 26250
rect 14188 25832 14240 25838
rect 14188 25774 14240 25780
rect 13820 25696 13872 25702
rect 13740 25656 13820 25684
rect 13544 25492 13596 25498
rect 13544 25434 13596 25440
rect 13636 25492 13688 25498
rect 13636 25434 13688 25440
rect 13740 25430 13768 25656
rect 13820 25638 13872 25644
rect 13830 25596 14138 25605
rect 13830 25594 13836 25596
rect 13892 25594 13916 25596
rect 13972 25594 13996 25596
rect 14052 25594 14076 25596
rect 14132 25594 14138 25596
rect 13892 25542 13894 25594
rect 14074 25542 14076 25594
rect 13830 25540 13836 25542
rect 13892 25540 13916 25542
rect 13972 25540 13996 25542
rect 14052 25540 14076 25542
rect 14132 25540 14138 25542
rect 13830 25531 14138 25540
rect 14200 25498 14228 25774
rect 14188 25492 14240 25498
rect 14188 25434 14240 25440
rect 13728 25424 13780 25430
rect 13728 25366 13780 25372
rect 14096 25356 14148 25362
rect 14096 25298 14148 25304
rect 13820 25220 13872 25226
rect 13820 25162 13872 25168
rect 13452 25152 13504 25158
rect 13452 25094 13504 25100
rect 13728 25152 13780 25158
rect 13728 25094 13780 25100
rect 13452 24812 13504 24818
rect 13452 24754 13504 24760
rect 13464 24070 13492 24754
rect 13740 24342 13768 25094
rect 13832 24818 13860 25162
rect 14004 25152 14056 25158
rect 14004 25094 14056 25100
rect 13820 24812 13872 24818
rect 13820 24754 13872 24760
rect 14016 24750 14044 25094
rect 14108 24954 14136 25298
rect 14096 24948 14148 24954
rect 14096 24890 14148 24896
rect 14292 24886 14320 26386
rect 14372 25832 14424 25838
rect 14372 25774 14424 25780
rect 14384 25294 14412 25774
rect 14372 25288 14424 25294
rect 14372 25230 14424 25236
rect 14476 24886 14504 29038
rect 14556 28688 14608 28694
rect 14556 28630 14608 28636
rect 14568 28014 14596 28630
rect 14556 28008 14608 28014
rect 14556 27950 14608 27956
rect 14568 27538 14596 27950
rect 14556 27532 14608 27538
rect 14556 27474 14608 27480
rect 14556 26240 14608 26246
rect 14556 26182 14608 26188
rect 14280 24880 14332 24886
rect 14280 24822 14332 24828
rect 14464 24880 14516 24886
rect 14464 24822 14516 24828
rect 14568 24818 14596 26182
rect 14660 25226 14688 29514
rect 15028 29170 15056 29786
rect 15016 29164 15068 29170
rect 15016 29106 15068 29112
rect 15120 29102 15148 30058
rect 15304 29850 15332 30738
rect 16396 30592 16448 30598
rect 16396 30534 16448 30540
rect 16408 30394 16436 30534
rect 15660 30388 15712 30394
rect 15660 30330 15712 30336
rect 16396 30388 16448 30394
rect 16396 30330 16448 30336
rect 15568 30116 15620 30122
rect 15568 30058 15620 30064
rect 15292 29844 15344 29850
rect 15292 29786 15344 29792
rect 15580 29782 15608 30058
rect 15384 29776 15436 29782
rect 15384 29718 15436 29724
rect 15568 29776 15620 29782
rect 15568 29718 15620 29724
rect 15108 29096 15160 29102
rect 15108 29038 15160 29044
rect 15016 28008 15068 28014
rect 15016 27950 15068 27956
rect 14832 27872 14884 27878
rect 14832 27814 14884 27820
rect 14844 27674 14872 27814
rect 14832 27668 14884 27674
rect 14832 27610 14884 27616
rect 15028 27402 15056 27950
rect 15120 27946 15148 29038
rect 15396 28762 15424 29718
rect 15568 29640 15620 29646
rect 15672 29628 15700 30330
rect 16408 30190 16436 30330
rect 16396 30184 16448 30190
rect 16396 30126 16448 30132
rect 16580 30116 16632 30122
rect 16580 30058 16632 30064
rect 16120 30048 16172 30054
rect 16120 29990 16172 29996
rect 16132 29850 16160 29990
rect 16120 29844 16172 29850
rect 16120 29786 16172 29792
rect 16212 29776 16264 29782
rect 16488 29776 16540 29782
rect 16264 29736 16488 29764
rect 16212 29718 16264 29724
rect 16488 29718 16540 29724
rect 15620 29600 15700 29628
rect 16592 29617 16620 30058
rect 16776 29850 16804 30738
rect 17776 30592 17828 30598
rect 17696 30552 17776 30580
rect 17188 30492 17496 30501
rect 17188 30490 17194 30492
rect 17250 30490 17274 30492
rect 17330 30490 17354 30492
rect 17410 30490 17434 30492
rect 17490 30490 17496 30492
rect 17250 30438 17252 30490
rect 17432 30438 17434 30490
rect 17188 30436 17194 30438
rect 17250 30436 17274 30438
rect 17330 30436 17354 30438
rect 17410 30436 17434 30438
rect 17490 30436 17496 30438
rect 17188 30427 17496 30436
rect 17040 30320 17092 30326
rect 17040 30262 17092 30268
rect 16948 30252 17000 30258
rect 16868 30212 16948 30240
rect 16764 29844 16816 29850
rect 16764 29786 16816 29792
rect 15568 29582 15620 29588
rect 15672 29510 15700 29600
rect 16578 29608 16634 29617
rect 16120 29572 16172 29578
rect 16578 29543 16634 29552
rect 16120 29514 16172 29520
rect 15660 29504 15712 29510
rect 15660 29446 15712 29452
rect 15936 29504 15988 29510
rect 15936 29446 15988 29452
rect 15568 28960 15620 28966
rect 15568 28902 15620 28908
rect 15384 28756 15436 28762
rect 15384 28698 15436 28704
rect 15292 28416 15344 28422
rect 15292 28358 15344 28364
rect 15304 28150 15332 28358
rect 15292 28144 15344 28150
rect 15292 28086 15344 28092
rect 15108 27940 15160 27946
rect 15108 27882 15160 27888
rect 15120 27538 15148 27882
rect 15108 27532 15160 27538
rect 15108 27474 15160 27480
rect 15016 27396 15068 27402
rect 15016 27338 15068 27344
rect 15200 27396 15252 27402
rect 15200 27338 15252 27344
rect 15212 27130 15240 27338
rect 15200 27124 15252 27130
rect 15200 27066 15252 27072
rect 15304 27062 15332 28086
rect 15580 27878 15608 28902
rect 15672 28626 15700 29446
rect 15752 29096 15804 29102
rect 15752 29038 15804 29044
rect 15660 28620 15712 28626
rect 15660 28562 15712 28568
rect 15764 28422 15792 29038
rect 15948 29034 15976 29446
rect 16132 29238 16160 29514
rect 16672 29504 16724 29510
rect 16672 29446 16724 29452
rect 16764 29504 16816 29510
rect 16764 29446 16816 29452
rect 16580 29300 16632 29306
rect 16580 29242 16632 29248
rect 16120 29232 16172 29238
rect 16120 29174 16172 29180
rect 15936 29028 15988 29034
rect 15936 28970 15988 28976
rect 15844 28960 15896 28966
rect 15844 28902 15896 28908
rect 15660 28416 15712 28422
rect 15660 28358 15712 28364
rect 15752 28416 15804 28422
rect 15752 28358 15804 28364
rect 15384 27872 15436 27878
rect 15384 27814 15436 27820
rect 15476 27872 15528 27878
rect 15476 27814 15528 27820
rect 15568 27872 15620 27878
rect 15568 27814 15620 27820
rect 15396 27334 15424 27814
rect 15488 27690 15516 27814
rect 15488 27662 15608 27690
rect 15580 27606 15608 27662
rect 15568 27600 15620 27606
rect 15568 27542 15620 27548
rect 15384 27328 15436 27334
rect 15384 27270 15436 27276
rect 15292 27056 15344 27062
rect 15292 26998 15344 27004
rect 15396 26790 15424 27270
rect 15580 26858 15608 27542
rect 15672 26926 15700 28358
rect 15856 28218 15884 28902
rect 15948 28762 15976 28970
rect 15936 28756 15988 28762
rect 15936 28698 15988 28704
rect 15936 28620 15988 28626
rect 15936 28562 15988 28568
rect 15844 28212 15896 28218
rect 15844 28154 15896 28160
rect 15948 27402 15976 28562
rect 16132 28422 16160 29174
rect 16396 28960 16448 28966
rect 16396 28902 16448 28908
rect 16408 28626 16436 28902
rect 16592 28642 16620 29242
rect 16684 29238 16712 29446
rect 16672 29232 16724 29238
rect 16672 29174 16724 29180
rect 16684 28694 16712 29174
rect 16776 28966 16804 29446
rect 16868 28994 16896 30212
rect 16948 30194 17000 30200
rect 17052 29850 17080 30262
rect 17316 30252 17368 30258
rect 17316 30194 17368 30200
rect 17040 29844 17092 29850
rect 17040 29786 17092 29792
rect 16948 29776 17000 29782
rect 16948 29718 17000 29724
rect 16960 29306 16988 29718
rect 17328 29714 17356 30194
rect 17316 29708 17368 29714
rect 17316 29650 17368 29656
rect 17040 29572 17092 29578
rect 17040 29514 17092 29520
rect 16948 29300 17000 29306
rect 16948 29242 17000 29248
rect 17052 29102 17080 29514
rect 17592 29504 17644 29510
rect 17592 29446 17644 29452
rect 17188 29404 17496 29413
rect 17188 29402 17194 29404
rect 17250 29402 17274 29404
rect 17330 29402 17354 29404
rect 17410 29402 17434 29404
rect 17490 29402 17496 29404
rect 17250 29350 17252 29402
rect 17432 29350 17434 29402
rect 17188 29348 17194 29350
rect 17250 29348 17274 29350
rect 17330 29348 17354 29350
rect 17410 29348 17434 29350
rect 17490 29348 17496 29350
rect 17188 29339 17496 29348
rect 17132 29300 17184 29306
rect 17132 29242 17184 29248
rect 17040 29096 17092 29102
rect 17040 29038 17092 29044
rect 16868 28966 17080 28994
rect 16764 28960 16816 28966
rect 16764 28902 16816 28908
rect 16396 28620 16448 28626
rect 16396 28562 16448 28568
rect 16500 28614 16620 28642
rect 16672 28688 16724 28694
rect 16672 28630 16724 28636
rect 16120 28416 16172 28422
rect 16120 28358 16172 28364
rect 16408 27878 16436 28562
rect 16396 27872 16448 27878
rect 16396 27814 16448 27820
rect 16408 27674 16436 27814
rect 16396 27668 16448 27674
rect 16396 27610 16448 27616
rect 15936 27396 15988 27402
rect 15936 27338 15988 27344
rect 16500 27334 16528 28614
rect 16580 28552 16632 28558
rect 16580 28494 16632 28500
rect 16592 28218 16620 28494
rect 16672 28484 16724 28490
rect 16672 28426 16724 28432
rect 16684 28218 16712 28426
rect 16764 28416 16816 28422
rect 16764 28358 16816 28364
rect 16580 28212 16632 28218
rect 16580 28154 16632 28160
rect 16672 28212 16724 28218
rect 16672 28154 16724 28160
rect 16592 27334 16620 28154
rect 16672 27872 16724 27878
rect 16670 27840 16672 27849
rect 16724 27840 16726 27849
rect 16776 27826 16804 28358
rect 16948 28076 17000 28082
rect 16948 28018 17000 28024
rect 16960 27860 16988 28018
rect 16868 27832 16988 27860
rect 16776 27798 16820 27826
rect 16670 27775 16726 27784
rect 16672 27668 16724 27674
rect 16672 27610 16724 27616
rect 16792 27614 16820 27798
rect 15844 27328 15896 27334
rect 15844 27270 15896 27276
rect 16488 27328 16540 27334
rect 16488 27270 16540 27276
rect 16580 27328 16632 27334
rect 16580 27270 16632 27276
rect 15660 26920 15712 26926
rect 15660 26862 15712 26868
rect 15568 26852 15620 26858
rect 15568 26794 15620 26800
rect 15384 26784 15436 26790
rect 15384 26726 15436 26732
rect 15660 26784 15712 26790
rect 15660 26726 15712 26732
rect 15752 26784 15804 26790
rect 15752 26726 15804 26732
rect 15672 26518 15700 26726
rect 15764 26586 15792 26726
rect 15856 26586 15884 27270
rect 16500 27146 16528 27270
rect 16500 27118 16620 27146
rect 15752 26580 15804 26586
rect 15752 26522 15804 26528
rect 15844 26580 15896 26586
rect 15844 26522 15896 26528
rect 15660 26512 15712 26518
rect 15660 26454 15712 26460
rect 15568 26444 15620 26450
rect 15568 26386 15620 26392
rect 15292 26308 15344 26314
rect 15292 26250 15344 26256
rect 15200 25696 15252 25702
rect 15200 25638 15252 25644
rect 14832 25492 14884 25498
rect 14832 25434 14884 25440
rect 14648 25220 14700 25226
rect 14648 25162 14700 25168
rect 14844 25158 14872 25434
rect 14924 25424 14976 25430
rect 14924 25366 14976 25372
rect 14832 25152 14884 25158
rect 14832 25094 14884 25100
rect 14936 24954 14964 25366
rect 15212 25242 15240 25638
rect 15016 25220 15068 25226
rect 15016 25162 15068 25168
rect 15120 25214 15240 25242
rect 15028 24954 15056 25162
rect 14924 24948 14976 24954
rect 14924 24890 14976 24896
rect 15016 24948 15068 24954
rect 15016 24890 15068 24896
rect 14832 24880 14884 24886
rect 14832 24822 14884 24828
rect 14188 24812 14240 24818
rect 14188 24754 14240 24760
rect 14556 24812 14608 24818
rect 14556 24754 14608 24760
rect 14004 24744 14056 24750
rect 14004 24686 14056 24692
rect 13830 24508 14138 24517
rect 13830 24506 13836 24508
rect 13892 24506 13916 24508
rect 13972 24506 13996 24508
rect 14052 24506 14076 24508
rect 14132 24506 14138 24508
rect 13892 24454 13894 24506
rect 14074 24454 14076 24506
rect 13830 24452 13836 24454
rect 13892 24452 13916 24454
rect 13972 24452 13996 24454
rect 14052 24452 14076 24454
rect 14132 24452 14138 24454
rect 13830 24443 14138 24452
rect 13728 24336 13780 24342
rect 13728 24278 13780 24284
rect 13820 24268 13872 24274
rect 13820 24210 13872 24216
rect 13452 24064 13504 24070
rect 13452 24006 13504 24012
rect 13464 22506 13492 24006
rect 13832 23798 13860 24210
rect 14200 24070 14228 24754
rect 14844 24732 14872 24822
rect 15120 24818 15148 25214
rect 15200 25152 15252 25158
rect 15200 25094 15252 25100
rect 15212 24818 15240 25094
rect 15108 24812 15160 24818
rect 15108 24754 15160 24760
rect 15200 24812 15252 24818
rect 15200 24754 15252 24760
rect 14844 24704 14964 24732
rect 14464 24676 14516 24682
rect 14464 24618 14516 24624
rect 14280 24200 14332 24206
rect 14280 24142 14332 24148
rect 14188 24064 14240 24070
rect 14188 24006 14240 24012
rect 13820 23792 13872 23798
rect 13820 23734 13872 23740
rect 13544 23520 13596 23526
rect 13832 23508 13860 23734
rect 13544 23462 13596 23468
rect 13740 23480 13860 23508
rect 13556 23186 13584 23462
rect 13544 23180 13596 23186
rect 13544 23122 13596 23128
rect 13740 22778 13768 23480
rect 13830 23420 14138 23429
rect 13830 23418 13836 23420
rect 13892 23418 13916 23420
rect 13972 23418 13996 23420
rect 14052 23418 14076 23420
rect 14132 23418 14138 23420
rect 13892 23366 13894 23418
rect 14074 23366 14076 23418
rect 13830 23364 13836 23366
rect 13892 23364 13916 23366
rect 13972 23364 13996 23366
rect 14052 23364 14076 23366
rect 14132 23364 14138 23366
rect 13830 23355 14138 23364
rect 14292 23186 14320 24142
rect 14476 24138 14504 24618
rect 14740 24608 14792 24614
rect 14740 24550 14792 24556
rect 14752 24206 14780 24550
rect 14740 24200 14792 24206
rect 14740 24142 14792 24148
rect 14464 24132 14516 24138
rect 14464 24074 14516 24080
rect 14476 23866 14504 24074
rect 14464 23860 14516 23866
rect 14464 23802 14516 23808
rect 14752 23798 14780 24142
rect 14740 23792 14792 23798
rect 14660 23752 14740 23780
rect 14280 23180 14332 23186
rect 14280 23122 14332 23128
rect 13820 23044 13872 23050
rect 13820 22986 13872 22992
rect 13728 22772 13780 22778
rect 13728 22714 13780 22720
rect 13832 22574 13860 22986
rect 14280 22704 14332 22710
rect 14280 22646 14332 22652
rect 13820 22568 13872 22574
rect 13740 22516 13820 22522
rect 13740 22510 13872 22516
rect 13452 22500 13504 22506
rect 13452 22442 13504 22448
rect 13740 22494 13860 22510
rect 13636 22432 13688 22438
rect 13636 22374 13688 22380
rect 13648 21690 13676 22374
rect 13740 22114 13768 22494
rect 13830 22332 14138 22341
rect 13830 22330 13836 22332
rect 13892 22330 13916 22332
rect 13972 22330 13996 22332
rect 14052 22330 14076 22332
rect 14132 22330 14138 22332
rect 13892 22278 13894 22330
rect 14074 22278 14076 22330
rect 13830 22276 13836 22278
rect 13892 22276 13916 22278
rect 13972 22276 13996 22278
rect 14052 22276 14076 22278
rect 14132 22276 14138 22278
rect 13830 22267 14138 22276
rect 13740 22086 13860 22114
rect 13832 21894 13860 22086
rect 14188 22092 14240 22098
rect 14188 22034 14240 22040
rect 13820 21888 13872 21894
rect 13820 21830 13872 21836
rect 13636 21684 13688 21690
rect 13636 21626 13688 21632
rect 13832 21486 13860 21830
rect 14200 21690 14228 22034
rect 14292 21842 14320 22646
rect 14660 22574 14688 23752
rect 14740 23734 14792 23740
rect 14740 23520 14792 23526
rect 14740 23462 14792 23468
rect 14752 23322 14780 23462
rect 14740 23316 14792 23322
rect 14740 23258 14792 23264
rect 14648 22568 14700 22574
rect 14648 22510 14700 22516
rect 14556 22500 14608 22506
rect 14556 22442 14608 22448
rect 14292 21814 14412 21842
rect 14188 21684 14240 21690
rect 14188 21626 14240 21632
rect 14384 21486 14412 21814
rect 13820 21480 13872 21486
rect 13820 21422 13872 21428
rect 14372 21480 14424 21486
rect 14372 21422 14424 21428
rect 14188 21412 14240 21418
rect 14188 21354 14240 21360
rect 13830 21244 14138 21253
rect 13830 21242 13836 21244
rect 13892 21242 13916 21244
rect 13972 21242 13996 21244
rect 14052 21242 14076 21244
rect 14132 21242 14138 21244
rect 13892 21190 13894 21242
rect 14074 21190 14076 21242
rect 13830 21188 13836 21190
rect 13892 21188 13916 21190
rect 13972 21188 13996 21190
rect 14052 21188 14076 21190
rect 14132 21188 14138 21190
rect 13830 21179 14138 21188
rect 13268 21072 13320 21078
rect 13268 21014 13320 21020
rect 13280 20466 13308 21014
rect 13636 20936 13688 20942
rect 13636 20878 13688 20884
rect 13268 20460 13320 20466
rect 13268 20402 13320 20408
rect 13648 20398 13676 20878
rect 14096 20800 14148 20806
rect 14096 20742 14148 20748
rect 14108 20398 14136 20742
rect 14200 20602 14228 21354
rect 14280 21344 14332 21350
rect 14280 21286 14332 21292
rect 14372 21344 14424 21350
rect 14372 21286 14424 21292
rect 14292 21146 14320 21286
rect 14280 21140 14332 21146
rect 14280 21082 14332 21088
rect 14188 20596 14240 20602
rect 14188 20538 14240 20544
rect 14384 20466 14412 21286
rect 14464 20528 14516 20534
rect 14464 20470 14516 20476
rect 14188 20460 14240 20466
rect 14188 20402 14240 20408
rect 14372 20460 14424 20466
rect 14372 20402 14424 20408
rect 13636 20392 13688 20398
rect 13636 20334 13688 20340
rect 14096 20392 14148 20398
rect 14096 20334 14148 20340
rect 13648 19922 13676 20334
rect 13830 20156 14138 20165
rect 13830 20154 13836 20156
rect 13892 20154 13916 20156
rect 13972 20154 13996 20156
rect 14052 20154 14076 20156
rect 14132 20154 14138 20156
rect 13892 20102 13894 20154
rect 14074 20102 14076 20154
rect 13830 20100 13836 20102
rect 13892 20100 13916 20102
rect 13972 20100 13996 20102
rect 14052 20100 14076 20102
rect 14132 20100 14138 20102
rect 13830 20091 14138 20100
rect 14200 20058 14228 20402
rect 14188 20052 14240 20058
rect 14188 19994 14240 20000
rect 14200 19922 14228 19994
rect 13636 19916 13688 19922
rect 13636 19858 13688 19864
rect 14188 19916 14240 19922
rect 14188 19858 14240 19864
rect 14096 19780 14148 19786
rect 14096 19722 14148 19728
rect 14108 19514 14136 19722
rect 13452 19508 13504 19514
rect 13452 19450 13504 19456
rect 14096 19508 14148 19514
rect 14096 19450 14148 19456
rect 13268 18216 13320 18222
rect 13268 18158 13320 18164
rect 13176 17876 13228 17882
rect 13176 17818 13228 17824
rect 13280 17746 13308 18158
rect 13464 17746 13492 19450
rect 13544 19304 13596 19310
rect 13544 19246 13596 19252
rect 13556 19174 13584 19246
rect 13544 19168 13596 19174
rect 13544 19110 13596 19116
rect 13728 19168 13780 19174
rect 13728 19110 13780 19116
rect 14280 19168 14332 19174
rect 14280 19110 14332 19116
rect 13740 18970 13768 19110
rect 13830 19068 14138 19077
rect 13830 19066 13836 19068
rect 13892 19066 13916 19068
rect 13972 19066 13996 19068
rect 14052 19066 14076 19068
rect 14132 19066 14138 19068
rect 13892 19014 13894 19066
rect 14074 19014 14076 19066
rect 13830 19012 13836 19014
rect 13892 19012 13916 19014
rect 13972 19012 13996 19014
rect 14052 19012 14076 19014
rect 14132 19012 14138 19014
rect 13830 19003 14138 19012
rect 14292 18970 14320 19110
rect 13728 18964 13780 18970
rect 13728 18906 13780 18912
rect 14280 18964 14332 18970
rect 14280 18906 14332 18912
rect 13740 17746 13768 18906
rect 14280 18624 14332 18630
rect 14280 18566 14332 18572
rect 14188 18148 14240 18154
rect 14188 18090 14240 18096
rect 13830 17980 14138 17989
rect 13830 17978 13836 17980
rect 13892 17978 13916 17980
rect 13972 17978 13996 17980
rect 14052 17978 14076 17980
rect 14132 17978 14138 17980
rect 13892 17926 13894 17978
rect 14074 17926 14076 17978
rect 13830 17924 13836 17926
rect 13892 17924 13916 17926
rect 13972 17924 13996 17926
rect 14052 17924 14076 17926
rect 14132 17924 14138 17926
rect 13830 17915 14138 17924
rect 14004 17808 14056 17814
rect 14004 17750 14056 17756
rect 13268 17740 13320 17746
rect 13268 17682 13320 17688
rect 13452 17740 13504 17746
rect 13452 17682 13504 17688
rect 13728 17740 13780 17746
rect 13728 17682 13780 17688
rect 13820 17740 13872 17746
rect 13820 17682 13872 17688
rect 13084 16788 13136 16794
rect 13084 16730 13136 16736
rect 12900 16176 12952 16182
rect 12900 16118 12952 16124
rect 12770 14334 12848 14362
rect 12714 14311 12770 14320
rect 12624 14272 12676 14278
rect 12624 14214 12676 14220
rect 12164 14068 12216 14074
rect 12164 14010 12216 14016
rect 12256 13796 12308 13802
rect 12256 13738 12308 13744
rect 12268 13530 12296 13738
rect 12636 13530 12664 14214
rect 12716 13864 12768 13870
rect 12716 13806 12768 13812
rect 12728 13734 12756 13806
rect 12716 13728 12768 13734
rect 12716 13670 12768 13676
rect 12256 13524 12308 13530
rect 11900 13484 12020 13512
rect 11796 13456 11848 13462
rect 11796 13398 11848 13404
rect 11888 13388 11940 13394
rect 11888 13330 11940 13336
rect 11900 12986 11928 13330
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 11992 12782 12020 13484
rect 12256 13466 12308 13472
rect 12624 13524 12676 13530
rect 12624 13466 12676 13472
rect 12072 12912 12124 12918
rect 12072 12854 12124 12860
rect 11980 12776 12032 12782
rect 11980 12718 12032 12724
rect 11612 12708 11664 12714
rect 11612 12650 11664 12656
rect 11980 12640 12032 12646
rect 11980 12582 12032 12588
rect 11992 12442 12020 12582
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 11520 12368 11572 12374
rect 11520 12310 11572 12316
rect 11532 6254 11560 12310
rect 11888 12300 11940 12306
rect 11888 12242 11940 12248
rect 11612 11552 11664 11558
rect 11612 11494 11664 11500
rect 11624 11286 11652 11494
rect 11612 11280 11664 11286
rect 11612 11222 11664 11228
rect 11900 11218 11928 12242
rect 12084 11694 12112 12854
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12348 12640 12400 12646
rect 12348 12582 12400 12588
rect 12360 11762 12388 12582
rect 12452 11898 12480 12718
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 12544 12102 12572 12582
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12348 11756 12400 11762
rect 12348 11698 12400 11704
rect 12072 11688 12124 11694
rect 12072 11630 12124 11636
rect 11888 11212 11940 11218
rect 11888 11154 11940 11160
rect 12164 10600 12216 10606
rect 12164 10542 12216 10548
rect 11980 10464 12032 10470
rect 11980 10406 12032 10412
rect 11888 7948 11940 7954
rect 11888 7890 11940 7896
rect 11704 7744 11756 7750
rect 11704 7686 11756 7692
rect 11716 7546 11744 7686
rect 11704 7540 11756 7546
rect 11704 7482 11756 7488
rect 11900 7177 11928 7890
rect 11886 7168 11942 7177
rect 11886 7103 11942 7112
rect 11900 7002 11928 7103
rect 11888 6996 11940 7002
rect 11888 6938 11940 6944
rect 11796 6860 11848 6866
rect 11796 6802 11848 6808
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11716 6458 11744 6598
rect 11704 6452 11756 6458
rect 11704 6394 11756 6400
rect 11808 6254 11836 6802
rect 11520 6248 11572 6254
rect 11520 6190 11572 6196
rect 11796 6248 11848 6254
rect 11796 6190 11848 6196
rect 11888 6248 11940 6254
rect 11888 6190 11940 6196
rect 11520 6112 11572 6118
rect 11520 6054 11572 6060
rect 11612 6112 11664 6118
rect 11612 6054 11664 6060
rect 11532 5574 11560 6054
rect 11624 5846 11652 6054
rect 11612 5840 11664 5846
rect 11612 5782 11664 5788
rect 11796 5772 11848 5778
rect 11796 5714 11848 5720
rect 11520 5568 11572 5574
rect 11520 5510 11572 5516
rect 11532 5098 11560 5510
rect 11520 5092 11572 5098
rect 11520 5034 11572 5040
rect 11336 5024 11388 5030
rect 11336 4966 11388 4972
rect 10784 4820 10836 4826
rect 10784 4762 10836 4768
rect 10692 4752 10744 4758
rect 10744 4700 10916 4706
rect 10692 4694 10916 4700
rect 10704 4678 10916 4694
rect 11808 4690 11836 5714
rect 11900 5370 11928 6190
rect 11992 5778 12020 10406
rect 12176 9586 12204 10542
rect 12728 9674 12756 13670
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 12820 12986 12848 13330
rect 12808 12980 12860 12986
rect 12808 12922 12860 12928
rect 12912 12646 12940 16118
rect 12992 15564 13044 15570
rect 12992 15506 13044 15512
rect 13004 15162 13032 15506
rect 12992 15156 13044 15162
rect 12992 15098 13044 15104
rect 13096 14958 13124 16730
rect 13464 16046 13492 17682
rect 13636 17672 13688 17678
rect 13636 17614 13688 17620
rect 13544 17060 13596 17066
rect 13544 17002 13596 17008
rect 13452 16040 13504 16046
rect 13452 15982 13504 15988
rect 13556 15638 13584 17002
rect 13544 15632 13596 15638
rect 13544 15574 13596 15580
rect 13452 15360 13504 15366
rect 13452 15302 13504 15308
rect 13464 14958 13492 15302
rect 13084 14952 13136 14958
rect 13084 14894 13136 14900
rect 13176 14952 13228 14958
rect 13176 14894 13228 14900
rect 13452 14952 13504 14958
rect 13452 14894 13504 14900
rect 13096 13938 13124 14894
rect 13084 13932 13136 13938
rect 13084 13874 13136 13880
rect 13096 13734 13124 13874
rect 13084 13728 13136 13734
rect 13084 13670 13136 13676
rect 13096 12850 13124 13670
rect 13084 12844 13136 12850
rect 13084 12786 13136 12792
rect 12900 12640 12952 12646
rect 12900 12582 12952 12588
rect 12912 11694 12940 12582
rect 12900 11688 12952 11694
rect 12900 11630 12952 11636
rect 12992 11552 13044 11558
rect 12992 11494 13044 11500
rect 13004 11354 13032 11494
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 12992 11008 13044 11014
rect 12992 10950 13044 10956
rect 13004 10606 13032 10950
rect 13084 10736 13136 10742
rect 13084 10678 13136 10684
rect 12992 10600 13044 10606
rect 12992 10542 13044 10548
rect 12900 10464 12952 10470
rect 12900 10406 12952 10412
rect 12544 9646 12756 9674
rect 12808 9648 12860 9654
rect 12164 9580 12216 9586
rect 12164 9522 12216 9528
rect 12348 9512 12400 9518
rect 12544 9500 12572 9646
rect 12808 9590 12860 9596
rect 12624 9512 12676 9518
rect 12544 9472 12624 9500
rect 12348 9454 12400 9460
rect 12624 9454 12676 9460
rect 12360 8430 12388 9454
rect 12532 9376 12584 9382
rect 12532 9318 12584 9324
rect 12440 8968 12492 8974
rect 12440 8910 12492 8916
rect 12348 8424 12400 8430
rect 12348 8366 12400 8372
rect 12360 7954 12388 8366
rect 12452 8022 12480 8910
rect 12544 8498 12572 9318
rect 12820 9178 12848 9590
rect 12912 9178 12940 10406
rect 13004 10130 13032 10542
rect 13096 10470 13124 10678
rect 13084 10464 13136 10470
rect 13084 10406 13136 10412
rect 13096 10130 13124 10406
rect 12992 10124 13044 10130
rect 12992 10066 13044 10072
rect 13084 10124 13136 10130
rect 13084 10066 13136 10072
rect 13004 9450 13032 10066
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 12992 9444 13044 9450
rect 12992 9386 13044 9392
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 12912 8566 12940 9114
rect 12900 8560 12952 8566
rect 12900 8502 12952 8508
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12624 8492 12676 8498
rect 12624 8434 12676 8440
rect 12544 8090 12572 8434
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12440 8016 12492 8022
rect 12440 7958 12492 7964
rect 12348 7948 12400 7954
rect 12348 7890 12400 7896
rect 12532 7948 12584 7954
rect 12636 7936 12664 8434
rect 12808 8356 12860 8362
rect 12808 8298 12860 8304
rect 12584 7908 12664 7936
rect 12532 7890 12584 7896
rect 12164 7880 12216 7886
rect 12164 7822 12216 7828
rect 12176 7002 12204 7822
rect 12348 7744 12400 7750
rect 12348 7686 12400 7692
rect 12164 6996 12216 7002
rect 12164 6938 12216 6944
rect 12072 6656 12124 6662
rect 12072 6598 12124 6604
rect 12084 6458 12112 6598
rect 12072 6452 12124 6458
rect 12072 6394 12124 6400
rect 12360 5778 12388 7686
rect 12624 7404 12676 7410
rect 12624 7346 12676 7352
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 12452 6730 12480 7278
rect 12532 6860 12584 6866
rect 12532 6802 12584 6808
rect 12440 6724 12492 6730
rect 12440 6666 12492 6672
rect 12544 6322 12572 6802
rect 12636 6322 12664 7346
rect 12716 6860 12768 6866
rect 12716 6802 12768 6808
rect 12728 6730 12756 6802
rect 12716 6724 12768 6730
rect 12716 6666 12768 6672
rect 12532 6316 12584 6322
rect 12532 6258 12584 6264
rect 12624 6316 12676 6322
rect 12624 6258 12676 6264
rect 12728 6186 12756 6666
rect 12716 6180 12768 6186
rect 12716 6122 12768 6128
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 12256 5772 12308 5778
rect 12256 5714 12308 5720
rect 12348 5772 12400 5778
rect 12348 5714 12400 5720
rect 12532 5772 12584 5778
rect 12532 5714 12584 5720
rect 12072 5568 12124 5574
rect 12072 5510 12124 5516
rect 11888 5364 11940 5370
rect 11888 5306 11940 5312
rect 11980 5364 12032 5370
rect 11980 5306 12032 5312
rect 11992 5250 12020 5306
rect 11900 5222 12020 5250
rect 11900 5030 11928 5222
rect 12084 5166 12112 5510
rect 12072 5160 12124 5166
rect 12072 5102 12124 5108
rect 12164 5092 12216 5098
rect 12164 5034 12216 5040
rect 11888 5024 11940 5030
rect 11888 4966 11940 4972
rect 12072 5024 12124 5030
rect 12072 4966 12124 4972
rect 12084 4758 12112 4966
rect 12072 4752 12124 4758
rect 12072 4694 12124 4700
rect 10472 4380 10780 4389
rect 10472 4378 10478 4380
rect 10534 4378 10558 4380
rect 10614 4378 10638 4380
rect 10694 4378 10718 4380
rect 10774 4378 10780 4380
rect 10534 4326 10536 4378
rect 10716 4326 10718 4378
rect 10472 4324 10478 4326
rect 10534 4324 10558 4326
rect 10614 4324 10638 4326
rect 10694 4324 10718 4326
rect 10774 4324 10780 4326
rect 10472 4315 10780 4324
rect 10888 4214 10916 4678
rect 11244 4684 11296 4690
rect 11244 4626 11296 4632
rect 11796 4684 11848 4690
rect 11796 4626 11848 4632
rect 10968 4480 11020 4486
rect 10968 4422 11020 4428
rect 10876 4208 10928 4214
rect 10876 4150 10928 4156
rect 10980 4146 11008 4422
rect 10968 4140 11020 4146
rect 10968 4082 11020 4088
rect 10600 4072 10652 4078
rect 10600 4014 10652 4020
rect 9956 4004 10008 4010
rect 9956 3946 10008 3952
rect 10324 4004 10376 4010
rect 10324 3946 10376 3952
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 9680 2916 9732 2922
rect 9680 2858 9732 2864
rect 9692 2650 9720 2858
rect 9680 2644 9732 2650
rect 9680 2586 9732 2592
rect 9496 2440 9548 2446
rect 9496 2382 9548 2388
rect 9128 2304 9180 2310
rect 9128 2246 9180 2252
rect 9220 1896 9272 1902
rect 9220 1838 9272 1844
rect 8944 1488 8996 1494
rect 8944 1430 8996 1436
rect 8300 1420 8352 1426
rect 8300 1362 8352 1368
rect 8024 1352 8076 1358
rect 8024 1294 8076 1300
rect 8036 1018 8064 1294
rect 8024 1012 8076 1018
rect 8024 954 8076 960
rect 8300 808 8352 814
rect 8352 768 8432 796
rect 8300 750 8352 756
rect 8404 400 8432 768
rect 8956 400 8984 1430
rect 9232 882 9260 1838
rect 9312 1420 9364 1426
rect 9364 1380 9536 1408
rect 9312 1362 9364 1368
rect 9220 876 9272 882
rect 9220 818 9272 824
rect 9508 400 9536 1380
rect 9680 808 9732 814
rect 9784 796 9812 3674
rect 9968 3058 9996 3946
rect 10612 3602 10640 4014
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 10796 3641 10824 3674
rect 10782 3632 10838 3641
rect 10232 3596 10284 3602
rect 10232 3538 10284 3544
rect 10600 3596 10652 3602
rect 10782 3567 10838 3576
rect 10600 3538 10652 3544
rect 10244 3194 10272 3538
rect 10472 3292 10780 3301
rect 10472 3290 10478 3292
rect 10534 3290 10558 3292
rect 10614 3290 10638 3292
rect 10694 3290 10718 3292
rect 10774 3290 10780 3292
rect 10534 3238 10536 3290
rect 10716 3238 10718 3290
rect 10472 3236 10478 3238
rect 10534 3236 10558 3238
rect 10614 3236 10638 3238
rect 10694 3236 10718 3238
rect 10774 3236 10780 3238
rect 10472 3227 10780 3236
rect 10232 3188 10284 3194
rect 10232 3130 10284 3136
rect 10692 3120 10744 3126
rect 10744 3080 10916 3108
rect 10692 3062 10744 3068
rect 9956 3052 10008 3058
rect 9956 2994 10008 3000
rect 10784 2984 10836 2990
rect 10784 2926 10836 2932
rect 10048 2848 10100 2854
rect 10048 2790 10100 2796
rect 9864 1420 9916 1426
rect 10060 1408 10088 2790
rect 10796 2650 10824 2926
rect 10784 2644 10836 2650
rect 10784 2586 10836 2592
rect 10140 2372 10192 2378
rect 10140 2314 10192 2320
rect 10152 1902 10180 2314
rect 10324 2304 10376 2310
rect 10324 2246 10376 2252
rect 10336 2106 10364 2246
rect 10472 2204 10780 2213
rect 10472 2202 10478 2204
rect 10534 2202 10558 2204
rect 10614 2202 10638 2204
rect 10694 2202 10718 2204
rect 10774 2202 10780 2204
rect 10534 2150 10536 2202
rect 10716 2150 10718 2202
rect 10472 2148 10478 2150
rect 10534 2148 10558 2150
rect 10614 2148 10638 2150
rect 10694 2148 10718 2150
rect 10774 2148 10780 2150
rect 10472 2139 10780 2148
rect 10324 2100 10376 2106
rect 10324 2042 10376 2048
rect 10140 1896 10192 1902
rect 10140 1838 10192 1844
rect 10784 1896 10836 1902
rect 10888 1884 10916 3080
rect 11072 2990 11100 3878
rect 11256 2990 11284 4626
rect 11808 4078 11836 4626
rect 12072 4616 12124 4622
rect 12176 4604 12204 5034
rect 12268 4826 12296 5714
rect 12256 4820 12308 4826
rect 12256 4762 12308 4768
rect 12124 4576 12204 4604
rect 12072 4558 12124 4564
rect 12084 4078 12112 4558
rect 11796 4072 11848 4078
rect 11796 4014 11848 4020
rect 12072 4072 12124 4078
rect 12072 4014 12124 4020
rect 11336 3528 11388 3534
rect 11336 3470 11388 3476
rect 11060 2984 11112 2990
rect 11060 2926 11112 2932
rect 11244 2984 11296 2990
rect 11244 2926 11296 2932
rect 11348 2922 11376 3470
rect 11808 3466 11836 4014
rect 12084 3738 12112 4014
rect 12072 3732 12124 3738
rect 12072 3674 12124 3680
rect 11796 3460 11848 3466
rect 11796 3402 11848 3408
rect 11428 3392 11480 3398
rect 11428 3334 11480 3340
rect 12256 3392 12308 3398
rect 12256 3334 12308 3340
rect 11336 2916 11388 2922
rect 11336 2858 11388 2864
rect 10968 2848 11020 2854
rect 10968 2790 11020 2796
rect 10980 2378 11008 2790
rect 11348 2650 11376 2858
rect 11336 2644 11388 2650
rect 11336 2586 11388 2592
rect 11440 2514 11468 3334
rect 11888 3188 11940 3194
rect 11888 3130 11940 3136
rect 11900 2514 11928 3130
rect 12268 2774 12296 3334
rect 12360 2990 12388 5714
rect 12544 4690 12572 5714
rect 12716 5568 12768 5574
rect 12716 5510 12768 5516
rect 12728 5166 12756 5510
rect 12716 5160 12768 5166
rect 12716 5102 12768 5108
rect 12532 4684 12584 4690
rect 12532 4626 12584 4632
rect 12820 4622 12848 8298
rect 12900 7880 12952 7886
rect 12900 7822 12952 7828
rect 12912 7546 12940 7822
rect 12900 7540 12952 7546
rect 12900 7482 12952 7488
rect 12992 7336 13044 7342
rect 12992 7278 13044 7284
rect 13004 7177 13032 7278
rect 12990 7168 13046 7177
rect 12990 7103 13046 7112
rect 12900 6928 12952 6934
rect 12900 6870 12952 6876
rect 12912 6458 12940 6870
rect 12900 6452 12952 6458
rect 12900 6394 12952 6400
rect 12900 5772 12952 5778
rect 12900 5714 12952 5720
rect 12912 5370 12940 5714
rect 12992 5704 13044 5710
rect 12992 5646 13044 5652
rect 13004 5370 13032 5646
rect 12900 5364 12952 5370
rect 12900 5306 12952 5312
rect 12992 5364 13044 5370
rect 12992 5306 13044 5312
rect 13096 5166 13124 9862
rect 13188 9518 13216 14894
rect 13556 14822 13584 15574
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 13556 13818 13584 14758
rect 13648 14618 13676 17614
rect 13740 16454 13768 17682
rect 13832 17066 13860 17682
rect 13912 17536 13964 17542
rect 13912 17478 13964 17484
rect 13924 17202 13952 17478
rect 14016 17202 14044 17750
rect 14200 17338 14228 18090
rect 14188 17332 14240 17338
rect 14188 17274 14240 17280
rect 13912 17196 13964 17202
rect 13912 17138 13964 17144
rect 14004 17196 14056 17202
rect 14004 17138 14056 17144
rect 14292 17134 14320 18566
rect 14384 17882 14412 20402
rect 14372 17876 14424 17882
rect 14372 17818 14424 17824
rect 14280 17128 14332 17134
rect 14280 17070 14332 17076
rect 13820 17060 13872 17066
rect 13820 17002 13872 17008
rect 13830 16892 14138 16901
rect 13830 16890 13836 16892
rect 13892 16890 13916 16892
rect 13972 16890 13996 16892
rect 14052 16890 14076 16892
rect 14132 16890 14138 16892
rect 13892 16838 13894 16890
rect 14074 16838 14076 16890
rect 13830 16836 13836 16838
rect 13892 16836 13916 16838
rect 13972 16836 13996 16838
rect 14052 16836 14076 16838
rect 14132 16836 14138 16838
rect 13830 16827 14138 16836
rect 14096 16652 14148 16658
rect 14096 16594 14148 16600
rect 13728 16448 13780 16454
rect 13728 16390 13780 16396
rect 14108 16250 14136 16594
rect 14096 16244 14148 16250
rect 14096 16186 14148 16192
rect 13830 15804 14138 15813
rect 13830 15802 13836 15804
rect 13892 15802 13916 15804
rect 13972 15802 13996 15804
rect 14052 15802 14076 15804
rect 14132 15802 14138 15804
rect 13892 15750 13894 15802
rect 14074 15750 14076 15802
rect 13830 15748 13836 15750
rect 13892 15748 13916 15750
rect 13972 15748 13996 15750
rect 14052 15748 14076 15750
rect 14132 15748 14138 15750
rect 13830 15739 14138 15748
rect 14280 15564 14332 15570
rect 14476 15552 14504 20470
rect 14568 19718 14596 22442
rect 14660 22234 14688 22510
rect 14648 22228 14700 22234
rect 14648 22170 14700 22176
rect 14660 21554 14688 22170
rect 14648 21548 14700 21554
rect 14648 21490 14700 21496
rect 14832 20596 14884 20602
rect 14832 20538 14884 20544
rect 14844 20262 14872 20538
rect 14648 20256 14700 20262
rect 14648 20198 14700 20204
rect 14740 20256 14792 20262
rect 14740 20198 14792 20204
rect 14832 20256 14884 20262
rect 14832 20198 14884 20204
rect 14660 20058 14688 20198
rect 14648 20052 14700 20058
rect 14648 19994 14700 20000
rect 14648 19848 14700 19854
rect 14648 19790 14700 19796
rect 14556 19712 14608 19718
rect 14556 19654 14608 19660
rect 14660 18766 14688 19790
rect 14752 19514 14780 20198
rect 14936 19836 14964 24704
rect 15200 24608 15252 24614
rect 15200 24550 15252 24556
rect 15212 24410 15240 24550
rect 15304 24410 15332 26250
rect 15580 26042 15608 26386
rect 15568 26036 15620 26042
rect 15568 25978 15620 25984
rect 15476 25424 15528 25430
rect 15476 25366 15528 25372
rect 15384 25152 15436 25158
rect 15384 25094 15436 25100
rect 15200 24404 15252 24410
rect 15200 24346 15252 24352
rect 15292 24404 15344 24410
rect 15292 24346 15344 24352
rect 15396 24274 15424 25094
rect 15488 24410 15516 25366
rect 15672 25158 15700 26454
rect 15936 26376 15988 26382
rect 15936 26318 15988 26324
rect 15844 25764 15896 25770
rect 15844 25706 15896 25712
rect 15660 25152 15712 25158
rect 15660 25094 15712 25100
rect 15752 25152 15804 25158
rect 15752 25094 15804 25100
rect 15764 24954 15792 25094
rect 15568 24948 15620 24954
rect 15568 24890 15620 24896
rect 15752 24948 15804 24954
rect 15752 24890 15804 24896
rect 15580 24857 15608 24890
rect 15566 24848 15622 24857
rect 15566 24783 15622 24792
rect 15660 24608 15712 24614
rect 15660 24550 15712 24556
rect 15476 24404 15528 24410
rect 15476 24346 15528 24352
rect 15016 24268 15068 24274
rect 15016 24210 15068 24216
rect 15384 24268 15436 24274
rect 15384 24210 15436 24216
rect 15568 24268 15620 24274
rect 15568 24210 15620 24216
rect 15028 23526 15056 24210
rect 15476 24200 15528 24206
rect 15476 24142 15528 24148
rect 15200 24064 15252 24070
rect 15200 24006 15252 24012
rect 15212 23798 15240 24006
rect 15200 23792 15252 23798
rect 15200 23734 15252 23740
rect 15488 23662 15516 24142
rect 15580 23866 15608 24210
rect 15568 23860 15620 23866
rect 15568 23802 15620 23808
rect 15476 23656 15528 23662
rect 15476 23598 15528 23604
rect 15016 23520 15068 23526
rect 15016 23462 15068 23468
rect 15488 23322 15516 23598
rect 15476 23316 15528 23322
rect 15476 23258 15528 23264
rect 15016 22976 15068 22982
rect 15016 22918 15068 22924
rect 15028 22574 15056 22918
rect 15016 22568 15068 22574
rect 15016 22510 15068 22516
rect 15200 21004 15252 21010
rect 15200 20946 15252 20952
rect 15108 20800 15160 20806
rect 15108 20742 15160 20748
rect 14844 19808 14964 19836
rect 14740 19508 14792 19514
rect 14740 19450 14792 19456
rect 14556 18760 14608 18766
rect 14556 18702 14608 18708
rect 14648 18760 14700 18766
rect 14648 18702 14700 18708
rect 14332 15524 14504 15552
rect 14280 15506 14332 15512
rect 13820 15496 13872 15502
rect 13820 15438 13872 15444
rect 13832 15162 13860 15438
rect 13912 15360 13964 15366
rect 13912 15302 13964 15308
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 13924 15026 13952 15302
rect 14568 15094 14596 18702
rect 14844 17626 14872 19808
rect 15016 19712 15068 19718
rect 15016 19654 15068 19660
rect 15120 19666 15148 20742
rect 15212 20058 15240 20946
rect 15672 20618 15700 24550
rect 15856 23866 15884 25706
rect 15948 24614 15976 26318
rect 16592 26314 16620 27118
rect 16684 26314 16712 27610
rect 16776 27586 16820 27614
rect 16868 27614 16896 27832
rect 16868 27586 16988 27614
rect 16776 26450 16804 27586
rect 16960 27538 16988 27586
rect 16948 27532 17000 27538
rect 16948 27474 17000 27480
rect 17052 27418 17080 28966
rect 17144 28422 17172 29242
rect 17604 29034 17632 29446
rect 17592 29028 17644 29034
rect 17592 28970 17644 28976
rect 17592 28620 17644 28626
rect 17592 28562 17644 28568
rect 17132 28416 17184 28422
rect 17132 28358 17184 28364
rect 17188 28316 17496 28325
rect 17188 28314 17194 28316
rect 17250 28314 17274 28316
rect 17330 28314 17354 28316
rect 17410 28314 17434 28316
rect 17490 28314 17496 28316
rect 17250 28262 17252 28314
rect 17432 28262 17434 28314
rect 17188 28260 17194 28262
rect 17250 28260 17274 28262
rect 17330 28260 17354 28262
rect 17410 28260 17434 28262
rect 17490 28260 17496 28262
rect 17188 28251 17496 28260
rect 17132 28008 17184 28014
rect 17132 27950 17184 27956
rect 16868 27390 17080 27418
rect 16764 26444 16816 26450
rect 16764 26386 16816 26392
rect 16868 26330 16896 27390
rect 16948 27328 17000 27334
rect 17144 27316 17172 27950
rect 17224 27872 17276 27878
rect 17222 27840 17224 27849
rect 17276 27840 17278 27849
rect 17222 27775 17278 27784
rect 17604 27713 17632 28562
rect 17222 27704 17278 27713
rect 17222 27639 17224 27648
rect 17276 27639 17278 27648
rect 17590 27704 17646 27713
rect 17590 27639 17646 27648
rect 17224 27610 17276 27616
rect 16948 27270 17000 27276
rect 17052 27288 17172 27316
rect 16960 27130 16988 27270
rect 16948 27124 17000 27130
rect 16948 27066 17000 27072
rect 16580 26308 16632 26314
rect 16580 26250 16632 26256
rect 16672 26308 16724 26314
rect 16672 26250 16724 26256
rect 16776 26302 16896 26330
rect 16304 25764 16356 25770
rect 16304 25706 16356 25712
rect 16316 24954 16344 25706
rect 16396 25356 16448 25362
rect 16396 25298 16448 25304
rect 16408 24954 16436 25298
rect 16672 25152 16724 25158
rect 16672 25094 16724 25100
rect 16304 24948 16356 24954
rect 16304 24890 16356 24896
rect 16396 24948 16448 24954
rect 16396 24890 16448 24896
rect 16304 24744 16356 24750
rect 16304 24686 16356 24692
rect 15936 24608 15988 24614
rect 15936 24550 15988 24556
rect 16316 24410 16344 24686
rect 16304 24404 16356 24410
rect 16304 24346 16356 24352
rect 16408 24206 16436 24890
rect 16684 24818 16712 25094
rect 16580 24812 16632 24818
rect 16580 24754 16632 24760
rect 16672 24812 16724 24818
rect 16672 24754 16724 24760
rect 16592 24410 16620 24754
rect 16776 24698 16804 26302
rect 16856 26240 16908 26246
rect 16856 26182 16908 26188
rect 16868 25498 16896 26182
rect 17052 25906 17080 27288
rect 17188 27228 17496 27237
rect 17188 27226 17194 27228
rect 17250 27226 17274 27228
rect 17330 27226 17354 27228
rect 17410 27226 17434 27228
rect 17490 27226 17496 27228
rect 17250 27174 17252 27226
rect 17432 27174 17434 27226
rect 17188 27172 17194 27174
rect 17250 27172 17274 27174
rect 17330 27172 17354 27174
rect 17410 27172 17434 27174
rect 17490 27172 17496 27174
rect 17188 27163 17496 27172
rect 17500 26920 17552 26926
rect 17500 26862 17552 26868
rect 17408 26852 17460 26858
rect 17408 26794 17460 26800
rect 17420 26382 17448 26794
rect 17512 26586 17540 26862
rect 17500 26580 17552 26586
rect 17500 26522 17552 26528
rect 17408 26376 17460 26382
rect 17408 26318 17460 26324
rect 17592 26308 17644 26314
rect 17592 26250 17644 26256
rect 17188 26140 17496 26149
rect 17188 26138 17194 26140
rect 17250 26138 17274 26140
rect 17330 26138 17354 26140
rect 17410 26138 17434 26140
rect 17490 26138 17496 26140
rect 17250 26086 17252 26138
rect 17432 26086 17434 26138
rect 17188 26084 17194 26086
rect 17250 26084 17274 26086
rect 17330 26084 17354 26086
rect 17410 26084 17434 26086
rect 17490 26084 17496 26086
rect 17188 26075 17496 26084
rect 17040 25900 17092 25906
rect 17040 25842 17092 25848
rect 16856 25492 16908 25498
rect 16856 25434 16908 25440
rect 16684 24670 16804 24698
rect 16580 24404 16632 24410
rect 16580 24346 16632 24352
rect 16396 24200 16448 24206
rect 16396 24142 16448 24148
rect 15844 23860 15896 23866
rect 15844 23802 15896 23808
rect 16580 23316 16632 23322
rect 16580 23258 16632 23264
rect 16592 22642 16620 23258
rect 16580 22636 16632 22642
rect 16580 22578 16632 22584
rect 16684 22438 16712 24670
rect 16764 24268 16816 24274
rect 16764 24210 16816 24216
rect 16672 22432 16724 22438
rect 16672 22374 16724 22380
rect 16580 22228 16632 22234
rect 16580 22170 16632 22176
rect 16592 22098 16620 22170
rect 16580 22092 16632 22098
rect 16580 22034 16632 22040
rect 16672 22092 16724 22098
rect 16672 22034 16724 22040
rect 16120 22024 16172 22030
rect 16120 21966 16172 21972
rect 16304 22024 16356 22030
rect 16304 21966 16356 21972
rect 15752 21888 15804 21894
rect 15752 21830 15804 21836
rect 15764 20788 15792 21830
rect 16132 21350 16160 21966
rect 16212 21888 16264 21894
rect 16212 21830 16264 21836
rect 16224 21622 16252 21830
rect 16316 21622 16344 21966
rect 16684 21690 16712 22034
rect 16672 21684 16724 21690
rect 16672 21626 16724 21632
rect 16212 21616 16264 21622
rect 16212 21558 16264 21564
rect 16304 21616 16356 21622
rect 16304 21558 16356 21564
rect 16120 21344 16172 21350
rect 16120 21286 16172 21292
rect 15936 20868 15988 20874
rect 15936 20810 15988 20816
rect 15844 20800 15896 20806
rect 15764 20760 15844 20788
rect 15844 20742 15896 20748
rect 15672 20590 15792 20618
rect 15292 20256 15344 20262
rect 15292 20198 15344 20204
rect 15200 20052 15252 20058
rect 15200 19994 15252 20000
rect 15304 19990 15332 20198
rect 15568 20052 15620 20058
rect 15620 20012 15700 20040
rect 15568 19994 15620 20000
rect 15292 19984 15344 19990
rect 15292 19926 15344 19932
rect 15028 19446 15056 19654
rect 15120 19638 15424 19666
rect 15292 19508 15344 19514
rect 15292 19450 15344 19456
rect 15016 19440 15068 19446
rect 14922 19408 14978 19417
rect 15016 19382 15068 19388
rect 15200 19440 15252 19446
rect 15200 19382 15252 19388
rect 14922 19343 14978 19352
rect 14936 19242 14964 19343
rect 14924 19236 14976 19242
rect 14924 19178 14976 19184
rect 14924 18896 14976 18902
rect 14924 18838 14976 18844
rect 14660 17598 14872 17626
rect 14660 16017 14688 17598
rect 14740 17536 14792 17542
rect 14740 17478 14792 17484
rect 14752 17066 14780 17478
rect 14740 17060 14792 17066
rect 14740 17002 14792 17008
rect 14832 16992 14884 16998
rect 14832 16934 14884 16940
rect 14646 16008 14702 16017
rect 14844 15978 14872 16934
rect 14936 16114 14964 18838
rect 15028 18290 15056 19382
rect 15108 19168 15160 19174
rect 15108 19110 15160 19116
rect 15120 18426 15148 19110
rect 15108 18420 15160 18426
rect 15108 18362 15160 18368
rect 15016 18284 15068 18290
rect 15016 18226 15068 18232
rect 15120 18154 15148 18362
rect 15212 18154 15240 19382
rect 15108 18148 15160 18154
rect 15108 18090 15160 18096
rect 15200 18148 15252 18154
rect 15200 18090 15252 18096
rect 15120 17882 15148 18090
rect 15108 17876 15160 17882
rect 15108 17818 15160 17824
rect 15212 17746 15240 18090
rect 15304 17882 15332 19450
rect 15396 19378 15424 19638
rect 15384 19372 15436 19378
rect 15384 19314 15436 19320
rect 15396 18834 15424 19314
rect 15476 19304 15528 19310
rect 15476 19246 15528 19252
rect 15568 19304 15620 19310
rect 15568 19246 15620 19252
rect 15384 18828 15436 18834
rect 15384 18770 15436 18776
rect 15488 18222 15516 19246
rect 15580 18970 15608 19246
rect 15568 18964 15620 18970
rect 15568 18906 15620 18912
rect 15476 18216 15528 18222
rect 15476 18158 15528 18164
rect 15292 17876 15344 17882
rect 15292 17818 15344 17824
rect 15200 17740 15252 17746
rect 15200 17682 15252 17688
rect 15292 17604 15344 17610
rect 15120 17564 15292 17592
rect 15016 17332 15068 17338
rect 15016 17274 15068 17280
rect 15028 17202 15056 17274
rect 15016 17196 15068 17202
rect 15016 17138 15068 17144
rect 15028 16674 15056 17138
rect 15120 16794 15148 17564
rect 15292 17546 15344 17552
rect 15108 16788 15160 16794
rect 15108 16730 15160 16736
rect 15028 16646 15148 16674
rect 14924 16108 14976 16114
rect 14924 16050 14976 16056
rect 14646 15943 14702 15952
rect 14832 15972 14884 15978
rect 14832 15914 14884 15920
rect 14832 15360 14884 15366
rect 14832 15302 14884 15308
rect 14740 15156 14792 15162
rect 14740 15098 14792 15104
rect 14096 15088 14148 15094
rect 14096 15030 14148 15036
rect 14556 15088 14608 15094
rect 14556 15030 14608 15036
rect 13912 15020 13964 15026
rect 13912 14962 13964 14968
rect 14108 14890 14136 15030
rect 14372 14952 14424 14958
rect 14372 14894 14424 14900
rect 14096 14884 14148 14890
rect 14096 14826 14148 14832
rect 13830 14716 14138 14725
rect 13830 14714 13836 14716
rect 13892 14714 13916 14716
rect 13972 14714 13996 14716
rect 14052 14714 14076 14716
rect 14132 14714 14138 14716
rect 13892 14662 13894 14714
rect 14074 14662 14076 14714
rect 13830 14660 13836 14662
rect 13892 14660 13916 14662
rect 13972 14660 13996 14662
rect 14052 14660 14076 14662
rect 14132 14660 14138 14662
rect 13830 14651 14138 14660
rect 13636 14612 13688 14618
rect 13636 14554 13688 14560
rect 14384 13938 14412 14894
rect 14568 14090 14596 15030
rect 14752 14958 14780 15098
rect 14740 14952 14792 14958
rect 14740 14894 14792 14900
rect 14844 14618 14872 15302
rect 14924 14952 14976 14958
rect 14924 14894 14976 14900
rect 14832 14612 14884 14618
rect 14832 14554 14884 14560
rect 14936 14482 14964 14894
rect 14924 14476 14976 14482
rect 14924 14418 14976 14424
rect 14648 14272 14700 14278
rect 14700 14232 14780 14260
rect 14648 14214 14700 14220
rect 14568 14062 14688 14090
rect 14372 13932 14424 13938
rect 14372 13874 14424 13880
rect 14556 13864 14608 13870
rect 13556 13790 13768 13818
rect 14556 13806 14608 13812
rect 13636 13728 13688 13734
rect 13636 13670 13688 13676
rect 13648 13190 13676 13670
rect 13740 13512 13768 13790
rect 14188 13728 14240 13734
rect 14188 13670 14240 13676
rect 14280 13728 14332 13734
rect 14280 13670 14332 13676
rect 14464 13728 14516 13734
rect 14464 13670 14516 13676
rect 13830 13628 14138 13637
rect 13830 13626 13836 13628
rect 13892 13626 13916 13628
rect 13972 13626 13996 13628
rect 14052 13626 14076 13628
rect 14132 13626 14138 13628
rect 13892 13574 13894 13626
rect 14074 13574 14076 13626
rect 13830 13572 13836 13574
rect 13892 13572 13916 13574
rect 13972 13572 13996 13574
rect 14052 13572 14076 13574
rect 14132 13572 14138 13574
rect 13830 13563 14138 13572
rect 13740 13484 13860 13512
rect 13636 13184 13688 13190
rect 13636 13126 13688 13132
rect 13360 12096 13412 12102
rect 13360 12038 13412 12044
rect 13268 10464 13320 10470
rect 13268 10406 13320 10412
rect 13280 10130 13308 10406
rect 13372 10130 13400 12038
rect 13648 10606 13676 13126
rect 13832 12850 13860 13484
rect 13912 13320 13964 13326
rect 13912 13262 13964 13268
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13832 12628 13860 12786
rect 13924 12714 13952 13262
rect 14200 12850 14228 13670
rect 14292 13394 14320 13670
rect 14476 13530 14504 13670
rect 14464 13524 14516 13530
rect 14464 13466 14516 13472
rect 14280 13388 14332 13394
rect 14280 13330 14332 13336
rect 14188 12844 14240 12850
rect 14188 12786 14240 12792
rect 13912 12708 13964 12714
rect 13912 12650 13964 12656
rect 13740 12600 13860 12628
rect 13740 11898 13768 12600
rect 13830 12540 14138 12549
rect 13830 12538 13836 12540
rect 13892 12538 13916 12540
rect 13972 12538 13996 12540
rect 14052 12538 14076 12540
rect 14132 12538 14138 12540
rect 13892 12486 13894 12538
rect 14074 12486 14076 12538
rect 13830 12484 13836 12486
rect 13892 12484 13916 12486
rect 13972 12484 13996 12486
rect 14052 12484 14076 12486
rect 14132 12484 14138 12486
rect 13830 12475 14138 12484
rect 14476 12288 14504 13466
rect 14568 12986 14596 13806
rect 14556 12980 14608 12986
rect 14556 12922 14608 12928
rect 14556 12300 14608 12306
rect 14476 12260 14556 12288
rect 14556 12242 14608 12248
rect 14372 12096 14424 12102
rect 14372 12038 14424 12044
rect 13728 11892 13780 11898
rect 13728 11834 13780 11840
rect 14188 11620 14240 11626
rect 14188 11562 14240 11568
rect 14280 11620 14332 11626
rect 14280 11562 14332 11568
rect 13830 11452 14138 11461
rect 13830 11450 13836 11452
rect 13892 11450 13916 11452
rect 13972 11450 13996 11452
rect 14052 11450 14076 11452
rect 14132 11450 14138 11452
rect 13892 11398 13894 11450
rect 14074 11398 14076 11450
rect 13830 11396 13836 11398
rect 13892 11396 13916 11398
rect 13972 11396 13996 11398
rect 14052 11396 14076 11398
rect 14132 11396 14138 11398
rect 13830 11387 14138 11396
rect 14200 11354 14228 11562
rect 14188 11348 14240 11354
rect 14188 11290 14240 11296
rect 14292 11218 14320 11562
rect 14188 11212 14240 11218
rect 14188 11154 14240 11160
rect 14280 11212 14332 11218
rect 14280 11154 14332 11160
rect 13636 10600 13688 10606
rect 13636 10542 13688 10548
rect 13452 10532 13504 10538
rect 13452 10474 13504 10480
rect 13464 10266 13492 10474
rect 13830 10364 14138 10373
rect 13830 10362 13836 10364
rect 13892 10362 13916 10364
rect 13972 10362 13996 10364
rect 14052 10362 14076 10364
rect 14132 10362 14138 10364
rect 13892 10310 13894 10362
rect 14074 10310 14076 10362
rect 13830 10308 13836 10310
rect 13892 10308 13916 10310
rect 13972 10308 13996 10310
rect 14052 10308 14076 10310
rect 14132 10308 14138 10310
rect 13830 10299 14138 10308
rect 13452 10260 13504 10266
rect 13452 10202 13504 10208
rect 14200 10130 14228 11154
rect 14280 11008 14332 11014
rect 14280 10950 14332 10956
rect 14292 10130 14320 10950
rect 13268 10124 13320 10130
rect 13268 10066 13320 10072
rect 13360 10124 13412 10130
rect 13360 10066 13412 10072
rect 14188 10124 14240 10130
rect 14188 10066 14240 10072
rect 14280 10124 14332 10130
rect 14280 10066 14332 10072
rect 14200 9518 14228 10066
rect 14384 9518 14412 12038
rect 14464 11688 14516 11694
rect 14464 11630 14516 11636
rect 14476 10062 14504 11630
rect 14568 11354 14596 12242
rect 14556 11348 14608 11354
rect 14556 11290 14608 11296
rect 14556 10260 14608 10266
rect 14556 10202 14608 10208
rect 14464 10056 14516 10062
rect 14464 9998 14516 10004
rect 14464 9920 14516 9926
rect 14464 9862 14516 9868
rect 14476 9518 14504 9862
rect 13176 9512 13228 9518
rect 13176 9454 13228 9460
rect 14188 9512 14240 9518
rect 14188 9454 14240 9460
rect 14372 9512 14424 9518
rect 14372 9454 14424 9460
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14568 9466 14596 10202
rect 14660 9602 14688 14062
rect 14752 13938 14780 14232
rect 14832 14000 14884 14006
rect 14832 13942 14884 13948
rect 14740 13932 14792 13938
rect 14740 13874 14792 13880
rect 14752 13394 14780 13874
rect 14740 13388 14792 13394
rect 14740 13330 14792 13336
rect 14752 12442 14780 13330
rect 14740 12436 14792 12442
rect 14740 12378 14792 12384
rect 14752 11762 14780 12378
rect 14844 12306 14872 13942
rect 15016 13728 15068 13734
rect 15016 13670 15068 13676
rect 15028 12782 15056 13670
rect 15016 12776 15068 12782
rect 15016 12718 15068 12724
rect 15120 12714 15148 16646
rect 15384 16652 15436 16658
rect 15384 16594 15436 16600
rect 15292 16448 15344 16454
rect 15292 16390 15344 16396
rect 15304 16046 15332 16390
rect 15292 16040 15344 16046
rect 15292 15982 15344 15988
rect 15200 15564 15252 15570
rect 15200 15506 15252 15512
rect 15212 15162 15240 15506
rect 15200 15156 15252 15162
rect 15200 15098 15252 15104
rect 15396 15026 15424 16594
rect 15568 16244 15620 16250
rect 15568 16186 15620 16192
rect 15476 16040 15528 16046
rect 15474 16008 15476 16017
rect 15528 16008 15530 16017
rect 15474 15943 15530 15952
rect 15476 15904 15528 15910
rect 15476 15846 15528 15852
rect 15488 15638 15516 15846
rect 15476 15632 15528 15638
rect 15476 15574 15528 15580
rect 15580 15502 15608 16186
rect 15672 15706 15700 20012
rect 15764 16114 15792 20590
rect 15856 20330 15884 20742
rect 15948 20330 15976 20810
rect 15844 20324 15896 20330
rect 15844 20266 15896 20272
rect 15936 20324 15988 20330
rect 15936 20266 15988 20272
rect 15856 19378 15884 20266
rect 16028 19916 16080 19922
rect 16028 19858 16080 19864
rect 16040 19514 16068 19858
rect 16120 19712 16172 19718
rect 16120 19654 16172 19660
rect 16028 19508 16080 19514
rect 16028 19450 16080 19456
rect 15844 19372 15896 19378
rect 15844 19314 15896 19320
rect 16132 19310 16160 19654
rect 16120 19304 16172 19310
rect 16120 19246 16172 19252
rect 16224 18426 16252 21558
rect 16316 21146 16344 21558
rect 16776 21332 16804 24210
rect 16868 22098 16896 25434
rect 17040 25356 17092 25362
rect 17040 25298 17092 25304
rect 16948 25288 17000 25294
rect 16948 25230 17000 25236
rect 16960 24274 16988 25230
rect 17052 24274 17080 25298
rect 17188 25052 17496 25061
rect 17188 25050 17194 25052
rect 17250 25050 17274 25052
rect 17330 25050 17354 25052
rect 17410 25050 17434 25052
rect 17490 25050 17496 25052
rect 17250 24998 17252 25050
rect 17432 24998 17434 25050
rect 17188 24996 17194 24998
rect 17250 24996 17274 24998
rect 17330 24996 17354 24998
rect 17410 24996 17434 24998
rect 17490 24996 17496 24998
rect 17188 24987 17496 24996
rect 17604 24834 17632 26250
rect 17512 24806 17632 24834
rect 17408 24744 17460 24750
rect 17408 24686 17460 24692
rect 17224 24608 17276 24614
rect 17224 24550 17276 24556
rect 17316 24608 17368 24614
rect 17316 24550 17368 24556
rect 17236 24410 17264 24550
rect 17328 24410 17356 24550
rect 17420 24410 17448 24686
rect 17224 24404 17276 24410
rect 17224 24346 17276 24352
rect 17316 24404 17368 24410
rect 17316 24346 17368 24352
rect 17408 24404 17460 24410
rect 17408 24346 17460 24352
rect 17512 24274 17540 24806
rect 17696 24698 17724 30552
rect 17776 30534 17828 30540
rect 18064 29306 18092 30738
rect 19076 30734 19104 31600
rect 20548 31226 20576 31600
rect 20456 31198 20576 31226
rect 21088 31204 21140 31210
rect 19432 31136 19484 31142
rect 19432 31078 19484 31084
rect 19444 30802 19472 31078
rect 19616 30864 19668 30870
rect 19616 30806 19668 30812
rect 19708 30864 19760 30870
rect 19760 30812 19840 30818
rect 19708 30806 19840 30812
rect 19432 30796 19484 30802
rect 19432 30738 19484 30744
rect 19064 30728 19116 30734
rect 19064 30670 19116 30676
rect 18144 30660 18196 30666
rect 18144 30602 18196 30608
rect 18156 30190 18184 30602
rect 18236 30592 18288 30598
rect 18236 30534 18288 30540
rect 18144 30184 18196 30190
rect 18144 30126 18196 30132
rect 18248 29782 18276 30534
rect 19444 30274 19472 30738
rect 19524 30592 19576 30598
rect 19524 30534 19576 30540
rect 19352 30246 19472 30274
rect 18236 29776 18288 29782
rect 18236 29718 18288 29724
rect 18972 29776 19024 29782
rect 18972 29718 19024 29724
rect 18984 29617 19012 29718
rect 19248 29640 19300 29646
rect 18970 29608 19026 29617
rect 19248 29582 19300 29588
rect 18970 29543 19026 29552
rect 18144 29504 18196 29510
rect 18144 29446 18196 29452
rect 19156 29504 19208 29510
rect 19156 29446 19208 29452
rect 18052 29300 18104 29306
rect 18052 29242 18104 29248
rect 18156 29102 18184 29446
rect 19168 29102 19196 29446
rect 19260 29102 19288 29582
rect 19352 29306 19380 30246
rect 19432 30184 19484 30190
rect 19432 30126 19484 30132
rect 19444 29696 19472 30126
rect 19536 30122 19564 30534
rect 19524 30116 19576 30122
rect 19524 30058 19576 30064
rect 19524 29708 19576 29714
rect 19444 29668 19524 29696
rect 19524 29650 19576 29656
rect 19340 29300 19392 29306
rect 19340 29242 19392 29248
rect 19352 29102 19380 29242
rect 18144 29096 18196 29102
rect 18144 29038 18196 29044
rect 18696 29096 18748 29102
rect 18696 29038 18748 29044
rect 19156 29096 19208 29102
rect 19156 29038 19208 29044
rect 19248 29096 19300 29102
rect 19248 29038 19300 29044
rect 19340 29096 19392 29102
rect 19340 29038 19392 29044
rect 18236 29028 18288 29034
rect 18236 28970 18288 28976
rect 17776 28008 17828 28014
rect 17776 27950 17828 27956
rect 17788 27674 17816 27950
rect 17776 27668 17828 27674
rect 17776 27610 17828 27616
rect 17776 27328 17828 27334
rect 17776 27270 17828 27276
rect 18052 27328 18104 27334
rect 18052 27270 18104 27276
rect 17788 25362 17816 27270
rect 18064 27130 18092 27270
rect 18052 27124 18104 27130
rect 18052 27066 18104 27072
rect 17868 27056 17920 27062
rect 17868 26998 17920 27004
rect 17880 26772 17908 26998
rect 17960 26784 18012 26790
rect 17880 26744 17960 26772
rect 17880 25838 17908 26744
rect 17960 26726 18012 26732
rect 17960 26240 18012 26246
rect 17960 26182 18012 26188
rect 18144 26240 18196 26246
rect 18144 26182 18196 26188
rect 17972 26042 18000 26182
rect 17960 26036 18012 26042
rect 17960 25978 18012 25984
rect 17868 25832 17920 25838
rect 17868 25774 17920 25780
rect 17972 25498 18000 25978
rect 18156 25838 18184 26182
rect 18144 25832 18196 25838
rect 18144 25774 18196 25780
rect 17960 25492 18012 25498
rect 17960 25434 18012 25440
rect 17776 25356 17828 25362
rect 17776 25298 17828 25304
rect 18144 25152 18196 25158
rect 18144 25094 18196 25100
rect 18156 24750 18184 25094
rect 17604 24670 17724 24698
rect 18144 24744 18196 24750
rect 18144 24686 18196 24692
rect 16948 24268 17000 24274
rect 16948 24210 17000 24216
rect 17040 24268 17092 24274
rect 17040 24210 17092 24216
rect 17500 24268 17552 24274
rect 17500 24210 17552 24216
rect 16960 23322 16988 24210
rect 17188 23964 17496 23973
rect 17188 23962 17194 23964
rect 17250 23962 17274 23964
rect 17330 23962 17354 23964
rect 17410 23962 17434 23964
rect 17490 23962 17496 23964
rect 17250 23910 17252 23962
rect 17432 23910 17434 23962
rect 17188 23908 17194 23910
rect 17250 23908 17274 23910
rect 17330 23908 17354 23910
rect 17410 23908 17434 23910
rect 17490 23908 17496 23910
rect 17188 23899 17496 23908
rect 16948 23316 17000 23322
rect 16948 23258 17000 23264
rect 17040 23248 17092 23254
rect 17040 23190 17092 23196
rect 17052 22778 17080 23190
rect 17188 22876 17496 22885
rect 17188 22874 17194 22876
rect 17250 22874 17274 22876
rect 17330 22874 17354 22876
rect 17410 22874 17434 22876
rect 17490 22874 17496 22876
rect 17250 22822 17252 22874
rect 17432 22822 17434 22874
rect 17188 22820 17194 22822
rect 17250 22820 17274 22822
rect 17330 22820 17354 22822
rect 17410 22820 17434 22822
rect 17490 22820 17496 22822
rect 17188 22811 17496 22820
rect 17040 22772 17092 22778
rect 17040 22714 17092 22720
rect 17408 22568 17460 22574
rect 17408 22510 17460 22516
rect 17040 22432 17092 22438
rect 17040 22374 17092 22380
rect 16856 22092 16908 22098
rect 16856 22034 16908 22040
rect 16856 21344 16908 21350
rect 16776 21304 16856 21332
rect 16856 21286 16908 21292
rect 16304 21140 16356 21146
rect 16304 21082 16356 21088
rect 16672 21004 16724 21010
rect 16672 20946 16724 20952
rect 16684 20874 16712 20946
rect 16672 20868 16724 20874
rect 16672 20810 16724 20816
rect 16488 19168 16540 19174
rect 16488 19110 16540 19116
rect 16500 18970 16528 19110
rect 16488 18964 16540 18970
rect 16488 18906 16540 18912
rect 16212 18420 16264 18426
rect 16212 18362 16264 18368
rect 16580 17672 16632 17678
rect 16580 17614 16632 17620
rect 15936 17536 15988 17542
rect 15936 17478 15988 17484
rect 16304 17536 16356 17542
rect 16304 17478 16356 17484
rect 15948 16794 15976 17478
rect 16316 17338 16344 17478
rect 16304 17332 16356 17338
rect 16304 17274 16356 17280
rect 16488 17264 16540 17270
rect 16488 17206 16540 17212
rect 16118 17096 16174 17105
rect 16118 17031 16120 17040
rect 16172 17031 16174 17040
rect 16120 17002 16172 17008
rect 16304 16992 16356 16998
rect 16304 16934 16356 16940
rect 15936 16788 15988 16794
rect 15936 16730 15988 16736
rect 15752 16108 15804 16114
rect 15752 16050 15804 16056
rect 16212 16040 16264 16046
rect 16212 15982 16264 15988
rect 16224 15706 16252 15982
rect 15660 15700 15712 15706
rect 15660 15642 15712 15648
rect 15936 15700 15988 15706
rect 15936 15642 15988 15648
rect 16212 15700 16264 15706
rect 16212 15642 16264 15648
rect 15568 15496 15620 15502
rect 15568 15438 15620 15444
rect 15568 15088 15620 15094
rect 15568 15030 15620 15036
rect 15384 15020 15436 15026
rect 15384 14962 15436 14968
rect 15292 14884 15344 14890
rect 15292 14826 15344 14832
rect 15304 14618 15332 14826
rect 15292 14612 15344 14618
rect 15292 14554 15344 14560
rect 15476 13864 15528 13870
rect 15476 13806 15528 13812
rect 15488 13530 15516 13806
rect 15476 13524 15528 13530
rect 15476 13466 15528 13472
rect 15200 13320 15252 13326
rect 15200 13262 15252 13268
rect 15108 12708 15160 12714
rect 15108 12650 15160 12656
rect 15212 12646 15240 13262
rect 15200 12640 15252 12646
rect 15200 12582 15252 12588
rect 14832 12300 14884 12306
rect 14832 12242 14884 12248
rect 14740 11756 14792 11762
rect 14740 11698 14792 11704
rect 14844 11082 14872 12242
rect 15016 11620 15068 11626
rect 15016 11562 15068 11568
rect 15028 11354 15056 11562
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 15120 11354 15148 11494
rect 15016 11348 15068 11354
rect 15016 11290 15068 11296
rect 15108 11348 15160 11354
rect 15108 11290 15160 11296
rect 14832 11076 14884 11082
rect 14832 11018 14884 11024
rect 14924 10600 14976 10606
rect 14924 10542 14976 10548
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14752 10198 14780 10406
rect 14740 10192 14792 10198
rect 14740 10134 14792 10140
rect 14936 9722 14964 10542
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 15476 10464 15528 10470
rect 15476 10406 15528 10412
rect 14924 9716 14976 9722
rect 14924 9658 14976 9664
rect 14660 9574 15056 9602
rect 13830 9276 14138 9285
rect 13830 9274 13836 9276
rect 13892 9274 13916 9276
rect 13972 9274 13996 9276
rect 14052 9274 14076 9276
rect 14132 9274 14138 9276
rect 13892 9222 13894 9274
rect 14074 9222 14076 9274
rect 13830 9220 13836 9222
rect 13892 9220 13916 9222
rect 13972 9220 13996 9222
rect 14052 9220 14076 9222
rect 14132 9220 14138 9222
rect 13830 9211 14138 9220
rect 14096 9172 14148 9178
rect 14096 9114 14148 9120
rect 13176 9036 13228 9042
rect 13176 8978 13228 8984
rect 13360 9036 13412 9042
rect 13360 8978 13412 8984
rect 13728 9036 13780 9042
rect 13728 8978 13780 8984
rect 13188 8430 13216 8978
rect 13176 8424 13228 8430
rect 13176 8366 13228 8372
rect 13372 8294 13400 8978
rect 13544 8832 13596 8838
rect 13544 8774 13596 8780
rect 13360 8288 13412 8294
rect 13360 8230 13412 8236
rect 13556 5846 13584 8774
rect 13740 8362 13768 8978
rect 14108 8548 14136 9114
rect 14200 9042 14228 9454
rect 14476 9042 14504 9454
rect 14568 9438 14872 9466
rect 14648 9376 14700 9382
rect 14648 9318 14700 9324
rect 14188 9036 14240 9042
rect 14188 8978 14240 8984
rect 14464 9036 14516 9042
rect 14464 8978 14516 8984
rect 14280 8832 14332 8838
rect 14280 8774 14332 8780
rect 14108 8520 14228 8548
rect 13728 8356 13780 8362
rect 13728 8298 13780 8304
rect 13636 8288 13688 8294
rect 13636 8230 13688 8236
rect 13648 7546 13676 8230
rect 13830 8188 14138 8197
rect 13830 8186 13836 8188
rect 13892 8186 13916 8188
rect 13972 8186 13996 8188
rect 14052 8186 14076 8188
rect 14132 8186 14138 8188
rect 13892 8134 13894 8186
rect 14074 8134 14076 8186
rect 13830 8132 13836 8134
rect 13892 8132 13916 8134
rect 13972 8132 13996 8134
rect 14052 8132 14076 8134
rect 14132 8132 14138 8134
rect 13830 8123 14138 8132
rect 14200 8090 14228 8520
rect 14188 8084 14240 8090
rect 14188 8026 14240 8032
rect 14188 7744 14240 7750
rect 14188 7686 14240 7692
rect 13636 7540 13688 7546
rect 13636 7482 13688 7488
rect 13830 7100 14138 7109
rect 13830 7098 13836 7100
rect 13892 7098 13916 7100
rect 13972 7098 13996 7100
rect 14052 7098 14076 7100
rect 14132 7098 14138 7100
rect 13892 7046 13894 7098
rect 14074 7046 14076 7098
rect 13830 7044 13836 7046
rect 13892 7044 13916 7046
rect 13972 7044 13996 7046
rect 14052 7044 14076 7046
rect 14132 7044 14138 7046
rect 13830 7035 14138 7044
rect 14096 6452 14148 6458
rect 14096 6394 14148 6400
rect 13728 6248 13780 6254
rect 14108 6225 14136 6394
rect 13728 6190 13780 6196
rect 14094 6216 14150 6225
rect 13740 5846 13768 6190
rect 14094 6151 14150 6160
rect 13830 6012 14138 6021
rect 13830 6010 13836 6012
rect 13892 6010 13916 6012
rect 13972 6010 13996 6012
rect 14052 6010 14076 6012
rect 14132 6010 14138 6012
rect 13892 5958 13894 6010
rect 14074 5958 14076 6010
rect 13830 5956 13836 5958
rect 13892 5956 13916 5958
rect 13972 5956 13996 5958
rect 14052 5956 14076 5958
rect 14132 5956 14138 5958
rect 13830 5947 14138 5956
rect 14200 5914 14228 7686
rect 14292 6118 14320 8774
rect 14372 8560 14424 8566
rect 14372 8502 14424 8508
rect 14384 6746 14412 8502
rect 14476 8430 14504 8978
rect 14464 8424 14516 8430
rect 14464 8366 14516 8372
rect 14476 7936 14504 8366
rect 14556 7948 14608 7954
rect 14476 7908 14556 7936
rect 14556 7890 14608 7896
rect 14556 7812 14608 7818
rect 14556 7754 14608 7760
rect 14568 7546 14596 7754
rect 14556 7540 14608 7546
rect 14556 7482 14608 7488
rect 14464 7336 14516 7342
rect 14464 7278 14516 7284
rect 14476 7002 14504 7278
rect 14464 6996 14516 7002
rect 14464 6938 14516 6944
rect 14660 6746 14688 9318
rect 14740 8832 14792 8838
rect 14740 8774 14792 8780
rect 14752 8498 14780 8774
rect 14740 8492 14792 8498
rect 14740 8434 14792 8440
rect 14844 8072 14872 9438
rect 14924 9036 14976 9042
rect 14924 8978 14976 8984
rect 14936 8430 14964 8978
rect 14924 8424 14976 8430
rect 14924 8366 14976 8372
rect 14936 8090 14964 8366
rect 15028 8294 15056 9574
rect 15212 9518 15240 10406
rect 15488 9926 15516 10406
rect 15580 10062 15608 15030
rect 15752 12844 15804 12850
rect 15752 12786 15804 12792
rect 15660 12436 15712 12442
rect 15660 12378 15712 12384
rect 15672 12306 15700 12378
rect 15660 12300 15712 12306
rect 15660 12242 15712 12248
rect 15764 11762 15792 12786
rect 15844 12640 15896 12646
rect 15844 12582 15896 12588
rect 15856 12442 15884 12582
rect 15844 12436 15896 12442
rect 15844 12378 15896 12384
rect 15752 11756 15804 11762
rect 15752 11698 15804 11704
rect 15660 10600 15712 10606
rect 15660 10542 15712 10548
rect 15568 10056 15620 10062
rect 15568 9998 15620 10004
rect 15476 9920 15528 9926
rect 15476 9862 15528 9868
rect 15200 9512 15252 9518
rect 15200 9454 15252 9460
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 15396 8974 15424 9318
rect 15488 9042 15516 9862
rect 15672 9042 15700 10542
rect 15764 10062 15792 11698
rect 15948 10266 15976 15642
rect 16224 15026 16252 15642
rect 16212 15020 16264 15026
rect 16212 14962 16264 14968
rect 16316 12850 16344 16934
rect 16500 16794 16528 17206
rect 16488 16788 16540 16794
rect 16488 16730 16540 16736
rect 16500 16250 16528 16730
rect 16488 16244 16540 16250
rect 16488 16186 16540 16192
rect 16488 14272 16540 14278
rect 16488 14214 16540 14220
rect 16500 13530 16528 14214
rect 16488 13524 16540 13530
rect 16488 13466 16540 13472
rect 16304 12844 16356 12850
rect 16304 12786 16356 12792
rect 16212 12776 16264 12782
rect 16212 12718 16264 12724
rect 16224 12442 16252 12718
rect 16212 12436 16264 12442
rect 16212 12378 16264 12384
rect 16592 11694 16620 17614
rect 16684 17134 16712 20810
rect 16868 20466 16896 21286
rect 16856 20460 16908 20466
rect 16856 20402 16908 20408
rect 16948 19916 17000 19922
rect 16948 19858 17000 19864
rect 16960 19514 16988 19858
rect 16948 19508 17000 19514
rect 16948 19450 17000 19456
rect 17052 18952 17080 22374
rect 17420 21962 17448 22510
rect 17408 21956 17460 21962
rect 17408 21898 17460 21904
rect 17188 21788 17496 21797
rect 17188 21786 17194 21788
rect 17250 21786 17274 21788
rect 17330 21786 17354 21788
rect 17410 21786 17434 21788
rect 17490 21786 17496 21788
rect 17250 21734 17252 21786
rect 17432 21734 17434 21786
rect 17188 21732 17194 21734
rect 17250 21732 17274 21734
rect 17330 21732 17354 21734
rect 17410 21732 17434 21734
rect 17490 21732 17496 21734
rect 17188 21723 17496 21732
rect 17188 20700 17496 20709
rect 17188 20698 17194 20700
rect 17250 20698 17274 20700
rect 17330 20698 17354 20700
rect 17410 20698 17434 20700
rect 17490 20698 17496 20700
rect 17250 20646 17252 20698
rect 17432 20646 17434 20698
rect 17188 20644 17194 20646
rect 17250 20644 17274 20646
rect 17330 20644 17354 20646
rect 17410 20644 17434 20646
rect 17490 20644 17496 20646
rect 17188 20635 17496 20644
rect 17188 19612 17496 19621
rect 17188 19610 17194 19612
rect 17250 19610 17274 19612
rect 17330 19610 17354 19612
rect 17410 19610 17434 19612
rect 17490 19610 17496 19612
rect 17250 19558 17252 19610
rect 17432 19558 17434 19610
rect 17188 19556 17194 19558
rect 17250 19556 17274 19558
rect 17330 19556 17354 19558
rect 17410 19556 17434 19558
rect 17490 19556 17496 19558
rect 17188 19547 17496 19556
rect 17604 19310 17632 24670
rect 17868 23180 17920 23186
rect 17868 23122 17920 23128
rect 17880 22778 17908 23122
rect 17960 23112 18012 23118
rect 17960 23054 18012 23060
rect 17868 22772 17920 22778
rect 17868 22714 17920 22720
rect 17868 22568 17920 22574
rect 17868 22510 17920 22516
rect 17684 22432 17736 22438
rect 17684 22374 17736 22380
rect 17696 22234 17724 22374
rect 17684 22228 17736 22234
rect 17684 22170 17736 22176
rect 17696 20398 17724 22170
rect 17776 22092 17828 22098
rect 17880 22080 17908 22510
rect 17828 22052 17908 22080
rect 17776 22034 17828 22040
rect 17684 20392 17736 20398
rect 17788 20380 17816 22034
rect 17868 21888 17920 21894
rect 17868 21830 17920 21836
rect 17880 21146 17908 21830
rect 17972 21486 18000 23054
rect 18248 22642 18276 28970
rect 18708 28762 18736 29038
rect 18880 28960 18932 28966
rect 18880 28902 18932 28908
rect 18696 28756 18748 28762
rect 18696 28698 18748 28704
rect 18892 28694 18920 28902
rect 18880 28688 18932 28694
rect 18880 28630 18932 28636
rect 19536 28558 19564 29650
rect 19628 29510 19656 30806
rect 19720 30790 19840 30806
rect 19708 29708 19760 29714
rect 19708 29650 19760 29656
rect 19616 29504 19668 29510
rect 19616 29446 19668 29452
rect 19720 29306 19748 29650
rect 19708 29300 19760 29306
rect 19708 29242 19760 29248
rect 19616 29232 19668 29238
rect 19812 29186 19840 30790
rect 20076 30592 20128 30598
rect 19616 29174 19668 29180
rect 19628 28626 19656 29174
rect 19720 29158 19840 29186
rect 19904 30552 20076 30580
rect 19616 28620 19668 28626
rect 19616 28562 19668 28568
rect 19524 28552 19576 28558
rect 19720 28506 19748 29158
rect 19800 29096 19852 29102
rect 19800 29038 19852 29044
rect 19524 28494 19576 28500
rect 19536 27878 19564 28494
rect 19628 28478 19748 28506
rect 18328 27872 18380 27878
rect 18328 27814 18380 27820
rect 18512 27872 18564 27878
rect 18512 27814 18564 27820
rect 19524 27872 19576 27878
rect 19524 27814 19576 27820
rect 18340 27130 18368 27814
rect 18524 27606 18552 27814
rect 18512 27600 18564 27606
rect 18512 27542 18564 27548
rect 19536 27538 19564 27814
rect 19340 27532 19392 27538
rect 19340 27474 19392 27480
rect 19524 27532 19576 27538
rect 19524 27474 19576 27480
rect 18420 27396 18472 27402
rect 18420 27338 18472 27344
rect 18432 27130 18460 27338
rect 19352 27130 19380 27474
rect 18328 27124 18380 27130
rect 18328 27066 18380 27072
rect 18420 27124 18472 27130
rect 18420 27066 18472 27072
rect 19340 27124 19392 27130
rect 19340 27066 19392 27072
rect 19536 26994 19564 27474
rect 19524 26988 19576 26994
rect 19524 26930 19576 26936
rect 18512 26920 18564 26926
rect 18512 26862 18564 26868
rect 18420 26240 18472 26246
rect 18420 26182 18472 26188
rect 18432 25906 18460 26182
rect 18524 26042 18552 26862
rect 18696 26784 18748 26790
rect 18696 26726 18748 26732
rect 18708 26586 18736 26726
rect 19536 26586 19564 26930
rect 18696 26580 18748 26586
rect 18696 26522 18748 26528
rect 19524 26580 19576 26586
rect 19524 26522 19576 26528
rect 19524 26444 19576 26450
rect 19524 26386 19576 26392
rect 19536 26042 19564 26386
rect 18512 26036 18564 26042
rect 18512 25978 18564 25984
rect 19524 26036 19576 26042
rect 19524 25978 19576 25984
rect 19628 25922 19656 28478
rect 19812 27538 19840 29038
rect 19800 27532 19852 27538
rect 19800 27474 19852 27480
rect 19812 27418 19840 27474
rect 18420 25900 18472 25906
rect 18420 25842 18472 25848
rect 19536 25894 19656 25922
rect 19720 27390 19840 27418
rect 18328 25424 18380 25430
rect 18328 25366 18380 25372
rect 18340 24274 18368 25366
rect 18432 24274 18460 25842
rect 18512 24608 18564 24614
rect 18512 24550 18564 24556
rect 18524 24410 18552 24550
rect 18512 24404 18564 24410
rect 18512 24346 18564 24352
rect 18328 24268 18380 24274
rect 18328 24210 18380 24216
rect 18420 24268 18472 24274
rect 18420 24210 18472 24216
rect 18420 24064 18472 24070
rect 18420 24006 18472 24012
rect 18432 23866 18460 24006
rect 18420 23860 18472 23866
rect 18420 23802 18472 23808
rect 18524 23798 18552 24346
rect 19340 24336 19392 24342
rect 19340 24278 19392 24284
rect 18788 24268 18840 24274
rect 18788 24210 18840 24216
rect 18696 24200 18748 24206
rect 18696 24142 18748 24148
rect 18512 23792 18564 23798
rect 18512 23734 18564 23740
rect 18708 23526 18736 24142
rect 18800 23662 18828 24210
rect 18788 23656 18840 23662
rect 18788 23598 18840 23604
rect 18696 23520 18748 23526
rect 18696 23462 18748 23468
rect 18708 22778 18736 23462
rect 19352 23322 19380 24278
rect 19432 23588 19484 23594
rect 19432 23530 19484 23536
rect 19340 23316 19392 23322
rect 19340 23258 19392 23264
rect 19444 23202 19472 23530
rect 19536 23526 19564 25894
rect 19720 25498 19748 27390
rect 19800 27328 19852 27334
rect 19800 27270 19852 27276
rect 19812 26926 19840 27270
rect 19800 26920 19852 26926
rect 19800 26862 19852 26868
rect 19800 26444 19852 26450
rect 19800 26386 19852 26392
rect 19812 25906 19840 26386
rect 19800 25900 19852 25906
rect 19800 25842 19852 25848
rect 19708 25492 19760 25498
rect 19708 25434 19760 25440
rect 19812 24818 19840 25842
rect 19800 24812 19852 24818
rect 19800 24754 19852 24760
rect 19708 24608 19760 24614
rect 19708 24550 19760 24556
rect 19720 24138 19748 24550
rect 19812 24274 19840 24754
rect 19800 24268 19852 24274
rect 19800 24210 19852 24216
rect 19708 24132 19760 24138
rect 19708 24074 19760 24080
rect 19904 23882 19932 30552
rect 20076 30534 20128 30540
rect 20456 30190 20484 31198
rect 21088 31146 21140 31152
rect 20546 31036 20854 31045
rect 20546 31034 20552 31036
rect 20608 31034 20632 31036
rect 20688 31034 20712 31036
rect 20768 31034 20792 31036
rect 20848 31034 20854 31036
rect 20608 30982 20610 31034
rect 20790 30982 20792 31034
rect 20546 30980 20552 30982
rect 20608 30980 20632 30982
rect 20688 30980 20712 30982
rect 20768 30980 20792 30982
rect 20848 30980 20854 30982
rect 20546 30971 20854 30980
rect 21100 30938 21128 31146
rect 21088 30932 21140 30938
rect 21088 30874 21140 30880
rect 20812 30728 20864 30734
rect 20812 30670 20864 30676
rect 20824 30394 20852 30670
rect 20812 30388 20864 30394
rect 20812 30330 20864 30336
rect 20444 30184 20496 30190
rect 20824 30161 20852 30330
rect 20444 30126 20496 30132
rect 20810 30152 20866 30161
rect 20810 30087 20866 30096
rect 20996 30048 21048 30054
rect 20996 29990 21048 29996
rect 20546 29948 20854 29957
rect 20546 29946 20552 29948
rect 20608 29946 20632 29948
rect 20688 29946 20712 29948
rect 20768 29946 20792 29948
rect 20848 29946 20854 29948
rect 20608 29894 20610 29946
rect 20790 29894 20792 29946
rect 20546 29892 20552 29894
rect 20608 29892 20632 29894
rect 20688 29892 20712 29894
rect 20768 29892 20792 29894
rect 20848 29892 20854 29894
rect 20546 29883 20854 29892
rect 20628 29844 20680 29850
rect 20628 29786 20680 29792
rect 20640 29510 20668 29786
rect 20076 29504 20128 29510
rect 20076 29446 20128 29452
rect 20628 29504 20680 29510
rect 20628 29446 20680 29452
rect 20088 27606 20116 29446
rect 20640 29170 20668 29446
rect 20628 29164 20680 29170
rect 20628 29106 20680 29112
rect 20546 28860 20854 28869
rect 20546 28858 20552 28860
rect 20608 28858 20632 28860
rect 20688 28858 20712 28860
rect 20768 28858 20792 28860
rect 20848 28858 20854 28860
rect 20608 28806 20610 28858
rect 20790 28806 20792 28858
rect 20546 28804 20552 28806
rect 20608 28804 20632 28806
rect 20688 28804 20712 28806
rect 20768 28804 20792 28806
rect 20848 28804 20854 28806
rect 20546 28795 20854 28804
rect 20546 27772 20854 27781
rect 20546 27770 20552 27772
rect 20608 27770 20632 27772
rect 20688 27770 20712 27772
rect 20768 27770 20792 27772
rect 20848 27770 20854 27772
rect 20608 27718 20610 27770
rect 20790 27718 20792 27770
rect 20546 27716 20552 27718
rect 20608 27716 20632 27718
rect 20688 27716 20712 27718
rect 20768 27716 20792 27718
rect 20848 27716 20854 27718
rect 20546 27707 20854 27716
rect 20076 27600 20128 27606
rect 20076 27542 20128 27548
rect 19984 27532 20036 27538
rect 19984 27474 20036 27480
rect 19996 24426 20024 27474
rect 20088 25498 20116 27542
rect 20904 27328 20956 27334
rect 20904 27270 20956 27276
rect 20916 27130 20944 27270
rect 20904 27124 20956 27130
rect 20904 27066 20956 27072
rect 20546 26684 20854 26693
rect 20546 26682 20552 26684
rect 20608 26682 20632 26684
rect 20688 26682 20712 26684
rect 20768 26682 20792 26684
rect 20848 26682 20854 26684
rect 20608 26630 20610 26682
rect 20790 26630 20792 26682
rect 20546 26628 20552 26630
rect 20608 26628 20632 26630
rect 20688 26628 20712 26630
rect 20768 26628 20792 26630
rect 20848 26628 20854 26630
rect 20546 26619 20854 26628
rect 20720 26240 20772 26246
rect 20720 26182 20772 26188
rect 20732 25770 20760 26182
rect 20720 25764 20772 25770
rect 20720 25706 20772 25712
rect 20546 25596 20854 25605
rect 20546 25594 20552 25596
rect 20608 25594 20632 25596
rect 20688 25594 20712 25596
rect 20768 25594 20792 25596
rect 20848 25594 20854 25596
rect 20608 25542 20610 25594
rect 20790 25542 20792 25594
rect 20546 25540 20552 25542
rect 20608 25540 20632 25542
rect 20688 25540 20712 25542
rect 20768 25540 20792 25542
rect 20848 25540 20854 25542
rect 20546 25531 20854 25540
rect 20076 25492 20128 25498
rect 20076 25434 20128 25440
rect 20536 25492 20588 25498
rect 20536 25434 20588 25440
rect 20352 25424 20404 25430
rect 20352 25366 20404 25372
rect 20076 25356 20128 25362
rect 20076 25298 20128 25304
rect 20088 24614 20116 25298
rect 20076 24608 20128 24614
rect 20076 24550 20128 24556
rect 19996 24398 20300 24426
rect 19984 24268 20036 24274
rect 19984 24210 20036 24216
rect 19720 23854 19932 23882
rect 19996 23866 20024 24210
rect 19984 23860 20036 23866
rect 19616 23656 19668 23662
rect 19616 23598 19668 23604
rect 19524 23520 19576 23526
rect 19524 23462 19576 23468
rect 19352 23174 19472 23202
rect 18972 22976 19024 22982
rect 18972 22918 19024 22924
rect 18696 22772 18748 22778
rect 18696 22714 18748 22720
rect 18984 22642 19012 22918
rect 19352 22710 19380 23174
rect 19340 22704 19392 22710
rect 19340 22646 19392 22652
rect 18236 22636 18288 22642
rect 18236 22578 18288 22584
rect 18972 22636 19024 22642
rect 18972 22578 19024 22584
rect 18248 22094 18276 22578
rect 19064 22568 19116 22574
rect 19064 22510 19116 22516
rect 19156 22568 19208 22574
rect 19156 22510 19208 22516
rect 19340 22568 19392 22574
rect 19340 22510 19392 22516
rect 19432 22568 19484 22574
rect 19432 22510 19484 22516
rect 19076 22098 19104 22510
rect 19168 22234 19196 22510
rect 19248 22500 19300 22506
rect 19248 22442 19300 22448
rect 19156 22228 19208 22234
rect 19156 22170 19208 22176
rect 18248 22066 18460 22094
rect 18052 22024 18104 22030
rect 18050 21992 18052 22001
rect 18104 21992 18106 22001
rect 18050 21927 18106 21936
rect 18328 21616 18380 21622
rect 18328 21558 18380 21564
rect 17960 21480 18012 21486
rect 17960 21422 18012 21428
rect 17868 21140 17920 21146
rect 17868 21082 17920 21088
rect 17972 20942 18000 21422
rect 18144 21412 18196 21418
rect 18144 21354 18196 21360
rect 18052 21004 18104 21010
rect 18052 20946 18104 20952
rect 17960 20936 18012 20942
rect 17960 20878 18012 20884
rect 17960 20392 18012 20398
rect 17788 20352 17960 20380
rect 17684 20334 17736 20340
rect 17960 20334 18012 20340
rect 18064 19990 18092 20946
rect 18156 20602 18184 21354
rect 18144 20596 18196 20602
rect 18144 20538 18196 20544
rect 18052 19984 18104 19990
rect 18052 19926 18104 19932
rect 17960 19712 18012 19718
rect 17960 19654 18012 19660
rect 17868 19372 17920 19378
rect 17868 19314 17920 19320
rect 17592 19304 17644 19310
rect 17592 19246 17644 19252
rect 17604 18970 17632 19246
rect 16960 18924 17080 18952
rect 17592 18964 17644 18970
rect 16856 18216 16908 18222
rect 16856 18158 16908 18164
rect 16764 18080 16816 18086
rect 16764 18022 16816 18028
rect 16776 17134 16804 18022
rect 16868 17746 16896 18158
rect 16856 17740 16908 17746
rect 16856 17682 16908 17688
rect 16960 17134 16988 18924
rect 17592 18906 17644 18912
rect 17040 18828 17092 18834
rect 17040 18770 17092 18776
rect 17052 18426 17080 18770
rect 17188 18524 17496 18533
rect 17188 18522 17194 18524
rect 17250 18522 17274 18524
rect 17330 18522 17354 18524
rect 17410 18522 17434 18524
rect 17490 18522 17496 18524
rect 17250 18470 17252 18522
rect 17432 18470 17434 18522
rect 17188 18468 17194 18470
rect 17250 18468 17274 18470
rect 17330 18468 17354 18470
rect 17410 18468 17434 18470
rect 17490 18468 17496 18470
rect 17188 18459 17496 18468
rect 17040 18420 17092 18426
rect 17040 18362 17092 18368
rect 17604 17746 17632 18906
rect 17880 18290 17908 19314
rect 17972 18902 18000 19654
rect 18064 19310 18092 19926
rect 18340 19417 18368 21558
rect 18432 21078 18460 22066
rect 19064 22092 19116 22098
rect 19064 22034 19116 22040
rect 18512 22024 18564 22030
rect 18512 21966 18564 21972
rect 18696 22024 18748 22030
rect 18696 21966 18748 21972
rect 18420 21072 18472 21078
rect 18420 21014 18472 21020
rect 18326 19408 18382 19417
rect 18326 19343 18382 19352
rect 18052 19304 18104 19310
rect 18052 19246 18104 19252
rect 18328 19304 18380 19310
rect 18328 19246 18380 19252
rect 17960 18896 18012 18902
rect 17960 18838 18012 18844
rect 18236 18624 18288 18630
rect 18236 18566 18288 18572
rect 17868 18284 17920 18290
rect 17868 18226 17920 18232
rect 18144 18080 18196 18086
rect 18144 18022 18196 18028
rect 18156 17882 18184 18022
rect 17684 17876 17736 17882
rect 17684 17818 17736 17824
rect 18144 17876 18196 17882
rect 18144 17818 18196 17824
rect 17592 17740 17644 17746
rect 17592 17682 17644 17688
rect 17188 17436 17496 17445
rect 17188 17434 17194 17436
rect 17250 17434 17274 17436
rect 17330 17434 17354 17436
rect 17410 17434 17434 17436
rect 17490 17434 17496 17436
rect 17250 17382 17252 17434
rect 17432 17382 17434 17434
rect 17188 17380 17194 17382
rect 17250 17380 17274 17382
rect 17330 17380 17354 17382
rect 17410 17380 17434 17382
rect 17490 17380 17496 17382
rect 17188 17371 17496 17380
rect 16672 17128 16724 17134
rect 16672 17070 16724 17076
rect 16764 17128 16816 17134
rect 16764 17070 16816 17076
rect 16948 17128 17000 17134
rect 16948 17070 17000 17076
rect 17132 17128 17184 17134
rect 17132 17070 17184 17076
rect 16948 16992 17000 16998
rect 16948 16934 17000 16940
rect 16856 16652 16908 16658
rect 16856 16594 16908 16600
rect 16868 14414 16896 16594
rect 16856 14408 16908 14414
rect 16856 14350 16908 14356
rect 16672 13796 16724 13802
rect 16672 13738 16724 13744
rect 16684 13326 16712 13738
rect 16672 13320 16724 13326
rect 16672 13262 16724 13268
rect 16672 12300 16724 12306
rect 16672 12242 16724 12248
rect 16580 11688 16632 11694
rect 16580 11630 16632 11636
rect 16580 11552 16632 11558
rect 16580 11494 16632 11500
rect 16592 11354 16620 11494
rect 16580 11348 16632 11354
rect 16580 11290 16632 11296
rect 16684 11150 16712 12242
rect 16960 11762 16988 16934
rect 17144 16658 17172 17070
rect 17696 16946 17724 17818
rect 18052 17808 18104 17814
rect 18052 17750 18104 17756
rect 17776 17740 17828 17746
rect 17776 17682 17828 17688
rect 17788 17338 17816 17682
rect 17960 17672 18012 17678
rect 17960 17614 18012 17620
rect 17776 17332 17828 17338
rect 17776 17274 17828 17280
rect 17972 17270 18000 17614
rect 18064 17610 18092 17750
rect 18052 17604 18104 17610
rect 18052 17546 18104 17552
rect 17960 17264 18012 17270
rect 17960 17206 18012 17212
rect 18052 17196 18104 17202
rect 18052 17138 18104 17144
rect 17604 16918 17724 16946
rect 17868 16992 17920 16998
rect 17868 16934 17920 16940
rect 17604 16658 17632 16918
rect 17880 16794 17908 16934
rect 17684 16788 17736 16794
rect 17684 16730 17736 16736
rect 17868 16788 17920 16794
rect 17868 16730 17920 16736
rect 17696 16658 17724 16730
rect 17132 16652 17184 16658
rect 17132 16594 17184 16600
rect 17592 16652 17644 16658
rect 17592 16594 17644 16600
rect 17684 16652 17736 16658
rect 17684 16594 17736 16600
rect 17188 16348 17496 16357
rect 17188 16346 17194 16348
rect 17250 16346 17274 16348
rect 17330 16346 17354 16348
rect 17410 16346 17434 16348
rect 17490 16346 17496 16348
rect 17250 16294 17252 16346
rect 17432 16294 17434 16346
rect 17188 16292 17194 16294
rect 17250 16292 17274 16294
rect 17330 16292 17354 16294
rect 17410 16292 17434 16294
rect 17490 16292 17496 16294
rect 17188 16283 17496 16292
rect 17776 16040 17828 16046
rect 17776 15982 17828 15988
rect 17684 15904 17736 15910
rect 17684 15846 17736 15852
rect 17696 15706 17724 15846
rect 17684 15700 17736 15706
rect 17684 15642 17736 15648
rect 17592 15496 17644 15502
rect 17592 15438 17644 15444
rect 17188 15260 17496 15269
rect 17188 15258 17194 15260
rect 17250 15258 17274 15260
rect 17330 15258 17354 15260
rect 17410 15258 17434 15260
rect 17490 15258 17496 15260
rect 17250 15206 17252 15258
rect 17432 15206 17434 15258
rect 17188 15204 17194 15206
rect 17250 15204 17274 15206
rect 17330 15204 17354 15206
rect 17410 15204 17434 15206
rect 17490 15204 17496 15206
rect 17188 15195 17496 15204
rect 17040 14408 17092 14414
rect 17040 14350 17092 14356
rect 17052 14074 17080 14350
rect 17188 14172 17496 14181
rect 17188 14170 17194 14172
rect 17250 14170 17274 14172
rect 17330 14170 17354 14172
rect 17410 14170 17434 14172
rect 17490 14170 17496 14172
rect 17250 14118 17252 14170
rect 17432 14118 17434 14170
rect 17188 14116 17194 14118
rect 17250 14116 17274 14118
rect 17330 14116 17354 14118
rect 17410 14116 17434 14118
rect 17490 14116 17496 14118
rect 17188 14107 17496 14116
rect 17040 14068 17092 14074
rect 17040 14010 17092 14016
rect 17316 13728 17368 13734
rect 17316 13670 17368 13676
rect 17328 13394 17356 13670
rect 17604 13394 17632 15438
rect 17788 15162 17816 15982
rect 17960 15904 18012 15910
rect 17960 15846 18012 15852
rect 17776 15156 17828 15162
rect 17776 15098 17828 15104
rect 17972 14958 18000 15846
rect 18064 15026 18092 17138
rect 18052 15020 18104 15026
rect 18052 14962 18104 14968
rect 17960 14952 18012 14958
rect 17960 14894 18012 14900
rect 18064 13938 18092 14962
rect 18248 14822 18276 18566
rect 18340 17678 18368 19246
rect 18328 17672 18380 17678
rect 18328 17614 18380 17620
rect 18432 17542 18460 21014
rect 18524 21010 18552 21966
rect 18512 21004 18564 21010
rect 18512 20946 18564 20952
rect 18708 20806 18736 21966
rect 19076 21622 19104 22034
rect 19260 22030 19288 22442
rect 19248 22024 19300 22030
rect 19248 21966 19300 21972
rect 19156 21956 19208 21962
rect 19156 21898 19208 21904
rect 19064 21616 19116 21622
rect 19064 21558 19116 21564
rect 19168 21554 19196 21898
rect 19156 21548 19208 21554
rect 19156 21490 19208 21496
rect 19260 21146 19288 21966
rect 19352 21690 19380 22510
rect 19340 21684 19392 21690
rect 19340 21626 19392 21632
rect 19352 21486 19380 21626
rect 19340 21480 19392 21486
rect 19340 21422 19392 21428
rect 19248 21140 19300 21146
rect 19248 21082 19300 21088
rect 19156 21004 19208 21010
rect 19156 20946 19208 20952
rect 18696 20800 18748 20806
rect 18696 20742 18748 20748
rect 18512 20392 18564 20398
rect 18512 20334 18564 20340
rect 18972 20392 19024 20398
rect 18972 20334 19024 20340
rect 18524 19825 18552 20334
rect 18984 20058 19012 20334
rect 18972 20052 19024 20058
rect 18972 19994 19024 20000
rect 18510 19816 18566 19825
rect 18510 19751 18566 19760
rect 18524 18222 18552 19751
rect 18604 19712 18656 19718
rect 18604 19654 18656 19660
rect 18616 19446 18644 19654
rect 18604 19440 18656 19446
rect 18604 19382 18656 19388
rect 18696 18624 18748 18630
rect 18696 18566 18748 18572
rect 18512 18216 18564 18222
rect 18512 18158 18564 18164
rect 18420 17536 18472 17542
rect 18420 17478 18472 17484
rect 18328 16040 18380 16046
rect 18328 15982 18380 15988
rect 18420 16040 18472 16046
rect 18420 15982 18472 15988
rect 18340 15706 18368 15982
rect 18328 15700 18380 15706
rect 18328 15642 18380 15648
rect 18432 14890 18460 15982
rect 18524 14940 18552 18158
rect 18708 18086 18736 18566
rect 18696 18080 18748 18086
rect 18696 18022 18748 18028
rect 18708 17746 18736 18022
rect 18696 17740 18748 17746
rect 18696 17682 18748 17688
rect 19064 17740 19116 17746
rect 19064 17682 19116 17688
rect 18880 17128 18932 17134
rect 18880 17070 18932 17076
rect 18892 16794 18920 17070
rect 18972 17060 19024 17066
rect 18972 17002 19024 17008
rect 18984 16794 19012 17002
rect 19076 16794 19104 17682
rect 18880 16788 18932 16794
rect 18880 16730 18932 16736
rect 18972 16788 19024 16794
rect 18972 16730 19024 16736
rect 19064 16788 19116 16794
rect 19064 16730 19116 16736
rect 18788 15972 18840 15978
rect 18788 15914 18840 15920
rect 18800 15638 18828 15914
rect 18788 15632 18840 15638
rect 18788 15574 18840 15580
rect 18524 14912 18644 14940
rect 18420 14884 18472 14890
rect 18472 14844 18552 14872
rect 18420 14826 18472 14832
rect 18236 14816 18288 14822
rect 18236 14758 18288 14764
rect 18328 14816 18380 14822
rect 18328 14758 18380 14764
rect 18144 14408 18196 14414
rect 18144 14350 18196 14356
rect 18052 13932 18104 13938
rect 18052 13874 18104 13880
rect 17776 13864 17828 13870
rect 17776 13806 17828 13812
rect 17316 13388 17368 13394
rect 17316 13330 17368 13336
rect 17592 13388 17644 13394
rect 17592 13330 17644 13336
rect 17188 13084 17496 13093
rect 17188 13082 17194 13084
rect 17250 13082 17274 13084
rect 17330 13082 17354 13084
rect 17410 13082 17434 13084
rect 17490 13082 17496 13084
rect 17250 13030 17252 13082
rect 17432 13030 17434 13082
rect 17188 13028 17194 13030
rect 17250 13028 17274 13030
rect 17330 13028 17354 13030
rect 17410 13028 17434 13030
rect 17490 13028 17496 13030
rect 17188 13019 17496 13028
rect 17788 12434 17816 13806
rect 17868 13728 17920 13734
rect 17868 13670 17920 13676
rect 17880 12986 17908 13670
rect 17868 12980 17920 12986
rect 17868 12922 17920 12928
rect 17788 12406 17908 12434
rect 17684 12096 17736 12102
rect 17684 12038 17736 12044
rect 17188 11996 17496 12005
rect 17188 11994 17194 11996
rect 17250 11994 17274 11996
rect 17330 11994 17354 11996
rect 17410 11994 17434 11996
rect 17490 11994 17496 11996
rect 17250 11942 17252 11994
rect 17432 11942 17434 11994
rect 17188 11940 17194 11942
rect 17250 11940 17274 11942
rect 17330 11940 17354 11942
rect 17410 11940 17434 11942
rect 17490 11940 17496 11942
rect 17188 11931 17496 11940
rect 17696 11762 17724 12038
rect 16948 11756 17000 11762
rect 16948 11698 17000 11704
rect 17684 11756 17736 11762
rect 17684 11698 17736 11704
rect 17408 11552 17460 11558
rect 17408 11494 17460 11500
rect 17420 11354 17448 11494
rect 17408 11348 17460 11354
rect 17408 11290 17460 11296
rect 16672 11144 16724 11150
rect 16672 11086 16724 11092
rect 16028 10600 16080 10606
rect 16028 10542 16080 10548
rect 16040 10266 16068 10542
rect 15936 10260 15988 10266
rect 15936 10202 15988 10208
rect 16028 10260 16080 10266
rect 16028 10202 16080 10208
rect 15948 10062 15976 10202
rect 16580 10192 16632 10198
rect 16580 10134 16632 10140
rect 15752 10056 15804 10062
rect 15752 9998 15804 10004
rect 15936 10056 15988 10062
rect 15936 9998 15988 10004
rect 15764 9586 15792 9998
rect 15752 9580 15804 9586
rect 15752 9522 15804 9528
rect 15844 9376 15896 9382
rect 15844 9318 15896 9324
rect 15856 9178 15884 9318
rect 16592 9178 16620 10134
rect 16684 9518 16712 11086
rect 17188 10908 17496 10917
rect 17188 10906 17194 10908
rect 17250 10906 17274 10908
rect 17330 10906 17354 10908
rect 17410 10906 17434 10908
rect 17490 10906 17496 10908
rect 17250 10854 17252 10906
rect 17432 10854 17434 10906
rect 17188 10852 17194 10854
rect 17250 10852 17274 10854
rect 17330 10852 17354 10854
rect 17410 10852 17434 10854
rect 17490 10852 17496 10854
rect 17188 10843 17496 10852
rect 16764 10464 16816 10470
rect 16764 10406 16816 10412
rect 16672 9512 16724 9518
rect 16672 9454 16724 9460
rect 16776 9450 16804 10406
rect 17696 9994 17724 11698
rect 17776 10124 17828 10130
rect 17776 10066 17828 10072
rect 17684 9988 17736 9994
rect 17684 9930 17736 9936
rect 17592 9920 17644 9926
rect 17592 9862 17644 9868
rect 17188 9820 17496 9829
rect 17188 9818 17194 9820
rect 17250 9818 17274 9820
rect 17330 9818 17354 9820
rect 17410 9818 17434 9820
rect 17490 9818 17496 9820
rect 17250 9766 17252 9818
rect 17432 9766 17434 9818
rect 17188 9764 17194 9766
rect 17250 9764 17274 9766
rect 17330 9764 17354 9766
rect 17410 9764 17434 9766
rect 17490 9764 17496 9766
rect 17188 9755 17496 9764
rect 17604 9518 17632 9862
rect 17788 9722 17816 10066
rect 17776 9716 17828 9722
rect 17776 9658 17828 9664
rect 17684 9648 17736 9654
rect 17880 9602 17908 12406
rect 17960 12300 18012 12306
rect 17960 12242 18012 12248
rect 17972 11898 18000 12242
rect 17960 11892 18012 11898
rect 17960 11834 18012 11840
rect 18156 10742 18184 14350
rect 18248 12782 18276 14758
rect 18340 14385 18368 14758
rect 18420 14476 18472 14482
rect 18420 14418 18472 14424
rect 18326 14376 18382 14385
rect 18326 14311 18382 14320
rect 18432 13530 18460 14418
rect 18420 13524 18472 13530
rect 18420 13466 18472 13472
rect 18432 12782 18460 13466
rect 18524 12850 18552 14844
rect 18616 14482 18644 14912
rect 18604 14476 18656 14482
rect 18604 14418 18656 14424
rect 18880 14476 18932 14482
rect 18880 14418 18932 14424
rect 18616 13938 18644 14418
rect 18696 14408 18748 14414
rect 18696 14350 18748 14356
rect 18604 13932 18656 13938
rect 18604 13874 18656 13880
rect 18512 12844 18564 12850
rect 18512 12786 18564 12792
rect 18236 12776 18288 12782
rect 18236 12718 18288 12724
rect 18420 12776 18472 12782
rect 18420 12718 18472 12724
rect 18708 11694 18736 14350
rect 18892 13530 18920 14418
rect 18880 13524 18932 13530
rect 18880 13466 18932 13472
rect 18788 12912 18840 12918
rect 18788 12854 18840 12860
rect 18800 12714 18828 12854
rect 18892 12850 18920 13466
rect 19168 12918 19196 20946
rect 19340 20800 19392 20806
rect 19340 20742 19392 20748
rect 19352 20330 19380 20742
rect 19340 20324 19392 20330
rect 19340 20266 19392 20272
rect 19444 20210 19472 22510
rect 19628 22234 19656 23598
rect 19616 22228 19668 22234
rect 19616 22170 19668 22176
rect 19616 21004 19668 21010
rect 19616 20946 19668 20952
rect 19352 20182 19472 20210
rect 19524 20256 19576 20262
rect 19524 20198 19576 20204
rect 19352 20058 19380 20182
rect 19536 20058 19564 20198
rect 19628 20058 19656 20946
rect 19340 20052 19392 20058
rect 19340 19994 19392 20000
rect 19524 20052 19576 20058
rect 19524 19994 19576 20000
rect 19616 20052 19668 20058
rect 19616 19994 19668 20000
rect 19352 19514 19380 19994
rect 19616 19848 19668 19854
rect 19616 19790 19668 19796
rect 19340 19508 19392 19514
rect 19340 19450 19392 19456
rect 19352 18902 19380 19450
rect 19628 19378 19656 19790
rect 19616 19372 19668 19378
rect 19616 19314 19668 19320
rect 19340 18896 19392 18902
rect 19392 18856 19472 18884
rect 19340 18838 19392 18844
rect 19444 18290 19472 18856
rect 19628 18408 19656 19314
rect 19720 19310 19748 23854
rect 19984 23802 20036 23808
rect 19800 23520 19852 23526
rect 19800 23462 19852 23468
rect 19812 19922 19840 23462
rect 19892 22500 19944 22506
rect 19892 22442 19944 22448
rect 19904 22234 19932 22442
rect 19892 22228 19944 22234
rect 19892 22170 19944 22176
rect 19892 22092 19944 22098
rect 19892 22034 19944 22040
rect 19904 21690 19932 22034
rect 19984 21956 20036 21962
rect 19984 21898 20036 21904
rect 19892 21684 19944 21690
rect 19892 21626 19944 21632
rect 19996 20602 20024 21898
rect 20272 20942 20300 24398
rect 20364 23866 20392 25366
rect 20444 25152 20496 25158
rect 20444 25094 20496 25100
rect 20456 24750 20484 25094
rect 20444 24744 20496 24750
rect 20444 24686 20496 24692
rect 20548 24596 20576 25434
rect 20904 25356 20956 25362
rect 20904 25298 20956 25304
rect 20456 24568 20576 24596
rect 20352 23860 20404 23866
rect 20352 23802 20404 23808
rect 20456 23662 20484 24568
rect 20546 24508 20854 24517
rect 20546 24506 20552 24508
rect 20608 24506 20632 24508
rect 20688 24506 20712 24508
rect 20768 24506 20792 24508
rect 20848 24506 20854 24508
rect 20608 24454 20610 24506
rect 20790 24454 20792 24506
rect 20546 24452 20552 24454
rect 20608 24452 20632 24454
rect 20688 24452 20712 24454
rect 20768 24452 20792 24454
rect 20848 24452 20854 24454
rect 20546 24443 20854 24452
rect 20444 23656 20496 23662
rect 20444 23598 20496 23604
rect 20352 23112 20404 23118
rect 20352 23054 20404 23060
rect 20364 22234 20392 23054
rect 20456 22778 20484 23598
rect 20546 23420 20854 23429
rect 20546 23418 20552 23420
rect 20608 23418 20632 23420
rect 20688 23418 20712 23420
rect 20768 23418 20792 23420
rect 20848 23418 20854 23420
rect 20608 23366 20610 23418
rect 20790 23366 20792 23418
rect 20546 23364 20552 23366
rect 20608 23364 20632 23366
rect 20688 23364 20712 23366
rect 20768 23364 20792 23366
rect 20848 23364 20854 23366
rect 20546 23355 20854 23364
rect 20444 22772 20496 22778
rect 20444 22714 20496 22720
rect 20546 22332 20854 22341
rect 20546 22330 20552 22332
rect 20608 22330 20632 22332
rect 20688 22330 20712 22332
rect 20768 22330 20792 22332
rect 20848 22330 20854 22332
rect 20608 22278 20610 22330
rect 20790 22278 20792 22330
rect 20546 22276 20552 22278
rect 20608 22276 20632 22278
rect 20688 22276 20712 22278
rect 20768 22276 20792 22278
rect 20848 22276 20854 22278
rect 20546 22267 20854 22276
rect 20352 22228 20404 22234
rect 20352 22170 20404 22176
rect 20364 21350 20392 22170
rect 20916 21962 20944 25298
rect 20904 21956 20956 21962
rect 20904 21898 20956 21904
rect 20352 21344 20404 21350
rect 20352 21286 20404 21292
rect 20444 21344 20496 21350
rect 20444 21286 20496 21292
rect 20456 21078 20484 21286
rect 20546 21244 20854 21253
rect 20546 21242 20552 21244
rect 20608 21242 20632 21244
rect 20688 21242 20712 21244
rect 20768 21242 20792 21244
rect 20848 21242 20854 21244
rect 20608 21190 20610 21242
rect 20790 21190 20792 21242
rect 20546 21188 20552 21190
rect 20608 21188 20632 21190
rect 20688 21188 20712 21190
rect 20768 21188 20792 21190
rect 20848 21188 20854 21190
rect 20546 21179 20854 21188
rect 21008 21162 21036 29990
rect 21100 22094 21128 30874
rect 22020 30802 22048 31600
rect 22744 31136 22796 31142
rect 22744 31078 22796 31084
rect 22756 30802 22784 31078
rect 23492 30938 23520 31600
rect 23480 30932 23532 30938
rect 23480 30874 23532 30880
rect 22008 30796 22060 30802
rect 22008 30738 22060 30744
rect 22744 30796 22796 30802
rect 22744 30738 22796 30744
rect 21732 30728 21784 30734
rect 21732 30670 21784 30676
rect 22468 30728 22520 30734
rect 22468 30670 22520 30676
rect 21364 30592 21416 30598
rect 21364 30534 21416 30540
rect 21272 30252 21324 30258
rect 21272 30194 21324 30200
rect 21180 29096 21232 29102
rect 21180 29038 21232 29044
rect 21192 28422 21220 29038
rect 21284 28626 21312 30194
rect 21272 28620 21324 28626
rect 21272 28562 21324 28568
rect 21180 28416 21232 28422
rect 21180 28358 21232 28364
rect 21284 28082 21312 28562
rect 21272 28076 21324 28082
rect 21272 28018 21324 28024
rect 21272 27056 21324 27062
rect 21270 27024 21272 27033
rect 21324 27024 21326 27033
rect 21270 26959 21326 26968
rect 21272 26920 21324 26926
rect 21272 26862 21324 26868
rect 21284 26586 21312 26862
rect 21272 26580 21324 26586
rect 21272 26522 21324 26528
rect 21376 24698 21404 30534
rect 21548 29776 21600 29782
rect 21548 29718 21600 29724
rect 21560 29238 21588 29718
rect 21744 29510 21772 30670
rect 22480 30394 22508 30670
rect 22468 30388 22520 30394
rect 22468 30330 22520 30336
rect 22652 30388 22704 30394
rect 22652 30330 22704 30336
rect 22664 30190 22692 30330
rect 22756 30258 22784 30738
rect 23204 30728 23256 30734
rect 23204 30670 23256 30676
rect 23020 30592 23072 30598
rect 23020 30534 23072 30540
rect 23112 30592 23164 30598
rect 23112 30534 23164 30540
rect 23032 30258 23060 30534
rect 22744 30252 22796 30258
rect 22744 30194 22796 30200
rect 23020 30252 23072 30258
rect 23020 30194 23072 30200
rect 22652 30184 22704 30190
rect 22652 30126 22704 30132
rect 23020 30116 23072 30122
rect 23020 30058 23072 30064
rect 22834 29744 22890 29753
rect 22834 29679 22890 29688
rect 22928 29708 22980 29714
rect 22652 29640 22704 29646
rect 22652 29582 22704 29588
rect 21732 29504 21784 29510
rect 21732 29446 21784 29452
rect 21548 29232 21600 29238
rect 21548 29174 21600 29180
rect 21560 28098 21588 29174
rect 21640 29096 21692 29102
rect 21640 29038 21692 29044
rect 21652 28218 21680 29038
rect 21732 28960 21784 28966
rect 21732 28902 21784 28908
rect 21744 28694 21772 28902
rect 21732 28688 21784 28694
rect 21732 28630 21784 28636
rect 22008 28416 22060 28422
rect 22008 28358 22060 28364
rect 21640 28212 21692 28218
rect 21640 28154 21692 28160
rect 21560 28070 21680 28098
rect 21548 27668 21600 27674
rect 21548 27610 21600 27616
rect 21456 27124 21508 27130
rect 21456 27066 21508 27072
rect 21468 26382 21496 27066
rect 21560 26994 21588 27610
rect 21548 26988 21600 26994
rect 21548 26930 21600 26936
rect 21548 26852 21600 26858
rect 21548 26794 21600 26800
rect 21560 26625 21588 26794
rect 21546 26616 21602 26625
rect 21546 26551 21602 26560
rect 21548 26512 21600 26518
rect 21548 26454 21600 26460
rect 21456 26376 21508 26382
rect 21456 26318 21508 26324
rect 21468 24954 21496 26318
rect 21560 26042 21588 26454
rect 21652 26058 21680 28070
rect 21824 27872 21876 27878
rect 21824 27814 21876 27820
rect 21836 27606 21864 27814
rect 21824 27600 21876 27606
rect 21824 27542 21876 27548
rect 22020 27554 22048 28358
rect 22664 28218 22692 29582
rect 22848 29510 22876 29679
rect 22928 29650 22980 29656
rect 22940 29617 22968 29650
rect 22926 29608 22982 29617
rect 22926 29543 22982 29552
rect 22836 29504 22888 29510
rect 22836 29446 22888 29452
rect 23032 29306 23060 30058
rect 23124 29646 23152 30534
rect 23216 30122 23244 30670
rect 23572 30592 23624 30598
rect 23572 30534 23624 30540
rect 23204 30116 23256 30122
rect 23204 30058 23256 30064
rect 23480 30116 23532 30122
rect 23480 30058 23532 30064
rect 23492 29866 23520 30058
rect 23400 29838 23520 29866
rect 23400 29714 23428 29838
rect 23584 29730 23612 30534
rect 23904 30492 24212 30501
rect 23904 30490 23910 30492
rect 23966 30490 23990 30492
rect 24046 30490 24070 30492
rect 24126 30490 24150 30492
rect 24206 30490 24212 30492
rect 23966 30438 23968 30490
rect 24148 30438 24150 30490
rect 23904 30436 23910 30438
rect 23966 30436 23990 30438
rect 24046 30436 24070 30438
rect 24126 30436 24150 30438
rect 24206 30436 24212 30438
rect 23904 30427 24212 30436
rect 23846 30152 23902 30161
rect 23846 30087 23902 30096
rect 24400 30116 24452 30122
rect 23664 30048 23716 30054
rect 23664 29990 23716 29996
rect 23388 29708 23440 29714
rect 23388 29650 23440 29656
rect 23492 29702 23612 29730
rect 23112 29640 23164 29646
rect 23112 29582 23164 29588
rect 23296 29504 23348 29510
rect 23296 29446 23348 29452
rect 23020 29300 23072 29306
rect 23020 29242 23072 29248
rect 23308 29102 23336 29446
rect 23296 29096 23348 29102
rect 23296 29038 23348 29044
rect 23112 28620 23164 28626
rect 23112 28562 23164 28568
rect 22836 28416 22888 28422
rect 22836 28358 22888 28364
rect 22928 28416 22980 28422
rect 22928 28358 22980 28364
rect 22192 28212 22244 28218
rect 22192 28154 22244 28160
rect 22652 28212 22704 28218
rect 22652 28154 22704 28160
rect 22204 27878 22232 28154
rect 22376 28008 22428 28014
rect 22376 27950 22428 27956
rect 22192 27872 22244 27878
rect 22192 27814 22244 27820
rect 22020 27538 22324 27554
rect 21732 27532 21784 27538
rect 22020 27532 22336 27538
rect 22020 27526 22284 27532
rect 21732 27474 21784 27480
rect 22284 27474 22336 27480
rect 21744 26586 21772 27474
rect 22284 27396 22336 27402
rect 22284 27338 22336 27344
rect 22192 27328 22244 27334
rect 22192 27270 22244 27276
rect 21916 27124 21968 27130
rect 21916 27066 21968 27072
rect 21928 26976 21956 27066
rect 22204 26994 22232 27270
rect 21836 26948 21956 26976
rect 22192 26988 22244 26994
rect 21836 26858 21864 26948
rect 22192 26930 22244 26936
rect 21824 26852 21876 26858
rect 21824 26794 21876 26800
rect 22100 26784 22152 26790
rect 22020 26744 22100 26772
rect 21822 26616 21878 26625
rect 21732 26580 21784 26586
rect 21822 26551 21878 26560
rect 21732 26522 21784 26528
rect 21836 26500 21864 26551
rect 21916 26512 21968 26518
rect 21836 26472 21916 26500
rect 21548 26036 21600 26042
rect 21652 26030 21772 26058
rect 21548 25978 21600 25984
rect 21640 25696 21692 25702
rect 21640 25638 21692 25644
rect 21456 24948 21508 24954
rect 21456 24890 21508 24896
rect 21376 24670 21588 24698
rect 21652 24682 21680 25638
rect 21272 24064 21324 24070
rect 21272 24006 21324 24012
rect 21284 23866 21312 24006
rect 21272 23860 21324 23866
rect 21272 23802 21324 23808
rect 21364 22500 21416 22506
rect 21364 22442 21416 22448
rect 21456 22500 21508 22506
rect 21456 22442 21508 22448
rect 21376 22386 21404 22442
rect 21284 22358 21404 22386
rect 21100 22066 21220 22094
rect 21088 21888 21140 21894
rect 21088 21830 21140 21836
rect 20916 21134 21036 21162
rect 20444 21072 20496 21078
rect 20444 21014 20496 21020
rect 20260 20936 20312 20942
rect 20916 20890 20944 21134
rect 20996 21004 21048 21010
rect 20996 20946 21048 20952
rect 20260 20878 20312 20884
rect 20824 20862 20944 20890
rect 19984 20596 20036 20602
rect 19984 20538 20036 20544
rect 19800 19916 19852 19922
rect 19800 19858 19852 19864
rect 19996 19802 20024 20538
rect 20824 20534 20852 20862
rect 20904 20800 20956 20806
rect 20904 20742 20956 20748
rect 20812 20528 20864 20534
rect 20812 20470 20864 20476
rect 20916 20398 20944 20742
rect 20812 20392 20864 20398
rect 20812 20334 20864 20340
rect 20904 20392 20956 20398
rect 20904 20334 20956 20340
rect 20824 20244 20852 20334
rect 20824 20216 20944 20244
rect 20546 20156 20854 20165
rect 20546 20154 20552 20156
rect 20608 20154 20632 20156
rect 20688 20154 20712 20156
rect 20768 20154 20792 20156
rect 20848 20154 20854 20156
rect 20608 20102 20610 20154
rect 20790 20102 20792 20154
rect 20546 20100 20552 20102
rect 20608 20100 20632 20102
rect 20688 20100 20712 20102
rect 20768 20100 20792 20102
rect 20848 20100 20854 20102
rect 20546 20091 20854 20100
rect 20916 19922 20944 20216
rect 21008 20058 21036 20946
rect 20996 20052 21048 20058
rect 20996 19994 21048 20000
rect 20076 19916 20128 19922
rect 20076 19858 20128 19864
rect 20168 19916 20220 19922
rect 20168 19858 20220 19864
rect 20904 19916 20956 19922
rect 20904 19858 20956 19864
rect 19812 19774 20024 19802
rect 19708 19304 19760 19310
rect 19708 19246 19760 19252
rect 19720 18630 19748 19246
rect 19708 18624 19760 18630
rect 19708 18566 19760 18572
rect 19708 18420 19760 18426
rect 19628 18380 19708 18408
rect 19708 18362 19760 18368
rect 19432 18284 19484 18290
rect 19432 18226 19484 18232
rect 19248 17536 19300 17542
rect 19248 17478 19300 17484
rect 19260 17066 19288 17478
rect 19444 17134 19472 18226
rect 19616 17536 19668 17542
rect 19616 17478 19668 17484
rect 19432 17128 19484 17134
rect 19432 17070 19484 17076
rect 19248 17060 19300 17066
rect 19248 17002 19300 17008
rect 19628 16794 19656 17478
rect 19616 16788 19668 16794
rect 19616 16730 19668 16736
rect 19432 16652 19484 16658
rect 19432 16594 19484 16600
rect 19444 15502 19472 16594
rect 19720 16590 19748 18362
rect 19708 16584 19760 16590
rect 19708 16526 19760 16532
rect 19708 16244 19760 16250
rect 19708 16186 19760 16192
rect 19616 15564 19668 15570
rect 19616 15506 19668 15512
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 19340 15428 19392 15434
rect 19340 15370 19392 15376
rect 19248 14884 19300 14890
rect 19248 14826 19300 14832
rect 19260 14618 19288 14826
rect 19248 14612 19300 14618
rect 19248 14554 19300 14560
rect 19156 12912 19208 12918
rect 19156 12854 19208 12860
rect 18880 12844 18932 12850
rect 18880 12786 18932 12792
rect 18788 12708 18840 12714
rect 18788 12650 18840 12656
rect 19064 12096 19116 12102
rect 19064 12038 19116 12044
rect 19156 12096 19208 12102
rect 19156 12038 19208 12044
rect 19076 11762 19104 12038
rect 19168 11830 19196 12038
rect 19156 11824 19208 11830
rect 19156 11766 19208 11772
rect 19064 11756 19116 11762
rect 19064 11698 19116 11704
rect 18236 11688 18288 11694
rect 18236 11630 18288 11636
rect 18696 11688 18748 11694
rect 18696 11630 18748 11636
rect 18248 11150 18276 11630
rect 18420 11212 18472 11218
rect 18420 11154 18472 11160
rect 18236 11144 18288 11150
rect 18236 11086 18288 11092
rect 18144 10736 18196 10742
rect 18144 10678 18196 10684
rect 17736 9596 17908 9602
rect 17684 9590 17908 9596
rect 17696 9574 17908 9590
rect 17132 9512 17184 9518
rect 17132 9454 17184 9460
rect 17592 9512 17644 9518
rect 17592 9454 17644 9460
rect 18052 9512 18104 9518
rect 18052 9454 18104 9460
rect 18144 9512 18196 9518
rect 18248 9500 18276 11086
rect 18432 10606 18460 11154
rect 19076 10606 19104 11698
rect 19248 11552 19300 11558
rect 19248 11494 19300 11500
rect 19260 11286 19288 11494
rect 19248 11280 19300 11286
rect 19248 11222 19300 11228
rect 19260 10606 19288 11222
rect 18420 10600 18472 10606
rect 18420 10542 18472 10548
rect 19064 10600 19116 10606
rect 19064 10542 19116 10548
rect 19248 10600 19300 10606
rect 19248 10542 19300 10548
rect 18604 10532 18656 10538
rect 18604 10474 18656 10480
rect 18616 10130 18644 10474
rect 18788 10464 18840 10470
rect 18788 10406 18840 10412
rect 18880 10464 18932 10470
rect 18880 10406 18932 10412
rect 18800 10266 18828 10406
rect 18788 10260 18840 10266
rect 18788 10202 18840 10208
rect 18604 10124 18656 10130
rect 18604 10066 18656 10072
rect 18196 9472 18276 9500
rect 18144 9454 18196 9460
rect 16764 9444 16816 9450
rect 16764 9386 16816 9392
rect 15844 9172 15896 9178
rect 15844 9114 15896 9120
rect 16580 9172 16632 9178
rect 16580 9114 16632 9120
rect 15476 9036 15528 9042
rect 15476 8978 15528 8984
rect 15660 9036 15712 9042
rect 15660 8978 15712 8984
rect 15384 8968 15436 8974
rect 15384 8910 15436 8916
rect 17040 8968 17092 8974
rect 17144 8956 17172 9454
rect 17408 9376 17460 9382
rect 17408 9318 17460 9324
rect 17420 9110 17448 9318
rect 18064 9178 18092 9454
rect 18052 9172 18104 9178
rect 18052 9114 18104 9120
rect 17408 9104 17460 9110
rect 17408 9046 17460 9052
rect 17092 8928 17172 8956
rect 17040 8910 17092 8916
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 15016 8288 15068 8294
rect 15016 8230 15068 8236
rect 14384 6718 14504 6746
rect 14372 6656 14424 6662
rect 14372 6598 14424 6604
rect 14384 6497 14412 6598
rect 14370 6488 14426 6497
rect 14370 6423 14372 6432
rect 14424 6423 14426 6432
rect 14372 6394 14424 6400
rect 14476 6338 14504 6718
rect 14384 6310 14504 6338
rect 14568 6718 14688 6746
rect 14752 8044 14872 8072
rect 14924 8084 14976 8090
rect 14280 6112 14332 6118
rect 14280 6054 14332 6060
rect 14188 5908 14240 5914
rect 14188 5850 14240 5856
rect 13544 5840 13596 5846
rect 13544 5782 13596 5788
rect 13728 5840 13780 5846
rect 13728 5782 13780 5788
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 12808 4616 12860 4622
rect 12860 4576 12940 4604
rect 12808 4558 12860 4564
rect 12808 4480 12860 4486
rect 12808 4422 12860 4428
rect 12820 3738 12848 4422
rect 12808 3732 12860 3738
rect 12808 3674 12860 3680
rect 12532 3596 12584 3602
rect 12532 3538 12584 3544
rect 12348 2984 12400 2990
rect 12348 2926 12400 2932
rect 12176 2746 12296 2774
rect 12176 2514 12204 2746
rect 12544 2514 12572 3538
rect 12820 3534 12848 3674
rect 12808 3528 12860 3534
rect 12808 3470 12860 3476
rect 12912 3126 12940 4576
rect 13096 4554 13124 5102
rect 13452 4684 13504 4690
rect 13452 4626 13504 4632
rect 13084 4548 13136 4554
rect 13084 4490 13136 4496
rect 13096 4282 13124 4490
rect 13176 4480 13228 4486
rect 13176 4422 13228 4428
rect 13084 4276 13136 4282
rect 13084 4218 13136 4224
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 13004 3738 13032 3878
rect 13096 3754 13124 4218
rect 13188 4010 13216 4422
rect 13464 4078 13492 4626
rect 13360 4072 13412 4078
rect 13360 4014 13412 4020
rect 13452 4072 13504 4078
rect 13452 4014 13504 4020
rect 13176 4004 13228 4010
rect 13176 3946 13228 3952
rect 12992 3732 13044 3738
rect 13096 3726 13216 3754
rect 12992 3674 13044 3680
rect 13188 3602 13216 3726
rect 13268 3664 13320 3670
rect 13268 3606 13320 3612
rect 13176 3596 13228 3602
rect 13176 3538 13228 3544
rect 12900 3120 12952 3126
rect 12900 3062 12952 3068
rect 12912 2990 12940 3062
rect 13280 3058 13308 3606
rect 13372 3602 13400 4014
rect 13556 3670 13584 5782
rect 14188 5568 14240 5574
rect 14188 5510 14240 5516
rect 14200 5234 14228 5510
rect 14188 5228 14240 5234
rect 14188 5170 14240 5176
rect 13830 4924 14138 4933
rect 13830 4922 13836 4924
rect 13892 4922 13916 4924
rect 13972 4922 13996 4924
rect 14052 4922 14076 4924
rect 14132 4922 14138 4924
rect 13892 4870 13894 4922
rect 14074 4870 14076 4922
rect 13830 4868 13836 4870
rect 13892 4868 13916 4870
rect 13972 4868 13996 4870
rect 14052 4868 14076 4870
rect 14132 4868 14138 4870
rect 13830 4859 14138 4868
rect 14188 4684 14240 4690
rect 14188 4626 14240 4632
rect 13636 3936 13688 3942
rect 13636 3878 13688 3884
rect 13544 3664 13596 3670
rect 13544 3606 13596 3612
rect 13360 3596 13412 3602
rect 13360 3538 13412 3544
rect 13268 3052 13320 3058
rect 13268 2994 13320 3000
rect 13556 2990 13584 3606
rect 12900 2984 12952 2990
rect 12900 2926 12952 2932
rect 13544 2984 13596 2990
rect 13544 2926 13596 2932
rect 12716 2848 12768 2854
rect 12900 2848 12952 2854
rect 12716 2790 12768 2796
rect 12820 2808 12900 2836
rect 12728 2650 12756 2790
rect 12716 2644 12768 2650
rect 12716 2586 12768 2592
rect 11428 2508 11480 2514
rect 11428 2450 11480 2456
rect 11888 2508 11940 2514
rect 11888 2450 11940 2456
rect 12164 2508 12216 2514
rect 12164 2450 12216 2456
rect 12532 2508 12584 2514
rect 12532 2450 12584 2456
rect 12716 2508 12768 2514
rect 12820 2496 12848 2808
rect 12900 2790 12952 2796
rect 12900 2644 12952 2650
rect 12900 2586 12952 2592
rect 12912 2514 12940 2586
rect 13648 2514 13676 3878
rect 13830 3836 14138 3845
rect 13830 3834 13836 3836
rect 13892 3834 13916 3836
rect 13972 3834 13996 3836
rect 14052 3834 14076 3836
rect 14132 3834 14138 3836
rect 13892 3782 13894 3834
rect 14074 3782 14076 3834
rect 13830 3780 13836 3782
rect 13892 3780 13916 3782
rect 13972 3780 13996 3782
rect 14052 3780 14076 3782
rect 14132 3780 14138 3782
rect 13830 3771 14138 3780
rect 13728 3732 13780 3738
rect 13728 3674 13780 3680
rect 13740 2990 13768 3674
rect 13912 3528 13964 3534
rect 13832 3488 13912 3516
rect 13832 3369 13860 3488
rect 13912 3470 13964 3476
rect 13818 3360 13874 3369
rect 13818 3295 13874 3304
rect 13832 3194 13860 3295
rect 14200 3194 14228 4626
rect 14280 4480 14332 4486
rect 14280 4422 14332 4428
rect 14292 3534 14320 4422
rect 14384 4049 14412 6310
rect 14464 6112 14516 6118
rect 14464 6054 14516 6060
rect 14476 5642 14504 6054
rect 14464 5636 14516 5642
rect 14464 5578 14516 5584
rect 14464 5160 14516 5166
rect 14464 5102 14516 5108
rect 14476 4826 14504 5102
rect 14464 4820 14516 4826
rect 14464 4762 14516 4768
rect 14370 4040 14426 4049
rect 14370 3975 14426 3984
rect 14568 3720 14596 6718
rect 14648 6656 14700 6662
rect 14648 6598 14700 6604
rect 14660 6458 14688 6598
rect 14648 6452 14700 6458
rect 14648 6394 14700 6400
rect 14752 4808 14780 8044
rect 14924 8026 14976 8032
rect 15120 7954 15148 8774
rect 16856 8560 16908 8566
rect 16856 8502 16908 8508
rect 16212 8424 16264 8430
rect 16212 8366 16264 8372
rect 14832 7948 14884 7954
rect 15108 7948 15160 7954
rect 14884 7908 14964 7936
rect 14832 7890 14884 7896
rect 14936 6338 14964 7908
rect 15108 7890 15160 7896
rect 15200 7948 15252 7954
rect 15200 7890 15252 7896
rect 15016 7812 15068 7818
rect 15016 7754 15068 7760
rect 15028 6458 15056 7754
rect 15212 7750 15240 7890
rect 15384 7880 15436 7886
rect 15384 7822 15436 7828
rect 15200 7744 15252 7750
rect 15200 7686 15252 7692
rect 15108 6792 15160 6798
rect 15108 6734 15160 6740
rect 15016 6452 15068 6458
rect 15016 6394 15068 6400
rect 14936 6310 15056 6338
rect 15028 6254 15056 6310
rect 15016 6248 15068 6254
rect 15120 6225 15148 6734
rect 15212 6730 15240 7686
rect 15396 7002 15424 7822
rect 15752 7744 15804 7750
rect 15752 7686 15804 7692
rect 15764 7546 15792 7686
rect 16224 7546 16252 8366
rect 16868 8022 16896 8502
rect 17052 8022 17080 8910
rect 17188 8732 17496 8741
rect 17188 8730 17194 8732
rect 17250 8730 17274 8732
rect 17330 8730 17354 8732
rect 17410 8730 17434 8732
rect 17490 8730 17496 8732
rect 17250 8678 17252 8730
rect 17432 8678 17434 8730
rect 17188 8676 17194 8678
rect 17250 8676 17274 8678
rect 17330 8676 17354 8678
rect 17410 8676 17434 8678
rect 17490 8676 17496 8678
rect 17188 8667 17496 8676
rect 18064 8634 18092 9114
rect 18156 9042 18184 9454
rect 18144 9036 18196 9042
rect 18144 8978 18196 8984
rect 18616 8906 18644 10066
rect 18696 10056 18748 10062
rect 18696 9998 18748 10004
rect 18708 9674 18736 9998
rect 18708 9646 18828 9674
rect 18800 9042 18828 9646
rect 18892 9178 18920 10406
rect 19352 10282 19380 15370
rect 19628 14550 19656 15506
rect 19616 14544 19668 14550
rect 19616 14486 19668 14492
rect 19720 14414 19748 16186
rect 19708 14408 19760 14414
rect 19708 14350 19760 14356
rect 19812 14278 19840 19774
rect 19892 19712 19944 19718
rect 19892 19654 19944 19660
rect 19904 18222 19932 19654
rect 19984 19236 20036 19242
rect 19984 19178 20036 19184
rect 19892 18216 19944 18222
rect 19892 18158 19944 18164
rect 19892 17604 19944 17610
rect 19892 17546 19944 17552
rect 19904 14550 19932 17546
rect 19996 16250 20024 19178
rect 20088 17814 20116 19858
rect 20180 18426 20208 19858
rect 20260 19848 20312 19854
rect 20260 19790 20312 19796
rect 20272 18766 20300 19790
rect 20352 19712 20404 19718
rect 20352 19654 20404 19660
rect 20364 18902 20392 19654
rect 20444 19168 20496 19174
rect 20444 19110 20496 19116
rect 20456 18970 20484 19110
rect 20546 19068 20854 19077
rect 20546 19066 20552 19068
rect 20608 19066 20632 19068
rect 20688 19066 20712 19068
rect 20768 19066 20792 19068
rect 20848 19066 20854 19068
rect 20608 19014 20610 19066
rect 20790 19014 20792 19066
rect 20546 19012 20552 19014
rect 20608 19012 20632 19014
rect 20688 19012 20712 19014
rect 20768 19012 20792 19014
rect 20848 19012 20854 19014
rect 20546 19003 20854 19012
rect 20444 18964 20496 18970
rect 20444 18906 20496 18912
rect 20352 18896 20404 18902
rect 20352 18838 20404 18844
rect 20916 18834 20944 19858
rect 21100 19718 21128 21830
rect 21192 19854 21220 22066
rect 21180 19848 21232 19854
rect 21180 19790 21232 19796
rect 21088 19712 21140 19718
rect 21088 19654 21140 19660
rect 20996 19168 21048 19174
rect 20996 19110 21048 19116
rect 21008 18970 21036 19110
rect 20996 18964 21048 18970
rect 20996 18906 21048 18912
rect 21100 18850 21128 19654
rect 20904 18828 20956 18834
rect 20904 18770 20956 18776
rect 21008 18822 21128 18850
rect 20260 18760 20312 18766
rect 20260 18702 20312 18708
rect 20444 18624 20496 18630
rect 20444 18566 20496 18572
rect 20168 18420 20220 18426
rect 20168 18362 20220 18368
rect 20456 18222 20484 18566
rect 20444 18216 20496 18222
rect 20444 18158 20496 18164
rect 20546 17980 20854 17989
rect 20546 17978 20552 17980
rect 20608 17978 20632 17980
rect 20688 17978 20712 17980
rect 20768 17978 20792 17980
rect 20848 17978 20854 17980
rect 20608 17926 20610 17978
rect 20790 17926 20792 17978
rect 20546 17924 20552 17926
rect 20608 17924 20632 17926
rect 20688 17924 20712 17926
rect 20768 17924 20792 17926
rect 20848 17924 20854 17926
rect 20546 17915 20854 17924
rect 20076 17808 20128 17814
rect 20076 17750 20128 17756
rect 20916 17746 20944 18770
rect 21008 18426 21036 18822
rect 21088 18760 21140 18766
rect 21088 18702 21140 18708
rect 21100 18426 21128 18702
rect 21180 18624 21232 18630
rect 21180 18566 21232 18572
rect 20996 18420 21048 18426
rect 20996 18362 21048 18368
rect 21088 18420 21140 18426
rect 21088 18362 21140 18368
rect 20444 17740 20496 17746
rect 20444 17682 20496 17688
rect 20904 17740 20956 17746
rect 20904 17682 20956 17688
rect 20260 17604 20312 17610
rect 20260 17546 20312 17552
rect 20272 17338 20300 17546
rect 20260 17332 20312 17338
rect 20260 17274 20312 17280
rect 20352 17060 20404 17066
rect 20352 17002 20404 17008
rect 20364 16794 20392 17002
rect 20352 16788 20404 16794
rect 20352 16730 20404 16736
rect 19984 16244 20036 16250
rect 19984 16186 20036 16192
rect 19892 14544 19944 14550
rect 19892 14486 19944 14492
rect 19892 14408 19944 14414
rect 19892 14350 19944 14356
rect 19524 14272 19576 14278
rect 19524 14214 19576 14220
rect 19708 14272 19760 14278
rect 19708 14214 19760 14220
rect 19800 14272 19852 14278
rect 19800 14214 19852 14220
rect 19536 12850 19564 14214
rect 19524 12844 19576 12850
rect 19524 12786 19576 12792
rect 19720 12782 19748 14214
rect 19904 14074 19932 14350
rect 19892 14068 19944 14074
rect 19892 14010 19944 14016
rect 19996 13870 20024 16186
rect 20456 16046 20484 17682
rect 20546 16892 20854 16901
rect 20546 16890 20552 16892
rect 20608 16890 20632 16892
rect 20688 16890 20712 16892
rect 20768 16890 20792 16892
rect 20848 16890 20854 16892
rect 20608 16838 20610 16890
rect 20790 16838 20792 16890
rect 20546 16836 20552 16838
rect 20608 16836 20632 16838
rect 20688 16836 20712 16838
rect 20768 16836 20792 16838
rect 20848 16836 20854 16838
rect 20546 16827 20854 16836
rect 20444 16040 20496 16046
rect 20444 15982 20496 15988
rect 20904 15904 20956 15910
rect 20904 15846 20956 15852
rect 20546 15804 20854 15813
rect 20546 15802 20552 15804
rect 20608 15802 20632 15804
rect 20688 15802 20712 15804
rect 20768 15802 20792 15804
rect 20848 15802 20854 15804
rect 20608 15750 20610 15802
rect 20790 15750 20792 15802
rect 20546 15748 20552 15750
rect 20608 15748 20632 15750
rect 20688 15748 20712 15750
rect 20768 15748 20792 15750
rect 20848 15748 20854 15750
rect 20546 15739 20854 15748
rect 20260 15496 20312 15502
rect 20260 15438 20312 15444
rect 20272 15162 20300 15438
rect 20260 15156 20312 15162
rect 20260 15098 20312 15104
rect 20916 15042 20944 15846
rect 21008 15570 21036 18362
rect 21192 18086 21220 18566
rect 21180 18080 21232 18086
rect 21180 18022 21232 18028
rect 21088 16040 21140 16046
rect 21088 15982 21140 15988
rect 20996 15564 21048 15570
rect 20996 15506 21048 15512
rect 21100 15162 21128 15982
rect 21284 15706 21312 22358
rect 21468 22250 21496 22442
rect 21376 22222 21496 22250
rect 21376 22098 21404 22222
rect 21364 22092 21416 22098
rect 21364 22034 21416 22040
rect 21456 22094 21508 22098
rect 21560 22094 21588 24670
rect 21640 24676 21692 24682
rect 21640 24618 21692 24624
rect 21652 24274 21680 24618
rect 21640 24268 21692 24274
rect 21640 24210 21692 24216
rect 21744 23202 21772 26030
rect 21836 25838 21864 26472
rect 21916 26454 21968 26460
rect 22020 26450 22048 26744
rect 22100 26726 22152 26732
rect 22008 26444 22060 26450
rect 22008 26386 22060 26392
rect 21916 26240 21968 26246
rect 21916 26182 21968 26188
rect 21824 25832 21876 25838
rect 21824 25774 21876 25780
rect 21836 24818 21864 25774
rect 21824 24812 21876 24818
rect 21824 24754 21876 24760
rect 21928 23662 21956 26182
rect 22020 25838 22048 26386
rect 22296 26246 22324 27338
rect 22388 26926 22416 27950
rect 22652 27872 22704 27878
rect 22652 27814 22704 27820
rect 22664 27334 22692 27814
rect 22848 27606 22876 28358
rect 22940 27946 22968 28358
rect 22928 27940 22980 27946
rect 22928 27882 22980 27888
rect 23124 27674 23152 28562
rect 23296 28212 23348 28218
rect 23296 28154 23348 28160
rect 23308 27878 23336 28154
rect 23296 27872 23348 27878
rect 23296 27814 23348 27820
rect 23388 27872 23440 27878
rect 23388 27814 23440 27820
rect 23112 27668 23164 27674
rect 23112 27610 23164 27616
rect 22744 27600 22796 27606
rect 22744 27542 22796 27548
rect 22836 27600 22888 27606
rect 22836 27542 22888 27548
rect 22652 27328 22704 27334
rect 22652 27270 22704 27276
rect 22468 27124 22520 27130
rect 22468 27066 22520 27072
rect 22376 26920 22428 26926
rect 22376 26862 22428 26868
rect 22480 26586 22508 27066
rect 22468 26580 22520 26586
rect 22468 26522 22520 26528
rect 22284 26240 22336 26246
rect 22284 26182 22336 26188
rect 22296 26042 22324 26182
rect 22480 26042 22508 26522
rect 22664 26382 22692 27270
rect 22756 27130 22784 27542
rect 22848 27130 22876 27542
rect 22928 27532 22980 27538
rect 22928 27474 22980 27480
rect 22744 27124 22796 27130
rect 22744 27066 22796 27072
rect 22836 27124 22888 27130
rect 22836 27066 22888 27072
rect 22940 26926 22968 27474
rect 23400 27130 23428 27814
rect 23388 27124 23440 27130
rect 23388 27066 23440 27072
rect 22928 26920 22980 26926
rect 22928 26862 22980 26868
rect 22836 26444 22888 26450
rect 22836 26386 22888 26392
rect 22652 26376 22704 26382
rect 22652 26318 22704 26324
rect 22848 26042 22876 26386
rect 22940 26042 22968 26862
rect 23400 26790 23428 27066
rect 23492 27033 23520 29702
rect 23676 28914 23704 29990
rect 23860 29850 23888 30087
rect 24400 30058 24452 30064
rect 23940 30048 23992 30054
rect 23940 29990 23992 29996
rect 24216 30048 24268 30054
rect 24216 29990 24268 29996
rect 23848 29844 23900 29850
rect 23848 29786 23900 29792
rect 23756 29640 23808 29646
rect 23808 29617 23888 29628
rect 23808 29608 23902 29617
rect 23808 29600 23846 29608
rect 23756 29582 23808 29588
rect 23846 29543 23902 29552
rect 23756 29504 23808 29510
rect 23952 29492 23980 29990
rect 24228 29510 24256 29990
rect 24412 29850 24440 30058
rect 24492 30048 24544 30054
rect 24492 29990 24544 29996
rect 24860 30048 24912 30054
rect 24860 29990 24912 29996
rect 24400 29844 24452 29850
rect 24400 29786 24452 29792
rect 23808 29464 23980 29492
rect 24216 29504 24268 29510
rect 23756 29446 23808 29452
rect 24268 29464 24348 29492
rect 24216 29446 24268 29452
rect 23768 29306 23796 29446
rect 23904 29404 24212 29413
rect 23904 29402 23910 29404
rect 23966 29402 23990 29404
rect 24046 29402 24070 29404
rect 24126 29402 24150 29404
rect 24206 29402 24212 29404
rect 23966 29350 23968 29402
rect 24148 29350 24150 29402
rect 23904 29348 23910 29350
rect 23966 29348 23990 29350
rect 24046 29348 24070 29350
rect 24126 29348 24150 29350
rect 24206 29348 24212 29350
rect 23904 29339 24212 29348
rect 24320 29306 24348 29464
rect 24412 29306 24440 29786
rect 23756 29300 23808 29306
rect 23756 29242 23808 29248
rect 24308 29300 24360 29306
rect 24308 29242 24360 29248
rect 24400 29300 24452 29306
rect 24400 29242 24452 29248
rect 24504 29186 24532 29990
rect 24872 29850 24900 29990
rect 24860 29844 24912 29850
rect 24860 29786 24912 29792
rect 24676 29776 24728 29782
rect 24676 29718 24728 29724
rect 24584 29572 24636 29578
rect 24584 29514 24636 29520
rect 24596 29238 24624 29514
rect 24320 29170 24532 29186
rect 24584 29232 24636 29238
rect 24584 29174 24636 29180
rect 24308 29164 24532 29170
rect 24360 29158 24532 29164
rect 24308 29106 24360 29112
rect 24504 29102 24532 29158
rect 24492 29096 24544 29102
rect 24492 29038 24544 29044
rect 23584 28886 23704 28914
rect 24400 28960 24452 28966
rect 24400 28902 24452 28908
rect 24492 28960 24544 28966
rect 24492 28902 24544 28908
rect 23584 27946 23612 28886
rect 23904 28316 24212 28325
rect 23904 28314 23910 28316
rect 23966 28314 23990 28316
rect 24046 28314 24070 28316
rect 24126 28314 24150 28316
rect 24206 28314 24212 28316
rect 23966 28262 23968 28314
rect 24148 28262 24150 28314
rect 23904 28260 23910 28262
rect 23966 28260 23990 28262
rect 24046 28260 24070 28262
rect 24126 28260 24150 28262
rect 24206 28260 24212 28262
rect 23904 28251 24212 28260
rect 24412 28014 24440 28902
rect 24504 28014 24532 28902
rect 24584 28416 24636 28422
rect 24584 28358 24636 28364
rect 23664 28008 23716 28014
rect 23664 27950 23716 27956
rect 24216 28008 24268 28014
rect 24216 27950 24268 27956
rect 24400 28008 24452 28014
rect 24400 27950 24452 27956
rect 24492 28008 24544 28014
rect 24492 27950 24544 27956
rect 23572 27940 23624 27946
rect 23572 27882 23624 27888
rect 23478 27024 23534 27033
rect 23478 26959 23534 26968
rect 23492 26926 23520 26959
rect 23480 26920 23532 26926
rect 23480 26862 23532 26868
rect 23020 26784 23072 26790
rect 23020 26726 23072 26732
rect 23388 26784 23440 26790
rect 23388 26726 23440 26732
rect 23480 26784 23532 26790
rect 23480 26726 23532 26732
rect 22284 26036 22336 26042
rect 22284 25978 22336 25984
rect 22468 26036 22520 26042
rect 22468 25978 22520 25984
rect 22836 26036 22888 26042
rect 22836 25978 22888 25984
rect 22928 26036 22980 26042
rect 22928 25978 22980 25984
rect 23032 25838 23060 26726
rect 23492 26450 23520 26726
rect 23480 26444 23532 26450
rect 23480 26386 23532 26392
rect 23112 26308 23164 26314
rect 23112 26250 23164 26256
rect 22008 25832 22060 25838
rect 22008 25774 22060 25780
rect 22284 25832 22336 25838
rect 22284 25774 22336 25780
rect 23020 25832 23072 25838
rect 23020 25774 23072 25780
rect 22008 25288 22060 25294
rect 22008 25230 22060 25236
rect 22020 24886 22048 25230
rect 22008 24880 22060 24886
rect 22008 24822 22060 24828
rect 22020 24070 22048 24822
rect 22008 24064 22060 24070
rect 22008 24006 22060 24012
rect 21824 23656 21876 23662
rect 21824 23598 21876 23604
rect 21916 23656 21968 23662
rect 21916 23598 21968 23604
rect 21836 23322 21864 23598
rect 22020 23594 22140 23610
rect 22020 23588 22152 23594
rect 22020 23582 22100 23588
rect 21824 23316 21876 23322
rect 21824 23258 21876 23264
rect 21744 23174 21864 23202
rect 22020 23186 22048 23582
rect 22100 23530 22152 23536
rect 22192 23520 22244 23526
rect 22192 23462 22244 23468
rect 22204 23254 22232 23462
rect 22296 23322 22324 25774
rect 22560 25288 22612 25294
rect 22560 25230 22612 25236
rect 22572 24818 22600 25230
rect 22928 25220 22980 25226
rect 22928 25162 22980 25168
rect 22560 24812 22612 24818
rect 22560 24754 22612 24760
rect 22652 24744 22704 24750
rect 22652 24686 22704 24692
rect 22664 24410 22692 24686
rect 22836 24608 22888 24614
rect 22836 24550 22888 24556
rect 22652 24404 22704 24410
rect 22652 24346 22704 24352
rect 22664 23730 22692 24346
rect 22848 24206 22876 24550
rect 22940 24410 22968 25162
rect 23020 25152 23072 25158
rect 23020 25094 23072 25100
rect 23032 24750 23060 25094
rect 23124 24750 23152 26250
rect 23492 25906 23520 26386
rect 23572 26308 23624 26314
rect 23572 26250 23624 26256
rect 23584 26042 23612 26250
rect 23572 26036 23624 26042
rect 23572 25978 23624 25984
rect 23480 25900 23532 25906
rect 23480 25842 23532 25848
rect 23296 24812 23348 24818
rect 23296 24754 23348 24760
rect 23020 24744 23072 24750
rect 23020 24686 23072 24692
rect 23112 24744 23164 24750
rect 23112 24686 23164 24692
rect 22928 24404 22980 24410
rect 22928 24346 22980 24352
rect 23308 24274 23336 24754
rect 23480 24744 23532 24750
rect 23480 24686 23532 24692
rect 23492 24410 23520 24686
rect 23676 24410 23704 27950
rect 24228 27316 24256 27950
rect 24596 27946 24624 28358
rect 24584 27940 24636 27946
rect 24584 27882 24636 27888
rect 24492 27872 24544 27878
rect 24492 27814 24544 27820
rect 24228 27288 24348 27316
rect 23904 27228 24212 27237
rect 23904 27226 23910 27228
rect 23966 27226 23990 27228
rect 24046 27226 24070 27228
rect 24126 27226 24150 27228
rect 24206 27226 24212 27228
rect 23966 27174 23968 27226
rect 24148 27174 24150 27226
rect 23904 27172 23910 27174
rect 23966 27172 23990 27174
rect 24046 27172 24070 27174
rect 24126 27172 24150 27174
rect 24206 27172 24212 27174
rect 23904 27163 24212 27172
rect 24320 26586 24348 27288
rect 24308 26580 24360 26586
rect 24308 26522 24360 26528
rect 24400 26512 24452 26518
rect 24400 26454 24452 26460
rect 24308 26444 24360 26450
rect 24308 26386 24360 26392
rect 23904 26140 24212 26149
rect 23904 26138 23910 26140
rect 23966 26138 23990 26140
rect 24046 26138 24070 26140
rect 24126 26138 24150 26140
rect 24206 26138 24212 26140
rect 23966 26086 23968 26138
rect 24148 26086 24150 26138
rect 23904 26084 23910 26086
rect 23966 26084 23990 26086
rect 24046 26084 24070 26086
rect 24126 26084 24150 26086
rect 24206 26084 24212 26086
rect 23904 26075 24212 26084
rect 24320 26042 24348 26386
rect 24308 26036 24360 26042
rect 24308 25978 24360 25984
rect 24308 25696 24360 25702
rect 24308 25638 24360 25644
rect 23756 25288 23808 25294
rect 23756 25230 23808 25236
rect 23768 24614 23796 25230
rect 23904 25052 24212 25061
rect 23904 25050 23910 25052
rect 23966 25050 23990 25052
rect 24046 25050 24070 25052
rect 24126 25050 24150 25052
rect 24206 25050 24212 25052
rect 23966 24998 23968 25050
rect 24148 24998 24150 25050
rect 23904 24996 23910 24998
rect 23966 24996 23990 24998
rect 24046 24996 24070 24998
rect 24126 24996 24150 24998
rect 24206 24996 24212 24998
rect 23904 24987 24212 24996
rect 24124 24948 24176 24954
rect 24124 24890 24176 24896
rect 24136 24750 24164 24890
rect 24320 24886 24348 25638
rect 24308 24880 24360 24886
rect 24308 24822 24360 24828
rect 24124 24744 24176 24750
rect 24124 24686 24176 24692
rect 24308 24744 24360 24750
rect 24308 24686 24360 24692
rect 23756 24608 23808 24614
rect 23756 24550 23808 24556
rect 23480 24404 23532 24410
rect 23480 24346 23532 24352
rect 23664 24404 23716 24410
rect 23664 24346 23716 24352
rect 23296 24268 23348 24274
rect 23296 24210 23348 24216
rect 22836 24200 22888 24206
rect 22836 24142 22888 24148
rect 22652 23724 22704 23730
rect 22652 23666 22704 23672
rect 22664 23322 22692 23666
rect 23480 23520 23532 23526
rect 23480 23462 23532 23468
rect 22284 23316 22336 23322
rect 22284 23258 22336 23264
rect 22652 23316 22704 23322
rect 22652 23258 22704 23264
rect 22192 23248 22244 23254
rect 22192 23190 22244 23196
rect 21640 22568 21692 22574
rect 21640 22510 21692 22516
rect 21652 22098 21680 22510
rect 21732 22432 21784 22438
rect 21732 22374 21784 22380
rect 21744 22098 21772 22374
rect 21456 22092 21588 22094
rect 21508 22066 21588 22092
rect 21640 22092 21692 22098
rect 21456 22034 21508 22040
rect 21640 22034 21692 22040
rect 21732 22092 21784 22098
rect 21836 22094 21864 23174
rect 22008 23180 22060 23186
rect 22008 23122 22060 23128
rect 21916 23112 21968 23118
rect 21916 23054 21968 23060
rect 21928 22642 21956 23054
rect 23492 22982 23520 23462
rect 23480 22976 23532 22982
rect 23480 22918 23532 22924
rect 23572 22976 23624 22982
rect 23572 22918 23624 22924
rect 23584 22710 23612 22918
rect 23572 22704 23624 22710
rect 23572 22646 23624 22652
rect 21916 22636 21968 22642
rect 21916 22578 21968 22584
rect 23584 22506 23612 22646
rect 23572 22500 23624 22506
rect 23572 22442 23624 22448
rect 21836 22066 22048 22094
rect 21732 22034 21784 22040
rect 21376 21486 21404 22034
rect 21548 21888 21600 21894
rect 21548 21830 21600 21836
rect 21560 21690 21588 21830
rect 21548 21684 21600 21690
rect 21548 21626 21600 21632
rect 21652 21486 21680 22034
rect 21824 21956 21876 21962
rect 21824 21898 21876 21904
rect 21364 21480 21416 21486
rect 21364 21422 21416 21428
rect 21640 21480 21692 21486
rect 21640 21422 21692 21428
rect 21376 21010 21404 21422
rect 21652 21010 21680 21422
rect 21732 21344 21784 21350
rect 21732 21286 21784 21292
rect 21744 21146 21772 21286
rect 21732 21140 21784 21146
rect 21732 21082 21784 21088
rect 21836 21026 21864 21898
rect 21916 21412 21968 21418
rect 21916 21354 21968 21360
rect 21928 21078 21956 21354
rect 21744 21010 21864 21026
rect 21916 21072 21968 21078
rect 21916 21014 21968 21020
rect 21364 21004 21416 21010
rect 21364 20946 21416 20952
rect 21640 21004 21692 21010
rect 21640 20946 21692 20952
rect 21732 21004 21864 21010
rect 21784 20998 21864 21004
rect 21732 20946 21784 20952
rect 21824 19848 21876 19854
rect 21824 19790 21876 19796
rect 21836 19378 21864 19790
rect 21824 19372 21876 19378
rect 21824 19314 21876 19320
rect 21916 18964 21968 18970
rect 21916 18906 21968 18912
rect 21928 18222 21956 18906
rect 21916 18216 21968 18222
rect 21916 18158 21968 18164
rect 21824 17672 21876 17678
rect 21824 17614 21876 17620
rect 21640 17536 21692 17542
rect 21640 17478 21692 17484
rect 21364 16992 21416 16998
rect 21364 16934 21416 16940
rect 21376 16658 21404 16934
rect 21652 16794 21680 17478
rect 21836 17338 21864 17614
rect 21824 17332 21876 17338
rect 21824 17274 21876 17280
rect 22020 16794 22048 22066
rect 22928 22024 22980 22030
rect 22928 21966 22980 21972
rect 23572 22024 23624 22030
rect 23572 21966 23624 21972
rect 22940 21418 22968 21966
rect 23584 21690 23612 21966
rect 23572 21684 23624 21690
rect 23572 21626 23624 21632
rect 22928 21412 22980 21418
rect 22928 21354 22980 21360
rect 22284 21344 22336 21350
rect 22284 21286 22336 21292
rect 22296 20806 22324 21286
rect 22940 21146 22968 21354
rect 22928 21140 22980 21146
rect 22928 21082 22980 21088
rect 22284 20800 22336 20806
rect 22284 20742 22336 20748
rect 22296 20398 22324 20742
rect 22284 20392 22336 20398
rect 22284 20334 22336 20340
rect 23020 20392 23072 20398
rect 23020 20334 23072 20340
rect 23664 20392 23716 20398
rect 23664 20334 23716 20340
rect 22100 20256 22152 20262
rect 22100 20198 22152 20204
rect 22192 20256 22244 20262
rect 22192 20198 22244 20204
rect 22112 19786 22140 20198
rect 22204 19922 22232 20198
rect 22192 19916 22244 19922
rect 22192 19858 22244 19864
rect 22100 19780 22152 19786
rect 22100 19722 22152 19728
rect 22376 19780 22428 19786
rect 22376 19722 22428 19728
rect 22100 19372 22152 19378
rect 22100 19314 22152 19320
rect 22112 16794 22140 19314
rect 22284 19304 22336 19310
rect 22284 19246 22336 19252
rect 22192 18828 22244 18834
rect 22192 18770 22244 18776
rect 22204 18630 22232 18770
rect 22192 18624 22244 18630
rect 22192 18566 22244 18572
rect 22204 18154 22232 18566
rect 22296 18426 22324 19246
rect 22284 18420 22336 18426
rect 22284 18362 22336 18368
rect 22388 18306 22416 19722
rect 23032 19718 23060 20334
rect 23480 20256 23532 20262
rect 23480 20198 23532 20204
rect 22652 19712 22704 19718
rect 22652 19654 22704 19660
rect 23020 19712 23072 19718
rect 23020 19654 23072 19660
rect 22468 19304 22520 19310
rect 22468 19246 22520 19252
rect 22560 19304 22612 19310
rect 22560 19246 22612 19252
rect 22480 18426 22508 19246
rect 22572 18970 22600 19246
rect 22560 18964 22612 18970
rect 22560 18906 22612 18912
rect 22468 18420 22520 18426
rect 22468 18362 22520 18368
rect 22296 18278 22416 18306
rect 22192 18148 22244 18154
rect 22192 18090 22244 18096
rect 21640 16788 21692 16794
rect 21640 16730 21692 16736
rect 22008 16788 22060 16794
rect 22008 16730 22060 16736
rect 22100 16788 22152 16794
rect 22100 16730 22152 16736
rect 21364 16652 21416 16658
rect 21364 16594 21416 16600
rect 21456 15904 21508 15910
rect 21456 15846 21508 15852
rect 21272 15700 21324 15706
rect 21272 15642 21324 15648
rect 21088 15156 21140 15162
rect 21088 15098 21140 15104
rect 20824 15014 20944 15042
rect 20824 14822 20852 15014
rect 20904 14952 20956 14958
rect 20904 14894 20956 14900
rect 20812 14816 20864 14822
rect 20812 14758 20864 14764
rect 20546 14716 20854 14725
rect 20546 14714 20552 14716
rect 20608 14714 20632 14716
rect 20688 14714 20712 14716
rect 20768 14714 20792 14716
rect 20848 14714 20854 14716
rect 20608 14662 20610 14714
rect 20790 14662 20792 14714
rect 20546 14660 20552 14662
rect 20608 14660 20632 14662
rect 20688 14660 20712 14662
rect 20768 14660 20792 14662
rect 20848 14660 20854 14662
rect 20546 14651 20854 14660
rect 20352 14476 20404 14482
rect 20352 14418 20404 14424
rect 20260 14272 20312 14278
rect 20260 14214 20312 14220
rect 19984 13864 20036 13870
rect 19984 13806 20036 13812
rect 20272 13394 20300 14214
rect 20364 13394 20392 14418
rect 20444 13864 20496 13870
rect 20444 13806 20496 13812
rect 19892 13388 19944 13394
rect 19892 13330 19944 13336
rect 20260 13388 20312 13394
rect 20260 13330 20312 13336
rect 20352 13388 20404 13394
rect 20352 13330 20404 13336
rect 19904 12986 19932 13330
rect 20260 13184 20312 13190
rect 20260 13126 20312 13132
rect 19892 12980 19944 12986
rect 19892 12922 19944 12928
rect 19616 12776 19668 12782
rect 19616 12718 19668 12724
rect 19708 12776 19760 12782
rect 19708 12718 19760 12724
rect 19628 12442 19656 12718
rect 19616 12436 19668 12442
rect 19616 12378 19668 12384
rect 20272 12374 20300 13126
rect 20352 12912 20404 12918
rect 20352 12854 20404 12860
rect 20260 12368 20312 12374
rect 20260 12310 20312 12316
rect 19524 12300 19576 12306
rect 19524 12242 19576 12248
rect 19800 12300 19852 12306
rect 19800 12242 19852 12248
rect 19536 11898 19564 12242
rect 19524 11892 19576 11898
rect 19524 11834 19576 11840
rect 19812 11354 19840 12242
rect 19984 12232 20036 12238
rect 19984 12174 20036 12180
rect 19800 11348 19852 11354
rect 19800 11290 19852 11296
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19444 10674 19472 11086
rect 19432 10668 19484 10674
rect 19432 10610 19484 10616
rect 19708 10600 19760 10606
rect 19708 10542 19760 10548
rect 19168 10254 19380 10282
rect 19168 10062 19196 10254
rect 19156 10056 19208 10062
rect 19156 9998 19208 10004
rect 19340 10056 19392 10062
rect 19340 9998 19392 10004
rect 19064 9920 19116 9926
rect 19064 9862 19116 9868
rect 19076 9518 19104 9862
rect 19352 9722 19380 9998
rect 19720 9722 19748 10542
rect 19892 10464 19944 10470
rect 19892 10406 19944 10412
rect 19904 10266 19932 10406
rect 19892 10260 19944 10266
rect 19892 10202 19944 10208
rect 19996 10062 20024 12174
rect 20364 11694 20392 12854
rect 20352 11688 20404 11694
rect 20352 11630 20404 11636
rect 20350 10568 20406 10577
rect 20350 10503 20352 10512
rect 20404 10503 20406 10512
rect 20352 10474 20404 10480
rect 19984 10056 20036 10062
rect 19984 9998 20036 10004
rect 19340 9716 19392 9722
rect 19340 9658 19392 9664
rect 19708 9716 19760 9722
rect 19708 9658 19760 9664
rect 20260 9716 20312 9722
rect 20260 9658 20312 9664
rect 19064 9512 19116 9518
rect 19064 9454 19116 9460
rect 18972 9376 19024 9382
rect 18972 9318 19024 9324
rect 18880 9172 18932 9178
rect 18880 9114 18932 9120
rect 18984 9042 19012 9318
rect 19340 9172 19392 9178
rect 19340 9114 19392 9120
rect 18788 9036 18840 9042
rect 18788 8978 18840 8984
rect 18972 9036 19024 9042
rect 18972 8978 19024 8984
rect 18604 8900 18656 8906
rect 18800 8888 18828 8978
rect 19248 8900 19300 8906
rect 18800 8860 19248 8888
rect 18604 8842 18656 8848
rect 19248 8842 19300 8848
rect 18052 8628 18104 8634
rect 18052 8570 18104 8576
rect 18144 8560 18196 8566
rect 18144 8502 18196 8508
rect 17592 8424 17644 8430
rect 17592 8366 17644 8372
rect 16856 8016 16908 8022
rect 16856 7958 16908 7964
rect 17040 8016 17092 8022
rect 17040 7958 17092 7964
rect 16856 7744 16908 7750
rect 16856 7686 16908 7692
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 16212 7540 16264 7546
rect 16212 7482 16264 7488
rect 15384 6996 15436 7002
rect 15384 6938 15436 6944
rect 16868 6934 16896 7686
rect 17188 7644 17496 7653
rect 17188 7642 17194 7644
rect 17250 7642 17274 7644
rect 17330 7642 17354 7644
rect 17410 7642 17434 7644
rect 17490 7642 17496 7644
rect 17250 7590 17252 7642
rect 17432 7590 17434 7642
rect 17188 7588 17194 7590
rect 17250 7588 17274 7590
rect 17330 7588 17354 7590
rect 17410 7588 17434 7590
rect 17490 7588 17496 7590
rect 17188 7579 17496 7588
rect 17604 7546 17632 8366
rect 18052 8288 18104 8294
rect 18052 8230 18104 8236
rect 18064 7546 18092 8230
rect 18156 7954 18184 8502
rect 18616 8430 18644 8842
rect 18604 8424 18656 8430
rect 18604 8366 18656 8372
rect 19156 8424 19208 8430
rect 19156 8366 19208 8372
rect 18420 8288 18472 8294
rect 18420 8230 18472 8236
rect 18432 8090 18460 8230
rect 19168 8090 19196 8366
rect 18420 8084 18472 8090
rect 18420 8026 18472 8032
rect 19156 8084 19208 8090
rect 19156 8026 19208 8032
rect 18144 7948 18196 7954
rect 18144 7890 18196 7896
rect 19064 7948 19116 7954
rect 19064 7890 19116 7896
rect 17592 7540 17644 7546
rect 17592 7482 17644 7488
rect 18052 7540 18104 7546
rect 18052 7482 18104 7488
rect 17040 7268 17092 7274
rect 17040 7210 17092 7216
rect 16856 6928 16908 6934
rect 16856 6870 16908 6876
rect 15384 6860 15436 6866
rect 15384 6802 15436 6808
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 15200 6724 15252 6730
rect 15200 6666 15252 6672
rect 15292 6656 15344 6662
rect 15292 6598 15344 6604
rect 15198 6488 15254 6497
rect 15198 6423 15254 6432
rect 15212 6390 15240 6423
rect 15200 6384 15252 6390
rect 15200 6326 15252 6332
rect 15016 6190 15068 6196
rect 15106 6216 15162 6225
rect 15028 5642 15056 6190
rect 15106 6151 15162 6160
rect 15120 5914 15148 6151
rect 15200 6112 15252 6118
rect 15200 6054 15252 6060
rect 15108 5908 15160 5914
rect 15108 5850 15160 5856
rect 15016 5636 15068 5642
rect 15016 5578 15068 5584
rect 15212 5370 15240 6054
rect 15304 5710 15332 6598
rect 15396 6458 15424 6802
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 15844 6112 15896 6118
rect 15844 6054 15896 6060
rect 15856 5914 15884 6054
rect 15844 5908 15896 5914
rect 15844 5850 15896 5856
rect 16592 5778 16620 6802
rect 16672 6656 16724 6662
rect 16672 6598 16724 6604
rect 16684 6390 16712 6598
rect 16672 6384 16724 6390
rect 16672 6326 16724 6332
rect 16868 5778 16896 6870
rect 17052 6458 17080 7210
rect 18064 6866 18092 7482
rect 19076 7410 19104 7890
rect 19064 7404 19116 7410
rect 19064 7346 19116 7352
rect 19168 7342 19196 8026
rect 19260 7954 19288 8842
rect 19352 7954 19380 9114
rect 19524 9104 19576 9110
rect 19524 9046 19576 9052
rect 19432 8288 19484 8294
rect 19432 8230 19484 8236
rect 19248 7948 19300 7954
rect 19248 7890 19300 7896
rect 19340 7948 19392 7954
rect 19340 7890 19392 7896
rect 19156 7336 19208 7342
rect 19156 7278 19208 7284
rect 19260 7274 19288 7890
rect 19352 7342 19380 7890
rect 19444 7818 19472 8230
rect 19432 7812 19484 7818
rect 19432 7754 19484 7760
rect 19340 7336 19392 7342
rect 19340 7278 19392 7284
rect 19248 7268 19300 7274
rect 19248 7210 19300 7216
rect 18052 6860 18104 6866
rect 18052 6802 18104 6808
rect 19064 6860 19116 6866
rect 19064 6802 19116 6808
rect 17960 6792 18012 6798
rect 17960 6734 18012 6740
rect 17188 6556 17496 6565
rect 17188 6554 17194 6556
rect 17250 6554 17274 6556
rect 17330 6554 17354 6556
rect 17410 6554 17434 6556
rect 17490 6554 17496 6556
rect 17250 6502 17252 6554
rect 17432 6502 17434 6554
rect 17188 6500 17194 6502
rect 17250 6500 17274 6502
rect 17330 6500 17354 6502
rect 17410 6500 17434 6502
rect 17490 6500 17496 6502
rect 17188 6491 17496 6500
rect 17040 6452 17092 6458
rect 17040 6394 17092 6400
rect 17592 6248 17644 6254
rect 17592 6190 17644 6196
rect 17604 5914 17632 6190
rect 17684 6180 17736 6186
rect 17684 6122 17736 6128
rect 17696 5914 17724 6122
rect 17592 5908 17644 5914
rect 17592 5850 17644 5856
rect 17684 5908 17736 5914
rect 17684 5850 17736 5856
rect 17972 5778 18000 6734
rect 18328 6724 18380 6730
rect 18328 6666 18380 6672
rect 18052 6248 18104 6254
rect 18052 6190 18104 6196
rect 18064 5778 18092 6190
rect 18340 5914 18368 6666
rect 18420 6656 18472 6662
rect 18420 6598 18472 6604
rect 18432 6458 18460 6598
rect 19076 6458 19104 6802
rect 18420 6452 18472 6458
rect 18420 6394 18472 6400
rect 19064 6452 19116 6458
rect 19064 6394 19116 6400
rect 19444 6254 19472 7754
rect 19536 6866 19564 9046
rect 20272 9042 20300 9658
rect 20260 9036 20312 9042
rect 20260 8978 20312 8984
rect 19616 8492 19668 8498
rect 19616 8434 19668 8440
rect 19628 7478 19656 8434
rect 20456 8430 20484 13806
rect 20916 13734 20944 14894
rect 21284 14550 21312 15642
rect 21272 14544 21324 14550
rect 21272 14486 21324 14492
rect 20996 14272 21048 14278
rect 20996 14214 21048 14220
rect 20904 13728 20956 13734
rect 20904 13670 20956 13676
rect 20546 13628 20854 13637
rect 20546 13626 20552 13628
rect 20608 13626 20632 13628
rect 20688 13626 20712 13628
rect 20768 13626 20792 13628
rect 20848 13626 20854 13628
rect 20608 13574 20610 13626
rect 20790 13574 20792 13626
rect 20546 13572 20552 13574
rect 20608 13572 20632 13574
rect 20688 13572 20712 13574
rect 20768 13572 20792 13574
rect 20848 13572 20854 13574
rect 20546 13563 20854 13572
rect 20916 13462 20944 13670
rect 20904 13456 20956 13462
rect 20904 13398 20956 13404
rect 21008 13410 21036 14214
rect 21088 13796 21140 13802
rect 21088 13738 21140 13744
rect 21100 13530 21128 13738
rect 21088 13524 21140 13530
rect 21088 13466 21140 13472
rect 20536 13388 20588 13394
rect 21008 13382 21128 13410
rect 20536 13330 20588 13336
rect 20548 12782 20576 13330
rect 21100 13258 21128 13382
rect 21272 13388 21324 13394
rect 21272 13330 21324 13336
rect 21088 13252 21140 13258
rect 21088 13194 21140 13200
rect 20628 13184 20680 13190
rect 20628 13126 20680 13132
rect 20640 12850 20668 13126
rect 20628 12844 20680 12850
rect 20628 12786 20680 12792
rect 20536 12776 20588 12782
rect 20536 12718 20588 12724
rect 20720 12776 20772 12782
rect 20772 12736 20944 12764
rect 20720 12718 20772 12724
rect 20546 12540 20854 12549
rect 20546 12538 20552 12540
rect 20608 12538 20632 12540
rect 20688 12538 20712 12540
rect 20768 12538 20792 12540
rect 20848 12538 20854 12540
rect 20608 12486 20610 12538
rect 20790 12486 20792 12538
rect 20546 12484 20552 12486
rect 20608 12484 20632 12486
rect 20688 12484 20712 12486
rect 20768 12484 20792 12486
rect 20848 12484 20854 12486
rect 20546 12475 20854 12484
rect 20916 12442 20944 12736
rect 21100 12714 21128 13194
rect 21088 12708 21140 12714
rect 21088 12650 21140 12656
rect 21180 12708 21232 12714
rect 21180 12650 21232 12656
rect 20996 12640 21048 12646
rect 21192 12594 21220 12650
rect 21048 12588 21220 12594
rect 20996 12582 21220 12588
rect 21008 12566 21220 12582
rect 20904 12436 20956 12442
rect 20904 12378 20956 12384
rect 21284 12306 21312 13330
rect 21468 13274 21496 15846
rect 21916 15360 21968 15366
rect 21916 15302 21968 15308
rect 21928 14958 21956 15302
rect 21916 14952 21968 14958
rect 21916 14894 21968 14900
rect 21548 14272 21600 14278
rect 21548 14214 21600 14220
rect 21560 13394 21588 14214
rect 21548 13388 21600 13394
rect 21548 13330 21600 13336
rect 21468 13246 21588 13274
rect 21456 12640 21508 12646
rect 21456 12582 21508 12588
rect 21468 12322 21496 12582
rect 21560 12434 21588 13246
rect 22020 12442 22048 16730
rect 22296 15434 22324 18278
rect 22468 17740 22520 17746
rect 22468 17682 22520 17688
rect 22480 17270 22508 17682
rect 22560 17536 22612 17542
rect 22560 17478 22612 17484
rect 22468 17264 22520 17270
rect 22468 17206 22520 17212
rect 22376 16992 22428 16998
rect 22376 16934 22428 16940
rect 22388 16794 22416 16934
rect 22572 16794 22600 17478
rect 22376 16788 22428 16794
rect 22376 16730 22428 16736
rect 22560 16788 22612 16794
rect 22560 16730 22612 16736
rect 22376 16448 22428 16454
rect 22376 16390 22428 16396
rect 22284 15428 22336 15434
rect 22284 15370 22336 15376
rect 22284 14816 22336 14822
rect 22284 14758 22336 14764
rect 22296 14618 22324 14758
rect 22388 14618 22416 16390
rect 22664 16046 22692 19654
rect 22744 19440 22796 19446
rect 22744 19382 22796 19388
rect 22756 18426 22784 19382
rect 22836 19168 22888 19174
rect 22836 19110 22888 19116
rect 22848 18698 22876 19110
rect 23032 18834 23060 19654
rect 23388 19236 23440 19242
rect 23388 19178 23440 19184
rect 23112 19168 23164 19174
rect 23112 19110 23164 19116
rect 23124 18970 23152 19110
rect 23112 18964 23164 18970
rect 23112 18906 23164 18912
rect 23020 18828 23072 18834
rect 23020 18770 23072 18776
rect 22836 18692 22888 18698
rect 22836 18634 22888 18640
rect 22848 18426 22876 18634
rect 22744 18420 22796 18426
rect 22744 18362 22796 18368
rect 22836 18420 22888 18426
rect 22836 18362 22888 18368
rect 22756 17898 22784 18362
rect 23124 18222 23152 18906
rect 23400 18714 23428 19178
rect 23492 18902 23520 20198
rect 23676 19514 23704 20334
rect 23572 19508 23624 19514
rect 23572 19450 23624 19456
rect 23664 19508 23716 19514
rect 23664 19450 23716 19456
rect 23480 18896 23532 18902
rect 23480 18838 23532 18844
rect 23400 18686 23520 18714
rect 23492 18306 23520 18686
rect 23584 18426 23612 19450
rect 23572 18420 23624 18426
rect 23572 18362 23624 18368
rect 23492 18278 23612 18306
rect 23112 18216 23164 18222
rect 23112 18158 23164 18164
rect 23204 18216 23256 18222
rect 23204 18158 23256 18164
rect 23296 18216 23348 18222
rect 23296 18158 23348 18164
rect 22756 17870 22876 17898
rect 23216 17882 23244 18158
rect 22744 17740 22796 17746
rect 22744 17682 22796 17688
rect 22756 17270 22784 17682
rect 22744 17264 22796 17270
rect 22744 17206 22796 17212
rect 22848 17134 22876 17870
rect 23204 17876 23256 17882
rect 23204 17818 23256 17824
rect 23216 17134 23244 17818
rect 23308 17626 23336 18158
rect 23584 17814 23612 18278
rect 23572 17808 23624 17814
rect 23572 17750 23624 17756
rect 23308 17598 23428 17626
rect 23296 17536 23348 17542
rect 23296 17478 23348 17484
rect 23308 17134 23336 17478
rect 22836 17128 22888 17134
rect 22836 17070 22888 17076
rect 23204 17128 23256 17134
rect 23204 17070 23256 17076
rect 23296 17128 23348 17134
rect 23296 17070 23348 17076
rect 23020 16992 23072 16998
rect 23020 16934 23072 16940
rect 23112 16992 23164 16998
rect 23112 16934 23164 16940
rect 23032 16794 23060 16934
rect 23020 16788 23072 16794
rect 23020 16730 23072 16736
rect 23020 16652 23072 16658
rect 23020 16594 23072 16600
rect 23032 16522 23060 16594
rect 23020 16516 23072 16522
rect 23020 16458 23072 16464
rect 23124 16454 23152 16934
rect 23400 16538 23428 17598
rect 23216 16510 23428 16538
rect 23112 16448 23164 16454
rect 23112 16390 23164 16396
rect 22652 16040 22704 16046
rect 22652 15982 22704 15988
rect 22664 15570 22692 15982
rect 22652 15564 22704 15570
rect 22652 15506 22704 15512
rect 22928 15496 22980 15502
rect 22928 15438 22980 15444
rect 22940 15094 22968 15438
rect 22928 15088 22980 15094
rect 22928 15030 22980 15036
rect 23216 15042 23244 16510
rect 23296 16448 23348 16454
rect 23296 16390 23348 16396
rect 23388 16448 23440 16454
rect 23388 16390 23440 16396
rect 23308 15706 23336 16390
rect 23296 15700 23348 15706
rect 23296 15642 23348 15648
rect 23296 15496 23348 15502
rect 23296 15438 23348 15444
rect 23308 15162 23336 15438
rect 23296 15156 23348 15162
rect 23296 15098 23348 15104
rect 23216 15014 23336 15042
rect 22836 14952 22888 14958
rect 22836 14894 22888 14900
rect 22284 14612 22336 14618
rect 22284 14554 22336 14560
rect 22376 14612 22428 14618
rect 22376 14554 22428 14560
rect 22284 14272 22336 14278
rect 22284 14214 22336 14220
rect 22468 14272 22520 14278
rect 22468 14214 22520 14220
rect 22008 12436 22060 12442
rect 21560 12406 21680 12434
rect 21548 12368 21600 12374
rect 21468 12316 21548 12322
rect 21468 12310 21600 12316
rect 21272 12300 21324 12306
rect 21468 12294 21588 12310
rect 21272 12242 21324 12248
rect 21284 11898 21312 12242
rect 21272 11892 21324 11898
rect 21272 11834 21324 11840
rect 20546 11452 20854 11461
rect 20546 11450 20552 11452
rect 20608 11450 20632 11452
rect 20688 11450 20712 11452
rect 20768 11450 20792 11452
rect 20848 11450 20854 11452
rect 20608 11398 20610 11450
rect 20790 11398 20792 11450
rect 20546 11396 20552 11398
rect 20608 11396 20632 11398
rect 20688 11396 20712 11398
rect 20768 11396 20792 11398
rect 20848 11396 20854 11398
rect 20546 11387 20854 11396
rect 21272 10668 21324 10674
rect 21272 10610 21324 10616
rect 20904 10600 20956 10606
rect 20904 10542 20956 10548
rect 20546 10364 20854 10373
rect 20546 10362 20552 10364
rect 20608 10362 20632 10364
rect 20688 10362 20712 10364
rect 20768 10362 20792 10364
rect 20848 10362 20854 10364
rect 20608 10310 20610 10362
rect 20790 10310 20792 10362
rect 20546 10308 20552 10310
rect 20608 10308 20632 10310
rect 20688 10308 20712 10310
rect 20768 10308 20792 10310
rect 20848 10308 20854 10310
rect 20546 10299 20854 10308
rect 20916 9722 20944 10542
rect 20996 10464 21048 10470
rect 20996 10406 21048 10412
rect 21088 10464 21140 10470
rect 21088 10406 21140 10412
rect 21008 9926 21036 10406
rect 21100 10062 21128 10406
rect 21284 10266 21312 10610
rect 21548 10600 21600 10606
rect 21652 10588 21680 12406
rect 22008 12378 22060 12384
rect 22296 10674 22324 14214
rect 22480 13394 22508 14214
rect 22744 14068 22796 14074
rect 22744 14010 22796 14016
rect 22468 13388 22520 13394
rect 22468 13330 22520 13336
rect 22468 12776 22520 12782
rect 22468 12718 22520 12724
rect 22480 12442 22508 12718
rect 22560 12640 22612 12646
rect 22560 12582 22612 12588
rect 22468 12436 22520 12442
rect 22468 12378 22520 12384
rect 22572 11694 22600 12582
rect 22560 11688 22612 11694
rect 22560 11630 22612 11636
rect 22284 10668 22336 10674
rect 22284 10610 22336 10616
rect 21600 10560 21680 10588
rect 21916 10600 21968 10606
rect 21548 10542 21600 10548
rect 21916 10542 21968 10548
rect 22192 10600 22244 10606
rect 22192 10542 22244 10548
rect 21272 10260 21324 10266
rect 21272 10202 21324 10208
rect 21180 10192 21232 10198
rect 21180 10134 21232 10140
rect 21088 10056 21140 10062
rect 21088 9998 21140 10004
rect 20996 9920 21048 9926
rect 20996 9862 21048 9868
rect 20904 9716 20956 9722
rect 20904 9658 20956 9664
rect 21008 9382 21036 9862
rect 21100 9722 21128 9998
rect 21088 9716 21140 9722
rect 21088 9658 21140 9664
rect 20996 9376 21048 9382
rect 20996 9318 21048 9324
rect 20546 9276 20854 9285
rect 20546 9274 20552 9276
rect 20608 9274 20632 9276
rect 20688 9274 20712 9276
rect 20768 9274 20792 9276
rect 20848 9274 20854 9276
rect 20608 9222 20610 9274
rect 20790 9222 20792 9274
rect 20546 9220 20552 9222
rect 20608 9220 20632 9222
rect 20688 9220 20712 9222
rect 20768 9220 20792 9222
rect 20848 9220 20854 9222
rect 20546 9211 20854 9220
rect 20628 8968 20680 8974
rect 20628 8910 20680 8916
rect 20640 8498 20668 8910
rect 20628 8492 20680 8498
rect 20628 8434 20680 8440
rect 20444 8424 20496 8430
rect 20444 8366 20496 8372
rect 20904 8288 20956 8294
rect 20904 8230 20956 8236
rect 20546 8188 20854 8197
rect 20546 8186 20552 8188
rect 20608 8186 20632 8188
rect 20688 8186 20712 8188
rect 20768 8186 20792 8188
rect 20848 8186 20854 8188
rect 20608 8134 20610 8186
rect 20790 8134 20792 8186
rect 20546 8132 20552 8134
rect 20608 8132 20632 8134
rect 20688 8132 20712 8134
rect 20768 8132 20792 8134
rect 20848 8132 20854 8134
rect 20546 8123 20854 8132
rect 20916 8090 20944 8230
rect 20904 8084 20956 8090
rect 20904 8026 20956 8032
rect 20444 7744 20496 7750
rect 20444 7686 20496 7692
rect 19616 7472 19668 7478
rect 19616 7414 19668 7420
rect 20352 7200 20404 7206
rect 20352 7142 20404 7148
rect 19892 6928 19944 6934
rect 19892 6870 19944 6876
rect 19524 6860 19576 6866
rect 19524 6802 19576 6808
rect 19800 6860 19852 6866
rect 19800 6802 19852 6808
rect 19524 6656 19576 6662
rect 19524 6598 19576 6604
rect 19432 6248 19484 6254
rect 19432 6190 19484 6196
rect 18880 6112 18932 6118
rect 18880 6054 18932 6060
rect 18892 5914 18920 6054
rect 18328 5908 18380 5914
rect 18328 5850 18380 5856
rect 18880 5908 18932 5914
rect 18880 5850 18932 5856
rect 16580 5772 16632 5778
rect 16580 5714 16632 5720
rect 16856 5772 16908 5778
rect 16856 5714 16908 5720
rect 17960 5772 18012 5778
rect 17960 5714 18012 5720
rect 18052 5772 18104 5778
rect 18052 5714 18104 5720
rect 18144 5772 18196 5778
rect 18144 5714 18196 5720
rect 15292 5704 15344 5710
rect 15292 5646 15344 5652
rect 15568 5568 15620 5574
rect 15568 5510 15620 5516
rect 15200 5364 15252 5370
rect 15200 5306 15252 5312
rect 15580 5166 15608 5510
rect 16592 5370 16620 5714
rect 17188 5468 17496 5477
rect 17188 5466 17194 5468
rect 17250 5466 17274 5468
rect 17330 5466 17354 5468
rect 17410 5466 17434 5468
rect 17490 5466 17496 5468
rect 17250 5414 17252 5466
rect 17432 5414 17434 5466
rect 17188 5412 17194 5414
rect 17250 5412 17274 5414
rect 17330 5412 17354 5414
rect 17410 5412 17434 5414
rect 17490 5412 17496 5414
rect 17188 5403 17496 5412
rect 16580 5364 16632 5370
rect 16580 5306 16632 5312
rect 15292 5160 15344 5166
rect 15292 5102 15344 5108
rect 15568 5160 15620 5166
rect 15568 5102 15620 5108
rect 15304 4826 15332 5102
rect 18064 4826 18092 5714
rect 18156 5642 18184 5714
rect 18144 5636 18196 5642
rect 18144 5578 18196 5584
rect 14476 3692 14596 3720
rect 14660 4780 14780 4808
rect 15292 4820 15344 4826
rect 14372 3596 14424 3602
rect 14372 3538 14424 3544
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 14384 3466 14412 3538
rect 14372 3460 14424 3466
rect 14372 3402 14424 3408
rect 13820 3188 13872 3194
rect 13820 3130 13872 3136
rect 14188 3188 14240 3194
rect 14188 3130 14240 3136
rect 14384 3126 14412 3402
rect 14476 3398 14504 3692
rect 14556 3596 14608 3602
rect 14556 3538 14608 3544
rect 14464 3392 14516 3398
rect 14464 3334 14516 3340
rect 14096 3120 14148 3126
rect 14372 3120 14424 3126
rect 14148 3068 14228 3074
rect 14096 3062 14228 3068
rect 14372 3062 14424 3068
rect 14108 3046 14228 3062
rect 13728 2984 13780 2990
rect 13728 2926 13780 2932
rect 13820 2984 13872 2990
rect 13820 2926 13872 2932
rect 13832 2836 13860 2926
rect 14200 2922 14228 3046
rect 14280 2984 14332 2990
rect 14280 2926 14332 2932
rect 14188 2916 14240 2922
rect 14188 2858 14240 2864
rect 13740 2808 13860 2836
rect 13740 2650 13768 2808
rect 13830 2748 14138 2757
rect 13830 2746 13836 2748
rect 13892 2746 13916 2748
rect 13972 2746 13996 2748
rect 14052 2746 14076 2748
rect 14132 2746 14138 2748
rect 13892 2694 13894 2746
rect 14074 2694 14076 2746
rect 13830 2692 13836 2694
rect 13892 2692 13916 2694
rect 13972 2692 13996 2694
rect 14052 2692 14076 2694
rect 14132 2692 14138 2694
rect 13830 2683 14138 2692
rect 13728 2644 13780 2650
rect 13780 2604 13860 2632
rect 13728 2586 13780 2592
rect 12768 2468 12848 2496
rect 12900 2508 12952 2514
rect 12716 2450 12768 2456
rect 12900 2450 12952 2456
rect 13636 2508 13688 2514
rect 13636 2450 13688 2456
rect 10968 2372 11020 2378
rect 10968 2314 11020 2320
rect 12624 2372 12676 2378
rect 12624 2314 12676 2320
rect 10980 2088 11008 2314
rect 11888 2304 11940 2310
rect 11888 2246 11940 2252
rect 11980 2304 12032 2310
rect 11980 2246 12032 2252
rect 11060 2100 11112 2106
rect 10980 2060 11060 2088
rect 11060 2042 11112 2048
rect 10836 1856 10916 1884
rect 11612 1896 11664 1902
rect 10784 1838 10836 1844
rect 11612 1838 11664 1844
rect 11704 1896 11756 1902
rect 11704 1838 11756 1844
rect 10324 1828 10376 1834
rect 10324 1770 10376 1776
rect 9916 1380 10088 1408
rect 9864 1362 9916 1368
rect 10336 1018 10364 1770
rect 11152 1760 11204 1766
rect 11152 1702 11204 1708
rect 10692 1420 10744 1426
rect 10744 1380 10916 1408
rect 10692 1362 10744 1368
rect 10472 1116 10780 1125
rect 10472 1114 10478 1116
rect 10534 1114 10558 1116
rect 10614 1114 10638 1116
rect 10694 1114 10718 1116
rect 10774 1114 10780 1116
rect 10534 1062 10536 1114
rect 10716 1062 10718 1114
rect 10472 1060 10478 1062
rect 10534 1060 10558 1062
rect 10614 1060 10638 1062
rect 10694 1060 10718 1062
rect 10774 1060 10780 1062
rect 10472 1051 10780 1060
rect 10324 1012 10376 1018
rect 10324 954 10376 960
rect 9732 768 9812 796
rect 10048 808 10100 814
rect 9680 750 9732 756
rect 10048 750 10100 756
rect 10060 400 10088 750
rect 10612 462 10732 490
rect 10612 400 10640 462
rect 7024 326 7236 354
rect 7286 0 7342 400
rect 7838 0 7894 400
rect 8390 0 8446 400
rect 8942 0 8998 400
rect 9494 0 9550 400
rect 10046 0 10102 400
rect 10598 0 10654 400
rect 10704 354 10732 462
rect 10888 354 10916 1380
rect 11060 1352 11112 1358
rect 11060 1294 11112 1300
rect 11072 1018 11100 1294
rect 11060 1012 11112 1018
rect 11060 954 11112 960
rect 11164 400 11192 1702
rect 11624 898 11652 1838
rect 11716 1018 11744 1838
rect 11900 1562 11928 2246
rect 11992 1902 12020 2246
rect 11980 1896 12032 1902
rect 11980 1838 12032 1844
rect 11888 1556 11940 1562
rect 11888 1498 11940 1504
rect 12636 1426 12664 2314
rect 12716 2304 12768 2310
rect 12716 2246 12768 2252
rect 12164 1420 12216 1426
rect 12624 1420 12676 1426
rect 12216 1380 12296 1408
rect 12164 1362 12216 1368
rect 11704 1012 11756 1018
rect 11704 954 11756 960
rect 11624 870 11744 898
rect 11716 400 11744 870
rect 12268 400 12296 1380
rect 12624 1362 12676 1368
rect 12728 814 12756 2246
rect 12808 1896 12860 1902
rect 12808 1838 12860 1844
rect 12900 1896 12952 1902
rect 12900 1838 12952 1844
rect 13176 1896 13228 1902
rect 13832 1850 13860 2604
rect 14200 2514 14228 2858
rect 14292 2514 14320 2926
rect 14568 2774 14596 3538
rect 14660 3505 14688 4780
rect 15292 4762 15344 4768
rect 18052 4820 18104 4826
rect 18052 4762 18104 4768
rect 14740 4684 14792 4690
rect 14740 4626 14792 4632
rect 14924 4684 14976 4690
rect 14924 4626 14976 4632
rect 16580 4684 16632 4690
rect 16580 4626 16632 4632
rect 17592 4684 17644 4690
rect 17592 4626 17644 4632
rect 17684 4684 17736 4690
rect 17684 4626 17736 4632
rect 14646 3496 14702 3505
rect 14646 3431 14702 3440
rect 14568 2746 14688 2774
rect 14188 2508 14240 2514
rect 14188 2450 14240 2456
rect 14280 2508 14332 2514
rect 14280 2450 14332 2456
rect 14660 2378 14688 2746
rect 14648 2372 14700 2378
rect 14648 2314 14700 2320
rect 14752 2310 14780 4626
rect 14936 3738 14964 4626
rect 15016 4208 15068 4214
rect 15016 4150 15068 4156
rect 14924 3732 14976 3738
rect 14924 3674 14976 3680
rect 14832 3596 14884 3602
rect 14832 3538 14884 3544
rect 14740 2304 14792 2310
rect 14740 2246 14792 2252
rect 13176 1838 13228 1844
rect 12716 808 12768 814
rect 12716 750 12768 756
rect 12820 400 12848 1838
rect 12912 1426 12940 1838
rect 12900 1420 12952 1426
rect 12900 1362 12952 1368
rect 13188 1018 13216 1838
rect 13740 1822 13860 1850
rect 14188 1896 14240 1902
rect 14188 1838 14240 1844
rect 14648 1896 14700 1902
rect 14648 1838 14700 1844
rect 13740 1426 13768 1822
rect 13830 1660 14138 1669
rect 13830 1658 13836 1660
rect 13892 1658 13916 1660
rect 13972 1658 13996 1660
rect 14052 1658 14076 1660
rect 14132 1658 14138 1660
rect 13892 1606 13894 1658
rect 14074 1606 14076 1658
rect 13830 1604 13836 1606
rect 13892 1604 13916 1606
rect 13972 1604 13996 1606
rect 14052 1604 14076 1606
rect 14132 1604 14138 1606
rect 13830 1595 14138 1604
rect 13636 1420 13688 1426
rect 13636 1362 13688 1368
rect 13728 1420 13780 1426
rect 13728 1362 13780 1368
rect 13452 1352 13504 1358
rect 13452 1294 13504 1300
rect 13464 1018 13492 1294
rect 13176 1012 13228 1018
rect 13176 954 13228 960
rect 13452 1012 13504 1018
rect 13452 954 13504 960
rect 13360 808 13412 814
rect 13360 750 13412 756
rect 13372 400 13400 750
rect 13648 456 13676 1362
rect 14200 1018 14228 1838
rect 14660 1426 14688 1838
rect 14556 1420 14608 1426
rect 14476 1380 14556 1408
rect 14188 1012 14240 1018
rect 14188 954 14240 960
rect 13830 572 14138 581
rect 13830 570 13836 572
rect 13892 570 13916 572
rect 13972 570 13996 572
rect 14052 570 14076 572
rect 14132 570 14138 572
rect 13892 518 13894 570
rect 14074 518 14076 570
rect 13830 516 13836 518
rect 13892 516 13916 518
rect 13972 516 13996 518
rect 14052 516 14076 518
rect 14132 516 14138 518
rect 13830 507 14138 516
rect 13648 428 13952 456
rect 13924 400 13952 428
rect 14476 400 14504 1380
rect 14556 1362 14608 1368
rect 14648 1420 14700 1426
rect 14648 1362 14700 1368
rect 14844 814 14872 3538
rect 14924 3528 14976 3534
rect 14924 3470 14976 3476
rect 14936 3369 14964 3470
rect 14922 3360 14978 3369
rect 14922 3295 14978 3304
rect 15028 2990 15056 4150
rect 16592 4078 16620 4626
rect 17188 4380 17496 4389
rect 17188 4378 17194 4380
rect 17250 4378 17274 4380
rect 17330 4378 17354 4380
rect 17410 4378 17434 4380
rect 17490 4378 17496 4380
rect 17250 4326 17252 4378
rect 17432 4326 17434 4378
rect 17188 4324 17194 4326
rect 17250 4324 17274 4326
rect 17330 4324 17354 4326
rect 17410 4324 17434 4326
rect 17490 4324 17496 4326
rect 17188 4315 17496 4324
rect 15292 4072 15344 4078
rect 15292 4014 15344 4020
rect 15568 4072 15620 4078
rect 15568 4014 15620 4020
rect 16580 4072 16632 4078
rect 16580 4014 16632 4020
rect 15304 3738 15332 4014
rect 15384 3936 15436 3942
rect 15384 3878 15436 3884
rect 15292 3732 15344 3738
rect 15292 3674 15344 3680
rect 15396 3602 15424 3878
rect 15384 3596 15436 3602
rect 15384 3538 15436 3544
rect 15108 3392 15160 3398
rect 15108 3334 15160 3340
rect 15476 3392 15528 3398
rect 15476 3334 15528 3340
rect 15120 3194 15148 3334
rect 15488 3194 15516 3334
rect 15580 3194 15608 4014
rect 17604 4010 17632 4626
rect 17696 4282 17724 4626
rect 17868 4616 17920 4622
rect 17868 4558 17920 4564
rect 17684 4276 17736 4282
rect 17684 4218 17736 4224
rect 17592 4004 17644 4010
rect 17592 3946 17644 3952
rect 15750 3632 15806 3641
rect 15660 3596 15712 3602
rect 15750 3567 15752 3576
rect 15660 3538 15712 3544
rect 15804 3567 15806 3576
rect 15752 3538 15804 3544
rect 15672 3380 15700 3538
rect 17604 3534 17632 3946
rect 17696 3738 17724 4218
rect 17880 4078 17908 4558
rect 18156 4554 18184 5578
rect 18696 5296 18748 5302
rect 18696 5238 18748 5244
rect 18144 4548 18196 4554
rect 18144 4490 18196 4496
rect 18236 4480 18288 4486
rect 18236 4422 18288 4428
rect 18248 4214 18276 4422
rect 18236 4208 18288 4214
rect 18236 4150 18288 4156
rect 17868 4072 17920 4078
rect 17868 4014 17920 4020
rect 17880 3942 17908 4014
rect 18708 4010 18736 5238
rect 19340 4684 19392 4690
rect 19340 4626 19392 4632
rect 19352 4282 19380 4626
rect 19444 4486 19472 6190
rect 19536 6186 19564 6598
rect 19524 6180 19576 6186
rect 19524 6122 19576 6128
rect 19812 5166 19840 6802
rect 19800 5160 19852 5166
rect 19800 5102 19852 5108
rect 19708 4684 19760 4690
rect 19708 4626 19760 4632
rect 19432 4480 19484 4486
rect 19432 4422 19484 4428
rect 19340 4276 19392 4282
rect 19340 4218 19392 4224
rect 18696 4004 18748 4010
rect 18696 3946 18748 3952
rect 17868 3936 17920 3942
rect 17868 3878 17920 3884
rect 18052 3936 18104 3942
rect 18052 3878 18104 3884
rect 17684 3732 17736 3738
rect 17684 3674 17736 3680
rect 17880 3602 17908 3878
rect 18064 3738 18092 3878
rect 18052 3732 18104 3738
rect 18052 3674 18104 3680
rect 17868 3596 17920 3602
rect 17868 3538 17920 3544
rect 17592 3528 17644 3534
rect 17592 3470 17644 3476
rect 16488 3392 16540 3398
rect 15672 3352 15976 3380
rect 15108 3188 15160 3194
rect 15108 3130 15160 3136
rect 15476 3188 15528 3194
rect 15476 3130 15528 3136
rect 15568 3188 15620 3194
rect 15568 3130 15620 3136
rect 15016 2984 15068 2990
rect 15016 2926 15068 2932
rect 15488 2650 15516 3130
rect 15844 2916 15896 2922
rect 15844 2858 15896 2864
rect 15476 2644 15528 2650
rect 15476 2586 15528 2592
rect 15384 2576 15436 2582
rect 15384 2518 15436 2524
rect 15016 2508 15068 2514
rect 15016 2450 15068 2456
rect 14924 2304 14976 2310
rect 14924 2246 14976 2252
rect 14936 1426 14964 2246
rect 15028 2106 15056 2450
rect 15016 2100 15068 2106
rect 15016 2042 15068 2048
rect 15396 1902 15424 2518
rect 15384 1896 15436 1902
rect 15384 1838 15436 1844
rect 15856 1426 15884 2858
rect 14924 1420 14976 1426
rect 15752 1420 15804 1426
rect 14924 1362 14976 1368
rect 15580 1380 15752 1408
rect 14832 808 14884 814
rect 14832 750 14884 756
rect 15016 808 15068 814
rect 15016 750 15068 756
rect 15028 400 15056 750
rect 15580 400 15608 1380
rect 15752 1362 15804 1368
rect 15844 1420 15896 1426
rect 15844 1362 15896 1368
rect 15948 746 15976 3352
rect 16488 3334 16540 3340
rect 17040 3392 17092 3398
rect 17040 3334 17092 3340
rect 16500 3194 16528 3334
rect 16488 3188 16540 3194
rect 16488 3130 16540 3136
rect 16212 2984 16264 2990
rect 16212 2926 16264 2932
rect 16224 2514 16252 2926
rect 16212 2508 16264 2514
rect 16212 2450 16264 2456
rect 16948 2508 17000 2514
rect 16948 2450 17000 2456
rect 16960 2106 16988 2450
rect 16948 2100 17000 2106
rect 16948 2042 17000 2048
rect 16304 1896 16356 1902
rect 16224 1856 16304 1884
rect 16120 1352 16172 1358
rect 16120 1294 16172 1300
rect 16132 1018 16160 1294
rect 16120 1012 16172 1018
rect 16120 954 16172 960
rect 16224 898 16252 1856
rect 16304 1838 16356 1844
rect 16396 1896 16448 1902
rect 16396 1838 16448 1844
rect 16132 870 16252 898
rect 15936 740 15988 746
rect 15936 682 15988 688
rect 16132 400 16160 870
rect 16408 814 16436 1838
rect 17052 1494 17080 3334
rect 17188 3292 17496 3301
rect 17188 3290 17194 3292
rect 17250 3290 17274 3292
rect 17330 3290 17354 3292
rect 17410 3290 17434 3292
rect 17490 3290 17496 3292
rect 17250 3238 17252 3290
rect 17432 3238 17434 3290
rect 17188 3236 17194 3238
rect 17250 3236 17274 3238
rect 17330 3236 17354 3238
rect 17410 3236 17434 3238
rect 17490 3236 17496 3238
rect 17188 3227 17496 3236
rect 17604 3194 17632 3470
rect 17684 3392 17736 3398
rect 17684 3334 17736 3340
rect 17592 3188 17644 3194
rect 17592 3130 17644 3136
rect 17696 3074 17724 3334
rect 18708 3194 18736 3946
rect 19340 3732 19392 3738
rect 19340 3674 19392 3680
rect 19352 3210 19380 3674
rect 19444 3398 19472 4422
rect 19720 3738 19748 4626
rect 19800 3936 19852 3942
rect 19800 3878 19852 3884
rect 19812 3738 19840 3878
rect 19708 3732 19760 3738
rect 19708 3674 19760 3680
rect 19800 3732 19852 3738
rect 19800 3674 19852 3680
rect 19524 3460 19576 3466
rect 19524 3402 19576 3408
rect 19432 3392 19484 3398
rect 19432 3334 19484 3340
rect 18696 3188 18748 3194
rect 18696 3130 18748 3136
rect 19260 3182 19380 3210
rect 17604 3046 17724 3074
rect 17604 2582 17632 3046
rect 18144 2984 18196 2990
rect 18328 2984 18380 2990
rect 18196 2944 18276 2972
rect 18144 2926 18196 2932
rect 17684 2848 17736 2854
rect 17684 2790 17736 2796
rect 18144 2848 18196 2854
rect 18144 2790 18196 2796
rect 17592 2576 17644 2582
rect 17592 2518 17644 2524
rect 17188 2204 17496 2213
rect 17188 2202 17194 2204
rect 17250 2202 17274 2204
rect 17330 2202 17354 2204
rect 17410 2202 17434 2204
rect 17490 2202 17496 2204
rect 17250 2150 17252 2202
rect 17432 2150 17434 2202
rect 17188 2148 17194 2150
rect 17250 2148 17274 2150
rect 17330 2148 17354 2150
rect 17410 2148 17434 2150
rect 17490 2148 17496 2150
rect 17188 2139 17496 2148
rect 17696 1902 17724 2790
rect 18156 2446 18184 2790
rect 18248 2514 18276 2944
rect 18328 2926 18380 2932
rect 18340 2582 18368 2926
rect 18708 2922 18736 3130
rect 19260 3126 19288 3182
rect 19248 3120 19300 3126
rect 19248 3062 19300 3068
rect 19340 3120 19392 3126
rect 19340 3062 19392 3068
rect 19352 2938 19380 3062
rect 19536 2938 19564 3402
rect 19708 3392 19760 3398
rect 19708 3334 19760 3340
rect 19720 2990 19748 3334
rect 19904 3126 19932 6870
rect 19984 6656 20036 6662
rect 19984 6598 20036 6604
rect 19996 6458 20024 6598
rect 19984 6452 20036 6458
rect 19984 6394 20036 6400
rect 19984 5364 20036 5370
rect 19984 5306 20036 5312
rect 19996 4078 20024 5306
rect 20364 5166 20392 7142
rect 20456 6934 20484 7686
rect 20546 7100 20854 7109
rect 20546 7098 20552 7100
rect 20608 7098 20632 7100
rect 20688 7098 20712 7100
rect 20768 7098 20792 7100
rect 20848 7098 20854 7100
rect 20608 7046 20610 7098
rect 20790 7046 20792 7098
rect 20546 7044 20552 7046
rect 20608 7044 20632 7046
rect 20688 7044 20712 7046
rect 20768 7044 20792 7046
rect 20848 7044 20854 7046
rect 20546 7035 20854 7044
rect 20444 6928 20496 6934
rect 20444 6870 20496 6876
rect 21008 6458 21036 9318
rect 21088 8832 21140 8838
rect 21088 8774 21140 8780
rect 21100 6730 21128 8774
rect 21192 6798 21220 10134
rect 21284 9450 21312 10202
rect 21928 9450 21956 10542
rect 22100 10124 22152 10130
rect 22100 10066 22152 10072
rect 22112 9654 22140 10066
rect 22100 9648 22152 9654
rect 22100 9590 22152 9596
rect 22204 9518 22232 10542
rect 22192 9512 22244 9518
rect 22192 9454 22244 9460
rect 21272 9444 21324 9450
rect 21272 9386 21324 9392
rect 21916 9444 21968 9450
rect 21916 9386 21968 9392
rect 21824 8628 21876 8634
rect 21824 8570 21876 8576
rect 21640 8424 21692 8430
rect 21640 8366 21692 8372
rect 21652 8294 21680 8366
rect 21640 8288 21692 8294
rect 21640 8230 21692 8236
rect 21652 7954 21680 8230
rect 21836 8090 21864 8570
rect 21928 8294 21956 9386
rect 22296 8974 22324 10610
rect 22652 9036 22704 9042
rect 22652 8978 22704 8984
rect 22284 8968 22336 8974
rect 22284 8910 22336 8916
rect 22008 8832 22060 8838
rect 22008 8774 22060 8780
rect 22020 8566 22048 8774
rect 22008 8560 22060 8566
rect 22008 8502 22060 8508
rect 22020 8430 22048 8502
rect 22100 8492 22152 8498
rect 22100 8434 22152 8440
rect 22008 8424 22060 8430
rect 22008 8366 22060 8372
rect 21916 8288 21968 8294
rect 21916 8230 21968 8236
rect 21824 8084 21876 8090
rect 21824 8026 21876 8032
rect 21640 7948 21692 7954
rect 21640 7890 21692 7896
rect 21916 7948 21968 7954
rect 22020 7936 22048 8366
rect 22112 8090 22140 8434
rect 22664 8090 22692 8978
rect 22100 8084 22152 8090
rect 22100 8026 22152 8032
rect 22652 8084 22704 8090
rect 22652 8026 22704 8032
rect 22756 7954 22784 14010
rect 22848 13870 22876 14894
rect 23020 14816 23072 14822
rect 23020 14758 23072 14764
rect 23032 14618 23060 14758
rect 23020 14612 23072 14618
rect 23020 14554 23072 14560
rect 23020 14476 23072 14482
rect 23020 14418 23072 14424
rect 23204 14476 23256 14482
rect 23204 14418 23256 14424
rect 22836 13864 22888 13870
rect 22836 13806 22888 13812
rect 22848 13530 22876 13806
rect 22928 13728 22980 13734
rect 22928 13670 22980 13676
rect 22836 13524 22888 13530
rect 22836 13466 22888 13472
rect 22848 13258 22876 13466
rect 22940 13462 22968 13670
rect 23032 13530 23060 14418
rect 23216 14006 23244 14418
rect 23204 14000 23256 14006
rect 23204 13942 23256 13948
rect 23020 13524 23072 13530
rect 23020 13466 23072 13472
rect 22928 13456 22980 13462
rect 22928 13398 22980 13404
rect 23308 13394 23336 15014
rect 23400 14550 23428 16390
rect 23584 15910 23612 17750
rect 23768 17660 23796 24550
rect 24136 24052 24164 24686
rect 24320 24410 24348 24686
rect 24308 24404 24360 24410
rect 24308 24346 24360 24352
rect 24412 24206 24440 26454
rect 24504 25974 24532 27814
rect 24596 27674 24624 27882
rect 24584 27668 24636 27674
rect 24584 27610 24636 27616
rect 24688 27606 24716 29718
rect 24768 29096 24820 29102
rect 24768 29038 24820 29044
rect 24780 27946 24808 29038
rect 24768 27940 24820 27946
rect 24768 27882 24820 27888
rect 24676 27600 24728 27606
rect 24676 27542 24728 27548
rect 24780 27554 24808 27882
rect 24964 27713 24992 31600
rect 26436 30938 26464 31600
rect 27262 31036 27570 31045
rect 27262 31034 27268 31036
rect 27324 31034 27348 31036
rect 27404 31034 27428 31036
rect 27484 31034 27508 31036
rect 27564 31034 27570 31036
rect 27324 30982 27326 31034
rect 27506 30982 27508 31034
rect 27262 30980 27268 30982
rect 27324 30980 27348 30982
rect 27404 30980 27428 30982
rect 27484 30980 27508 30982
rect 27564 30980 27570 30982
rect 27262 30971 27570 30980
rect 26424 30932 26476 30938
rect 26424 30874 26476 30880
rect 26516 30592 26568 30598
rect 26516 30534 26568 30540
rect 26528 30394 26556 30534
rect 26516 30388 26568 30394
rect 26516 30330 26568 30336
rect 25228 30048 25280 30054
rect 25228 29990 25280 29996
rect 25240 29753 25268 29990
rect 27262 29948 27570 29957
rect 27262 29946 27268 29948
rect 27324 29946 27348 29948
rect 27404 29946 27428 29948
rect 27484 29946 27508 29948
rect 27564 29946 27570 29948
rect 27324 29894 27326 29946
rect 27506 29894 27508 29946
rect 27262 29892 27268 29894
rect 27324 29892 27348 29894
rect 27404 29892 27428 29894
rect 27484 29892 27508 29894
rect 27564 29892 27570 29894
rect 27262 29883 27570 29892
rect 25226 29744 25282 29753
rect 25226 29679 25282 29688
rect 25964 29708 26016 29714
rect 25240 29510 25268 29679
rect 25964 29650 26016 29656
rect 25686 29608 25742 29617
rect 25686 29543 25742 29552
rect 25228 29504 25280 29510
rect 25228 29446 25280 29452
rect 25320 29096 25372 29102
rect 25320 29038 25372 29044
rect 25332 28762 25360 29038
rect 25700 28762 25728 29543
rect 25320 28756 25372 28762
rect 25320 28698 25372 28704
rect 25688 28756 25740 28762
rect 25688 28698 25740 28704
rect 25044 28688 25096 28694
rect 25228 28688 25280 28694
rect 25096 28636 25176 28642
rect 25044 28630 25176 28636
rect 25228 28630 25280 28636
rect 25056 28614 25176 28630
rect 25148 28422 25176 28614
rect 25044 28416 25096 28422
rect 25044 28358 25096 28364
rect 25136 28416 25188 28422
rect 25136 28358 25188 28364
rect 25056 28218 25084 28358
rect 25044 28212 25096 28218
rect 25044 28154 25096 28160
rect 25240 28150 25268 28630
rect 25596 28620 25648 28626
rect 25596 28562 25648 28568
rect 25228 28144 25280 28150
rect 25228 28086 25280 28092
rect 25228 28008 25280 28014
rect 25228 27950 25280 27956
rect 24950 27704 25006 27713
rect 24950 27639 25006 27648
rect 24780 27538 24900 27554
rect 24584 27532 24636 27538
rect 24780 27532 24912 27538
rect 24780 27526 24860 27532
rect 24584 27474 24636 27480
rect 24860 27474 24912 27480
rect 24596 26246 24624 27474
rect 25240 27334 25268 27950
rect 25320 27940 25372 27946
rect 25320 27882 25372 27888
rect 25136 27328 25188 27334
rect 25136 27270 25188 27276
rect 25228 27328 25280 27334
rect 25228 27270 25280 27276
rect 24676 26920 24728 26926
rect 24676 26862 24728 26868
rect 24584 26240 24636 26246
rect 24584 26182 24636 26188
rect 24492 25968 24544 25974
rect 24492 25910 24544 25916
rect 24596 25838 24624 26182
rect 24584 25832 24636 25838
rect 24584 25774 24636 25780
rect 24492 25696 24544 25702
rect 24492 25638 24544 25644
rect 24504 25498 24532 25638
rect 24596 25498 24624 25774
rect 24492 25492 24544 25498
rect 24492 25434 24544 25440
rect 24584 25492 24636 25498
rect 24584 25434 24636 25440
rect 24688 25226 24716 26862
rect 24952 26512 25004 26518
rect 24952 26454 25004 26460
rect 24860 26376 24912 26382
rect 24860 26318 24912 26324
rect 24768 25968 24820 25974
rect 24768 25910 24820 25916
rect 24676 25220 24728 25226
rect 24676 25162 24728 25168
rect 24400 24200 24452 24206
rect 24400 24142 24452 24148
rect 24584 24064 24636 24070
rect 24136 24024 24348 24052
rect 23904 23964 24212 23973
rect 23904 23962 23910 23964
rect 23966 23962 23990 23964
rect 24046 23962 24070 23964
rect 24126 23962 24150 23964
rect 24206 23962 24212 23964
rect 23966 23910 23968 23962
rect 24148 23910 24150 23962
rect 23904 23908 23910 23910
rect 23966 23908 23990 23910
rect 24046 23908 24070 23910
rect 24126 23908 24150 23910
rect 24206 23908 24212 23910
rect 23904 23899 24212 23908
rect 23904 22876 24212 22885
rect 23904 22874 23910 22876
rect 23966 22874 23990 22876
rect 24046 22874 24070 22876
rect 24126 22874 24150 22876
rect 24206 22874 24212 22876
rect 23966 22822 23968 22874
rect 24148 22822 24150 22874
rect 23904 22820 23910 22822
rect 23966 22820 23990 22822
rect 24046 22820 24070 22822
rect 24126 22820 24150 22822
rect 24206 22820 24212 22822
rect 23904 22811 24212 22820
rect 23904 21788 24212 21797
rect 23904 21786 23910 21788
rect 23966 21786 23990 21788
rect 24046 21786 24070 21788
rect 24126 21786 24150 21788
rect 24206 21786 24212 21788
rect 23966 21734 23968 21786
rect 24148 21734 24150 21786
rect 23904 21732 23910 21734
rect 23966 21732 23990 21734
rect 24046 21732 24070 21734
rect 24126 21732 24150 21734
rect 24206 21732 24212 21734
rect 23904 21723 24212 21732
rect 24032 21548 24084 21554
rect 24032 21490 24084 21496
rect 23848 21480 23900 21486
rect 23848 21422 23900 21428
rect 23860 21146 23888 21422
rect 24044 21146 24072 21490
rect 23848 21140 23900 21146
rect 23848 21082 23900 21088
rect 24032 21140 24084 21146
rect 24032 21082 24084 21088
rect 23904 20700 24212 20709
rect 23904 20698 23910 20700
rect 23966 20698 23990 20700
rect 24046 20698 24070 20700
rect 24126 20698 24150 20700
rect 24206 20698 24212 20700
rect 23966 20646 23968 20698
rect 24148 20646 24150 20698
rect 23904 20644 23910 20646
rect 23966 20644 23990 20646
rect 24046 20644 24070 20646
rect 24126 20644 24150 20646
rect 24206 20644 24212 20646
rect 23904 20635 24212 20644
rect 23904 19612 24212 19621
rect 23904 19610 23910 19612
rect 23966 19610 23990 19612
rect 24046 19610 24070 19612
rect 24126 19610 24150 19612
rect 24206 19610 24212 19612
rect 23966 19558 23968 19610
rect 24148 19558 24150 19610
rect 23904 19556 23910 19558
rect 23966 19556 23990 19558
rect 24046 19556 24070 19558
rect 24126 19556 24150 19558
rect 24206 19556 24212 19558
rect 23904 19547 24212 19556
rect 24032 19304 24084 19310
rect 24032 19246 24084 19252
rect 24044 18970 24072 19246
rect 24032 18964 24084 18970
rect 24032 18906 24084 18912
rect 24320 18834 24348 24024
rect 24584 24006 24636 24012
rect 24492 23656 24544 23662
rect 24492 23598 24544 23604
rect 24400 23588 24452 23594
rect 24400 23530 24452 23536
rect 24412 23322 24440 23530
rect 24504 23322 24532 23598
rect 24400 23316 24452 23322
rect 24400 23258 24452 23264
rect 24492 23316 24544 23322
rect 24492 23258 24544 23264
rect 24596 23254 24624 24006
rect 24688 23746 24716 25162
rect 24780 24954 24808 25910
rect 24768 24948 24820 24954
rect 24768 24890 24820 24896
rect 24768 24676 24820 24682
rect 24768 24618 24820 24624
rect 24780 24342 24808 24618
rect 24872 24410 24900 26318
rect 24964 26042 24992 26454
rect 25148 26450 25176 27270
rect 25240 26450 25268 27270
rect 25332 26858 25360 27882
rect 25608 27878 25636 28562
rect 25504 27872 25556 27878
rect 25504 27814 25556 27820
rect 25596 27872 25648 27878
rect 25596 27814 25648 27820
rect 25516 27674 25544 27814
rect 25504 27668 25556 27674
rect 25504 27610 25556 27616
rect 25608 27606 25636 27814
rect 25596 27600 25648 27606
rect 25596 27542 25648 27548
rect 25700 27538 25728 28698
rect 25872 28620 25924 28626
rect 25872 28562 25924 28568
rect 25780 28416 25832 28422
rect 25780 28358 25832 28364
rect 25792 27538 25820 28358
rect 25884 28218 25912 28562
rect 25872 28212 25924 28218
rect 25872 28154 25924 28160
rect 25688 27532 25740 27538
rect 25688 27474 25740 27480
rect 25780 27532 25832 27538
rect 25780 27474 25832 27480
rect 25320 26852 25372 26858
rect 25320 26794 25372 26800
rect 25136 26444 25188 26450
rect 25136 26386 25188 26392
rect 25228 26444 25280 26450
rect 25228 26386 25280 26392
rect 24952 26036 25004 26042
rect 24952 25978 25004 25984
rect 25240 25838 25268 26386
rect 25228 25832 25280 25838
rect 25228 25774 25280 25780
rect 24860 24404 24912 24410
rect 24860 24346 24912 24352
rect 24768 24336 24820 24342
rect 24768 24278 24820 24284
rect 24780 23866 24808 24278
rect 25044 24200 25096 24206
rect 25044 24142 25096 24148
rect 24768 23860 24820 23866
rect 24768 23802 24820 23808
rect 24688 23718 24808 23746
rect 24584 23248 24636 23254
rect 24584 23190 24636 23196
rect 24400 23180 24452 23186
rect 24400 23122 24452 23128
rect 24412 22710 24440 23122
rect 24492 23112 24544 23118
rect 24492 23054 24544 23060
rect 24676 23112 24728 23118
rect 24676 23054 24728 23060
rect 24400 22704 24452 22710
rect 24400 22646 24452 22652
rect 24412 22098 24440 22646
rect 24504 22438 24532 23054
rect 24584 22568 24636 22574
rect 24584 22510 24636 22516
rect 24492 22432 24544 22438
rect 24492 22374 24544 22380
rect 24492 22228 24544 22234
rect 24492 22170 24544 22176
rect 24400 22092 24452 22098
rect 24400 22034 24452 22040
rect 24400 21956 24452 21962
rect 24400 21898 24452 21904
rect 24412 21486 24440 21898
rect 24400 21480 24452 21486
rect 24400 21422 24452 21428
rect 24504 19310 24532 22170
rect 24596 20874 24624 22510
rect 24688 22506 24716 23054
rect 24676 22500 24728 22506
rect 24676 22442 24728 22448
rect 24688 21690 24716 22442
rect 24676 21684 24728 21690
rect 24676 21626 24728 21632
rect 24584 20868 24636 20874
rect 24584 20810 24636 20816
rect 24780 19334 24808 23718
rect 24952 23656 25004 23662
rect 24952 23598 25004 23604
rect 24964 23254 24992 23598
rect 24952 23248 25004 23254
rect 24952 23190 25004 23196
rect 24964 22778 24992 23190
rect 25056 22982 25084 24142
rect 25136 23180 25188 23186
rect 25136 23122 25188 23128
rect 25044 22976 25096 22982
rect 25044 22918 25096 22924
rect 24952 22772 25004 22778
rect 24952 22714 25004 22720
rect 24860 22704 24912 22710
rect 24860 22646 24912 22652
rect 24872 22574 24900 22646
rect 24860 22568 24912 22574
rect 24860 22510 24912 22516
rect 25148 21690 25176 23122
rect 25136 21684 25188 21690
rect 25136 21626 25188 21632
rect 25148 21078 25176 21626
rect 25332 21486 25360 26794
rect 25976 26518 26004 29650
rect 26424 29028 26476 29034
rect 26424 28970 26476 28976
rect 26240 28960 26292 28966
rect 26240 28902 26292 28908
rect 26056 28416 26108 28422
rect 26056 28358 26108 28364
rect 26068 28218 26096 28358
rect 26056 28212 26108 28218
rect 26056 28154 26108 28160
rect 26252 28014 26280 28902
rect 26436 28626 26464 28970
rect 27262 28860 27570 28869
rect 27262 28858 27268 28860
rect 27324 28858 27348 28860
rect 27404 28858 27428 28860
rect 27484 28858 27508 28860
rect 27564 28858 27570 28860
rect 27324 28806 27326 28858
rect 27506 28806 27508 28858
rect 27262 28804 27268 28806
rect 27324 28804 27348 28806
rect 27404 28804 27428 28806
rect 27484 28804 27508 28806
rect 27564 28804 27570 28806
rect 27262 28795 27570 28804
rect 26424 28620 26476 28626
rect 26424 28562 26476 28568
rect 26240 28008 26292 28014
rect 26240 27950 26292 27956
rect 26252 26790 26280 27950
rect 27262 27772 27570 27781
rect 27262 27770 27268 27772
rect 27324 27770 27348 27772
rect 27404 27770 27428 27772
rect 27484 27770 27508 27772
rect 27564 27770 27570 27772
rect 27324 27718 27326 27770
rect 27506 27718 27508 27770
rect 27262 27716 27268 27718
rect 27324 27716 27348 27718
rect 27404 27716 27428 27718
rect 27484 27716 27508 27718
rect 27564 27716 27570 27718
rect 27262 27707 27570 27716
rect 26240 26784 26292 26790
rect 26240 26726 26292 26732
rect 25964 26512 26016 26518
rect 25964 26454 26016 26460
rect 25412 26240 25464 26246
rect 25412 26182 25464 26188
rect 25504 26240 25556 26246
rect 25504 26182 25556 26188
rect 25424 26042 25452 26182
rect 25412 26036 25464 26042
rect 25412 25978 25464 25984
rect 25412 25832 25464 25838
rect 25516 25786 25544 26182
rect 25976 26042 26004 26454
rect 26148 26376 26200 26382
rect 26148 26318 26200 26324
rect 26056 26240 26108 26246
rect 26056 26182 26108 26188
rect 25964 26036 26016 26042
rect 25964 25978 26016 25984
rect 25464 25780 25544 25786
rect 25412 25774 25544 25780
rect 25424 25758 25544 25774
rect 25424 24886 25452 25758
rect 25504 25696 25556 25702
rect 25504 25638 25556 25644
rect 25596 25696 25648 25702
rect 25596 25638 25648 25644
rect 25516 25158 25544 25638
rect 25608 25498 25636 25638
rect 25596 25492 25648 25498
rect 25596 25434 25648 25440
rect 25976 25276 26004 25978
rect 26068 25430 26096 26182
rect 26160 25430 26188 26318
rect 26252 25838 26280 26726
rect 27262 26684 27570 26693
rect 27262 26682 27268 26684
rect 27324 26682 27348 26684
rect 27404 26682 27428 26684
rect 27484 26682 27508 26684
rect 27564 26682 27570 26684
rect 27324 26630 27326 26682
rect 27506 26630 27508 26682
rect 27262 26628 27268 26630
rect 27324 26628 27348 26630
rect 27404 26628 27428 26630
rect 27484 26628 27508 26630
rect 27564 26628 27570 26630
rect 27262 26619 27570 26628
rect 26240 25832 26292 25838
rect 26240 25774 26292 25780
rect 26056 25424 26108 25430
rect 26056 25366 26108 25372
rect 26148 25424 26200 25430
rect 26148 25366 26200 25372
rect 26252 25362 26280 25774
rect 26792 25764 26844 25770
rect 26792 25706 26844 25712
rect 26804 25498 26832 25706
rect 27262 25596 27570 25605
rect 27262 25594 27268 25596
rect 27324 25594 27348 25596
rect 27404 25594 27428 25596
rect 27484 25594 27508 25596
rect 27564 25594 27570 25596
rect 27324 25542 27326 25594
rect 27506 25542 27508 25594
rect 27262 25540 27268 25542
rect 27324 25540 27348 25542
rect 27404 25540 27428 25542
rect 27484 25540 27508 25542
rect 27564 25540 27570 25542
rect 27262 25531 27570 25540
rect 26792 25492 26844 25498
rect 26792 25434 26844 25440
rect 26240 25356 26292 25362
rect 26240 25298 26292 25304
rect 26332 25356 26384 25362
rect 26332 25298 26384 25304
rect 25976 25248 26096 25276
rect 25504 25152 25556 25158
rect 25504 25094 25556 25100
rect 25872 24948 25924 24954
rect 25872 24890 25924 24896
rect 25412 24880 25464 24886
rect 25412 24822 25464 24828
rect 25504 24744 25556 24750
rect 25504 24686 25556 24692
rect 25412 24676 25464 24682
rect 25412 24618 25464 24624
rect 25424 24410 25452 24618
rect 25412 24404 25464 24410
rect 25412 24346 25464 24352
rect 25516 23662 25544 24686
rect 25504 23656 25556 23662
rect 25504 23598 25556 23604
rect 25780 23656 25832 23662
rect 25884 23644 25912 24890
rect 25976 24070 26004 25248
rect 26068 25242 26096 25248
rect 26344 25242 26372 25298
rect 26068 25214 26372 25242
rect 26424 24608 26476 24614
rect 26424 24550 26476 24556
rect 26976 24608 27028 24614
rect 26976 24550 27028 24556
rect 26436 24410 26464 24550
rect 26988 24410 27016 24550
rect 27262 24508 27570 24517
rect 27262 24506 27268 24508
rect 27324 24506 27348 24508
rect 27404 24506 27428 24508
rect 27484 24506 27508 24508
rect 27564 24506 27570 24508
rect 27324 24454 27326 24506
rect 27506 24454 27508 24506
rect 27262 24452 27268 24454
rect 27324 24452 27348 24454
rect 27404 24452 27428 24454
rect 27484 24452 27508 24454
rect 27564 24452 27570 24454
rect 27262 24443 27570 24452
rect 26424 24404 26476 24410
rect 26424 24346 26476 24352
rect 26976 24404 27028 24410
rect 26976 24346 27028 24352
rect 26240 24268 26292 24274
rect 26240 24210 26292 24216
rect 25964 24064 26016 24070
rect 25964 24006 26016 24012
rect 26056 24064 26108 24070
rect 26056 24006 26108 24012
rect 25832 23616 25912 23644
rect 25780 23598 25832 23604
rect 25412 22976 25464 22982
rect 25412 22918 25464 22924
rect 25424 22574 25452 22918
rect 25516 22642 25544 23598
rect 25596 23588 25648 23594
rect 25596 23530 25648 23536
rect 25608 22778 25636 23530
rect 25884 23254 25912 23616
rect 26068 23322 26096 24006
rect 26252 23526 26280 24210
rect 26424 24064 26476 24070
rect 26424 24006 26476 24012
rect 26240 23520 26292 23526
rect 26240 23462 26292 23468
rect 26252 23322 26280 23462
rect 26056 23316 26108 23322
rect 26056 23258 26108 23264
rect 26240 23316 26292 23322
rect 26240 23258 26292 23264
rect 25872 23248 25924 23254
rect 25872 23190 25924 23196
rect 25688 23112 25740 23118
rect 25688 23054 25740 23060
rect 25700 22778 25728 23054
rect 25596 22772 25648 22778
rect 25596 22714 25648 22720
rect 25688 22772 25740 22778
rect 25688 22714 25740 22720
rect 25504 22636 25556 22642
rect 25504 22578 25556 22584
rect 25412 22568 25464 22574
rect 25412 22510 25464 22516
rect 25504 22024 25556 22030
rect 25504 21966 25556 21972
rect 25516 21690 25544 21966
rect 25700 21690 25728 22714
rect 25884 22166 25912 23190
rect 25872 22160 25924 22166
rect 25872 22102 25924 22108
rect 26068 22094 26096 23258
rect 26436 23186 26464 24006
rect 27262 23420 27570 23429
rect 27262 23418 27268 23420
rect 27324 23418 27348 23420
rect 27404 23418 27428 23420
rect 27484 23418 27508 23420
rect 27564 23418 27570 23420
rect 27324 23366 27326 23418
rect 27506 23366 27508 23418
rect 27262 23364 27268 23366
rect 27324 23364 27348 23366
rect 27404 23364 27428 23366
rect 27484 23364 27508 23366
rect 27564 23364 27570 23366
rect 27262 23355 27570 23364
rect 26424 23180 26476 23186
rect 26424 23122 26476 23128
rect 26148 22976 26200 22982
rect 26148 22918 26200 22924
rect 26976 22976 27028 22982
rect 26976 22918 27028 22924
rect 26160 22506 26188 22918
rect 26516 22568 26568 22574
rect 26988 22522 27016 22918
rect 26516 22510 26568 22516
rect 26148 22500 26200 22506
rect 26148 22442 26200 22448
rect 26068 22066 26188 22094
rect 25872 21888 25924 21894
rect 25872 21830 25924 21836
rect 25504 21684 25556 21690
rect 25504 21626 25556 21632
rect 25688 21684 25740 21690
rect 25688 21626 25740 21632
rect 25320 21480 25372 21486
rect 25320 21422 25372 21428
rect 25136 21072 25188 21078
rect 25136 21014 25188 21020
rect 25332 19990 25360 21422
rect 25516 21146 25544 21626
rect 25884 21146 25912 21830
rect 25504 21140 25556 21146
rect 25504 21082 25556 21088
rect 25872 21140 25924 21146
rect 25872 21082 25924 21088
rect 26160 21078 26188 22066
rect 26424 21888 26476 21894
rect 26424 21830 26476 21836
rect 26436 21146 26464 21830
rect 26528 21690 26556 22510
rect 26792 22500 26844 22506
rect 26792 22442 26844 22448
rect 26896 22494 27016 22522
rect 26804 22234 26832 22442
rect 26792 22228 26844 22234
rect 26792 22170 26844 22176
rect 26516 21684 26568 21690
rect 26516 21626 26568 21632
rect 26424 21140 26476 21146
rect 26424 21082 26476 21088
rect 26148 21072 26200 21078
rect 26148 21014 26200 21020
rect 26528 21010 26556 21626
rect 26516 21004 26568 21010
rect 26516 20946 26568 20952
rect 26700 21004 26752 21010
rect 26896 20992 26924 22494
rect 27262 22332 27570 22341
rect 27262 22330 27268 22332
rect 27324 22330 27348 22332
rect 27404 22330 27428 22332
rect 27484 22330 27508 22332
rect 27564 22330 27570 22332
rect 27324 22278 27326 22330
rect 27506 22278 27508 22330
rect 27262 22276 27268 22278
rect 27324 22276 27348 22278
rect 27404 22276 27428 22278
rect 27484 22276 27508 22278
rect 27564 22276 27570 22278
rect 27262 22267 27570 22276
rect 26976 22160 27028 22166
rect 26976 22102 27028 22108
rect 26988 21146 27016 22102
rect 27262 21244 27570 21253
rect 27262 21242 27268 21244
rect 27324 21242 27348 21244
rect 27404 21242 27428 21244
rect 27484 21242 27508 21244
rect 27564 21242 27570 21244
rect 27324 21190 27326 21242
rect 27506 21190 27508 21242
rect 27262 21188 27268 21190
rect 27324 21188 27348 21190
rect 27404 21188 27428 21190
rect 27484 21188 27508 21190
rect 27564 21188 27570 21190
rect 27262 21179 27570 21188
rect 26976 21140 27028 21146
rect 26976 21082 27028 21088
rect 26976 21004 27028 21010
rect 26752 20964 26976 20992
rect 26700 20946 26752 20952
rect 26976 20946 27028 20952
rect 26528 20398 26556 20946
rect 26240 20392 26292 20398
rect 26240 20334 26292 20340
rect 26516 20392 26568 20398
rect 26516 20334 26568 20340
rect 25596 20324 25648 20330
rect 25596 20266 25648 20272
rect 25320 19984 25372 19990
rect 25320 19926 25372 19932
rect 25504 19712 25556 19718
rect 25504 19654 25556 19660
rect 24492 19304 24544 19310
rect 24688 19306 24808 19334
rect 24688 19258 24716 19306
rect 24492 19246 24544 19252
rect 24596 19230 24716 19258
rect 25228 19304 25280 19310
rect 25228 19246 25280 19252
rect 24308 18828 24360 18834
rect 24308 18770 24360 18776
rect 23904 18524 24212 18533
rect 23904 18522 23910 18524
rect 23966 18522 23990 18524
rect 24046 18522 24070 18524
rect 24126 18522 24150 18524
rect 24206 18522 24212 18524
rect 23966 18470 23968 18522
rect 24148 18470 24150 18522
rect 23904 18468 23910 18470
rect 23966 18468 23990 18470
rect 24046 18468 24070 18470
rect 24126 18468 24150 18470
rect 24206 18468 24212 18470
rect 23904 18459 24212 18468
rect 24124 18420 24176 18426
rect 24124 18362 24176 18368
rect 24136 18222 24164 18362
rect 24320 18358 24348 18770
rect 24492 18760 24544 18766
rect 24492 18702 24544 18708
rect 24504 18358 24532 18702
rect 24308 18352 24360 18358
rect 24308 18294 24360 18300
rect 24492 18352 24544 18358
rect 24492 18294 24544 18300
rect 24124 18216 24176 18222
rect 24124 18158 24176 18164
rect 24308 17808 24360 17814
rect 24308 17750 24360 17756
rect 23676 17632 23796 17660
rect 23572 15904 23624 15910
rect 23572 15846 23624 15852
rect 23480 15564 23532 15570
rect 23480 15506 23532 15512
rect 23492 14958 23520 15506
rect 23572 15360 23624 15366
rect 23572 15302 23624 15308
rect 23480 14952 23532 14958
rect 23480 14894 23532 14900
rect 23388 14544 23440 14550
rect 23388 14486 23440 14492
rect 23480 13728 23532 13734
rect 23480 13670 23532 13676
rect 23492 13394 23520 13670
rect 23296 13388 23348 13394
rect 23296 13330 23348 13336
rect 23480 13388 23532 13394
rect 23480 13330 23532 13336
rect 23112 13320 23164 13326
rect 23112 13262 23164 13268
rect 22836 13252 22888 13258
rect 22836 13194 22888 13200
rect 23124 12986 23152 13262
rect 23584 13190 23612 15302
rect 23676 15026 23704 17632
rect 23756 17536 23808 17542
rect 23756 17478 23808 17484
rect 23768 16726 23796 17478
rect 23904 17436 24212 17445
rect 23904 17434 23910 17436
rect 23966 17434 23990 17436
rect 24046 17434 24070 17436
rect 24126 17434 24150 17436
rect 24206 17434 24212 17436
rect 23966 17382 23968 17434
rect 24148 17382 24150 17434
rect 23904 17380 23910 17382
rect 23966 17380 23990 17382
rect 24046 17380 24070 17382
rect 24126 17380 24150 17382
rect 24206 17380 24212 17382
rect 23904 17371 24212 17380
rect 23940 17264 23992 17270
rect 23938 17232 23940 17241
rect 23992 17232 23994 17241
rect 23938 17167 23994 17176
rect 24124 16992 24176 16998
rect 24216 16992 24268 16998
rect 24124 16934 24176 16940
rect 24214 16960 24216 16969
rect 24268 16960 24270 16969
rect 23756 16720 23808 16726
rect 23756 16662 23808 16668
rect 24136 16658 24164 16934
rect 24214 16895 24270 16904
rect 24320 16794 24348 17750
rect 24492 17672 24544 17678
rect 24492 17614 24544 17620
rect 24400 17536 24452 17542
rect 24400 17478 24452 17484
rect 24412 17338 24440 17478
rect 24400 17332 24452 17338
rect 24400 17274 24452 17280
rect 24504 17082 24532 17614
rect 24412 17054 24532 17082
rect 24412 16998 24440 17054
rect 24400 16992 24452 16998
rect 24400 16934 24452 16940
rect 24308 16788 24360 16794
rect 24308 16730 24360 16736
rect 24124 16652 24176 16658
rect 24124 16594 24176 16600
rect 24596 16590 24624 19230
rect 24676 19168 24728 19174
rect 24676 19110 24728 19116
rect 24860 19168 24912 19174
rect 24860 19110 24912 19116
rect 24688 18970 24716 19110
rect 24676 18964 24728 18970
rect 24676 18906 24728 18912
rect 24872 18902 24900 19110
rect 24860 18896 24912 18902
rect 24860 18838 24912 18844
rect 24860 18692 24912 18698
rect 24860 18634 24912 18640
rect 24768 18624 24820 18630
rect 24768 18566 24820 18572
rect 24676 17740 24728 17746
rect 24676 17682 24728 17688
rect 24688 16969 24716 17682
rect 24674 16960 24730 16969
rect 24674 16895 24730 16904
rect 24780 16794 24808 18566
rect 24872 17814 24900 18634
rect 25044 18080 25096 18086
rect 25044 18022 25096 18028
rect 25056 17814 25084 18022
rect 25240 17814 25268 19246
rect 25412 18624 25464 18630
rect 25412 18566 25464 18572
rect 25424 18426 25452 18566
rect 25412 18420 25464 18426
rect 25412 18362 25464 18368
rect 24860 17808 24912 17814
rect 24860 17750 24912 17756
rect 25044 17808 25096 17814
rect 25044 17750 25096 17756
rect 25228 17808 25280 17814
rect 25228 17750 25280 17756
rect 24860 17604 24912 17610
rect 24860 17546 24912 17552
rect 24872 17202 24900 17546
rect 25136 17536 25188 17542
rect 25136 17478 25188 17484
rect 24950 17232 25006 17241
rect 24860 17196 24912 17202
rect 25006 17190 25084 17218
rect 24950 17167 25006 17176
rect 24860 17138 24912 17144
rect 25056 17134 25084 17190
rect 25044 17128 25096 17134
rect 25044 17070 25096 17076
rect 24952 17060 25004 17066
rect 24952 17002 25004 17008
rect 24964 16794 24992 17002
rect 25044 16992 25096 16998
rect 25044 16934 25096 16940
rect 24768 16788 24820 16794
rect 24768 16730 24820 16736
rect 24952 16788 25004 16794
rect 24952 16730 25004 16736
rect 24308 16584 24360 16590
rect 24308 16526 24360 16532
rect 24584 16584 24636 16590
rect 24584 16526 24636 16532
rect 23904 16348 24212 16357
rect 23904 16346 23910 16348
rect 23966 16346 23990 16348
rect 24046 16346 24070 16348
rect 24126 16346 24150 16348
rect 24206 16346 24212 16348
rect 23966 16294 23968 16346
rect 24148 16294 24150 16346
rect 23904 16292 23910 16294
rect 23966 16292 23990 16294
rect 24046 16292 24070 16294
rect 24126 16292 24150 16294
rect 24206 16292 24212 16294
rect 23904 16283 24212 16292
rect 23756 16040 23808 16046
rect 23756 15982 23808 15988
rect 24124 16040 24176 16046
rect 24124 15982 24176 15988
rect 23768 15570 23796 15982
rect 24136 15638 24164 15982
rect 24320 15638 24348 16526
rect 24596 15722 24624 16526
rect 24780 16046 24808 16730
rect 24964 16658 24992 16730
rect 25056 16658 25084 16934
rect 25148 16794 25176 17478
rect 25516 17202 25544 19654
rect 25608 19514 25636 20266
rect 25596 19508 25648 19514
rect 25596 19450 25648 19456
rect 26252 19310 26280 20334
rect 27068 20256 27120 20262
rect 27068 20198 27120 20204
rect 27080 19922 27108 20198
rect 27262 20156 27570 20165
rect 27262 20154 27268 20156
rect 27324 20154 27348 20156
rect 27404 20154 27428 20156
rect 27484 20154 27508 20156
rect 27564 20154 27570 20156
rect 27324 20102 27326 20154
rect 27506 20102 27508 20154
rect 27262 20100 27268 20102
rect 27324 20100 27348 20102
rect 27404 20100 27428 20102
rect 27484 20100 27508 20102
rect 27564 20100 27570 20102
rect 27262 20091 27570 20100
rect 27068 19916 27120 19922
rect 27068 19858 27120 19864
rect 26424 19712 26476 19718
rect 26424 19654 26476 19660
rect 25780 19304 25832 19310
rect 25780 19246 25832 19252
rect 26240 19304 26292 19310
rect 26240 19246 26292 19252
rect 25792 18222 25820 19246
rect 25872 19236 25924 19242
rect 25872 19178 25924 19184
rect 25884 18970 25912 19178
rect 26436 19174 26464 19654
rect 26424 19168 26476 19174
rect 26424 19110 26476 19116
rect 25872 18964 25924 18970
rect 25872 18906 25924 18912
rect 27080 18766 27108 19858
rect 27262 19068 27570 19077
rect 27262 19066 27268 19068
rect 27324 19066 27348 19068
rect 27404 19066 27428 19068
rect 27484 19066 27508 19068
rect 27564 19066 27570 19068
rect 27324 19014 27326 19066
rect 27506 19014 27508 19066
rect 27262 19012 27268 19014
rect 27324 19012 27348 19014
rect 27404 19012 27428 19014
rect 27484 19012 27508 19014
rect 27564 19012 27570 19014
rect 27262 19003 27570 19012
rect 27068 18760 27120 18766
rect 27068 18702 27120 18708
rect 25780 18216 25832 18222
rect 25780 18158 25832 18164
rect 25964 18148 26016 18154
rect 25964 18090 26016 18096
rect 25976 17882 26004 18090
rect 27262 17980 27570 17989
rect 27262 17978 27268 17980
rect 27324 17978 27348 17980
rect 27404 17978 27428 17980
rect 27484 17978 27508 17980
rect 27564 17978 27570 17980
rect 27324 17926 27326 17978
rect 27506 17926 27508 17978
rect 27262 17924 27268 17926
rect 27324 17924 27348 17926
rect 27404 17924 27428 17926
rect 27484 17924 27508 17926
rect 27564 17924 27570 17926
rect 27262 17915 27570 17924
rect 25964 17876 26016 17882
rect 25964 17818 26016 17824
rect 25504 17196 25556 17202
rect 25504 17138 25556 17144
rect 25320 17128 25372 17134
rect 25320 17070 25372 17076
rect 25228 16992 25280 16998
rect 25228 16934 25280 16940
rect 25136 16788 25188 16794
rect 25136 16730 25188 16736
rect 24952 16652 25004 16658
rect 24952 16594 25004 16600
rect 25044 16652 25096 16658
rect 25044 16594 25096 16600
rect 25240 16454 25268 16934
rect 25228 16448 25280 16454
rect 25228 16390 25280 16396
rect 25332 16250 25360 17070
rect 25780 17060 25832 17066
rect 25780 17002 25832 17008
rect 25792 16794 25820 17002
rect 27262 16892 27570 16901
rect 27262 16890 27268 16892
rect 27324 16890 27348 16892
rect 27404 16890 27428 16892
rect 27484 16890 27508 16892
rect 27564 16890 27570 16892
rect 27324 16838 27326 16890
rect 27506 16838 27508 16890
rect 27262 16836 27268 16838
rect 27324 16836 27348 16838
rect 27404 16836 27428 16838
rect 27484 16836 27508 16838
rect 27564 16836 27570 16838
rect 27262 16827 27570 16836
rect 25780 16788 25832 16794
rect 25780 16730 25832 16736
rect 26240 16720 26292 16726
rect 26240 16662 26292 16668
rect 25320 16244 25372 16250
rect 25320 16186 25372 16192
rect 26252 16046 26280 16662
rect 24768 16040 24820 16046
rect 24768 15982 24820 15988
rect 26240 16040 26292 16046
rect 26240 15982 26292 15988
rect 26884 16040 26936 16046
rect 26884 15982 26936 15988
rect 24676 15904 24728 15910
rect 24676 15846 24728 15852
rect 24504 15694 24624 15722
rect 24124 15632 24176 15638
rect 24124 15574 24176 15580
rect 24308 15632 24360 15638
rect 24308 15574 24360 15580
rect 23756 15564 23808 15570
rect 23756 15506 23808 15512
rect 23904 15260 24212 15269
rect 23904 15258 23910 15260
rect 23966 15258 23990 15260
rect 24046 15258 24070 15260
rect 24126 15258 24150 15260
rect 24206 15258 24212 15260
rect 23966 15206 23968 15258
rect 24148 15206 24150 15258
rect 23904 15204 23910 15206
rect 23966 15204 23990 15206
rect 24046 15204 24070 15206
rect 24126 15204 24150 15206
rect 24206 15204 24212 15206
rect 23904 15195 24212 15204
rect 23664 15020 23716 15026
rect 23664 14962 23716 14968
rect 24320 14940 24348 15574
rect 24504 15570 24532 15694
rect 24584 15632 24636 15638
rect 24584 15574 24636 15580
rect 24492 15564 24544 15570
rect 24492 15506 24544 15512
rect 24596 14958 24624 15574
rect 24400 14952 24452 14958
rect 24320 14912 24400 14940
rect 24124 14816 24176 14822
rect 24124 14758 24176 14764
rect 24136 14618 24164 14758
rect 24320 14618 24348 14912
rect 24400 14894 24452 14900
rect 24584 14952 24636 14958
rect 24584 14894 24636 14900
rect 24400 14816 24452 14822
rect 24400 14758 24452 14764
rect 24124 14612 24176 14618
rect 24124 14554 24176 14560
rect 24308 14612 24360 14618
rect 24308 14554 24360 14560
rect 24412 14550 24440 14758
rect 24596 14618 24624 14894
rect 24688 14890 24716 15846
rect 25412 15564 25464 15570
rect 25412 15506 25464 15512
rect 24768 15360 24820 15366
rect 24768 15302 24820 15308
rect 24780 15162 24808 15302
rect 25424 15162 25452 15506
rect 26240 15360 26292 15366
rect 26240 15302 26292 15308
rect 24768 15156 24820 15162
rect 24768 15098 24820 15104
rect 25412 15156 25464 15162
rect 25412 15098 25464 15104
rect 26252 14958 26280 15302
rect 26896 14958 26924 15982
rect 27262 15804 27570 15813
rect 27262 15802 27268 15804
rect 27324 15802 27348 15804
rect 27404 15802 27428 15804
rect 27484 15802 27508 15804
rect 27564 15802 27570 15804
rect 27324 15750 27326 15802
rect 27506 15750 27508 15802
rect 27262 15748 27268 15750
rect 27324 15748 27348 15750
rect 27404 15748 27428 15750
rect 27484 15748 27508 15750
rect 27564 15748 27570 15750
rect 27262 15739 27570 15748
rect 26240 14952 26292 14958
rect 26240 14894 26292 14900
rect 26884 14952 26936 14958
rect 26884 14894 26936 14900
rect 24676 14884 24728 14890
rect 24676 14826 24728 14832
rect 24688 14618 24716 14826
rect 25228 14816 25280 14822
rect 25228 14758 25280 14764
rect 25240 14618 25268 14758
rect 24584 14612 24636 14618
rect 24584 14554 24636 14560
rect 24676 14612 24728 14618
rect 24676 14554 24728 14560
rect 25228 14612 25280 14618
rect 25228 14554 25280 14560
rect 24400 14544 24452 14550
rect 24400 14486 24452 14492
rect 25044 14476 25096 14482
rect 25044 14418 25096 14424
rect 24768 14340 24820 14346
rect 24768 14282 24820 14288
rect 24860 14340 24912 14346
rect 24860 14282 24912 14288
rect 23756 14272 23808 14278
rect 23756 14214 23808 14220
rect 23768 13938 23796 14214
rect 23904 14172 24212 14181
rect 23904 14170 23910 14172
rect 23966 14170 23990 14172
rect 24046 14170 24070 14172
rect 24126 14170 24150 14172
rect 24206 14170 24212 14172
rect 23966 14118 23968 14170
rect 24148 14118 24150 14170
rect 23904 14116 23910 14118
rect 23966 14116 23990 14118
rect 24046 14116 24070 14118
rect 24126 14116 24150 14118
rect 24206 14116 24212 14118
rect 23904 14107 24212 14116
rect 24216 14068 24268 14074
rect 24216 14010 24268 14016
rect 23848 14000 23900 14006
rect 23848 13942 23900 13948
rect 23756 13932 23808 13938
rect 23756 13874 23808 13880
rect 23664 13796 23716 13802
rect 23664 13738 23716 13744
rect 23676 13394 23704 13738
rect 23768 13394 23796 13874
rect 23860 13394 23888 13942
rect 24228 13870 24256 14010
rect 24780 13938 24808 14282
rect 24768 13932 24820 13938
rect 24596 13892 24768 13920
rect 24216 13864 24268 13870
rect 24216 13806 24268 13812
rect 24400 13796 24452 13802
rect 24400 13738 24452 13744
rect 23664 13388 23716 13394
rect 23664 13330 23716 13336
rect 23756 13388 23808 13394
rect 23756 13330 23808 13336
rect 23848 13388 23900 13394
rect 23848 13330 23900 13336
rect 23572 13184 23624 13190
rect 23572 13126 23624 13132
rect 23112 12980 23164 12986
rect 23112 12922 23164 12928
rect 23676 12782 23704 13330
rect 24412 13258 24440 13738
rect 24400 13252 24452 13258
rect 24400 13194 24452 13200
rect 24308 13184 24360 13190
rect 24308 13126 24360 13132
rect 23904 13084 24212 13093
rect 23904 13082 23910 13084
rect 23966 13082 23990 13084
rect 24046 13082 24070 13084
rect 24126 13082 24150 13084
rect 24206 13082 24212 13084
rect 23966 13030 23968 13082
rect 24148 13030 24150 13082
rect 23904 13028 23910 13030
rect 23966 13028 23990 13030
rect 24046 13028 24070 13030
rect 24126 13028 24150 13030
rect 24206 13028 24212 13030
rect 23904 13019 24212 13028
rect 23848 12980 23900 12986
rect 23848 12922 23900 12928
rect 23112 12776 23164 12782
rect 23112 12718 23164 12724
rect 23664 12776 23716 12782
rect 23664 12718 23716 12724
rect 23124 12442 23152 12718
rect 23388 12708 23440 12714
rect 23388 12650 23440 12656
rect 23572 12708 23624 12714
rect 23572 12650 23624 12656
rect 22928 12436 22980 12442
rect 22928 12378 22980 12384
rect 23112 12436 23164 12442
rect 23400 12434 23428 12650
rect 23584 12434 23612 12650
rect 23112 12378 23164 12384
rect 23308 12406 23428 12434
rect 23492 12406 23612 12434
rect 22836 12232 22888 12238
rect 22836 12174 22888 12180
rect 22848 11898 22876 12174
rect 22940 11898 22968 12378
rect 22836 11892 22888 11898
rect 22836 11834 22888 11840
rect 22928 11892 22980 11898
rect 22928 11834 22980 11840
rect 22848 11354 22876 11834
rect 23020 11620 23072 11626
rect 23020 11562 23072 11568
rect 22836 11348 22888 11354
rect 22836 11290 22888 11296
rect 23032 11218 23060 11562
rect 23308 11558 23336 12406
rect 23388 12096 23440 12102
rect 23388 12038 23440 12044
rect 23400 11762 23428 12038
rect 23492 11898 23520 12406
rect 23664 12368 23716 12374
rect 23664 12310 23716 12316
rect 23572 12232 23624 12238
rect 23572 12174 23624 12180
rect 23480 11892 23532 11898
rect 23480 11834 23532 11840
rect 23388 11756 23440 11762
rect 23388 11698 23440 11704
rect 23388 11620 23440 11626
rect 23388 11562 23440 11568
rect 23296 11552 23348 11558
rect 23296 11494 23348 11500
rect 23020 11212 23072 11218
rect 23020 11154 23072 11160
rect 23400 11082 23428 11562
rect 23492 11286 23520 11834
rect 23584 11830 23612 12174
rect 23572 11824 23624 11830
rect 23572 11766 23624 11772
rect 23572 11688 23624 11694
rect 23572 11630 23624 11636
rect 23584 11354 23612 11630
rect 23572 11348 23624 11354
rect 23572 11290 23624 11296
rect 23480 11280 23532 11286
rect 23480 11222 23532 11228
rect 23676 11150 23704 12310
rect 23860 12306 23888 12922
rect 24320 12918 24348 13126
rect 24308 12912 24360 12918
rect 24308 12854 24360 12860
rect 23848 12300 23900 12306
rect 23848 12242 23900 12248
rect 23756 12096 23808 12102
rect 23756 12038 23808 12044
rect 23768 11286 23796 12038
rect 23904 11996 24212 12005
rect 23904 11994 23910 11996
rect 23966 11994 23990 11996
rect 24046 11994 24070 11996
rect 24126 11994 24150 11996
rect 24206 11994 24212 11996
rect 23966 11942 23968 11994
rect 24148 11942 24150 11994
rect 23904 11940 23910 11942
rect 23966 11940 23990 11942
rect 24046 11940 24070 11942
rect 24126 11940 24150 11942
rect 24206 11940 24212 11942
rect 23904 11931 24212 11940
rect 24320 11642 24348 12854
rect 24596 11898 24624 13892
rect 24768 13874 24820 13880
rect 24872 13734 24900 14282
rect 25056 14074 25084 14418
rect 25136 14340 25188 14346
rect 25136 14282 25188 14288
rect 24952 14068 25004 14074
rect 24952 14010 25004 14016
rect 25044 14068 25096 14074
rect 25044 14010 25096 14016
rect 24860 13728 24912 13734
rect 24860 13670 24912 13676
rect 24872 13530 24900 13670
rect 24964 13530 24992 14010
rect 24860 13524 24912 13530
rect 24860 13466 24912 13472
rect 24952 13524 25004 13530
rect 24952 13466 25004 13472
rect 25148 13326 25176 14282
rect 25044 13320 25096 13326
rect 25044 13262 25096 13268
rect 25136 13320 25188 13326
rect 25136 13262 25188 13268
rect 24676 12980 24728 12986
rect 24676 12922 24728 12928
rect 24688 12646 24716 12922
rect 24952 12708 25004 12714
rect 24952 12650 25004 12656
rect 24676 12640 24728 12646
rect 24676 12582 24728 12588
rect 24768 12640 24820 12646
rect 24768 12582 24820 12588
rect 24780 12434 24808 12582
rect 24688 12406 24808 12434
rect 24584 11892 24636 11898
rect 24584 11834 24636 11840
rect 24320 11614 24532 11642
rect 24504 11558 24532 11614
rect 24688 11558 24716 12406
rect 24768 12232 24820 12238
rect 24768 12174 24820 12180
rect 24780 11898 24808 12174
rect 24860 12096 24912 12102
rect 24860 12038 24912 12044
rect 24768 11892 24820 11898
rect 24768 11834 24820 11840
rect 24872 11778 24900 12038
rect 24964 11898 24992 12650
rect 25056 12646 25084 13262
rect 25044 12640 25096 12646
rect 25044 12582 25096 12588
rect 24952 11892 25004 11898
rect 24952 11834 25004 11840
rect 24872 11762 24992 11778
rect 24872 11756 25004 11762
rect 24872 11750 24952 11756
rect 24952 11698 25004 11704
rect 24492 11552 24544 11558
rect 24492 11494 24544 11500
rect 24676 11552 24728 11558
rect 24676 11494 24728 11500
rect 24768 11552 24820 11558
rect 24768 11494 24820 11500
rect 23756 11280 23808 11286
rect 23756 11222 23808 11228
rect 23664 11144 23716 11150
rect 23664 11086 23716 11092
rect 23388 11076 23440 11082
rect 23388 11018 23440 11024
rect 23676 10130 23704 11086
rect 23904 10908 24212 10917
rect 23904 10906 23910 10908
rect 23966 10906 23990 10908
rect 24046 10906 24070 10908
rect 24126 10906 24150 10908
rect 24206 10906 24212 10908
rect 23966 10854 23968 10906
rect 24148 10854 24150 10906
rect 23904 10852 23910 10854
rect 23966 10852 23990 10854
rect 24046 10852 24070 10854
rect 24126 10852 24150 10854
rect 24206 10852 24212 10854
rect 23904 10843 24212 10852
rect 24504 10674 24532 11494
rect 24492 10668 24544 10674
rect 24492 10610 24544 10616
rect 24688 10606 24716 11494
rect 24676 10600 24728 10606
rect 24676 10542 24728 10548
rect 23664 10124 23716 10130
rect 23664 10066 23716 10072
rect 24676 10124 24728 10130
rect 24676 10066 24728 10072
rect 23904 9820 24212 9829
rect 23904 9818 23910 9820
rect 23966 9818 23990 9820
rect 24046 9818 24070 9820
rect 24126 9818 24150 9820
rect 24206 9818 24212 9820
rect 23966 9766 23968 9818
rect 24148 9766 24150 9818
rect 23904 9764 23910 9766
rect 23966 9764 23990 9766
rect 24046 9764 24070 9766
rect 24126 9764 24150 9766
rect 24206 9764 24212 9766
rect 23904 9755 24212 9764
rect 23480 9648 23532 9654
rect 23480 9590 23532 9596
rect 23020 9512 23072 9518
rect 23020 9454 23072 9460
rect 23032 9058 23060 9454
rect 23112 9376 23164 9382
rect 23112 9318 23164 9324
rect 23124 9178 23152 9318
rect 23492 9178 23520 9590
rect 24308 9580 24360 9586
rect 24308 9522 24360 9528
rect 23112 9172 23164 9178
rect 23112 9114 23164 9120
rect 23480 9172 23532 9178
rect 23480 9114 23532 9120
rect 23492 9058 23520 9114
rect 23032 9042 23152 9058
rect 23032 9036 23164 9042
rect 23032 9030 23112 9036
rect 23112 8978 23164 8984
rect 23400 9030 23520 9058
rect 23572 9036 23624 9042
rect 22836 8900 22888 8906
rect 22836 8842 22888 8848
rect 22848 8498 22876 8842
rect 22928 8832 22980 8838
rect 22928 8774 22980 8780
rect 23020 8832 23072 8838
rect 23020 8774 23072 8780
rect 22940 8634 22968 8774
rect 22928 8628 22980 8634
rect 22928 8570 22980 8576
rect 22836 8492 22888 8498
rect 22836 8434 22888 8440
rect 22848 7954 22876 8434
rect 23032 8378 23060 8774
rect 23124 8430 23152 8978
rect 23400 8498 23428 9030
rect 23572 8978 23624 8984
rect 23480 8900 23532 8906
rect 23480 8842 23532 8848
rect 23388 8492 23440 8498
rect 23388 8434 23440 8440
rect 23492 8430 23520 8842
rect 23584 8430 23612 8978
rect 23904 8732 24212 8741
rect 23904 8730 23910 8732
rect 23966 8730 23990 8732
rect 24046 8730 24070 8732
rect 24126 8730 24150 8732
rect 24206 8730 24212 8732
rect 23966 8678 23968 8730
rect 24148 8678 24150 8730
rect 23904 8676 23910 8678
rect 23966 8676 23990 8678
rect 24046 8676 24070 8678
rect 24126 8676 24150 8678
rect 24206 8676 24212 8678
rect 23904 8667 24212 8676
rect 24216 8628 24268 8634
rect 24320 8616 24348 9522
rect 24400 9376 24452 9382
rect 24400 9318 24452 9324
rect 24412 9178 24440 9318
rect 24688 9178 24716 10066
rect 24400 9172 24452 9178
rect 24400 9114 24452 9120
rect 24676 9172 24728 9178
rect 24676 9114 24728 9120
rect 24400 8968 24452 8974
rect 24400 8910 24452 8916
rect 24412 8634 24440 8910
rect 24268 8588 24348 8616
rect 24400 8628 24452 8634
rect 24216 8570 24268 8576
rect 24400 8570 24452 8576
rect 22940 8362 23060 8378
rect 23112 8424 23164 8430
rect 23112 8366 23164 8372
rect 23480 8424 23532 8430
rect 23480 8366 23532 8372
rect 23572 8424 23624 8430
rect 23572 8366 23624 8372
rect 23756 8424 23808 8430
rect 23756 8366 23808 8372
rect 24216 8424 24268 8430
rect 24216 8366 24268 8372
rect 22928 8356 23060 8362
rect 22980 8350 23060 8356
rect 22928 8298 22980 8304
rect 21968 7908 22048 7936
rect 22468 7948 22520 7954
rect 21916 7890 21968 7896
rect 22468 7890 22520 7896
rect 22744 7948 22796 7954
rect 22744 7890 22796 7896
rect 22836 7948 22888 7954
rect 22836 7890 22888 7896
rect 21640 7336 21692 7342
rect 21640 7278 21692 7284
rect 21652 6866 21680 7278
rect 21640 6860 21692 6866
rect 21640 6802 21692 6808
rect 21180 6792 21232 6798
rect 21180 6734 21232 6740
rect 21548 6792 21600 6798
rect 21548 6734 21600 6740
rect 21088 6724 21140 6730
rect 21088 6666 21140 6672
rect 20996 6452 21048 6458
rect 20996 6394 21048 6400
rect 20444 6112 20496 6118
rect 20444 6054 20496 6060
rect 20352 5160 20404 5166
rect 20352 5102 20404 5108
rect 20076 5024 20128 5030
rect 20076 4966 20128 4972
rect 20168 5024 20220 5030
rect 20168 4966 20220 4972
rect 20088 4758 20116 4966
rect 20076 4752 20128 4758
rect 20076 4694 20128 4700
rect 19984 4072 20036 4078
rect 19984 4014 20036 4020
rect 20180 3602 20208 4966
rect 20260 4072 20312 4078
rect 20260 4014 20312 4020
rect 20168 3596 20220 3602
rect 20168 3538 20220 3544
rect 19892 3120 19944 3126
rect 19892 3062 19944 3068
rect 18696 2916 18748 2922
rect 19352 2910 19564 2938
rect 19708 2984 19760 2990
rect 19708 2926 19760 2932
rect 20180 2922 20208 3538
rect 18696 2858 18748 2864
rect 19156 2848 19208 2854
rect 19156 2790 19208 2796
rect 18328 2576 18380 2582
rect 18328 2518 18380 2524
rect 18236 2508 18288 2514
rect 18236 2450 18288 2456
rect 18144 2440 18196 2446
rect 18144 2382 18196 2388
rect 17316 1896 17368 1902
rect 17316 1838 17368 1844
rect 17684 1896 17736 1902
rect 17684 1838 17736 1844
rect 17040 1488 17092 1494
rect 17040 1430 17092 1436
rect 17328 1426 17356 1838
rect 16764 1420 16816 1426
rect 16684 1380 16764 1408
rect 16396 808 16448 814
rect 16396 750 16448 756
rect 16684 400 16712 1380
rect 16764 1362 16816 1368
rect 17316 1420 17368 1426
rect 17316 1362 17368 1368
rect 17776 1420 17828 1426
rect 18512 1420 18564 1426
rect 17776 1362 17828 1368
rect 18340 1380 18512 1408
rect 17188 1116 17496 1125
rect 17188 1114 17194 1116
rect 17250 1114 17274 1116
rect 17330 1114 17354 1116
rect 17410 1114 17434 1116
rect 17490 1114 17496 1116
rect 17250 1062 17252 1114
rect 17432 1062 17434 1114
rect 17188 1060 17194 1062
rect 17250 1060 17274 1062
rect 17330 1060 17354 1062
rect 17410 1060 17434 1062
rect 17490 1060 17496 1062
rect 17188 1051 17496 1060
rect 17316 808 17368 814
rect 17236 768 17316 796
rect 17236 400 17264 768
rect 17316 750 17368 756
rect 17788 400 17816 1362
rect 17868 1216 17920 1222
rect 17868 1158 17920 1164
rect 17880 1018 17908 1158
rect 17868 1012 17920 1018
rect 17868 954 17920 960
rect 18340 400 18368 1380
rect 18512 1362 18564 1368
rect 18972 808 19024 814
rect 19168 796 19196 2790
rect 19340 1420 19392 1426
rect 19536 1408 19564 2910
rect 20168 2916 20220 2922
rect 20168 2858 20220 2864
rect 19708 2848 19760 2854
rect 19984 2848 20036 2854
rect 19708 2790 19760 2796
rect 19812 2808 19984 2836
rect 19720 2378 19748 2790
rect 19708 2372 19760 2378
rect 19708 2314 19760 2320
rect 19720 1562 19748 2314
rect 19812 1902 19840 2808
rect 19984 2790 20036 2796
rect 20272 2514 20300 4014
rect 20364 2990 20392 5102
rect 20456 4554 20484 6054
rect 20546 6012 20854 6021
rect 20546 6010 20552 6012
rect 20608 6010 20632 6012
rect 20688 6010 20712 6012
rect 20768 6010 20792 6012
rect 20848 6010 20854 6012
rect 20608 5958 20610 6010
rect 20790 5958 20792 6010
rect 20546 5956 20552 5958
rect 20608 5956 20632 5958
rect 20688 5956 20712 5958
rect 20768 5956 20792 5958
rect 20848 5956 20854 5958
rect 20546 5947 20854 5956
rect 20720 5568 20772 5574
rect 20720 5510 20772 5516
rect 20732 5370 20760 5510
rect 20720 5364 20772 5370
rect 20720 5306 20772 5312
rect 20720 5160 20772 5166
rect 20720 5102 20772 5108
rect 20732 5030 20760 5102
rect 21100 5098 21128 6666
rect 21456 6248 21508 6254
rect 21456 6190 21508 6196
rect 21468 5914 21496 6190
rect 21456 5908 21508 5914
rect 21456 5850 21508 5856
rect 21560 5574 21588 6734
rect 22480 6458 22508 7890
rect 22560 7744 22612 7750
rect 22560 7686 22612 7692
rect 22572 7274 22600 7686
rect 22560 7268 22612 7274
rect 22560 7210 22612 7216
rect 22756 7002 22784 7890
rect 22744 6996 22796 7002
rect 22744 6938 22796 6944
rect 23124 6730 23152 8366
rect 23492 8022 23520 8366
rect 23480 8016 23532 8022
rect 23480 7958 23532 7964
rect 23492 7546 23520 7958
rect 23584 7954 23612 8366
rect 23768 8090 23796 8366
rect 24228 8090 24256 8366
rect 23756 8084 23808 8090
rect 23756 8026 23808 8032
rect 24216 8084 24268 8090
rect 24216 8026 24268 8032
rect 23572 7948 23624 7954
rect 23572 7890 23624 7896
rect 23480 7540 23532 7546
rect 23480 7482 23532 7488
rect 23112 6724 23164 6730
rect 23112 6666 23164 6672
rect 23584 6458 23612 7890
rect 24308 7880 24360 7886
rect 24308 7822 24360 7828
rect 23904 7644 24212 7653
rect 23904 7642 23910 7644
rect 23966 7642 23990 7644
rect 24046 7642 24070 7644
rect 24126 7642 24150 7644
rect 24206 7642 24212 7644
rect 23966 7590 23968 7642
rect 24148 7590 24150 7642
rect 23904 7588 23910 7590
rect 23966 7588 23990 7590
rect 24046 7588 24070 7590
rect 24126 7588 24150 7590
rect 24206 7588 24212 7590
rect 23904 7579 24212 7588
rect 24320 7410 24348 7822
rect 24412 7478 24440 8570
rect 24780 8498 24808 11494
rect 24964 10810 24992 11698
rect 25056 11626 25084 12582
rect 25148 11694 25176 13262
rect 25240 12782 25268 14554
rect 25504 14544 25556 14550
rect 25504 14486 25556 14492
rect 25412 14476 25464 14482
rect 25412 14418 25464 14424
rect 25424 14362 25452 14418
rect 25332 14334 25452 14362
rect 25332 14278 25360 14334
rect 25320 14272 25372 14278
rect 25320 14214 25372 14220
rect 25332 12918 25360 14214
rect 25320 12912 25372 12918
rect 25320 12854 25372 12860
rect 25516 12850 25544 14486
rect 26148 14340 26200 14346
rect 26148 14282 26200 14288
rect 26160 13462 26188 14282
rect 26240 14272 26292 14278
rect 26240 14214 26292 14220
rect 26252 13870 26280 14214
rect 26896 13870 26924 14894
rect 27262 14716 27570 14725
rect 27262 14714 27268 14716
rect 27324 14714 27348 14716
rect 27404 14714 27428 14716
rect 27484 14714 27508 14716
rect 27564 14714 27570 14716
rect 27324 14662 27326 14714
rect 27506 14662 27508 14714
rect 27262 14660 27268 14662
rect 27324 14660 27348 14662
rect 27404 14660 27428 14662
rect 27484 14660 27508 14662
rect 27564 14660 27570 14662
rect 27262 14651 27570 14660
rect 26240 13864 26292 13870
rect 26240 13806 26292 13812
rect 26884 13864 26936 13870
rect 26884 13806 26936 13812
rect 26148 13456 26200 13462
rect 26148 13398 26200 13404
rect 26896 13394 26924 13806
rect 27262 13628 27570 13637
rect 27262 13626 27268 13628
rect 27324 13626 27348 13628
rect 27404 13626 27428 13628
rect 27484 13626 27508 13628
rect 27564 13626 27570 13628
rect 27324 13574 27326 13626
rect 27506 13574 27508 13626
rect 27262 13572 27268 13574
rect 27324 13572 27348 13574
rect 27404 13572 27428 13574
rect 27484 13572 27508 13574
rect 27564 13572 27570 13574
rect 27262 13563 27570 13572
rect 26884 13388 26936 13394
rect 26884 13330 26936 13336
rect 26240 12980 26292 12986
rect 26240 12922 26292 12928
rect 25504 12844 25556 12850
rect 25504 12786 25556 12792
rect 25228 12776 25280 12782
rect 25228 12718 25280 12724
rect 25320 12776 25372 12782
rect 25320 12718 25372 12724
rect 25332 12442 25360 12718
rect 25320 12436 25372 12442
rect 26252 12434 26280 12922
rect 26896 12850 26924 13330
rect 26884 12844 26936 12850
rect 26884 12786 26936 12792
rect 26608 12708 26660 12714
rect 26608 12650 26660 12656
rect 26620 12442 26648 12650
rect 26608 12436 26660 12442
rect 26252 12406 26464 12434
rect 25320 12378 25372 12384
rect 25136 11688 25188 11694
rect 25136 11630 25188 11636
rect 25044 11620 25096 11626
rect 25044 11562 25096 11568
rect 25332 11218 25360 12378
rect 25964 12368 26016 12374
rect 25964 12310 26016 12316
rect 25320 11212 25372 11218
rect 25320 11154 25372 11160
rect 24952 10804 25004 10810
rect 24952 10746 25004 10752
rect 24860 9920 24912 9926
rect 24860 9862 24912 9868
rect 24872 9518 24900 9862
rect 25976 9586 26004 12310
rect 26436 12306 26464 12406
rect 26608 12378 26660 12384
rect 26896 12374 26924 12786
rect 27262 12540 27570 12549
rect 27262 12538 27268 12540
rect 27324 12538 27348 12540
rect 27404 12538 27428 12540
rect 27484 12538 27508 12540
rect 27564 12538 27570 12540
rect 27324 12486 27326 12538
rect 27506 12486 27508 12538
rect 27262 12484 27268 12486
rect 27324 12484 27348 12486
rect 27404 12484 27428 12486
rect 27484 12484 27508 12486
rect 27564 12484 27570 12486
rect 27262 12475 27570 12484
rect 26884 12368 26936 12374
rect 26884 12310 26936 12316
rect 26424 12300 26476 12306
rect 26424 12242 26476 12248
rect 26896 11898 26924 12310
rect 26884 11892 26936 11898
rect 26884 11834 26936 11840
rect 27262 11452 27570 11461
rect 27262 11450 27268 11452
rect 27324 11450 27348 11452
rect 27404 11450 27428 11452
rect 27484 11450 27508 11452
rect 27564 11450 27570 11452
rect 27324 11398 27326 11450
rect 27506 11398 27508 11450
rect 27262 11396 27268 11398
rect 27324 11396 27348 11398
rect 27404 11396 27428 11398
rect 27484 11396 27508 11398
rect 27564 11396 27570 11398
rect 27262 11387 27570 11396
rect 27262 10364 27570 10373
rect 27262 10362 27268 10364
rect 27324 10362 27348 10364
rect 27404 10362 27428 10364
rect 27484 10362 27508 10364
rect 27564 10362 27570 10364
rect 27324 10310 27326 10362
rect 27506 10310 27508 10362
rect 27262 10308 27268 10310
rect 27324 10308 27348 10310
rect 27404 10308 27428 10310
rect 27484 10308 27508 10310
rect 27564 10308 27570 10310
rect 27262 10299 27570 10308
rect 25964 9580 26016 9586
rect 25964 9522 26016 9528
rect 24860 9512 24912 9518
rect 24860 9454 24912 9460
rect 25136 8560 25188 8566
rect 25136 8502 25188 8508
rect 24768 8492 24820 8498
rect 24768 8434 24820 8440
rect 24584 8356 24636 8362
rect 24584 8298 24636 8304
rect 24768 8356 24820 8362
rect 24768 8298 24820 8304
rect 24400 7472 24452 7478
rect 24400 7414 24452 7420
rect 24308 7404 24360 7410
rect 24308 7346 24360 7352
rect 23756 7336 23808 7342
rect 23756 7278 23808 7284
rect 22468 6452 22520 6458
rect 22468 6394 22520 6400
rect 23572 6452 23624 6458
rect 23572 6394 23624 6400
rect 23768 6322 23796 7278
rect 23904 6556 24212 6565
rect 23904 6554 23910 6556
rect 23966 6554 23990 6556
rect 24046 6554 24070 6556
rect 24126 6554 24150 6556
rect 24206 6554 24212 6556
rect 23966 6502 23968 6554
rect 24148 6502 24150 6554
rect 23904 6500 23910 6502
rect 23966 6500 23990 6502
rect 24046 6500 24070 6502
rect 24126 6500 24150 6502
rect 24206 6500 24212 6502
rect 23904 6491 24212 6500
rect 23756 6316 23808 6322
rect 23756 6258 23808 6264
rect 22560 6248 22612 6254
rect 22560 6190 22612 6196
rect 22836 6248 22888 6254
rect 22836 6190 22888 6196
rect 23480 6248 23532 6254
rect 23480 6190 23532 6196
rect 21732 6112 21784 6118
rect 21732 6054 21784 6060
rect 21548 5568 21600 5574
rect 21548 5510 21600 5516
rect 21560 5302 21588 5510
rect 21744 5370 21772 6054
rect 22572 5914 22600 6190
rect 22848 5914 22876 6190
rect 22560 5908 22612 5914
rect 22560 5850 22612 5856
rect 22836 5908 22888 5914
rect 22836 5850 22888 5856
rect 23020 5772 23072 5778
rect 23020 5714 23072 5720
rect 23204 5772 23256 5778
rect 23204 5714 23256 5720
rect 21732 5364 21784 5370
rect 21732 5306 21784 5312
rect 21548 5296 21600 5302
rect 21376 5244 21548 5250
rect 21376 5238 21600 5244
rect 21180 5228 21232 5234
rect 21180 5170 21232 5176
rect 21376 5222 21588 5238
rect 20904 5092 20956 5098
rect 20904 5034 20956 5040
rect 21088 5092 21140 5098
rect 21088 5034 21140 5040
rect 20720 5024 20772 5030
rect 20720 4966 20772 4972
rect 20546 4924 20854 4933
rect 20546 4922 20552 4924
rect 20608 4922 20632 4924
rect 20688 4922 20712 4924
rect 20768 4922 20792 4924
rect 20848 4922 20854 4924
rect 20608 4870 20610 4922
rect 20790 4870 20792 4922
rect 20546 4868 20552 4870
rect 20608 4868 20632 4870
rect 20688 4868 20712 4870
rect 20768 4868 20792 4870
rect 20848 4868 20854 4870
rect 20546 4859 20854 4868
rect 20444 4548 20496 4554
rect 20444 4490 20496 4496
rect 20916 4078 20944 5034
rect 21192 4758 21220 5170
rect 21180 4752 21232 4758
rect 21180 4694 21232 4700
rect 21192 4214 21220 4694
rect 21376 4486 21404 5222
rect 21456 5160 21508 5166
rect 21456 5102 21508 5108
rect 22744 5160 22796 5166
rect 22744 5102 22796 5108
rect 22928 5160 22980 5166
rect 22928 5102 22980 5108
rect 21468 4826 21496 5102
rect 22100 5024 22152 5030
rect 22100 4966 22152 4972
rect 22192 5024 22244 5030
rect 22192 4966 22244 4972
rect 22112 4826 22140 4966
rect 21456 4820 21508 4826
rect 21456 4762 21508 4768
rect 22100 4820 22152 4826
rect 22100 4762 22152 4768
rect 21364 4480 21416 4486
rect 21364 4422 21416 4428
rect 21376 4214 21404 4422
rect 21180 4208 21232 4214
rect 21180 4150 21232 4156
rect 21364 4208 21416 4214
rect 21364 4150 21416 4156
rect 21192 4078 21220 4150
rect 20904 4072 20956 4078
rect 20904 4014 20956 4020
rect 21180 4072 21232 4078
rect 21232 4032 21312 4060
rect 21180 4014 21232 4020
rect 21180 3936 21232 3942
rect 21180 3878 21232 3884
rect 20546 3836 20854 3845
rect 20546 3834 20552 3836
rect 20608 3834 20632 3836
rect 20688 3834 20712 3836
rect 20768 3834 20792 3836
rect 20848 3834 20854 3836
rect 20608 3782 20610 3834
rect 20790 3782 20792 3834
rect 20546 3780 20552 3782
rect 20608 3780 20632 3782
rect 20688 3780 20712 3782
rect 20768 3780 20792 3782
rect 20848 3780 20854 3782
rect 20546 3771 20854 3780
rect 21088 3528 21140 3534
rect 21088 3470 21140 3476
rect 21100 3126 21128 3470
rect 21088 3120 21140 3126
rect 21088 3062 21140 3068
rect 20996 3052 21048 3058
rect 20996 2994 21048 3000
rect 20352 2984 20404 2990
rect 20352 2926 20404 2932
rect 20720 2848 20772 2854
rect 20772 2808 20944 2836
rect 20720 2790 20772 2796
rect 20546 2748 20854 2757
rect 20546 2746 20552 2748
rect 20608 2746 20632 2748
rect 20688 2746 20712 2748
rect 20768 2746 20792 2748
rect 20848 2746 20854 2748
rect 20608 2694 20610 2746
rect 20790 2694 20792 2746
rect 20546 2692 20552 2694
rect 20608 2692 20632 2694
rect 20688 2692 20712 2694
rect 20768 2692 20792 2694
rect 20848 2692 20854 2694
rect 20546 2683 20854 2692
rect 20916 2582 20944 2808
rect 20904 2576 20956 2582
rect 20904 2518 20956 2524
rect 21008 2514 21036 2994
rect 21192 2514 21220 3878
rect 21284 3602 21312 4032
rect 21376 3618 21404 4150
rect 21468 3942 21496 4762
rect 21824 4072 21876 4078
rect 21744 4032 21824 4060
rect 21456 3936 21508 3942
rect 21456 3878 21508 3884
rect 21376 3602 21496 3618
rect 21272 3596 21324 3602
rect 21376 3596 21508 3602
rect 21376 3590 21456 3596
rect 21272 3538 21324 3544
rect 21456 3538 21508 3544
rect 21744 3534 21772 4032
rect 21824 4014 21876 4020
rect 22008 4004 22060 4010
rect 22008 3946 22060 3952
rect 21824 3936 21876 3942
rect 21824 3878 21876 3884
rect 21836 3738 21864 3878
rect 21824 3732 21876 3738
rect 21824 3674 21876 3680
rect 21916 3732 21968 3738
rect 21916 3674 21968 3680
rect 21732 3528 21784 3534
rect 21732 3470 21784 3476
rect 21456 3392 21508 3398
rect 21456 3334 21508 3340
rect 21468 3126 21496 3334
rect 21456 3120 21508 3126
rect 21456 3062 21508 3068
rect 21744 2922 21772 3470
rect 21824 3392 21876 3398
rect 21928 3380 21956 3674
rect 22020 3398 22048 3946
rect 22100 3596 22152 3602
rect 22100 3538 22152 3544
rect 21876 3352 21956 3380
rect 22008 3392 22060 3398
rect 21824 3334 21876 3340
rect 22008 3334 22060 3340
rect 21732 2916 21784 2922
rect 21732 2858 21784 2864
rect 21836 2514 21864 3334
rect 22112 3058 22140 3538
rect 22100 3052 22152 3058
rect 22100 2994 22152 3000
rect 20260 2508 20312 2514
rect 20260 2450 20312 2456
rect 20996 2508 21048 2514
rect 20996 2450 21048 2456
rect 21180 2508 21232 2514
rect 21180 2450 21232 2456
rect 21824 2508 21876 2514
rect 21824 2450 21876 2456
rect 20352 2372 20404 2378
rect 20352 2314 20404 2320
rect 19800 1896 19852 1902
rect 20076 1896 20128 1902
rect 19800 1838 19852 1844
rect 19996 1856 20076 1884
rect 19708 1556 19760 1562
rect 19708 1498 19760 1504
rect 19892 1488 19944 1494
rect 19892 1430 19944 1436
rect 19392 1380 19564 1408
rect 19340 1362 19392 1368
rect 19708 1352 19760 1358
rect 19708 1294 19760 1300
rect 19720 1018 19748 1294
rect 19708 1012 19760 1018
rect 19708 954 19760 960
rect 19024 768 19196 796
rect 19340 808 19392 814
rect 18972 750 19024 756
rect 19340 750 19392 756
rect 18892 462 19012 490
rect 18892 400 18920 462
rect 10704 326 10916 354
rect 11150 0 11206 400
rect 11702 0 11758 400
rect 12254 0 12310 400
rect 12806 0 12862 400
rect 13358 0 13414 400
rect 13910 0 13966 400
rect 14462 0 14518 400
rect 15014 0 15070 400
rect 15566 0 15622 400
rect 16118 0 16174 400
rect 16670 0 16726 400
rect 17222 0 17278 400
rect 17774 0 17830 400
rect 18326 0 18382 400
rect 18878 0 18934 400
rect 18984 354 19012 462
rect 19352 354 19380 750
rect 19444 462 19564 490
rect 19444 400 19472 462
rect 18984 326 19380 354
rect 19430 0 19486 400
rect 19536 354 19564 462
rect 19904 354 19932 1430
rect 19996 400 20024 1856
rect 20076 1838 20128 1844
rect 20364 814 20392 2314
rect 20444 2304 20496 2310
rect 20444 2246 20496 2252
rect 20996 2304 21048 2310
rect 20996 2246 21048 2252
rect 21548 2304 21600 2310
rect 21548 2246 21600 2252
rect 20456 1902 20484 2246
rect 20444 1896 20496 1902
rect 20444 1838 20496 1844
rect 20546 1660 20854 1669
rect 20546 1658 20552 1660
rect 20608 1658 20632 1660
rect 20688 1658 20712 1660
rect 20768 1658 20792 1660
rect 20848 1658 20854 1660
rect 20608 1606 20610 1658
rect 20790 1606 20792 1658
rect 20546 1604 20552 1606
rect 20608 1604 20632 1606
rect 20688 1604 20712 1606
rect 20768 1604 20792 1606
rect 20848 1604 20854 1606
rect 20546 1595 20854 1604
rect 21008 1562 21036 2246
rect 21272 1896 21324 1902
rect 21192 1856 21272 1884
rect 20996 1556 21048 1562
rect 20996 1498 21048 1504
rect 21088 1216 21140 1222
rect 21088 1158 21140 1164
rect 21100 1018 21128 1158
rect 21088 1012 21140 1018
rect 21088 954 21140 960
rect 21192 898 21220 1856
rect 21272 1838 21324 1844
rect 21456 1896 21508 1902
rect 21456 1838 21508 1844
rect 21468 1426 21496 1838
rect 21456 1420 21508 1426
rect 21456 1362 21508 1368
rect 21100 870 21220 898
rect 20260 808 20312 814
rect 20260 750 20312 756
rect 20352 808 20404 814
rect 20352 750 20404 756
rect 19536 326 19932 354
rect 19982 0 20038 400
rect 20272 354 20300 750
rect 20546 572 20854 581
rect 20546 570 20552 572
rect 20608 570 20632 572
rect 20688 570 20712 572
rect 20768 570 20792 572
rect 20848 570 20854 572
rect 20608 518 20610 570
rect 20790 518 20792 570
rect 20546 516 20552 518
rect 20608 516 20632 518
rect 20688 516 20712 518
rect 20768 516 20792 518
rect 20848 516 20854 518
rect 20546 507 20854 516
rect 20456 428 20576 456
rect 20456 354 20484 428
rect 20548 400 20576 428
rect 21100 400 21128 870
rect 21560 814 21588 2246
rect 21916 1896 21968 1902
rect 21916 1838 21968 1844
rect 21928 1018 21956 1838
rect 22112 1494 22140 2994
rect 22204 2990 22232 4966
rect 22560 4616 22612 4622
rect 22560 4558 22612 4564
rect 22284 4480 22336 4486
rect 22284 4422 22336 4428
rect 22468 4480 22520 4486
rect 22468 4422 22520 4428
rect 22296 4214 22324 4422
rect 22284 4208 22336 4214
rect 22284 4150 22336 4156
rect 22480 3602 22508 4422
rect 22572 4282 22600 4558
rect 22560 4276 22612 4282
rect 22560 4218 22612 4224
rect 22572 4078 22600 4218
rect 22652 4208 22704 4214
rect 22652 4150 22704 4156
rect 22664 4078 22692 4150
rect 22560 4072 22612 4078
rect 22560 4014 22612 4020
rect 22652 4072 22704 4078
rect 22652 4014 22704 4020
rect 22560 3936 22612 3942
rect 22560 3878 22612 3884
rect 22572 3738 22600 3878
rect 22560 3732 22612 3738
rect 22560 3674 22612 3680
rect 22468 3596 22520 3602
rect 22468 3538 22520 3544
rect 22560 3120 22612 3126
rect 22560 3062 22612 3068
rect 22192 2984 22244 2990
rect 22192 2926 22244 2932
rect 22204 2514 22232 2926
rect 22572 2514 22600 3062
rect 22192 2508 22244 2514
rect 22192 2450 22244 2456
rect 22560 2508 22612 2514
rect 22560 2450 22612 2456
rect 22664 1902 22692 4014
rect 22756 3924 22784 5102
rect 22940 4282 22968 5102
rect 22928 4276 22980 4282
rect 22928 4218 22980 4224
rect 22756 3896 22876 3924
rect 22744 3596 22796 3602
rect 22744 3538 22796 3544
rect 22756 3126 22784 3538
rect 22744 3120 22796 3126
rect 22744 3062 22796 3068
rect 22848 2650 22876 3896
rect 22940 3738 22968 4218
rect 22928 3732 22980 3738
rect 22928 3674 22980 3680
rect 23032 3534 23060 5714
rect 23216 5370 23244 5714
rect 23492 5710 23520 6190
rect 23480 5704 23532 5710
rect 23480 5646 23532 5652
rect 23768 5370 23796 6258
rect 24320 5914 24348 7346
rect 24492 6656 24544 6662
rect 24492 6598 24544 6604
rect 24504 6254 24532 6598
rect 24492 6248 24544 6254
rect 24492 6190 24544 6196
rect 24308 5908 24360 5914
rect 24308 5850 24360 5856
rect 24308 5636 24360 5642
rect 24308 5578 24360 5584
rect 23904 5468 24212 5477
rect 23904 5466 23910 5468
rect 23966 5466 23990 5468
rect 24046 5466 24070 5468
rect 24126 5466 24150 5468
rect 24206 5466 24212 5468
rect 23966 5414 23968 5466
rect 24148 5414 24150 5466
rect 23904 5412 23910 5414
rect 23966 5412 23990 5414
rect 24046 5412 24070 5414
rect 24126 5412 24150 5414
rect 24206 5412 24212 5414
rect 23904 5403 24212 5412
rect 23204 5364 23256 5370
rect 23204 5306 23256 5312
rect 23756 5364 23808 5370
rect 23756 5306 23808 5312
rect 23756 5160 23808 5166
rect 23756 5102 23808 5108
rect 23388 4684 23440 4690
rect 23388 4626 23440 4632
rect 23112 4480 23164 4486
rect 23112 4422 23164 4428
rect 23020 3528 23072 3534
rect 23020 3470 23072 3476
rect 23124 3398 23152 4422
rect 23204 4276 23256 4282
rect 23204 4218 23256 4224
rect 23112 3392 23164 3398
rect 23112 3334 23164 3340
rect 23124 2650 23152 3334
rect 23216 2854 23244 4218
rect 23400 4128 23428 4626
rect 23768 4146 23796 5102
rect 24320 4486 24348 5578
rect 24492 5364 24544 5370
rect 24492 5306 24544 5312
rect 24308 4480 24360 4486
rect 24308 4422 24360 4428
rect 23904 4380 24212 4389
rect 23904 4378 23910 4380
rect 23966 4378 23990 4380
rect 24046 4378 24070 4380
rect 24126 4378 24150 4380
rect 24206 4378 24212 4380
rect 23966 4326 23968 4378
rect 24148 4326 24150 4378
rect 23904 4324 23910 4326
rect 23966 4324 23990 4326
rect 24046 4324 24070 4326
rect 24126 4324 24150 4326
rect 24206 4324 24212 4326
rect 23904 4315 24212 4324
rect 23756 4140 23808 4146
rect 23400 4100 23612 4128
rect 23296 4072 23348 4078
rect 23296 4014 23348 4020
rect 23308 3738 23336 4014
rect 23480 3936 23532 3942
rect 23480 3878 23532 3884
rect 23492 3738 23520 3878
rect 23296 3732 23348 3738
rect 23296 3674 23348 3680
rect 23480 3732 23532 3738
rect 23480 3674 23532 3680
rect 23388 2984 23440 2990
rect 23388 2926 23440 2932
rect 23204 2848 23256 2854
rect 23204 2790 23256 2796
rect 23400 2774 23428 2926
rect 23584 2922 23612 4100
rect 23756 4082 23808 4088
rect 24216 4072 24268 4078
rect 24216 4014 24268 4020
rect 24228 3738 24256 4014
rect 24216 3732 24268 3738
rect 24216 3674 24268 3680
rect 24308 3460 24360 3466
rect 24308 3402 24360 3408
rect 23756 3392 23808 3398
rect 23756 3334 23808 3340
rect 23768 3194 23796 3334
rect 23904 3292 24212 3301
rect 23904 3290 23910 3292
rect 23966 3290 23990 3292
rect 24046 3290 24070 3292
rect 24126 3290 24150 3292
rect 24206 3290 24212 3292
rect 23966 3238 23968 3290
rect 24148 3238 24150 3290
rect 23904 3236 23910 3238
rect 23966 3236 23990 3238
rect 24046 3236 24070 3238
rect 24126 3236 24150 3238
rect 24206 3236 24212 3238
rect 23904 3227 24212 3236
rect 23756 3188 23808 3194
rect 23756 3130 23808 3136
rect 24320 2990 24348 3402
rect 24308 2984 24360 2990
rect 24308 2926 24360 2932
rect 23572 2916 23624 2922
rect 23572 2858 23624 2864
rect 23308 2746 23428 2774
rect 22836 2644 22888 2650
rect 22836 2586 22888 2592
rect 23112 2644 23164 2650
rect 23112 2586 23164 2592
rect 22560 1896 22612 1902
rect 22560 1838 22612 1844
rect 22652 1896 22704 1902
rect 22652 1838 22704 1844
rect 22100 1488 22152 1494
rect 22100 1430 22152 1436
rect 22008 1420 22060 1426
rect 22008 1362 22060 1368
rect 21916 1012 21968 1018
rect 21916 954 21968 960
rect 21548 808 21600 814
rect 21548 750 21600 756
rect 21652 462 21772 490
rect 21652 400 21680 462
rect 20272 326 20484 354
rect 20534 0 20590 400
rect 21086 0 21142 400
rect 21638 0 21694 400
rect 21744 354 21772 462
rect 22020 354 22048 1362
rect 22468 1352 22520 1358
rect 22468 1294 22520 1300
rect 22480 1018 22508 1294
rect 22572 1018 22600 1838
rect 22848 1562 22876 2586
rect 23308 2446 23336 2746
rect 23296 2440 23348 2446
rect 23296 2382 23348 2388
rect 23296 1896 23348 1902
rect 23296 1838 23348 1844
rect 22836 1556 22888 1562
rect 22836 1498 22888 1504
rect 22836 1420 22888 1426
rect 22836 1362 22888 1368
rect 22468 1012 22520 1018
rect 22468 954 22520 960
rect 22560 1012 22612 1018
rect 22560 954 22612 960
rect 22376 808 22428 814
rect 22204 768 22376 796
rect 22204 400 22232 768
rect 22848 762 22876 1362
rect 22376 750 22428 756
rect 22756 734 22876 762
rect 22756 400 22784 734
rect 23308 400 23336 1838
rect 23584 814 23612 2858
rect 24504 2514 24532 5306
rect 24596 5166 24624 8298
rect 24780 8022 24808 8298
rect 24768 8016 24820 8022
rect 24768 7958 24820 7964
rect 24780 7750 24808 7958
rect 25148 7954 25176 8502
rect 25596 8424 25648 8430
rect 25596 8366 25648 8372
rect 25228 8288 25280 8294
rect 25228 8230 25280 8236
rect 25136 7948 25188 7954
rect 25136 7890 25188 7896
rect 25044 7880 25096 7886
rect 25044 7822 25096 7828
rect 24768 7744 24820 7750
rect 24768 7686 24820 7692
rect 25056 7342 25084 7822
rect 25240 7410 25268 8230
rect 25504 7948 25556 7954
rect 25504 7890 25556 7896
rect 25320 7744 25372 7750
rect 25320 7686 25372 7692
rect 25332 7410 25360 7686
rect 25228 7404 25280 7410
rect 25228 7346 25280 7352
rect 25320 7404 25372 7410
rect 25320 7346 25372 7352
rect 25044 7336 25096 7342
rect 25044 7278 25096 7284
rect 25412 7336 25464 7342
rect 25412 7278 25464 7284
rect 25044 6860 25096 6866
rect 25044 6802 25096 6808
rect 24952 6792 25004 6798
rect 24952 6734 25004 6740
rect 24964 6458 24992 6734
rect 24952 6452 25004 6458
rect 24952 6394 25004 6400
rect 24584 5160 24636 5166
rect 24584 5102 24636 5108
rect 25056 4826 25084 6802
rect 25424 5914 25452 7278
rect 25516 7206 25544 7890
rect 25608 7546 25636 8366
rect 25976 8090 26004 9522
rect 27262 9276 27570 9285
rect 27262 9274 27268 9276
rect 27324 9274 27348 9276
rect 27404 9274 27428 9276
rect 27484 9274 27508 9276
rect 27564 9274 27570 9276
rect 27324 9222 27326 9274
rect 27506 9222 27508 9274
rect 27262 9220 27268 9222
rect 27324 9220 27348 9222
rect 27404 9220 27428 9222
rect 27484 9220 27508 9222
rect 27564 9220 27570 9222
rect 27262 9211 27570 9220
rect 26240 8356 26292 8362
rect 26240 8298 26292 8304
rect 26252 8090 26280 8298
rect 27262 8188 27570 8197
rect 27262 8186 27268 8188
rect 27324 8186 27348 8188
rect 27404 8186 27428 8188
rect 27484 8186 27508 8188
rect 27564 8186 27570 8188
rect 27324 8134 27326 8186
rect 27506 8134 27508 8186
rect 27262 8132 27268 8134
rect 27324 8132 27348 8134
rect 27404 8132 27428 8134
rect 27484 8132 27508 8134
rect 27564 8132 27570 8134
rect 27262 8123 27570 8132
rect 25964 8084 26016 8090
rect 25964 8026 26016 8032
rect 26240 8084 26292 8090
rect 26240 8026 26292 8032
rect 25596 7540 25648 7546
rect 25596 7482 25648 7488
rect 25504 7200 25556 7206
rect 25504 7142 25556 7148
rect 27262 7100 27570 7109
rect 27262 7098 27268 7100
rect 27324 7098 27348 7100
rect 27404 7098 27428 7100
rect 27484 7098 27508 7100
rect 27564 7098 27570 7100
rect 27324 7046 27326 7098
rect 27506 7046 27508 7098
rect 27262 7044 27268 7046
rect 27324 7044 27348 7046
rect 27404 7044 27428 7046
rect 27484 7044 27508 7046
rect 27564 7044 27570 7046
rect 27262 7035 27570 7044
rect 25596 6656 25648 6662
rect 25596 6598 25648 6604
rect 25688 6656 25740 6662
rect 25688 6598 25740 6604
rect 25780 6656 25832 6662
rect 25780 6598 25832 6604
rect 25608 6458 25636 6598
rect 25596 6452 25648 6458
rect 25596 6394 25648 6400
rect 25700 6186 25728 6598
rect 25792 6390 25820 6598
rect 25780 6384 25832 6390
rect 25780 6326 25832 6332
rect 25688 6180 25740 6186
rect 25688 6122 25740 6128
rect 25412 5908 25464 5914
rect 25412 5850 25464 5856
rect 25700 5710 25728 6122
rect 25792 5778 25820 6326
rect 26148 6248 26200 6254
rect 26148 6190 26200 6196
rect 25780 5772 25832 5778
rect 25780 5714 25832 5720
rect 26160 5710 26188 6190
rect 27262 6012 27570 6021
rect 27262 6010 27268 6012
rect 27324 6010 27348 6012
rect 27404 6010 27428 6012
rect 27484 6010 27508 6012
rect 27564 6010 27570 6012
rect 27324 5958 27326 6010
rect 27506 5958 27508 6010
rect 27262 5956 27268 5958
rect 27324 5956 27348 5958
rect 27404 5956 27428 5958
rect 27484 5956 27508 5958
rect 27564 5956 27570 5958
rect 27262 5947 27570 5956
rect 25688 5704 25740 5710
rect 25688 5646 25740 5652
rect 26148 5704 26200 5710
rect 26148 5646 26200 5652
rect 25780 5296 25832 5302
rect 25780 5238 25832 5244
rect 25596 5160 25648 5166
rect 25596 5102 25648 5108
rect 25044 4820 25096 4826
rect 25044 4762 25096 4768
rect 25608 4690 25636 5102
rect 25792 4826 25820 5238
rect 26056 5160 26108 5166
rect 26056 5102 26108 5108
rect 25780 4820 25832 4826
rect 25780 4762 25832 4768
rect 25792 4690 25820 4762
rect 26068 4690 26096 5102
rect 26160 4826 26188 5646
rect 26332 5364 26384 5370
rect 26332 5306 26384 5312
rect 26148 4820 26200 4826
rect 26148 4762 26200 4768
rect 25596 4684 25648 4690
rect 25596 4626 25648 4632
rect 25780 4684 25832 4690
rect 25780 4626 25832 4632
rect 26056 4684 26108 4690
rect 26056 4626 26108 4632
rect 25504 4548 25556 4554
rect 25504 4490 25556 4496
rect 25516 4282 25544 4490
rect 25504 4276 25556 4282
rect 25504 4218 25556 4224
rect 24952 3936 25004 3942
rect 24952 3878 25004 3884
rect 24964 3738 24992 3878
rect 24952 3732 25004 3738
rect 24952 3674 25004 3680
rect 24584 3392 24636 3398
rect 24584 3334 24636 3340
rect 24596 3194 24624 3334
rect 25608 3194 25636 4626
rect 25688 3936 25740 3942
rect 25688 3878 25740 3884
rect 25700 3738 25728 3878
rect 25688 3732 25740 3738
rect 25688 3674 25740 3680
rect 25792 3534 25820 4626
rect 26344 4282 26372 5306
rect 26792 5024 26844 5030
rect 26792 4966 26844 4972
rect 26424 4752 26476 4758
rect 26424 4694 26476 4700
rect 26332 4276 26384 4282
rect 26332 4218 26384 4224
rect 25780 3528 25832 3534
rect 25780 3470 25832 3476
rect 26436 3466 26464 4694
rect 26804 4622 26832 4966
rect 27262 4924 27570 4933
rect 27262 4922 27268 4924
rect 27324 4922 27348 4924
rect 27404 4922 27428 4924
rect 27484 4922 27508 4924
rect 27564 4922 27570 4924
rect 27324 4870 27326 4922
rect 27506 4870 27508 4922
rect 27262 4868 27268 4870
rect 27324 4868 27348 4870
rect 27404 4868 27428 4870
rect 27484 4868 27508 4870
rect 27564 4868 27570 4870
rect 27262 4859 27570 4868
rect 26792 4616 26844 4622
rect 26792 4558 26844 4564
rect 26884 4480 26936 4486
rect 26884 4422 26936 4428
rect 26896 4010 26924 4422
rect 26884 4004 26936 4010
rect 26884 3946 26936 3952
rect 27262 3836 27570 3845
rect 27262 3834 27268 3836
rect 27324 3834 27348 3836
rect 27404 3834 27428 3836
rect 27484 3834 27508 3836
rect 27564 3834 27570 3836
rect 27324 3782 27326 3834
rect 27506 3782 27508 3834
rect 27262 3780 27268 3782
rect 27324 3780 27348 3782
rect 27404 3780 27428 3782
rect 27484 3780 27508 3782
rect 27564 3780 27570 3782
rect 27262 3771 27570 3780
rect 25688 3460 25740 3466
rect 25688 3402 25740 3408
rect 26424 3460 26476 3466
rect 26424 3402 26476 3408
rect 24584 3188 24636 3194
rect 24584 3130 24636 3136
rect 25596 3188 25648 3194
rect 25596 3130 25648 3136
rect 25136 2984 25188 2990
rect 25136 2926 25188 2932
rect 24860 2848 24912 2854
rect 24860 2790 24912 2796
rect 25044 2848 25096 2854
rect 25044 2790 25096 2796
rect 24400 2508 24452 2514
rect 24400 2450 24452 2456
rect 24492 2508 24544 2514
rect 24492 2450 24544 2456
rect 23904 2204 24212 2213
rect 23904 2202 23910 2204
rect 23966 2202 23990 2204
rect 24046 2202 24070 2204
rect 24126 2202 24150 2204
rect 24206 2202 24212 2204
rect 23966 2150 23968 2202
rect 24148 2150 24150 2202
rect 23904 2148 23910 2150
rect 23966 2148 23990 2150
rect 24046 2148 24070 2150
rect 24126 2148 24150 2150
rect 24206 2148 24212 2150
rect 23904 2139 24212 2148
rect 23756 1896 23808 1902
rect 23756 1838 23808 1844
rect 23664 1352 23716 1358
rect 23664 1294 23716 1300
rect 23676 1018 23704 1294
rect 23664 1012 23716 1018
rect 23664 954 23716 960
rect 23768 882 23796 1838
rect 24308 1420 24360 1426
rect 24308 1362 24360 1368
rect 23904 1116 24212 1125
rect 23904 1114 23910 1116
rect 23966 1114 23990 1116
rect 24046 1114 24070 1116
rect 24126 1114 24150 1116
rect 24206 1114 24212 1116
rect 23966 1062 23968 1114
rect 24148 1062 24150 1114
rect 23904 1060 23910 1062
rect 23966 1060 23990 1062
rect 24046 1060 24070 1062
rect 24126 1060 24150 1062
rect 24206 1060 24212 1062
rect 23904 1051 24212 1060
rect 23756 876 23808 882
rect 23756 818 23808 824
rect 23572 808 23624 814
rect 23572 750 23624 756
rect 23860 462 23980 490
rect 23860 400 23888 462
rect 21744 326 22048 354
rect 22190 0 22246 400
rect 22742 0 22798 400
rect 23294 0 23350 400
rect 23846 0 23902 400
rect 23952 354 23980 462
rect 24320 354 24348 1362
rect 24412 400 24440 2450
rect 24872 1902 24900 2790
rect 25056 2582 25084 2790
rect 25044 2576 25096 2582
rect 25044 2518 25096 2524
rect 24860 1896 24912 1902
rect 24860 1838 24912 1844
rect 25148 1426 25176 2926
rect 25700 2922 25728 3402
rect 25688 2916 25740 2922
rect 25688 2858 25740 2864
rect 26056 2916 26108 2922
rect 26056 2858 26108 2864
rect 26068 2650 26096 2858
rect 27262 2748 27570 2757
rect 27262 2746 27268 2748
rect 27324 2746 27348 2748
rect 27404 2746 27428 2748
rect 27484 2746 27508 2748
rect 27564 2746 27570 2748
rect 27324 2694 27326 2746
rect 27506 2694 27508 2746
rect 27262 2692 27268 2694
rect 27324 2692 27348 2694
rect 27404 2692 27428 2694
rect 27484 2692 27508 2694
rect 27564 2692 27570 2694
rect 27262 2683 27570 2692
rect 26056 2644 26108 2650
rect 26056 2586 26108 2592
rect 26056 1896 26108 1902
rect 26056 1838 26108 1844
rect 25320 1828 25372 1834
rect 25320 1770 25372 1776
rect 25136 1420 25188 1426
rect 25136 1362 25188 1368
rect 24860 1352 24912 1358
rect 24860 1294 24912 1300
rect 24872 1018 24900 1294
rect 25332 1018 25360 1770
rect 25504 1420 25556 1426
rect 25504 1362 25556 1368
rect 24860 1012 24912 1018
rect 24860 954 24912 960
rect 25320 1012 25372 1018
rect 25320 954 25372 960
rect 24952 808 25004 814
rect 24952 750 25004 756
rect 24964 400 24992 750
rect 25516 400 25544 1362
rect 26068 400 26096 1838
rect 27262 1660 27570 1669
rect 27262 1658 27268 1660
rect 27324 1658 27348 1660
rect 27404 1658 27428 1660
rect 27484 1658 27508 1660
rect 27564 1658 27570 1660
rect 27324 1606 27326 1658
rect 27506 1606 27508 1658
rect 27262 1604 27268 1606
rect 27324 1604 27348 1606
rect 27404 1604 27428 1606
rect 27484 1604 27508 1606
rect 27564 1604 27570 1606
rect 27262 1595 27570 1604
rect 27262 572 27570 581
rect 27262 570 27268 572
rect 27324 570 27348 572
rect 27404 570 27428 572
rect 27484 570 27508 572
rect 27564 570 27570 572
rect 27324 518 27326 570
rect 27506 518 27508 570
rect 27262 516 27268 518
rect 27324 516 27348 518
rect 27404 516 27428 518
rect 27484 516 27508 518
rect 27564 516 27570 518
rect 27262 507 27570 516
rect 23952 326 24348 354
rect 24398 0 24454 400
rect 24950 0 25006 400
rect 25502 0 25558 400
rect 26054 0 26110 400
<< via2 >>
rect 2042 30368 2098 30424
rect 3762 30490 3818 30492
rect 3842 30490 3898 30492
rect 3922 30490 3978 30492
rect 4002 30490 4058 30492
rect 3762 30438 3808 30490
rect 3808 30438 3818 30490
rect 3842 30438 3872 30490
rect 3872 30438 3884 30490
rect 3884 30438 3898 30490
rect 3922 30438 3936 30490
rect 3936 30438 3948 30490
rect 3948 30438 3978 30490
rect 4002 30438 4012 30490
rect 4012 30438 4058 30490
rect 3762 30436 3818 30438
rect 3842 30436 3898 30438
rect 3922 30436 3978 30438
rect 4002 30436 4058 30438
rect 1858 29688 1914 29744
rect 3762 29402 3818 29404
rect 3842 29402 3898 29404
rect 3922 29402 3978 29404
rect 4002 29402 4058 29404
rect 3762 29350 3808 29402
rect 3808 29350 3818 29402
rect 3842 29350 3872 29402
rect 3872 29350 3884 29402
rect 3884 29350 3898 29402
rect 3922 29350 3936 29402
rect 3936 29350 3948 29402
rect 3948 29350 3978 29402
rect 4002 29350 4012 29402
rect 4012 29350 4058 29402
rect 3762 29348 3818 29350
rect 3842 29348 3898 29350
rect 3922 29348 3978 29350
rect 4002 29348 4058 29350
rect 7120 31034 7176 31036
rect 7200 31034 7256 31036
rect 7280 31034 7336 31036
rect 7360 31034 7416 31036
rect 7120 30982 7166 31034
rect 7166 30982 7176 31034
rect 7200 30982 7230 31034
rect 7230 30982 7242 31034
rect 7242 30982 7256 31034
rect 7280 30982 7294 31034
rect 7294 30982 7306 31034
rect 7306 30982 7336 31034
rect 7360 30982 7370 31034
rect 7370 30982 7416 31034
rect 7120 30980 7176 30982
rect 7200 30980 7256 30982
rect 7280 30980 7336 30982
rect 7360 30980 7416 30982
rect 4158 29008 4214 29064
rect 3762 28314 3818 28316
rect 3842 28314 3898 28316
rect 3922 28314 3978 28316
rect 4002 28314 4058 28316
rect 3762 28262 3808 28314
rect 3808 28262 3818 28314
rect 3842 28262 3872 28314
rect 3872 28262 3884 28314
rect 3884 28262 3898 28314
rect 3922 28262 3936 28314
rect 3936 28262 3948 28314
rect 3948 28262 3978 28314
rect 4002 28262 4012 28314
rect 4012 28262 4058 28314
rect 3762 28260 3818 28262
rect 3842 28260 3898 28262
rect 3922 28260 3978 28262
rect 4002 28260 4058 28262
rect 4618 29044 4620 29064
rect 4620 29044 4672 29064
rect 4672 29044 4674 29064
rect 4618 29008 4674 29044
rect 3762 27226 3818 27228
rect 3842 27226 3898 27228
rect 3922 27226 3978 27228
rect 4002 27226 4058 27228
rect 3762 27174 3808 27226
rect 3808 27174 3818 27226
rect 3842 27174 3872 27226
rect 3872 27174 3884 27226
rect 3884 27174 3898 27226
rect 3922 27174 3936 27226
rect 3936 27174 3948 27226
rect 3948 27174 3978 27226
rect 4002 27174 4012 27226
rect 4012 27174 4058 27226
rect 3762 27172 3818 27174
rect 3842 27172 3898 27174
rect 3922 27172 3978 27174
rect 4002 27172 4058 27174
rect 3762 26138 3818 26140
rect 3842 26138 3898 26140
rect 3922 26138 3978 26140
rect 4002 26138 4058 26140
rect 3762 26086 3808 26138
rect 3808 26086 3818 26138
rect 3842 26086 3872 26138
rect 3872 26086 3884 26138
rect 3884 26086 3898 26138
rect 3922 26086 3936 26138
rect 3936 26086 3948 26138
rect 3948 26086 3978 26138
rect 4002 26086 4012 26138
rect 4012 26086 4058 26138
rect 3762 26084 3818 26086
rect 3842 26084 3898 26086
rect 3922 26084 3978 26086
rect 4002 26084 4058 26086
rect 3762 25050 3818 25052
rect 3842 25050 3898 25052
rect 3922 25050 3978 25052
rect 4002 25050 4058 25052
rect 3762 24998 3808 25050
rect 3808 24998 3818 25050
rect 3842 24998 3872 25050
rect 3872 24998 3884 25050
rect 3884 24998 3898 25050
rect 3922 24998 3936 25050
rect 3936 24998 3948 25050
rect 3948 24998 3978 25050
rect 4002 24998 4012 25050
rect 4012 24998 4058 25050
rect 3762 24996 3818 24998
rect 3842 24996 3898 24998
rect 3922 24996 3978 24998
rect 4002 24996 4058 24998
rect 3762 23962 3818 23964
rect 3842 23962 3898 23964
rect 3922 23962 3978 23964
rect 4002 23962 4058 23964
rect 3762 23910 3808 23962
rect 3808 23910 3818 23962
rect 3842 23910 3872 23962
rect 3872 23910 3884 23962
rect 3884 23910 3898 23962
rect 3922 23910 3936 23962
rect 3936 23910 3948 23962
rect 3948 23910 3978 23962
rect 4002 23910 4012 23962
rect 4012 23910 4058 23962
rect 3762 23908 3818 23910
rect 3842 23908 3898 23910
rect 3922 23908 3978 23910
rect 4002 23908 4058 23910
rect 3762 22874 3818 22876
rect 3842 22874 3898 22876
rect 3922 22874 3978 22876
rect 4002 22874 4058 22876
rect 3762 22822 3808 22874
rect 3808 22822 3818 22874
rect 3842 22822 3872 22874
rect 3872 22822 3884 22874
rect 3884 22822 3898 22874
rect 3922 22822 3936 22874
rect 3936 22822 3948 22874
rect 3948 22822 3978 22874
rect 4002 22822 4012 22874
rect 4012 22822 4058 22874
rect 3762 22820 3818 22822
rect 3842 22820 3898 22822
rect 3922 22820 3978 22822
rect 4002 22820 4058 22822
rect 3762 21786 3818 21788
rect 3842 21786 3898 21788
rect 3922 21786 3978 21788
rect 4002 21786 4058 21788
rect 3762 21734 3808 21786
rect 3808 21734 3818 21786
rect 3842 21734 3872 21786
rect 3872 21734 3884 21786
rect 3884 21734 3898 21786
rect 3922 21734 3936 21786
rect 3936 21734 3948 21786
rect 3948 21734 3978 21786
rect 4002 21734 4012 21786
rect 4012 21734 4058 21786
rect 3762 21732 3818 21734
rect 3842 21732 3898 21734
rect 3922 21732 3978 21734
rect 4002 21732 4058 21734
rect 3762 20698 3818 20700
rect 3842 20698 3898 20700
rect 3922 20698 3978 20700
rect 4002 20698 4058 20700
rect 3762 20646 3808 20698
rect 3808 20646 3818 20698
rect 3842 20646 3872 20698
rect 3872 20646 3884 20698
rect 3884 20646 3898 20698
rect 3922 20646 3936 20698
rect 3936 20646 3948 20698
rect 3948 20646 3978 20698
rect 4002 20646 4012 20698
rect 4012 20646 4058 20698
rect 3762 20644 3818 20646
rect 3842 20644 3898 20646
rect 3922 20644 3978 20646
rect 4002 20644 4058 20646
rect 3762 19610 3818 19612
rect 3842 19610 3898 19612
rect 3922 19610 3978 19612
rect 4002 19610 4058 19612
rect 3762 19558 3808 19610
rect 3808 19558 3818 19610
rect 3842 19558 3872 19610
rect 3872 19558 3884 19610
rect 3884 19558 3898 19610
rect 3922 19558 3936 19610
rect 3936 19558 3948 19610
rect 3948 19558 3978 19610
rect 4002 19558 4012 19610
rect 4012 19558 4058 19610
rect 3762 19556 3818 19558
rect 3842 19556 3898 19558
rect 3922 19556 3978 19558
rect 4002 19556 4058 19558
rect 3762 18522 3818 18524
rect 3842 18522 3898 18524
rect 3922 18522 3978 18524
rect 4002 18522 4058 18524
rect 3762 18470 3808 18522
rect 3808 18470 3818 18522
rect 3842 18470 3872 18522
rect 3872 18470 3884 18522
rect 3884 18470 3898 18522
rect 3922 18470 3936 18522
rect 3936 18470 3948 18522
rect 3948 18470 3978 18522
rect 4002 18470 4012 18522
rect 4012 18470 4058 18522
rect 3762 18468 3818 18470
rect 3842 18468 3898 18470
rect 3922 18468 3978 18470
rect 4002 18468 4058 18470
rect 3762 17434 3818 17436
rect 3842 17434 3898 17436
rect 3922 17434 3978 17436
rect 4002 17434 4058 17436
rect 3762 17382 3808 17434
rect 3808 17382 3818 17434
rect 3842 17382 3872 17434
rect 3872 17382 3884 17434
rect 3884 17382 3898 17434
rect 3922 17382 3936 17434
rect 3936 17382 3948 17434
rect 3948 17382 3978 17434
rect 4002 17382 4012 17434
rect 4012 17382 4058 17434
rect 3762 17380 3818 17382
rect 3842 17380 3898 17382
rect 3922 17380 3978 17382
rect 4002 17380 4058 17382
rect 3762 16346 3818 16348
rect 3842 16346 3898 16348
rect 3922 16346 3978 16348
rect 4002 16346 4058 16348
rect 3762 16294 3808 16346
rect 3808 16294 3818 16346
rect 3842 16294 3872 16346
rect 3872 16294 3884 16346
rect 3884 16294 3898 16346
rect 3922 16294 3936 16346
rect 3936 16294 3948 16346
rect 3948 16294 3978 16346
rect 4002 16294 4012 16346
rect 4012 16294 4058 16346
rect 3762 16292 3818 16294
rect 3842 16292 3898 16294
rect 3922 16292 3978 16294
rect 4002 16292 4058 16294
rect 6458 29416 6514 29472
rect 7120 29946 7176 29948
rect 7200 29946 7256 29948
rect 7280 29946 7336 29948
rect 7360 29946 7416 29948
rect 7120 29894 7166 29946
rect 7166 29894 7176 29946
rect 7200 29894 7230 29946
rect 7230 29894 7242 29946
rect 7242 29894 7256 29946
rect 7280 29894 7294 29946
rect 7294 29894 7306 29946
rect 7306 29894 7336 29946
rect 7360 29894 7370 29946
rect 7370 29894 7416 29946
rect 7120 29892 7176 29894
rect 7200 29892 7256 29894
rect 7280 29892 7336 29894
rect 7360 29892 7416 29894
rect 6366 24792 6422 24848
rect 6366 24656 6422 24712
rect 6366 24248 6422 24304
rect 7120 28858 7176 28860
rect 7200 28858 7256 28860
rect 7280 28858 7336 28860
rect 7360 28858 7416 28860
rect 7120 28806 7166 28858
rect 7166 28806 7176 28858
rect 7200 28806 7230 28858
rect 7230 28806 7242 28858
rect 7242 28806 7256 28858
rect 7280 28806 7294 28858
rect 7294 28806 7306 28858
rect 7306 28806 7336 28858
rect 7360 28806 7370 28858
rect 7370 28806 7416 28858
rect 7120 28804 7176 28806
rect 7200 28804 7256 28806
rect 7280 28804 7336 28806
rect 7360 28804 7416 28806
rect 7746 29416 7802 29472
rect 10478 30490 10534 30492
rect 10558 30490 10614 30492
rect 10638 30490 10694 30492
rect 10718 30490 10774 30492
rect 10478 30438 10524 30490
rect 10524 30438 10534 30490
rect 10558 30438 10588 30490
rect 10588 30438 10600 30490
rect 10600 30438 10614 30490
rect 10638 30438 10652 30490
rect 10652 30438 10664 30490
rect 10664 30438 10694 30490
rect 10718 30438 10728 30490
rect 10728 30438 10774 30490
rect 10478 30436 10534 30438
rect 10558 30436 10614 30438
rect 10638 30436 10694 30438
rect 10718 30436 10774 30438
rect 10478 29402 10534 29404
rect 10558 29402 10614 29404
rect 10638 29402 10694 29404
rect 10718 29402 10774 29404
rect 10478 29350 10524 29402
rect 10524 29350 10534 29402
rect 10558 29350 10588 29402
rect 10588 29350 10600 29402
rect 10600 29350 10614 29402
rect 10638 29350 10652 29402
rect 10652 29350 10664 29402
rect 10664 29350 10694 29402
rect 10718 29350 10728 29402
rect 10728 29350 10774 29402
rect 10478 29348 10534 29350
rect 10558 29348 10614 29350
rect 10638 29348 10694 29350
rect 10718 29348 10774 29350
rect 7120 27770 7176 27772
rect 7200 27770 7256 27772
rect 7280 27770 7336 27772
rect 7360 27770 7416 27772
rect 7120 27718 7166 27770
rect 7166 27718 7176 27770
rect 7200 27718 7230 27770
rect 7230 27718 7242 27770
rect 7242 27718 7256 27770
rect 7280 27718 7294 27770
rect 7294 27718 7306 27770
rect 7306 27718 7336 27770
rect 7360 27718 7370 27770
rect 7370 27718 7416 27770
rect 7120 27716 7176 27718
rect 7200 27716 7256 27718
rect 7280 27716 7336 27718
rect 7360 27716 7416 27718
rect 7120 26682 7176 26684
rect 7200 26682 7256 26684
rect 7280 26682 7336 26684
rect 7360 26682 7416 26684
rect 7120 26630 7166 26682
rect 7166 26630 7176 26682
rect 7200 26630 7230 26682
rect 7230 26630 7242 26682
rect 7242 26630 7256 26682
rect 7280 26630 7294 26682
rect 7294 26630 7306 26682
rect 7306 26630 7336 26682
rect 7360 26630 7370 26682
rect 7370 26630 7416 26682
rect 7120 26628 7176 26630
rect 7200 26628 7256 26630
rect 7280 26628 7336 26630
rect 7360 26628 7416 26630
rect 11978 29552 12034 29608
rect 7120 25594 7176 25596
rect 7200 25594 7256 25596
rect 7280 25594 7336 25596
rect 7360 25594 7416 25596
rect 7120 25542 7166 25594
rect 7166 25542 7176 25594
rect 7200 25542 7230 25594
rect 7230 25542 7242 25594
rect 7242 25542 7256 25594
rect 7280 25542 7294 25594
rect 7294 25542 7306 25594
rect 7306 25542 7336 25594
rect 7360 25542 7370 25594
rect 7370 25542 7416 25594
rect 7120 25540 7176 25542
rect 7200 25540 7256 25542
rect 7280 25540 7336 25542
rect 7360 25540 7416 25542
rect 7120 24506 7176 24508
rect 7200 24506 7256 24508
rect 7280 24506 7336 24508
rect 7360 24506 7416 24508
rect 7120 24454 7166 24506
rect 7166 24454 7176 24506
rect 7200 24454 7230 24506
rect 7230 24454 7242 24506
rect 7242 24454 7256 24506
rect 7280 24454 7294 24506
rect 7294 24454 7306 24506
rect 7306 24454 7336 24506
rect 7360 24454 7370 24506
rect 7370 24454 7416 24506
rect 7120 24452 7176 24454
rect 7200 24452 7256 24454
rect 7280 24452 7336 24454
rect 7360 24452 7416 24454
rect 6918 24012 6920 24032
rect 6920 24012 6972 24032
rect 6972 24012 6974 24032
rect 6918 23976 6974 24012
rect 7654 24676 7710 24712
rect 7654 24656 7656 24676
rect 7656 24656 7708 24676
rect 7708 24656 7710 24676
rect 7120 23418 7176 23420
rect 7200 23418 7256 23420
rect 7280 23418 7336 23420
rect 7360 23418 7416 23420
rect 7120 23366 7166 23418
rect 7166 23366 7176 23418
rect 7200 23366 7230 23418
rect 7230 23366 7242 23418
rect 7242 23366 7256 23418
rect 7280 23366 7294 23418
rect 7294 23366 7306 23418
rect 7306 23366 7336 23418
rect 7360 23366 7370 23418
rect 7370 23366 7416 23418
rect 7120 23364 7176 23366
rect 7200 23364 7256 23366
rect 7280 23364 7336 23366
rect 7360 23364 7416 23366
rect 7930 24268 7986 24304
rect 7930 24248 7932 24268
rect 7932 24248 7984 24268
rect 7984 24248 7986 24268
rect 7838 23976 7894 24032
rect 7120 22330 7176 22332
rect 7200 22330 7256 22332
rect 7280 22330 7336 22332
rect 7360 22330 7416 22332
rect 7120 22278 7166 22330
rect 7166 22278 7176 22330
rect 7200 22278 7230 22330
rect 7230 22278 7242 22330
rect 7242 22278 7256 22330
rect 7280 22278 7294 22330
rect 7294 22278 7306 22330
rect 7306 22278 7336 22330
rect 7360 22278 7370 22330
rect 7370 22278 7416 22330
rect 7120 22276 7176 22278
rect 7200 22276 7256 22278
rect 7280 22276 7336 22278
rect 7360 22276 7416 22278
rect 7120 21242 7176 21244
rect 7200 21242 7256 21244
rect 7280 21242 7336 21244
rect 7360 21242 7416 21244
rect 7120 21190 7166 21242
rect 7166 21190 7176 21242
rect 7200 21190 7230 21242
rect 7230 21190 7242 21242
rect 7242 21190 7256 21242
rect 7280 21190 7294 21242
rect 7294 21190 7306 21242
rect 7306 21190 7336 21242
rect 7360 21190 7370 21242
rect 7370 21190 7416 21242
rect 7120 21188 7176 21190
rect 7200 21188 7256 21190
rect 7280 21188 7336 21190
rect 7360 21188 7416 21190
rect 7120 20154 7176 20156
rect 7200 20154 7256 20156
rect 7280 20154 7336 20156
rect 7360 20154 7416 20156
rect 7120 20102 7166 20154
rect 7166 20102 7176 20154
rect 7200 20102 7230 20154
rect 7230 20102 7242 20154
rect 7242 20102 7256 20154
rect 7280 20102 7294 20154
rect 7294 20102 7306 20154
rect 7306 20102 7336 20154
rect 7360 20102 7370 20154
rect 7370 20102 7416 20154
rect 7120 20100 7176 20102
rect 7200 20100 7256 20102
rect 7280 20100 7336 20102
rect 7360 20100 7416 20102
rect 8114 24792 8170 24848
rect 7120 19066 7176 19068
rect 7200 19066 7256 19068
rect 7280 19066 7336 19068
rect 7360 19066 7416 19068
rect 7120 19014 7166 19066
rect 7166 19014 7176 19066
rect 7200 19014 7230 19066
rect 7230 19014 7242 19066
rect 7242 19014 7256 19066
rect 7280 19014 7294 19066
rect 7294 19014 7306 19066
rect 7306 19014 7336 19066
rect 7360 19014 7370 19066
rect 7370 19014 7416 19066
rect 7120 19012 7176 19014
rect 7200 19012 7256 19014
rect 7280 19012 7336 19014
rect 7360 19012 7416 19014
rect 7120 17978 7176 17980
rect 7200 17978 7256 17980
rect 7280 17978 7336 17980
rect 7360 17978 7416 17980
rect 7120 17926 7166 17978
rect 7166 17926 7176 17978
rect 7200 17926 7230 17978
rect 7230 17926 7242 17978
rect 7242 17926 7256 17978
rect 7280 17926 7294 17978
rect 7294 17926 7306 17978
rect 7306 17926 7336 17978
rect 7360 17926 7370 17978
rect 7370 17926 7416 17978
rect 7120 17924 7176 17926
rect 7200 17924 7256 17926
rect 7280 17924 7336 17926
rect 7360 17924 7416 17926
rect 7120 16890 7176 16892
rect 7200 16890 7256 16892
rect 7280 16890 7336 16892
rect 7360 16890 7416 16892
rect 7120 16838 7166 16890
rect 7166 16838 7176 16890
rect 7200 16838 7230 16890
rect 7230 16838 7242 16890
rect 7242 16838 7256 16890
rect 7280 16838 7294 16890
rect 7294 16838 7306 16890
rect 7306 16838 7336 16890
rect 7360 16838 7370 16890
rect 7370 16838 7416 16890
rect 7120 16836 7176 16838
rect 7200 16836 7256 16838
rect 7280 16836 7336 16838
rect 7360 16836 7416 16838
rect 10478 28314 10534 28316
rect 10558 28314 10614 28316
rect 10638 28314 10694 28316
rect 10718 28314 10774 28316
rect 10478 28262 10524 28314
rect 10524 28262 10534 28314
rect 10558 28262 10588 28314
rect 10588 28262 10600 28314
rect 10600 28262 10614 28314
rect 10638 28262 10652 28314
rect 10652 28262 10664 28314
rect 10664 28262 10694 28314
rect 10718 28262 10728 28314
rect 10728 28262 10774 28314
rect 10478 28260 10534 28262
rect 10558 28260 10614 28262
rect 10638 28260 10694 28262
rect 10718 28260 10774 28262
rect 8482 17176 8538 17232
rect 3762 15258 3818 15260
rect 3842 15258 3898 15260
rect 3922 15258 3978 15260
rect 4002 15258 4058 15260
rect 3762 15206 3808 15258
rect 3808 15206 3818 15258
rect 3842 15206 3872 15258
rect 3872 15206 3884 15258
rect 3884 15206 3898 15258
rect 3922 15206 3936 15258
rect 3936 15206 3948 15258
rect 3948 15206 3978 15258
rect 4002 15206 4012 15258
rect 4012 15206 4058 15258
rect 3762 15204 3818 15206
rect 3842 15204 3898 15206
rect 3922 15204 3978 15206
rect 4002 15204 4058 15206
rect 3762 14170 3818 14172
rect 3842 14170 3898 14172
rect 3922 14170 3978 14172
rect 4002 14170 4058 14172
rect 3762 14118 3808 14170
rect 3808 14118 3818 14170
rect 3842 14118 3872 14170
rect 3872 14118 3884 14170
rect 3884 14118 3898 14170
rect 3922 14118 3936 14170
rect 3936 14118 3948 14170
rect 3948 14118 3978 14170
rect 4002 14118 4012 14170
rect 4012 14118 4058 14170
rect 3762 14116 3818 14118
rect 3842 14116 3898 14118
rect 3922 14116 3978 14118
rect 4002 14116 4058 14118
rect 3762 13082 3818 13084
rect 3842 13082 3898 13084
rect 3922 13082 3978 13084
rect 4002 13082 4058 13084
rect 3762 13030 3808 13082
rect 3808 13030 3818 13082
rect 3842 13030 3872 13082
rect 3872 13030 3884 13082
rect 3884 13030 3898 13082
rect 3922 13030 3936 13082
rect 3936 13030 3948 13082
rect 3948 13030 3978 13082
rect 4002 13030 4012 13082
rect 4012 13030 4058 13082
rect 3762 13028 3818 13030
rect 3842 13028 3898 13030
rect 3922 13028 3978 13030
rect 4002 13028 4058 13030
rect 3762 11994 3818 11996
rect 3842 11994 3898 11996
rect 3922 11994 3978 11996
rect 4002 11994 4058 11996
rect 3762 11942 3808 11994
rect 3808 11942 3818 11994
rect 3842 11942 3872 11994
rect 3872 11942 3884 11994
rect 3884 11942 3898 11994
rect 3922 11942 3936 11994
rect 3936 11942 3948 11994
rect 3948 11942 3978 11994
rect 4002 11942 4012 11994
rect 4012 11942 4058 11994
rect 3762 11940 3818 11942
rect 3842 11940 3898 11942
rect 3922 11940 3978 11942
rect 4002 11940 4058 11942
rect 3762 10906 3818 10908
rect 3842 10906 3898 10908
rect 3922 10906 3978 10908
rect 4002 10906 4058 10908
rect 3762 10854 3808 10906
rect 3808 10854 3818 10906
rect 3842 10854 3872 10906
rect 3872 10854 3884 10906
rect 3884 10854 3898 10906
rect 3922 10854 3936 10906
rect 3936 10854 3948 10906
rect 3948 10854 3978 10906
rect 4002 10854 4012 10906
rect 4012 10854 4058 10906
rect 3762 10852 3818 10854
rect 3842 10852 3898 10854
rect 3922 10852 3978 10854
rect 4002 10852 4058 10854
rect 3762 9818 3818 9820
rect 3842 9818 3898 9820
rect 3922 9818 3978 9820
rect 4002 9818 4058 9820
rect 3762 9766 3808 9818
rect 3808 9766 3818 9818
rect 3842 9766 3872 9818
rect 3872 9766 3884 9818
rect 3884 9766 3898 9818
rect 3922 9766 3936 9818
rect 3936 9766 3948 9818
rect 3948 9766 3978 9818
rect 4002 9766 4012 9818
rect 4012 9766 4058 9818
rect 3762 9764 3818 9766
rect 3842 9764 3898 9766
rect 3922 9764 3978 9766
rect 4002 9764 4058 9766
rect 7120 15802 7176 15804
rect 7200 15802 7256 15804
rect 7280 15802 7336 15804
rect 7360 15802 7416 15804
rect 7120 15750 7166 15802
rect 7166 15750 7176 15802
rect 7200 15750 7230 15802
rect 7230 15750 7242 15802
rect 7242 15750 7256 15802
rect 7280 15750 7294 15802
rect 7294 15750 7306 15802
rect 7306 15750 7336 15802
rect 7360 15750 7370 15802
rect 7370 15750 7416 15802
rect 7120 15748 7176 15750
rect 7200 15748 7256 15750
rect 7280 15748 7336 15750
rect 7360 15748 7416 15750
rect 10478 27226 10534 27228
rect 10558 27226 10614 27228
rect 10638 27226 10694 27228
rect 10718 27226 10774 27228
rect 10478 27174 10524 27226
rect 10524 27174 10534 27226
rect 10558 27174 10588 27226
rect 10588 27174 10600 27226
rect 10600 27174 10614 27226
rect 10638 27174 10652 27226
rect 10652 27174 10664 27226
rect 10664 27174 10694 27226
rect 10718 27174 10728 27226
rect 10728 27174 10774 27226
rect 10478 27172 10534 27174
rect 10558 27172 10614 27174
rect 10638 27172 10694 27174
rect 10718 27172 10774 27174
rect 10478 26138 10534 26140
rect 10558 26138 10614 26140
rect 10638 26138 10694 26140
rect 10718 26138 10774 26140
rect 10478 26086 10524 26138
rect 10524 26086 10534 26138
rect 10558 26086 10588 26138
rect 10588 26086 10600 26138
rect 10600 26086 10614 26138
rect 10638 26086 10652 26138
rect 10652 26086 10664 26138
rect 10664 26086 10694 26138
rect 10718 26086 10728 26138
rect 10728 26086 10774 26138
rect 10478 26084 10534 26086
rect 10558 26084 10614 26086
rect 10638 26084 10694 26086
rect 10718 26084 10774 26086
rect 10478 25050 10534 25052
rect 10558 25050 10614 25052
rect 10638 25050 10694 25052
rect 10718 25050 10774 25052
rect 10478 24998 10524 25050
rect 10524 24998 10534 25050
rect 10558 24998 10588 25050
rect 10588 24998 10600 25050
rect 10600 24998 10614 25050
rect 10638 24998 10652 25050
rect 10652 24998 10664 25050
rect 10664 24998 10694 25050
rect 10718 24998 10728 25050
rect 10728 24998 10774 25050
rect 10478 24996 10534 24998
rect 10558 24996 10614 24998
rect 10638 24996 10694 24998
rect 10718 24996 10774 24998
rect 10478 23962 10534 23964
rect 10558 23962 10614 23964
rect 10638 23962 10694 23964
rect 10718 23962 10774 23964
rect 10478 23910 10524 23962
rect 10524 23910 10534 23962
rect 10558 23910 10588 23962
rect 10588 23910 10600 23962
rect 10600 23910 10614 23962
rect 10638 23910 10652 23962
rect 10652 23910 10664 23962
rect 10664 23910 10694 23962
rect 10718 23910 10728 23962
rect 10728 23910 10774 23962
rect 10478 23908 10534 23910
rect 10558 23908 10614 23910
rect 10638 23908 10694 23910
rect 10718 23908 10774 23910
rect 10478 22874 10534 22876
rect 10558 22874 10614 22876
rect 10638 22874 10694 22876
rect 10718 22874 10774 22876
rect 10478 22822 10524 22874
rect 10524 22822 10534 22874
rect 10558 22822 10588 22874
rect 10588 22822 10600 22874
rect 10600 22822 10614 22874
rect 10638 22822 10652 22874
rect 10652 22822 10664 22874
rect 10664 22822 10694 22874
rect 10718 22822 10728 22874
rect 10728 22822 10774 22874
rect 10478 22820 10534 22822
rect 10558 22820 10614 22822
rect 10638 22820 10694 22822
rect 10718 22820 10774 22822
rect 10478 21786 10534 21788
rect 10558 21786 10614 21788
rect 10638 21786 10694 21788
rect 10718 21786 10774 21788
rect 10478 21734 10524 21786
rect 10524 21734 10534 21786
rect 10558 21734 10588 21786
rect 10588 21734 10600 21786
rect 10600 21734 10614 21786
rect 10638 21734 10652 21786
rect 10652 21734 10664 21786
rect 10664 21734 10694 21786
rect 10718 21734 10728 21786
rect 10728 21734 10774 21786
rect 10478 21732 10534 21734
rect 10558 21732 10614 21734
rect 10638 21732 10694 21734
rect 10718 21732 10774 21734
rect 10478 20698 10534 20700
rect 10558 20698 10614 20700
rect 10638 20698 10694 20700
rect 10718 20698 10774 20700
rect 10478 20646 10524 20698
rect 10524 20646 10534 20698
rect 10558 20646 10588 20698
rect 10588 20646 10600 20698
rect 10600 20646 10614 20698
rect 10638 20646 10652 20698
rect 10652 20646 10664 20698
rect 10664 20646 10694 20698
rect 10718 20646 10728 20698
rect 10728 20646 10774 20698
rect 10478 20644 10534 20646
rect 10558 20644 10614 20646
rect 10638 20644 10694 20646
rect 10718 20644 10774 20646
rect 7120 14714 7176 14716
rect 7200 14714 7256 14716
rect 7280 14714 7336 14716
rect 7360 14714 7416 14716
rect 7120 14662 7166 14714
rect 7166 14662 7176 14714
rect 7200 14662 7230 14714
rect 7230 14662 7242 14714
rect 7242 14662 7256 14714
rect 7280 14662 7294 14714
rect 7294 14662 7306 14714
rect 7306 14662 7336 14714
rect 7360 14662 7370 14714
rect 7370 14662 7416 14714
rect 7120 14660 7176 14662
rect 7200 14660 7256 14662
rect 7280 14660 7336 14662
rect 7360 14660 7416 14662
rect 7120 13626 7176 13628
rect 7200 13626 7256 13628
rect 7280 13626 7336 13628
rect 7360 13626 7416 13628
rect 7120 13574 7166 13626
rect 7166 13574 7176 13626
rect 7200 13574 7230 13626
rect 7230 13574 7242 13626
rect 7242 13574 7256 13626
rect 7280 13574 7294 13626
rect 7294 13574 7306 13626
rect 7306 13574 7336 13626
rect 7360 13574 7370 13626
rect 7370 13574 7416 13626
rect 7120 13572 7176 13574
rect 7200 13572 7256 13574
rect 7280 13572 7336 13574
rect 7360 13572 7416 13574
rect 7120 12538 7176 12540
rect 7200 12538 7256 12540
rect 7280 12538 7336 12540
rect 7360 12538 7416 12540
rect 7120 12486 7166 12538
rect 7166 12486 7176 12538
rect 7200 12486 7230 12538
rect 7230 12486 7242 12538
rect 7242 12486 7256 12538
rect 7280 12486 7294 12538
rect 7294 12486 7306 12538
rect 7306 12486 7336 12538
rect 7360 12486 7370 12538
rect 7370 12486 7416 12538
rect 7120 12484 7176 12486
rect 7200 12484 7256 12486
rect 7280 12484 7336 12486
rect 7360 12484 7416 12486
rect 7120 11450 7176 11452
rect 7200 11450 7256 11452
rect 7280 11450 7336 11452
rect 7360 11450 7416 11452
rect 7120 11398 7166 11450
rect 7166 11398 7176 11450
rect 7200 11398 7230 11450
rect 7230 11398 7242 11450
rect 7242 11398 7256 11450
rect 7280 11398 7294 11450
rect 7294 11398 7306 11450
rect 7306 11398 7336 11450
rect 7360 11398 7370 11450
rect 7370 11398 7416 11450
rect 7120 11396 7176 11398
rect 7200 11396 7256 11398
rect 7280 11396 7336 11398
rect 7360 11396 7416 11398
rect 7120 10362 7176 10364
rect 7200 10362 7256 10364
rect 7280 10362 7336 10364
rect 7360 10362 7416 10364
rect 7120 10310 7166 10362
rect 7166 10310 7176 10362
rect 7200 10310 7230 10362
rect 7230 10310 7242 10362
rect 7242 10310 7256 10362
rect 7280 10310 7294 10362
rect 7294 10310 7306 10362
rect 7306 10310 7336 10362
rect 7360 10310 7370 10362
rect 7370 10310 7416 10362
rect 7120 10308 7176 10310
rect 7200 10308 7256 10310
rect 7280 10308 7336 10310
rect 7360 10308 7416 10310
rect 10478 19610 10534 19612
rect 10558 19610 10614 19612
rect 10638 19610 10694 19612
rect 10718 19610 10774 19612
rect 10478 19558 10524 19610
rect 10524 19558 10534 19610
rect 10558 19558 10588 19610
rect 10588 19558 10600 19610
rect 10600 19558 10614 19610
rect 10638 19558 10652 19610
rect 10652 19558 10664 19610
rect 10664 19558 10694 19610
rect 10718 19558 10728 19610
rect 10728 19558 10774 19610
rect 10478 19556 10534 19558
rect 10558 19556 10614 19558
rect 10638 19556 10694 19558
rect 10718 19556 10774 19558
rect 10478 18522 10534 18524
rect 10558 18522 10614 18524
rect 10638 18522 10694 18524
rect 10718 18522 10774 18524
rect 10478 18470 10524 18522
rect 10524 18470 10534 18522
rect 10558 18470 10588 18522
rect 10588 18470 10600 18522
rect 10600 18470 10614 18522
rect 10638 18470 10652 18522
rect 10652 18470 10664 18522
rect 10664 18470 10694 18522
rect 10718 18470 10728 18522
rect 10728 18470 10774 18522
rect 10478 18468 10534 18470
rect 10558 18468 10614 18470
rect 10638 18468 10694 18470
rect 10718 18468 10774 18470
rect 10966 21936 11022 21992
rect 10478 17434 10534 17436
rect 10558 17434 10614 17436
rect 10638 17434 10694 17436
rect 10718 17434 10774 17436
rect 10478 17382 10524 17434
rect 10524 17382 10534 17434
rect 10558 17382 10588 17434
rect 10588 17382 10600 17434
rect 10600 17382 10614 17434
rect 10638 17382 10652 17434
rect 10652 17382 10664 17434
rect 10664 17382 10694 17434
rect 10718 17382 10728 17434
rect 10728 17382 10774 17434
rect 10478 17380 10534 17382
rect 10558 17380 10614 17382
rect 10638 17380 10694 17382
rect 10718 17380 10774 17382
rect 10506 17176 10562 17232
rect 10478 16346 10534 16348
rect 10558 16346 10614 16348
rect 10638 16346 10694 16348
rect 10718 16346 10774 16348
rect 10478 16294 10524 16346
rect 10524 16294 10534 16346
rect 10558 16294 10588 16346
rect 10588 16294 10600 16346
rect 10600 16294 10614 16346
rect 10638 16294 10652 16346
rect 10652 16294 10664 16346
rect 10664 16294 10694 16346
rect 10718 16294 10728 16346
rect 10728 16294 10774 16346
rect 10478 16292 10534 16294
rect 10558 16292 10614 16294
rect 10638 16292 10694 16294
rect 10718 16292 10774 16294
rect 10690 15972 10746 16008
rect 10690 15952 10692 15972
rect 10692 15952 10744 15972
rect 10744 15952 10746 15972
rect 9862 14320 9918 14376
rect 7120 9274 7176 9276
rect 7200 9274 7256 9276
rect 7280 9274 7336 9276
rect 7360 9274 7416 9276
rect 7120 9222 7166 9274
rect 7166 9222 7176 9274
rect 7200 9222 7230 9274
rect 7230 9222 7242 9274
rect 7242 9222 7256 9274
rect 7280 9222 7294 9274
rect 7294 9222 7306 9274
rect 7306 9222 7336 9274
rect 7360 9222 7370 9274
rect 7370 9222 7416 9274
rect 7120 9220 7176 9222
rect 7200 9220 7256 9222
rect 7280 9220 7336 9222
rect 7360 9220 7416 9222
rect 3762 8730 3818 8732
rect 3842 8730 3898 8732
rect 3922 8730 3978 8732
rect 4002 8730 4058 8732
rect 3762 8678 3808 8730
rect 3808 8678 3818 8730
rect 3842 8678 3872 8730
rect 3872 8678 3884 8730
rect 3884 8678 3898 8730
rect 3922 8678 3936 8730
rect 3936 8678 3948 8730
rect 3948 8678 3978 8730
rect 4002 8678 4012 8730
rect 4012 8678 4058 8730
rect 3762 8676 3818 8678
rect 3842 8676 3898 8678
rect 3922 8676 3978 8678
rect 4002 8676 4058 8678
rect 3762 7642 3818 7644
rect 3842 7642 3898 7644
rect 3922 7642 3978 7644
rect 4002 7642 4058 7644
rect 3762 7590 3808 7642
rect 3808 7590 3818 7642
rect 3842 7590 3872 7642
rect 3872 7590 3884 7642
rect 3884 7590 3898 7642
rect 3922 7590 3936 7642
rect 3936 7590 3948 7642
rect 3948 7590 3978 7642
rect 4002 7590 4012 7642
rect 4012 7590 4058 7642
rect 3762 7588 3818 7590
rect 3842 7588 3898 7590
rect 3922 7588 3978 7590
rect 4002 7588 4058 7590
rect 3762 6554 3818 6556
rect 3842 6554 3898 6556
rect 3922 6554 3978 6556
rect 4002 6554 4058 6556
rect 3762 6502 3808 6554
rect 3808 6502 3818 6554
rect 3842 6502 3872 6554
rect 3872 6502 3884 6554
rect 3884 6502 3898 6554
rect 3922 6502 3936 6554
rect 3936 6502 3948 6554
rect 3948 6502 3978 6554
rect 4002 6502 4012 6554
rect 4012 6502 4058 6554
rect 3762 6500 3818 6502
rect 3842 6500 3898 6502
rect 3922 6500 3978 6502
rect 4002 6500 4058 6502
rect 10230 14320 10286 14376
rect 10478 15258 10534 15260
rect 10558 15258 10614 15260
rect 10638 15258 10694 15260
rect 10718 15258 10774 15260
rect 10478 15206 10524 15258
rect 10524 15206 10534 15258
rect 10558 15206 10588 15258
rect 10588 15206 10600 15258
rect 10600 15206 10614 15258
rect 10638 15206 10652 15258
rect 10652 15206 10664 15258
rect 10664 15206 10694 15258
rect 10718 15206 10728 15258
rect 10728 15206 10774 15258
rect 10478 15204 10534 15206
rect 10558 15204 10614 15206
rect 10638 15204 10694 15206
rect 10718 15204 10774 15206
rect 10478 14170 10534 14172
rect 10558 14170 10614 14172
rect 10638 14170 10694 14172
rect 10718 14170 10774 14172
rect 10478 14118 10524 14170
rect 10524 14118 10534 14170
rect 10558 14118 10588 14170
rect 10588 14118 10600 14170
rect 10600 14118 10614 14170
rect 10638 14118 10652 14170
rect 10652 14118 10664 14170
rect 10664 14118 10694 14170
rect 10718 14118 10728 14170
rect 10728 14118 10774 14170
rect 10478 14116 10534 14118
rect 10558 14116 10614 14118
rect 10638 14116 10694 14118
rect 10718 14116 10774 14118
rect 10478 13082 10534 13084
rect 10558 13082 10614 13084
rect 10638 13082 10694 13084
rect 10718 13082 10774 13084
rect 10478 13030 10524 13082
rect 10524 13030 10534 13082
rect 10558 13030 10588 13082
rect 10588 13030 10600 13082
rect 10600 13030 10614 13082
rect 10638 13030 10652 13082
rect 10652 13030 10664 13082
rect 10664 13030 10694 13082
rect 10718 13030 10728 13082
rect 10728 13030 10774 13082
rect 10478 13028 10534 13030
rect 10558 13028 10614 13030
rect 10638 13028 10694 13030
rect 10718 13028 10774 13030
rect 10478 11994 10534 11996
rect 10558 11994 10614 11996
rect 10638 11994 10694 11996
rect 10718 11994 10774 11996
rect 10478 11942 10524 11994
rect 10524 11942 10534 11994
rect 10558 11942 10588 11994
rect 10588 11942 10600 11994
rect 10600 11942 10614 11994
rect 10638 11942 10652 11994
rect 10652 11942 10664 11994
rect 10664 11942 10694 11994
rect 10718 11942 10728 11994
rect 10728 11942 10774 11994
rect 10478 11940 10534 11942
rect 10558 11940 10614 11942
rect 10638 11940 10694 11942
rect 10718 11940 10774 11942
rect 10478 10906 10534 10908
rect 10558 10906 10614 10908
rect 10638 10906 10694 10908
rect 10718 10906 10774 10908
rect 10478 10854 10524 10906
rect 10524 10854 10534 10906
rect 10558 10854 10588 10906
rect 10588 10854 10600 10906
rect 10600 10854 10614 10906
rect 10638 10854 10652 10906
rect 10652 10854 10664 10906
rect 10664 10854 10694 10906
rect 10718 10854 10728 10906
rect 10728 10854 10774 10906
rect 10478 10852 10534 10854
rect 10558 10852 10614 10854
rect 10638 10852 10694 10854
rect 10718 10852 10774 10854
rect 10478 9818 10534 9820
rect 10558 9818 10614 9820
rect 10638 9818 10694 9820
rect 10718 9818 10774 9820
rect 10478 9766 10524 9818
rect 10524 9766 10534 9818
rect 10558 9766 10588 9818
rect 10588 9766 10600 9818
rect 10600 9766 10614 9818
rect 10638 9766 10652 9818
rect 10652 9766 10664 9818
rect 10664 9766 10694 9818
rect 10718 9766 10728 9818
rect 10728 9766 10774 9818
rect 10478 9764 10534 9766
rect 10558 9764 10614 9766
rect 10638 9764 10694 9766
rect 10718 9764 10774 9766
rect 7120 8186 7176 8188
rect 7200 8186 7256 8188
rect 7280 8186 7336 8188
rect 7360 8186 7416 8188
rect 7120 8134 7166 8186
rect 7166 8134 7176 8186
rect 7200 8134 7230 8186
rect 7230 8134 7242 8186
rect 7242 8134 7256 8186
rect 7280 8134 7294 8186
rect 7294 8134 7306 8186
rect 7306 8134 7336 8186
rect 7360 8134 7370 8186
rect 7370 8134 7416 8186
rect 7120 8132 7176 8134
rect 7200 8132 7256 8134
rect 7280 8132 7336 8134
rect 7360 8132 7416 8134
rect 7120 7098 7176 7100
rect 7200 7098 7256 7100
rect 7280 7098 7336 7100
rect 7360 7098 7416 7100
rect 7120 7046 7166 7098
rect 7166 7046 7176 7098
rect 7200 7046 7230 7098
rect 7230 7046 7242 7098
rect 7242 7046 7256 7098
rect 7280 7046 7294 7098
rect 7294 7046 7306 7098
rect 7306 7046 7336 7098
rect 7360 7046 7370 7098
rect 7370 7046 7416 7098
rect 7120 7044 7176 7046
rect 7200 7044 7256 7046
rect 7280 7044 7336 7046
rect 7360 7044 7416 7046
rect 7120 6010 7176 6012
rect 7200 6010 7256 6012
rect 7280 6010 7336 6012
rect 7360 6010 7416 6012
rect 7120 5958 7166 6010
rect 7166 5958 7176 6010
rect 7200 5958 7230 6010
rect 7230 5958 7242 6010
rect 7242 5958 7256 6010
rect 7280 5958 7294 6010
rect 7294 5958 7306 6010
rect 7306 5958 7336 6010
rect 7360 5958 7370 6010
rect 7370 5958 7416 6010
rect 7120 5956 7176 5958
rect 7200 5956 7256 5958
rect 7280 5956 7336 5958
rect 7360 5956 7416 5958
rect 9862 7268 9918 7304
rect 9862 7248 9864 7268
rect 9864 7248 9916 7268
rect 9916 7248 9918 7268
rect 10478 8730 10534 8732
rect 10558 8730 10614 8732
rect 10638 8730 10694 8732
rect 10718 8730 10774 8732
rect 10478 8678 10524 8730
rect 10524 8678 10534 8730
rect 10558 8678 10588 8730
rect 10588 8678 10600 8730
rect 10600 8678 10614 8730
rect 10638 8678 10652 8730
rect 10652 8678 10664 8730
rect 10664 8678 10694 8730
rect 10718 8678 10728 8730
rect 10728 8678 10774 8730
rect 10478 8676 10534 8678
rect 10558 8676 10614 8678
rect 10638 8676 10694 8678
rect 10718 8676 10774 8678
rect 10478 7642 10534 7644
rect 10558 7642 10614 7644
rect 10638 7642 10694 7644
rect 10718 7642 10774 7644
rect 10478 7590 10524 7642
rect 10524 7590 10534 7642
rect 10558 7590 10588 7642
rect 10588 7590 10600 7642
rect 10600 7590 10614 7642
rect 10638 7590 10652 7642
rect 10652 7590 10664 7642
rect 10664 7590 10694 7642
rect 10718 7590 10728 7642
rect 10728 7590 10774 7642
rect 10478 7588 10534 7590
rect 10558 7588 10614 7590
rect 10638 7588 10694 7590
rect 10718 7588 10774 7590
rect 2962 3984 3018 4040
rect 3762 5466 3818 5468
rect 3842 5466 3898 5468
rect 3922 5466 3978 5468
rect 4002 5466 4058 5468
rect 3762 5414 3808 5466
rect 3808 5414 3818 5466
rect 3842 5414 3872 5466
rect 3872 5414 3884 5466
rect 3884 5414 3898 5466
rect 3922 5414 3936 5466
rect 3936 5414 3948 5466
rect 3948 5414 3978 5466
rect 4002 5414 4012 5466
rect 4012 5414 4058 5466
rect 3762 5412 3818 5414
rect 3842 5412 3898 5414
rect 3922 5412 3978 5414
rect 4002 5412 4058 5414
rect 3762 4378 3818 4380
rect 3842 4378 3898 4380
rect 3922 4378 3978 4380
rect 4002 4378 4058 4380
rect 3762 4326 3808 4378
rect 3808 4326 3818 4378
rect 3842 4326 3872 4378
rect 3872 4326 3884 4378
rect 3884 4326 3898 4378
rect 3922 4326 3936 4378
rect 3936 4326 3948 4378
rect 3948 4326 3978 4378
rect 4002 4326 4012 4378
rect 4012 4326 4058 4378
rect 3762 4324 3818 4326
rect 3842 4324 3898 4326
rect 3922 4324 3978 4326
rect 4002 4324 4058 4326
rect 3606 3984 3662 4040
rect 3762 3290 3818 3292
rect 3842 3290 3898 3292
rect 3922 3290 3978 3292
rect 4002 3290 4058 3292
rect 3762 3238 3808 3290
rect 3808 3238 3818 3290
rect 3842 3238 3872 3290
rect 3872 3238 3884 3290
rect 3884 3238 3898 3290
rect 3922 3238 3936 3290
rect 3936 3238 3948 3290
rect 3948 3238 3978 3290
rect 4002 3238 4012 3290
rect 4012 3238 4058 3290
rect 3762 3236 3818 3238
rect 3842 3236 3898 3238
rect 3922 3236 3978 3238
rect 4002 3236 4058 3238
rect 4434 2488 4490 2544
rect 4986 3440 5042 3496
rect 3762 2202 3818 2204
rect 3842 2202 3898 2204
rect 3922 2202 3978 2204
rect 4002 2202 4058 2204
rect 3762 2150 3808 2202
rect 3808 2150 3818 2202
rect 3842 2150 3872 2202
rect 3872 2150 3884 2202
rect 3884 2150 3898 2202
rect 3922 2150 3936 2202
rect 3936 2150 3948 2202
rect 3948 2150 3978 2202
rect 4002 2150 4012 2202
rect 4012 2150 4058 2202
rect 3762 2148 3818 2150
rect 3842 2148 3898 2150
rect 3922 2148 3978 2150
rect 4002 2148 4058 2150
rect 3762 1114 3818 1116
rect 3842 1114 3898 1116
rect 3922 1114 3978 1116
rect 4002 1114 4058 1116
rect 3762 1062 3808 1114
rect 3808 1062 3818 1114
rect 3842 1062 3872 1114
rect 3872 1062 3884 1114
rect 3884 1062 3898 1114
rect 3922 1062 3936 1114
rect 3936 1062 3948 1114
rect 3948 1062 3978 1114
rect 4002 1062 4012 1114
rect 4012 1062 4058 1114
rect 3762 1060 3818 1062
rect 3842 1060 3898 1062
rect 3922 1060 3978 1062
rect 4002 1060 4058 1062
rect 5446 2488 5502 2544
rect 7120 4922 7176 4924
rect 7200 4922 7256 4924
rect 7280 4922 7336 4924
rect 7360 4922 7416 4924
rect 7120 4870 7166 4922
rect 7166 4870 7176 4922
rect 7200 4870 7230 4922
rect 7230 4870 7242 4922
rect 7242 4870 7256 4922
rect 7280 4870 7294 4922
rect 7294 4870 7306 4922
rect 7306 4870 7336 4922
rect 7360 4870 7370 4922
rect 7370 4870 7416 4922
rect 7120 4868 7176 4870
rect 7200 4868 7256 4870
rect 7280 4868 7336 4870
rect 7360 4868 7416 4870
rect 7654 3984 7710 4040
rect 7120 3834 7176 3836
rect 7200 3834 7256 3836
rect 7280 3834 7336 3836
rect 7360 3834 7416 3836
rect 7120 3782 7166 3834
rect 7166 3782 7176 3834
rect 7200 3782 7230 3834
rect 7230 3782 7242 3834
rect 7242 3782 7256 3834
rect 7280 3782 7294 3834
rect 7294 3782 7306 3834
rect 7306 3782 7336 3834
rect 7360 3782 7370 3834
rect 7370 3782 7416 3834
rect 7120 3780 7176 3782
rect 7200 3780 7256 3782
rect 7280 3780 7336 3782
rect 7360 3780 7416 3782
rect 6458 2508 6514 2544
rect 6458 2488 6460 2508
rect 6460 2488 6512 2508
rect 6512 2488 6514 2508
rect 7194 3440 7250 3496
rect 7120 2746 7176 2748
rect 7200 2746 7256 2748
rect 7280 2746 7336 2748
rect 7360 2746 7416 2748
rect 7120 2694 7166 2746
rect 7166 2694 7176 2746
rect 7200 2694 7230 2746
rect 7230 2694 7242 2746
rect 7242 2694 7256 2746
rect 7280 2694 7294 2746
rect 7294 2694 7306 2746
rect 7306 2694 7336 2746
rect 7360 2694 7370 2746
rect 7370 2694 7416 2746
rect 7120 2692 7176 2694
rect 7200 2692 7256 2694
rect 7280 2692 7336 2694
rect 7360 2692 7416 2694
rect 7120 1658 7176 1660
rect 7200 1658 7256 1660
rect 7280 1658 7336 1660
rect 7360 1658 7416 1660
rect 7120 1606 7166 1658
rect 7166 1606 7176 1658
rect 7200 1606 7230 1658
rect 7230 1606 7242 1658
rect 7242 1606 7256 1658
rect 7280 1606 7294 1658
rect 7294 1606 7306 1658
rect 7306 1606 7336 1658
rect 7360 1606 7370 1658
rect 7370 1606 7416 1658
rect 7120 1604 7176 1606
rect 7200 1604 7256 1606
rect 7280 1604 7336 1606
rect 7360 1604 7416 1606
rect 7120 570 7176 572
rect 7200 570 7256 572
rect 7280 570 7336 572
rect 7360 570 7416 572
rect 7120 518 7166 570
rect 7166 518 7176 570
rect 7200 518 7230 570
rect 7230 518 7242 570
rect 7242 518 7256 570
rect 7280 518 7294 570
rect 7294 518 7306 570
rect 7306 518 7336 570
rect 7360 518 7370 570
rect 7370 518 7416 570
rect 7120 516 7176 518
rect 7200 516 7256 518
rect 7280 516 7336 518
rect 7360 516 7416 518
rect 10478 6554 10534 6556
rect 10558 6554 10614 6556
rect 10638 6554 10694 6556
rect 10718 6554 10774 6556
rect 10478 6502 10524 6554
rect 10524 6502 10534 6554
rect 10558 6502 10588 6554
rect 10588 6502 10600 6554
rect 10600 6502 10614 6554
rect 10638 6502 10652 6554
rect 10652 6502 10664 6554
rect 10664 6502 10694 6554
rect 10718 6502 10728 6554
rect 10728 6502 10774 6554
rect 10478 6500 10534 6502
rect 10558 6500 10614 6502
rect 10638 6500 10694 6502
rect 10718 6500 10774 6502
rect 10478 5466 10534 5468
rect 10558 5466 10614 5468
rect 10638 5466 10694 5468
rect 10718 5466 10774 5468
rect 10478 5414 10524 5466
rect 10524 5414 10534 5466
rect 10558 5414 10588 5466
rect 10588 5414 10600 5466
rect 10600 5414 10614 5466
rect 10638 5414 10652 5466
rect 10652 5414 10664 5466
rect 10664 5414 10694 5466
rect 10718 5414 10728 5466
rect 10728 5414 10774 5466
rect 10478 5412 10534 5414
rect 10558 5412 10614 5414
rect 10638 5412 10694 5414
rect 10718 5412 10774 5414
rect 13836 31034 13892 31036
rect 13916 31034 13972 31036
rect 13996 31034 14052 31036
rect 14076 31034 14132 31036
rect 13836 30982 13882 31034
rect 13882 30982 13892 31034
rect 13916 30982 13946 31034
rect 13946 30982 13958 31034
rect 13958 30982 13972 31034
rect 13996 30982 14010 31034
rect 14010 30982 14022 31034
rect 14022 30982 14052 31034
rect 14076 30982 14086 31034
rect 14086 30982 14132 31034
rect 13836 30980 13892 30982
rect 13916 30980 13972 30982
rect 13996 30980 14052 30982
rect 14076 30980 14132 30982
rect 12990 19760 13046 19816
rect 12714 14320 12770 14376
rect 13836 29946 13892 29948
rect 13916 29946 13972 29948
rect 13996 29946 14052 29948
rect 14076 29946 14132 29948
rect 13836 29894 13882 29946
rect 13882 29894 13892 29946
rect 13916 29894 13946 29946
rect 13946 29894 13958 29946
rect 13958 29894 13972 29946
rect 13996 29894 14010 29946
rect 14010 29894 14022 29946
rect 14022 29894 14052 29946
rect 14076 29894 14086 29946
rect 14086 29894 14132 29946
rect 13836 29892 13892 29894
rect 13916 29892 13972 29894
rect 13996 29892 14052 29894
rect 14076 29892 14132 29894
rect 13836 28858 13892 28860
rect 13916 28858 13972 28860
rect 13996 28858 14052 28860
rect 14076 28858 14132 28860
rect 13836 28806 13882 28858
rect 13882 28806 13892 28858
rect 13916 28806 13946 28858
rect 13946 28806 13958 28858
rect 13958 28806 13972 28858
rect 13996 28806 14010 28858
rect 14010 28806 14022 28858
rect 14022 28806 14052 28858
rect 14076 28806 14086 28858
rect 14086 28806 14132 28858
rect 13836 28804 13892 28806
rect 13916 28804 13972 28806
rect 13996 28804 14052 28806
rect 14076 28804 14132 28806
rect 13836 27770 13892 27772
rect 13916 27770 13972 27772
rect 13996 27770 14052 27772
rect 14076 27770 14132 27772
rect 13836 27718 13882 27770
rect 13882 27718 13892 27770
rect 13916 27718 13946 27770
rect 13946 27718 13958 27770
rect 13958 27718 13972 27770
rect 13996 27718 14010 27770
rect 14010 27718 14022 27770
rect 14022 27718 14052 27770
rect 14076 27718 14086 27770
rect 14086 27718 14132 27770
rect 13836 27716 13892 27718
rect 13916 27716 13972 27718
rect 13996 27716 14052 27718
rect 14076 27716 14132 27718
rect 13836 26682 13892 26684
rect 13916 26682 13972 26684
rect 13996 26682 14052 26684
rect 14076 26682 14132 26684
rect 13836 26630 13882 26682
rect 13882 26630 13892 26682
rect 13916 26630 13946 26682
rect 13946 26630 13958 26682
rect 13958 26630 13972 26682
rect 13996 26630 14010 26682
rect 14010 26630 14022 26682
rect 14022 26630 14052 26682
rect 14076 26630 14086 26682
rect 14086 26630 14132 26682
rect 13836 26628 13892 26630
rect 13916 26628 13972 26630
rect 13996 26628 14052 26630
rect 14076 26628 14132 26630
rect 13836 25594 13892 25596
rect 13916 25594 13972 25596
rect 13996 25594 14052 25596
rect 14076 25594 14132 25596
rect 13836 25542 13882 25594
rect 13882 25542 13892 25594
rect 13916 25542 13946 25594
rect 13946 25542 13958 25594
rect 13958 25542 13972 25594
rect 13996 25542 14010 25594
rect 14010 25542 14022 25594
rect 14022 25542 14052 25594
rect 14076 25542 14086 25594
rect 14086 25542 14132 25594
rect 13836 25540 13892 25542
rect 13916 25540 13972 25542
rect 13996 25540 14052 25542
rect 14076 25540 14132 25542
rect 17194 30490 17250 30492
rect 17274 30490 17330 30492
rect 17354 30490 17410 30492
rect 17434 30490 17490 30492
rect 17194 30438 17240 30490
rect 17240 30438 17250 30490
rect 17274 30438 17304 30490
rect 17304 30438 17316 30490
rect 17316 30438 17330 30490
rect 17354 30438 17368 30490
rect 17368 30438 17380 30490
rect 17380 30438 17410 30490
rect 17434 30438 17444 30490
rect 17444 30438 17490 30490
rect 17194 30436 17250 30438
rect 17274 30436 17330 30438
rect 17354 30436 17410 30438
rect 17434 30436 17490 30438
rect 16578 29552 16634 29608
rect 17194 29402 17250 29404
rect 17274 29402 17330 29404
rect 17354 29402 17410 29404
rect 17434 29402 17490 29404
rect 17194 29350 17240 29402
rect 17240 29350 17250 29402
rect 17274 29350 17304 29402
rect 17304 29350 17316 29402
rect 17316 29350 17330 29402
rect 17354 29350 17368 29402
rect 17368 29350 17380 29402
rect 17380 29350 17410 29402
rect 17434 29350 17444 29402
rect 17444 29350 17490 29402
rect 17194 29348 17250 29350
rect 17274 29348 17330 29350
rect 17354 29348 17410 29350
rect 17434 29348 17490 29350
rect 16670 27820 16672 27840
rect 16672 27820 16724 27840
rect 16724 27820 16726 27840
rect 16670 27784 16726 27820
rect 13836 24506 13892 24508
rect 13916 24506 13972 24508
rect 13996 24506 14052 24508
rect 14076 24506 14132 24508
rect 13836 24454 13882 24506
rect 13882 24454 13892 24506
rect 13916 24454 13946 24506
rect 13946 24454 13958 24506
rect 13958 24454 13972 24506
rect 13996 24454 14010 24506
rect 14010 24454 14022 24506
rect 14022 24454 14052 24506
rect 14076 24454 14086 24506
rect 14086 24454 14132 24506
rect 13836 24452 13892 24454
rect 13916 24452 13972 24454
rect 13996 24452 14052 24454
rect 14076 24452 14132 24454
rect 13836 23418 13892 23420
rect 13916 23418 13972 23420
rect 13996 23418 14052 23420
rect 14076 23418 14132 23420
rect 13836 23366 13882 23418
rect 13882 23366 13892 23418
rect 13916 23366 13946 23418
rect 13946 23366 13958 23418
rect 13958 23366 13972 23418
rect 13996 23366 14010 23418
rect 14010 23366 14022 23418
rect 14022 23366 14052 23418
rect 14076 23366 14086 23418
rect 14086 23366 14132 23418
rect 13836 23364 13892 23366
rect 13916 23364 13972 23366
rect 13996 23364 14052 23366
rect 14076 23364 14132 23366
rect 13836 22330 13892 22332
rect 13916 22330 13972 22332
rect 13996 22330 14052 22332
rect 14076 22330 14132 22332
rect 13836 22278 13882 22330
rect 13882 22278 13892 22330
rect 13916 22278 13946 22330
rect 13946 22278 13958 22330
rect 13958 22278 13972 22330
rect 13996 22278 14010 22330
rect 14010 22278 14022 22330
rect 14022 22278 14052 22330
rect 14076 22278 14086 22330
rect 14086 22278 14132 22330
rect 13836 22276 13892 22278
rect 13916 22276 13972 22278
rect 13996 22276 14052 22278
rect 14076 22276 14132 22278
rect 13836 21242 13892 21244
rect 13916 21242 13972 21244
rect 13996 21242 14052 21244
rect 14076 21242 14132 21244
rect 13836 21190 13882 21242
rect 13882 21190 13892 21242
rect 13916 21190 13946 21242
rect 13946 21190 13958 21242
rect 13958 21190 13972 21242
rect 13996 21190 14010 21242
rect 14010 21190 14022 21242
rect 14022 21190 14052 21242
rect 14076 21190 14086 21242
rect 14086 21190 14132 21242
rect 13836 21188 13892 21190
rect 13916 21188 13972 21190
rect 13996 21188 14052 21190
rect 14076 21188 14132 21190
rect 13836 20154 13892 20156
rect 13916 20154 13972 20156
rect 13996 20154 14052 20156
rect 14076 20154 14132 20156
rect 13836 20102 13882 20154
rect 13882 20102 13892 20154
rect 13916 20102 13946 20154
rect 13946 20102 13958 20154
rect 13958 20102 13972 20154
rect 13996 20102 14010 20154
rect 14010 20102 14022 20154
rect 14022 20102 14052 20154
rect 14076 20102 14086 20154
rect 14086 20102 14132 20154
rect 13836 20100 13892 20102
rect 13916 20100 13972 20102
rect 13996 20100 14052 20102
rect 14076 20100 14132 20102
rect 13836 19066 13892 19068
rect 13916 19066 13972 19068
rect 13996 19066 14052 19068
rect 14076 19066 14132 19068
rect 13836 19014 13882 19066
rect 13882 19014 13892 19066
rect 13916 19014 13946 19066
rect 13946 19014 13958 19066
rect 13958 19014 13972 19066
rect 13996 19014 14010 19066
rect 14010 19014 14022 19066
rect 14022 19014 14052 19066
rect 14076 19014 14086 19066
rect 14086 19014 14132 19066
rect 13836 19012 13892 19014
rect 13916 19012 13972 19014
rect 13996 19012 14052 19014
rect 14076 19012 14132 19014
rect 13836 17978 13892 17980
rect 13916 17978 13972 17980
rect 13996 17978 14052 17980
rect 14076 17978 14132 17980
rect 13836 17926 13882 17978
rect 13882 17926 13892 17978
rect 13916 17926 13946 17978
rect 13946 17926 13958 17978
rect 13958 17926 13972 17978
rect 13996 17926 14010 17978
rect 14010 17926 14022 17978
rect 14022 17926 14052 17978
rect 14076 17926 14086 17978
rect 14086 17926 14132 17978
rect 13836 17924 13892 17926
rect 13916 17924 13972 17926
rect 13996 17924 14052 17926
rect 14076 17924 14132 17926
rect 11886 7112 11942 7168
rect 10478 4378 10534 4380
rect 10558 4378 10614 4380
rect 10638 4378 10694 4380
rect 10718 4378 10774 4380
rect 10478 4326 10524 4378
rect 10524 4326 10534 4378
rect 10558 4326 10588 4378
rect 10588 4326 10600 4378
rect 10600 4326 10614 4378
rect 10638 4326 10652 4378
rect 10652 4326 10664 4378
rect 10664 4326 10694 4378
rect 10718 4326 10728 4378
rect 10728 4326 10774 4378
rect 10478 4324 10534 4326
rect 10558 4324 10614 4326
rect 10638 4324 10694 4326
rect 10718 4324 10774 4326
rect 10782 3576 10838 3632
rect 10478 3290 10534 3292
rect 10558 3290 10614 3292
rect 10638 3290 10694 3292
rect 10718 3290 10774 3292
rect 10478 3238 10524 3290
rect 10524 3238 10534 3290
rect 10558 3238 10588 3290
rect 10588 3238 10600 3290
rect 10600 3238 10614 3290
rect 10638 3238 10652 3290
rect 10652 3238 10664 3290
rect 10664 3238 10694 3290
rect 10718 3238 10728 3290
rect 10728 3238 10774 3290
rect 10478 3236 10534 3238
rect 10558 3236 10614 3238
rect 10638 3236 10694 3238
rect 10718 3236 10774 3238
rect 10478 2202 10534 2204
rect 10558 2202 10614 2204
rect 10638 2202 10694 2204
rect 10718 2202 10774 2204
rect 10478 2150 10524 2202
rect 10524 2150 10534 2202
rect 10558 2150 10588 2202
rect 10588 2150 10600 2202
rect 10600 2150 10614 2202
rect 10638 2150 10652 2202
rect 10652 2150 10664 2202
rect 10664 2150 10694 2202
rect 10718 2150 10728 2202
rect 10728 2150 10774 2202
rect 10478 2148 10534 2150
rect 10558 2148 10614 2150
rect 10638 2148 10694 2150
rect 10718 2148 10774 2150
rect 12990 7112 13046 7168
rect 13836 16890 13892 16892
rect 13916 16890 13972 16892
rect 13996 16890 14052 16892
rect 14076 16890 14132 16892
rect 13836 16838 13882 16890
rect 13882 16838 13892 16890
rect 13916 16838 13946 16890
rect 13946 16838 13958 16890
rect 13958 16838 13972 16890
rect 13996 16838 14010 16890
rect 14010 16838 14022 16890
rect 14022 16838 14052 16890
rect 14076 16838 14086 16890
rect 14086 16838 14132 16890
rect 13836 16836 13892 16838
rect 13916 16836 13972 16838
rect 13996 16836 14052 16838
rect 14076 16836 14132 16838
rect 13836 15802 13892 15804
rect 13916 15802 13972 15804
rect 13996 15802 14052 15804
rect 14076 15802 14132 15804
rect 13836 15750 13882 15802
rect 13882 15750 13892 15802
rect 13916 15750 13946 15802
rect 13946 15750 13958 15802
rect 13958 15750 13972 15802
rect 13996 15750 14010 15802
rect 14010 15750 14022 15802
rect 14022 15750 14052 15802
rect 14076 15750 14086 15802
rect 14086 15750 14132 15802
rect 13836 15748 13892 15750
rect 13916 15748 13972 15750
rect 13996 15748 14052 15750
rect 14076 15748 14132 15750
rect 15566 24792 15622 24848
rect 17194 28314 17250 28316
rect 17274 28314 17330 28316
rect 17354 28314 17410 28316
rect 17434 28314 17490 28316
rect 17194 28262 17240 28314
rect 17240 28262 17250 28314
rect 17274 28262 17304 28314
rect 17304 28262 17316 28314
rect 17316 28262 17330 28314
rect 17354 28262 17368 28314
rect 17368 28262 17380 28314
rect 17380 28262 17410 28314
rect 17434 28262 17444 28314
rect 17444 28262 17490 28314
rect 17194 28260 17250 28262
rect 17274 28260 17330 28262
rect 17354 28260 17410 28262
rect 17434 28260 17490 28262
rect 17222 27820 17224 27840
rect 17224 27820 17276 27840
rect 17276 27820 17278 27840
rect 17222 27784 17278 27820
rect 17222 27668 17278 27704
rect 17222 27648 17224 27668
rect 17224 27648 17276 27668
rect 17276 27648 17278 27668
rect 17590 27648 17646 27704
rect 17194 27226 17250 27228
rect 17274 27226 17330 27228
rect 17354 27226 17410 27228
rect 17434 27226 17490 27228
rect 17194 27174 17240 27226
rect 17240 27174 17250 27226
rect 17274 27174 17304 27226
rect 17304 27174 17316 27226
rect 17316 27174 17330 27226
rect 17354 27174 17368 27226
rect 17368 27174 17380 27226
rect 17380 27174 17410 27226
rect 17434 27174 17444 27226
rect 17444 27174 17490 27226
rect 17194 27172 17250 27174
rect 17274 27172 17330 27174
rect 17354 27172 17410 27174
rect 17434 27172 17490 27174
rect 17194 26138 17250 26140
rect 17274 26138 17330 26140
rect 17354 26138 17410 26140
rect 17434 26138 17490 26140
rect 17194 26086 17240 26138
rect 17240 26086 17250 26138
rect 17274 26086 17304 26138
rect 17304 26086 17316 26138
rect 17316 26086 17330 26138
rect 17354 26086 17368 26138
rect 17368 26086 17380 26138
rect 17380 26086 17410 26138
rect 17434 26086 17444 26138
rect 17444 26086 17490 26138
rect 17194 26084 17250 26086
rect 17274 26084 17330 26086
rect 17354 26084 17410 26086
rect 17434 26084 17490 26086
rect 14922 19352 14978 19408
rect 14646 15952 14702 16008
rect 13836 14714 13892 14716
rect 13916 14714 13972 14716
rect 13996 14714 14052 14716
rect 14076 14714 14132 14716
rect 13836 14662 13882 14714
rect 13882 14662 13892 14714
rect 13916 14662 13946 14714
rect 13946 14662 13958 14714
rect 13958 14662 13972 14714
rect 13996 14662 14010 14714
rect 14010 14662 14022 14714
rect 14022 14662 14052 14714
rect 14076 14662 14086 14714
rect 14086 14662 14132 14714
rect 13836 14660 13892 14662
rect 13916 14660 13972 14662
rect 13996 14660 14052 14662
rect 14076 14660 14132 14662
rect 13836 13626 13892 13628
rect 13916 13626 13972 13628
rect 13996 13626 14052 13628
rect 14076 13626 14132 13628
rect 13836 13574 13882 13626
rect 13882 13574 13892 13626
rect 13916 13574 13946 13626
rect 13946 13574 13958 13626
rect 13958 13574 13972 13626
rect 13996 13574 14010 13626
rect 14010 13574 14022 13626
rect 14022 13574 14052 13626
rect 14076 13574 14086 13626
rect 14086 13574 14132 13626
rect 13836 13572 13892 13574
rect 13916 13572 13972 13574
rect 13996 13572 14052 13574
rect 14076 13572 14132 13574
rect 13836 12538 13892 12540
rect 13916 12538 13972 12540
rect 13996 12538 14052 12540
rect 14076 12538 14132 12540
rect 13836 12486 13882 12538
rect 13882 12486 13892 12538
rect 13916 12486 13946 12538
rect 13946 12486 13958 12538
rect 13958 12486 13972 12538
rect 13996 12486 14010 12538
rect 14010 12486 14022 12538
rect 14022 12486 14052 12538
rect 14076 12486 14086 12538
rect 14086 12486 14132 12538
rect 13836 12484 13892 12486
rect 13916 12484 13972 12486
rect 13996 12484 14052 12486
rect 14076 12484 14132 12486
rect 13836 11450 13892 11452
rect 13916 11450 13972 11452
rect 13996 11450 14052 11452
rect 14076 11450 14132 11452
rect 13836 11398 13882 11450
rect 13882 11398 13892 11450
rect 13916 11398 13946 11450
rect 13946 11398 13958 11450
rect 13958 11398 13972 11450
rect 13996 11398 14010 11450
rect 14010 11398 14022 11450
rect 14022 11398 14052 11450
rect 14076 11398 14086 11450
rect 14086 11398 14132 11450
rect 13836 11396 13892 11398
rect 13916 11396 13972 11398
rect 13996 11396 14052 11398
rect 14076 11396 14132 11398
rect 13836 10362 13892 10364
rect 13916 10362 13972 10364
rect 13996 10362 14052 10364
rect 14076 10362 14132 10364
rect 13836 10310 13882 10362
rect 13882 10310 13892 10362
rect 13916 10310 13946 10362
rect 13946 10310 13958 10362
rect 13958 10310 13972 10362
rect 13996 10310 14010 10362
rect 14010 10310 14022 10362
rect 14022 10310 14052 10362
rect 14076 10310 14086 10362
rect 14086 10310 14132 10362
rect 13836 10308 13892 10310
rect 13916 10308 13972 10310
rect 13996 10308 14052 10310
rect 14076 10308 14132 10310
rect 15474 15988 15476 16008
rect 15476 15988 15528 16008
rect 15528 15988 15530 16008
rect 15474 15952 15530 15988
rect 17194 25050 17250 25052
rect 17274 25050 17330 25052
rect 17354 25050 17410 25052
rect 17434 25050 17490 25052
rect 17194 24998 17240 25050
rect 17240 24998 17250 25050
rect 17274 24998 17304 25050
rect 17304 24998 17316 25050
rect 17316 24998 17330 25050
rect 17354 24998 17368 25050
rect 17368 24998 17380 25050
rect 17380 24998 17410 25050
rect 17434 24998 17444 25050
rect 17444 24998 17490 25050
rect 17194 24996 17250 24998
rect 17274 24996 17330 24998
rect 17354 24996 17410 24998
rect 17434 24996 17490 24998
rect 18970 29552 19026 29608
rect 17194 23962 17250 23964
rect 17274 23962 17330 23964
rect 17354 23962 17410 23964
rect 17434 23962 17490 23964
rect 17194 23910 17240 23962
rect 17240 23910 17250 23962
rect 17274 23910 17304 23962
rect 17304 23910 17316 23962
rect 17316 23910 17330 23962
rect 17354 23910 17368 23962
rect 17368 23910 17380 23962
rect 17380 23910 17410 23962
rect 17434 23910 17444 23962
rect 17444 23910 17490 23962
rect 17194 23908 17250 23910
rect 17274 23908 17330 23910
rect 17354 23908 17410 23910
rect 17434 23908 17490 23910
rect 17194 22874 17250 22876
rect 17274 22874 17330 22876
rect 17354 22874 17410 22876
rect 17434 22874 17490 22876
rect 17194 22822 17240 22874
rect 17240 22822 17250 22874
rect 17274 22822 17304 22874
rect 17304 22822 17316 22874
rect 17316 22822 17330 22874
rect 17354 22822 17368 22874
rect 17368 22822 17380 22874
rect 17380 22822 17410 22874
rect 17434 22822 17444 22874
rect 17444 22822 17490 22874
rect 17194 22820 17250 22822
rect 17274 22820 17330 22822
rect 17354 22820 17410 22822
rect 17434 22820 17490 22822
rect 16118 17060 16174 17096
rect 16118 17040 16120 17060
rect 16120 17040 16172 17060
rect 16172 17040 16174 17060
rect 13836 9274 13892 9276
rect 13916 9274 13972 9276
rect 13996 9274 14052 9276
rect 14076 9274 14132 9276
rect 13836 9222 13882 9274
rect 13882 9222 13892 9274
rect 13916 9222 13946 9274
rect 13946 9222 13958 9274
rect 13958 9222 13972 9274
rect 13996 9222 14010 9274
rect 14010 9222 14022 9274
rect 14022 9222 14052 9274
rect 14076 9222 14086 9274
rect 14086 9222 14132 9274
rect 13836 9220 13892 9222
rect 13916 9220 13972 9222
rect 13996 9220 14052 9222
rect 14076 9220 14132 9222
rect 13836 8186 13892 8188
rect 13916 8186 13972 8188
rect 13996 8186 14052 8188
rect 14076 8186 14132 8188
rect 13836 8134 13882 8186
rect 13882 8134 13892 8186
rect 13916 8134 13946 8186
rect 13946 8134 13958 8186
rect 13958 8134 13972 8186
rect 13996 8134 14010 8186
rect 14010 8134 14022 8186
rect 14022 8134 14052 8186
rect 14076 8134 14086 8186
rect 14086 8134 14132 8186
rect 13836 8132 13892 8134
rect 13916 8132 13972 8134
rect 13996 8132 14052 8134
rect 14076 8132 14132 8134
rect 13836 7098 13892 7100
rect 13916 7098 13972 7100
rect 13996 7098 14052 7100
rect 14076 7098 14132 7100
rect 13836 7046 13882 7098
rect 13882 7046 13892 7098
rect 13916 7046 13946 7098
rect 13946 7046 13958 7098
rect 13958 7046 13972 7098
rect 13996 7046 14010 7098
rect 14010 7046 14022 7098
rect 14022 7046 14052 7098
rect 14076 7046 14086 7098
rect 14086 7046 14132 7098
rect 13836 7044 13892 7046
rect 13916 7044 13972 7046
rect 13996 7044 14052 7046
rect 14076 7044 14132 7046
rect 14094 6160 14150 6216
rect 13836 6010 13892 6012
rect 13916 6010 13972 6012
rect 13996 6010 14052 6012
rect 14076 6010 14132 6012
rect 13836 5958 13882 6010
rect 13882 5958 13892 6010
rect 13916 5958 13946 6010
rect 13946 5958 13958 6010
rect 13958 5958 13972 6010
rect 13996 5958 14010 6010
rect 14010 5958 14022 6010
rect 14022 5958 14052 6010
rect 14076 5958 14086 6010
rect 14086 5958 14132 6010
rect 13836 5956 13892 5958
rect 13916 5956 13972 5958
rect 13996 5956 14052 5958
rect 14076 5956 14132 5958
rect 17194 21786 17250 21788
rect 17274 21786 17330 21788
rect 17354 21786 17410 21788
rect 17434 21786 17490 21788
rect 17194 21734 17240 21786
rect 17240 21734 17250 21786
rect 17274 21734 17304 21786
rect 17304 21734 17316 21786
rect 17316 21734 17330 21786
rect 17354 21734 17368 21786
rect 17368 21734 17380 21786
rect 17380 21734 17410 21786
rect 17434 21734 17444 21786
rect 17444 21734 17490 21786
rect 17194 21732 17250 21734
rect 17274 21732 17330 21734
rect 17354 21732 17410 21734
rect 17434 21732 17490 21734
rect 17194 20698 17250 20700
rect 17274 20698 17330 20700
rect 17354 20698 17410 20700
rect 17434 20698 17490 20700
rect 17194 20646 17240 20698
rect 17240 20646 17250 20698
rect 17274 20646 17304 20698
rect 17304 20646 17316 20698
rect 17316 20646 17330 20698
rect 17354 20646 17368 20698
rect 17368 20646 17380 20698
rect 17380 20646 17410 20698
rect 17434 20646 17444 20698
rect 17444 20646 17490 20698
rect 17194 20644 17250 20646
rect 17274 20644 17330 20646
rect 17354 20644 17410 20646
rect 17434 20644 17490 20646
rect 17194 19610 17250 19612
rect 17274 19610 17330 19612
rect 17354 19610 17410 19612
rect 17434 19610 17490 19612
rect 17194 19558 17240 19610
rect 17240 19558 17250 19610
rect 17274 19558 17304 19610
rect 17304 19558 17316 19610
rect 17316 19558 17330 19610
rect 17354 19558 17368 19610
rect 17368 19558 17380 19610
rect 17380 19558 17410 19610
rect 17434 19558 17444 19610
rect 17444 19558 17490 19610
rect 17194 19556 17250 19558
rect 17274 19556 17330 19558
rect 17354 19556 17410 19558
rect 17434 19556 17490 19558
rect 20552 31034 20608 31036
rect 20632 31034 20688 31036
rect 20712 31034 20768 31036
rect 20792 31034 20848 31036
rect 20552 30982 20598 31034
rect 20598 30982 20608 31034
rect 20632 30982 20662 31034
rect 20662 30982 20674 31034
rect 20674 30982 20688 31034
rect 20712 30982 20726 31034
rect 20726 30982 20738 31034
rect 20738 30982 20768 31034
rect 20792 30982 20802 31034
rect 20802 30982 20848 31034
rect 20552 30980 20608 30982
rect 20632 30980 20688 30982
rect 20712 30980 20768 30982
rect 20792 30980 20848 30982
rect 20810 30096 20866 30152
rect 20552 29946 20608 29948
rect 20632 29946 20688 29948
rect 20712 29946 20768 29948
rect 20792 29946 20848 29948
rect 20552 29894 20598 29946
rect 20598 29894 20608 29946
rect 20632 29894 20662 29946
rect 20662 29894 20674 29946
rect 20674 29894 20688 29946
rect 20712 29894 20726 29946
rect 20726 29894 20738 29946
rect 20738 29894 20768 29946
rect 20792 29894 20802 29946
rect 20802 29894 20848 29946
rect 20552 29892 20608 29894
rect 20632 29892 20688 29894
rect 20712 29892 20768 29894
rect 20792 29892 20848 29894
rect 20552 28858 20608 28860
rect 20632 28858 20688 28860
rect 20712 28858 20768 28860
rect 20792 28858 20848 28860
rect 20552 28806 20598 28858
rect 20598 28806 20608 28858
rect 20632 28806 20662 28858
rect 20662 28806 20674 28858
rect 20674 28806 20688 28858
rect 20712 28806 20726 28858
rect 20726 28806 20738 28858
rect 20738 28806 20768 28858
rect 20792 28806 20802 28858
rect 20802 28806 20848 28858
rect 20552 28804 20608 28806
rect 20632 28804 20688 28806
rect 20712 28804 20768 28806
rect 20792 28804 20848 28806
rect 20552 27770 20608 27772
rect 20632 27770 20688 27772
rect 20712 27770 20768 27772
rect 20792 27770 20848 27772
rect 20552 27718 20598 27770
rect 20598 27718 20608 27770
rect 20632 27718 20662 27770
rect 20662 27718 20674 27770
rect 20674 27718 20688 27770
rect 20712 27718 20726 27770
rect 20726 27718 20738 27770
rect 20738 27718 20768 27770
rect 20792 27718 20802 27770
rect 20802 27718 20848 27770
rect 20552 27716 20608 27718
rect 20632 27716 20688 27718
rect 20712 27716 20768 27718
rect 20792 27716 20848 27718
rect 20552 26682 20608 26684
rect 20632 26682 20688 26684
rect 20712 26682 20768 26684
rect 20792 26682 20848 26684
rect 20552 26630 20598 26682
rect 20598 26630 20608 26682
rect 20632 26630 20662 26682
rect 20662 26630 20674 26682
rect 20674 26630 20688 26682
rect 20712 26630 20726 26682
rect 20726 26630 20738 26682
rect 20738 26630 20768 26682
rect 20792 26630 20802 26682
rect 20802 26630 20848 26682
rect 20552 26628 20608 26630
rect 20632 26628 20688 26630
rect 20712 26628 20768 26630
rect 20792 26628 20848 26630
rect 20552 25594 20608 25596
rect 20632 25594 20688 25596
rect 20712 25594 20768 25596
rect 20792 25594 20848 25596
rect 20552 25542 20598 25594
rect 20598 25542 20608 25594
rect 20632 25542 20662 25594
rect 20662 25542 20674 25594
rect 20674 25542 20688 25594
rect 20712 25542 20726 25594
rect 20726 25542 20738 25594
rect 20738 25542 20768 25594
rect 20792 25542 20802 25594
rect 20802 25542 20848 25594
rect 20552 25540 20608 25542
rect 20632 25540 20688 25542
rect 20712 25540 20768 25542
rect 20792 25540 20848 25542
rect 18050 21972 18052 21992
rect 18052 21972 18104 21992
rect 18104 21972 18106 21992
rect 18050 21936 18106 21972
rect 17194 18522 17250 18524
rect 17274 18522 17330 18524
rect 17354 18522 17410 18524
rect 17434 18522 17490 18524
rect 17194 18470 17240 18522
rect 17240 18470 17250 18522
rect 17274 18470 17304 18522
rect 17304 18470 17316 18522
rect 17316 18470 17330 18522
rect 17354 18470 17368 18522
rect 17368 18470 17380 18522
rect 17380 18470 17410 18522
rect 17434 18470 17444 18522
rect 17444 18470 17490 18522
rect 17194 18468 17250 18470
rect 17274 18468 17330 18470
rect 17354 18468 17410 18470
rect 17434 18468 17490 18470
rect 18326 19352 18382 19408
rect 17194 17434 17250 17436
rect 17274 17434 17330 17436
rect 17354 17434 17410 17436
rect 17434 17434 17490 17436
rect 17194 17382 17240 17434
rect 17240 17382 17250 17434
rect 17274 17382 17304 17434
rect 17304 17382 17316 17434
rect 17316 17382 17330 17434
rect 17354 17382 17368 17434
rect 17368 17382 17380 17434
rect 17380 17382 17410 17434
rect 17434 17382 17444 17434
rect 17444 17382 17490 17434
rect 17194 17380 17250 17382
rect 17274 17380 17330 17382
rect 17354 17380 17410 17382
rect 17434 17380 17490 17382
rect 17194 16346 17250 16348
rect 17274 16346 17330 16348
rect 17354 16346 17410 16348
rect 17434 16346 17490 16348
rect 17194 16294 17240 16346
rect 17240 16294 17250 16346
rect 17274 16294 17304 16346
rect 17304 16294 17316 16346
rect 17316 16294 17330 16346
rect 17354 16294 17368 16346
rect 17368 16294 17380 16346
rect 17380 16294 17410 16346
rect 17434 16294 17444 16346
rect 17444 16294 17490 16346
rect 17194 16292 17250 16294
rect 17274 16292 17330 16294
rect 17354 16292 17410 16294
rect 17434 16292 17490 16294
rect 17194 15258 17250 15260
rect 17274 15258 17330 15260
rect 17354 15258 17410 15260
rect 17434 15258 17490 15260
rect 17194 15206 17240 15258
rect 17240 15206 17250 15258
rect 17274 15206 17304 15258
rect 17304 15206 17316 15258
rect 17316 15206 17330 15258
rect 17354 15206 17368 15258
rect 17368 15206 17380 15258
rect 17380 15206 17410 15258
rect 17434 15206 17444 15258
rect 17444 15206 17490 15258
rect 17194 15204 17250 15206
rect 17274 15204 17330 15206
rect 17354 15204 17410 15206
rect 17434 15204 17490 15206
rect 17194 14170 17250 14172
rect 17274 14170 17330 14172
rect 17354 14170 17410 14172
rect 17434 14170 17490 14172
rect 17194 14118 17240 14170
rect 17240 14118 17250 14170
rect 17274 14118 17304 14170
rect 17304 14118 17316 14170
rect 17316 14118 17330 14170
rect 17354 14118 17368 14170
rect 17368 14118 17380 14170
rect 17380 14118 17410 14170
rect 17434 14118 17444 14170
rect 17444 14118 17490 14170
rect 17194 14116 17250 14118
rect 17274 14116 17330 14118
rect 17354 14116 17410 14118
rect 17434 14116 17490 14118
rect 18510 19760 18566 19816
rect 17194 13082 17250 13084
rect 17274 13082 17330 13084
rect 17354 13082 17410 13084
rect 17434 13082 17490 13084
rect 17194 13030 17240 13082
rect 17240 13030 17250 13082
rect 17274 13030 17304 13082
rect 17304 13030 17316 13082
rect 17316 13030 17330 13082
rect 17354 13030 17368 13082
rect 17368 13030 17380 13082
rect 17380 13030 17410 13082
rect 17434 13030 17444 13082
rect 17444 13030 17490 13082
rect 17194 13028 17250 13030
rect 17274 13028 17330 13030
rect 17354 13028 17410 13030
rect 17434 13028 17490 13030
rect 17194 11994 17250 11996
rect 17274 11994 17330 11996
rect 17354 11994 17410 11996
rect 17434 11994 17490 11996
rect 17194 11942 17240 11994
rect 17240 11942 17250 11994
rect 17274 11942 17304 11994
rect 17304 11942 17316 11994
rect 17316 11942 17330 11994
rect 17354 11942 17368 11994
rect 17368 11942 17380 11994
rect 17380 11942 17410 11994
rect 17434 11942 17444 11994
rect 17444 11942 17490 11994
rect 17194 11940 17250 11942
rect 17274 11940 17330 11942
rect 17354 11940 17410 11942
rect 17434 11940 17490 11942
rect 17194 10906 17250 10908
rect 17274 10906 17330 10908
rect 17354 10906 17410 10908
rect 17434 10906 17490 10908
rect 17194 10854 17240 10906
rect 17240 10854 17250 10906
rect 17274 10854 17304 10906
rect 17304 10854 17316 10906
rect 17316 10854 17330 10906
rect 17354 10854 17368 10906
rect 17368 10854 17380 10906
rect 17380 10854 17410 10906
rect 17434 10854 17444 10906
rect 17444 10854 17490 10906
rect 17194 10852 17250 10854
rect 17274 10852 17330 10854
rect 17354 10852 17410 10854
rect 17434 10852 17490 10854
rect 17194 9818 17250 9820
rect 17274 9818 17330 9820
rect 17354 9818 17410 9820
rect 17434 9818 17490 9820
rect 17194 9766 17240 9818
rect 17240 9766 17250 9818
rect 17274 9766 17304 9818
rect 17304 9766 17316 9818
rect 17316 9766 17330 9818
rect 17354 9766 17368 9818
rect 17368 9766 17380 9818
rect 17380 9766 17410 9818
rect 17434 9766 17444 9818
rect 17444 9766 17490 9818
rect 17194 9764 17250 9766
rect 17274 9764 17330 9766
rect 17354 9764 17410 9766
rect 17434 9764 17490 9766
rect 18326 14320 18382 14376
rect 20552 24506 20608 24508
rect 20632 24506 20688 24508
rect 20712 24506 20768 24508
rect 20792 24506 20848 24508
rect 20552 24454 20598 24506
rect 20598 24454 20608 24506
rect 20632 24454 20662 24506
rect 20662 24454 20674 24506
rect 20674 24454 20688 24506
rect 20712 24454 20726 24506
rect 20726 24454 20738 24506
rect 20738 24454 20768 24506
rect 20792 24454 20802 24506
rect 20802 24454 20848 24506
rect 20552 24452 20608 24454
rect 20632 24452 20688 24454
rect 20712 24452 20768 24454
rect 20792 24452 20848 24454
rect 20552 23418 20608 23420
rect 20632 23418 20688 23420
rect 20712 23418 20768 23420
rect 20792 23418 20848 23420
rect 20552 23366 20598 23418
rect 20598 23366 20608 23418
rect 20632 23366 20662 23418
rect 20662 23366 20674 23418
rect 20674 23366 20688 23418
rect 20712 23366 20726 23418
rect 20726 23366 20738 23418
rect 20738 23366 20768 23418
rect 20792 23366 20802 23418
rect 20802 23366 20848 23418
rect 20552 23364 20608 23366
rect 20632 23364 20688 23366
rect 20712 23364 20768 23366
rect 20792 23364 20848 23366
rect 20552 22330 20608 22332
rect 20632 22330 20688 22332
rect 20712 22330 20768 22332
rect 20792 22330 20848 22332
rect 20552 22278 20598 22330
rect 20598 22278 20608 22330
rect 20632 22278 20662 22330
rect 20662 22278 20674 22330
rect 20674 22278 20688 22330
rect 20712 22278 20726 22330
rect 20726 22278 20738 22330
rect 20738 22278 20768 22330
rect 20792 22278 20802 22330
rect 20802 22278 20848 22330
rect 20552 22276 20608 22278
rect 20632 22276 20688 22278
rect 20712 22276 20768 22278
rect 20792 22276 20848 22278
rect 20552 21242 20608 21244
rect 20632 21242 20688 21244
rect 20712 21242 20768 21244
rect 20792 21242 20848 21244
rect 20552 21190 20598 21242
rect 20598 21190 20608 21242
rect 20632 21190 20662 21242
rect 20662 21190 20674 21242
rect 20674 21190 20688 21242
rect 20712 21190 20726 21242
rect 20726 21190 20738 21242
rect 20738 21190 20768 21242
rect 20792 21190 20802 21242
rect 20802 21190 20848 21242
rect 20552 21188 20608 21190
rect 20632 21188 20688 21190
rect 20712 21188 20768 21190
rect 20792 21188 20848 21190
rect 21270 27004 21272 27024
rect 21272 27004 21324 27024
rect 21324 27004 21326 27024
rect 21270 26968 21326 27004
rect 22834 29688 22890 29744
rect 21546 26560 21602 26616
rect 22926 29552 22982 29608
rect 23910 30490 23966 30492
rect 23990 30490 24046 30492
rect 24070 30490 24126 30492
rect 24150 30490 24206 30492
rect 23910 30438 23956 30490
rect 23956 30438 23966 30490
rect 23990 30438 24020 30490
rect 24020 30438 24032 30490
rect 24032 30438 24046 30490
rect 24070 30438 24084 30490
rect 24084 30438 24096 30490
rect 24096 30438 24126 30490
rect 24150 30438 24160 30490
rect 24160 30438 24206 30490
rect 23910 30436 23966 30438
rect 23990 30436 24046 30438
rect 24070 30436 24126 30438
rect 24150 30436 24206 30438
rect 23846 30096 23902 30152
rect 21822 26560 21878 26616
rect 20552 20154 20608 20156
rect 20632 20154 20688 20156
rect 20712 20154 20768 20156
rect 20792 20154 20848 20156
rect 20552 20102 20598 20154
rect 20598 20102 20608 20154
rect 20632 20102 20662 20154
rect 20662 20102 20674 20154
rect 20674 20102 20688 20154
rect 20712 20102 20726 20154
rect 20726 20102 20738 20154
rect 20738 20102 20768 20154
rect 20792 20102 20802 20154
rect 20802 20102 20848 20154
rect 20552 20100 20608 20102
rect 20632 20100 20688 20102
rect 20712 20100 20768 20102
rect 20792 20100 20848 20102
rect 14370 6452 14426 6488
rect 14370 6432 14372 6452
rect 14372 6432 14424 6452
rect 14424 6432 14426 6452
rect 13836 4922 13892 4924
rect 13916 4922 13972 4924
rect 13996 4922 14052 4924
rect 14076 4922 14132 4924
rect 13836 4870 13882 4922
rect 13882 4870 13892 4922
rect 13916 4870 13946 4922
rect 13946 4870 13958 4922
rect 13958 4870 13972 4922
rect 13996 4870 14010 4922
rect 14010 4870 14022 4922
rect 14022 4870 14052 4922
rect 14076 4870 14086 4922
rect 14086 4870 14132 4922
rect 13836 4868 13892 4870
rect 13916 4868 13972 4870
rect 13996 4868 14052 4870
rect 14076 4868 14132 4870
rect 13836 3834 13892 3836
rect 13916 3834 13972 3836
rect 13996 3834 14052 3836
rect 14076 3834 14132 3836
rect 13836 3782 13882 3834
rect 13882 3782 13892 3834
rect 13916 3782 13946 3834
rect 13946 3782 13958 3834
rect 13958 3782 13972 3834
rect 13996 3782 14010 3834
rect 14010 3782 14022 3834
rect 14022 3782 14052 3834
rect 14076 3782 14086 3834
rect 14086 3782 14132 3834
rect 13836 3780 13892 3782
rect 13916 3780 13972 3782
rect 13996 3780 14052 3782
rect 14076 3780 14132 3782
rect 13818 3304 13874 3360
rect 14370 3984 14426 4040
rect 17194 8730 17250 8732
rect 17274 8730 17330 8732
rect 17354 8730 17410 8732
rect 17434 8730 17490 8732
rect 17194 8678 17240 8730
rect 17240 8678 17250 8730
rect 17274 8678 17304 8730
rect 17304 8678 17316 8730
rect 17316 8678 17330 8730
rect 17354 8678 17368 8730
rect 17368 8678 17380 8730
rect 17380 8678 17410 8730
rect 17434 8678 17444 8730
rect 17444 8678 17490 8730
rect 17194 8676 17250 8678
rect 17274 8676 17330 8678
rect 17354 8676 17410 8678
rect 17434 8676 17490 8678
rect 20552 19066 20608 19068
rect 20632 19066 20688 19068
rect 20712 19066 20768 19068
rect 20792 19066 20848 19068
rect 20552 19014 20598 19066
rect 20598 19014 20608 19066
rect 20632 19014 20662 19066
rect 20662 19014 20674 19066
rect 20674 19014 20688 19066
rect 20712 19014 20726 19066
rect 20726 19014 20738 19066
rect 20738 19014 20768 19066
rect 20792 19014 20802 19066
rect 20802 19014 20848 19066
rect 20552 19012 20608 19014
rect 20632 19012 20688 19014
rect 20712 19012 20768 19014
rect 20792 19012 20848 19014
rect 20552 17978 20608 17980
rect 20632 17978 20688 17980
rect 20712 17978 20768 17980
rect 20792 17978 20848 17980
rect 20552 17926 20598 17978
rect 20598 17926 20608 17978
rect 20632 17926 20662 17978
rect 20662 17926 20674 17978
rect 20674 17926 20688 17978
rect 20712 17926 20726 17978
rect 20726 17926 20738 17978
rect 20738 17926 20768 17978
rect 20792 17926 20802 17978
rect 20802 17926 20848 17978
rect 20552 17924 20608 17926
rect 20632 17924 20688 17926
rect 20712 17924 20768 17926
rect 20792 17924 20848 17926
rect 20552 16890 20608 16892
rect 20632 16890 20688 16892
rect 20712 16890 20768 16892
rect 20792 16890 20848 16892
rect 20552 16838 20598 16890
rect 20598 16838 20608 16890
rect 20632 16838 20662 16890
rect 20662 16838 20674 16890
rect 20674 16838 20688 16890
rect 20712 16838 20726 16890
rect 20726 16838 20738 16890
rect 20738 16838 20768 16890
rect 20792 16838 20802 16890
rect 20802 16838 20848 16890
rect 20552 16836 20608 16838
rect 20632 16836 20688 16838
rect 20712 16836 20768 16838
rect 20792 16836 20848 16838
rect 20552 15802 20608 15804
rect 20632 15802 20688 15804
rect 20712 15802 20768 15804
rect 20792 15802 20848 15804
rect 20552 15750 20598 15802
rect 20598 15750 20608 15802
rect 20632 15750 20662 15802
rect 20662 15750 20674 15802
rect 20674 15750 20688 15802
rect 20712 15750 20726 15802
rect 20726 15750 20738 15802
rect 20738 15750 20768 15802
rect 20792 15750 20802 15802
rect 20802 15750 20848 15802
rect 20552 15748 20608 15750
rect 20632 15748 20688 15750
rect 20712 15748 20768 15750
rect 20792 15748 20848 15750
rect 23846 29552 23902 29608
rect 23910 29402 23966 29404
rect 23990 29402 24046 29404
rect 24070 29402 24126 29404
rect 24150 29402 24206 29404
rect 23910 29350 23956 29402
rect 23956 29350 23966 29402
rect 23990 29350 24020 29402
rect 24020 29350 24032 29402
rect 24032 29350 24046 29402
rect 24070 29350 24084 29402
rect 24084 29350 24096 29402
rect 24096 29350 24126 29402
rect 24150 29350 24160 29402
rect 24160 29350 24206 29402
rect 23910 29348 23966 29350
rect 23990 29348 24046 29350
rect 24070 29348 24126 29350
rect 24150 29348 24206 29350
rect 23910 28314 23966 28316
rect 23990 28314 24046 28316
rect 24070 28314 24126 28316
rect 24150 28314 24206 28316
rect 23910 28262 23956 28314
rect 23956 28262 23966 28314
rect 23990 28262 24020 28314
rect 24020 28262 24032 28314
rect 24032 28262 24046 28314
rect 24070 28262 24084 28314
rect 24084 28262 24096 28314
rect 24096 28262 24126 28314
rect 24150 28262 24160 28314
rect 24160 28262 24206 28314
rect 23910 28260 23966 28262
rect 23990 28260 24046 28262
rect 24070 28260 24126 28262
rect 24150 28260 24206 28262
rect 23478 26968 23534 27024
rect 23910 27226 23966 27228
rect 23990 27226 24046 27228
rect 24070 27226 24126 27228
rect 24150 27226 24206 27228
rect 23910 27174 23956 27226
rect 23956 27174 23966 27226
rect 23990 27174 24020 27226
rect 24020 27174 24032 27226
rect 24032 27174 24046 27226
rect 24070 27174 24084 27226
rect 24084 27174 24096 27226
rect 24096 27174 24126 27226
rect 24150 27174 24160 27226
rect 24160 27174 24206 27226
rect 23910 27172 23966 27174
rect 23990 27172 24046 27174
rect 24070 27172 24126 27174
rect 24150 27172 24206 27174
rect 23910 26138 23966 26140
rect 23990 26138 24046 26140
rect 24070 26138 24126 26140
rect 24150 26138 24206 26140
rect 23910 26086 23956 26138
rect 23956 26086 23966 26138
rect 23990 26086 24020 26138
rect 24020 26086 24032 26138
rect 24032 26086 24046 26138
rect 24070 26086 24084 26138
rect 24084 26086 24096 26138
rect 24096 26086 24126 26138
rect 24150 26086 24160 26138
rect 24160 26086 24206 26138
rect 23910 26084 23966 26086
rect 23990 26084 24046 26086
rect 24070 26084 24126 26086
rect 24150 26084 24206 26086
rect 23910 25050 23966 25052
rect 23990 25050 24046 25052
rect 24070 25050 24126 25052
rect 24150 25050 24206 25052
rect 23910 24998 23956 25050
rect 23956 24998 23966 25050
rect 23990 24998 24020 25050
rect 24020 24998 24032 25050
rect 24032 24998 24046 25050
rect 24070 24998 24084 25050
rect 24084 24998 24096 25050
rect 24096 24998 24126 25050
rect 24150 24998 24160 25050
rect 24160 24998 24206 25050
rect 23910 24996 23966 24998
rect 23990 24996 24046 24998
rect 24070 24996 24126 24998
rect 24150 24996 24206 24998
rect 20552 14714 20608 14716
rect 20632 14714 20688 14716
rect 20712 14714 20768 14716
rect 20792 14714 20848 14716
rect 20552 14662 20598 14714
rect 20598 14662 20608 14714
rect 20632 14662 20662 14714
rect 20662 14662 20674 14714
rect 20674 14662 20688 14714
rect 20712 14662 20726 14714
rect 20726 14662 20738 14714
rect 20738 14662 20768 14714
rect 20792 14662 20802 14714
rect 20802 14662 20848 14714
rect 20552 14660 20608 14662
rect 20632 14660 20688 14662
rect 20712 14660 20768 14662
rect 20792 14660 20848 14662
rect 20350 10532 20406 10568
rect 20350 10512 20352 10532
rect 20352 10512 20404 10532
rect 20404 10512 20406 10532
rect 17194 7642 17250 7644
rect 17274 7642 17330 7644
rect 17354 7642 17410 7644
rect 17434 7642 17490 7644
rect 17194 7590 17240 7642
rect 17240 7590 17250 7642
rect 17274 7590 17304 7642
rect 17304 7590 17316 7642
rect 17316 7590 17330 7642
rect 17354 7590 17368 7642
rect 17368 7590 17380 7642
rect 17380 7590 17410 7642
rect 17434 7590 17444 7642
rect 17444 7590 17490 7642
rect 17194 7588 17250 7590
rect 17274 7588 17330 7590
rect 17354 7588 17410 7590
rect 17434 7588 17490 7590
rect 15198 6432 15254 6488
rect 15106 6160 15162 6216
rect 17194 6554 17250 6556
rect 17274 6554 17330 6556
rect 17354 6554 17410 6556
rect 17434 6554 17490 6556
rect 17194 6502 17240 6554
rect 17240 6502 17250 6554
rect 17274 6502 17304 6554
rect 17304 6502 17316 6554
rect 17316 6502 17330 6554
rect 17354 6502 17368 6554
rect 17368 6502 17380 6554
rect 17380 6502 17410 6554
rect 17434 6502 17444 6554
rect 17444 6502 17490 6554
rect 17194 6500 17250 6502
rect 17274 6500 17330 6502
rect 17354 6500 17410 6502
rect 17434 6500 17490 6502
rect 20552 13626 20608 13628
rect 20632 13626 20688 13628
rect 20712 13626 20768 13628
rect 20792 13626 20848 13628
rect 20552 13574 20598 13626
rect 20598 13574 20608 13626
rect 20632 13574 20662 13626
rect 20662 13574 20674 13626
rect 20674 13574 20688 13626
rect 20712 13574 20726 13626
rect 20726 13574 20738 13626
rect 20738 13574 20768 13626
rect 20792 13574 20802 13626
rect 20802 13574 20848 13626
rect 20552 13572 20608 13574
rect 20632 13572 20688 13574
rect 20712 13572 20768 13574
rect 20792 13572 20848 13574
rect 20552 12538 20608 12540
rect 20632 12538 20688 12540
rect 20712 12538 20768 12540
rect 20792 12538 20848 12540
rect 20552 12486 20598 12538
rect 20598 12486 20608 12538
rect 20632 12486 20662 12538
rect 20662 12486 20674 12538
rect 20674 12486 20688 12538
rect 20712 12486 20726 12538
rect 20726 12486 20738 12538
rect 20738 12486 20768 12538
rect 20792 12486 20802 12538
rect 20802 12486 20848 12538
rect 20552 12484 20608 12486
rect 20632 12484 20688 12486
rect 20712 12484 20768 12486
rect 20792 12484 20848 12486
rect 20552 11450 20608 11452
rect 20632 11450 20688 11452
rect 20712 11450 20768 11452
rect 20792 11450 20848 11452
rect 20552 11398 20598 11450
rect 20598 11398 20608 11450
rect 20632 11398 20662 11450
rect 20662 11398 20674 11450
rect 20674 11398 20688 11450
rect 20712 11398 20726 11450
rect 20726 11398 20738 11450
rect 20738 11398 20768 11450
rect 20792 11398 20802 11450
rect 20802 11398 20848 11450
rect 20552 11396 20608 11398
rect 20632 11396 20688 11398
rect 20712 11396 20768 11398
rect 20792 11396 20848 11398
rect 20552 10362 20608 10364
rect 20632 10362 20688 10364
rect 20712 10362 20768 10364
rect 20792 10362 20848 10364
rect 20552 10310 20598 10362
rect 20598 10310 20608 10362
rect 20632 10310 20662 10362
rect 20662 10310 20674 10362
rect 20674 10310 20688 10362
rect 20712 10310 20726 10362
rect 20726 10310 20738 10362
rect 20738 10310 20768 10362
rect 20792 10310 20802 10362
rect 20802 10310 20848 10362
rect 20552 10308 20608 10310
rect 20632 10308 20688 10310
rect 20712 10308 20768 10310
rect 20792 10308 20848 10310
rect 20552 9274 20608 9276
rect 20632 9274 20688 9276
rect 20712 9274 20768 9276
rect 20792 9274 20848 9276
rect 20552 9222 20598 9274
rect 20598 9222 20608 9274
rect 20632 9222 20662 9274
rect 20662 9222 20674 9274
rect 20674 9222 20688 9274
rect 20712 9222 20726 9274
rect 20726 9222 20738 9274
rect 20738 9222 20768 9274
rect 20792 9222 20802 9274
rect 20802 9222 20848 9274
rect 20552 9220 20608 9222
rect 20632 9220 20688 9222
rect 20712 9220 20768 9222
rect 20792 9220 20848 9222
rect 20552 8186 20608 8188
rect 20632 8186 20688 8188
rect 20712 8186 20768 8188
rect 20792 8186 20848 8188
rect 20552 8134 20598 8186
rect 20598 8134 20608 8186
rect 20632 8134 20662 8186
rect 20662 8134 20674 8186
rect 20674 8134 20688 8186
rect 20712 8134 20726 8186
rect 20726 8134 20738 8186
rect 20738 8134 20768 8186
rect 20792 8134 20802 8186
rect 20802 8134 20848 8186
rect 20552 8132 20608 8134
rect 20632 8132 20688 8134
rect 20712 8132 20768 8134
rect 20792 8132 20848 8134
rect 17194 5466 17250 5468
rect 17274 5466 17330 5468
rect 17354 5466 17410 5468
rect 17434 5466 17490 5468
rect 17194 5414 17240 5466
rect 17240 5414 17250 5466
rect 17274 5414 17304 5466
rect 17304 5414 17316 5466
rect 17316 5414 17330 5466
rect 17354 5414 17368 5466
rect 17368 5414 17380 5466
rect 17380 5414 17410 5466
rect 17434 5414 17444 5466
rect 17444 5414 17490 5466
rect 17194 5412 17250 5414
rect 17274 5412 17330 5414
rect 17354 5412 17410 5414
rect 17434 5412 17490 5414
rect 13836 2746 13892 2748
rect 13916 2746 13972 2748
rect 13996 2746 14052 2748
rect 14076 2746 14132 2748
rect 13836 2694 13882 2746
rect 13882 2694 13892 2746
rect 13916 2694 13946 2746
rect 13946 2694 13958 2746
rect 13958 2694 13972 2746
rect 13996 2694 14010 2746
rect 14010 2694 14022 2746
rect 14022 2694 14052 2746
rect 14076 2694 14086 2746
rect 14086 2694 14132 2746
rect 13836 2692 13892 2694
rect 13916 2692 13972 2694
rect 13996 2692 14052 2694
rect 14076 2692 14132 2694
rect 10478 1114 10534 1116
rect 10558 1114 10614 1116
rect 10638 1114 10694 1116
rect 10718 1114 10774 1116
rect 10478 1062 10524 1114
rect 10524 1062 10534 1114
rect 10558 1062 10588 1114
rect 10588 1062 10600 1114
rect 10600 1062 10614 1114
rect 10638 1062 10652 1114
rect 10652 1062 10664 1114
rect 10664 1062 10694 1114
rect 10718 1062 10728 1114
rect 10728 1062 10774 1114
rect 10478 1060 10534 1062
rect 10558 1060 10614 1062
rect 10638 1060 10694 1062
rect 10718 1060 10774 1062
rect 14646 3440 14702 3496
rect 13836 1658 13892 1660
rect 13916 1658 13972 1660
rect 13996 1658 14052 1660
rect 14076 1658 14132 1660
rect 13836 1606 13882 1658
rect 13882 1606 13892 1658
rect 13916 1606 13946 1658
rect 13946 1606 13958 1658
rect 13958 1606 13972 1658
rect 13996 1606 14010 1658
rect 14010 1606 14022 1658
rect 14022 1606 14052 1658
rect 14076 1606 14086 1658
rect 14086 1606 14132 1658
rect 13836 1604 13892 1606
rect 13916 1604 13972 1606
rect 13996 1604 14052 1606
rect 14076 1604 14132 1606
rect 13836 570 13892 572
rect 13916 570 13972 572
rect 13996 570 14052 572
rect 14076 570 14132 572
rect 13836 518 13882 570
rect 13882 518 13892 570
rect 13916 518 13946 570
rect 13946 518 13958 570
rect 13958 518 13972 570
rect 13996 518 14010 570
rect 14010 518 14022 570
rect 14022 518 14052 570
rect 14076 518 14086 570
rect 14086 518 14132 570
rect 13836 516 13892 518
rect 13916 516 13972 518
rect 13996 516 14052 518
rect 14076 516 14132 518
rect 14922 3304 14978 3360
rect 17194 4378 17250 4380
rect 17274 4378 17330 4380
rect 17354 4378 17410 4380
rect 17434 4378 17490 4380
rect 17194 4326 17240 4378
rect 17240 4326 17250 4378
rect 17274 4326 17304 4378
rect 17304 4326 17316 4378
rect 17316 4326 17330 4378
rect 17354 4326 17368 4378
rect 17368 4326 17380 4378
rect 17380 4326 17410 4378
rect 17434 4326 17444 4378
rect 17444 4326 17490 4378
rect 17194 4324 17250 4326
rect 17274 4324 17330 4326
rect 17354 4324 17410 4326
rect 17434 4324 17490 4326
rect 15750 3596 15806 3632
rect 15750 3576 15752 3596
rect 15752 3576 15804 3596
rect 15804 3576 15806 3596
rect 17194 3290 17250 3292
rect 17274 3290 17330 3292
rect 17354 3290 17410 3292
rect 17434 3290 17490 3292
rect 17194 3238 17240 3290
rect 17240 3238 17250 3290
rect 17274 3238 17304 3290
rect 17304 3238 17316 3290
rect 17316 3238 17330 3290
rect 17354 3238 17368 3290
rect 17368 3238 17380 3290
rect 17380 3238 17410 3290
rect 17434 3238 17444 3290
rect 17444 3238 17490 3290
rect 17194 3236 17250 3238
rect 17274 3236 17330 3238
rect 17354 3236 17410 3238
rect 17434 3236 17490 3238
rect 17194 2202 17250 2204
rect 17274 2202 17330 2204
rect 17354 2202 17410 2204
rect 17434 2202 17490 2204
rect 17194 2150 17240 2202
rect 17240 2150 17250 2202
rect 17274 2150 17304 2202
rect 17304 2150 17316 2202
rect 17316 2150 17330 2202
rect 17354 2150 17368 2202
rect 17368 2150 17380 2202
rect 17380 2150 17410 2202
rect 17434 2150 17444 2202
rect 17444 2150 17490 2202
rect 17194 2148 17250 2150
rect 17274 2148 17330 2150
rect 17354 2148 17410 2150
rect 17434 2148 17490 2150
rect 20552 7098 20608 7100
rect 20632 7098 20688 7100
rect 20712 7098 20768 7100
rect 20792 7098 20848 7100
rect 20552 7046 20598 7098
rect 20598 7046 20608 7098
rect 20632 7046 20662 7098
rect 20662 7046 20674 7098
rect 20674 7046 20688 7098
rect 20712 7046 20726 7098
rect 20726 7046 20738 7098
rect 20738 7046 20768 7098
rect 20792 7046 20802 7098
rect 20802 7046 20848 7098
rect 20552 7044 20608 7046
rect 20632 7044 20688 7046
rect 20712 7044 20768 7046
rect 20792 7044 20848 7046
rect 27268 31034 27324 31036
rect 27348 31034 27404 31036
rect 27428 31034 27484 31036
rect 27508 31034 27564 31036
rect 27268 30982 27314 31034
rect 27314 30982 27324 31034
rect 27348 30982 27378 31034
rect 27378 30982 27390 31034
rect 27390 30982 27404 31034
rect 27428 30982 27442 31034
rect 27442 30982 27454 31034
rect 27454 30982 27484 31034
rect 27508 30982 27518 31034
rect 27518 30982 27564 31034
rect 27268 30980 27324 30982
rect 27348 30980 27404 30982
rect 27428 30980 27484 30982
rect 27508 30980 27564 30982
rect 27268 29946 27324 29948
rect 27348 29946 27404 29948
rect 27428 29946 27484 29948
rect 27508 29946 27564 29948
rect 27268 29894 27314 29946
rect 27314 29894 27324 29946
rect 27348 29894 27378 29946
rect 27378 29894 27390 29946
rect 27390 29894 27404 29946
rect 27428 29894 27442 29946
rect 27442 29894 27454 29946
rect 27454 29894 27484 29946
rect 27508 29894 27518 29946
rect 27518 29894 27564 29946
rect 27268 29892 27324 29894
rect 27348 29892 27404 29894
rect 27428 29892 27484 29894
rect 27508 29892 27564 29894
rect 25226 29688 25282 29744
rect 25686 29552 25742 29608
rect 24950 27648 25006 27704
rect 23910 23962 23966 23964
rect 23990 23962 24046 23964
rect 24070 23962 24126 23964
rect 24150 23962 24206 23964
rect 23910 23910 23956 23962
rect 23956 23910 23966 23962
rect 23990 23910 24020 23962
rect 24020 23910 24032 23962
rect 24032 23910 24046 23962
rect 24070 23910 24084 23962
rect 24084 23910 24096 23962
rect 24096 23910 24126 23962
rect 24150 23910 24160 23962
rect 24160 23910 24206 23962
rect 23910 23908 23966 23910
rect 23990 23908 24046 23910
rect 24070 23908 24126 23910
rect 24150 23908 24206 23910
rect 23910 22874 23966 22876
rect 23990 22874 24046 22876
rect 24070 22874 24126 22876
rect 24150 22874 24206 22876
rect 23910 22822 23956 22874
rect 23956 22822 23966 22874
rect 23990 22822 24020 22874
rect 24020 22822 24032 22874
rect 24032 22822 24046 22874
rect 24070 22822 24084 22874
rect 24084 22822 24096 22874
rect 24096 22822 24126 22874
rect 24150 22822 24160 22874
rect 24160 22822 24206 22874
rect 23910 22820 23966 22822
rect 23990 22820 24046 22822
rect 24070 22820 24126 22822
rect 24150 22820 24206 22822
rect 23910 21786 23966 21788
rect 23990 21786 24046 21788
rect 24070 21786 24126 21788
rect 24150 21786 24206 21788
rect 23910 21734 23956 21786
rect 23956 21734 23966 21786
rect 23990 21734 24020 21786
rect 24020 21734 24032 21786
rect 24032 21734 24046 21786
rect 24070 21734 24084 21786
rect 24084 21734 24096 21786
rect 24096 21734 24126 21786
rect 24150 21734 24160 21786
rect 24160 21734 24206 21786
rect 23910 21732 23966 21734
rect 23990 21732 24046 21734
rect 24070 21732 24126 21734
rect 24150 21732 24206 21734
rect 23910 20698 23966 20700
rect 23990 20698 24046 20700
rect 24070 20698 24126 20700
rect 24150 20698 24206 20700
rect 23910 20646 23956 20698
rect 23956 20646 23966 20698
rect 23990 20646 24020 20698
rect 24020 20646 24032 20698
rect 24032 20646 24046 20698
rect 24070 20646 24084 20698
rect 24084 20646 24096 20698
rect 24096 20646 24126 20698
rect 24150 20646 24160 20698
rect 24160 20646 24206 20698
rect 23910 20644 23966 20646
rect 23990 20644 24046 20646
rect 24070 20644 24126 20646
rect 24150 20644 24206 20646
rect 23910 19610 23966 19612
rect 23990 19610 24046 19612
rect 24070 19610 24126 19612
rect 24150 19610 24206 19612
rect 23910 19558 23956 19610
rect 23956 19558 23966 19610
rect 23990 19558 24020 19610
rect 24020 19558 24032 19610
rect 24032 19558 24046 19610
rect 24070 19558 24084 19610
rect 24084 19558 24096 19610
rect 24096 19558 24126 19610
rect 24150 19558 24160 19610
rect 24160 19558 24206 19610
rect 23910 19556 23966 19558
rect 23990 19556 24046 19558
rect 24070 19556 24126 19558
rect 24150 19556 24206 19558
rect 27268 28858 27324 28860
rect 27348 28858 27404 28860
rect 27428 28858 27484 28860
rect 27508 28858 27564 28860
rect 27268 28806 27314 28858
rect 27314 28806 27324 28858
rect 27348 28806 27378 28858
rect 27378 28806 27390 28858
rect 27390 28806 27404 28858
rect 27428 28806 27442 28858
rect 27442 28806 27454 28858
rect 27454 28806 27484 28858
rect 27508 28806 27518 28858
rect 27518 28806 27564 28858
rect 27268 28804 27324 28806
rect 27348 28804 27404 28806
rect 27428 28804 27484 28806
rect 27508 28804 27564 28806
rect 27268 27770 27324 27772
rect 27348 27770 27404 27772
rect 27428 27770 27484 27772
rect 27508 27770 27564 27772
rect 27268 27718 27314 27770
rect 27314 27718 27324 27770
rect 27348 27718 27378 27770
rect 27378 27718 27390 27770
rect 27390 27718 27404 27770
rect 27428 27718 27442 27770
rect 27442 27718 27454 27770
rect 27454 27718 27484 27770
rect 27508 27718 27518 27770
rect 27518 27718 27564 27770
rect 27268 27716 27324 27718
rect 27348 27716 27404 27718
rect 27428 27716 27484 27718
rect 27508 27716 27564 27718
rect 27268 26682 27324 26684
rect 27348 26682 27404 26684
rect 27428 26682 27484 26684
rect 27508 26682 27564 26684
rect 27268 26630 27314 26682
rect 27314 26630 27324 26682
rect 27348 26630 27378 26682
rect 27378 26630 27390 26682
rect 27390 26630 27404 26682
rect 27428 26630 27442 26682
rect 27442 26630 27454 26682
rect 27454 26630 27484 26682
rect 27508 26630 27518 26682
rect 27518 26630 27564 26682
rect 27268 26628 27324 26630
rect 27348 26628 27404 26630
rect 27428 26628 27484 26630
rect 27508 26628 27564 26630
rect 27268 25594 27324 25596
rect 27348 25594 27404 25596
rect 27428 25594 27484 25596
rect 27508 25594 27564 25596
rect 27268 25542 27314 25594
rect 27314 25542 27324 25594
rect 27348 25542 27378 25594
rect 27378 25542 27390 25594
rect 27390 25542 27404 25594
rect 27428 25542 27442 25594
rect 27442 25542 27454 25594
rect 27454 25542 27484 25594
rect 27508 25542 27518 25594
rect 27518 25542 27564 25594
rect 27268 25540 27324 25542
rect 27348 25540 27404 25542
rect 27428 25540 27484 25542
rect 27508 25540 27564 25542
rect 27268 24506 27324 24508
rect 27348 24506 27404 24508
rect 27428 24506 27484 24508
rect 27508 24506 27564 24508
rect 27268 24454 27314 24506
rect 27314 24454 27324 24506
rect 27348 24454 27378 24506
rect 27378 24454 27390 24506
rect 27390 24454 27404 24506
rect 27428 24454 27442 24506
rect 27442 24454 27454 24506
rect 27454 24454 27484 24506
rect 27508 24454 27518 24506
rect 27518 24454 27564 24506
rect 27268 24452 27324 24454
rect 27348 24452 27404 24454
rect 27428 24452 27484 24454
rect 27508 24452 27564 24454
rect 27268 23418 27324 23420
rect 27348 23418 27404 23420
rect 27428 23418 27484 23420
rect 27508 23418 27564 23420
rect 27268 23366 27314 23418
rect 27314 23366 27324 23418
rect 27348 23366 27378 23418
rect 27378 23366 27390 23418
rect 27390 23366 27404 23418
rect 27428 23366 27442 23418
rect 27442 23366 27454 23418
rect 27454 23366 27484 23418
rect 27508 23366 27518 23418
rect 27518 23366 27564 23418
rect 27268 23364 27324 23366
rect 27348 23364 27404 23366
rect 27428 23364 27484 23366
rect 27508 23364 27564 23366
rect 27268 22330 27324 22332
rect 27348 22330 27404 22332
rect 27428 22330 27484 22332
rect 27508 22330 27564 22332
rect 27268 22278 27314 22330
rect 27314 22278 27324 22330
rect 27348 22278 27378 22330
rect 27378 22278 27390 22330
rect 27390 22278 27404 22330
rect 27428 22278 27442 22330
rect 27442 22278 27454 22330
rect 27454 22278 27484 22330
rect 27508 22278 27518 22330
rect 27518 22278 27564 22330
rect 27268 22276 27324 22278
rect 27348 22276 27404 22278
rect 27428 22276 27484 22278
rect 27508 22276 27564 22278
rect 27268 21242 27324 21244
rect 27348 21242 27404 21244
rect 27428 21242 27484 21244
rect 27508 21242 27564 21244
rect 27268 21190 27314 21242
rect 27314 21190 27324 21242
rect 27348 21190 27378 21242
rect 27378 21190 27390 21242
rect 27390 21190 27404 21242
rect 27428 21190 27442 21242
rect 27442 21190 27454 21242
rect 27454 21190 27484 21242
rect 27508 21190 27518 21242
rect 27518 21190 27564 21242
rect 27268 21188 27324 21190
rect 27348 21188 27404 21190
rect 27428 21188 27484 21190
rect 27508 21188 27564 21190
rect 23910 18522 23966 18524
rect 23990 18522 24046 18524
rect 24070 18522 24126 18524
rect 24150 18522 24206 18524
rect 23910 18470 23956 18522
rect 23956 18470 23966 18522
rect 23990 18470 24020 18522
rect 24020 18470 24032 18522
rect 24032 18470 24046 18522
rect 24070 18470 24084 18522
rect 24084 18470 24096 18522
rect 24096 18470 24126 18522
rect 24150 18470 24160 18522
rect 24160 18470 24206 18522
rect 23910 18468 23966 18470
rect 23990 18468 24046 18470
rect 24070 18468 24126 18470
rect 24150 18468 24206 18470
rect 23910 17434 23966 17436
rect 23990 17434 24046 17436
rect 24070 17434 24126 17436
rect 24150 17434 24206 17436
rect 23910 17382 23956 17434
rect 23956 17382 23966 17434
rect 23990 17382 24020 17434
rect 24020 17382 24032 17434
rect 24032 17382 24046 17434
rect 24070 17382 24084 17434
rect 24084 17382 24096 17434
rect 24096 17382 24126 17434
rect 24150 17382 24160 17434
rect 24160 17382 24206 17434
rect 23910 17380 23966 17382
rect 23990 17380 24046 17382
rect 24070 17380 24126 17382
rect 24150 17380 24206 17382
rect 23938 17212 23940 17232
rect 23940 17212 23992 17232
rect 23992 17212 23994 17232
rect 23938 17176 23994 17212
rect 24214 16940 24216 16960
rect 24216 16940 24268 16960
rect 24268 16940 24270 16960
rect 24214 16904 24270 16940
rect 24674 16904 24730 16960
rect 24950 17176 25006 17232
rect 23910 16346 23966 16348
rect 23990 16346 24046 16348
rect 24070 16346 24126 16348
rect 24150 16346 24206 16348
rect 23910 16294 23956 16346
rect 23956 16294 23966 16346
rect 23990 16294 24020 16346
rect 24020 16294 24032 16346
rect 24032 16294 24046 16346
rect 24070 16294 24084 16346
rect 24084 16294 24096 16346
rect 24096 16294 24126 16346
rect 24150 16294 24160 16346
rect 24160 16294 24206 16346
rect 23910 16292 23966 16294
rect 23990 16292 24046 16294
rect 24070 16292 24126 16294
rect 24150 16292 24206 16294
rect 27268 20154 27324 20156
rect 27348 20154 27404 20156
rect 27428 20154 27484 20156
rect 27508 20154 27564 20156
rect 27268 20102 27314 20154
rect 27314 20102 27324 20154
rect 27348 20102 27378 20154
rect 27378 20102 27390 20154
rect 27390 20102 27404 20154
rect 27428 20102 27442 20154
rect 27442 20102 27454 20154
rect 27454 20102 27484 20154
rect 27508 20102 27518 20154
rect 27518 20102 27564 20154
rect 27268 20100 27324 20102
rect 27348 20100 27404 20102
rect 27428 20100 27484 20102
rect 27508 20100 27564 20102
rect 27268 19066 27324 19068
rect 27348 19066 27404 19068
rect 27428 19066 27484 19068
rect 27508 19066 27564 19068
rect 27268 19014 27314 19066
rect 27314 19014 27324 19066
rect 27348 19014 27378 19066
rect 27378 19014 27390 19066
rect 27390 19014 27404 19066
rect 27428 19014 27442 19066
rect 27442 19014 27454 19066
rect 27454 19014 27484 19066
rect 27508 19014 27518 19066
rect 27518 19014 27564 19066
rect 27268 19012 27324 19014
rect 27348 19012 27404 19014
rect 27428 19012 27484 19014
rect 27508 19012 27564 19014
rect 27268 17978 27324 17980
rect 27348 17978 27404 17980
rect 27428 17978 27484 17980
rect 27508 17978 27564 17980
rect 27268 17926 27314 17978
rect 27314 17926 27324 17978
rect 27348 17926 27378 17978
rect 27378 17926 27390 17978
rect 27390 17926 27404 17978
rect 27428 17926 27442 17978
rect 27442 17926 27454 17978
rect 27454 17926 27484 17978
rect 27508 17926 27518 17978
rect 27518 17926 27564 17978
rect 27268 17924 27324 17926
rect 27348 17924 27404 17926
rect 27428 17924 27484 17926
rect 27508 17924 27564 17926
rect 27268 16890 27324 16892
rect 27348 16890 27404 16892
rect 27428 16890 27484 16892
rect 27508 16890 27564 16892
rect 27268 16838 27314 16890
rect 27314 16838 27324 16890
rect 27348 16838 27378 16890
rect 27378 16838 27390 16890
rect 27390 16838 27404 16890
rect 27428 16838 27442 16890
rect 27442 16838 27454 16890
rect 27454 16838 27484 16890
rect 27508 16838 27518 16890
rect 27518 16838 27564 16890
rect 27268 16836 27324 16838
rect 27348 16836 27404 16838
rect 27428 16836 27484 16838
rect 27508 16836 27564 16838
rect 23910 15258 23966 15260
rect 23990 15258 24046 15260
rect 24070 15258 24126 15260
rect 24150 15258 24206 15260
rect 23910 15206 23956 15258
rect 23956 15206 23966 15258
rect 23990 15206 24020 15258
rect 24020 15206 24032 15258
rect 24032 15206 24046 15258
rect 24070 15206 24084 15258
rect 24084 15206 24096 15258
rect 24096 15206 24126 15258
rect 24150 15206 24160 15258
rect 24160 15206 24206 15258
rect 23910 15204 23966 15206
rect 23990 15204 24046 15206
rect 24070 15204 24126 15206
rect 24150 15204 24206 15206
rect 27268 15802 27324 15804
rect 27348 15802 27404 15804
rect 27428 15802 27484 15804
rect 27508 15802 27564 15804
rect 27268 15750 27314 15802
rect 27314 15750 27324 15802
rect 27348 15750 27378 15802
rect 27378 15750 27390 15802
rect 27390 15750 27404 15802
rect 27428 15750 27442 15802
rect 27442 15750 27454 15802
rect 27454 15750 27484 15802
rect 27508 15750 27518 15802
rect 27518 15750 27564 15802
rect 27268 15748 27324 15750
rect 27348 15748 27404 15750
rect 27428 15748 27484 15750
rect 27508 15748 27564 15750
rect 23910 14170 23966 14172
rect 23990 14170 24046 14172
rect 24070 14170 24126 14172
rect 24150 14170 24206 14172
rect 23910 14118 23956 14170
rect 23956 14118 23966 14170
rect 23990 14118 24020 14170
rect 24020 14118 24032 14170
rect 24032 14118 24046 14170
rect 24070 14118 24084 14170
rect 24084 14118 24096 14170
rect 24096 14118 24126 14170
rect 24150 14118 24160 14170
rect 24160 14118 24206 14170
rect 23910 14116 23966 14118
rect 23990 14116 24046 14118
rect 24070 14116 24126 14118
rect 24150 14116 24206 14118
rect 23910 13082 23966 13084
rect 23990 13082 24046 13084
rect 24070 13082 24126 13084
rect 24150 13082 24206 13084
rect 23910 13030 23956 13082
rect 23956 13030 23966 13082
rect 23990 13030 24020 13082
rect 24020 13030 24032 13082
rect 24032 13030 24046 13082
rect 24070 13030 24084 13082
rect 24084 13030 24096 13082
rect 24096 13030 24126 13082
rect 24150 13030 24160 13082
rect 24160 13030 24206 13082
rect 23910 13028 23966 13030
rect 23990 13028 24046 13030
rect 24070 13028 24126 13030
rect 24150 13028 24206 13030
rect 23910 11994 23966 11996
rect 23990 11994 24046 11996
rect 24070 11994 24126 11996
rect 24150 11994 24206 11996
rect 23910 11942 23956 11994
rect 23956 11942 23966 11994
rect 23990 11942 24020 11994
rect 24020 11942 24032 11994
rect 24032 11942 24046 11994
rect 24070 11942 24084 11994
rect 24084 11942 24096 11994
rect 24096 11942 24126 11994
rect 24150 11942 24160 11994
rect 24160 11942 24206 11994
rect 23910 11940 23966 11942
rect 23990 11940 24046 11942
rect 24070 11940 24126 11942
rect 24150 11940 24206 11942
rect 23910 10906 23966 10908
rect 23990 10906 24046 10908
rect 24070 10906 24126 10908
rect 24150 10906 24206 10908
rect 23910 10854 23956 10906
rect 23956 10854 23966 10906
rect 23990 10854 24020 10906
rect 24020 10854 24032 10906
rect 24032 10854 24046 10906
rect 24070 10854 24084 10906
rect 24084 10854 24096 10906
rect 24096 10854 24126 10906
rect 24150 10854 24160 10906
rect 24160 10854 24206 10906
rect 23910 10852 23966 10854
rect 23990 10852 24046 10854
rect 24070 10852 24126 10854
rect 24150 10852 24206 10854
rect 23910 9818 23966 9820
rect 23990 9818 24046 9820
rect 24070 9818 24126 9820
rect 24150 9818 24206 9820
rect 23910 9766 23956 9818
rect 23956 9766 23966 9818
rect 23990 9766 24020 9818
rect 24020 9766 24032 9818
rect 24032 9766 24046 9818
rect 24070 9766 24084 9818
rect 24084 9766 24096 9818
rect 24096 9766 24126 9818
rect 24150 9766 24160 9818
rect 24160 9766 24206 9818
rect 23910 9764 23966 9766
rect 23990 9764 24046 9766
rect 24070 9764 24126 9766
rect 24150 9764 24206 9766
rect 23910 8730 23966 8732
rect 23990 8730 24046 8732
rect 24070 8730 24126 8732
rect 24150 8730 24206 8732
rect 23910 8678 23956 8730
rect 23956 8678 23966 8730
rect 23990 8678 24020 8730
rect 24020 8678 24032 8730
rect 24032 8678 24046 8730
rect 24070 8678 24084 8730
rect 24084 8678 24096 8730
rect 24096 8678 24126 8730
rect 24150 8678 24160 8730
rect 24160 8678 24206 8730
rect 23910 8676 23966 8678
rect 23990 8676 24046 8678
rect 24070 8676 24126 8678
rect 24150 8676 24206 8678
rect 17194 1114 17250 1116
rect 17274 1114 17330 1116
rect 17354 1114 17410 1116
rect 17434 1114 17490 1116
rect 17194 1062 17240 1114
rect 17240 1062 17250 1114
rect 17274 1062 17304 1114
rect 17304 1062 17316 1114
rect 17316 1062 17330 1114
rect 17354 1062 17368 1114
rect 17368 1062 17380 1114
rect 17380 1062 17410 1114
rect 17434 1062 17444 1114
rect 17444 1062 17490 1114
rect 17194 1060 17250 1062
rect 17274 1060 17330 1062
rect 17354 1060 17410 1062
rect 17434 1060 17490 1062
rect 20552 6010 20608 6012
rect 20632 6010 20688 6012
rect 20712 6010 20768 6012
rect 20792 6010 20848 6012
rect 20552 5958 20598 6010
rect 20598 5958 20608 6010
rect 20632 5958 20662 6010
rect 20662 5958 20674 6010
rect 20674 5958 20688 6010
rect 20712 5958 20726 6010
rect 20726 5958 20738 6010
rect 20738 5958 20768 6010
rect 20792 5958 20802 6010
rect 20802 5958 20848 6010
rect 20552 5956 20608 5958
rect 20632 5956 20688 5958
rect 20712 5956 20768 5958
rect 20792 5956 20848 5958
rect 23910 7642 23966 7644
rect 23990 7642 24046 7644
rect 24070 7642 24126 7644
rect 24150 7642 24206 7644
rect 23910 7590 23956 7642
rect 23956 7590 23966 7642
rect 23990 7590 24020 7642
rect 24020 7590 24032 7642
rect 24032 7590 24046 7642
rect 24070 7590 24084 7642
rect 24084 7590 24096 7642
rect 24096 7590 24126 7642
rect 24150 7590 24160 7642
rect 24160 7590 24206 7642
rect 23910 7588 23966 7590
rect 23990 7588 24046 7590
rect 24070 7588 24126 7590
rect 24150 7588 24206 7590
rect 27268 14714 27324 14716
rect 27348 14714 27404 14716
rect 27428 14714 27484 14716
rect 27508 14714 27564 14716
rect 27268 14662 27314 14714
rect 27314 14662 27324 14714
rect 27348 14662 27378 14714
rect 27378 14662 27390 14714
rect 27390 14662 27404 14714
rect 27428 14662 27442 14714
rect 27442 14662 27454 14714
rect 27454 14662 27484 14714
rect 27508 14662 27518 14714
rect 27518 14662 27564 14714
rect 27268 14660 27324 14662
rect 27348 14660 27404 14662
rect 27428 14660 27484 14662
rect 27508 14660 27564 14662
rect 27268 13626 27324 13628
rect 27348 13626 27404 13628
rect 27428 13626 27484 13628
rect 27508 13626 27564 13628
rect 27268 13574 27314 13626
rect 27314 13574 27324 13626
rect 27348 13574 27378 13626
rect 27378 13574 27390 13626
rect 27390 13574 27404 13626
rect 27428 13574 27442 13626
rect 27442 13574 27454 13626
rect 27454 13574 27484 13626
rect 27508 13574 27518 13626
rect 27518 13574 27564 13626
rect 27268 13572 27324 13574
rect 27348 13572 27404 13574
rect 27428 13572 27484 13574
rect 27508 13572 27564 13574
rect 27268 12538 27324 12540
rect 27348 12538 27404 12540
rect 27428 12538 27484 12540
rect 27508 12538 27564 12540
rect 27268 12486 27314 12538
rect 27314 12486 27324 12538
rect 27348 12486 27378 12538
rect 27378 12486 27390 12538
rect 27390 12486 27404 12538
rect 27428 12486 27442 12538
rect 27442 12486 27454 12538
rect 27454 12486 27484 12538
rect 27508 12486 27518 12538
rect 27518 12486 27564 12538
rect 27268 12484 27324 12486
rect 27348 12484 27404 12486
rect 27428 12484 27484 12486
rect 27508 12484 27564 12486
rect 27268 11450 27324 11452
rect 27348 11450 27404 11452
rect 27428 11450 27484 11452
rect 27508 11450 27564 11452
rect 27268 11398 27314 11450
rect 27314 11398 27324 11450
rect 27348 11398 27378 11450
rect 27378 11398 27390 11450
rect 27390 11398 27404 11450
rect 27428 11398 27442 11450
rect 27442 11398 27454 11450
rect 27454 11398 27484 11450
rect 27508 11398 27518 11450
rect 27518 11398 27564 11450
rect 27268 11396 27324 11398
rect 27348 11396 27404 11398
rect 27428 11396 27484 11398
rect 27508 11396 27564 11398
rect 27268 10362 27324 10364
rect 27348 10362 27404 10364
rect 27428 10362 27484 10364
rect 27508 10362 27564 10364
rect 27268 10310 27314 10362
rect 27314 10310 27324 10362
rect 27348 10310 27378 10362
rect 27378 10310 27390 10362
rect 27390 10310 27404 10362
rect 27428 10310 27442 10362
rect 27442 10310 27454 10362
rect 27454 10310 27484 10362
rect 27508 10310 27518 10362
rect 27518 10310 27564 10362
rect 27268 10308 27324 10310
rect 27348 10308 27404 10310
rect 27428 10308 27484 10310
rect 27508 10308 27564 10310
rect 23910 6554 23966 6556
rect 23990 6554 24046 6556
rect 24070 6554 24126 6556
rect 24150 6554 24206 6556
rect 23910 6502 23956 6554
rect 23956 6502 23966 6554
rect 23990 6502 24020 6554
rect 24020 6502 24032 6554
rect 24032 6502 24046 6554
rect 24070 6502 24084 6554
rect 24084 6502 24096 6554
rect 24096 6502 24126 6554
rect 24150 6502 24160 6554
rect 24160 6502 24206 6554
rect 23910 6500 23966 6502
rect 23990 6500 24046 6502
rect 24070 6500 24126 6502
rect 24150 6500 24206 6502
rect 20552 4922 20608 4924
rect 20632 4922 20688 4924
rect 20712 4922 20768 4924
rect 20792 4922 20848 4924
rect 20552 4870 20598 4922
rect 20598 4870 20608 4922
rect 20632 4870 20662 4922
rect 20662 4870 20674 4922
rect 20674 4870 20688 4922
rect 20712 4870 20726 4922
rect 20726 4870 20738 4922
rect 20738 4870 20768 4922
rect 20792 4870 20802 4922
rect 20802 4870 20848 4922
rect 20552 4868 20608 4870
rect 20632 4868 20688 4870
rect 20712 4868 20768 4870
rect 20792 4868 20848 4870
rect 20552 3834 20608 3836
rect 20632 3834 20688 3836
rect 20712 3834 20768 3836
rect 20792 3834 20848 3836
rect 20552 3782 20598 3834
rect 20598 3782 20608 3834
rect 20632 3782 20662 3834
rect 20662 3782 20674 3834
rect 20674 3782 20688 3834
rect 20712 3782 20726 3834
rect 20726 3782 20738 3834
rect 20738 3782 20768 3834
rect 20792 3782 20802 3834
rect 20802 3782 20848 3834
rect 20552 3780 20608 3782
rect 20632 3780 20688 3782
rect 20712 3780 20768 3782
rect 20792 3780 20848 3782
rect 20552 2746 20608 2748
rect 20632 2746 20688 2748
rect 20712 2746 20768 2748
rect 20792 2746 20848 2748
rect 20552 2694 20598 2746
rect 20598 2694 20608 2746
rect 20632 2694 20662 2746
rect 20662 2694 20674 2746
rect 20674 2694 20688 2746
rect 20712 2694 20726 2746
rect 20726 2694 20738 2746
rect 20738 2694 20768 2746
rect 20792 2694 20802 2746
rect 20802 2694 20848 2746
rect 20552 2692 20608 2694
rect 20632 2692 20688 2694
rect 20712 2692 20768 2694
rect 20792 2692 20848 2694
rect 20552 1658 20608 1660
rect 20632 1658 20688 1660
rect 20712 1658 20768 1660
rect 20792 1658 20848 1660
rect 20552 1606 20598 1658
rect 20598 1606 20608 1658
rect 20632 1606 20662 1658
rect 20662 1606 20674 1658
rect 20674 1606 20688 1658
rect 20712 1606 20726 1658
rect 20726 1606 20738 1658
rect 20738 1606 20768 1658
rect 20792 1606 20802 1658
rect 20802 1606 20848 1658
rect 20552 1604 20608 1606
rect 20632 1604 20688 1606
rect 20712 1604 20768 1606
rect 20792 1604 20848 1606
rect 20552 570 20608 572
rect 20632 570 20688 572
rect 20712 570 20768 572
rect 20792 570 20848 572
rect 20552 518 20598 570
rect 20598 518 20608 570
rect 20632 518 20662 570
rect 20662 518 20674 570
rect 20674 518 20688 570
rect 20712 518 20726 570
rect 20726 518 20738 570
rect 20738 518 20768 570
rect 20792 518 20802 570
rect 20802 518 20848 570
rect 20552 516 20608 518
rect 20632 516 20688 518
rect 20712 516 20768 518
rect 20792 516 20848 518
rect 23910 5466 23966 5468
rect 23990 5466 24046 5468
rect 24070 5466 24126 5468
rect 24150 5466 24206 5468
rect 23910 5414 23956 5466
rect 23956 5414 23966 5466
rect 23990 5414 24020 5466
rect 24020 5414 24032 5466
rect 24032 5414 24046 5466
rect 24070 5414 24084 5466
rect 24084 5414 24096 5466
rect 24096 5414 24126 5466
rect 24150 5414 24160 5466
rect 24160 5414 24206 5466
rect 23910 5412 23966 5414
rect 23990 5412 24046 5414
rect 24070 5412 24126 5414
rect 24150 5412 24206 5414
rect 23910 4378 23966 4380
rect 23990 4378 24046 4380
rect 24070 4378 24126 4380
rect 24150 4378 24206 4380
rect 23910 4326 23956 4378
rect 23956 4326 23966 4378
rect 23990 4326 24020 4378
rect 24020 4326 24032 4378
rect 24032 4326 24046 4378
rect 24070 4326 24084 4378
rect 24084 4326 24096 4378
rect 24096 4326 24126 4378
rect 24150 4326 24160 4378
rect 24160 4326 24206 4378
rect 23910 4324 23966 4326
rect 23990 4324 24046 4326
rect 24070 4324 24126 4326
rect 24150 4324 24206 4326
rect 23910 3290 23966 3292
rect 23990 3290 24046 3292
rect 24070 3290 24126 3292
rect 24150 3290 24206 3292
rect 23910 3238 23956 3290
rect 23956 3238 23966 3290
rect 23990 3238 24020 3290
rect 24020 3238 24032 3290
rect 24032 3238 24046 3290
rect 24070 3238 24084 3290
rect 24084 3238 24096 3290
rect 24096 3238 24126 3290
rect 24150 3238 24160 3290
rect 24160 3238 24206 3290
rect 23910 3236 23966 3238
rect 23990 3236 24046 3238
rect 24070 3236 24126 3238
rect 24150 3236 24206 3238
rect 27268 9274 27324 9276
rect 27348 9274 27404 9276
rect 27428 9274 27484 9276
rect 27508 9274 27564 9276
rect 27268 9222 27314 9274
rect 27314 9222 27324 9274
rect 27348 9222 27378 9274
rect 27378 9222 27390 9274
rect 27390 9222 27404 9274
rect 27428 9222 27442 9274
rect 27442 9222 27454 9274
rect 27454 9222 27484 9274
rect 27508 9222 27518 9274
rect 27518 9222 27564 9274
rect 27268 9220 27324 9222
rect 27348 9220 27404 9222
rect 27428 9220 27484 9222
rect 27508 9220 27564 9222
rect 27268 8186 27324 8188
rect 27348 8186 27404 8188
rect 27428 8186 27484 8188
rect 27508 8186 27564 8188
rect 27268 8134 27314 8186
rect 27314 8134 27324 8186
rect 27348 8134 27378 8186
rect 27378 8134 27390 8186
rect 27390 8134 27404 8186
rect 27428 8134 27442 8186
rect 27442 8134 27454 8186
rect 27454 8134 27484 8186
rect 27508 8134 27518 8186
rect 27518 8134 27564 8186
rect 27268 8132 27324 8134
rect 27348 8132 27404 8134
rect 27428 8132 27484 8134
rect 27508 8132 27564 8134
rect 27268 7098 27324 7100
rect 27348 7098 27404 7100
rect 27428 7098 27484 7100
rect 27508 7098 27564 7100
rect 27268 7046 27314 7098
rect 27314 7046 27324 7098
rect 27348 7046 27378 7098
rect 27378 7046 27390 7098
rect 27390 7046 27404 7098
rect 27428 7046 27442 7098
rect 27442 7046 27454 7098
rect 27454 7046 27484 7098
rect 27508 7046 27518 7098
rect 27518 7046 27564 7098
rect 27268 7044 27324 7046
rect 27348 7044 27404 7046
rect 27428 7044 27484 7046
rect 27508 7044 27564 7046
rect 27268 6010 27324 6012
rect 27348 6010 27404 6012
rect 27428 6010 27484 6012
rect 27508 6010 27564 6012
rect 27268 5958 27314 6010
rect 27314 5958 27324 6010
rect 27348 5958 27378 6010
rect 27378 5958 27390 6010
rect 27390 5958 27404 6010
rect 27428 5958 27442 6010
rect 27442 5958 27454 6010
rect 27454 5958 27484 6010
rect 27508 5958 27518 6010
rect 27518 5958 27564 6010
rect 27268 5956 27324 5958
rect 27348 5956 27404 5958
rect 27428 5956 27484 5958
rect 27508 5956 27564 5958
rect 27268 4922 27324 4924
rect 27348 4922 27404 4924
rect 27428 4922 27484 4924
rect 27508 4922 27564 4924
rect 27268 4870 27314 4922
rect 27314 4870 27324 4922
rect 27348 4870 27378 4922
rect 27378 4870 27390 4922
rect 27390 4870 27404 4922
rect 27428 4870 27442 4922
rect 27442 4870 27454 4922
rect 27454 4870 27484 4922
rect 27508 4870 27518 4922
rect 27518 4870 27564 4922
rect 27268 4868 27324 4870
rect 27348 4868 27404 4870
rect 27428 4868 27484 4870
rect 27508 4868 27564 4870
rect 27268 3834 27324 3836
rect 27348 3834 27404 3836
rect 27428 3834 27484 3836
rect 27508 3834 27564 3836
rect 27268 3782 27314 3834
rect 27314 3782 27324 3834
rect 27348 3782 27378 3834
rect 27378 3782 27390 3834
rect 27390 3782 27404 3834
rect 27428 3782 27442 3834
rect 27442 3782 27454 3834
rect 27454 3782 27484 3834
rect 27508 3782 27518 3834
rect 27518 3782 27564 3834
rect 27268 3780 27324 3782
rect 27348 3780 27404 3782
rect 27428 3780 27484 3782
rect 27508 3780 27564 3782
rect 23910 2202 23966 2204
rect 23990 2202 24046 2204
rect 24070 2202 24126 2204
rect 24150 2202 24206 2204
rect 23910 2150 23956 2202
rect 23956 2150 23966 2202
rect 23990 2150 24020 2202
rect 24020 2150 24032 2202
rect 24032 2150 24046 2202
rect 24070 2150 24084 2202
rect 24084 2150 24096 2202
rect 24096 2150 24126 2202
rect 24150 2150 24160 2202
rect 24160 2150 24206 2202
rect 23910 2148 23966 2150
rect 23990 2148 24046 2150
rect 24070 2148 24126 2150
rect 24150 2148 24206 2150
rect 23910 1114 23966 1116
rect 23990 1114 24046 1116
rect 24070 1114 24126 1116
rect 24150 1114 24206 1116
rect 23910 1062 23956 1114
rect 23956 1062 23966 1114
rect 23990 1062 24020 1114
rect 24020 1062 24032 1114
rect 24032 1062 24046 1114
rect 24070 1062 24084 1114
rect 24084 1062 24096 1114
rect 24096 1062 24126 1114
rect 24150 1062 24160 1114
rect 24160 1062 24206 1114
rect 23910 1060 23966 1062
rect 23990 1060 24046 1062
rect 24070 1060 24126 1062
rect 24150 1060 24206 1062
rect 27268 2746 27324 2748
rect 27348 2746 27404 2748
rect 27428 2746 27484 2748
rect 27508 2746 27564 2748
rect 27268 2694 27314 2746
rect 27314 2694 27324 2746
rect 27348 2694 27378 2746
rect 27378 2694 27390 2746
rect 27390 2694 27404 2746
rect 27428 2694 27442 2746
rect 27442 2694 27454 2746
rect 27454 2694 27484 2746
rect 27508 2694 27518 2746
rect 27518 2694 27564 2746
rect 27268 2692 27324 2694
rect 27348 2692 27404 2694
rect 27428 2692 27484 2694
rect 27508 2692 27564 2694
rect 27268 1658 27324 1660
rect 27348 1658 27404 1660
rect 27428 1658 27484 1660
rect 27508 1658 27564 1660
rect 27268 1606 27314 1658
rect 27314 1606 27324 1658
rect 27348 1606 27378 1658
rect 27378 1606 27390 1658
rect 27390 1606 27404 1658
rect 27428 1606 27442 1658
rect 27442 1606 27454 1658
rect 27454 1606 27484 1658
rect 27508 1606 27518 1658
rect 27518 1606 27564 1658
rect 27268 1604 27324 1606
rect 27348 1604 27404 1606
rect 27428 1604 27484 1606
rect 27508 1604 27564 1606
rect 27268 570 27324 572
rect 27348 570 27404 572
rect 27428 570 27484 572
rect 27508 570 27564 572
rect 27268 518 27314 570
rect 27314 518 27324 570
rect 27348 518 27378 570
rect 27378 518 27390 570
rect 27390 518 27404 570
rect 27428 518 27442 570
rect 27442 518 27454 570
rect 27454 518 27484 570
rect 27508 518 27518 570
rect 27518 518 27564 570
rect 27268 516 27324 518
rect 27348 516 27404 518
rect 27428 516 27484 518
rect 27508 516 27564 518
<< metal3 >>
rect 7110 31040 7426 31041
rect 7110 30976 7116 31040
rect 7180 30976 7196 31040
rect 7260 30976 7276 31040
rect 7340 30976 7356 31040
rect 7420 30976 7426 31040
rect 7110 30975 7426 30976
rect 13826 31040 14142 31041
rect 13826 30976 13832 31040
rect 13896 30976 13912 31040
rect 13976 30976 13992 31040
rect 14056 30976 14072 31040
rect 14136 30976 14142 31040
rect 13826 30975 14142 30976
rect 20542 31040 20858 31041
rect 20542 30976 20548 31040
rect 20612 30976 20628 31040
rect 20692 30976 20708 31040
rect 20772 30976 20788 31040
rect 20852 30976 20858 31040
rect 20542 30975 20858 30976
rect 27258 31040 27574 31041
rect 27258 30976 27264 31040
rect 27328 30976 27344 31040
rect 27408 30976 27424 31040
rect 27488 30976 27504 31040
rect 27568 30976 27574 31040
rect 27258 30975 27574 30976
rect 3752 30496 4068 30497
rect 3752 30432 3758 30496
rect 3822 30432 3838 30496
rect 3902 30432 3918 30496
rect 3982 30432 3998 30496
rect 4062 30432 4068 30496
rect 3752 30431 4068 30432
rect 10468 30496 10784 30497
rect 10468 30432 10474 30496
rect 10538 30432 10554 30496
rect 10618 30432 10634 30496
rect 10698 30432 10714 30496
rect 10778 30432 10784 30496
rect 10468 30431 10784 30432
rect 17184 30496 17500 30497
rect 17184 30432 17190 30496
rect 17254 30432 17270 30496
rect 17334 30432 17350 30496
rect 17414 30432 17430 30496
rect 17494 30432 17500 30496
rect 17184 30431 17500 30432
rect 23900 30496 24216 30497
rect 23900 30432 23906 30496
rect 23970 30432 23986 30496
rect 24050 30432 24066 30496
rect 24130 30432 24146 30496
rect 24210 30432 24216 30496
rect 23900 30431 24216 30432
rect 2037 30428 2103 30429
rect 2037 30424 2084 30428
rect 2148 30426 2154 30428
rect 2037 30368 2042 30424
rect 2037 30364 2084 30368
rect 2148 30366 2194 30426
rect 2148 30364 2154 30366
rect 2037 30363 2103 30364
rect 20805 30154 20871 30157
rect 23841 30154 23907 30157
rect 20805 30152 23907 30154
rect 20805 30096 20810 30152
rect 20866 30096 23846 30152
rect 23902 30096 23907 30152
rect 20805 30094 23907 30096
rect 20805 30091 20871 30094
rect 23841 30091 23907 30094
rect 7110 29952 7426 29953
rect 7110 29888 7116 29952
rect 7180 29888 7196 29952
rect 7260 29888 7276 29952
rect 7340 29888 7356 29952
rect 7420 29888 7426 29952
rect 7110 29887 7426 29888
rect 13826 29952 14142 29953
rect 13826 29888 13832 29952
rect 13896 29888 13912 29952
rect 13976 29888 13992 29952
rect 14056 29888 14072 29952
rect 14136 29888 14142 29952
rect 13826 29887 14142 29888
rect 20542 29952 20858 29953
rect 20542 29888 20548 29952
rect 20612 29888 20628 29952
rect 20692 29888 20708 29952
rect 20772 29888 20788 29952
rect 20852 29888 20858 29952
rect 20542 29887 20858 29888
rect 27258 29952 27574 29953
rect 27258 29888 27264 29952
rect 27328 29888 27344 29952
rect 27408 29888 27424 29952
rect 27488 29888 27504 29952
rect 27568 29888 27574 29952
rect 27258 29887 27574 29888
rect 1853 29748 1919 29749
rect 1853 29744 1900 29748
rect 1964 29746 1970 29748
rect 22829 29746 22895 29749
rect 25221 29746 25287 29749
rect 1853 29688 1858 29744
rect 1853 29684 1900 29688
rect 1964 29686 2010 29746
rect 22829 29744 25287 29746
rect 22829 29688 22834 29744
rect 22890 29688 25226 29744
rect 25282 29688 25287 29744
rect 22829 29686 25287 29688
rect 1964 29684 1970 29686
rect 1853 29683 1919 29684
rect 22829 29683 22895 29686
rect 25221 29683 25287 29686
rect 11973 29610 12039 29613
rect 16573 29610 16639 29613
rect 18965 29610 19031 29613
rect 11973 29608 19031 29610
rect 11973 29552 11978 29608
rect 12034 29552 16578 29608
rect 16634 29552 18970 29608
rect 19026 29552 19031 29608
rect 11973 29550 19031 29552
rect 11973 29547 12039 29550
rect 16573 29547 16639 29550
rect 18965 29547 19031 29550
rect 22921 29610 22987 29613
rect 23841 29610 23907 29613
rect 25681 29610 25747 29613
rect 22921 29608 25747 29610
rect 22921 29552 22926 29608
rect 22982 29552 23846 29608
rect 23902 29552 25686 29608
rect 25742 29552 25747 29608
rect 22921 29550 25747 29552
rect 22921 29547 22987 29550
rect 23841 29547 23907 29550
rect 25681 29547 25747 29550
rect 6453 29474 6519 29477
rect 7741 29474 7807 29477
rect 6453 29472 7807 29474
rect 6453 29416 6458 29472
rect 6514 29416 7746 29472
rect 7802 29416 7807 29472
rect 6453 29414 7807 29416
rect 6453 29411 6519 29414
rect 7741 29411 7807 29414
rect 3752 29408 4068 29409
rect 3752 29344 3758 29408
rect 3822 29344 3838 29408
rect 3902 29344 3918 29408
rect 3982 29344 3998 29408
rect 4062 29344 4068 29408
rect 3752 29343 4068 29344
rect 10468 29408 10784 29409
rect 10468 29344 10474 29408
rect 10538 29344 10554 29408
rect 10618 29344 10634 29408
rect 10698 29344 10714 29408
rect 10778 29344 10784 29408
rect 10468 29343 10784 29344
rect 17184 29408 17500 29409
rect 17184 29344 17190 29408
rect 17254 29344 17270 29408
rect 17334 29344 17350 29408
rect 17414 29344 17430 29408
rect 17494 29344 17500 29408
rect 17184 29343 17500 29344
rect 23900 29408 24216 29409
rect 23900 29344 23906 29408
rect 23970 29344 23986 29408
rect 24050 29344 24066 29408
rect 24130 29344 24146 29408
rect 24210 29344 24216 29408
rect 23900 29343 24216 29344
rect 4153 29066 4219 29069
rect 4613 29066 4679 29069
rect 4153 29064 4679 29066
rect 4153 29008 4158 29064
rect 4214 29008 4618 29064
rect 4674 29008 4679 29064
rect 4153 29006 4679 29008
rect 4153 29003 4219 29006
rect 4613 29003 4679 29006
rect 7110 28864 7426 28865
rect 7110 28800 7116 28864
rect 7180 28800 7196 28864
rect 7260 28800 7276 28864
rect 7340 28800 7356 28864
rect 7420 28800 7426 28864
rect 7110 28799 7426 28800
rect 13826 28864 14142 28865
rect 13826 28800 13832 28864
rect 13896 28800 13912 28864
rect 13976 28800 13992 28864
rect 14056 28800 14072 28864
rect 14136 28800 14142 28864
rect 13826 28799 14142 28800
rect 20542 28864 20858 28865
rect 20542 28800 20548 28864
rect 20612 28800 20628 28864
rect 20692 28800 20708 28864
rect 20772 28800 20788 28864
rect 20852 28800 20858 28864
rect 20542 28799 20858 28800
rect 27258 28864 27574 28865
rect 27258 28800 27264 28864
rect 27328 28800 27344 28864
rect 27408 28800 27424 28864
rect 27488 28800 27504 28864
rect 27568 28800 27574 28864
rect 27258 28799 27574 28800
rect 3752 28320 4068 28321
rect 3752 28256 3758 28320
rect 3822 28256 3838 28320
rect 3902 28256 3918 28320
rect 3982 28256 3998 28320
rect 4062 28256 4068 28320
rect 3752 28255 4068 28256
rect 10468 28320 10784 28321
rect 10468 28256 10474 28320
rect 10538 28256 10554 28320
rect 10618 28256 10634 28320
rect 10698 28256 10714 28320
rect 10778 28256 10784 28320
rect 10468 28255 10784 28256
rect 17184 28320 17500 28321
rect 17184 28256 17190 28320
rect 17254 28256 17270 28320
rect 17334 28256 17350 28320
rect 17414 28256 17430 28320
rect 17494 28256 17500 28320
rect 17184 28255 17500 28256
rect 23900 28320 24216 28321
rect 23900 28256 23906 28320
rect 23970 28256 23986 28320
rect 24050 28256 24066 28320
rect 24130 28256 24146 28320
rect 24210 28256 24216 28320
rect 23900 28255 24216 28256
rect 16665 27842 16731 27845
rect 17217 27842 17283 27845
rect 16665 27840 17283 27842
rect 16665 27784 16670 27840
rect 16726 27784 17222 27840
rect 17278 27784 17283 27840
rect 16665 27782 17283 27784
rect 16665 27779 16731 27782
rect 17217 27779 17283 27782
rect 7110 27776 7426 27777
rect 7110 27712 7116 27776
rect 7180 27712 7196 27776
rect 7260 27712 7276 27776
rect 7340 27712 7356 27776
rect 7420 27712 7426 27776
rect 7110 27711 7426 27712
rect 13826 27776 14142 27777
rect 13826 27712 13832 27776
rect 13896 27712 13912 27776
rect 13976 27712 13992 27776
rect 14056 27712 14072 27776
rect 14136 27712 14142 27776
rect 13826 27711 14142 27712
rect 20542 27776 20858 27777
rect 20542 27712 20548 27776
rect 20612 27712 20628 27776
rect 20692 27712 20708 27776
rect 20772 27712 20788 27776
rect 20852 27712 20858 27776
rect 20542 27711 20858 27712
rect 27258 27776 27574 27777
rect 27258 27712 27264 27776
rect 27328 27712 27344 27776
rect 27408 27712 27424 27776
rect 27488 27712 27504 27776
rect 27568 27712 27574 27776
rect 27258 27711 27574 27712
rect 17217 27706 17283 27709
rect 17585 27706 17651 27709
rect 24945 27708 25011 27709
rect 24894 27706 24900 27708
rect 17217 27704 17651 27706
rect 17217 27648 17222 27704
rect 17278 27648 17590 27704
rect 17646 27648 17651 27704
rect 17217 27646 17651 27648
rect 24854 27646 24900 27706
rect 24964 27704 25011 27708
rect 25006 27648 25011 27704
rect 17217 27643 17283 27646
rect 17585 27643 17651 27646
rect 24894 27644 24900 27646
rect 24964 27644 25011 27648
rect 24945 27643 25011 27644
rect 3752 27232 4068 27233
rect 3752 27168 3758 27232
rect 3822 27168 3838 27232
rect 3902 27168 3918 27232
rect 3982 27168 3998 27232
rect 4062 27168 4068 27232
rect 3752 27167 4068 27168
rect 10468 27232 10784 27233
rect 10468 27168 10474 27232
rect 10538 27168 10554 27232
rect 10618 27168 10634 27232
rect 10698 27168 10714 27232
rect 10778 27168 10784 27232
rect 10468 27167 10784 27168
rect 17184 27232 17500 27233
rect 17184 27168 17190 27232
rect 17254 27168 17270 27232
rect 17334 27168 17350 27232
rect 17414 27168 17430 27232
rect 17494 27168 17500 27232
rect 17184 27167 17500 27168
rect 23900 27232 24216 27233
rect 23900 27168 23906 27232
rect 23970 27168 23986 27232
rect 24050 27168 24066 27232
rect 24130 27168 24146 27232
rect 24210 27168 24216 27232
rect 23900 27167 24216 27168
rect 21265 27026 21331 27029
rect 23473 27026 23539 27029
rect 21265 27024 23539 27026
rect 21265 26968 21270 27024
rect 21326 26968 23478 27024
rect 23534 26968 23539 27024
rect 21265 26966 23539 26968
rect 21265 26963 21331 26966
rect 23473 26963 23539 26966
rect 7110 26688 7426 26689
rect 7110 26624 7116 26688
rect 7180 26624 7196 26688
rect 7260 26624 7276 26688
rect 7340 26624 7356 26688
rect 7420 26624 7426 26688
rect 7110 26623 7426 26624
rect 13826 26688 14142 26689
rect 13826 26624 13832 26688
rect 13896 26624 13912 26688
rect 13976 26624 13992 26688
rect 14056 26624 14072 26688
rect 14136 26624 14142 26688
rect 13826 26623 14142 26624
rect 20542 26688 20858 26689
rect 20542 26624 20548 26688
rect 20612 26624 20628 26688
rect 20692 26624 20708 26688
rect 20772 26624 20788 26688
rect 20852 26624 20858 26688
rect 20542 26623 20858 26624
rect 27258 26688 27574 26689
rect 27258 26624 27264 26688
rect 27328 26624 27344 26688
rect 27408 26624 27424 26688
rect 27488 26624 27504 26688
rect 27568 26624 27574 26688
rect 27258 26623 27574 26624
rect 21541 26618 21607 26621
rect 21817 26618 21883 26621
rect 21541 26616 21883 26618
rect 21541 26560 21546 26616
rect 21602 26560 21822 26616
rect 21878 26560 21883 26616
rect 21541 26558 21883 26560
rect 21541 26555 21607 26558
rect 21817 26555 21883 26558
rect 3752 26144 4068 26145
rect 3752 26080 3758 26144
rect 3822 26080 3838 26144
rect 3902 26080 3918 26144
rect 3982 26080 3998 26144
rect 4062 26080 4068 26144
rect 3752 26079 4068 26080
rect 10468 26144 10784 26145
rect 10468 26080 10474 26144
rect 10538 26080 10554 26144
rect 10618 26080 10634 26144
rect 10698 26080 10714 26144
rect 10778 26080 10784 26144
rect 10468 26079 10784 26080
rect 17184 26144 17500 26145
rect 17184 26080 17190 26144
rect 17254 26080 17270 26144
rect 17334 26080 17350 26144
rect 17414 26080 17430 26144
rect 17494 26080 17500 26144
rect 17184 26079 17500 26080
rect 23900 26144 24216 26145
rect 23900 26080 23906 26144
rect 23970 26080 23986 26144
rect 24050 26080 24066 26144
rect 24130 26080 24146 26144
rect 24210 26080 24216 26144
rect 23900 26079 24216 26080
rect 7110 25600 7426 25601
rect 7110 25536 7116 25600
rect 7180 25536 7196 25600
rect 7260 25536 7276 25600
rect 7340 25536 7356 25600
rect 7420 25536 7426 25600
rect 7110 25535 7426 25536
rect 13826 25600 14142 25601
rect 13826 25536 13832 25600
rect 13896 25536 13912 25600
rect 13976 25536 13992 25600
rect 14056 25536 14072 25600
rect 14136 25536 14142 25600
rect 13826 25535 14142 25536
rect 20542 25600 20858 25601
rect 20542 25536 20548 25600
rect 20612 25536 20628 25600
rect 20692 25536 20708 25600
rect 20772 25536 20788 25600
rect 20852 25536 20858 25600
rect 20542 25535 20858 25536
rect 27258 25600 27574 25601
rect 27258 25536 27264 25600
rect 27328 25536 27344 25600
rect 27408 25536 27424 25600
rect 27488 25536 27504 25600
rect 27568 25536 27574 25600
rect 27258 25535 27574 25536
rect 3752 25056 4068 25057
rect 3752 24992 3758 25056
rect 3822 24992 3838 25056
rect 3902 24992 3918 25056
rect 3982 24992 3998 25056
rect 4062 24992 4068 25056
rect 3752 24991 4068 24992
rect 10468 25056 10784 25057
rect 10468 24992 10474 25056
rect 10538 24992 10554 25056
rect 10618 24992 10634 25056
rect 10698 24992 10714 25056
rect 10778 24992 10784 25056
rect 10468 24991 10784 24992
rect 17184 25056 17500 25057
rect 17184 24992 17190 25056
rect 17254 24992 17270 25056
rect 17334 24992 17350 25056
rect 17414 24992 17430 25056
rect 17494 24992 17500 25056
rect 17184 24991 17500 24992
rect 23900 25056 24216 25057
rect 23900 24992 23906 25056
rect 23970 24992 23986 25056
rect 24050 24992 24066 25056
rect 24130 24992 24146 25056
rect 24210 24992 24216 25056
rect 23900 24991 24216 24992
rect 6361 24850 6427 24853
rect 8109 24850 8175 24853
rect 15561 24850 15627 24853
rect 6361 24848 15627 24850
rect 6361 24792 6366 24848
rect 6422 24792 8114 24848
rect 8170 24792 15566 24848
rect 15622 24792 15627 24848
rect 6361 24790 15627 24792
rect 6361 24787 6427 24790
rect 8109 24787 8175 24790
rect 15561 24787 15627 24790
rect 6361 24714 6427 24717
rect 7649 24714 7715 24717
rect 6361 24712 7715 24714
rect 6361 24656 6366 24712
rect 6422 24656 7654 24712
rect 7710 24656 7715 24712
rect 6361 24654 7715 24656
rect 6361 24651 6427 24654
rect 7649 24651 7715 24654
rect 7110 24512 7426 24513
rect 7110 24448 7116 24512
rect 7180 24448 7196 24512
rect 7260 24448 7276 24512
rect 7340 24448 7356 24512
rect 7420 24448 7426 24512
rect 7110 24447 7426 24448
rect 13826 24512 14142 24513
rect 13826 24448 13832 24512
rect 13896 24448 13912 24512
rect 13976 24448 13992 24512
rect 14056 24448 14072 24512
rect 14136 24448 14142 24512
rect 13826 24447 14142 24448
rect 20542 24512 20858 24513
rect 20542 24448 20548 24512
rect 20612 24448 20628 24512
rect 20692 24448 20708 24512
rect 20772 24448 20788 24512
rect 20852 24448 20858 24512
rect 20542 24447 20858 24448
rect 27258 24512 27574 24513
rect 27258 24448 27264 24512
rect 27328 24448 27344 24512
rect 27408 24448 27424 24512
rect 27488 24448 27504 24512
rect 27568 24448 27574 24512
rect 27258 24447 27574 24448
rect 6361 24306 6427 24309
rect 7925 24306 7991 24309
rect 6361 24304 7991 24306
rect 6361 24248 6366 24304
rect 6422 24248 7930 24304
rect 7986 24248 7991 24304
rect 6361 24246 7991 24248
rect 6361 24243 6427 24246
rect 7925 24243 7991 24246
rect 6913 24034 6979 24037
rect 7833 24034 7899 24037
rect 6913 24032 7899 24034
rect 6913 23976 6918 24032
rect 6974 23976 7838 24032
rect 7894 23976 7899 24032
rect 6913 23974 7899 23976
rect 6913 23971 6979 23974
rect 7833 23971 7899 23974
rect 3752 23968 4068 23969
rect 3752 23904 3758 23968
rect 3822 23904 3838 23968
rect 3902 23904 3918 23968
rect 3982 23904 3998 23968
rect 4062 23904 4068 23968
rect 3752 23903 4068 23904
rect 10468 23968 10784 23969
rect 10468 23904 10474 23968
rect 10538 23904 10554 23968
rect 10618 23904 10634 23968
rect 10698 23904 10714 23968
rect 10778 23904 10784 23968
rect 10468 23903 10784 23904
rect 17184 23968 17500 23969
rect 17184 23904 17190 23968
rect 17254 23904 17270 23968
rect 17334 23904 17350 23968
rect 17414 23904 17430 23968
rect 17494 23904 17500 23968
rect 17184 23903 17500 23904
rect 23900 23968 24216 23969
rect 23900 23904 23906 23968
rect 23970 23904 23986 23968
rect 24050 23904 24066 23968
rect 24130 23904 24146 23968
rect 24210 23904 24216 23968
rect 23900 23903 24216 23904
rect 7110 23424 7426 23425
rect 7110 23360 7116 23424
rect 7180 23360 7196 23424
rect 7260 23360 7276 23424
rect 7340 23360 7356 23424
rect 7420 23360 7426 23424
rect 7110 23359 7426 23360
rect 13826 23424 14142 23425
rect 13826 23360 13832 23424
rect 13896 23360 13912 23424
rect 13976 23360 13992 23424
rect 14056 23360 14072 23424
rect 14136 23360 14142 23424
rect 13826 23359 14142 23360
rect 20542 23424 20858 23425
rect 20542 23360 20548 23424
rect 20612 23360 20628 23424
rect 20692 23360 20708 23424
rect 20772 23360 20788 23424
rect 20852 23360 20858 23424
rect 20542 23359 20858 23360
rect 27258 23424 27574 23425
rect 27258 23360 27264 23424
rect 27328 23360 27344 23424
rect 27408 23360 27424 23424
rect 27488 23360 27504 23424
rect 27568 23360 27574 23424
rect 27258 23359 27574 23360
rect 3752 22880 4068 22881
rect 3752 22816 3758 22880
rect 3822 22816 3838 22880
rect 3902 22816 3918 22880
rect 3982 22816 3998 22880
rect 4062 22816 4068 22880
rect 3752 22815 4068 22816
rect 10468 22880 10784 22881
rect 10468 22816 10474 22880
rect 10538 22816 10554 22880
rect 10618 22816 10634 22880
rect 10698 22816 10714 22880
rect 10778 22816 10784 22880
rect 10468 22815 10784 22816
rect 17184 22880 17500 22881
rect 17184 22816 17190 22880
rect 17254 22816 17270 22880
rect 17334 22816 17350 22880
rect 17414 22816 17430 22880
rect 17494 22816 17500 22880
rect 17184 22815 17500 22816
rect 23900 22880 24216 22881
rect 23900 22816 23906 22880
rect 23970 22816 23986 22880
rect 24050 22816 24066 22880
rect 24130 22816 24146 22880
rect 24210 22816 24216 22880
rect 23900 22815 24216 22816
rect 7110 22336 7426 22337
rect 7110 22272 7116 22336
rect 7180 22272 7196 22336
rect 7260 22272 7276 22336
rect 7340 22272 7356 22336
rect 7420 22272 7426 22336
rect 7110 22271 7426 22272
rect 13826 22336 14142 22337
rect 13826 22272 13832 22336
rect 13896 22272 13912 22336
rect 13976 22272 13992 22336
rect 14056 22272 14072 22336
rect 14136 22272 14142 22336
rect 13826 22271 14142 22272
rect 20542 22336 20858 22337
rect 20542 22272 20548 22336
rect 20612 22272 20628 22336
rect 20692 22272 20708 22336
rect 20772 22272 20788 22336
rect 20852 22272 20858 22336
rect 20542 22271 20858 22272
rect 27258 22336 27574 22337
rect 27258 22272 27264 22336
rect 27328 22272 27344 22336
rect 27408 22272 27424 22336
rect 27488 22272 27504 22336
rect 27568 22272 27574 22336
rect 27258 22271 27574 22272
rect 10961 21994 11027 21997
rect 18045 21994 18111 21997
rect 10961 21992 18111 21994
rect 10961 21936 10966 21992
rect 11022 21936 18050 21992
rect 18106 21936 18111 21992
rect 10961 21934 18111 21936
rect 10961 21931 11027 21934
rect 18045 21931 18111 21934
rect 3752 21792 4068 21793
rect 3752 21728 3758 21792
rect 3822 21728 3838 21792
rect 3902 21728 3918 21792
rect 3982 21728 3998 21792
rect 4062 21728 4068 21792
rect 3752 21727 4068 21728
rect 10468 21792 10784 21793
rect 10468 21728 10474 21792
rect 10538 21728 10554 21792
rect 10618 21728 10634 21792
rect 10698 21728 10714 21792
rect 10778 21728 10784 21792
rect 10468 21727 10784 21728
rect 17184 21792 17500 21793
rect 17184 21728 17190 21792
rect 17254 21728 17270 21792
rect 17334 21728 17350 21792
rect 17414 21728 17430 21792
rect 17494 21728 17500 21792
rect 17184 21727 17500 21728
rect 23900 21792 24216 21793
rect 23900 21728 23906 21792
rect 23970 21728 23986 21792
rect 24050 21728 24066 21792
rect 24130 21728 24146 21792
rect 24210 21728 24216 21792
rect 23900 21727 24216 21728
rect 7110 21248 7426 21249
rect 7110 21184 7116 21248
rect 7180 21184 7196 21248
rect 7260 21184 7276 21248
rect 7340 21184 7356 21248
rect 7420 21184 7426 21248
rect 7110 21183 7426 21184
rect 13826 21248 14142 21249
rect 13826 21184 13832 21248
rect 13896 21184 13912 21248
rect 13976 21184 13992 21248
rect 14056 21184 14072 21248
rect 14136 21184 14142 21248
rect 13826 21183 14142 21184
rect 20542 21248 20858 21249
rect 20542 21184 20548 21248
rect 20612 21184 20628 21248
rect 20692 21184 20708 21248
rect 20772 21184 20788 21248
rect 20852 21184 20858 21248
rect 20542 21183 20858 21184
rect 27258 21248 27574 21249
rect 27258 21184 27264 21248
rect 27328 21184 27344 21248
rect 27408 21184 27424 21248
rect 27488 21184 27504 21248
rect 27568 21184 27574 21248
rect 27258 21183 27574 21184
rect 3752 20704 4068 20705
rect 3752 20640 3758 20704
rect 3822 20640 3838 20704
rect 3902 20640 3918 20704
rect 3982 20640 3998 20704
rect 4062 20640 4068 20704
rect 3752 20639 4068 20640
rect 10468 20704 10784 20705
rect 10468 20640 10474 20704
rect 10538 20640 10554 20704
rect 10618 20640 10634 20704
rect 10698 20640 10714 20704
rect 10778 20640 10784 20704
rect 10468 20639 10784 20640
rect 17184 20704 17500 20705
rect 17184 20640 17190 20704
rect 17254 20640 17270 20704
rect 17334 20640 17350 20704
rect 17414 20640 17430 20704
rect 17494 20640 17500 20704
rect 17184 20639 17500 20640
rect 23900 20704 24216 20705
rect 23900 20640 23906 20704
rect 23970 20640 23986 20704
rect 24050 20640 24066 20704
rect 24130 20640 24146 20704
rect 24210 20640 24216 20704
rect 23900 20639 24216 20640
rect 7110 20160 7426 20161
rect 7110 20096 7116 20160
rect 7180 20096 7196 20160
rect 7260 20096 7276 20160
rect 7340 20096 7356 20160
rect 7420 20096 7426 20160
rect 7110 20095 7426 20096
rect 13826 20160 14142 20161
rect 13826 20096 13832 20160
rect 13896 20096 13912 20160
rect 13976 20096 13992 20160
rect 14056 20096 14072 20160
rect 14136 20096 14142 20160
rect 13826 20095 14142 20096
rect 20542 20160 20858 20161
rect 20542 20096 20548 20160
rect 20612 20096 20628 20160
rect 20692 20096 20708 20160
rect 20772 20096 20788 20160
rect 20852 20096 20858 20160
rect 20542 20095 20858 20096
rect 27258 20160 27574 20161
rect 27258 20096 27264 20160
rect 27328 20096 27344 20160
rect 27408 20096 27424 20160
rect 27488 20096 27504 20160
rect 27568 20096 27574 20160
rect 27258 20095 27574 20096
rect 12985 19818 13051 19821
rect 18505 19818 18571 19821
rect 12985 19816 18571 19818
rect 12985 19760 12990 19816
rect 13046 19760 18510 19816
rect 18566 19760 18571 19816
rect 12985 19758 18571 19760
rect 12985 19755 13051 19758
rect 18505 19755 18571 19758
rect 3752 19616 4068 19617
rect 3752 19552 3758 19616
rect 3822 19552 3838 19616
rect 3902 19552 3918 19616
rect 3982 19552 3998 19616
rect 4062 19552 4068 19616
rect 3752 19551 4068 19552
rect 10468 19616 10784 19617
rect 10468 19552 10474 19616
rect 10538 19552 10554 19616
rect 10618 19552 10634 19616
rect 10698 19552 10714 19616
rect 10778 19552 10784 19616
rect 10468 19551 10784 19552
rect 17184 19616 17500 19617
rect 17184 19552 17190 19616
rect 17254 19552 17270 19616
rect 17334 19552 17350 19616
rect 17414 19552 17430 19616
rect 17494 19552 17500 19616
rect 17184 19551 17500 19552
rect 23900 19616 24216 19617
rect 23900 19552 23906 19616
rect 23970 19552 23986 19616
rect 24050 19552 24066 19616
rect 24130 19552 24146 19616
rect 24210 19552 24216 19616
rect 23900 19551 24216 19552
rect 14917 19410 14983 19413
rect 18321 19410 18387 19413
rect 14917 19408 18387 19410
rect 14917 19352 14922 19408
rect 14978 19352 18326 19408
rect 18382 19352 18387 19408
rect 14917 19350 18387 19352
rect 14917 19347 14983 19350
rect 18321 19347 18387 19350
rect 7110 19072 7426 19073
rect 7110 19008 7116 19072
rect 7180 19008 7196 19072
rect 7260 19008 7276 19072
rect 7340 19008 7356 19072
rect 7420 19008 7426 19072
rect 7110 19007 7426 19008
rect 13826 19072 14142 19073
rect 13826 19008 13832 19072
rect 13896 19008 13912 19072
rect 13976 19008 13992 19072
rect 14056 19008 14072 19072
rect 14136 19008 14142 19072
rect 13826 19007 14142 19008
rect 20542 19072 20858 19073
rect 20542 19008 20548 19072
rect 20612 19008 20628 19072
rect 20692 19008 20708 19072
rect 20772 19008 20788 19072
rect 20852 19008 20858 19072
rect 20542 19007 20858 19008
rect 27258 19072 27574 19073
rect 27258 19008 27264 19072
rect 27328 19008 27344 19072
rect 27408 19008 27424 19072
rect 27488 19008 27504 19072
rect 27568 19008 27574 19072
rect 27258 19007 27574 19008
rect 3752 18528 4068 18529
rect 3752 18464 3758 18528
rect 3822 18464 3838 18528
rect 3902 18464 3918 18528
rect 3982 18464 3998 18528
rect 4062 18464 4068 18528
rect 3752 18463 4068 18464
rect 10468 18528 10784 18529
rect 10468 18464 10474 18528
rect 10538 18464 10554 18528
rect 10618 18464 10634 18528
rect 10698 18464 10714 18528
rect 10778 18464 10784 18528
rect 10468 18463 10784 18464
rect 17184 18528 17500 18529
rect 17184 18464 17190 18528
rect 17254 18464 17270 18528
rect 17334 18464 17350 18528
rect 17414 18464 17430 18528
rect 17494 18464 17500 18528
rect 17184 18463 17500 18464
rect 23900 18528 24216 18529
rect 23900 18464 23906 18528
rect 23970 18464 23986 18528
rect 24050 18464 24066 18528
rect 24130 18464 24146 18528
rect 24210 18464 24216 18528
rect 23900 18463 24216 18464
rect 7110 17984 7426 17985
rect 7110 17920 7116 17984
rect 7180 17920 7196 17984
rect 7260 17920 7276 17984
rect 7340 17920 7356 17984
rect 7420 17920 7426 17984
rect 7110 17919 7426 17920
rect 13826 17984 14142 17985
rect 13826 17920 13832 17984
rect 13896 17920 13912 17984
rect 13976 17920 13992 17984
rect 14056 17920 14072 17984
rect 14136 17920 14142 17984
rect 13826 17919 14142 17920
rect 20542 17984 20858 17985
rect 20542 17920 20548 17984
rect 20612 17920 20628 17984
rect 20692 17920 20708 17984
rect 20772 17920 20788 17984
rect 20852 17920 20858 17984
rect 20542 17919 20858 17920
rect 27258 17984 27574 17985
rect 27258 17920 27264 17984
rect 27328 17920 27344 17984
rect 27408 17920 27424 17984
rect 27488 17920 27504 17984
rect 27568 17920 27574 17984
rect 27258 17919 27574 17920
rect 3752 17440 4068 17441
rect 3752 17376 3758 17440
rect 3822 17376 3838 17440
rect 3902 17376 3918 17440
rect 3982 17376 3998 17440
rect 4062 17376 4068 17440
rect 3752 17375 4068 17376
rect 10468 17440 10784 17441
rect 10468 17376 10474 17440
rect 10538 17376 10554 17440
rect 10618 17376 10634 17440
rect 10698 17376 10714 17440
rect 10778 17376 10784 17440
rect 10468 17375 10784 17376
rect 17184 17440 17500 17441
rect 17184 17376 17190 17440
rect 17254 17376 17270 17440
rect 17334 17376 17350 17440
rect 17414 17376 17430 17440
rect 17494 17376 17500 17440
rect 17184 17375 17500 17376
rect 23900 17440 24216 17441
rect 23900 17376 23906 17440
rect 23970 17376 23986 17440
rect 24050 17376 24066 17440
rect 24130 17376 24146 17440
rect 24210 17376 24216 17440
rect 23900 17375 24216 17376
rect 8477 17234 8543 17237
rect 10501 17234 10567 17237
rect 8477 17232 10567 17234
rect 8477 17176 8482 17232
rect 8538 17176 10506 17232
rect 10562 17176 10567 17232
rect 8477 17174 10567 17176
rect 8477 17171 8543 17174
rect 10501 17171 10567 17174
rect 23933 17234 23999 17237
rect 24945 17234 25011 17237
rect 23933 17232 25011 17234
rect 23933 17176 23938 17232
rect 23994 17176 24950 17232
rect 25006 17176 25011 17232
rect 23933 17174 25011 17176
rect 23933 17171 23999 17174
rect 24945 17171 25011 17174
rect 16113 17098 16179 17101
rect 24894 17098 24900 17100
rect 16113 17096 24900 17098
rect 16113 17040 16118 17096
rect 16174 17040 24900 17096
rect 16113 17038 24900 17040
rect 16113 17035 16179 17038
rect 24894 17036 24900 17038
rect 24964 17036 24970 17100
rect 24209 16962 24275 16965
rect 24669 16962 24735 16965
rect 24209 16960 24735 16962
rect 24209 16904 24214 16960
rect 24270 16904 24674 16960
rect 24730 16904 24735 16960
rect 24209 16902 24735 16904
rect 24209 16899 24275 16902
rect 24669 16899 24735 16902
rect 7110 16896 7426 16897
rect 7110 16832 7116 16896
rect 7180 16832 7196 16896
rect 7260 16832 7276 16896
rect 7340 16832 7356 16896
rect 7420 16832 7426 16896
rect 7110 16831 7426 16832
rect 13826 16896 14142 16897
rect 13826 16832 13832 16896
rect 13896 16832 13912 16896
rect 13976 16832 13992 16896
rect 14056 16832 14072 16896
rect 14136 16832 14142 16896
rect 13826 16831 14142 16832
rect 20542 16896 20858 16897
rect 20542 16832 20548 16896
rect 20612 16832 20628 16896
rect 20692 16832 20708 16896
rect 20772 16832 20788 16896
rect 20852 16832 20858 16896
rect 20542 16831 20858 16832
rect 27258 16896 27574 16897
rect 27258 16832 27264 16896
rect 27328 16832 27344 16896
rect 27408 16832 27424 16896
rect 27488 16832 27504 16896
rect 27568 16832 27574 16896
rect 27258 16831 27574 16832
rect 3752 16352 4068 16353
rect 3752 16288 3758 16352
rect 3822 16288 3838 16352
rect 3902 16288 3918 16352
rect 3982 16288 3998 16352
rect 4062 16288 4068 16352
rect 3752 16287 4068 16288
rect 10468 16352 10784 16353
rect 10468 16288 10474 16352
rect 10538 16288 10554 16352
rect 10618 16288 10634 16352
rect 10698 16288 10714 16352
rect 10778 16288 10784 16352
rect 10468 16287 10784 16288
rect 17184 16352 17500 16353
rect 17184 16288 17190 16352
rect 17254 16288 17270 16352
rect 17334 16288 17350 16352
rect 17414 16288 17430 16352
rect 17494 16288 17500 16352
rect 17184 16287 17500 16288
rect 23900 16352 24216 16353
rect 23900 16288 23906 16352
rect 23970 16288 23986 16352
rect 24050 16288 24066 16352
rect 24130 16288 24146 16352
rect 24210 16288 24216 16352
rect 23900 16287 24216 16288
rect 10685 16010 10751 16013
rect 14641 16010 14707 16013
rect 15469 16010 15535 16013
rect 10685 16008 15535 16010
rect 10685 15952 10690 16008
rect 10746 15952 14646 16008
rect 14702 15952 15474 16008
rect 15530 15952 15535 16008
rect 10685 15950 15535 15952
rect 10685 15947 10751 15950
rect 14641 15947 14707 15950
rect 15469 15947 15535 15950
rect 7110 15808 7426 15809
rect 7110 15744 7116 15808
rect 7180 15744 7196 15808
rect 7260 15744 7276 15808
rect 7340 15744 7356 15808
rect 7420 15744 7426 15808
rect 7110 15743 7426 15744
rect 13826 15808 14142 15809
rect 13826 15744 13832 15808
rect 13896 15744 13912 15808
rect 13976 15744 13992 15808
rect 14056 15744 14072 15808
rect 14136 15744 14142 15808
rect 13826 15743 14142 15744
rect 20542 15808 20858 15809
rect 20542 15744 20548 15808
rect 20612 15744 20628 15808
rect 20692 15744 20708 15808
rect 20772 15744 20788 15808
rect 20852 15744 20858 15808
rect 20542 15743 20858 15744
rect 27258 15808 27574 15809
rect 27258 15744 27264 15808
rect 27328 15744 27344 15808
rect 27408 15744 27424 15808
rect 27488 15744 27504 15808
rect 27568 15744 27574 15808
rect 27258 15743 27574 15744
rect 3752 15264 4068 15265
rect 3752 15200 3758 15264
rect 3822 15200 3838 15264
rect 3902 15200 3918 15264
rect 3982 15200 3998 15264
rect 4062 15200 4068 15264
rect 3752 15199 4068 15200
rect 10468 15264 10784 15265
rect 10468 15200 10474 15264
rect 10538 15200 10554 15264
rect 10618 15200 10634 15264
rect 10698 15200 10714 15264
rect 10778 15200 10784 15264
rect 10468 15199 10784 15200
rect 17184 15264 17500 15265
rect 17184 15200 17190 15264
rect 17254 15200 17270 15264
rect 17334 15200 17350 15264
rect 17414 15200 17430 15264
rect 17494 15200 17500 15264
rect 17184 15199 17500 15200
rect 23900 15264 24216 15265
rect 23900 15200 23906 15264
rect 23970 15200 23986 15264
rect 24050 15200 24066 15264
rect 24130 15200 24146 15264
rect 24210 15200 24216 15264
rect 23900 15199 24216 15200
rect 7110 14720 7426 14721
rect 7110 14656 7116 14720
rect 7180 14656 7196 14720
rect 7260 14656 7276 14720
rect 7340 14656 7356 14720
rect 7420 14656 7426 14720
rect 7110 14655 7426 14656
rect 13826 14720 14142 14721
rect 13826 14656 13832 14720
rect 13896 14656 13912 14720
rect 13976 14656 13992 14720
rect 14056 14656 14072 14720
rect 14136 14656 14142 14720
rect 13826 14655 14142 14656
rect 20542 14720 20858 14721
rect 20542 14656 20548 14720
rect 20612 14656 20628 14720
rect 20692 14656 20708 14720
rect 20772 14656 20788 14720
rect 20852 14656 20858 14720
rect 20542 14655 20858 14656
rect 27258 14720 27574 14721
rect 27258 14656 27264 14720
rect 27328 14656 27344 14720
rect 27408 14656 27424 14720
rect 27488 14656 27504 14720
rect 27568 14656 27574 14720
rect 27258 14655 27574 14656
rect 9857 14378 9923 14381
rect 10225 14378 10291 14381
rect 12709 14378 12775 14381
rect 18321 14378 18387 14381
rect 9857 14376 18387 14378
rect 9857 14320 9862 14376
rect 9918 14320 10230 14376
rect 10286 14320 12714 14376
rect 12770 14320 18326 14376
rect 18382 14320 18387 14376
rect 9857 14318 18387 14320
rect 9857 14315 9923 14318
rect 10225 14315 10291 14318
rect 12709 14315 12775 14318
rect 18321 14315 18387 14318
rect 3752 14176 4068 14177
rect 3752 14112 3758 14176
rect 3822 14112 3838 14176
rect 3902 14112 3918 14176
rect 3982 14112 3998 14176
rect 4062 14112 4068 14176
rect 3752 14111 4068 14112
rect 10468 14176 10784 14177
rect 10468 14112 10474 14176
rect 10538 14112 10554 14176
rect 10618 14112 10634 14176
rect 10698 14112 10714 14176
rect 10778 14112 10784 14176
rect 10468 14111 10784 14112
rect 17184 14176 17500 14177
rect 17184 14112 17190 14176
rect 17254 14112 17270 14176
rect 17334 14112 17350 14176
rect 17414 14112 17430 14176
rect 17494 14112 17500 14176
rect 17184 14111 17500 14112
rect 23900 14176 24216 14177
rect 23900 14112 23906 14176
rect 23970 14112 23986 14176
rect 24050 14112 24066 14176
rect 24130 14112 24146 14176
rect 24210 14112 24216 14176
rect 23900 14111 24216 14112
rect 7110 13632 7426 13633
rect 7110 13568 7116 13632
rect 7180 13568 7196 13632
rect 7260 13568 7276 13632
rect 7340 13568 7356 13632
rect 7420 13568 7426 13632
rect 7110 13567 7426 13568
rect 13826 13632 14142 13633
rect 13826 13568 13832 13632
rect 13896 13568 13912 13632
rect 13976 13568 13992 13632
rect 14056 13568 14072 13632
rect 14136 13568 14142 13632
rect 13826 13567 14142 13568
rect 20542 13632 20858 13633
rect 20542 13568 20548 13632
rect 20612 13568 20628 13632
rect 20692 13568 20708 13632
rect 20772 13568 20788 13632
rect 20852 13568 20858 13632
rect 20542 13567 20858 13568
rect 27258 13632 27574 13633
rect 27258 13568 27264 13632
rect 27328 13568 27344 13632
rect 27408 13568 27424 13632
rect 27488 13568 27504 13632
rect 27568 13568 27574 13632
rect 27258 13567 27574 13568
rect 3752 13088 4068 13089
rect 3752 13024 3758 13088
rect 3822 13024 3838 13088
rect 3902 13024 3918 13088
rect 3982 13024 3998 13088
rect 4062 13024 4068 13088
rect 3752 13023 4068 13024
rect 10468 13088 10784 13089
rect 10468 13024 10474 13088
rect 10538 13024 10554 13088
rect 10618 13024 10634 13088
rect 10698 13024 10714 13088
rect 10778 13024 10784 13088
rect 10468 13023 10784 13024
rect 17184 13088 17500 13089
rect 17184 13024 17190 13088
rect 17254 13024 17270 13088
rect 17334 13024 17350 13088
rect 17414 13024 17430 13088
rect 17494 13024 17500 13088
rect 17184 13023 17500 13024
rect 23900 13088 24216 13089
rect 23900 13024 23906 13088
rect 23970 13024 23986 13088
rect 24050 13024 24066 13088
rect 24130 13024 24146 13088
rect 24210 13024 24216 13088
rect 23900 13023 24216 13024
rect 7110 12544 7426 12545
rect 7110 12480 7116 12544
rect 7180 12480 7196 12544
rect 7260 12480 7276 12544
rect 7340 12480 7356 12544
rect 7420 12480 7426 12544
rect 7110 12479 7426 12480
rect 13826 12544 14142 12545
rect 13826 12480 13832 12544
rect 13896 12480 13912 12544
rect 13976 12480 13992 12544
rect 14056 12480 14072 12544
rect 14136 12480 14142 12544
rect 13826 12479 14142 12480
rect 20542 12544 20858 12545
rect 20542 12480 20548 12544
rect 20612 12480 20628 12544
rect 20692 12480 20708 12544
rect 20772 12480 20788 12544
rect 20852 12480 20858 12544
rect 20542 12479 20858 12480
rect 27258 12544 27574 12545
rect 27258 12480 27264 12544
rect 27328 12480 27344 12544
rect 27408 12480 27424 12544
rect 27488 12480 27504 12544
rect 27568 12480 27574 12544
rect 27258 12479 27574 12480
rect 3752 12000 4068 12001
rect 3752 11936 3758 12000
rect 3822 11936 3838 12000
rect 3902 11936 3918 12000
rect 3982 11936 3998 12000
rect 4062 11936 4068 12000
rect 3752 11935 4068 11936
rect 10468 12000 10784 12001
rect 10468 11936 10474 12000
rect 10538 11936 10554 12000
rect 10618 11936 10634 12000
rect 10698 11936 10714 12000
rect 10778 11936 10784 12000
rect 10468 11935 10784 11936
rect 17184 12000 17500 12001
rect 17184 11936 17190 12000
rect 17254 11936 17270 12000
rect 17334 11936 17350 12000
rect 17414 11936 17430 12000
rect 17494 11936 17500 12000
rect 17184 11935 17500 11936
rect 23900 12000 24216 12001
rect 23900 11936 23906 12000
rect 23970 11936 23986 12000
rect 24050 11936 24066 12000
rect 24130 11936 24146 12000
rect 24210 11936 24216 12000
rect 23900 11935 24216 11936
rect 7110 11456 7426 11457
rect 7110 11392 7116 11456
rect 7180 11392 7196 11456
rect 7260 11392 7276 11456
rect 7340 11392 7356 11456
rect 7420 11392 7426 11456
rect 7110 11391 7426 11392
rect 13826 11456 14142 11457
rect 13826 11392 13832 11456
rect 13896 11392 13912 11456
rect 13976 11392 13992 11456
rect 14056 11392 14072 11456
rect 14136 11392 14142 11456
rect 13826 11391 14142 11392
rect 20542 11456 20858 11457
rect 20542 11392 20548 11456
rect 20612 11392 20628 11456
rect 20692 11392 20708 11456
rect 20772 11392 20788 11456
rect 20852 11392 20858 11456
rect 20542 11391 20858 11392
rect 27258 11456 27574 11457
rect 27258 11392 27264 11456
rect 27328 11392 27344 11456
rect 27408 11392 27424 11456
rect 27488 11392 27504 11456
rect 27568 11392 27574 11456
rect 27258 11391 27574 11392
rect 3752 10912 4068 10913
rect 3752 10848 3758 10912
rect 3822 10848 3838 10912
rect 3902 10848 3918 10912
rect 3982 10848 3998 10912
rect 4062 10848 4068 10912
rect 3752 10847 4068 10848
rect 10468 10912 10784 10913
rect 10468 10848 10474 10912
rect 10538 10848 10554 10912
rect 10618 10848 10634 10912
rect 10698 10848 10714 10912
rect 10778 10848 10784 10912
rect 10468 10847 10784 10848
rect 17184 10912 17500 10913
rect 17184 10848 17190 10912
rect 17254 10848 17270 10912
rect 17334 10848 17350 10912
rect 17414 10848 17430 10912
rect 17494 10848 17500 10912
rect 17184 10847 17500 10848
rect 23900 10912 24216 10913
rect 23900 10848 23906 10912
rect 23970 10848 23986 10912
rect 24050 10848 24066 10912
rect 24130 10848 24146 10912
rect 24210 10848 24216 10912
rect 23900 10847 24216 10848
rect 2078 10508 2084 10572
rect 2148 10570 2154 10572
rect 20345 10570 20411 10573
rect 2148 10568 20411 10570
rect 2148 10512 20350 10568
rect 20406 10512 20411 10568
rect 2148 10510 20411 10512
rect 2148 10508 2154 10510
rect 20345 10507 20411 10510
rect 7110 10368 7426 10369
rect 7110 10304 7116 10368
rect 7180 10304 7196 10368
rect 7260 10304 7276 10368
rect 7340 10304 7356 10368
rect 7420 10304 7426 10368
rect 7110 10303 7426 10304
rect 13826 10368 14142 10369
rect 13826 10304 13832 10368
rect 13896 10304 13912 10368
rect 13976 10304 13992 10368
rect 14056 10304 14072 10368
rect 14136 10304 14142 10368
rect 13826 10303 14142 10304
rect 20542 10368 20858 10369
rect 20542 10304 20548 10368
rect 20612 10304 20628 10368
rect 20692 10304 20708 10368
rect 20772 10304 20788 10368
rect 20852 10304 20858 10368
rect 20542 10303 20858 10304
rect 27258 10368 27574 10369
rect 27258 10304 27264 10368
rect 27328 10304 27344 10368
rect 27408 10304 27424 10368
rect 27488 10304 27504 10368
rect 27568 10304 27574 10368
rect 27258 10303 27574 10304
rect 3752 9824 4068 9825
rect 3752 9760 3758 9824
rect 3822 9760 3838 9824
rect 3902 9760 3918 9824
rect 3982 9760 3998 9824
rect 4062 9760 4068 9824
rect 3752 9759 4068 9760
rect 10468 9824 10784 9825
rect 10468 9760 10474 9824
rect 10538 9760 10554 9824
rect 10618 9760 10634 9824
rect 10698 9760 10714 9824
rect 10778 9760 10784 9824
rect 10468 9759 10784 9760
rect 17184 9824 17500 9825
rect 17184 9760 17190 9824
rect 17254 9760 17270 9824
rect 17334 9760 17350 9824
rect 17414 9760 17430 9824
rect 17494 9760 17500 9824
rect 17184 9759 17500 9760
rect 23900 9824 24216 9825
rect 23900 9760 23906 9824
rect 23970 9760 23986 9824
rect 24050 9760 24066 9824
rect 24130 9760 24146 9824
rect 24210 9760 24216 9824
rect 23900 9759 24216 9760
rect 7110 9280 7426 9281
rect 7110 9216 7116 9280
rect 7180 9216 7196 9280
rect 7260 9216 7276 9280
rect 7340 9216 7356 9280
rect 7420 9216 7426 9280
rect 7110 9215 7426 9216
rect 13826 9280 14142 9281
rect 13826 9216 13832 9280
rect 13896 9216 13912 9280
rect 13976 9216 13992 9280
rect 14056 9216 14072 9280
rect 14136 9216 14142 9280
rect 13826 9215 14142 9216
rect 20542 9280 20858 9281
rect 20542 9216 20548 9280
rect 20612 9216 20628 9280
rect 20692 9216 20708 9280
rect 20772 9216 20788 9280
rect 20852 9216 20858 9280
rect 20542 9215 20858 9216
rect 27258 9280 27574 9281
rect 27258 9216 27264 9280
rect 27328 9216 27344 9280
rect 27408 9216 27424 9280
rect 27488 9216 27504 9280
rect 27568 9216 27574 9280
rect 27258 9215 27574 9216
rect 3752 8736 4068 8737
rect 3752 8672 3758 8736
rect 3822 8672 3838 8736
rect 3902 8672 3918 8736
rect 3982 8672 3998 8736
rect 4062 8672 4068 8736
rect 3752 8671 4068 8672
rect 10468 8736 10784 8737
rect 10468 8672 10474 8736
rect 10538 8672 10554 8736
rect 10618 8672 10634 8736
rect 10698 8672 10714 8736
rect 10778 8672 10784 8736
rect 10468 8671 10784 8672
rect 17184 8736 17500 8737
rect 17184 8672 17190 8736
rect 17254 8672 17270 8736
rect 17334 8672 17350 8736
rect 17414 8672 17430 8736
rect 17494 8672 17500 8736
rect 17184 8671 17500 8672
rect 23900 8736 24216 8737
rect 23900 8672 23906 8736
rect 23970 8672 23986 8736
rect 24050 8672 24066 8736
rect 24130 8672 24146 8736
rect 24210 8672 24216 8736
rect 23900 8671 24216 8672
rect 7110 8192 7426 8193
rect 7110 8128 7116 8192
rect 7180 8128 7196 8192
rect 7260 8128 7276 8192
rect 7340 8128 7356 8192
rect 7420 8128 7426 8192
rect 7110 8127 7426 8128
rect 13826 8192 14142 8193
rect 13826 8128 13832 8192
rect 13896 8128 13912 8192
rect 13976 8128 13992 8192
rect 14056 8128 14072 8192
rect 14136 8128 14142 8192
rect 13826 8127 14142 8128
rect 20542 8192 20858 8193
rect 20542 8128 20548 8192
rect 20612 8128 20628 8192
rect 20692 8128 20708 8192
rect 20772 8128 20788 8192
rect 20852 8128 20858 8192
rect 20542 8127 20858 8128
rect 27258 8192 27574 8193
rect 27258 8128 27264 8192
rect 27328 8128 27344 8192
rect 27408 8128 27424 8192
rect 27488 8128 27504 8192
rect 27568 8128 27574 8192
rect 27258 8127 27574 8128
rect 3752 7648 4068 7649
rect 3752 7584 3758 7648
rect 3822 7584 3838 7648
rect 3902 7584 3918 7648
rect 3982 7584 3998 7648
rect 4062 7584 4068 7648
rect 3752 7583 4068 7584
rect 10468 7648 10784 7649
rect 10468 7584 10474 7648
rect 10538 7584 10554 7648
rect 10618 7584 10634 7648
rect 10698 7584 10714 7648
rect 10778 7584 10784 7648
rect 10468 7583 10784 7584
rect 17184 7648 17500 7649
rect 17184 7584 17190 7648
rect 17254 7584 17270 7648
rect 17334 7584 17350 7648
rect 17414 7584 17430 7648
rect 17494 7584 17500 7648
rect 17184 7583 17500 7584
rect 23900 7648 24216 7649
rect 23900 7584 23906 7648
rect 23970 7584 23986 7648
rect 24050 7584 24066 7648
rect 24130 7584 24146 7648
rect 24210 7584 24216 7648
rect 23900 7583 24216 7584
rect 1894 7244 1900 7308
rect 1964 7306 1970 7308
rect 9857 7306 9923 7309
rect 1964 7304 9923 7306
rect 1964 7248 9862 7304
rect 9918 7248 9923 7304
rect 1964 7246 9923 7248
rect 1964 7244 1970 7246
rect 9857 7243 9923 7246
rect 11881 7170 11947 7173
rect 12985 7170 13051 7173
rect 11881 7168 13051 7170
rect 11881 7112 11886 7168
rect 11942 7112 12990 7168
rect 13046 7112 13051 7168
rect 11881 7110 13051 7112
rect 11881 7107 11947 7110
rect 12985 7107 13051 7110
rect 7110 7104 7426 7105
rect 7110 7040 7116 7104
rect 7180 7040 7196 7104
rect 7260 7040 7276 7104
rect 7340 7040 7356 7104
rect 7420 7040 7426 7104
rect 7110 7039 7426 7040
rect 13826 7104 14142 7105
rect 13826 7040 13832 7104
rect 13896 7040 13912 7104
rect 13976 7040 13992 7104
rect 14056 7040 14072 7104
rect 14136 7040 14142 7104
rect 13826 7039 14142 7040
rect 20542 7104 20858 7105
rect 20542 7040 20548 7104
rect 20612 7040 20628 7104
rect 20692 7040 20708 7104
rect 20772 7040 20788 7104
rect 20852 7040 20858 7104
rect 20542 7039 20858 7040
rect 27258 7104 27574 7105
rect 27258 7040 27264 7104
rect 27328 7040 27344 7104
rect 27408 7040 27424 7104
rect 27488 7040 27504 7104
rect 27568 7040 27574 7104
rect 27258 7039 27574 7040
rect 3752 6560 4068 6561
rect 3752 6496 3758 6560
rect 3822 6496 3838 6560
rect 3902 6496 3918 6560
rect 3982 6496 3998 6560
rect 4062 6496 4068 6560
rect 3752 6495 4068 6496
rect 10468 6560 10784 6561
rect 10468 6496 10474 6560
rect 10538 6496 10554 6560
rect 10618 6496 10634 6560
rect 10698 6496 10714 6560
rect 10778 6496 10784 6560
rect 10468 6495 10784 6496
rect 17184 6560 17500 6561
rect 17184 6496 17190 6560
rect 17254 6496 17270 6560
rect 17334 6496 17350 6560
rect 17414 6496 17430 6560
rect 17494 6496 17500 6560
rect 17184 6495 17500 6496
rect 23900 6560 24216 6561
rect 23900 6496 23906 6560
rect 23970 6496 23986 6560
rect 24050 6496 24066 6560
rect 24130 6496 24146 6560
rect 24210 6496 24216 6560
rect 23900 6495 24216 6496
rect 14365 6490 14431 6493
rect 15193 6490 15259 6493
rect 14365 6488 15259 6490
rect 14365 6432 14370 6488
rect 14426 6432 15198 6488
rect 15254 6432 15259 6488
rect 14365 6430 15259 6432
rect 14365 6427 14431 6430
rect 15193 6427 15259 6430
rect 14089 6218 14155 6221
rect 15101 6218 15167 6221
rect 14089 6216 15167 6218
rect 14089 6160 14094 6216
rect 14150 6160 15106 6216
rect 15162 6160 15167 6216
rect 14089 6158 15167 6160
rect 14089 6155 14155 6158
rect 15101 6155 15167 6158
rect 7110 6016 7426 6017
rect 7110 5952 7116 6016
rect 7180 5952 7196 6016
rect 7260 5952 7276 6016
rect 7340 5952 7356 6016
rect 7420 5952 7426 6016
rect 7110 5951 7426 5952
rect 13826 6016 14142 6017
rect 13826 5952 13832 6016
rect 13896 5952 13912 6016
rect 13976 5952 13992 6016
rect 14056 5952 14072 6016
rect 14136 5952 14142 6016
rect 13826 5951 14142 5952
rect 20542 6016 20858 6017
rect 20542 5952 20548 6016
rect 20612 5952 20628 6016
rect 20692 5952 20708 6016
rect 20772 5952 20788 6016
rect 20852 5952 20858 6016
rect 20542 5951 20858 5952
rect 27258 6016 27574 6017
rect 27258 5952 27264 6016
rect 27328 5952 27344 6016
rect 27408 5952 27424 6016
rect 27488 5952 27504 6016
rect 27568 5952 27574 6016
rect 27258 5951 27574 5952
rect 3752 5472 4068 5473
rect 3752 5408 3758 5472
rect 3822 5408 3838 5472
rect 3902 5408 3918 5472
rect 3982 5408 3998 5472
rect 4062 5408 4068 5472
rect 3752 5407 4068 5408
rect 10468 5472 10784 5473
rect 10468 5408 10474 5472
rect 10538 5408 10554 5472
rect 10618 5408 10634 5472
rect 10698 5408 10714 5472
rect 10778 5408 10784 5472
rect 10468 5407 10784 5408
rect 17184 5472 17500 5473
rect 17184 5408 17190 5472
rect 17254 5408 17270 5472
rect 17334 5408 17350 5472
rect 17414 5408 17430 5472
rect 17494 5408 17500 5472
rect 17184 5407 17500 5408
rect 23900 5472 24216 5473
rect 23900 5408 23906 5472
rect 23970 5408 23986 5472
rect 24050 5408 24066 5472
rect 24130 5408 24146 5472
rect 24210 5408 24216 5472
rect 23900 5407 24216 5408
rect 7110 4928 7426 4929
rect 7110 4864 7116 4928
rect 7180 4864 7196 4928
rect 7260 4864 7276 4928
rect 7340 4864 7356 4928
rect 7420 4864 7426 4928
rect 7110 4863 7426 4864
rect 13826 4928 14142 4929
rect 13826 4864 13832 4928
rect 13896 4864 13912 4928
rect 13976 4864 13992 4928
rect 14056 4864 14072 4928
rect 14136 4864 14142 4928
rect 13826 4863 14142 4864
rect 20542 4928 20858 4929
rect 20542 4864 20548 4928
rect 20612 4864 20628 4928
rect 20692 4864 20708 4928
rect 20772 4864 20788 4928
rect 20852 4864 20858 4928
rect 20542 4863 20858 4864
rect 27258 4928 27574 4929
rect 27258 4864 27264 4928
rect 27328 4864 27344 4928
rect 27408 4864 27424 4928
rect 27488 4864 27504 4928
rect 27568 4864 27574 4928
rect 27258 4863 27574 4864
rect 3752 4384 4068 4385
rect 3752 4320 3758 4384
rect 3822 4320 3838 4384
rect 3902 4320 3918 4384
rect 3982 4320 3998 4384
rect 4062 4320 4068 4384
rect 3752 4319 4068 4320
rect 10468 4384 10784 4385
rect 10468 4320 10474 4384
rect 10538 4320 10554 4384
rect 10618 4320 10634 4384
rect 10698 4320 10714 4384
rect 10778 4320 10784 4384
rect 10468 4319 10784 4320
rect 17184 4384 17500 4385
rect 17184 4320 17190 4384
rect 17254 4320 17270 4384
rect 17334 4320 17350 4384
rect 17414 4320 17430 4384
rect 17494 4320 17500 4384
rect 17184 4319 17500 4320
rect 23900 4384 24216 4385
rect 23900 4320 23906 4384
rect 23970 4320 23986 4384
rect 24050 4320 24066 4384
rect 24130 4320 24146 4384
rect 24210 4320 24216 4384
rect 23900 4319 24216 4320
rect 2957 4042 3023 4045
rect 3601 4042 3667 4045
rect 7649 4042 7715 4045
rect 14365 4042 14431 4045
rect 2957 4040 14431 4042
rect 2957 3984 2962 4040
rect 3018 3984 3606 4040
rect 3662 3984 7654 4040
rect 7710 3984 14370 4040
rect 14426 3984 14431 4040
rect 2957 3982 14431 3984
rect 2957 3979 3023 3982
rect 3601 3979 3667 3982
rect 7649 3979 7715 3982
rect 14365 3979 14431 3982
rect 7110 3840 7426 3841
rect 7110 3776 7116 3840
rect 7180 3776 7196 3840
rect 7260 3776 7276 3840
rect 7340 3776 7356 3840
rect 7420 3776 7426 3840
rect 7110 3775 7426 3776
rect 13826 3840 14142 3841
rect 13826 3776 13832 3840
rect 13896 3776 13912 3840
rect 13976 3776 13992 3840
rect 14056 3776 14072 3840
rect 14136 3776 14142 3840
rect 13826 3775 14142 3776
rect 20542 3840 20858 3841
rect 20542 3776 20548 3840
rect 20612 3776 20628 3840
rect 20692 3776 20708 3840
rect 20772 3776 20788 3840
rect 20852 3776 20858 3840
rect 20542 3775 20858 3776
rect 27258 3840 27574 3841
rect 27258 3776 27264 3840
rect 27328 3776 27344 3840
rect 27408 3776 27424 3840
rect 27488 3776 27504 3840
rect 27568 3776 27574 3840
rect 27258 3775 27574 3776
rect 10777 3634 10843 3637
rect 15745 3634 15811 3637
rect 10777 3632 15811 3634
rect 10777 3576 10782 3632
rect 10838 3576 15750 3632
rect 15806 3576 15811 3632
rect 10777 3574 15811 3576
rect 10777 3571 10843 3574
rect 15745 3571 15811 3574
rect 4981 3498 5047 3501
rect 7189 3498 7255 3501
rect 14641 3498 14707 3501
rect 4981 3496 14707 3498
rect 4981 3440 4986 3496
rect 5042 3440 7194 3496
rect 7250 3440 14646 3496
rect 14702 3440 14707 3496
rect 4981 3438 14707 3440
rect 4981 3435 5047 3438
rect 7189 3435 7255 3438
rect 14641 3435 14707 3438
rect 13813 3362 13879 3365
rect 14917 3362 14983 3365
rect 13813 3360 14983 3362
rect 13813 3304 13818 3360
rect 13874 3304 14922 3360
rect 14978 3304 14983 3360
rect 13813 3302 14983 3304
rect 13813 3299 13879 3302
rect 14917 3299 14983 3302
rect 3752 3296 4068 3297
rect 3752 3232 3758 3296
rect 3822 3232 3838 3296
rect 3902 3232 3918 3296
rect 3982 3232 3998 3296
rect 4062 3232 4068 3296
rect 3752 3231 4068 3232
rect 10468 3296 10784 3297
rect 10468 3232 10474 3296
rect 10538 3232 10554 3296
rect 10618 3232 10634 3296
rect 10698 3232 10714 3296
rect 10778 3232 10784 3296
rect 10468 3231 10784 3232
rect 17184 3296 17500 3297
rect 17184 3232 17190 3296
rect 17254 3232 17270 3296
rect 17334 3232 17350 3296
rect 17414 3232 17430 3296
rect 17494 3232 17500 3296
rect 17184 3231 17500 3232
rect 23900 3296 24216 3297
rect 23900 3232 23906 3296
rect 23970 3232 23986 3296
rect 24050 3232 24066 3296
rect 24130 3232 24146 3296
rect 24210 3232 24216 3296
rect 23900 3231 24216 3232
rect 7110 2752 7426 2753
rect 7110 2688 7116 2752
rect 7180 2688 7196 2752
rect 7260 2688 7276 2752
rect 7340 2688 7356 2752
rect 7420 2688 7426 2752
rect 7110 2687 7426 2688
rect 13826 2752 14142 2753
rect 13826 2688 13832 2752
rect 13896 2688 13912 2752
rect 13976 2688 13992 2752
rect 14056 2688 14072 2752
rect 14136 2688 14142 2752
rect 13826 2687 14142 2688
rect 20542 2752 20858 2753
rect 20542 2688 20548 2752
rect 20612 2688 20628 2752
rect 20692 2688 20708 2752
rect 20772 2688 20788 2752
rect 20852 2688 20858 2752
rect 20542 2687 20858 2688
rect 27258 2752 27574 2753
rect 27258 2688 27264 2752
rect 27328 2688 27344 2752
rect 27408 2688 27424 2752
rect 27488 2688 27504 2752
rect 27568 2688 27574 2752
rect 27258 2687 27574 2688
rect 4429 2546 4495 2549
rect 5441 2546 5507 2549
rect 6453 2546 6519 2549
rect 4429 2544 6519 2546
rect 4429 2488 4434 2544
rect 4490 2488 5446 2544
rect 5502 2488 6458 2544
rect 6514 2488 6519 2544
rect 4429 2486 6519 2488
rect 4429 2483 4495 2486
rect 5441 2483 5507 2486
rect 6453 2483 6519 2486
rect 3752 2208 4068 2209
rect 3752 2144 3758 2208
rect 3822 2144 3838 2208
rect 3902 2144 3918 2208
rect 3982 2144 3998 2208
rect 4062 2144 4068 2208
rect 3752 2143 4068 2144
rect 10468 2208 10784 2209
rect 10468 2144 10474 2208
rect 10538 2144 10554 2208
rect 10618 2144 10634 2208
rect 10698 2144 10714 2208
rect 10778 2144 10784 2208
rect 10468 2143 10784 2144
rect 17184 2208 17500 2209
rect 17184 2144 17190 2208
rect 17254 2144 17270 2208
rect 17334 2144 17350 2208
rect 17414 2144 17430 2208
rect 17494 2144 17500 2208
rect 17184 2143 17500 2144
rect 23900 2208 24216 2209
rect 23900 2144 23906 2208
rect 23970 2144 23986 2208
rect 24050 2144 24066 2208
rect 24130 2144 24146 2208
rect 24210 2144 24216 2208
rect 23900 2143 24216 2144
rect 7110 1664 7426 1665
rect 7110 1600 7116 1664
rect 7180 1600 7196 1664
rect 7260 1600 7276 1664
rect 7340 1600 7356 1664
rect 7420 1600 7426 1664
rect 7110 1599 7426 1600
rect 13826 1664 14142 1665
rect 13826 1600 13832 1664
rect 13896 1600 13912 1664
rect 13976 1600 13992 1664
rect 14056 1600 14072 1664
rect 14136 1600 14142 1664
rect 13826 1599 14142 1600
rect 20542 1664 20858 1665
rect 20542 1600 20548 1664
rect 20612 1600 20628 1664
rect 20692 1600 20708 1664
rect 20772 1600 20788 1664
rect 20852 1600 20858 1664
rect 20542 1599 20858 1600
rect 27258 1664 27574 1665
rect 27258 1600 27264 1664
rect 27328 1600 27344 1664
rect 27408 1600 27424 1664
rect 27488 1600 27504 1664
rect 27568 1600 27574 1664
rect 27258 1599 27574 1600
rect 3752 1120 4068 1121
rect 3752 1056 3758 1120
rect 3822 1056 3838 1120
rect 3902 1056 3918 1120
rect 3982 1056 3998 1120
rect 4062 1056 4068 1120
rect 3752 1055 4068 1056
rect 10468 1120 10784 1121
rect 10468 1056 10474 1120
rect 10538 1056 10554 1120
rect 10618 1056 10634 1120
rect 10698 1056 10714 1120
rect 10778 1056 10784 1120
rect 10468 1055 10784 1056
rect 17184 1120 17500 1121
rect 17184 1056 17190 1120
rect 17254 1056 17270 1120
rect 17334 1056 17350 1120
rect 17414 1056 17430 1120
rect 17494 1056 17500 1120
rect 17184 1055 17500 1056
rect 23900 1120 24216 1121
rect 23900 1056 23906 1120
rect 23970 1056 23986 1120
rect 24050 1056 24066 1120
rect 24130 1056 24146 1120
rect 24210 1056 24216 1120
rect 23900 1055 24216 1056
rect 7110 576 7426 577
rect 7110 512 7116 576
rect 7180 512 7196 576
rect 7260 512 7276 576
rect 7340 512 7356 576
rect 7420 512 7426 576
rect 7110 511 7426 512
rect 13826 576 14142 577
rect 13826 512 13832 576
rect 13896 512 13912 576
rect 13976 512 13992 576
rect 14056 512 14072 576
rect 14136 512 14142 576
rect 13826 511 14142 512
rect 20542 576 20858 577
rect 20542 512 20548 576
rect 20612 512 20628 576
rect 20692 512 20708 576
rect 20772 512 20788 576
rect 20852 512 20858 576
rect 20542 511 20858 512
rect 27258 576 27574 577
rect 27258 512 27264 576
rect 27328 512 27344 576
rect 27408 512 27424 576
rect 27488 512 27504 576
rect 27568 512 27574 576
rect 27258 511 27574 512
<< via3 >>
rect 7116 31036 7180 31040
rect 7116 30980 7120 31036
rect 7120 30980 7176 31036
rect 7176 30980 7180 31036
rect 7116 30976 7180 30980
rect 7196 31036 7260 31040
rect 7196 30980 7200 31036
rect 7200 30980 7256 31036
rect 7256 30980 7260 31036
rect 7196 30976 7260 30980
rect 7276 31036 7340 31040
rect 7276 30980 7280 31036
rect 7280 30980 7336 31036
rect 7336 30980 7340 31036
rect 7276 30976 7340 30980
rect 7356 31036 7420 31040
rect 7356 30980 7360 31036
rect 7360 30980 7416 31036
rect 7416 30980 7420 31036
rect 7356 30976 7420 30980
rect 13832 31036 13896 31040
rect 13832 30980 13836 31036
rect 13836 30980 13892 31036
rect 13892 30980 13896 31036
rect 13832 30976 13896 30980
rect 13912 31036 13976 31040
rect 13912 30980 13916 31036
rect 13916 30980 13972 31036
rect 13972 30980 13976 31036
rect 13912 30976 13976 30980
rect 13992 31036 14056 31040
rect 13992 30980 13996 31036
rect 13996 30980 14052 31036
rect 14052 30980 14056 31036
rect 13992 30976 14056 30980
rect 14072 31036 14136 31040
rect 14072 30980 14076 31036
rect 14076 30980 14132 31036
rect 14132 30980 14136 31036
rect 14072 30976 14136 30980
rect 20548 31036 20612 31040
rect 20548 30980 20552 31036
rect 20552 30980 20608 31036
rect 20608 30980 20612 31036
rect 20548 30976 20612 30980
rect 20628 31036 20692 31040
rect 20628 30980 20632 31036
rect 20632 30980 20688 31036
rect 20688 30980 20692 31036
rect 20628 30976 20692 30980
rect 20708 31036 20772 31040
rect 20708 30980 20712 31036
rect 20712 30980 20768 31036
rect 20768 30980 20772 31036
rect 20708 30976 20772 30980
rect 20788 31036 20852 31040
rect 20788 30980 20792 31036
rect 20792 30980 20848 31036
rect 20848 30980 20852 31036
rect 20788 30976 20852 30980
rect 27264 31036 27328 31040
rect 27264 30980 27268 31036
rect 27268 30980 27324 31036
rect 27324 30980 27328 31036
rect 27264 30976 27328 30980
rect 27344 31036 27408 31040
rect 27344 30980 27348 31036
rect 27348 30980 27404 31036
rect 27404 30980 27408 31036
rect 27344 30976 27408 30980
rect 27424 31036 27488 31040
rect 27424 30980 27428 31036
rect 27428 30980 27484 31036
rect 27484 30980 27488 31036
rect 27424 30976 27488 30980
rect 27504 31036 27568 31040
rect 27504 30980 27508 31036
rect 27508 30980 27564 31036
rect 27564 30980 27568 31036
rect 27504 30976 27568 30980
rect 3758 30492 3822 30496
rect 3758 30436 3762 30492
rect 3762 30436 3818 30492
rect 3818 30436 3822 30492
rect 3758 30432 3822 30436
rect 3838 30492 3902 30496
rect 3838 30436 3842 30492
rect 3842 30436 3898 30492
rect 3898 30436 3902 30492
rect 3838 30432 3902 30436
rect 3918 30492 3982 30496
rect 3918 30436 3922 30492
rect 3922 30436 3978 30492
rect 3978 30436 3982 30492
rect 3918 30432 3982 30436
rect 3998 30492 4062 30496
rect 3998 30436 4002 30492
rect 4002 30436 4058 30492
rect 4058 30436 4062 30492
rect 3998 30432 4062 30436
rect 10474 30492 10538 30496
rect 10474 30436 10478 30492
rect 10478 30436 10534 30492
rect 10534 30436 10538 30492
rect 10474 30432 10538 30436
rect 10554 30492 10618 30496
rect 10554 30436 10558 30492
rect 10558 30436 10614 30492
rect 10614 30436 10618 30492
rect 10554 30432 10618 30436
rect 10634 30492 10698 30496
rect 10634 30436 10638 30492
rect 10638 30436 10694 30492
rect 10694 30436 10698 30492
rect 10634 30432 10698 30436
rect 10714 30492 10778 30496
rect 10714 30436 10718 30492
rect 10718 30436 10774 30492
rect 10774 30436 10778 30492
rect 10714 30432 10778 30436
rect 17190 30492 17254 30496
rect 17190 30436 17194 30492
rect 17194 30436 17250 30492
rect 17250 30436 17254 30492
rect 17190 30432 17254 30436
rect 17270 30492 17334 30496
rect 17270 30436 17274 30492
rect 17274 30436 17330 30492
rect 17330 30436 17334 30492
rect 17270 30432 17334 30436
rect 17350 30492 17414 30496
rect 17350 30436 17354 30492
rect 17354 30436 17410 30492
rect 17410 30436 17414 30492
rect 17350 30432 17414 30436
rect 17430 30492 17494 30496
rect 17430 30436 17434 30492
rect 17434 30436 17490 30492
rect 17490 30436 17494 30492
rect 17430 30432 17494 30436
rect 23906 30492 23970 30496
rect 23906 30436 23910 30492
rect 23910 30436 23966 30492
rect 23966 30436 23970 30492
rect 23906 30432 23970 30436
rect 23986 30492 24050 30496
rect 23986 30436 23990 30492
rect 23990 30436 24046 30492
rect 24046 30436 24050 30492
rect 23986 30432 24050 30436
rect 24066 30492 24130 30496
rect 24066 30436 24070 30492
rect 24070 30436 24126 30492
rect 24126 30436 24130 30492
rect 24066 30432 24130 30436
rect 24146 30492 24210 30496
rect 24146 30436 24150 30492
rect 24150 30436 24206 30492
rect 24206 30436 24210 30492
rect 24146 30432 24210 30436
rect 2084 30424 2148 30428
rect 2084 30368 2098 30424
rect 2098 30368 2148 30424
rect 2084 30364 2148 30368
rect 7116 29948 7180 29952
rect 7116 29892 7120 29948
rect 7120 29892 7176 29948
rect 7176 29892 7180 29948
rect 7116 29888 7180 29892
rect 7196 29948 7260 29952
rect 7196 29892 7200 29948
rect 7200 29892 7256 29948
rect 7256 29892 7260 29948
rect 7196 29888 7260 29892
rect 7276 29948 7340 29952
rect 7276 29892 7280 29948
rect 7280 29892 7336 29948
rect 7336 29892 7340 29948
rect 7276 29888 7340 29892
rect 7356 29948 7420 29952
rect 7356 29892 7360 29948
rect 7360 29892 7416 29948
rect 7416 29892 7420 29948
rect 7356 29888 7420 29892
rect 13832 29948 13896 29952
rect 13832 29892 13836 29948
rect 13836 29892 13892 29948
rect 13892 29892 13896 29948
rect 13832 29888 13896 29892
rect 13912 29948 13976 29952
rect 13912 29892 13916 29948
rect 13916 29892 13972 29948
rect 13972 29892 13976 29948
rect 13912 29888 13976 29892
rect 13992 29948 14056 29952
rect 13992 29892 13996 29948
rect 13996 29892 14052 29948
rect 14052 29892 14056 29948
rect 13992 29888 14056 29892
rect 14072 29948 14136 29952
rect 14072 29892 14076 29948
rect 14076 29892 14132 29948
rect 14132 29892 14136 29948
rect 14072 29888 14136 29892
rect 20548 29948 20612 29952
rect 20548 29892 20552 29948
rect 20552 29892 20608 29948
rect 20608 29892 20612 29948
rect 20548 29888 20612 29892
rect 20628 29948 20692 29952
rect 20628 29892 20632 29948
rect 20632 29892 20688 29948
rect 20688 29892 20692 29948
rect 20628 29888 20692 29892
rect 20708 29948 20772 29952
rect 20708 29892 20712 29948
rect 20712 29892 20768 29948
rect 20768 29892 20772 29948
rect 20708 29888 20772 29892
rect 20788 29948 20852 29952
rect 20788 29892 20792 29948
rect 20792 29892 20848 29948
rect 20848 29892 20852 29948
rect 20788 29888 20852 29892
rect 27264 29948 27328 29952
rect 27264 29892 27268 29948
rect 27268 29892 27324 29948
rect 27324 29892 27328 29948
rect 27264 29888 27328 29892
rect 27344 29948 27408 29952
rect 27344 29892 27348 29948
rect 27348 29892 27404 29948
rect 27404 29892 27408 29948
rect 27344 29888 27408 29892
rect 27424 29948 27488 29952
rect 27424 29892 27428 29948
rect 27428 29892 27484 29948
rect 27484 29892 27488 29948
rect 27424 29888 27488 29892
rect 27504 29948 27568 29952
rect 27504 29892 27508 29948
rect 27508 29892 27564 29948
rect 27564 29892 27568 29948
rect 27504 29888 27568 29892
rect 1900 29744 1964 29748
rect 1900 29688 1914 29744
rect 1914 29688 1964 29744
rect 1900 29684 1964 29688
rect 3758 29404 3822 29408
rect 3758 29348 3762 29404
rect 3762 29348 3818 29404
rect 3818 29348 3822 29404
rect 3758 29344 3822 29348
rect 3838 29404 3902 29408
rect 3838 29348 3842 29404
rect 3842 29348 3898 29404
rect 3898 29348 3902 29404
rect 3838 29344 3902 29348
rect 3918 29404 3982 29408
rect 3918 29348 3922 29404
rect 3922 29348 3978 29404
rect 3978 29348 3982 29404
rect 3918 29344 3982 29348
rect 3998 29404 4062 29408
rect 3998 29348 4002 29404
rect 4002 29348 4058 29404
rect 4058 29348 4062 29404
rect 3998 29344 4062 29348
rect 10474 29404 10538 29408
rect 10474 29348 10478 29404
rect 10478 29348 10534 29404
rect 10534 29348 10538 29404
rect 10474 29344 10538 29348
rect 10554 29404 10618 29408
rect 10554 29348 10558 29404
rect 10558 29348 10614 29404
rect 10614 29348 10618 29404
rect 10554 29344 10618 29348
rect 10634 29404 10698 29408
rect 10634 29348 10638 29404
rect 10638 29348 10694 29404
rect 10694 29348 10698 29404
rect 10634 29344 10698 29348
rect 10714 29404 10778 29408
rect 10714 29348 10718 29404
rect 10718 29348 10774 29404
rect 10774 29348 10778 29404
rect 10714 29344 10778 29348
rect 17190 29404 17254 29408
rect 17190 29348 17194 29404
rect 17194 29348 17250 29404
rect 17250 29348 17254 29404
rect 17190 29344 17254 29348
rect 17270 29404 17334 29408
rect 17270 29348 17274 29404
rect 17274 29348 17330 29404
rect 17330 29348 17334 29404
rect 17270 29344 17334 29348
rect 17350 29404 17414 29408
rect 17350 29348 17354 29404
rect 17354 29348 17410 29404
rect 17410 29348 17414 29404
rect 17350 29344 17414 29348
rect 17430 29404 17494 29408
rect 17430 29348 17434 29404
rect 17434 29348 17490 29404
rect 17490 29348 17494 29404
rect 17430 29344 17494 29348
rect 23906 29404 23970 29408
rect 23906 29348 23910 29404
rect 23910 29348 23966 29404
rect 23966 29348 23970 29404
rect 23906 29344 23970 29348
rect 23986 29404 24050 29408
rect 23986 29348 23990 29404
rect 23990 29348 24046 29404
rect 24046 29348 24050 29404
rect 23986 29344 24050 29348
rect 24066 29404 24130 29408
rect 24066 29348 24070 29404
rect 24070 29348 24126 29404
rect 24126 29348 24130 29404
rect 24066 29344 24130 29348
rect 24146 29404 24210 29408
rect 24146 29348 24150 29404
rect 24150 29348 24206 29404
rect 24206 29348 24210 29404
rect 24146 29344 24210 29348
rect 7116 28860 7180 28864
rect 7116 28804 7120 28860
rect 7120 28804 7176 28860
rect 7176 28804 7180 28860
rect 7116 28800 7180 28804
rect 7196 28860 7260 28864
rect 7196 28804 7200 28860
rect 7200 28804 7256 28860
rect 7256 28804 7260 28860
rect 7196 28800 7260 28804
rect 7276 28860 7340 28864
rect 7276 28804 7280 28860
rect 7280 28804 7336 28860
rect 7336 28804 7340 28860
rect 7276 28800 7340 28804
rect 7356 28860 7420 28864
rect 7356 28804 7360 28860
rect 7360 28804 7416 28860
rect 7416 28804 7420 28860
rect 7356 28800 7420 28804
rect 13832 28860 13896 28864
rect 13832 28804 13836 28860
rect 13836 28804 13892 28860
rect 13892 28804 13896 28860
rect 13832 28800 13896 28804
rect 13912 28860 13976 28864
rect 13912 28804 13916 28860
rect 13916 28804 13972 28860
rect 13972 28804 13976 28860
rect 13912 28800 13976 28804
rect 13992 28860 14056 28864
rect 13992 28804 13996 28860
rect 13996 28804 14052 28860
rect 14052 28804 14056 28860
rect 13992 28800 14056 28804
rect 14072 28860 14136 28864
rect 14072 28804 14076 28860
rect 14076 28804 14132 28860
rect 14132 28804 14136 28860
rect 14072 28800 14136 28804
rect 20548 28860 20612 28864
rect 20548 28804 20552 28860
rect 20552 28804 20608 28860
rect 20608 28804 20612 28860
rect 20548 28800 20612 28804
rect 20628 28860 20692 28864
rect 20628 28804 20632 28860
rect 20632 28804 20688 28860
rect 20688 28804 20692 28860
rect 20628 28800 20692 28804
rect 20708 28860 20772 28864
rect 20708 28804 20712 28860
rect 20712 28804 20768 28860
rect 20768 28804 20772 28860
rect 20708 28800 20772 28804
rect 20788 28860 20852 28864
rect 20788 28804 20792 28860
rect 20792 28804 20848 28860
rect 20848 28804 20852 28860
rect 20788 28800 20852 28804
rect 27264 28860 27328 28864
rect 27264 28804 27268 28860
rect 27268 28804 27324 28860
rect 27324 28804 27328 28860
rect 27264 28800 27328 28804
rect 27344 28860 27408 28864
rect 27344 28804 27348 28860
rect 27348 28804 27404 28860
rect 27404 28804 27408 28860
rect 27344 28800 27408 28804
rect 27424 28860 27488 28864
rect 27424 28804 27428 28860
rect 27428 28804 27484 28860
rect 27484 28804 27488 28860
rect 27424 28800 27488 28804
rect 27504 28860 27568 28864
rect 27504 28804 27508 28860
rect 27508 28804 27564 28860
rect 27564 28804 27568 28860
rect 27504 28800 27568 28804
rect 3758 28316 3822 28320
rect 3758 28260 3762 28316
rect 3762 28260 3818 28316
rect 3818 28260 3822 28316
rect 3758 28256 3822 28260
rect 3838 28316 3902 28320
rect 3838 28260 3842 28316
rect 3842 28260 3898 28316
rect 3898 28260 3902 28316
rect 3838 28256 3902 28260
rect 3918 28316 3982 28320
rect 3918 28260 3922 28316
rect 3922 28260 3978 28316
rect 3978 28260 3982 28316
rect 3918 28256 3982 28260
rect 3998 28316 4062 28320
rect 3998 28260 4002 28316
rect 4002 28260 4058 28316
rect 4058 28260 4062 28316
rect 3998 28256 4062 28260
rect 10474 28316 10538 28320
rect 10474 28260 10478 28316
rect 10478 28260 10534 28316
rect 10534 28260 10538 28316
rect 10474 28256 10538 28260
rect 10554 28316 10618 28320
rect 10554 28260 10558 28316
rect 10558 28260 10614 28316
rect 10614 28260 10618 28316
rect 10554 28256 10618 28260
rect 10634 28316 10698 28320
rect 10634 28260 10638 28316
rect 10638 28260 10694 28316
rect 10694 28260 10698 28316
rect 10634 28256 10698 28260
rect 10714 28316 10778 28320
rect 10714 28260 10718 28316
rect 10718 28260 10774 28316
rect 10774 28260 10778 28316
rect 10714 28256 10778 28260
rect 17190 28316 17254 28320
rect 17190 28260 17194 28316
rect 17194 28260 17250 28316
rect 17250 28260 17254 28316
rect 17190 28256 17254 28260
rect 17270 28316 17334 28320
rect 17270 28260 17274 28316
rect 17274 28260 17330 28316
rect 17330 28260 17334 28316
rect 17270 28256 17334 28260
rect 17350 28316 17414 28320
rect 17350 28260 17354 28316
rect 17354 28260 17410 28316
rect 17410 28260 17414 28316
rect 17350 28256 17414 28260
rect 17430 28316 17494 28320
rect 17430 28260 17434 28316
rect 17434 28260 17490 28316
rect 17490 28260 17494 28316
rect 17430 28256 17494 28260
rect 23906 28316 23970 28320
rect 23906 28260 23910 28316
rect 23910 28260 23966 28316
rect 23966 28260 23970 28316
rect 23906 28256 23970 28260
rect 23986 28316 24050 28320
rect 23986 28260 23990 28316
rect 23990 28260 24046 28316
rect 24046 28260 24050 28316
rect 23986 28256 24050 28260
rect 24066 28316 24130 28320
rect 24066 28260 24070 28316
rect 24070 28260 24126 28316
rect 24126 28260 24130 28316
rect 24066 28256 24130 28260
rect 24146 28316 24210 28320
rect 24146 28260 24150 28316
rect 24150 28260 24206 28316
rect 24206 28260 24210 28316
rect 24146 28256 24210 28260
rect 7116 27772 7180 27776
rect 7116 27716 7120 27772
rect 7120 27716 7176 27772
rect 7176 27716 7180 27772
rect 7116 27712 7180 27716
rect 7196 27772 7260 27776
rect 7196 27716 7200 27772
rect 7200 27716 7256 27772
rect 7256 27716 7260 27772
rect 7196 27712 7260 27716
rect 7276 27772 7340 27776
rect 7276 27716 7280 27772
rect 7280 27716 7336 27772
rect 7336 27716 7340 27772
rect 7276 27712 7340 27716
rect 7356 27772 7420 27776
rect 7356 27716 7360 27772
rect 7360 27716 7416 27772
rect 7416 27716 7420 27772
rect 7356 27712 7420 27716
rect 13832 27772 13896 27776
rect 13832 27716 13836 27772
rect 13836 27716 13892 27772
rect 13892 27716 13896 27772
rect 13832 27712 13896 27716
rect 13912 27772 13976 27776
rect 13912 27716 13916 27772
rect 13916 27716 13972 27772
rect 13972 27716 13976 27772
rect 13912 27712 13976 27716
rect 13992 27772 14056 27776
rect 13992 27716 13996 27772
rect 13996 27716 14052 27772
rect 14052 27716 14056 27772
rect 13992 27712 14056 27716
rect 14072 27772 14136 27776
rect 14072 27716 14076 27772
rect 14076 27716 14132 27772
rect 14132 27716 14136 27772
rect 14072 27712 14136 27716
rect 20548 27772 20612 27776
rect 20548 27716 20552 27772
rect 20552 27716 20608 27772
rect 20608 27716 20612 27772
rect 20548 27712 20612 27716
rect 20628 27772 20692 27776
rect 20628 27716 20632 27772
rect 20632 27716 20688 27772
rect 20688 27716 20692 27772
rect 20628 27712 20692 27716
rect 20708 27772 20772 27776
rect 20708 27716 20712 27772
rect 20712 27716 20768 27772
rect 20768 27716 20772 27772
rect 20708 27712 20772 27716
rect 20788 27772 20852 27776
rect 20788 27716 20792 27772
rect 20792 27716 20848 27772
rect 20848 27716 20852 27772
rect 20788 27712 20852 27716
rect 27264 27772 27328 27776
rect 27264 27716 27268 27772
rect 27268 27716 27324 27772
rect 27324 27716 27328 27772
rect 27264 27712 27328 27716
rect 27344 27772 27408 27776
rect 27344 27716 27348 27772
rect 27348 27716 27404 27772
rect 27404 27716 27408 27772
rect 27344 27712 27408 27716
rect 27424 27772 27488 27776
rect 27424 27716 27428 27772
rect 27428 27716 27484 27772
rect 27484 27716 27488 27772
rect 27424 27712 27488 27716
rect 27504 27772 27568 27776
rect 27504 27716 27508 27772
rect 27508 27716 27564 27772
rect 27564 27716 27568 27772
rect 27504 27712 27568 27716
rect 24900 27704 24964 27708
rect 24900 27648 24950 27704
rect 24950 27648 24964 27704
rect 24900 27644 24964 27648
rect 3758 27228 3822 27232
rect 3758 27172 3762 27228
rect 3762 27172 3818 27228
rect 3818 27172 3822 27228
rect 3758 27168 3822 27172
rect 3838 27228 3902 27232
rect 3838 27172 3842 27228
rect 3842 27172 3898 27228
rect 3898 27172 3902 27228
rect 3838 27168 3902 27172
rect 3918 27228 3982 27232
rect 3918 27172 3922 27228
rect 3922 27172 3978 27228
rect 3978 27172 3982 27228
rect 3918 27168 3982 27172
rect 3998 27228 4062 27232
rect 3998 27172 4002 27228
rect 4002 27172 4058 27228
rect 4058 27172 4062 27228
rect 3998 27168 4062 27172
rect 10474 27228 10538 27232
rect 10474 27172 10478 27228
rect 10478 27172 10534 27228
rect 10534 27172 10538 27228
rect 10474 27168 10538 27172
rect 10554 27228 10618 27232
rect 10554 27172 10558 27228
rect 10558 27172 10614 27228
rect 10614 27172 10618 27228
rect 10554 27168 10618 27172
rect 10634 27228 10698 27232
rect 10634 27172 10638 27228
rect 10638 27172 10694 27228
rect 10694 27172 10698 27228
rect 10634 27168 10698 27172
rect 10714 27228 10778 27232
rect 10714 27172 10718 27228
rect 10718 27172 10774 27228
rect 10774 27172 10778 27228
rect 10714 27168 10778 27172
rect 17190 27228 17254 27232
rect 17190 27172 17194 27228
rect 17194 27172 17250 27228
rect 17250 27172 17254 27228
rect 17190 27168 17254 27172
rect 17270 27228 17334 27232
rect 17270 27172 17274 27228
rect 17274 27172 17330 27228
rect 17330 27172 17334 27228
rect 17270 27168 17334 27172
rect 17350 27228 17414 27232
rect 17350 27172 17354 27228
rect 17354 27172 17410 27228
rect 17410 27172 17414 27228
rect 17350 27168 17414 27172
rect 17430 27228 17494 27232
rect 17430 27172 17434 27228
rect 17434 27172 17490 27228
rect 17490 27172 17494 27228
rect 17430 27168 17494 27172
rect 23906 27228 23970 27232
rect 23906 27172 23910 27228
rect 23910 27172 23966 27228
rect 23966 27172 23970 27228
rect 23906 27168 23970 27172
rect 23986 27228 24050 27232
rect 23986 27172 23990 27228
rect 23990 27172 24046 27228
rect 24046 27172 24050 27228
rect 23986 27168 24050 27172
rect 24066 27228 24130 27232
rect 24066 27172 24070 27228
rect 24070 27172 24126 27228
rect 24126 27172 24130 27228
rect 24066 27168 24130 27172
rect 24146 27228 24210 27232
rect 24146 27172 24150 27228
rect 24150 27172 24206 27228
rect 24206 27172 24210 27228
rect 24146 27168 24210 27172
rect 7116 26684 7180 26688
rect 7116 26628 7120 26684
rect 7120 26628 7176 26684
rect 7176 26628 7180 26684
rect 7116 26624 7180 26628
rect 7196 26684 7260 26688
rect 7196 26628 7200 26684
rect 7200 26628 7256 26684
rect 7256 26628 7260 26684
rect 7196 26624 7260 26628
rect 7276 26684 7340 26688
rect 7276 26628 7280 26684
rect 7280 26628 7336 26684
rect 7336 26628 7340 26684
rect 7276 26624 7340 26628
rect 7356 26684 7420 26688
rect 7356 26628 7360 26684
rect 7360 26628 7416 26684
rect 7416 26628 7420 26684
rect 7356 26624 7420 26628
rect 13832 26684 13896 26688
rect 13832 26628 13836 26684
rect 13836 26628 13892 26684
rect 13892 26628 13896 26684
rect 13832 26624 13896 26628
rect 13912 26684 13976 26688
rect 13912 26628 13916 26684
rect 13916 26628 13972 26684
rect 13972 26628 13976 26684
rect 13912 26624 13976 26628
rect 13992 26684 14056 26688
rect 13992 26628 13996 26684
rect 13996 26628 14052 26684
rect 14052 26628 14056 26684
rect 13992 26624 14056 26628
rect 14072 26684 14136 26688
rect 14072 26628 14076 26684
rect 14076 26628 14132 26684
rect 14132 26628 14136 26684
rect 14072 26624 14136 26628
rect 20548 26684 20612 26688
rect 20548 26628 20552 26684
rect 20552 26628 20608 26684
rect 20608 26628 20612 26684
rect 20548 26624 20612 26628
rect 20628 26684 20692 26688
rect 20628 26628 20632 26684
rect 20632 26628 20688 26684
rect 20688 26628 20692 26684
rect 20628 26624 20692 26628
rect 20708 26684 20772 26688
rect 20708 26628 20712 26684
rect 20712 26628 20768 26684
rect 20768 26628 20772 26684
rect 20708 26624 20772 26628
rect 20788 26684 20852 26688
rect 20788 26628 20792 26684
rect 20792 26628 20848 26684
rect 20848 26628 20852 26684
rect 20788 26624 20852 26628
rect 27264 26684 27328 26688
rect 27264 26628 27268 26684
rect 27268 26628 27324 26684
rect 27324 26628 27328 26684
rect 27264 26624 27328 26628
rect 27344 26684 27408 26688
rect 27344 26628 27348 26684
rect 27348 26628 27404 26684
rect 27404 26628 27408 26684
rect 27344 26624 27408 26628
rect 27424 26684 27488 26688
rect 27424 26628 27428 26684
rect 27428 26628 27484 26684
rect 27484 26628 27488 26684
rect 27424 26624 27488 26628
rect 27504 26684 27568 26688
rect 27504 26628 27508 26684
rect 27508 26628 27564 26684
rect 27564 26628 27568 26684
rect 27504 26624 27568 26628
rect 3758 26140 3822 26144
rect 3758 26084 3762 26140
rect 3762 26084 3818 26140
rect 3818 26084 3822 26140
rect 3758 26080 3822 26084
rect 3838 26140 3902 26144
rect 3838 26084 3842 26140
rect 3842 26084 3898 26140
rect 3898 26084 3902 26140
rect 3838 26080 3902 26084
rect 3918 26140 3982 26144
rect 3918 26084 3922 26140
rect 3922 26084 3978 26140
rect 3978 26084 3982 26140
rect 3918 26080 3982 26084
rect 3998 26140 4062 26144
rect 3998 26084 4002 26140
rect 4002 26084 4058 26140
rect 4058 26084 4062 26140
rect 3998 26080 4062 26084
rect 10474 26140 10538 26144
rect 10474 26084 10478 26140
rect 10478 26084 10534 26140
rect 10534 26084 10538 26140
rect 10474 26080 10538 26084
rect 10554 26140 10618 26144
rect 10554 26084 10558 26140
rect 10558 26084 10614 26140
rect 10614 26084 10618 26140
rect 10554 26080 10618 26084
rect 10634 26140 10698 26144
rect 10634 26084 10638 26140
rect 10638 26084 10694 26140
rect 10694 26084 10698 26140
rect 10634 26080 10698 26084
rect 10714 26140 10778 26144
rect 10714 26084 10718 26140
rect 10718 26084 10774 26140
rect 10774 26084 10778 26140
rect 10714 26080 10778 26084
rect 17190 26140 17254 26144
rect 17190 26084 17194 26140
rect 17194 26084 17250 26140
rect 17250 26084 17254 26140
rect 17190 26080 17254 26084
rect 17270 26140 17334 26144
rect 17270 26084 17274 26140
rect 17274 26084 17330 26140
rect 17330 26084 17334 26140
rect 17270 26080 17334 26084
rect 17350 26140 17414 26144
rect 17350 26084 17354 26140
rect 17354 26084 17410 26140
rect 17410 26084 17414 26140
rect 17350 26080 17414 26084
rect 17430 26140 17494 26144
rect 17430 26084 17434 26140
rect 17434 26084 17490 26140
rect 17490 26084 17494 26140
rect 17430 26080 17494 26084
rect 23906 26140 23970 26144
rect 23906 26084 23910 26140
rect 23910 26084 23966 26140
rect 23966 26084 23970 26140
rect 23906 26080 23970 26084
rect 23986 26140 24050 26144
rect 23986 26084 23990 26140
rect 23990 26084 24046 26140
rect 24046 26084 24050 26140
rect 23986 26080 24050 26084
rect 24066 26140 24130 26144
rect 24066 26084 24070 26140
rect 24070 26084 24126 26140
rect 24126 26084 24130 26140
rect 24066 26080 24130 26084
rect 24146 26140 24210 26144
rect 24146 26084 24150 26140
rect 24150 26084 24206 26140
rect 24206 26084 24210 26140
rect 24146 26080 24210 26084
rect 7116 25596 7180 25600
rect 7116 25540 7120 25596
rect 7120 25540 7176 25596
rect 7176 25540 7180 25596
rect 7116 25536 7180 25540
rect 7196 25596 7260 25600
rect 7196 25540 7200 25596
rect 7200 25540 7256 25596
rect 7256 25540 7260 25596
rect 7196 25536 7260 25540
rect 7276 25596 7340 25600
rect 7276 25540 7280 25596
rect 7280 25540 7336 25596
rect 7336 25540 7340 25596
rect 7276 25536 7340 25540
rect 7356 25596 7420 25600
rect 7356 25540 7360 25596
rect 7360 25540 7416 25596
rect 7416 25540 7420 25596
rect 7356 25536 7420 25540
rect 13832 25596 13896 25600
rect 13832 25540 13836 25596
rect 13836 25540 13892 25596
rect 13892 25540 13896 25596
rect 13832 25536 13896 25540
rect 13912 25596 13976 25600
rect 13912 25540 13916 25596
rect 13916 25540 13972 25596
rect 13972 25540 13976 25596
rect 13912 25536 13976 25540
rect 13992 25596 14056 25600
rect 13992 25540 13996 25596
rect 13996 25540 14052 25596
rect 14052 25540 14056 25596
rect 13992 25536 14056 25540
rect 14072 25596 14136 25600
rect 14072 25540 14076 25596
rect 14076 25540 14132 25596
rect 14132 25540 14136 25596
rect 14072 25536 14136 25540
rect 20548 25596 20612 25600
rect 20548 25540 20552 25596
rect 20552 25540 20608 25596
rect 20608 25540 20612 25596
rect 20548 25536 20612 25540
rect 20628 25596 20692 25600
rect 20628 25540 20632 25596
rect 20632 25540 20688 25596
rect 20688 25540 20692 25596
rect 20628 25536 20692 25540
rect 20708 25596 20772 25600
rect 20708 25540 20712 25596
rect 20712 25540 20768 25596
rect 20768 25540 20772 25596
rect 20708 25536 20772 25540
rect 20788 25596 20852 25600
rect 20788 25540 20792 25596
rect 20792 25540 20848 25596
rect 20848 25540 20852 25596
rect 20788 25536 20852 25540
rect 27264 25596 27328 25600
rect 27264 25540 27268 25596
rect 27268 25540 27324 25596
rect 27324 25540 27328 25596
rect 27264 25536 27328 25540
rect 27344 25596 27408 25600
rect 27344 25540 27348 25596
rect 27348 25540 27404 25596
rect 27404 25540 27408 25596
rect 27344 25536 27408 25540
rect 27424 25596 27488 25600
rect 27424 25540 27428 25596
rect 27428 25540 27484 25596
rect 27484 25540 27488 25596
rect 27424 25536 27488 25540
rect 27504 25596 27568 25600
rect 27504 25540 27508 25596
rect 27508 25540 27564 25596
rect 27564 25540 27568 25596
rect 27504 25536 27568 25540
rect 3758 25052 3822 25056
rect 3758 24996 3762 25052
rect 3762 24996 3818 25052
rect 3818 24996 3822 25052
rect 3758 24992 3822 24996
rect 3838 25052 3902 25056
rect 3838 24996 3842 25052
rect 3842 24996 3898 25052
rect 3898 24996 3902 25052
rect 3838 24992 3902 24996
rect 3918 25052 3982 25056
rect 3918 24996 3922 25052
rect 3922 24996 3978 25052
rect 3978 24996 3982 25052
rect 3918 24992 3982 24996
rect 3998 25052 4062 25056
rect 3998 24996 4002 25052
rect 4002 24996 4058 25052
rect 4058 24996 4062 25052
rect 3998 24992 4062 24996
rect 10474 25052 10538 25056
rect 10474 24996 10478 25052
rect 10478 24996 10534 25052
rect 10534 24996 10538 25052
rect 10474 24992 10538 24996
rect 10554 25052 10618 25056
rect 10554 24996 10558 25052
rect 10558 24996 10614 25052
rect 10614 24996 10618 25052
rect 10554 24992 10618 24996
rect 10634 25052 10698 25056
rect 10634 24996 10638 25052
rect 10638 24996 10694 25052
rect 10694 24996 10698 25052
rect 10634 24992 10698 24996
rect 10714 25052 10778 25056
rect 10714 24996 10718 25052
rect 10718 24996 10774 25052
rect 10774 24996 10778 25052
rect 10714 24992 10778 24996
rect 17190 25052 17254 25056
rect 17190 24996 17194 25052
rect 17194 24996 17250 25052
rect 17250 24996 17254 25052
rect 17190 24992 17254 24996
rect 17270 25052 17334 25056
rect 17270 24996 17274 25052
rect 17274 24996 17330 25052
rect 17330 24996 17334 25052
rect 17270 24992 17334 24996
rect 17350 25052 17414 25056
rect 17350 24996 17354 25052
rect 17354 24996 17410 25052
rect 17410 24996 17414 25052
rect 17350 24992 17414 24996
rect 17430 25052 17494 25056
rect 17430 24996 17434 25052
rect 17434 24996 17490 25052
rect 17490 24996 17494 25052
rect 17430 24992 17494 24996
rect 23906 25052 23970 25056
rect 23906 24996 23910 25052
rect 23910 24996 23966 25052
rect 23966 24996 23970 25052
rect 23906 24992 23970 24996
rect 23986 25052 24050 25056
rect 23986 24996 23990 25052
rect 23990 24996 24046 25052
rect 24046 24996 24050 25052
rect 23986 24992 24050 24996
rect 24066 25052 24130 25056
rect 24066 24996 24070 25052
rect 24070 24996 24126 25052
rect 24126 24996 24130 25052
rect 24066 24992 24130 24996
rect 24146 25052 24210 25056
rect 24146 24996 24150 25052
rect 24150 24996 24206 25052
rect 24206 24996 24210 25052
rect 24146 24992 24210 24996
rect 7116 24508 7180 24512
rect 7116 24452 7120 24508
rect 7120 24452 7176 24508
rect 7176 24452 7180 24508
rect 7116 24448 7180 24452
rect 7196 24508 7260 24512
rect 7196 24452 7200 24508
rect 7200 24452 7256 24508
rect 7256 24452 7260 24508
rect 7196 24448 7260 24452
rect 7276 24508 7340 24512
rect 7276 24452 7280 24508
rect 7280 24452 7336 24508
rect 7336 24452 7340 24508
rect 7276 24448 7340 24452
rect 7356 24508 7420 24512
rect 7356 24452 7360 24508
rect 7360 24452 7416 24508
rect 7416 24452 7420 24508
rect 7356 24448 7420 24452
rect 13832 24508 13896 24512
rect 13832 24452 13836 24508
rect 13836 24452 13892 24508
rect 13892 24452 13896 24508
rect 13832 24448 13896 24452
rect 13912 24508 13976 24512
rect 13912 24452 13916 24508
rect 13916 24452 13972 24508
rect 13972 24452 13976 24508
rect 13912 24448 13976 24452
rect 13992 24508 14056 24512
rect 13992 24452 13996 24508
rect 13996 24452 14052 24508
rect 14052 24452 14056 24508
rect 13992 24448 14056 24452
rect 14072 24508 14136 24512
rect 14072 24452 14076 24508
rect 14076 24452 14132 24508
rect 14132 24452 14136 24508
rect 14072 24448 14136 24452
rect 20548 24508 20612 24512
rect 20548 24452 20552 24508
rect 20552 24452 20608 24508
rect 20608 24452 20612 24508
rect 20548 24448 20612 24452
rect 20628 24508 20692 24512
rect 20628 24452 20632 24508
rect 20632 24452 20688 24508
rect 20688 24452 20692 24508
rect 20628 24448 20692 24452
rect 20708 24508 20772 24512
rect 20708 24452 20712 24508
rect 20712 24452 20768 24508
rect 20768 24452 20772 24508
rect 20708 24448 20772 24452
rect 20788 24508 20852 24512
rect 20788 24452 20792 24508
rect 20792 24452 20848 24508
rect 20848 24452 20852 24508
rect 20788 24448 20852 24452
rect 27264 24508 27328 24512
rect 27264 24452 27268 24508
rect 27268 24452 27324 24508
rect 27324 24452 27328 24508
rect 27264 24448 27328 24452
rect 27344 24508 27408 24512
rect 27344 24452 27348 24508
rect 27348 24452 27404 24508
rect 27404 24452 27408 24508
rect 27344 24448 27408 24452
rect 27424 24508 27488 24512
rect 27424 24452 27428 24508
rect 27428 24452 27484 24508
rect 27484 24452 27488 24508
rect 27424 24448 27488 24452
rect 27504 24508 27568 24512
rect 27504 24452 27508 24508
rect 27508 24452 27564 24508
rect 27564 24452 27568 24508
rect 27504 24448 27568 24452
rect 3758 23964 3822 23968
rect 3758 23908 3762 23964
rect 3762 23908 3818 23964
rect 3818 23908 3822 23964
rect 3758 23904 3822 23908
rect 3838 23964 3902 23968
rect 3838 23908 3842 23964
rect 3842 23908 3898 23964
rect 3898 23908 3902 23964
rect 3838 23904 3902 23908
rect 3918 23964 3982 23968
rect 3918 23908 3922 23964
rect 3922 23908 3978 23964
rect 3978 23908 3982 23964
rect 3918 23904 3982 23908
rect 3998 23964 4062 23968
rect 3998 23908 4002 23964
rect 4002 23908 4058 23964
rect 4058 23908 4062 23964
rect 3998 23904 4062 23908
rect 10474 23964 10538 23968
rect 10474 23908 10478 23964
rect 10478 23908 10534 23964
rect 10534 23908 10538 23964
rect 10474 23904 10538 23908
rect 10554 23964 10618 23968
rect 10554 23908 10558 23964
rect 10558 23908 10614 23964
rect 10614 23908 10618 23964
rect 10554 23904 10618 23908
rect 10634 23964 10698 23968
rect 10634 23908 10638 23964
rect 10638 23908 10694 23964
rect 10694 23908 10698 23964
rect 10634 23904 10698 23908
rect 10714 23964 10778 23968
rect 10714 23908 10718 23964
rect 10718 23908 10774 23964
rect 10774 23908 10778 23964
rect 10714 23904 10778 23908
rect 17190 23964 17254 23968
rect 17190 23908 17194 23964
rect 17194 23908 17250 23964
rect 17250 23908 17254 23964
rect 17190 23904 17254 23908
rect 17270 23964 17334 23968
rect 17270 23908 17274 23964
rect 17274 23908 17330 23964
rect 17330 23908 17334 23964
rect 17270 23904 17334 23908
rect 17350 23964 17414 23968
rect 17350 23908 17354 23964
rect 17354 23908 17410 23964
rect 17410 23908 17414 23964
rect 17350 23904 17414 23908
rect 17430 23964 17494 23968
rect 17430 23908 17434 23964
rect 17434 23908 17490 23964
rect 17490 23908 17494 23964
rect 17430 23904 17494 23908
rect 23906 23964 23970 23968
rect 23906 23908 23910 23964
rect 23910 23908 23966 23964
rect 23966 23908 23970 23964
rect 23906 23904 23970 23908
rect 23986 23964 24050 23968
rect 23986 23908 23990 23964
rect 23990 23908 24046 23964
rect 24046 23908 24050 23964
rect 23986 23904 24050 23908
rect 24066 23964 24130 23968
rect 24066 23908 24070 23964
rect 24070 23908 24126 23964
rect 24126 23908 24130 23964
rect 24066 23904 24130 23908
rect 24146 23964 24210 23968
rect 24146 23908 24150 23964
rect 24150 23908 24206 23964
rect 24206 23908 24210 23964
rect 24146 23904 24210 23908
rect 7116 23420 7180 23424
rect 7116 23364 7120 23420
rect 7120 23364 7176 23420
rect 7176 23364 7180 23420
rect 7116 23360 7180 23364
rect 7196 23420 7260 23424
rect 7196 23364 7200 23420
rect 7200 23364 7256 23420
rect 7256 23364 7260 23420
rect 7196 23360 7260 23364
rect 7276 23420 7340 23424
rect 7276 23364 7280 23420
rect 7280 23364 7336 23420
rect 7336 23364 7340 23420
rect 7276 23360 7340 23364
rect 7356 23420 7420 23424
rect 7356 23364 7360 23420
rect 7360 23364 7416 23420
rect 7416 23364 7420 23420
rect 7356 23360 7420 23364
rect 13832 23420 13896 23424
rect 13832 23364 13836 23420
rect 13836 23364 13892 23420
rect 13892 23364 13896 23420
rect 13832 23360 13896 23364
rect 13912 23420 13976 23424
rect 13912 23364 13916 23420
rect 13916 23364 13972 23420
rect 13972 23364 13976 23420
rect 13912 23360 13976 23364
rect 13992 23420 14056 23424
rect 13992 23364 13996 23420
rect 13996 23364 14052 23420
rect 14052 23364 14056 23420
rect 13992 23360 14056 23364
rect 14072 23420 14136 23424
rect 14072 23364 14076 23420
rect 14076 23364 14132 23420
rect 14132 23364 14136 23420
rect 14072 23360 14136 23364
rect 20548 23420 20612 23424
rect 20548 23364 20552 23420
rect 20552 23364 20608 23420
rect 20608 23364 20612 23420
rect 20548 23360 20612 23364
rect 20628 23420 20692 23424
rect 20628 23364 20632 23420
rect 20632 23364 20688 23420
rect 20688 23364 20692 23420
rect 20628 23360 20692 23364
rect 20708 23420 20772 23424
rect 20708 23364 20712 23420
rect 20712 23364 20768 23420
rect 20768 23364 20772 23420
rect 20708 23360 20772 23364
rect 20788 23420 20852 23424
rect 20788 23364 20792 23420
rect 20792 23364 20848 23420
rect 20848 23364 20852 23420
rect 20788 23360 20852 23364
rect 27264 23420 27328 23424
rect 27264 23364 27268 23420
rect 27268 23364 27324 23420
rect 27324 23364 27328 23420
rect 27264 23360 27328 23364
rect 27344 23420 27408 23424
rect 27344 23364 27348 23420
rect 27348 23364 27404 23420
rect 27404 23364 27408 23420
rect 27344 23360 27408 23364
rect 27424 23420 27488 23424
rect 27424 23364 27428 23420
rect 27428 23364 27484 23420
rect 27484 23364 27488 23420
rect 27424 23360 27488 23364
rect 27504 23420 27568 23424
rect 27504 23364 27508 23420
rect 27508 23364 27564 23420
rect 27564 23364 27568 23420
rect 27504 23360 27568 23364
rect 3758 22876 3822 22880
rect 3758 22820 3762 22876
rect 3762 22820 3818 22876
rect 3818 22820 3822 22876
rect 3758 22816 3822 22820
rect 3838 22876 3902 22880
rect 3838 22820 3842 22876
rect 3842 22820 3898 22876
rect 3898 22820 3902 22876
rect 3838 22816 3902 22820
rect 3918 22876 3982 22880
rect 3918 22820 3922 22876
rect 3922 22820 3978 22876
rect 3978 22820 3982 22876
rect 3918 22816 3982 22820
rect 3998 22876 4062 22880
rect 3998 22820 4002 22876
rect 4002 22820 4058 22876
rect 4058 22820 4062 22876
rect 3998 22816 4062 22820
rect 10474 22876 10538 22880
rect 10474 22820 10478 22876
rect 10478 22820 10534 22876
rect 10534 22820 10538 22876
rect 10474 22816 10538 22820
rect 10554 22876 10618 22880
rect 10554 22820 10558 22876
rect 10558 22820 10614 22876
rect 10614 22820 10618 22876
rect 10554 22816 10618 22820
rect 10634 22876 10698 22880
rect 10634 22820 10638 22876
rect 10638 22820 10694 22876
rect 10694 22820 10698 22876
rect 10634 22816 10698 22820
rect 10714 22876 10778 22880
rect 10714 22820 10718 22876
rect 10718 22820 10774 22876
rect 10774 22820 10778 22876
rect 10714 22816 10778 22820
rect 17190 22876 17254 22880
rect 17190 22820 17194 22876
rect 17194 22820 17250 22876
rect 17250 22820 17254 22876
rect 17190 22816 17254 22820
rect 17270 22876 17334 22880
rect 17270 22820 17274 22876
rect 17274 22820 17330 22876
rect 17330 22820 17334 22876
rect 17270 22816 17334 22820
rect 17350 22876 17414 22880
rect 17350 22820 17354 22876
rect 17354 22820 17410 22876
rect 17410 22820 17414 22876
rect 17350 22816 17414 22820
rect 17430 22876 17494 22880
rect 17430 22820 17434 22876
rect 17434 22820 17490 22876
rect 17490 22820 17494 22876
rect 17430 22816 17494 22820
rect 23906 22876 23970 22880
rect 23906 22820 23910 22876
rect 23910 22820 23966 22876
rect 23966 22820 23970 22876
rect 23906 22816 23970 22820
rect 23986 22876 24050 22880
rect 23986 22820 23990 22876
rect 23990 22820 24046 22876
rect 24046 22820 24050 22876
rect 23986 22816 24050 22820
rect 24066 22876 24130 22880
rect 24066 22820 24070 22876
rect 24070 22820 24126 22876
rect 24126 22820 24130 22876
rect 24066 22816 24130 22820
rect 24146 22876 24210 22880
rect 24146 22820 24150 22876
rect 24150 22820 24206 22876
rect 24206 22820 24210 22876
rect 24146 22816 24210 22820
rect 7116 22332 7180 22336
rect 7116 22276 7120 22332
rect 7120 22276 7176 22332
rect 7176 22276 7180 22332
rect 7116 22272 7180 22276
rect 7196 22332 7260 22336
rect 7196 22276 7200 22332
rect 7200 22276 7256 22332
rect 7256 22276 7260 22332
rect 7196 22272 7260 22276
rect 7276 22332 7340 22336
rect 7276 22276 7280 22332
rect 7280 22276 7336 22332
rect 7336 22276 7340 22332
rect 7276 22272 7340 22276
rect 7356 22332 7420 22336
rect 7356 22276 7360 22332
rect 7360 22276 7416 22332
rect 7416 22276 7420 22332
rect 7356 22272 7420 22276
rect 13832 22332 13896 22336
rect 13832 22276 13836 22332
rect 13836 22276 13892 22332
rect 13892 22276 13896 22332
rect 13832 22272 13896 22276
rect 13912 22332 13976 22336
rect 13912 22276 13916 22332
rect 13916 22276 13972 22332
rect 13972 22276 13976 22332
rect 13912 22272 13976 22276
rect 13992 22332 14056 22336
rect 13992 22276 13996 22332
rect 13996 22276 14052 22332
rect 14052 22276 14056 22332
rect 13992 22272 14056 22276
rect 14072 22332 14136 22336
rect 14072 22276 14076 22332
rect 14076 22276 14132 22332
rect 14132 22276 14136 22332
rect 14072 22272 14136 22276
rect 20548 22332 20612 22336
rect 20548 22276 20552 22332
rect 20552 22276 20608 22332
rect 20608 22276 20612 22332
rect 20548 22272 20612 22276
rect 20628 22332 20692 22336
rect 20628 22276 20632 22332
rect 20632 22276 20688 22332
rect 20688 22276 20692 22332
rect 20628 22272 20692 22276
rect 20708 22332 20772 22336
rect 20708 22276 20712 22332
rect 20712 22276 20768 22332
rect 20768 22276 20772 22332
rect 20708 22272 20772 22276
rect 20788 22332 20852 22336
rect 20788 22276 20792 22332
rect 20792 22276 20848 22332
rect 20848 22276 20852 22332
rect 20788 22272 20852 22276
rect 27264 22332 27328 22336
rect 27264 22276 27268 22332
rect 27268 22276 27324 22332
rect 27324 22276 27328 22332
rect 27264 22272 27328 22276
rect 27344 22332 27408 22336
rect 27344 22276 27348 22332
rect 27348 22276 27404 22332
rect 27404 22276 27408 22332
rect 27344 22272 27408 22276
rect 27424 22332 27488 22336
rect 27424 22276 27428 22332
rect 27428 22276 27484 22332
rect 27484 22276 27488 22332
rect 27424 22272 27488 22276
rect 27504 22332 27568 22336
rect 27504 22276 27508 22332
rect 27508 22276 27564 22332
rect 27564 22276 27568 22332
rect 27504 22272 27568 22276
rect 3758 21788 3822 21792
rect 3758 21732 3762 21788
rect 3762 21732 3818 21788
rect 3818 21732 3822 21788
rect 3758 21728 3822 21732
rect 3838 21788 3902 21792
rect 3838 21732 3842 21788
rect 3842 21732 3898 21788
rect 3898 21732 3902 21788
rect 3838 21728 3902 21732
rect 3918 21788 3982 21792
rect 3918 21732 3922 21788
rect 3922 21732 3978 21788
rect 3978 21732 3982 21788
rect 3918 21728 3982 21732
rect 3998 21788 4062 21792
rect 3998 21732 4002 21788
rect 4002 21732 4058 21788
rect 4058 21732 4062 21788
rect 3998 21728 4062 21732
rect 10474 21788 10538 21792
rect 10474 21732 10478 21788
rect 10478 21732 10534 21788
rect 10534 21732 10538 21788
rect 10474 21728 10538 21732
rect 10554 21788 10618 21792
rect 10554 21732 10558 21788
rect 10558 21732 10614 21788
rect 10614 21732 10618 21788
rect 10554 21728 10618 21732
rect 10634 21788 10698 21792
rect 10634 21732 10638 21788
rect 10638 21732 10694 21788
rect 10694 21732 10698 21788
rect 10634 21728 10698 21732
rect 10714 21788 10778 21792
rect 10714 21732 10718 21788
rect 10718 21732 10774 21788
rect 10774 21732 10778 21788
rect 10714 21728 10778 21732
rect 17190 21788 17254 21792
rect 17190 21732 17194 21788
rect 17194 21732 17250 21788
rect 17250 21732 17254 21788
rect 17190 21728 17254 21732
rect 17270 21788 17334 21792
rect 17270 21732 17274 21788
rect 17274 21732 17330 21788
rect 17330 21732 17334 21788
rect 17270 21728 17334 21732
rect 17350 21788 17414 21792
rect 17350 21732 17354 21788
rect 17354 21732 17410 21788
rect 17410 21732 17414 21788
rect 17350 21728 17414 21732
rect 17430 21788 17494 21792
rect 17430 21732 17434 21788
rect 17434 21732 17490 21788
rect 17490 21732 17494 21788
rect 17430 21728 17494 21732
rect 23906 21788 23970 21792
rect 23906 21732 23910 21788
rect 23910 21732 23966 21788
rect 23966 21732 23970 21788
rect 23906 21728 23970 21732
rect 23986 21788 24050 21792
rect 23986 21732 23990 21788
rect 23990 21732 24046 21788
rect 24046 21732 24050 21788
rect 23986 21728 24050 21732
rect 24066 21788 24130 21792
rect 24066 21732 24070 21788
rect 24070 21732 24126 21788
rect 24126 21732 24130 21788
rect 24066 21728 24130 21732
rect 24146 21788 24210 21792
rect 24146 21732 24150 21788
rect 24150 21732 24206 21788
rect 24206 21732 24210 21788
rect 24146 21728 24210 21732
rect 7116 21244 7180 21248
rect 7116 21188 7120 21244
rect 7120 21188 7176 21244
rect 7176 21188 7180 21244
rect 7116 21184 7180 21188
rect 7196 21244 7260 21248
rect 7196 21188 7200 21244
rect 7200 21188 7256 21244
rect 7256 21188 7260 21244
rect 7196 21184 7260 21188
rect 7276 21244 7340 21248
rect 7276 21188 7280 21244
rect 7280 21188 7336 21244
rect 7336 21188 7340 21244
rect 7276 21184 7340 21188
rect 7356 21244 7420 21248
rect 7356 21188 7360 21244
rect 7360 21188 7416 21244
rect 7416 21188 7420 21244
rect 7356 21184 7420 21188
rect 13832 21244 13896 21248
rect 13832 21188 13836 21244
rect 13836 21188 13892 21244
rect 13892 21188 13896 21244
rect 13832 21184 13896 21188
rect 13912 21244 13976 21248
rect 13912 21188 13916 21244
rect 13916 21188 13972 21244
rect 13972 21188 13976 21244
rect 13912 21184 13976 21188
rect 13992 21244 14056 21248
rect 13992 21188 13996 21244
rect 13996 21188 14052 21244
rect 14052 21188 14056 21244
rect 13992 21184 14056 21188
rect 14072 21244 14136 21248
rect 14072 21188 14076 21244
rect 14076 21188 14132 21244
rect 14132 21188 14136 21244
rect 14072 21184 14136 21188
rect 20548 21244 20612 21248
rect 20548 21188 20552 21244
rect 20552 21188 20608 21244
rect 20608 21188 20612 21244
rect 20548 21184 20612 21188
rect 20628 21244 20692 21248
rect 20628 21188 20632 21244
rect 20632 21188 20688 21244
rect 20688 21188 20692 21244
rect 20628 21184 20692 21188
rect 20708 21244 20772 21248
rect 20708 21188 20712 21244
rect 20712 21188 20768 21244
rect 20768 21188 20772 21244
rect 20708 21184 20772 21188
rect 20788 21244 20852 21248
rect 20788 21188 20792 21244
rect 20792 21188 20848 21244
rect 20848 21188 20852 21244
rect 20788 21184 20852 21188
rect 27264 21244 27328 21248
rect 27264 21188 27268 21244
rect 27268 21188 27324 21244
rect 27324 21188 27328 21244
rect 27264 21184 27328 21188
rect 27344 21244 27408 21248
rect 27344 21188 27348 21244
rect 27348 21188 27404 21244
rect 27404 21188 27408 21244
rect 27344 21184 27408 21188
rect 27424 21244 27488 21248
rect 27424 21188 27428 21244
rect 27428 21188 27484 21244
rect 27484 21188 27488 21244
rect 27424 21184 27488 21188
rect 27504 21244 27568 21248
rect 27504 21188 27508 21244
rect 27508 21188 27564 21244
rect 27564 21188 27568 21244
rect 27504 21184 27568 21188
rect 3758 20700 3822 20704
rect 3758 20644 3762 20700
rect 3762 20644 3818 20700
rect 3818 20644 3822 20700
rect 3758 20640 3822 20644
rect 3838 20700 3902 20704
rect 3838 20644 3842 20700
rect 3842 20644 3898 20700
rect 3898 20644 3902 20700
rect 3838 20640 3902 20644
rect 3918 20700 3982 20704
rect 3918 20644 3922 20700
rect 3922 20644 3978 20700
rect 3978 20644 3982 20700
rect 3918 20640 3982 20644
rect 3998 20700 4062 20704
rect 3998 20644 4002 20700
rect 4002 20644 4058 20700
rect 4058 20644 4062 20700
rect 3998 20640 4062 20644
rect 10474 20700 10538 20704
rect 10474 20644 10478 20700
rect 10478 20644 10534 20700
rect 10534 20644 10538 20700
rect 10474 20640 10538 20644
rect 10554 20700 10618 20704
rect 10554 20644 10558 20700
rect 10558 20644 10614 20700
rect 10614 20644 10618 20700
rect 10554 20640 10618 20644
rect 10634 20700 10698 20704
rect 10634 20644 10638 20700
rect 10638 20644 10694 20700
rect 10694 20644 10698 20700
rect 10634 20640 10698 20644
rect 10714 20700 10778 20704
rect 10714 20644 10718 20700
rect 10718 20644 10774 20700
rect 10774 20644 10778 20700
rect 10714 20640 10778 20644
rect 17190 20700 17254 20704
rect 17190 20644 17194 20700
rect 17194 20644 17250 20700
rect 17250 20644 17254 20700
rect 17190 20640 17254 20644
rect 17270 20700 17334 20704
rect 17270 20644 17274 20700
rect 17274 20644 17330 20700
rect 17330 20644 17334 20700
rect 17270 20640 17334 20644
rect 17350 20700 17414 20704
rect 17350 20644 17354 20700
rect 17354 20644 17410 20700
rect 17410 20644 17414 20700
rect 17350 20640 17414 20644
rect 17430 20700 17494 20704
rect 17430 20644 17434 20700
rect 17434 20644 17490 20700
rect 17490 20644 17494 20700
rect 17430 20640 17494 20644
rect 23906 20700 23970 20704
rect 23906 20644 23910 20700
rect 23910 20644 23966 20700
rect 23966 20644 23970 20700
rect 23906 20640 23970 20644
rect 23986 20700 24050 20704
rect 23986 20644 23990 20700
rect 23990 20644 24046 20700
rect 24046 20644 24050 20700
rect 23986 20640 24050 20644
rect 24066 20700 24130 20704
rect 24066 20644 24070 20700
rect 24070 20644 24126 20700
rect 24126 20644 24130 20700
rect 24066 20640 24130 20644
rect 24146 20700 24210 20704
rect 24146 20644 24150 20700
rect 24150 20644 24206 20700
rect 24206 20644 24210 20700
rect 24146 20640 24210 20644
rect 7116 20156 7180 20160
rect 7116 20100 7120 20156
rect 7120 20100 7176 20156
rect 7176 20100 7180 20156
rect 7116 20096 7180 20100
rect 7196 20156 7260 20160
rect 7196 20100 7200 20156
rect 7200 20100 7256 20156
rect 7256 20100 7260 20156
rect 7196 20096 7260 20100
rect 7276 20156 7340 20160
rect 7276 20100 7280 20156
rect 7280 20100 7336 20156
rect 7336 20100 7340 20156
rect 7276 20096 7340 20100
rect 7356 20156 7420 20160
rect 7356 20100 7360 20156
rect 7360 20100 7416 20156
rect 7416 20100 7420 20156
rect 7356 20096 7420 20100
rect 13832 20156 13896 20160
rect 13832 20100 13836 20156
rect 13836 20100 13892 20156
rect 13892 20100 13896 20156
rect 13832 20096 13896 20100
rect 13912 20156 13976 20160
rect 13912 20100 13916 20156
rect 13916 20100 13972 20156
rect 13972 20100 13976 20156
rect 13912 20096 13976 20100
rect 13992 20156 14056 20160
rect 13992 20100 13996 20156
rect 13996 20100 14052 20156
rect 14052 20100 14056 20156
rect 13992 20096 14056 20100
rect 14072 20156 14136 20160
rect 14072 20100 14076 20156
rect 14076 20100 14132 20156
rect 14132 20100 14136 20156
rect 14072 20096 14136 20100
rect 20548 20156 20612 20160
rect 20548 20100 20552 20156
rect 20552 20100 20608 20156
rect 20608 20100 20612 20156
rect 20548 20096 20612 20100
rect 20628 20156 20692 20160
rect 20628 20100 20632 20156
rect 20632 20100 20688 20156
rect 20688 20100 20692 20156
rect 20628 20096 20692 20100
rect 20708 20156 20772 20160
rect 20708 20100 20712 20156
rect 20712 20100 20768 20156
rect 20768 20100 20772 20156
rect 20708 20096 20772 20100
rect 20788 20156 20852 20160
rect 20788 20100 20792 20156
rect 20792 20100 20848 20156
rect 20848 20100 20852 20156
rect 20788 20096 20852 20100
rect 27264 20156 27328 20160
rect 27264 20100 27268 20156
rect 27268 20100 27324 20156
rect 27324 20100 27328 20156
rect 27264 20096 27328 20100
rect 27344 20156 27408 20160
rect 27344 20100 27348 20156
rect 27348 20100 27404 20156
rect 27404 20100 27408 20156
rect 27344 20096 27408 20100
rect 27424 20156 27488 20160
rect 27424 20100 27428 20156
rect 27428 20100 27484 20156
rect 27484 20100 27488 20156
rect 27424 20096 27488 20100
rect 27504 20156 27568 20160
rect 27504 20100 27508 20156
rect 27508 20100 27564 20156
rect 27564 20100 27568 20156
rect 27504 20096 27568 20100
rect 3758 19612 3822 19616
rect 3758 19556 3762 19612
rect 3762 19556 3818 19612
rect 3818 19556 3822 19612
rect 3758 19552 3822 19556
rect 3838 19612 3902 19616
rect 3838 19556 3842 19612
rect 3842 19556 3898 19612
rect 3898 19556 3902 19612
rect 3838 19552 3902 19556
rect 3918 19612 3982 19616
rect 3918 19556 3922 19612
rect 3922 19556 3978 19612
rect 3978 19556 3982 19612
rect 3918 19552 3982 19556
rect 3998 19612 4062 19616
rect 3998 19556 4002 19612
rect 4002 19556 4058 19612
rect 4058 19556 4062 19612
rect 3998 19552 4062 19556
rect 10474 19612 10538 19616
rect 10474 19556 10478 19612
rect 10478 19556 10534 19612
rect 10534 19556 10538 19612
rect 10474 19552 10538 19556
rect 10554 19612 10618 19616
rect 10554 19556 10558 19612
rect 10558 19556 10614 19612
rect 10614 19556 10618 19612
rect 10554 19552 10618 19556
rect 10634 19612 10698 19616
rect 10634 19556 10638 19612
rect 10638 19556 10694 19612
rect 10694 19556 10698 19612
rect 10634 19552 10698 19556
rect 10714 19612 10778 19616
rect 10714 19556 10718 19612
rect 10718 19556 10774 19612
rect 10774 19556 10778 19612
rect 10714 19552 10778 19556
rect 17190 19612 17254 19616
rect 17190 19556 17194 19612
rect 17194 19556 17250 19612
rect 17250 19556 17254 19612
rect 17190 19552 17254 19556
rect 17270 19612 17334 19616
rect 17270 19556 17274 19612
rect 17274 19556 17330 19612
rect 17330 19556 17334 19612
rect 17270 19552 17334 19556
rect 17350 19612 17414 19616
rect 17350 19556 17354 19612
rect 17354 19556 17410 19612
rect 17410 19556 17414 19612
rect 17350 19552 17414 19556
rect 17430 19612 17494 19616
rect 17430 19556 17434 19612
rect 17434 19556 17490 19612
rect 17490 19556 17494 19612
rect 17430 19552 17494 19556
rect 23906 19612 23970 19616
rect 23906 19556 23910 19612
rect 23910 19556 23966 19612
rect 23966 19556 23970 19612
rect 23906 19552 23970 19556
rect 23986 19612 24050 19616
rect 23986 19556 23990 19612
rect 23990 19556 24046 19612
rect 24046 19556 24050 19612
rect 23986 19552 24050 19556
rect 24066 19612 24130 19616
rect 24066 19556 24070 19612
rect 24070 19556 24126 19612
rect 24126 19556 24130 19612
rect 24066 19552 24130 19556
rect 24146 19612 24210 19616
rect 24146 19556 24150 19612
rect 24150 19556 24206 19612
rect 24206 19556 24210 19612
rect 24146 19552 24210 19556
rect 7116 19068 7180 19072
rect 7116 19012 7120 19068
rect 7120 19012 7176 19068
rect 7176 19012 7180 19068
rect 7116 19008 7180 19012
rect 7196 19068 7260 19072
rect 7196 19012 7200 19068
rect 7200 19012 7256 19068
rect 7256 19012 7260 19068
rect 7196 19008 7260 19012
rect 7276 19068 7340 19072
rect 7276 19012 7280 19068
rect 7280 19012 7336 19068
rect 7336 19012 7340 19068
rect 7276 19008 7340 19012
rect 7356 19068 7420 19072
rect 7356 19012 7360 19068
rect 7360 19012 7416 19068
rect 7416 19012 7420 19068
rect 7356 19008 7420 19012
rect 13832 19068 13896 19072
rect 13832 19012 13836 19068
rect 13836 19012 13892 19068
rect 13892 19012 13896 19068
rect 13832 19008 13896 19012
rect 13912 19068 13976 19072
rect 13912 19012 13916 19068
rect 13916 19012 13972 19068
rect 13972 19012 13976 19068
rect 13912 19008 13976 19012
rect 13992 19068 14056 19072
rect 13992 19012 13996 19068
rect 13996 19012 14052 19068
rect 14052 19012 14056 19068
rect 13992 19008 14056 19012
rect 14072 19068 14136 19072
rect 14072 19012 14076 19068
rect 14076 19012 14132 19068
rect 14132 19012 14136 19068
rect 14072 19008 14136 19012
rect 20548 19068 20612 19072
rect 20548 19012 20552 19068
rect 20552 19012 20608 19068
rect 20608 19012 20612 19068
rect 20548 19008 20612 19012
rect 20628 19068 20692 19072
rect 20628 19012 20632 19068
rect 20632 19012 20688 19068
rect 20688 19012 20692 19068
rect 20628 19008 20692 19012
rect 20708 19068 20772 19072
rect 20708 19012 20712 19068
rect 20712 19012 20768 19068
rect 20768 19012 20772 19068
rect 20708 19008 20772 19012
rect 20788 19068 20852 19072
rect 20788 19012 20792 19068
rect 20792 19012 20848 19068
rect 20848 19012 20852 19068
rect 20788 19008 20852 19012
rect 27264 19068 27328 19072
rect 27264 19012 27268 19068
rect 27268 19012 27324 19068
rect 27324 19012 27328 19068
rect 27264 19008 27328 19012
rect 27344 19068 27408 19072
rect 27344 19012 27348 19068
rect 27348 19012 27404 19068
rect 27404 19012 27408 19068
rect 27344 19008 27408 19012
rect 27424 19068 27488 19072
rect 27424 19012 27428 19068
rect 27428 19012 27484 19068
rect 27484 19012 27488 19068
rect 27424 19008 27488 19012
rect 27504 19068 27568 19072
rect 27504 19012 27508 19068
rect 27508 19012 27564 19068
rect 27564 19012 27568 19068
rect 27504 19008 27568 19012
rect 3758 18524 3822 18528
rect 3758 18468 3762 18524
rect 3762 18468 3818 18524
rect 3818 18468 3822 18524
rect 3758 18464 3822 18468
rect 3838 18524 3902 18528
rect 3838 18468 3842 18524
rect 3842 18468 3898 18524
rect 3898 18468 3902 18524
rect 3838 18464 3902 18468
rect 3918 18524 3982 18528
rect 3918 18468 3922 18524
rect 3922 18468 3978 18524
rect 3978 18468 3982 18524
rect 3918 18464 3982 18468
rect 3998 18524 4062 18528
rect 3998 18468 4002 18524
rect 4002 18468 4058 18524
rect 4058 18468 4062 18524
rect 3998 18464 4062 18468
rect 10474 18524 10538 18528
rect 10474 18468 10478 18524
rect 10478 18468 10534 18524
rect 10534 18468 10538 18524
rect 10474 18464 10538 18468
rect 10554 18524 10618 18528
rect 10554 18468 10558 18524
rect 10558 18468 10614 18524
rect 10614 18468 10618 18524
rect 10554 18464 10618 18468
rect 10634 18524 10698 18528
rect 10634 18468 10638 18524
rect 10638 18468 10694 18524
rect 10694 18468 10698 18524
rect 10634 18464 10698 18468
rect 10714 18524 10778 18528
rect 10714 18468 10718 18524
rect 10718 18468 10774 18524
rect 10774 18468 10778 18524
rect 10714 18464 10778 18468
rect 17190 18524 17254 18528
rect 17190 18468 17194 18524
rect 17194 18468 17250 18524
rect 17250 18468 17254 18524
rect 17190 18464 17254 18468
rect 17270 18524 17334 18528
rect 17270 18468 17274 18524
rect 17274 18468 17330 18524
rect 17330 18468 17334 18524
rect 17270 18464 17334 18468
rect 17350 18524 17414 18528
rect 17350 18468 17354 18524
rect 17354 18468 17410 18524
rect 17410 18468 17414 18524
rect 17350 18464 17414 18468
rect 17430 18524 17494 18528
rect 17430 18468 17434 18524
rect 17434 18468 17490 18524
rect 17490 18468 17494 18524
rect 17430 18464 17494 18468
rect 23906 18524 23970 18528
rect 23906 18468 23910 18524
rect 23910 18468 23966 18524
rect 23966 18468 23970 18524
rect 23906 18464 23970 18468
rect 23986 18524 24050 18528
rect 23986 18468 23990 18524
rect 23990 18468 24046 18524
rect 24046 18468 24050 18524
rect 23986 18464 24050 18468
rect 24066 18524 24130 18528
rect 24066 18468 24070 18524
rect 24070 18468 24126 18524
rect 24126 18468 24130 18524
rect 24066 18464 24130 18468
rect 24146 18524 24210 18528
rect 24146 18468 24150 18524
rect 24150 18468 24206 18524
rect 24206 18468 24210 18524
rect 24146 18464 24210 18468
rect 7116 17980 7180 17984
rect 7116 17924 7120 17980
rect 7120 17924 7176 17980
rect 7176 17924 7180 17980
rect 7116 17920 7180 17924
rect 7196 17980 7260 17984
rect 7196 17924 7200 17980
rect 7200 17924 7256 17980
rect 7256 17924 7260 17980
rect 7196 17920 7260 17924
rect 7276 17980 7340 17984
rect 7276 17924 7280 17980
rect 7280 17924 7336 17980
rect 7336 17924 7340 17980
rect 7276 17920 7340 17924
rect 7356 17980 7420 17984
rect 7356 17924 7360 17980
rect 7360 17924 7416 17980
rect 7416 17924 7420 17980
rect 7356 17920 7420 17924
rect 13832 17980 13896 17984
rect 13832 17924 13836 17980
rect 13836 17924 13892 17980
rect 13892 17924 13896 17980
rect 13832 17920 13896 17924
rect 13912 17980 13976 17984
rect 13912 17924 13916 17980
rect 13916 17924 13972 17980
rect 13972 17924 13976 17980
rect 13912 17920 13976 17924
rect 13992 17980 14056 17984
rect 13992 17924 13996 17980
rect 13996 17924 14052 17980
rect 14052 17924 14056 17980
rect 13992 17920 14056 17924
rect 14072 17980 14136 17984
rect 14072 17924 14076 17980
rect 14076 17924 14132 17980
rect 14132 17924 14136 17980
rect 14072 17920 14136 17924
rect 20548 17980 20612 17984
rect 20548 17924 20552 17980
rect 20552 17924 20608 17980
rect 20608 17924 20612 17980
rect 20548 17920 20612 17924
rect 20628 17980 20692 17984
rect 20628 17924 20632 17980
rect 20632 17924 20688 17980
rect 20688 17924 20692 17980
rect 20628 17920 20692 17924
rect 20708 17980 20772 17984
rect 20708 17924 20712 17980
rect 20712 17924 20768 17980
rect 20768 17924 20772 17980
rect 20708 17920 20772 17924
rect 20788 17980 20852 17984
rect 20788 17924 20792 17980
rect 20792 17924 20848 17980
rect 20848 17924 20852 17980
rect 20788 17920 20852 17924
rect 27264 17980 27328 17984
rect 27264 17924 27268 17980
rect 27268 17924 27324 17980
rect 27324 17924 27328 17980
rect 27264 17920 27328 17924
rect 27344 17980 27408 17984
rect 27344 17924 27348 17980
rect 27348 17924 27404 17980
rect 27404 17924 27408 17980
rect 27344 17920 27408 17924
rect 27424 17980 27488 17984
rect 27424 17924 27428 17980
rect 27428 17924 27484 17980
rect 27484 17924 27488 17980
rect 27424 17920 27488 17924
rect 27504 17980 27568 17984
rect 27504 17924 27508 17980
rect 27508 17924 27564 17980
rect 27564 17924 27568 17980
rect 27504 17920 27568 17924
rect 3758 17436 3822 17440
rect 3758 17380 3762 17436
rect 3762 17380 3818 17436
rect 3818 17380 3822 17436
rect 3758 17376 3822 17380
rect 3838 17436 3902 17440
rect 3838 17380 3842 17436
rect 3842 17380 3898 17436
rect 3898 17380 3902 17436
rect 3838 17376 3902 17380
rect 3918 17436 3982 17440
rect 3918 17380 3922 17436
rect 3922 17380 3978 17436
rect 3978 17380 3982 17436
rect 3918 17376 3982 17380
rect 3998 17436 4062 17440
rect 3998 17380 4002 17436
rect 4002 17380 4058 17436
rect 4058 17380 4062 17436
rect 3998 17376 4062 17380
rect 10474 17436 10538 17440
rect 10474 17380 10478 17436
rect 10478 17380 10534 17436
rect 10534 17380 10538 17436
rect 10474 17376 10538 17380
rect 10554 17436 10618 17440
rect 10554 17380 10558 17436
rect 10558 17380 10614 17436
rect 10614 17380 10618 17436
rect 10554 17376 10618 17380
rect 10634 17436 10698 17440
rect 10634 17380 10638 17436
rect 10638 17380 10694 17436
rect 10694 17380 10698 17436
rect 10634 17376 10698 17380
rect 10714 17436 10778 17440
rect 10714 17380 10718 17436
rect 10718 17380 10774 17436
rect 10774 17380 10778 17436
rect 10714 17376 10778 17380
rect 17190 17436 17254 17440
rect 17190 17380 17194 17436
rect 17194 17380 17250 17436
rect 17250 17380 17254 17436
rect 17190 17376 17254 17380
rect 17270 17436 17334 17440
rect 17270 17380 17274 17436
rect 17274 17380 17330 17436
rect 17330 17380 17334 17436
rect 17270 17376 17334 17380
rect 17350 17436 17414 17440
rect 17350 17380 17354 17436
rect 17354 17380 17410 17436
rect 17410 17380 17414 17436
rect 17350 17376 17414 17380
rect 17430 17436 17494 17440
rect 17430 17380 17434 17436
rect 17434 17380 17490 17436
rect 17490 17380 17494 17436
rect 17430 17376 17494 17380
rect 23906 17436 23970 17440
rect 23906 17380 23910 17436
rect 23910 17380 23966 17436
rect 23966 17380 23970 17436
rect 23906 17376 23970 17380
rect 23986 17436 24050 17440
rect 23986 17380 23990 17436
rect 23990 17380 24046 17436
rect 24046 17380 24050 17436
rect 23986 17376 24050 17380
rect 24066 17436 24130 17440
rect 24066 17380 24070 17436
rect 24070 17380 24126 17436
rect 24126 17380 24130 17436
rect 24066 17376 24130 17380
rect 24146 17436 24210 17440
rect 24146 17380 24150 17436
rect 24150 17380 24206 17436
rect 24206 17380 24210 17436
rect 24146 17376 24210 17380
rect 24900 17036 24964 17100
rect 7116 16892 7180 16896
rect 7116 16836 7120 16892
rect 7120 16836 7176 16892
rect 7176 16836 7180 16892
rect 7116 16832 7180 16836
rect 7196 16892 7260 16896
rect 7196 16836 7200 16892
rect 7200 16836 7256 16892
rect 7256 16836 7260 16892
rect 7196 16832 7260 16836
rect 7276 16892 7340 16896
rect 7276 16836 7280 16892
rect 7280 16836 7336 16892
rect 7336 16836 7340 16892
rect 7276 16832 7340 16836
rect 7356 16892 7420 16896
rect 7356 16836 7360 16892
rect 7360 16836 7416 16892
rect 7416 16836 7420 16892
rect 7356 16832 7420 16836
rect 13832 16892 13896 16896
rect 13832 16836 13836 16892
rect 13836 16836 13892 16892
rect 13892 16836 13896 16892
rect 13832 16832 13896 16836
rect 13912 16892 13976 16896
rect 13912 16836 13916 16892
rect 13916 16836 13972 16892
rect 13972 16836 13976 16892
rect 13912 16832 13976 16836
rect 13992 16892 14056 16896
rect 13992 16836 13996 16892
rect 13996 16836 14052 16892
rect 14052 16836 14056 16892
rect 13992 16832 14056 16836
rect 14072 16892 14136 16896
rect 14072 16836 14076 16892
rect 14076 16836 14132 16892
rect 14132 16836 14136 16892
rect 14072 16832 14136 16836
rect 20548 16892 20612 16896
rect 20548 16836 20552 16892
rect 20552 16836 20608 16892
rect 20608 16836 20612 16892
rect 20548 16832 20612 16836
rect 20628 16892 20692 16896
rect 20628 16836 20632 16892
rect 20632 16836 20688 16892
rect 20688 16836 20692 16892
rect 20628 16832 20692 16836
rect 20708 16892 20772 16896
rect 20708 16836 20712 16892
rect 20712 16836 20768 16892
rect 20768 16836 20772 16892
rect 20708 16832 20772 16836
rect 20788 16892 20852 16896
rect 20788 16836 20792 16892
rect 20792 16836 20848 16892
rect 20848 16836 20852 16892
rect 20788 16832 20852 16836
rect 27264 16892 27328 16896
rect 27264 16836 27268 16892
rect 27268 16836 27324 16892
rect 27324 16836 27328 16892
rect 27264 16832 27328 16836
rect 27344 16892 27408 16896
rect 27344 16836 27348 16892
rect 27348 16836 27404 16892
rect 27404 16836 27408 16892
rect 27344 16832 27408 16836
rect 27424 16892 27488 16896
rect 27424 16836 27428 16892
rect 27428 16836 27484 16892
rect 27484 16836 27488 16892
rect 27424 16832 27488 16836
rect 27504 16892 27568 16896
rect 27504 16836 27508 16892
rect 27508 16836 27564 16892
rect 27564 16836 27568 16892
rect 27504 16832 27568 16836
rect 3758 16348 3822 16352
rect 3758 16292 3762 16348
rect 3762 16292 3818 16348
rect 3818 16292 3822 16348
rect 3758 16288 3822 16292
rect 3838 16348 3902 16352
rect 3838 16292 3842 16348
rect 3842 16292 3898 16348
rect 3898 16292 3902 16348
rect 3838 16288 3902 16292
rect 3918 16348 3982 16352
rect 3918 16292 3922 16348
rect 3922 16292 3978 16348
rect 3978 16292 3982 16348
rect 3918 16288 3982 16292
rect 3998 16348 4062 16352
rect 3998 16292 4002 16348
rect 4002 16292 4058 16348
rect 4058 16292 4062 16348
rect 3998 16288 4062 16292
rect 10474 16348 10538 16352
rect 10474 16292 10478 16348
rect 10478 16292 10534 16348
rect 10534 16292 10538 16348
rect 10474 16288 10538 16292
rect 10554 16348 10618 16352
rect 10554 16292 10558 16348
rect 10558 16292 10614 16348
rect 10614 16292 10618 16348
rect 10554 16288 10618 16292
rect 10634 16348 10698 16352
rect 10634 16292 10638 16348
rect 10638 16292 10694 16348
rect 10694 16292 10698 16348
rect 10634 16288 10698 16292
rect 10714 16348 10778 16352
rect 10714 16292 10718 16348
rect 10718 16292 10774 16348
rect 10774 16292 10778 16348
rect 10714 16288 10778 16292
rect 17190 16348 17254 16352
rect 17190 16292 17194 16348
rect 17194 16292 17250 16348
rect 17250 16292 17254 16348
rect 17190 16288 17254 16292
rect 17270 16348 17334 16352
rect 17270 16292 17274 16348
rect 17274 16292 17330 16348
rect 17330 16292 17334 16348
rect 17270 16288 17334 16292
rect 17350 16348 17414 16352
rect 17350 16292 17354 16348
rect 17354 16292 17410 16348
rect 17410 16292 17414 16348
rect 17350 16288 17414 16292
rect 17430 16348 17494 16352
rect 17430 16292 17434 16348
rect 17434 16292 17490 16348
rect 17490 16292 17494 16348
rect 17430 16288 17494 16292
rect 23906 16348 23970 16352
rect 23906 16292 23910 16348
rect 23910 16292 23966 16348
rect 23966 16292 23970 16348
rect 23906 16288 23970 16292
rect 23986 16348 24050 16352
rect 23986 16292 23990 16348
rect 23990 16292 24046 16348
rect 24046 16292 24050 16348
rect 23986 16288 24050 16292
rect 24066 16348 24130 16352
rect 24066 16292 24070 16348
rect 24070 16292 24126 16348
rect 24126 16292 24130 16348
rect 24066 16288 24130 16292
rect 24146 16348 24210 16352
rect 24146 16292 24150 16348
rect 24150 16292 24206 16348
rect 24206 16292 24210 16348
rect 24146 16288 24210 16292
rect 7116 15804 7180 15808
rect 7116 15748 7120 15804
rect 7120 15748 7176 15804
rect 7176 15748 7180 15804
rect 7116 15744 7180 15748
rect 7196 15804 7260 15808
rect 7196 15748 7200 15804
rect 7200 15748 7256 15804
rect 7256 15748 7260 15804
rect 7196 15744 7260 15748
rect 7276 15804 7340 15808
rect 7276 15748 7280 15804
rect 7280 15748 7336 15804
rect 7336 15748 7340 15804
rect 7276 15744 7340 15748
rect 7356 15804 7420 15808
rect 7356 15748 7360 15804
rect 7360 15748 7416 15804
rect 7416 15748 7420 15804
rect 7356 15744 7420 15748
rect 13832 15804 13896 15808
rect 13832 15748 13836 15804
rect 13836 15748 13892 15804
rect 13892 15748 13896 15804
rect 13832 15744 13896 15748
rect 13912 15804 13976 15808
rect 13912 15748 13916 15804
rect 13916 15748 13972 15804
rect 13972 15748 13976 15804
rect 13912 15744 13976 15748
rect 13992 15804 14056 15808
rect 13992 15748 13996 15804
rect 13996 15748 14052 15804
rect 14052 15748 14056 15804
rect 13992 15744 14056 15748
rect 14072 15804 14136 15808
rect 14072 15748 14076 15804
rect 14076 15748 14132 15804
rect 14132 15748 14136 15804
rect 14072 15744 14136 15748
rect 20548 15804 20612 15808
rect 20548 15748 20552 15804
rect 20552 15748 20608 15804
rect 20608 15748 20612 15804
rect 20548 15744 20612 15748
rect 20628 15804 20692 15808
rect 20628 15748 20632 15804
rect 20632 15748 20688 15804
rect 20688 15748 20692 15804
rect 20628 15744 20692 15748
rect 20708 15804 20772 15808
rect 20708 15748 20712 15804
rect 20712 15748 20768 15804
rect 20768 15748 20772 15804
rect 20708 15744 20772 15748
rect 20788 15804 20852 15808
rect 20788 15748 20792 15804
rect 20792 15748 20848 15804
rect 20848 15748 20852 15804
rect 20788 15744 20852 15748
rect 27264 15804 27328 15808
rect 27264 15748 27268 15804
rect 27268 15748 27324 15804
rect 27324 15748 27328 15804
rect 27264 15744 27328 15748
rect 27344 15804 27408 15808
rect 27344 15748 27348 15804
rect 27348 15748 27404 15804
rect 27404 15748 27408 15804
rect 27344 15744 27408 15748
rect 27424 15804 27488 15808
rect 27424 15748 27428 15804
rect 27428 15748 27484 15804
rect 27484 15748 27488 15804
rect 27424 15744 27488 15748
rect 27504 15804 27568 15808
rect 27504 15748 27508 15804
rect 27508 15748 27564 15804
rect 27564 15748 27568 15804
rect 27504 15744 27568 15748
rect 3758 15260 3822 15264
rect 3758 15204 3762 15260
rect 3762 15204 3818 15260
rect 3818 15204 3822 15260
rect 3758 15200 3822 15204
rect 3838 15260 3902 15264
rect 3838 15204 3842 15260
rect 3842 15204 3898 15260
rect 3898 15204 3902 15260
rect 3838 15200 3902 15204
rect 3918 15260 3982 15264
rect 3918 15204 3922 15260
rect 3922 15204 3978 15260
rect 3978 15204 3982 15260
rect 3918 15200 3982 15204
rect 3998 15260 4062 15264
rect 3998 15204 4002 15260
rect 4002 15204 4058 15260
rect 4058 15204 4062 15260
rect 3998 15200 4062 15204
rect 10474 15260 10538 15264
rect 10474 15204 10478 15260
rect 10478 15204 10534 15260
rect 10534 15204 10538 15260
rect 10474 15200 10538 15204
rect 10554 15260 10618 15264
rect 10554 15204 10558 15260
rect 10558 15204 10614 15260
rect 10614 15204 10618 15260
rect 10554 15200 10618 15204
rect 10634 15260 10698 15264
rect 10634 15204 10638 15260
rect 10638 15204 10694 15260
rect 10694 15204 10698 15260
rect 10634 15200 10698 15204
rect 10714 15260 10778 15264
rect 10714 15204 10718 15260
rect 10718 15204 10774 15260
rect 10774 15204 10778 15260
rect 10714 15200 10778 15204
rect 17190 15260 17254 15264
rect 17190 15204 17194 15260
rect 17194 15204 17250 15260
rect 17250 15204 17254 15260
rect 17190 15200 17254 15204
rect 17270 15260 17334 15264
rect 17270 15204 17274 15260
rect 17274 15204 17330 15260
rect 17330 15204 17334 15260
rect 17270 15200 17334 15204
rect 17350 15260 17414 15264
rect 17350 15204 17354 15260
rect 17354 15204 17410 15260
rect 17410 15204 17414 15260
rect 17350 15200 17414 15204
rect 17430 15260 17494 15264
rect 17430 15204 17434 15260
rect 17434 15204 17490 15260
rect 17490 15204 17494 15260
rect 17430 15200 17494 15204
rect 23906 15260 23970 15264
rect 23906 15204 23910 15260
rect 23910 15204 23966 15260
rect 23966 15204 23970 15260
rect 23906 15200 23970 15204
rect 23986 15260 24050 15264
rect 23986 15204 23990 15260
rect 23990 15204 24046 15260
rect 24046 15204 24050 15260
rect 23986 15200 24050 15204
rect 24066 15260 24130 15264
rect 24066 15204 24070 15260
rect 24070 15204 24126 15260
rect 24126 15204 24130 15260
rect 24066 15200 24130 15204
rect 24146 15260 24210 15264
rect 24146 15204 24150 15260
rect 24150 15204 24206 15260
rect 24206 15204 24210 15260
rect 24146 15200 24210 15204
rect 7116 14716 7180 14720
rect 7116 14660 7120 14716
rect 7120 14660 7176 14716
rect 7176 14660 7180 14716
rect 7116 14656 7180 14660
rect 7196 14716 7260 14720
rect 7196 14660 7200 14716
rect 7200 14660 7256 14716
rect 7256 14660 7260 14716
rect 7196 14656 7260 14660
rect 7276 14716 7340 14720
rect 7276 14660 7280 14716
rect 7280 14660 7336 14716
rect 7336 14660 7340 14716
rect 7276 14656 7340 14660
rect 7356 14716 7420 14720
rect 7356 14660 7360 14716
rect 7360 14660 7416 14716
rect 7416 14660 7420 14716
rect 7356 14656 7420 14660
rect 13832 14716 13896 14720
rect 13832 14660 13836 14716
rect 13836 14660 13892 14716
rect 13892 14660 13896 14716
rect 13832 14656 13896 14660
rect 13912 14716 13976 14720
rect 13912 14660 13916 14716
rect 13916 14660 13972 14716
rect 13972 14660 13976 14716
rect 13912 14656 13976 14660
rect 13992 14716 14056 14720
rect 13992 14660 13996 14716
rect 13996 14660 14052 14716
rect 14052 14660 14056 14716
rect 13992 14656 14056 14660
rect 14072 14716 14136 14720
rect 14072 14660 14076 14716
rect 14076 14660 14132 14716
rect 14132 14660 14136 14716
rect 14072 14656 14136 14660
rect 20548 14716 20612 14720
rect 20548 14660 20552 14716
rect 20552 14660 20608 14716
rect 20608 14660 20612 14716
rect 20548 14656 20612 14660
rect 20628 14716 20692 14720
rect 20628 14660 20632 14716
rect 20632 14660 20688 14716
rect 20688 14660 20692 14716
rect 20628 14656 20692 14660
rect 20708 14716 20772 14720
rect 20708 14660 20712 14716
rect 20712 14660 20768 14716
rect 20768 14660 20772 14716
rect 20708 14656 20772 14660
rect 20788 14716 20852 14720
rect 20788 14660 20792 14716
rect 20792 14660 20848 14716
rect 20848 14660 20852 14716
rect 20788 14656 20852 14660
rect 27264 14716 27328 14720
rect 27264 14660 27268 14716
rect 27268 14660 27324 14716
rect 27324 14660 27328 14716
rect 27264 14656 27328 14660
rect 27344 14716 27408 14720
rect 27344 14660 27348 14716
rect 27348 14660 27404 14716
rect 27404 14660 27408 14716
rect 27344 14656 27408 14660
rect 27424 14716 27488 14720
rect 27424 14660 27428 14716
rect 27428 14660 27484 14716
rect 27484 14660 27488 14716
rect 27424 14656 27488 14660
rect 27504 14716 27568 14720
rect 27504 14660 27508 14716
rect 27508 14660 27564 14716
rect 27564 14660 27568 14716
rect 27504 14656 27568 14660
rect 3758 14172 3822 14176
rect 3758 14116 3762 14172
rect 3762 14116 3818 14172
rect 3818 14116 3822 14172
rect 3758 14112 3822 14116
rect 3838 14172 3902 14176
rect 3838 14116 3842 14172
rect 3842 14116 3898 14172
rect 3898 14116 3902 14172
rect 3838 14112 3902 14116
rect 3918 14172 3982 14176
rect 3918 14116 3922 14172
rect 3922 14116 3978 14172
rect 3978 14116 3982 14172
rect 3918 14112 3982 14116
rect 3998 14172 4062 14176
rect 3998 14116 4002 14172
rect 4002 14116 4058 14172
rect 4058 14116 4062 14172
rect 3998 14112 4062 14116
rect 10474 14172 10538 14176
rect 10474 14116 10478 14172
rect 10478 14116 10534 14172
rect 10534 14116 10538 14172
rect 10474 14112 10538 14116
rect 10554 14172 10618 14176
rect 10554 14116 10558 14172
rect 10558 14116 10614 14172
rect 10614 14116 10618 14172
rect 10554 14112 10618 14116
rect 10634 14172 10698 14176
rect 10634 14116 10638 14172
rect 10638 14116 10694 14172
rect 10694 14116 10698 14172
rect 10634 14112 10698 14116
rect 10714 14172 10778 14176
rect 10714 14116 10718 14172
rect 10718 14116 10774 14172
rect 10774 14116 10778 14172
rect 10714 14112 10778 14116
rect 17190 14172 17254 14176
rect 17190 14116 17194 14172
rect 17194 14116 17250 14172
rect 17250 14116 17254 14172
rect 17190 14112 17254 14116
rect 17270 14172 17334 14176
rect 17270 14116 17274 14172
rect 17274 14116 17330 14172
rect 17330 14116 17334 14172
rect 17270 14112 17334 14116
rect 17350 14172 17414 14176
rect 17350 14116 17354 14172
rect 17354 14116 17410 14172
rect 17410 14116 17414 14172
rect 17350 14112 17414 14116
rect 17430 14172 17494 14176
rect 17430 14116 17434 14172
rect 17434 14116 17490 14172
rect 17490 14116 17494 14172
rect 17430 14112 17494 14116
rect 23906 14172 23970 14176
rect 23906 14116 23910 14172
rect 23910 14116 23966 14172
rect 23966 14116 23970 14172
rect 23906 14112 23970 14116
rect 23986 14172 24050 14176
rect 23986 14116 23990 14172
rect 23990 14116 24046 14172
rect 24046 14116 24050 14172
rect 23986 14112 24050 14116
rect 24066 14172 24130 14176
rect 24066 14116 24070 14172
rect 24070 14116 24126 14172
rect 24126 14116 24130 14172
rect 24066 14112 24130 14116
rect 24146 14172 24210 14176
rect 24146 14116 24150 14172
rect 24150 14116 24206 14172
rect 24206 14116 24210 14172
rect 24146 14112 24210 14116
rect 7116 13628 7180 13632
rect 7116 13572 7120 13628
rect 7120 13572 7176 13628
rect 7176 13572 7180 13628
rect 7116 13568 7180 13572
rect 7196 13628 7260 13632
rect 7196 13572 7200 13628
rect 7200 13572 7256 13628
rect 7256 13572 7260 13628
rect 7196 13568 7260 13572
rect 7276 13628 7340 13632
rect 7276 13572 7280 13628
rect 7280 13572 7336 13628
rect 7336 13572 7340 13628
rect 7276 13568 7340 13572
rect 7356 13628 7420 13632
rect 7356 13572 7360 13628
rect 7360 13572 7416 13628
rect 7416 13572 7420 13628
rect 7356 13568 7420 13572
rect 13832 13628 13896 13632
rect 13832 13572 13836 13628
rect 13836 13572 13892 13628
rect 13892 13572 13896 13628
rect 13832 13568 13896 13572
rect 13912 13628 13976 13632
rect 13912 13572 13916 13628
rect 13916 13572 13972 13628
rect 13972 13572 13976 13628
rect 13912 13568 13976 13572
rect 13992 13628 14056 13632
rect 13992 13572 13996 13628
rect 13996 13572 14052 13628
rect 14052 13572 14056 13628
rect 13992 13568 14056 13572
rect 14072 13628 14136 13632
rect 14072 13572 14076 13628
rect 14076 13572 14132 13628
rect 14132 13572 14136 13628
rect 14072 13568 14136 13572
rect 20548 13628 20612 13632
rect 20548 13572 20552 13628
rect 20552 13572 20608 13628
rect 20608 13572 20612 13628
rect 20548 13568 20612 13572
rect 20628 13628 20692 13632
rect 20628 13572 20632 13628
rect 20632 13572 20688 13628
rect 20688 13572 20692 13628
rect 20628 13568 20692 13572
rect 20708 13628 20772 13632
rect 20708 13572 20712 13628
rect 20712 13572 20768 13628
rect 20768 13572 20772 13628
rect 20708 13568 20772 13572
rect 20788 13628 20852 13632
rect 20788 13572 20792 13628
rect 20792 13572 20848 13628
rect 20848 13572 20852 13628
rect 20788 13568 20852 13572
rect 27264 13628 27328 13632
rect 27264 13572 27268 13628
rect 27268 13572 27324 13628
rect 27324 13572 27328 13628
rect 27264 13568 27328 13572
rect 27344 13628 27408 13632
rect 27344 13572 27348 13628
rect 27348 13572 27404 13628
rect 27404 13572 27408 13628
rect 27344 13568 27408 13572
rect 27424 13628 27488 13632
rect 27424 13572 27428 13628
rect 27428 13572 27484 13628
rect 27484 13572 27488 13628
rect 27424 13568 27488 13572
rect 27504 13628 27568 13632
rect 27504 13572 27508 13628
rect 27508 13572 27564 13628
rect 27564 13572 27568 13628
rect 27504 13568 27568 13572
rect 3758 13084 3822 13088
rect 3758 13028 3762 13084
rect 3762 13028 3818 13084
rect 3818 13028 3822 13084
rect 3758 13024 3822 13028
rect 3838 13084 3902 13088
rect 3838 13028 3842 13084
rect 3842 13028 3898 13084
rect 3898 13028 3902 13084
rect 3838 13024 3902 13028
rect 3918 13084 3982 13088
rect 3918 13028 3922 13084
rect 3922 13028 3978 13084
rect 3978 13028 3982 13084
rect 3918 13024 3982 13028
rect 3998 13084 4062 13088
rect 3998 13028 4002 13084
rect 4002 13028 4058 13084
rect 4058 13028 4062 13084
rect 3998 13024 4062 13028
rect 10474 13084 10538 13088
rect 10474 13028 10478 13084
rect 10478 13028 10534 13084
rect 10534 13028 10538 13084
rect 10474 13024 10538 13028
rect 10554 13084 10618 13088
rect 10554 13028 10558 13084
rect 10558 13028 10614 13084
rect 10614 13028 10618 13084
rect 10554 13024 10618 13028
rect 10634 13084 10698 13088
rect 10634 13028 10638 13084
rect 10638 13028 10694 13084
rect 10694 13028 10698 13084
rect 10634 13024 10698 13028
rect 10714 13084 10778 13088
rect 10714 13028 10718 13084
rect 10718 13028 10774 13084
rect 10774 13028 10778 13084
rect 10714 13024 10778 13028
rect 17190 13084 17254 13088
rect 17190 13028 17194 13084
rect 17194 13028 17250 13084
rect 17250 13028 17254 13084
rect 17190 13024 17254 13028
rect 17270 13084 17334 13088
rect 17270 13028 17274 13084
rect 17274 13028 17330 13084
rect 17330 13028 17334 13084
rect 17270 13024 17334 13028
rect 17350 13084 17414 13088
rect 17350 13028 17354 13084
rect 17354 13028 17410 13084
rect 17410 13028 17414 13084
rect 17350 13024 17414 13028
rect 17430 13084 17494 13088
rect 17430 13028 17434 13084
rect 17434 13028 17490 13084
rect 17490 13028 17494 13084
rect 17430 13024 17494 13028
rect 23906 13084 23970 13088
rect 23906 13028 23910 13084
rect 23910 13028 23966 13084
rect 23966 13028 23970 13084
rect 23906 13024 23970 13028
rect 23986 13084 24050 13088
rect 23986 13028 23990 13084
rect 23990 13028 24046 13084
rect 24046 13028 24050 13084
rect 23986 13024 24050 13028
rect 24066 13084 24130 13088
rect 24066 13028 24070 13084
rect 24070 13028 24126 13084
rect 24126 13028 24130 13084
rect 24066 13024 24130 13028
rect 24146 13084 24210 13088
rect 24146 13028 24150 13084
rect 24150 13028 24206 13084
rect 24206 13028 24210 13084
rect 24146 13024 24210 13028
rect 7116 12540 7180 12544
rect 7116 12484 7120 12540
rect 7120 12484 7176 12540
rect 7176 12484 7180 12540
rect 7116 12480 7180 12484
rect 7196 12540 7260 12544
rect 7196 12484 7200 12540
rect 7200 12484 7256 12540
rect 7256 12484 7260 12540
rect 7196 12480 7260 12484
rect 7276 12540 7340 12544
rect 7276 12484 7280 12540
rect 7280 12484 7336 12540
rect 7336 12484 7340 12540
rect 7276 12480 7340 12484
rect 7356 12540 7420 12544
rect 7356 12484 7360 12540
rect 7360 12484 7416 12540
rect 7416 12484 7420 12540
rect 7356 12480 7420 12484
rect 13832 12540 13896 12544
rect 13832 12484 13836 12540
rect 13836 12484 13892 12540
rect 13892 12484 13896 12540
rect 13832 12480 13896 12484
rect 13912 12540 13976 12544
rect 13912 12484 13916 12540
rect 13916 12484 13972 12540
rect 13972 12484 13976 12540
rect 13912 12480 13976 12484
rect 13992 12540 14056 12544
rect 13992 12484 13996 12540
rect 13996 12484 14052 12540
rect 14052 12484 14056 12540
rect 13992 12480 14056 12484
rect 14072 12540 14136 12544
rect 14072 12484 14076 12540
rect 14076 12484 14132 12540
rect 14132 12484 14136 12540
rect 14072 12480 14136 12484
rect 20548 12540 20612 12544
rect 20548 12484 20552 12540
rect 20552 12484 20608 12540
rect 20608 12484 20612 12540
rect 20548 12480 20612 12484
rect 20628 12540 20692 12544
rect 20628 12484 20632 12540
rect 20632 12484 20688 12540
rect 20688 12484 20692 12540
rect 20628 12480 20692 12484
rect 20708 12540 20772 12544
rect 20708 12484 20712 12540
rect 20712 12484 20768 12540
rect 20768 12484 20772 12540
rect 20708 12480 20772 12484
rect 20788 12540 20852 12544
rect 20788 12484 20792 12540
rect 20792 12484 20848 12540
rect 20848 12484 20852 12540
rect 20788 12480 20852 12484
rect 27264 12540 27328 12544
rect 27264 12484 27268 12540
rect 27268 12484 27324 12540
rect 27324 12484 27328 12540
rect 27264 12480 27328 12484
rect 27344 12540 27408 12544
rect 27344 12484 27348 12540
rect 27348 12484 27404 12540
rect 27404 12484 27408 12540
rect 27344 12480 27408 12484
rect 27424 12540 27488 12544
rect 27424 12484 27428 12540
rect 27428 12484 27484 12540
rect 27484 12484 27488 12540
rect 27424 12480 27488 12484
rect 27504 12540 27568 12544
rect 27504 12484 27508 12540
rect 27508 12484 27564 12540
rect 27564 12484 27568 12540
rect 27504 12480 27568 12484
rect 3758 11996 3822 12000
rect 3758 11940 3762 11996
rect 3762 11940 3818 11996
rect 3818 11940 3822 11996
rect 3758 11936 3822 11940
rect 3838 11996 3902 12000
rect 3838 11940 3842 11996
rect 3842 11940 3898 11996
rect 3898 11940 3902 11996
rect 3838 11936 3902 11940
rect 3918 11996 3982 12000
rect 3918 11940 3922 11996
rect 3922 11940 3978 11996
rect 3978 11940 3982 11996
rect 3918 11936 3982 11940
rect 3998 11996 4062 12000
rect 3998 11940 4002 11996
rect 4002 11940 4058 11996
rect 4058 11940 4062 11996
rect 3998 11936 4062 11940
rect 10474 11996 10538 12000
rect 10474 11940 10478 11996
rect 10478 11940 10534 11996
rect 10534 11940 10538 11996
rect 10474 11936 10538 11940
rect 10554 11996 10618 12000
rect 10554 11940 10558 11996
rect 10558 11940 10614 11996
rect 10614 11940 10618 11996
rect 10554 11936 10618 11940
rect 10634 11996 10698 12000
rect 10634 11940 10638 11996
rect 10638 11940 10694 11996
rect 10694 11940 10698 11996
rect 10634 11936 10698 11940
rect 10714 11996 10778 12000
rect 10714 11940 10718 11996
rect 10718 11940 10774 11996
rect 10774 11940 10778 11996
rect 10714 11936 10778 11940
rect 17190 11996 17254 12000
rect 17190 11940 17194 11996
rect 17194 11940 17250 11996
rect 17250 11940 17254 11996
rect 17190 11936 17254 11940
rect 17270 11996 17334 12000
rect 17270 11940 17274 11996
rect 17274 11940 17330 11996
rect 17330 11940 17334 11996
rect 17270 11936 17334 11940
rect 17350 11996 17414 12000
rect 17350 11940 17354 11996
rect 17354 11940 17410 11996
rect 17410 11940 17414 11996
rect 17350 11936 17414 11940
rect 17430 11996 17494 12000
rect 17430 11940 17434 11996
rect 17434 11940 17490 11996
rect 17490 11940 17494 11996
rect 17430 11936 17494 11940
rect 23906 11996 23970 12000
rect 23906 11940 23910 11996
rect 23910 11940 23966 11996
rect 23966 11940 23970 11996
rect 23906 11936 23970 11940
rect 23986 11996 24050 12000
rect 23986 11940 23990 11996
rect 23990 11940 24046 11996
rect 24046 11940 24050 11996
rect 23986 11936 24050 11940
rect 24066 11996 24130 12000
rect 24066 11940 24070 11996
rect 24070 11940 24126 11996
rect 24126 11940 24130 11996
rect 24066 11936 24130 11940
rect 24146 11996 24210 12000
rect 24146 11940 24150 11996
rect 24150 11940 24206 11996
rect 24206 11940 24210 11996
rect 24146 11936 24210 11940
rect 7116 11452 7180 11456
rect 7116 11396 7120 11452
rect 7120 11396 7176 11452
rect 7176 11396 7180 11452
rect 7116 11392 7180 11396
rect 7196 11452 7260 11456
rect 7196 11396 7200 11452
rect 7200 11396 7256 11452
rect 7256 11396 7260 11452
rect 7196 11392 7260 11396
rect 7276 11452 7340 11456
rect 7276 11396 7280 11452
rect 7280 11396 7336 11452
rect 7336 11396 7340 11452
rect 7276 11392 7340 11396
rect 7356 11452 7420 11456
rect 7356 11396 7360 11452
rect 7360 11396 7416 11452
rect 7416 11396 7420 11452
rect 7356 11392 7420 11396
rect 13832 11452 13896 11456
rect 13832 11396 13836 11452
rect 13836 11396 13892 11452
rect 13892 11396 13896 11452
rect 13832 11392 13896 11396
rect 13912 11452 13976 11456
rect 13912 11396 13916 11452
rect 13916 11396 13972 11452
rect 13972 11396 13976 11452
rect 13912 11392 13976 11396
rect 13992 11452 14056 11456
rect 13992 11396 13996 11452
rect 13996 11396 14052 11452
rect 14052 11396 14056 11452
rect 13992 11392 14056 11396
rect 14072 11452 14136 11456
rect 14072 11396 14076 11452
rect 14076 11396 14132 11452
rect 14132 11396 14136 11452
rect 14072 11392 14136 11396
rect 20548 11452 20612 11456
rect 20548 11396 20552 11452
rect 20552 11396 20608 11452
rect 20608 11396 20612 11452
rect 20548 11392 20612 11396
rect 20628 11452 20692 11456
rect 20628 11396 20632 11452
rect 20632 11396 20688 11452
rect 20688 11396 20692 11452
rect 20628 11392 20692 11396
rect 20708 11452 20772 11456
rect 20708 11396 20712 11452
rect 20712 11396 20768 11452
rect 20768 11396 20772 11452
rect 20708 11392 20772 11396
rect 20788 11452 20852 11456
rect 20788 11396 20792 11452
rect 20792 11396 20848 11452
rect 20848 11396 20852 11452
rect 20788 11392 20852 11396
rect 27264 11452 27328 11456
rect 27264 11396 27268 11452
rect 27268 11396 27324 11452
rect 27324 11396 27328 11452
rect 27264 11392 27328 11396
rect 27344 11452 27408 11456
rect 27344 11396 27348 11452
rect 27348 11396 27404 11452
rect 27404 11396 27408 11452
rect 27344 11392 27408 11396
rect 27424 11452 27488 11456
rect 27424 11396 27428 11452
rect 27428 11396 27484 11452
rect 27484 11396 27488 11452
rect 27424 11392 27488 11396
rect 27504 11452 27568 11456
rect 27504 11396 27508 11452
rect 27508 11396 27564 11452
rect 27564 11396 27568 11452
rect 27504 11392 27568 11396
rect 3758 10908 3822 10912
rect 3758 10852 3762 10908
rect 3762 10852 3818 10908
rect 3818 10852 3822 10908
rect 3758 10848 3822 10852
rect 3838 10908 3902 10912
rect 3838 10852 3842 10908
rect 3842 10852 3898 10908
rect 3898 10852 3902 10908
rect 3838 10848 3902 10852
rect 3918 10908 3982 10912
rect 3918 10852 3922 10908
rect 3922 10852 3978 10908
rect 3978 10852 3982 10908
rect 3918 10848 3982 10852
rect 3998 10908 4062 10912
rect 3998 10852 4002 10908
rect 4002 10852 4058 10908
rect 4058 10852 4062 10908
rect 3998 10848 4062 10852
rect 10474 10908 10538 10912
rect 10474 10852 10478 10908
rect 10478 10852 10534 10908
rect 10534 10852 10538 10908
rect 10474 10848 10538 10852
rect 10554 10908 10618 10912
rect 10554 10852 10558 10908
rect 10558 10852 10614 10908
rect 10614 10852 10618 10908
rect 10554 10848 10618 10852
rect 10634 10908 10698 10912
rect 10634 10852 10638 10908
rect 10638 10852 10694 10908
rect 10694 10852 10698 10908
rect 10634 10848 10698 10852
rect 10714 10908 10778 10912
rect 10714 10852 10718 10908
rect 10718 10852 10774 10908
rect 10774 10852 10778 10908
rect 10714 10848 10778 10852
rect 17190 10908 17254 10912
rect 17190 10852 17194 10908
rect 17194 10852 17250 10908
rect 17250 10852 17254 10908
rect 17190 10848 17254 10852
rect 17270 10908 17334 10912
rect 17270 10852 17274 10908
rect 17274 10852 17330 10908
rect 17330 10852 17334 10908
rect 17270 10848 17334 10852
rect 17350 10908 17414 10912
rect 17350 10852 17354 10908
rect 17354 10852 17410 10908
rect 17410 10852 17414 10908
rect 17350 10848 17414 10852
rect 17430 10908 17494 10912
rect 17430 10852 17434 10908
rect 17434 10852 17490 10908
rect 17490 10852 17494 10908
rect 17430 10848 17494 10852
rect 23906 10908 23970 10912
rect 23906 10852 23910 10908
rect 23910 10852 23966 10908
rect 23966 10852 23970 10908
rect 23906 10848 23970 10852
rect 23986 10908 24050 10912
rect 23986 10852 23990 10908
rect 23990 10852 24046 10908
rect 24046 10852 24050 10908
rect 23986 10848 24050 10852
rect 24066 10908 24130 10912
rect 24066 10852 24070 10908
rect 24070 10852 24126 10908
rect 24126 10852 24130 10908
rect 24066 10848 24130 10852
rect 24146 10908 24210 10912
rect 24146 10852 24150 10908
rect 24150 10852 24206 10908
rect 24206 10852 24210 10908
rect 24146 10848 24210 10852
rect 2084 10508 2148 10572
rect 7116 10364 7180 10368
rect 7116 10308 7120 10364
rect 7120 10308 7176 10364
rect 7176 10308 7180 10364
rect 7116 10304 7180 10308
rect 7196 10364 7260 10368
rect 7196 10308 7200 10364
rect 7200 10308 7256 10364
rect 7256 10308 7260 10364
rect 7196 10304 7260 10308
rect 7276 10364 7340 10368
rect 7276 10308 7280 10364
rect 7280 10308 7336 10364
rect 7336 10308 7340 10364
rect 7276 10304 7340 10308
rect 7356 10364 7420 10368
rect 7356 10308 7360 10364
rect 7360 10308 7416 10364
rect 7416 10308 7420 10364
rect 7356 10304 7420 10308
rect 13832 10364 13896 10368
rect 13832 10308 13836 10364
rect 13836 10308 13892 10364
rect 13892 10308 13896 10364
rect 13832 10304 13896 10308
rect 13912 10364 13976 10368
rect 13912 10308 13916 10364
rect 13916 10308 13972 10364
rect 13972 10308 13976 10364
rect 13912 10304 13976 10308
rect 13992 10364 14056 10368
rect 13992 10308 13996 10364
rect 13996 10308 14052 10364
rect 14052 10308 14056 10364
rect 13992 10304 14056 10308
rect 14072 10364 14136 10368
rect 14072 10308 14076 10364
rect 14076 10308 14132 10364
rect 14132 10308 14136 10364
rect 14072 10304 14136 10308
rect 20548 10364 20612 10368
rect 20548 10308 20552 10364
rect 20552 10308 20608 10364
rect 20608 10308 20612 10364
rect 20548 10304 20612 10308
rect 20628 10364 20692 10368
rect 20628 10308 20632 10364
rect 20632 10308 20688 10364
rect 20688 10308 20692 10364
rect 20628 10304 20692 10308
rect 20708 10364 20772 10368
rect 20708 10308 20712 10364
rect 20712 10308 20768 10364
rect 20768 10308 20772 10364
rect 20708 10304 20772 10308
rect 20788 10364 20852 10368
rect 20788 10308 20792 10364
rect 20792 10308 20848 10364
rect 20848 10308 20852 10364
rect 20788 10304 20852 10308
rect 27264 10364 27328 10368
rect 27264 10308 27268 10364
rect 27268 10308 27324 10364
rect 27324 10308 27328 10364
rect 27264 10304 27328 10308
rect 27344 10364 27408 10368
rect 27344 10308 27348 10364
rect 27348 10308 27404 10364
rect 27404 10308 27408 10364
rect 27344 10304 27408 10308
rect 27424 10364 27488 10368
rect 27424 10308 27428 10364
rect 27428 10308 27484 10364
rect 27484 10308 27488 10364
rect 27424 10304 27488 10308
rect 27504 10364 27568 10368
rect 27504 10308 27508 10364
rect 27508 10308 27564 10364
rect 27564 10308 27568 10364
rect 27504 10304 27568 10308
rect 3758 9820 3822 9824
rect 3758 9764 3762 9820
rect 3762 9764 3818 9820
rect 3818 9764 3822 9820
rect 3758 9760 3822 9764
rect 3838 9820 3902 9824
rect 3838 9764 3842 9820
rect 3842 9764 3898 9820
rect 3898 9764 3902 9820
rect 3838 9760 3902 9764
rect 3918 9820 3982 9824
rect 3918 9764 3922 9820
rect 3922 9764 3978 9820
rect 3978 9764 3982 9820
rect 3918 9760 3982 9764
rect 3998 9820 4062 9824
rect 3998 9764 4002 9820
rect 4002 9764 4058 9820
rect 4058 9764 4062 9820
rect 3998 9760 4062 9764
rect 10474 9820 10538 9824
rect 10474 9764 10478 9820
rect 10478 9764 10534 9820
rect 10534 9764 10538 9820
rect 10474 9760 10538 9764
rect 10554 9820 10618 9824
rect 10554 9764 10558 9820
rect 10558 9764 10614 9820
rect 10614 9764 10618 9820
rect 10554 9760 10618 9764
rect 10634 9820 10698 9824
rect 10634 9764 10638 9820
rect 10638 9764 10694 9820
rect 10694 9764 10698 9820
rect 10634 9760 10698 9764
rect 10714 9820 10778 9824
rect 10714 9764 10718 9820
rect 10718 9764 10774 9820
rect 10774 9764 10778 9820
rect 10714 9760 10778 9764
rect 17190 9820 17254 9824
rect 17190 9764 17194 9820
rect 17194 9764 17250 9820
rect 17250 9764 17254 9820
rect 17190 9760 17254 9764
rect 17270 9820 17334 9824
rect 17270 9764 17274 9820
rect 17274 9764 17330 9820
rect 17330 9764 17334 9820
rect 17270 9760 17334 9764
rect 17350 9820 17414 9824
rect 17350 9764 17354 9820
rect 17354 9764 17410 9820
rect 17410 9764 17414 9820
rect 17350 9760 17414 9764
rect 17430 9820 17494 9824
rect 17430 9764 17434 9820
rect 17434 9764 17490 9820
rect 17490 9764 17494 9820
rect 17430 9760 17494 9764
rect 23906 9820 23970 9824
rect 23906 9764 23910 9820
rect 23910 9764 23966 9820
rect 23966 9764 23970 9820
rect 23906 9760 23970 9764
rect 23986 9820 24050 9824
rect 23986 9764 23990 9820
rect 23990 9764 24046 9820
rect 24046 9764 24050 9820
rect 23986 9760 24050 9764
rect 24066 9820 24130 9824
rect 24066 9764 24070 9820
rect 24070 9764 24126 9820
rect 24126 9764 24130 9820
rect 24066 9760 24130 9764
rect 24146 9820 24210 9824
rect 24146 9764 24150 9820
rect 24150 9764 24206 9820
rect 24206 9764 24210 9820
rect 24146 9760 24210 9764
rect 7116 9276 7180 9280
rect 7116 9220 7120 9276
rect 7120 9220 7176 9276
rect 7176 9220 7180 9276
rect 7116 9216 7180 9220
rect 7196 9276 7260 9280
rect 7196 9220 7200 9276
rect 7200 9220 7256 9276
rect 7256 9220 7260 9276
rect 7196 9216 7260 9220
rect 7276 9276 7340 9280
rect 7276 9220 7280 9276
rect 7280 9220 7336 9276
rect 7336 9220 7340 9276
rect 7276 9216 7340 9220
rect 7356 9276 7420 9280
rect 7356 9220 7360 9276
rect 7360 9220 7416 9276
rect 7416 9220 7420 9276
rect 7356 9216 7420 9220
rect 13832 9276 13896 9280
rect 13832 9220 13836 9276
rect 13836 9220 13892 9276
rect 13892 9220 13896 9276
rect 13832 9216 13896 9220
rect 13912 9276 13976 9280
rect 13912 9220 13916 9276
rect 13916 9220 13972 9276
rect 13972 9220 13976 9276
rect 13912 9216 13976 9220
rect 13992 9276 14056 9280
rect 13992 9220 13996 9276
rect 13996 9220 14052 9276
rect 14052 9220 14056 9276
rect 13992 9216 14056 9220
rect 14072 9276 14136 9280
rect 14072 9220 14076 9276
rect 14076 9220 14132 9276
rect 14132 9220 14136 9276
rect 14072 9216 14136 9220
rect 20548 9276 20612 9280
rect 20548 9220 20552 9276
rect 20552 9220 20608 9276
rect 20608 9220 20612 9276
rect 20548 9216 20612 9220
rect 20628 9276 20692 9280
rect 20628 9220 20632 9276
rect 20632 9220 20688 9276
rect 20688 9220 20692 9276
rect 20628 9216 20692 9220
rect 20708 9276 20772 9280
rect 20708 9220 20712 9276
rect 20712 9220 20768 9276
rect 20768 9220 20772 9276
rect 20708 9216 20772 9220
rect 20788 9276 20852 9280
rect 20788 9220 20792 9276
rect 20792 9220 20848 9276
rect 20848 9220 20852 9276
rect 20788 9216 20852 9220
rect 27264 9276 27328 9280
rect 27264 9220 27268 9276
rect 27268 9220 27324 9276
rect 27324 9220 27328 9276
rect 27264 9216 27328 9220
rect 27344 9276 27408 9280
rect 27344 9220 27348 9276
rect 27348 9220 27404 9276
rect 27404 9220 27408 9276
rect 27344 9216 27408 9220
rect 27424 9276 27488 9280
rect 27424 9220 27428 9276
rect 27428 9220 27484 9276
rect 27484 9220 27488 9276
rect 27424 9216 27488 9220
rect 27504 9276 27568 9280
rect 27504 9220 27508 9276
rect 27508 9220 27564 9276
rect 27564 9220 27568 9276
rect 27504 9216 27568 9220
rect 3758 8732 3822 8736
rect 3758 8676 3762 8732
rect 3762 8676 3818 8732
rect 3818 8676 3822 8732
rect 3758 8672 3822 8676
rect 3838 8732 3902 8736
rect 3838 8676 3842 8732
rect 3842 8676 3898 8732
rect 3898 8676 3902 8732
rect 3838 8672 3902 8676
rect 3918 8732 3982 8736
rect 3918 8676 3922 8732
rect 3922 8676 3978 8732
rect 3978 8676 3982 8732
rect 3918 8672 3982 8676
rect 3998 8732 4062 8736
rect 3998 8676 4002 8732
rect 4002 8676 4058 8732
rect 4058 8676 4062 8732
rect 3998 8672 4062 8676
rect 10474 8732 10538 8736
rect 10474 8676 10478 8732
rect 10478 8676 10534 8732
rect 10534 8676 10538 8732
rect 10474 8672 10538 8676
rect 10554 8732 10618 8736
rect 10554 8676 10558 8732
rect 10558 8676 10614 8732
rect 10614 8676 10618 8732
rect 10554 8672 10618 8676
rect 10634 8732 10698 8736
rect 10634 8676 10638 8732
rect 10638 8676 10694 8732
rect 10694 8676 10698 8732
rect 10634 8672 10698 8676
rect 10714 8732 10778 8736
rect 10714 8676 10718 8732
rect 10718 8676 10774 8732
rect 10774 8676 10778 8732
rect 10714 8672 10778 8676
rect 17190 8732 17254 8736
rect 17190 8676 17194 8732
rect 17194 8676 17250 8732
rect 17250 8676 17254 8732
rect 17190 8672 17254 8676
rect 17270 8732 17334 8736
rect 17270 8676 17274 8732
rect 17274 8676 17330 8732
rect 17330 8676 17334 8732
rect 17270 8672 17334 8676
rect 17350 8732 17414 8736
rect 17350 8676 17354 8732
rect 17354 8676 17410 8732
rect 17410 8676 17414 8732
rect 17350 8672 17414 8676
rect 17430 8732 17494 8736
rect 17430 8676 17434 8732
rect 17434 8676 17490 8732
rect 17490 8676 17494 8732
rect 17430 8672 17494 8676
rect 23906 8732 23970 8736
rect 23906 8676 23910 8732
rect 23910 8676 23966 8732
rect 23966 8676 23970 8732
rect 23906 8672 23970 8676
rect 23986 8732 24050 8736
rect 23986 8676 23990 8732
rect 23990 8676 24046 8732
rect 24046 8676 24050 8732
rect 23986 8672 24050 8676
rect 24066 8732 24130 8736
rect 24066 8676 24070 8732
rect 24070 8676 24126 8732
rect 24126 8676 24130 8732
rect 24066 8672 24130 8676
rect 24146 8732 24210 8736
rect 24146 8676 24150 8732
rect 24150 8676 24206 8732
rect 24206 8676 24210 8732
rect 24146 8672 24210 8676
rect 7116 8188 7180 8192
rect 7116 8132 7120 8188
rect 7120 8132 7176 8188
rect 7176 8132 7180 8188
rect 7116 8128 7180 8132
rect 7196 8188 7260 8192
rect 7196 8132 7200 8188
rect 7200 8132 7256 8188
rect 7256 8132 7260 8188
rect 7196 8128 7260 8132
rect 7276 8188 7340 8192
rect 7276 8132 7280 8188
rect 7280 8132 7336 8188
rect 7336 8132 7340 8188
rect 7276 8128 7340 8132
rect 7356 8188 7420 8192
rect 7356 8132 7360 8188
rect 7360 8132 7416 8188
rect 7416 8132 7420 8188
rect 7356 8128 7420 8132
rect 13832 8188 13896 8192
rect 13832 8132 13836 8188
rect 13836 8132 13892 8188
rect 13892 8132 13896 8188
rect 13832 8128 13896 8132
rect 13912 8188 13976 8192
rect 13912 8132 13916 8188
rect 13916 8132 13972 8188
rect 13972 8132 13976 8188
rect 13912 8128 13976 8132
rect 13992 8188 14056 8192
rect 13992 8132 13996 8188
rect 13996 8132 14052 8188
rect 14052 8132 14056 8188
rect 13992 8128 14056 8132
rect 14072 8188 14136 8192
rect 14072 8132 14076 8188
rect 14076 8132 14132 8188
rect 14132 8132 14136 8188
rect 14072 8128 14136 8132
rect 20548 8188 20612 8192
rect 20548 8132 20552 8188
rect 20552 8132 20608 8188
rect 20608 8132 20612 8188
rect 20548 8128 20612 8132
rect 20628 8188 20692 8192
rect 20628 8132 20632 8188
rect 20632 8132 20688 8188
rect 20688 8132 20692 8188
rect 20628 8128 20692 8132
rect 20708 8188 20772 8192
rect 20708 8132 20712 8188
rect 20712 8132 20768 8188
rect 20768 8132 20772 8188
rect 20708 8128 20772 8132
rect 20788 8188 20852 8192
rect 20788 8132 20792 8188
rect 20792 8132 20848 8188
rect 20848 8132 20852 8188
rect 20788 8128 20852 8132
rect 27264 8188 27328 8192
rect 27264 8132 27268 8188
rect 27268 8132 27324 8188
rect 27324 8132 27328 8188
rect 27264 8128 27328 8132
rect 27344 8188 27408 8192
rect 27344 8132 27348 8188
rect 27348 8132 27404 8188
rect 27404 8132 27408 8188
rect 27344 8128 27408 8132
rect 27424 8188 27488 8192
rect 27424 8132 27428 8188
rect 27428 8132 27484 8188
rect 27484 8132 27488 8188
rect 27424 8128 27488 8132
rect 27504 8188 27568 8192
rect 27504 8132 27508 8188
rect 27508 8132 27564 8188
rect 27564 8132 27568 8188
rect 27504 8128 27568 8132
rect 3758 7644 3822 7648
rect 3758 7588 3762 7644
rect 3762 7588 3818 7644
rect 3818 7588 3822 7644
rect 3758 7584 3822 7588
rect 3838 7644 3902 7648
rect 3838 7588 3842 7644
rect 3842 7588 3898 7644
rect 3898 7588 3902 7644
rect 3838 7584 3902 7588
rect 3918 7644 3982 7648
rect 3918 7588 3922 7644
rect 3922 7588 3978 7644
rect 3978 7588 3982 7644
rect 3918 7584 3982 7588
rect 3998 7644 4062 7648
rect 3998 7588 4002 7644
rect 4002 7588 4058 7644
rect 4058 7588 4062 7644
rect 3998 7584 4062 7588
rect 10474 7644 10538 7648
rect 10474 7588 10478 7644
rect 10478 7588 10534 7644
rect 10534 7588 10538 7644
rect 10474 7584 10538 7588
rect 10554 7644 10618 7648
rect 10554 7588 10558 7644
rect 10558 7588 10614 7644
rect 10614 7588 10618 7644
rect 10554 7584 10618 7588
rect 10634 7644 10698 7648
rect 10634 7588 10638 7644
rect 10638 7588 10694 7644
rect 10694 7588 10698 7644
rect 10634 7584 10698 7588
rect 10714 7644 10778 7648
rect 10714 7588 10718 7644
rect 10718 7588 10774 7644
rect 10774 7588 10778 7644
rect 10714 7584 10778 7588
rect 17190 7644 17254 7648
rect 17190 7588 17194 7644
rect 17194 7588 17250 7644
rect 17250 7588 17254 7644
rect 17190 7584 17254 7588
rect 17270 7644 17334 7648
rect 17270 7588 17274 7644
rect 17274 7588 17330 7644
rect 17330 7588 17334 7644
rect 17270 7584 17334 7588
rect 17350 7644 17414 7648
rect 17350 7588 17354 7644
rect 17354 7588 17410 7644
rect 17410 7588 17414 7644
rect 17350 7584 17414 7588
rect 17430 7644 17494 7648
rect 17430 7588 17434 7644
rect 17434 7588 17490 7644
rect 17490 7588 17494 7644
rect 17430 7584 17494 7588
rect 23906 7644 23970 7648
rect 23906 7588 23910 7644
rect 23910 7588 23966 7644
rect 23966 7588 23970 7644
rect 23906 7584 23970 7588
rect 23986 7644 24050 7648
rect 23986 7588 23990 7644
rect 23990 7588 24046 7644
rect 24046 7588 24050 7644
rect 23986 7584 24050 7588
rect 24066 7644 24130 7648
rect 24066 7588 24070 7644
rect 24070 7588 24126 7644
rect 24126 7588 24130 7644
rect 24066 7584 24130 7588
rect 24146 7644 24210 7648
rect 24146 7588 24150 7644
rect 24150 7588 24206 7644
rect 24206 7588 24210 7644
rect 24146 7584 24210 7588
rect 1900 7244 1964 7308
rect 7116 7100 7180 7104
rect 7116 7044 7120 7100
rect 7120 7044 7176 7100
rect 7176 7044 7180 7100
rect 7116 7040 7180 7044
rect 7196 7100 7260 7104
rect 7196 7044 7200 7100
rect 7200 7044 7256 7100
rect 7256 7044 7260 7100
rect 7196 7040 7260 7044
rect 7276 7100 7340 7104
rect 7276 7044 7280 7100
rect 7280 7044 7336 7100
rect 7336 7044 7340 7100
rect 7276 7040 7340 7044
rect 7356 7100 7420 7104
rect 7356 7044 7360 7100
rect 7360 7044 7416 7100
rect 7416 7044 7420 7100
rect 7356 7040 7420 7044
rect 13832 7100 13896 7104
rect 13832 7044 13836 7100
rect 13836 7044 13892 7100
rect 13892 7044 13896 7100
rect 13832 7040 13896 7044
rect 13912 7100 13976 7104
rect 13912 7044 13916 7100
rect 13916 7044 13972 7100
rect 13972 7044 13976 7100
rect 13912 7040 13976 7044
rect 13992 7100 14056 7104
rect 13992 7044 13996 7100
rect 13996 7044 14052 7100
rect 14052 7044 14056 7100
rect 13992 7040 14056 7044
rect 14072 7100 14136 7104
rect 14072 7044 14076 7100
rect 14076 7044 14132 7100
rect 14132 7044 14136 7100
rect 14072 7040 14136 7044
rect 20548 7100 20612 7104
rect 20548 7044 20552 7100
rect 20552 7044 20608 7100
rect 20608 7044 20612 7100
rect 20548 7040 20612 7044
rect 20628 7100 20692 7104
rect 20628 7044 20632 7100
rect 20632 7044 20688 7100
rect 20688 7044 20692 7100
rect 20628 7040 20692 7044
rect 20708 7100 20772 7104
rect 20708 7044 20712 7100
rect 20712 7044 20768 7100
rect 20768 7044 20772 7100
rect 20708 7040 20772 7044
rect 20788 7100 20852 7104
rect 20788 7044 20792 7100
rect 20792 7044 20848 7100
rect 20848 7044 20852 7100
rect 20788 7040 20852 7044
rect 27264 7100 27328 7104
rect 27264 7044 27268 7100
rect 27268 7044 27324 7100
rect 27324 7044 27328 7100
rect 27264 7040 27328 7044
rect 27344 7100 27408 7104
rect 27344 7044 27348 7100
rect 27348 7044 27404 7100
rect 27404 7044 27408 7100
rect 27344 7040 27408 7044
rect 27424 7100 27488 7104
rect 27424 7044 27428 7100
rect 27428 7044 27484 7100
rect 27484 7044 27488 7100
rect 27424 7040 27488 7044
rect 27504 7100 27568 7104
rect 27504 7044 27508 7100
rect 27508 7044 27564 7100
rect 27564 7044 27568 7100
rect 27504 7040 27568 7044
rect 3758 6556 3822 6560
rect 3758 6500 3762 6556
rect 3762 6500 3818 6556
rect 3818 6500 3822 6556
rect 3758 6496 3822 6500
rect 3838 6556 3902 6560
rect 3838 6500 3842 6556
rect 3842 6500 3898 6556
rect 3898 6500 3902 6556
rect 3838 6496 3902 6500
rect 3918 6556 3982 6560
rect 3918 6500 3922 6556
rect 3922 6500 3978 6556
rect 3978 6500 3982 6556
rect 3918 6496 3982 6500
rect 3998 6556 4062 6560
rect 3998 6500 4002 6556
rect 4002 6500 4058 6556
rect 4058 6500 4062 6556
rect 3998 6496 4062 6500
rect 10474 6556 10538 6560
rect 10474 6500 10478 6556
rect 10478 6500 10534 6556
rect 10534 6500 10538 6556
rect 10474 6496 10538 6500
rect 10554 6556 10618 6560
rect 10554 6500 10558 6556
rect 10558 6500 10614 6556
rect 10614 6500 10618 6556
rect 10554 6496 10618 6500
rect 10634 6556 10698 6560
rect 10634 6500 10638 6556
rect 10638 6500 10694 6556
rect 10694 6500 10698 6556
rect 10634 6496 10698 6500
rect 10714 6556 10778 6560
rect 10714 6500 10718 6556
rect 10718 6500 10774 6556
rect 10774 6500 10778 6556
rect 10714 6496 10778 6500
rect 17190 6556 17254 6560
rect 17190 6500 17194 6556
rect 17194 6500 17250 6556
rect 17250 6500 17254 6556
rect 17190 6496 17254 6500
rect 17270 6556 17334 6560
rect 17270 6500 17274 6556
rect 17274 6500 17330 6556
rect 17330 6500 17334 6556
rect 17270 6496 17334 6500
rect 17350 6556 17414 6560
rect 17350 6500 17354 6556
rect 17354 6500 17410 6556
rect 17410 6500 17414 6556
rect 17350 6496 17414 6500
rect 17430 6556 17494 6560
rect 17430 6500 17434 6556
rect 17434 6500 17490 6556
rect 17490 6500 17494 6556
rect 17430 6496 17494 6500
rect 23906 6556 23970 6560
rect 23906 6500 23910 6556
rect 23910 6500 23966 6556
rect 23966 6500 23970 6556
rect 23906 6496 23970 6500
rect 23986 6556 24050 6560
rect 23986 6500 23990 6556
rect 23990 6500 24046 6556
rect 24046 6500 24050 6556
rect 23986 6496 24050 6500
rect 24066 6556 24130 6560
rect 24066 6500 24070 6556
rect 24070 6500 24126 6556
rect 24126 6500 24130 6556
rect 24066 6496 24130 6500
rect 24146 6556 24210 6560
rect 24146 6500 24150 6556
rect 24150 6500 24206 6556
rect 24206 6500 24210 6556
rect 24146 6496 24210 6500
rect 7116 6012 7180 6016
rect 7116 5956 7120 6012
rect 7120 5956 7176 6012
rect 7176 5956 7180 6012
rect 7116 5952 7180 5956
rect 7196 6012 7260 6016
rect 7196 5956 7200 6012
rect 7200 5956 7256 6012
rect 7256 5956 7260 6012
rect 7196 5952 7260 5956
rect 7276 6012 7340 6016
rect 7276 5956 7280 6012
rect 7280 5956 7336 6012
rect 7336 5956 7340 6012
rect 7276 5952 7340 5956
rect 7356 6012 7420 6016
rect 7356 5956 7360 6012
rect 7360 5956 7416 6012
rect 7416 5956 7420 6012
rect 7356 5952 7420 5956
rect 13832 6012 13896 6016
rect 13832 5956 13836 6012
rect 13836 5956 13892 6012
rect 13892 5956 13896 6012
rect 13832 5952 13896 5956
rect 13912 6012 13976 6016
rect 13912 5956 13916 6012
rect 13916 5956 13972 6012
rect 13972 5956 13976 6012
rect 13912 5952 13976 5956
rect 13992 6012 14056 6016
rect 13992 5956 13996 6012
rect 13996 5956 14052 6012
rect 14052 5956 14056 6012
rect 13992 5952 14056 5956
rect 14072 6012 14136 6016
rect 14072 5956 14076 6012
rect 14076 5956 14132 6012
rect 14132 5956 14136 6012
rect 14072 5952 14136 5956
rect 20548 6012 20612 6016
rect 20548 5956 20552 6012
rect 20552 5956 20608 6012
rect 20608 5956 20612 6012
rect 20548 5952 20612 5956
rect 20628 6012 20692 6016
rect 20628 5956 20632 6012
rect 20632 5956 20688 6012
rect 20688 5956 20692 6012
rect 20628 5952 20692 5956
rect 20708 6012 20772 6016
rect 20708 5956 20712 6012
rect 20712 5956 20768 6012
rect 20768 5956 20772 6012
rect 20708 5952 20772 5956
rect 20788 6012 20852 6016
rect 20788 5956 20792 6012
rect 20792 5956 20848 6012
rect 20848 5956 20852 6012
rect 20788 5952 20852 5956
rect 27264 6012 27328 6016
rect 27264 5956 27268 6012
rect 27268 5956 27324 6012
rect 27324 5956 27328 6012
rect 27264 5952 27328 5956
rect 27344 6012 27408 6016
rect 27344 5956 27348 6012
rect 27348 5956 27404 6012
rect 27404 5956 27408 6012
rect 27344 5952 27408 5956
rect 27424 6012 27488 6016
rect 27424 5956 27428 6012
rect 27428 5956 27484 6012
rect 27484 5956 27488 6012
rect 27424 5952 27488 5956
rect 27504 6012 27568 6016
rect 27504 5956 27508 6012
rect 27508 5956 27564 6012
rect 27564 5956 27568 6012
rect 27504 5952 27568 5956
rect 3758 5468 3822 5472
rect 3758 5412 3762 5468
rect 3762 5412 3818 5468
rect 3818 5412 3822 5468
rect 3758 5408 3822 5412
rect 3838 5468 3902 5472
rect 3838 5412 3842 5468
rect 3842 5412 3898 5468
rect 3898 5412 3902 5468
rect 3838 5408 3902 5412
rect 3918 5468 3982 5472
rect 3918 5412 3922 5468
rect 3922 5412 3978 5468
rect 3978 5412 3982 5468
rect 3918 5408 3982 5412
rect 3998 5468 4062 5472
rect 3998 5412 4002 5468
rect 4002 5412 4058 5468
rect 4058 5412 4062 5468
rect 3998 5408 4062 5412
rect 10474 5468 10538 5472
rect 10474 5412 10478 5468
rect 10478 5412 10534 5468
rect 10534 5412 10538 5468
rect 10474 5408 10538 5412
rect 10554 5468 10618 5472
rect 10554 5412 10558 5468
rect 10558 5412 10614 5468
rect 10614 5412 10618 5468
rect 10554 5408 10618 5412
rect 10634 5468 10698 5472
rect 10634 5412 10638 5468
rect 10638 5412 10694 5468
rect 10694 5412 10698 5468
rect 10634 5408 10698 5412
rect 10714 5468 10778 5472
rect 10714 5412 10718 5468
rect 10718 5412 10774 5468
rect 10774 5412 10778 5468
rect 10714 5408 10778 5412
rect 17190 5468 17254 5472
rect 17190 5412 17194 5468
rect 17194 5412 17250 5468
rect 17250 5412 17254 5468
rect 17190 5408 17254 5412
rect 17270 5468 17334 5472
rect 17270 5412 17274 5468
rect 17274 5412 17330 5468
rect 17330 5412 17334 5468
rect 17270 5408 17334 5412
rect 17350 5468 17414 5472
rect 17350 5412 17354 5468
rect 17354 5412 17410 5468
rect 17410 5412 17414 5468
rect 17350 5408 17414 5412
rect 17430 5468 17494 5472
rect 17430 5412 17434 5468
rect 17434 5412 17490 5468
rect 17490 5412 17494 5468
rect 17430 5408 17494 5412
rect 23906 5468 23970 5472
rect 23906 5412 23910 5468
rect 23910 5412 23966 5468
rect 23966 5412 23970 5468
rect 23906 5408 23970 5412
rect 23986 5468 24050 5472
rect 23986 5412 23990 5468
rect 23990 5412 24046 5468
rect 24046 5412 24050 5468
rect 23986 5408 24050 5412
rect 24066 5468 24130 5472
rect 24066 5412 24070 5468
rect 24070 5412 24126 5468
rect 24126 5412 24130 5468
rect 24066 5408 24130 5412
rect 24146 5468 24210 5472
rect 24146 5412 24150 5468
rect 24150 5412 24206 5468
rect 24206 5412 24210 5468
rect 24146 5408 24210 5412
rect 7116 4924 7180 4928
rect 7116 4868 7120 4924
rect 7120 4868 7176 4924
rect 7176 4868 7180 4924
rect 7116 4864 7180 4868
rect 7196 4924 7260 4928
rect 7196 4868 7200 4924
rect 7200 4868 7256 4924
rect 7256 4868 7260 4924
rect 7196 4864 7260 4868
rect 7276 4924 7340 4928
rect 7276 4868 7280 4924
rect 7280 4868 7336 4924
rect 7336 4868 7340 4924
rect 7276 4864 7340 4868
rect 7356 4924 7420 4928
rect 7356 4868 7360 4924
rect 7360 4868 7416 4924
rect 7416 4868 7420 4924
rect 7356 4864 7420 4868
rect 13832 4924 13896 4928
rect 13832 4868 13836 4924
rect 13836 4868 13892 4924
rect 13892 4868 13896 4924
rect 13832 4864 13896 4868
rect 13912 4924 13976 4928
rect 13912 4868 13916 4924
rect 13916 4868 13972 4924
rect 13972 4868 13976 4924
rect 13912 4864 13976 4868
rect 13992 4924 14056 4928
rect 13992 4868 13996 4924
rect 13996 4868 14052 4924
rect 14052 4868 14056 4924
rect 13992 4864 14056 4868
rect 14072 4924 14136 4928
rect 14072 4868 14076 4924
rect 14076 4868 14132 4924
rect 14132 4868 14136 4924
rect 14072 4864 14136 4868
rect 20548 4924 20612 4928
rect 20548 4868 20552 4924
rect 20552 4868 20608 4924
rect 20608 4868 20612 4924
rect 20548 4864 20612 4868
rect 20628 4924 20692 4928
rect 20628 4868 20632 4924
rect 20632 4868 20688 4924
rect 20688 4868 20692 4924
rect 20628 4864 20692 4868
rect 20708 4924 20772 4928
rect 20708 4868 20712 4924
rect 20712 4868 20768 4924
rect 20768 4868 20772 4924
rect 20708 4864 20772 4868
rect 20788 4924 20852 4928
rect 20788 4868 20792 4924
rect 20792 4868 20848 4924
rect 20848 4868 20852 4924
rect 20788 4864 20852 4868
rect 27264 4924 27328 4928
rect 27264 4868 27268 4924
rect 27268 4868 27324 4924
rect 27324 4868 27328 4924
rect 27264 4864 27328 4868
rect 27344 4924 27408 4928
rect 27344 4868 27348 4924
rect 27348 4868 27404 4924
rect 27404 4868 27408 4924
rect 27344 4864 27408 4868
rect 27424 4924 27488 4928
rect 27424 4868 27428 4924
rect 27428 4868 27484 4924
rect 27484 4868 27488 4924
rect 27424 4864 27488 4868
rect 27504 4924 27568 4928
rect 27504 4868 27508 4924
rect 27508 4868 27564 4924
rect 27564 4868 27568 4924
rect 27504 4864 27568 4868
rect 3758 4380 3822 4384
rect 3758 4324 3762 4380
rect 3762 4324 3818 4380
rect 3818 4324 3822 4380
rect 3758 4320 3822 4324
rect 3838 4380 3902 4384
rect 3838 4324 3842 4380
rect 3842 4324 3898 4380
rect 3898 4324 3902 4380
rect 3838 4320 3902 4324
rect 3918 4380 3982 4384
rect 3918 4324 3922 4380
rect 3922 4324 3978 4380
rect 3978 4324 3982 4380
rect 3918 4320 3982 4324
rect 3998 4380 4062 4384
rect 3998 4324 4002 4380
rect 4002 4324 4058 4380
rect 4058 4324 4062 4380
rect 3998 4320 4062 4324
rect 10474 4380 10538 4384
rect 10474 4324 10478 4380
rect 10478 4324 10534 4380
rect 10534 4324 10538 4380
rect 10474 4320 10538 4324
rect 10554 4380 10618 4384
rect 10554 4324 10558 4380
rect 10558 4324 10614 4380
rect 10614 4324 10618 4380
rect 10554 4320 10618 4324
rect 10634 4380 10698 4384
rect 10634 4324 10638 4380
rect 10638 4324 10694 4380
rect 10694 4324 10698 4380
rect 10634 4320 10698 4324
rect 10714 4380 10778 4384
rect 10714 4324 10718 4380
rect 10718 4324 10774 4380
rect 10774 4324 10778 4380
rect 10714 4320 10778 4324
rect 17190 4380 17254 4384
rect 17190 4324 17194 4380
rect 17194 4324 17250 4380
rect 17250 4324 17254 4380
rect 17190 4320 17254 4324
rect 17270 4380 17334 4384
rect 17270 4324 17274 4380
rect 17274 4324 17330 4380
rect 17330 4324 17334 4380
rect 17270 4320 17334 4324
rect 17350 4380 17414 4384
rect 17350 4324 17354 4380
rect 17354 4324 17410 4380
rect 17410 4324 17414 4380
rect 17350 4320 17414 4324
rect 17430 4380 17494 4384
rect 17430 4324 17434 4380
rect 17434 4324 17490 4380
rect 17490 4324 17494 4380
rect 17430 4320 17494 4324
rect 23906 4380 23970 4384
rect 23906 4324 23910 4380
rect 23910 4324 23966 4380
rect 23966 4324 23970 4380
rect 23906 4320 23970 4324
rect 23986 4380 24050 4384
rect 23986 4324 23990 4380
rect 23990 4324 24046 4380
rect 24046 4324 24050 4380
rect 23986 4320 24050 4324
rect 24066 4380 24130 4384
rect 24066 4324 24070 4380
rect 24070 4324 24126 4380
rect 24126 4324 24130 4380
rect 24066 4320 24130 4324
rect 24146 4380 24210 4384
rect 24146 4324 24150 4380
rect 24150 4324 24206 4380
rect 24206 4324 24210 4380
rect 24146 4320 24210 4324
rect 7116 3836 7180 3840
rect 7116 3780 7120 3836
rect 7120 3780 7176 3836
rect 7176 3780 7180 3836
rect 7116 3776 7180 3780
rect 7196 3836 7260 3840
rect 7196 3780 7200 3836
rect 7200 3780 7256 3836
rect 7256 3780 7260 3836
rect 7196 3776 7260 3780
rect 7276 3836 7340 3840
rect 7276 3780 7280 3836
rect 7280 3780 7336 3836
rect 7336 3780 7340 3836
rect 7276 3776 7340 3780
rect 7356 3836 7420 3840
rect 7356 3780 7360 3836
rect 7360 3780 7416 3836
rect 7416 3780 7420 3836
rect 7356 3776 7420 3780
rect 13832 3836 13896 3840
rect 13832 3780 13836 3836
rect 13836 3780 13892 3836
rect 13892 3780 13896 3836
rect 13832 3776 13896 3780
rect 13912 3836 13976 3840
rect 13912 3780 13916 3836
rect 13916 3780 13972 3836
rect 13972 3780 13976 3836
rect 13912 3776 13976 3780
rect 13992 3836 14056 3840
rect 13992 3780 13996 3836
rect 13996 3780 14052 3836
rect 14052 3780 14056 3836
rect 13992 3776 14056 3780
rect 14072 3836 14136 3840
rect 14072 3780 14076 3836
rect 14076 3780 14132 3836
rect 14132 3780 14136 3836
rect 14072 3776 14136 3780
rect 20548 3836 20612 3840
rect 20548 3780 20552 3836
rect 20552 3780 20608 3836
rect 20608 3780 20612 3836
rect 20548 3776 20612 3780
rect 20628 3836 20692 3840
rect 20628 3780 20632 3836
rect 20632 3780 20688 3836
rect 20688 3780 20692 3836
rect 20628 3776 20692 3780
rect 20708 3836 20772 3840
rect 20708 3780 20712 3836
rect 20712 3780 20768 3836
rect 20768 3780 20772 3836
rect 20708 3776 20772 3780
rect 20788 3836 20852 3840
rect 20788 3780 20792 3836
rect 20792 3780 20848 3836
rect 20848 3780 20852 3836
rect 20788 3776 20852 3780
rect 27264 3836 27328 3840
rect 27264 3780 27268 3836
rect 27268 3780 27324 3836
rect 27324 3780 27328 3836
rect 27264 3776 27328 3780
rect 27344 3836 27408 3840
rect 27344 3780 27348 3836
rect 27348 3780 27404 3836
rect 27404 3780 27408 3836
rect 27344 3776 27408 3780
rect 27424 3836 27488 3840
rect 27424 3780 27428 3836
rect 27428 3780 27484 3836
rect 27484 3780 27488 3836
rect 27424 3776 27488 3780
rect 27504 3836 27568 3840
rect 27504 3780 27508 3836
rect 27508 3780 27564 3836
rect 27564 3780 27568 3836
rect 27504 3776 27568 3780
rect 3758 3292 3822 3296
rect 3758 3236 3762 3292
rect 3762 3236 3818 3292
rect 3818 3236 3822 3292
rect 3758 3232 3822 3236
rect 3838 3292 3902 3296
rect 3838 3236 3842 3292
rect 3842 3236 3898 3292
rect 3898 3236 3902 3292
rect 3838 3232 3902 3236
rect 3918 3292 3982 3296
rect 3918 3236 3922 3292
rect 3922 3236 3978 3292
rect 3978 3236 3982 3292
rect 3918 3232 3982 3236
rect 3998 3292 4062 3296
rect 3998 3236 4002 3292
rect 4002 3236 4058 3292
rect 4058 3236 4062 3292
rect 3998 3232 4062 3236
rect 10474 3292 10538 3296
rect 10474 3236 10478 3292
rect 10478 3236 10534 3292
rect 10534 3236 10538 3292
rect 10474 3232 10538 3236
rect 10554 3292 10618 3296
rect 10554 3236 10558 3292
rect 10558 3236 10614 3292
rect 10614 3236 10618 3292
rect 10554 3232 10618 3236
rect 10634 3292 10698 3296
rect 10634 3236 10638 3292
rect 10638 3236 10694 3292
rect 10694 3236 10698 3292
rect 10634 3232 10698 3236
rect 10714 3292 10778 3296
rect 10714 3236 10718 3292
rect 10718 3236 10774 3292
rect 10774 3236 10778 3292
rect 10714 3232 10778 3236
rect 17190 3292 17254 3296
rect 17190 3236 17194 3292
rect 17194 3236 17250 3292
rect 17250 3236 17254 3292
rect 17190 3232 17254 3236
rect 17270 3292 17334 3296
rect 17270 3236 17274 3292
rect 17274 3236 17330 3292
rect 17330 3236 17334 3292
rect 17270 3232 17334 3236
rect 17350 3292 17414 3296
rect 17350 3236 17354 3292
rect 17354 3236 17410 3292
rect 17410 3236 17414 3292
rect 17350 3232 17414 3236
rect 17430 3292 17494 3296
rect 17430 3236 17434 3292
rect 17434 3236 17490 3292
rect 17490 3236 17494 3292
rect 17430 3232 17494 3236
rect 23906 3292 23970 3296
rect 23906 3236 23910 3292
rect 23910 3236 23966 3292
rect 23966 3236 23970 3292
rect 23906 3232 23970 3236
rect 23986 3292 24050 3296
rect 23986 3236 23990 3292
rect 23990 3236 24046 3292
rect 24046 3236 24050 3292
rect 23986 3232 24050 3236
rect 24066 3292 24130 3296
rect 24066 3236 24070 3292
rect 24070 3236 24126 3292
rect 24126 3236 24130 3292
rect 24066 3232 24130 3236
rect 24146 3292 24210 3296
rect 24146 3236 24150 3292
rect 24150 3236 24206 3292
rect 24206 3236 24210 3292
rect 24146 3232 24210 3236
rect 7116 2748 7180 2752
rect 7116 2692 7120 2748
rect 7120 2692 7176 2748
rect 7176 2692 7180 2748
rect 7116 2688 7180 2692
rect 7196 2748 7260 2752
rect 7196 2692 7200 2748
rect 7200 2692 7256 2748
rect 7256 2692 7260 2748
rect 7196 2688 7260 2692
rect 7276 2748 7340 2752
rect 7276 2692 7280 2748
rect 7280 2692 7336 2748
rect 7336 2692 7340 2748
rect 7276 2688 7340 2692
rect 7356 2748 7420 2752
rect 7356 2692 7360 2748
rect 7360 2692 7416 2748
rect 7416 2692 7420 2748
rect 7356 2688 7420 2692
rect 13832 2748 13896 2752
rect 13832 2692 13836 2748
rect 13836 2692 13892 2748
rect 13892 2692 13896 2748
rect 13832 2688 13896 2692
rect 13912 2748 13976 2752
rect 13912 2692 13916 2748
rect 13916 2692 13972 2748
rect 13972 2692 13976 2748
rect 13912 2688 13976 2692
rect 13992 2748 14056 2752
rect 13992 2692 13996 2748
rect 13996 2692 14052 2748
rect 14052 2692 14056 2748
rect 13992 2688 14056 2692
rect 14072 2748 14136 2752
rect 14072 2692 14076 2748
rect 14076 2692 14132 2748
rect 14132 2692 14136 2748
rect 14072 2688 14136 2692
rect 20548 2748 20612 2752
rect 20548 2692 20552 2748
rect 20552 2692 20608 2748
rect 20608 2692 20612 2748
rect 20548 2688 20612 2692
rect 20628 2748 20692 2752
rect 20628 2692 20632 2748
rect 20632 2692 20688 2748
rect 20688 2692 20692 2748
rect 20628 2688 20692 2692
rect 20708 2748 20772 2752
rect 20708 2692 20712 2748
rect 20712 2692 20768 2748
rect 20768 2692 20772 2748
rect 20708 2688 20772 2692
rect 20788 2748 20852 2752
rect 20788 2692 20792 2748
rect 20792 2692 20848 2748
rect 20848 2692 20852 2748
rect 20788 2688 20852 2692
rect 27264 2748 27328 2752
rect 27264 2692 27268 2748
rect 27268 2692 27324 2748
rect 27324 2692 27328 2748
rect 27264 2688 27328 2692
rect 27344 2748 27408 2752
rect 27344 2692 27348 2748
rect 27348 2692 27404 2748
rect 27404 2692 27408 2748
rect 27344 2688 27408 2692
rect 27424 2748 27488 2752
rect 27424 2692 27428 2748
rect 27428 2692 27484 2748
rect 27484 2692 27488 2748
rect 27424 2688 27488 2692
rect 27504 2748 27568 2752
rect 27504 2692 27508 2748
rect 27508 2692 27564 2748
rect 27564 2692 27568 2748
rect 27504 2688 27568 2692
rect 3758 2204 3822 2208
rect 3758 2148 3762 2204
rect 3762 2148 3818 2204
rect 3818 2148 3822 2204
rect 3758 2144 3822 2148
rect 3838 2204 3902 2208
rect 3838 2148 3842 2204
rect 3842 2148 3898 2204
rect 3898 2148 3902 2204
rect 3838 2144 3902 2148
rect 3918 2204 3982 2208
rect 3918 2148 3922 2204
rect 3922 2148 3978 2204
rect 3978 2148 3982 2204
rect 3918 2144 3982 2148
rect 3998 2204 4062 2208
rect 3998 2148 4002 2204
rect 4002 2148 4058 2204
rect 4058 2148 4062 2204
rect 3998 2144 4062 2148
rect 10474 2204 10538 2208
rect 10474 2148 10478 2204
rect 10478 2148 10534 2204
rect 10534 2148 10538 2204
rect 10474 2144 10538 2148
rect 10554 2204 10618 2208
rect 10554 2148 10558 2204
rect 10558 2148 10614 2204
rect 10614 2148 10618 2204
rect 10554 2144 10618 2148
rect 10634 2204 10698 2208
rect 10634 2148 10638 2204
rect 10638 2148 10694 2204
rect 10694 2148 10698 2204
rect 10634 2144 10698 2148
rect 10714 2204 10778 2208
rect 10714 2148 10718 2204
rect 10718 2148 10774 2204
rect 10774 2148 10778 2204
rect 10714 2144 10778 2148
rect 17190 2204 17254 2208
rect 17190 2148 17194 2204
rect 17194 2148 17250 2204
rect 17250 2148 17254 2204
rect 17190 2144 17254 2148
rect 17270 2204 17334 2208
rect 17270 2148 17274 2204
rect 17274 2148 17330 2204
rect 17330 2148 17334 2204
rect 17270 2144 17334 2148
rect 17350 2204 17414 2208
rect 17350 2148 17354 2204
rect 17354 2148 17410 2204
rect 17410 2148 17414 2204
rect 17350 2144 17414 2148
rect 17430 2204 17494 2208
rect 17430 2148 17434 2204
rect 17434 2148 17490 2204
rect 17490 2148 17494 2204
rect 17430 2144 17494 2148
rect 23906 2204 23970 2208
rect 23906 2148 23910 2204
rect 23910 2148 23966 2204
rect 23966 2148 23970 2204
rect 23906 2144 23970 2148
rect 23986 2204 24050 2208
rect 23986 2148 23990 2204
rect 23990 2148 24046 2204
rect 24046 2148 24050 2204
rect 23986 2144 24050 2148
rect 24066 2204 24130 2208
rect 24066 2148 24070 2204
rect 24070 2148 24126 2204
rect 24126 2148 24130 2204
rect 24066 2144 24130 2148
rect 24146 2204 24210 2208
rect 24146 2148 24150 2204
rect 24150 2148 24206 2204
rect 24206 2148 24210 2204
rect 24146 2144 24210 2148
rect 7116 1660 7180 1664
rect 7116 1604 7120 1660
rect 7120 1604 7176 1660
rect 7176 1604 7180 1660
rect 7116 1600 7180 1604
rect 7196 1660 7260 1664
rect 7196 1604 7200 1660
rect 7200 1604 7256 1660
rect 7256 1604 7260 1660
rect 7196 1600 7260 1604
rect 7276 1660 7340 1664
rect 7276 1604 7280 1660
rect 7280 1604 7336 1660
rect 7336 1604 7340 1660
rect 7276 1600 7340 1604
rect 7356 1660 7420 1664
rect 7356 1604 7360 1660
rect 7360 1604 7416 1660
rect 7416 1604 7420 1660
rect 7356 1600 7420 1604
rect 13832 1660 13896 1664
rect 13832 1604 13836 1660
rect 13836 1604 13892 1660
rect 13892 1604 13896 1660
rect 13832 1600 13896 1604
rect 13912 1660 13976 1664
rect 13912 1604 13916 1660
rect 13916 1604 13972 1660
rect 13972 1604 13976 1660
rect 13912 1600 13976 1604
rect 13992 1660 14056 1664
rect 13992 1604 13996 1660
rect 13996 1604 14052 1660
rect 14052 1604 14056 1660
rect 13992 1600 14056 1604
rect 14072 1660 14136 1664
rect 14072 1604 14076 1660
rect 14076 1604 14132 1660
rect 14132 1604 14136 1660
rect 14072 1600 14136 1604
rect 20548 1660 20612 1664
rect 20548 1604 20552 1660
rect 20552 1604 20608 1660
rect 20608 1604 20612 1660
rect 20548 1600 20612 1604
rect 20628 1660 20692 1664
rect 20628 1604 20632 1660
rect 20632 1604 20688 1660
rect 20688 1604 20692 1660
rect 20628 1600 20692 1604
rect 20708 1660 20772 1664
rect 20708 1604 20712 1660
rect 20712 1604 20768 1660
rect 20768 1604 20772 1660
rect 20708 1600 20772 1604
rect 20788 1660 20852 1664
rect 20788 1604 20792 1660
rect 20792 1604 20848 1660
rect 20848 1604 20852 1660
rect 20788 1600 20852 1604
rect 27264 1660 27328 1664
rect 27264 1604 27268 1660
rect 27268 1604 27324 1660
rect 27324 1604 27328 1660
rect 27264 1600 27328 1604
rect 27344 1660 27408 1664
rect 27344 1604 27348 1660
rect 27348 1604 27404 1660
rect 27404 1604 27408 1660
rect 27344 1600 27408 1604
rect 27424 1660 27488 1664
rect 27424 1604 27428 1660
rect 27428 1604 27484 1660
rect 27484 1604 27488 1660
rect 27424 1600 27488 1604
rect 27504 1660 27568 1664
rect 27504 1604 27508 1660
rect 27508 1604 27564 1660
rect 27564 1604 27568 1660
rect 27504 1600 27568 1604
rect 3758 1116 3822 1120
rect 3758 1060 3762 1116
rect 3762 1060 3818 1116
rect 3818 1060 3822 1116
rect 3758 1056 3822 1060
rect 3838 1116 3902 1120
rect 3838 1060 3842 1116
rect 3842 1060 3898 1116
rect 3898 1060 3902 1116
rect 3838 1056 3902 1060
rect 3918 1116 3982 1120
rect 3918 1060 3922 1116
rect 3922 1060 3978 1116
rect 3978 1060 3982 1116
rect 3918 1056 3982 1060
rect 3998 1116 4062 1120
rect 3998 1060 4002 1116
rect 4002 1060 4058 1116
rect 4058 1060 4062 1116
rect 3998 1056 4062 1060
rect 10474 1116 10538 1120
rect 10474 1060 10478 1116
rect 10478 1060 10534 1116
rect 10534 1060 10538 1116
rect 10474 1056 10538 1060
rect 10554 1116 10618 1120
rect 10554 1060 10558 1116
rect 10558 1060 10614 1116
rect 10614 1060 10618 1116
rect 10554 1056 10618 1060
rect 10634 1116 10698 1120
rect 10634 1060 10638 1116
rect 10638 1060 10694 1116
rect 10694 1060 10698 1116
rect 10634 1056 10698 1060
rect 10714 1116 10778 1120
rect 10714 1060 10718 1116
rect 10718 1060 10774 1116
rect 10774 1060 10778 1116
rect 10714 1056 10778 1060
rect 17190 1116 17254 1120
rect 17190 1060 17194 1116
rect 17194 1060 17250 1116
rect 17250 1060 17254 1116
rect 17190 1056 17254 1060
rect 17270 1116 17334 1120
rect 17270 1060 17274 1116
rect 17274 1060 17330 1116
rect 17330 1060 17334 1116
rect 17270 1056 17334 1060
rect 17350 1116 17414 1120
rect 17350 1060 17354 1116
rect 17354 1060 17410 1116
rect 17410 1060 17414 1116
rect 17350 1056 17414 1060
rect 17430 1116 17494 1120
rect 17430 1060 17434 1116
rect 17434 1060 17490 1116
rect 17490 1060 17494 1116
rect 17430 1056 17494 1060
rect 23906 1116 23970 1120
rect 23906 1060 23910 1116
rect 23910 1060 23966 1116
rect 23966 1060 23970 1116
rect 23906 1056 23970 1060
rect 23986 1116 24050 1120
rect 23986 1060 23990 1116
rect 23990 1060 24046 1116
rect 24046 1060 24050 1116
rect 23986 1056 24050 1060
rect 24066 1116 24130 1120
rect 24066 1060 24070 1116
rect 24070 1060 24126 1116
rect 24126 1060 24130 1116
rect 24066 1056 24130 1060
rect 24146 1116 24210 1120
rect 24146 1060 24150 1116
rect 24150 1060 24206 1116
rect 24206 1060 24210 1116
rect 24146 1056 24210 1060
rect 7116 572 7180 576
rect 7116 516 7120 572
rect 7120 516 7176 572
rect 7176 516 7180 572
rect 7116 512 7180 516
rect 7196 572 7260 576
rect 7196 516 7200 572
rect 7200 516 7256 572
rect 7256 516 7260 572
rect 7196 512 7260 516
rect 7276 572 7340 576
rect 7276 516 7280 572
rect 7280 516 7336 572
rect 7336 516 7340 572
rect 7276 512 7340 516
rect 7356 572 7420 576
rect 7356 516 7360 572
rect 7360 516 7416 572
rect 7416 516 7420 572
rect 7356 512 7420 516
rect 13832 572 13896 576
rect 13832 516 13836 572
rect 13836 516 13892 572
rect 13892 516 13896 572
rect 13832 512 13896 516
rect 13912 572 13976 576
rect 13912 516 13916 572
rect 13916 516 13972 572
rect 13972 516 13976 572
rect 13912 512 13976 516
rect 13992 572 14056 576
rect 13992 516 13996 572
rect 13996 516 14052 572
rect 14052 516 14056 572
rect 13992 512 14056 516
rect 14072 572 14136 576
rect 14072 516 14076 572
rect 14076 516 14132 572
rect 14132 516 14136 572
rect 14072 512 14136 516
rect 20548 572 20612 576
rect 20548 516 20552 572
rect 20552 516 20608 572
rect 20608 516 20612 572
rect 20548 512 20612 516
rect 20628 572 20692 576
rect 20628 516 20632 572
rect 20632 516 20688 572
rect 20688 516 20692 572
rect 20628 512 20692 516
rect 20708 572 20772 576
rect 20708 516 20712 572
rect 20712 516 20768 572
rect 20768 516 20772 572
rect 20708 512 20772 516
rect 20788 572 20852 576
rect 20788 516 20792 572
rect 20792 516 20848 572
rect 20848 516 20852 572
rect 20788 512 20852 516
rect 27264 572 27328 576
rect 27264 516 27268 572
rect 27268 516 27324 572
rect 27324 516 27328 572
rect 27264 512 27328 516
rect 27344 572 27408 576
rect 27344 516 27348 572
rect 27348 516 27404 572
rect 27404 516 27408 572
rect 27344 512 27408 516
rect 27424 572 27488 576
rect 27424 516 27428 572
rect 27428 516 27484 572
rect 27484 516 27488 572
rect 27424 512 27488 516
rect 27504 572 27568 576
rect 27504 516 27508 572
rect 27508 516 27564 572
rect 27564 516 27568 572
rect 27504 512 27568 516
<< metal4 >>
rect 3750 30496 4070 31056
rect 3750 30432 3758 30496
rect 3822 30432 3838 30496
rect 3902 30432 3918 30496
rect 3982 30432 3998 30496
rect 4062 30432 4070 30496
rect 2083 30428 2149 30429
rect 2083 30364 2084 30428
rect 2148 30364 2149 30428
rect 2083 30363 2149 30364
rect 1899 29748 1965 29749
rect 1899 29684 1900 29748
rect 1964 29684 1965 29748
rect 1899 29683 1965 29684
rect 1902 7309 1962 29683
rect 2086 10573 2146 30363
rect 3750 29408 4070 30432
rect 3750 29344 3758 29408
rect 3822 29344 3838 29408
rect 3902 29344 3918 29408
rect 3982 29344 3998 29408
rect 4062 29344 4070 29408
rect 3750 28320 4070 29344
rect 3750 28256 3758 28320
rect 3822 28256 3838 28320
rect 3902 28256 3918 28320
rect 3982 28256 3998 28320
rect 4062 28256 4070 28320
rect 3750 27232 4070 28256
rect 3750 27168 3758 27232
rect 3822 27168 3838 27232
rect 3902 27168 3918 27232
rect 3982 27168 3998 27232
rect 4062 27168 4070 27232
rect 3750 26144 4070 27168
rect 3750 26080 3758 26144
rect 3822 26080 3838 26144
rect 3902 26080 3918 26144
rect 3982 26080 3998 26144
rect 4062 26080 4070 26144
rect 3750 25056 4070 26080
rect 3750 24992 3758 25056
rect 3822 24992 3838 25056
rect 3902 24992 3918 25056
rect 3982 24992 3998 25056
rect 4062 24992 4070 25056
rect 3750 23968 4070 24992
rect 3750 23904 3758 23968
rect 3822 23904 3838 23968
rect 3902 23904 3918 23968
rect 3982 23904 3998 23968
rect 4062 23904 4070 23968
rect 3750 22880 4070 23904
rect 3750 22816 3758 22880
rect 3822 22816 3838 22880
rect 3902 22816 3918 22880
rect 3982 22816 3998 22880
rect 4062 22816 4070 22880
rect 3750 21792 4070 22816
rect 3750 21728 3758 21792
rect 3822 21728 3838 21792
rect 3902 21728 3918 21792
rect 3982 21728 3998 21792
rect 4062 21728 4070 21792
rect 3750 20704 4070 21728
rect 3750 20640 3758 20704
rect 3822 20640 3838 20704
rect 3902 20640 3918 20704
rect 3982 20640 3998 20704
rect 4062 20640 4070 20704
rect 3750 19616 4070 20640
rect 3750 19552 3758 19616
rect 3822 19552 3838 19616
rect 3902 19552 3918 19616
rect 3982 19552 3998 19616
rect 4062 19552 4070 19616
rect 3750 18528 4070 19552
rect 3750 18464 3758 18528
rect 3822 18464 3838 18528
rect 3902 18464 3918 18528
rect 3982 18464 3998 18528
rect 4062 18464 4070 18528
rect 3750 17440 4070 18464
rect 3750 17376 3758 17440
rect 3822 17376 3838 17440
rect 3902 17376 3918 17440
rect 3982 17376 3998 17440
rect 4062 17376 4070 17440
rect 3750 16352 4070 17376
rect 3750 16288 3758 16352
rect 3822 16288 3838 16352
rect 3902 16288 3918 16352
rect 3982 16288 3998 16352
rect 4062 16288 4070 16352
rect 3750 15264 4070 16288
rect 3750 15200 3758 15264
rect 3822 15200 3838 15264
rect 3902 15200 3918 15264
rect 3982 15200 3998 15264
rect 4062 15200 4070 15264
rect 3750 14176 4070 15200
rect 3750 14112 3758 14176
rect 3822 14112 3838 14176
rect 3902 14112 3918 14176
rect 3982 14112 3998 14176
rect 4062 14112 4070 14176
rect 3750 13088 4070 14112
rect 3750 13024 3758 13088
rect 3822 13024 3838 13088
rect 3902 13024 3918 13088
rect 3982 13024 3998 13088
rect 4062 13024 4070 13088
rect 3750 12000 4070 13024
rect 3750 11936 3758 12000
rect 3822 11936 3838 12000
rect 3902 11936 3918 12000
rect 3982 11936 3998 12000
rect 4062 11936 4070 12000
rect 3750 10912 4070 11936
rect 3750 10848 3758 10912
rect 3822 10848 3838 10912
rect 3902 10848 3918 10912
rect 3982 10848 3998 10912
rect 4062 10848 4070 10912
rect 2083 10572 2149 10573
rect 2083 10508 2084 10572
rect 2148 10508 2149 10572
rect 2083 10507 2149 10508
rect 3750 9824 4070 10848
rect 3750 9760 3758 9824
rect 3822 9760 3838 9824
rect 3902 9760 3918 9824
rect 3982 9760 3998 9824
rect 4062 9760 4070 9824
rect 3750 8736 4070 9760
rect 3750 8672 3758 8736
rect 3822 8672 3838 8736
rect 3902 8672 3918 8736
rect 3982 8672 3998 8736
rect 4062 8672 4070 8736
rect 3750 7648 4070 8672
rect 3750 7584 3758 7648
rect 3822 7584 3838 7648
rect 3902 7584 3918 7648
rect 3982 7584 3998 7648
rect 4062 7584 4070 7648
rect 1899 7308 1965 7309
rect 1899 7244 1900 7308
rect 1964 7244 1965 7308
rect 1899 7243 1965 7244
rect 3750 6560 4070 7584
rect 3750 6496 3758 6560
rect 3822 6496 3838 6560
rect 3902 6496 3918 6560
rect 3982 6496 3998 6560
rect 4062 6496 4070 6560
rect 3750 5472 4070 6496
rect 3750 5408 3758 5472
rect 3822 5408 3838 5472
rect 3902 5408 3918 5472
rect 3982 5408 3998 5472
rect 4062 5408 4070 5472
rect 3750 4384 4070 5408
rect 3750 4320 3758 4384
rect 3822 4320 3838 4384
rect 3902 4320 3918 4384
rect 3982 4320 3998 4384
rect 4062 4320 4070 4384
rect 3750 3296 4070 4320
rect 3750 3232 3758 3296
rect 3822 3232 3838 3296
rect 3902 3232 3918 3296
rect 3982 3232 3998 3296
rect 4062 3232 4070 3296
rect 3750 2208 4070 3232
rect 3750 2144 3758 2208
rect 3822 2144 3838 2208
rect 3902 2144 3918 2208
rect 3982 2144 3998 2208
rect 4062 2144 4070 2208
rect 3750 1120 4070 2144
rect 3750 1056 3758 1120
rect 3822 1056 3838 1120
rect 3902 1056 3918 1120
rect 3982 1056 3998 1120
rect 4062 1056 4070 1120
rect 3750 496 4070 1056
rect 7108 31040 7428 31056
rect 7108 30976 7116 31040
rect 7180 30976 7196 31040
rect 7260 30976 7276 31040
rect 7340 30976 7356 31040
rect 7420 30976 7428 31040
rect 7108 29952 7428 30976
rect 7108 29888 7116 29952
rect 7180 29888 7196 29952
rect 7260 29888 7276 29952
rect 7340 29888 7356 29952
rect 7420 29888 7428 29952
rect 7108 28864 7428 29888
rect 7108 28800 7116 28864
rect 7180 28800 7196 28864
rect 7260 28800 7276 28864
rect 7340 28800 7356 28864
rect 7420 28800 7428 28864
rect 7108 27776 7428 28800
rect 7108 27712 7116 27776
rect 7180 27712 7196 27776
rect 7260 27712 7276 27776
rect 7340 27712 7356 27776
rect 7420 27712 7428 27776
rect 7108 26688 7428 27712
rect 7108 26624 7116 26688
rect 7180 26624 7196 26688
rect 7260 26624 7276 26688
rect 7340 26624 7356 26688
rect 7420 26624 7428 26688
rect 7108 25600 7428 26624
rect 7108 25536 7116 25600
rect 7180 25536 7196 25600
rect 7260 25536 7276 25600
rect 7340 25536 7356 25600
rect 7420 25536 7428 25600
rect 7108 24512 7428 25536
rect 7108 24448 7116 24512
rect 7180 24448 7196 24512
rect 7260 24448 7276 24512
rect 7340 24448 7356 24512
rect 7420 24448 7428 24512
rect 7108 23424 7428 24448
rect 7108 23360 7116 23424
rect 7180 23360 7196 23424
rect 7260 23360 7276 23424
rect 7340 23360 7356 23424
rect 7420 23360 7428 23424
rect 7108 22336 7428 23360
rect 7108 22272 7116 22336
rect 7180 22272 7196 22336
rect 7260 22272 7276 22336
rect 7340 22272 7356 22336
rect 7420 22272 7428 22336
rect 7108 21248 7428 22272
rect 7108 21184 7116 21248
rect 7180 21184 7196 21248
rect 7260 21184 7276 21248
rect 7340 21184 7356 21248
rect 7420 21184 7428 21248
rect 7108 20160 7428 21184
rect 7108 20096 7116 20160
rect 7180 20096 7196 20160
rect 7260 20096 7276 20160
rect 7340 20096 7356 20160
rect 7420 20096 7428 20160
rect 7108 19072 7428 20096
rect 7108 19008 7116 19072
rect 7180 19008 7196 19072
rect 7260 19008 7276 19072
rect 7340 19008 7356 19072
rect 7420 19008 7428 19072
rect 7108 17984 7428 19008
rect 7108 17920 7116 17984
rect 7180 17920 7196 17984
rect 7260 17920 7276 17984
rect 7340 17920 7356 17984
rect 7420 17920 7428 17984
rect 7108 16896 7428 17920
rect 7108 16832 7116 16896
rect 7180 16832 7196 16896
rect 7260 16832 7276 16896
rect 7340 16832 7356 16896
rect 7420 16832 7428 16896
rect 7108 15808 7428 16832
rect 7108 15744 7116 15808
rect 7180 15744 7196 15808
rect 7260 15744 7276 15808
rect 7340 15744 7356 15808
rect 7420 15744 7428 15808
rect 7108 14720 7428 15744
rect 7108 14656 7116 14720
rect 7180 14656 7196 14720
rect 7260 14656 7276 14720
rect 7340 14656 7356 14720
rect 7420 14656 7428 14720
rect 7108 13632 7428 14656
rect 7108 13568 7116 13632
rect 7180 13568 7196 13632
rect 7260 13568 7276 13632
rect 7340 13568 7356 13632
rect 7420 13568 7428 13632
rect 7108 12544 7428 13568
rect 7108 12480 7116 12544
rect 7180 12480 7196 12544
rect 7260 12480 7276 12544
rect 7340 12480 7356 12544
rect 7420 12480 7428 12544
rect 7108 11456 7428 12480
rect 7108 11392 7116 11456
rect 7180 11392 7196 11456
rect 7260 11392 7276 11456
rect 7340 11392 7356 11456
rect 7420 11392 7428 11456
rect 7108 10368 7428 11392
rect 7108 10304 7116 10368
rect 7180 10304 7196 10368
rect 7260 10304 7276 10368
rect 7340 10304 7356 10368
rect 7420 10304 7428 10368
rect 7108 9280 7428 10304
rect 7108 9216 7116 9280
rect 7180 9216 7196 9280
rect 7260 9216 7276 9280
rect 7340 9216 7356 9280
rect 7420 9216 7428 9280
rect 7108 8192 7428 9216
rect 7108 8128 7116 8192
rect 7180 8128 7196 8192
rect 7260 8128 7276 8192
rect 7340 8128 7356 8192
rect 7420 8128 7428 8192
rect 7108 7104 7428 8128
rect 7108 7040 7116 7104
rect 7180 7040 7196 7104
rect 7260 7040 7276 7104
rect 7340 7040 7356 7104
rect 7420 7040 7428 7104
rect 7108 6016 7428 7040
rect 7108 5952 7116 6016
rect 7180 5952 7196 6016
rect 7260 5952 7276 6016
rect 7340 5952 7356 6016
rect 7420 5952 7428 6016
rect 7108 4928 7428 5952
rect 7108 4864 7116 4928
rect 7180 4864 7196 4928
rect 7260 4864 7276 4928
rect 7340 4864 7356 4928
rect 7420 4864 7428 4928
rect 7108 3840 7428 4864
rect 7108 3776 7116 3840
rect 7180 3776 7196 3840
rect 7260 3776 7276 3840
rect 7340 3776 7356 3840
rect 7420 3776 7428 3840
rect 7108 2752 7428 3776
rect 7108 2688 7116 2752
rect 7180 2688 7196 2752
rect 7260 2688 7276 2752
rect 7340 2688 7356 2752
rect 7420 2688 7428 2752
rect 7108 1664 7428 2688
rect 7108 1600 7116 1664
rect 7180 1600 7196 1664
rect 7260 1600 7276 1664
rect 7340 1600 7356 1664
rect 7420 1600 7428 1664
rect 7108 576 7428 1600
rect 7108 512 7116 576
rect 7180 512 7196 576
rect 7260 512 7276 576
rect 7340 512 7356 576
rect 7420 512 7428 576
rect 7108 496 7428 512
rect 10466 30496 10786 31056
rect 10466 30432 10474 30496
rect 10538 30432 10554 30496
rect 10618 30432 10634 30496
rect 10698 30432 10714 30496
rect 10778 30432 10786 30496
rect 10466 29408 10786 30432
rect 10466 29344 10474 29408
rect 10538 29344 10554 29408
rect 10618 29344 10634 29408
rect 10698 29344 10714 29408
rect 10778 29344 10786 29408
rect 10466 28320 10786 29344
rect 10466 28256 10474 28320
rect 10538 28256 10554 28320
rect 10618 28256 10634 28320
rect 10698 28256 10714 28320
rect 10778 28256 10786 28320
rect 10466 27232 10786 28256
rect 10466 27168 10474 27232
rect 10538 27168 10554 27232
rect 10618 27168 10634 27232
rect 10698 27168 10714 27232
rect 10778 27168 10786 27232
rect 10466 26144 10786 27168
rect 10466 26080 10474 26144
rect 10538 26080 10554 26144
rect 10618 26080 10634 26144
rect 10698 26080 10714 26144
rect 10778 26080 10786 26144
rect 10466 25056 10786 26080
rect 10466 24992 10474 25056
rect 10538 24992 10554 25056
rect 10618 24992 10634 25056
rect 10698 24992 10714 25056
rect 10778 24992 10786 25056
rect 10466 23968 10786 24992
rect 10466 23904 10474 23968
rect 10538 23904 10554 23968
rect 10618 23904 10634 23968
rect 10698 23904 10714 23968
rect 10778 23904 10786 23968
rect 10466 22880 10786 23904
rect 10466 22816 10474 22880
rect 10538 22816 10554 22880
rect 10618 22816 10634 22880
rect 10698 22816 10714 22880
rect 10778 22816 10786 22880
rect 10466 21792 10786 22816
rect 10466 21728 10474 21792
rect 10538 21728 10554 21792
rect 10618 21728 10634 21792
rect 10698 21728 10714 21792
rect 10778 21728 10786 21792
rect 10466 20704 10786 21728
rect 10466 20640 10474 20704
rect 10538 20640 10554 20704
rect 10618 20640 10634 20704
rect 10698 20640 10714 20704
rect 10778 20640 10786 20704
rect 10466 19616 10786 20640
rect 10466 19552 10474 19616
rect 10538 19552 10554 19616
rect 10618 19552 10634 19616
rect 10698 19552 10714 19616
rect 10778 19552 10786 19616
rect 10466 18528 10786 19552
rect 10466 18464 10474 18528
rect 10538 18464 10554 18528
rect 10618 18464 10634 18528
rect 10698 18464 10714 18528
rect 10778 18464 10786 18528
rect 10466 17440 10786 18464
rect 10466 17376 10474 17440
rect 10538 17376 10554 17440
rect 10618 17376 10634 17440
rect 10698 17376 10714 17440
rect 10778 17376 10786 17440
rect 10466 16352 10786 17376
rect 10466 16288 10474 16352
rect 10538 16288 10554 16352
rect 10618 16288 10634 16352
rect 10698 16288 10714 16352
rect 10778 16288 10786 16352
rect 10466 15264 10786 16288
rect 10466 15200 10474 15264
rect 10538 15200 10554 15264
rect 10618 15200 10634 15264
rect 10698 15200 10714 15264
rect 10778 15200 10786 15264
rect 10466 14176 10786 15200
rect 10466 14112 10474 14176
rect 10538 14112 10554 14176
rect 10618 14112 10634 14176
rect 10698 14112 10714 14176
rect 10778 14112 10786 14176
rect 10466 13088 10786 14112
rect 10466 13024 10474 13088
rect 10538 13024 10554 13088
rect 10618 13024 10634 13088
rect 10698 13024 10714 13088
rect 10778 13024 10786 13088
rect 10466 12000 10786 13024
rect 10466 11936 10474 12000
rect 10538 11936 10554 12000
rect 10618 11936 10634 12000
rect 10698 11936 10714 12000
rect 10778 11936 10786 12000
rect 10466 10912 10786 11936
rect 10466 10848 10474 10912
rect 10538 10848 10554 10912
rect 10618 10848 10634 10912
rect 10698 10848 10714 10912
rect 10778 10848 10786 10912
rect 10466 9824 10786 10848
rect 10466 9760 10474 9824
rect 10538 9760 10554 9824
rect 10618 9760 10634 9824
rect 10698 9760 10714 9824
rect 10778 9760 10786 9824
rect 10466 8736 10786 9760
rect 10466 8672 10474 8736
rect 10538 8672 10554 8736
rect 10618 8672 10634 8736
rect 10698 8672 10714 8736
rect 10778 8672 10786 8736
rect 10466 7648 10786 8672
rect 10466 7584 10474 7648
rect 10538 7584 10554 7648
rect 10618 7584 10634 7648
rect 10698 7584 10714 7648
rect 10778 7584 10786 7648
rect 10466 6560 10786 7584
rect 10466 6496 10474 6560
rect 10538 6496 10554 6560
rect 10618 6496 10634 6560
rect 10698 6496 10714 6560
rect 10778 6496 10786 6560
rect 10466 5472 10786 6496
rect 10466 5408 10474 5472
rect 10538 5408 10554 5472
rect 10618 5408 10634 5472
rect 10698 5408 10714 5472
rect 10778 5408 10786 5472
rect 10466 4384 10786 5408
rect 10466 4320 10474 4384
rect 10538 4320 10554 4384
rect 10618 4320 10634 4384
rect 10698 4320 10714 4384
rect 10778 4320 10786 4384
rect 10466 3296 10786 4320
rect 10466 3232 10474 3296
rect 10538 3232 10554 3296
rect 10618 3232 10634 3296
rect 10698 3232 10714 3296
rect 10778 3232 10786 3296
rect 10466 2208 10786 3232
rect 10466 2144 10474 2208
rect 10538 2144 10554 2208
rect 10618 2144 10634 2208
rect 10698 2144 10714 2208
rect 10778 2144 10786 2208
rect 10466 1120 10786 2144
rect 10466 1056 10474 1120
rect 10538 1056 10554 1120
rect 10618 1056 10634 1120
rect 10698 1056 10714 1120
rect 10778 1056 10786 1120
rect 10466 496 10786 1056
rect 13824 31040 14144 31056
rect 13824 30976 13832 31040
rect 13896 30976 13912 31040
rect 13976 30976 13992 31040
rect 14056 30976 14072 31040
rect 14136 30976 14144 31040
rect 13824 29952 14144 30976
rect 13824 29888 13832 29952
rect 13896 29888 13912 29952
rect 13976 29888 13992 29952
rect 14056 29888 14072 29952
rect 14136 29888 14144 29952
rect 13824 28864 14144 29888
rect 13824 28800 13832 28864
rect 13896 28800 13912 28864
rect 13976 28800 13992 28864
rect 14056 28800 14072 28864
rect 14136 28800 14144 28864
rect 13824 27776 14144 28800
rect 13824 27712 13832 27776
rect 13896 27712 13912 27776
rect 13976 27712 13992 27776
rect 14056 27712 14072 27776
rect 14136 27712 14144 27776
rect 13824 26688 14144 27712
rect 13824 26624 13832 26688
rect 13896 26624 13912 26688
rect 13976 26624 13992 26688
rect 14056 26624 14072 26688
rect 14136 26624 14144 26688
rect 13824 25600 14144 26624
rect 13824 25536 13832 25600
rect 13896 25536 13912 25600
rect 13976 25536 13992 25600
rect 14056 25536 14072 25600
rect 14136 25536 14144 25600
rect 13824 24512 14144 25536
rect 13824 24448 13832 24512
rect 13896 24448 13912 24512
rect 13976 24448 13992 24512
rect 14056 24448 14072 24512
rect 14136 24448 14144 24512
rect 13824 23424 14144 24448
rect 13824 23360 13832 23424
rect 13896 23360 13912 23424
rect 13976 23360 13992 23424
rect 14056 23360 14072 23424
rect 14136 23360 14144 23424
rect 13824 22336 14144 23360
rect 13824 22272 13832 22336
rect 13896 22272 13912 22336
rect 13976 22272 13992 22336
rect 14056 22272 14072 22336
rect 14136 22272 14144 22336
rect 13824 21248 14144 22272
rect 13824 21184 13832 21248
rect 13896 21184 13912 21248
rect 13976 21184 13992 21248
rect 14056 21184 14072 21248
rect 14136 21184 14144 21248
rect 13824 20160 14144 21184
rect 13824 20096 13832 20160
rect 13896 20096 13912 20160
rect 13976 20096 13992 20160
rect 14056 20096 14072 20160
rect 14136 20096 14144 20160
rect 13824 19072 14144 20096
rect 13824 19008 13832 19072
rect 13896 19008 13912 19072
rect 13976 19008 13992 19072
rect 14056 19008 14072 19072
rect 14136 19008 14144 19072
rect 13824 17984 14144 19008
rect 13824 17920 13832 17984
rect 13896 17920 13912 17984
rect 13976 17920 13992 17984
rect 14056 17920 14072 17984
rect 14136 17920 14144 17984
rect 13824 16896 14144 17920
rect 13824 16832 13832 16896
rect 13896 16832 13912 16896
rect 13976 16832 13992 16896
rect 14056 16832 14072 16896
rect 14136 16832 14144 16896
rect 13824 15808 14144 16832
rect 13824 15744 13832 15808
rect 13896 15744 13912 15808
rect 13976 15744 13992 15808
rect 14056 15744 14072 15808
rect 14136 15744 14144 15808
rect 13824 14720 14144 15744
rect 13824 14656 13832 14720
rect 13896 14656 13912 14720
rect 13976 14656 13992 14720
rect 14056 14656 14072 14720
rect 14136 14656 14144 14720
rect 13824 13632 14144 14656
rect 13824 13568 13832 13632
rect 13896 13568 13912 13632
rect 13976 13568 13992 13632
rect 14056 13568 14072 13632
rect 14136 13568 14144 13632
rect 13824 12544 14144 13568
rect 13824 12480 13832 12544
rect 13896 12480 13912 12544
rect 13976 12480 13992 12544
rect 14056 12480 14072 12544
rect 14136 12480 14144 12544
rect 13824 11456 14144 12480
rect 13824 11392 13832 11456
rect 13896 11392 13912 11456
rect 13976 11392 13992 11456
rect 14056 11392 14072 11456
rect 14136 11392 14144 11456
rect 13824 10368 14144 11392
rect 13824 10304 13832 10368
rect 13896 10304 13912 10368
rect 13976 10304 13992 10368
rect 14056 10304 14072 10368
rect 14136 10304 14144 10368
rect 13824 9280 14144 10304
rect 13824 9216 13832 9280
rect 13896 9216 13912 9280
rect 13976 9216 13992 9280
rect 14056 9216 14072 9280
rect 14136 9216 14144 9280
rect 13824 8192 14144 9216
rect 13824 8128 13832 8192
rect 13896 8128 13912 8192
rect 13976 8128 13992 8192
rect 14056 8128 14072 8192
rect 14136 8128 14144 8192
rect 13824 7104 14144 8128
rect 13824 7040 13832 7104
rect 13896 7040 13912 7104
rect 13976 7040 13992 7104
rect 14056 7040 14072 7104
rect 14136 7040 14144 7104
rect 13824 6016 14144 7040
rect 13824 5952 13832 6016
rect 13896 5952 13912 6016
rect 13976 5952 13992 6016
rect 14056 5952 14072 6016
rect 14136 5952 14144 6016
rect 13824 4928 14144 5952
rect 13824 4864 13832 4928
rect 13896 4864 13912 4928
rect 13976 4864 13992 4928
rect 14056 4864 14072 4928
rect 14136 4864 14144 4928
rect 13824 3840 14144 4864
rect 13824 3776 13832 3840
rect 13896 3776 13912 3840
rect 13976 3776 13992 3840
rect 14056 3776 14072 3840
rect 14136 3776 14144 3840
rect 13824 2752 14144 3776
rect 13824 2688 13832 2752
rect 13896 2688 13912 2752
rect 13976 2688 13992 2752
rect 14056 2688 14072 2752
rect 14136 2688 14144 2752
rect 13824 1664 14144 2688
rect 13824 1600 13832 1664
rect 13896 1600 13912 1664
rect 13976 1600 13992 1664
rect 14056 1600 14072 1664
rect 14136 1600 14144 1664
rect 13824 576 14144 1600
rect 13824 512 13832 576
rect 13896 512 13912 576
rect 13976 512 13992 576
rect 14056 512 14072 576
rect 14136 512 14144 576
rect 13824 496 14144 512
rect 17182 30496 17502 31056
rect 17182 30432 17190 30496
rect 17254 30432 17270 30496
rect 17334 30432 17350 30496
rect 17414 30432 17430 30496
rect 17494 30432 17502 30496
rect 17182 29408 17502 30432
rect 17182 29344 17190 29408
rect 17254 29344 17270 29408
rect 17334 29344 17350 29408
rect 17414 29344 17430 29408
rect 17494 29344 17502 29408
rect 17182 28320 17502 29344
rect 17182 28256 17190 28320
rect 17254 28256 17270 28320
rect 17334 28256 17350 28320
rect 17414 28256 17430 28320
rect 17494 28256 17502 28320
rect 17182 27232 17502 28256
rect 17182 27168 17190 27232
rect 17254 27168 17270 27232
rect 17334 27168 17350 27232
rect 17414 27168 17430 27232
rect 17494 27168 17502 27232
rect 17182 26144 17502 27168
rect 17182 26080 17190 26144
rect 17254 26080 17270 26144
rect 17334 26080 17350 26144
rect 17414 26080 17430 26144
rect 17494 26080 17502 26144
rect 17182 25056 17502 26080
rect 17182 24992 17190 25056
rect 17254 24992 17270 25056
rect 17334 24992 17350 25056
rect 17414 24992 17430 25056
rect 17494 24992 17502 25056
rect 17182 23968 17502 24992
rect 17182 23904 17190 23968
rect 17254 23904 17270 23968
rect 17334 23904 17350 23968
rect 17414 23904 17430 23968
rect 17494 23904 17502 23968
rect 17182 22880 17502 23904
rect 17182 22816 17190 22880
rect 17254 22816 17270 22880
rect 17334 22816 17350 22880
rect 17414 22816 17430 22880
rect 17494 22816 17502 22880
rect 17182 21792 17502 22816
rect 17182 21728 17190 21792
rect 17254 21728 17270 21792
rect 17334 21728 17350 21792
rect 17414 21728 17430 21792
rect 17494 21728 17502 21792
rect 17182 20704 17502 21728
rect 17182 20640 17190 20704
rect 17254 20640 17270 20704
rect 17334 20640 17350 20704
rect 17414 20640 17430 20704
rect 17494 20640 17502 20704
rect 17182 19616 17502 20640
rect 17182 19552 17190 19616
rect 17254 19552 17270 19616
rect 17334 19552 17350 19616
rect 17414 19552 17430 19616
rect 17494 19552 17502 19616
rect 17182 18528 17502 19552
rect 17182 18464 17190 18528
rect 17254 18464 17270 18528
rect 17334 18464 17350 18528
rect 17414 18464 17430 18528
rect 17494 18464 17502 18528
rect 17182 17440 17502 18464
rect 17182 17376 17190 17440
rect 17254 17376 17270 17440
rect 17334 17376 17350 17440
rect 17414 17376 17430 17440
rect 17494 17376 17502 17440
rect 17182 16352 17502 17376
rect 17182 16288 17190 16352
rect 17254 16288 17270 16352
rect 17334 16288 17350 16352
rect 17414 16288 17430 16352
rect 17494 16288 17502 16352
rect 17182 15264 17502 16288
rect 17182 15200 17190 15264
rect 17254 15200 17270 15264
rect 17334 15200 17350 15264
rect 17414 15200 17430 15264
rect 17494 15200 17502 15264
rect 17182 14176 17502 15200
rect 17182 14112 17190 14176
rect 17254 14112 17270 14176
rect 17334 14112 17350 14176
rect 17414 14112 17430 14176
rect 17494 14112 17502 14176
rect 17182 13088 17502 14112
rect 17182 13024 17190 13088
rect 17254 13024 17270 13088
rect 17334 13024 17350 13088
rect 17414 13024 17430 13088
rect 17494 13024 17502 13088
rect 17182 12000 17502 13024
rect 17182 11936 17190 12000
rect 17254 11936 17270 12000
rect 17334 11936 17350 12000
rect 17414 11936 17430 12000
rect 17494 11936 17502 12000
rect 17182 10912 17502 11936
rect 17182 10848 17190 10912
rect 17254 10848 17270 10912
rect 17334 10848 17350 10912
rect 17414 10848 17430 10912
rect 17494 10848 17502 10912
rect 17182 9824 17502 10848
rect 17182 9760 17190 9824
rect 17254 9760 17270 9824
rect 17334 9760 17350 9824
rect 17414 9760 17430 9824
rect 17494 9760 17502 9824
rect 17182 8736 17502 9760
rect 17182 8672 17190 8736
rect 17254 8672 17270 8736
rect 17334 8672 17350 8736
rect 17414 8672 17430 8736
rect 17494 8672 17502 8736
rect 17182 7648 17502 8672
rect 17182 7584 17190 7648
rect 17254 7584 17270 7648
rect 17334 7584 17350 7648
rect 17414 7584 17430 7648
rect 17494 7584 17502 7648
rect 17182 6560 17502 7584
rect 17182 6496 17190 6560
rect 17254 6496 17270 6560
rect 17334 6496 17350 6560
rect 17414 6496 17430 6560
rect 17494 6496 17502 6560
rect 17182 5472 17502 6496
rect 17182 5408 17190 5472
rect 17254 5408 17270 5472
rect 17334 5408 17350 5472
rect 17414 5408 17430 5472
rect 17494 5408 17502 5472
rect 17182 4384 17502 5408
rect 17182 4320 17190 4384
rect 17254 4320 17270 4384
rect 17334 4320 17350 4384
rect 17414 4320 17430 4384
rect 17494 4320 17502 4384
rect 17182 3296 17502 4320
rect 17182 3232 17190 3296
rect 17254 3232 17270 3296
rect 17334 3232 17350 3296
rect 17414 3232 17430 3296
rect 17494 3232 17502 3296
rect 17182 2208 17502 3232
rect 17182 2144 17190 2208
rect 17254 2144 17270 2208
rect 17334 2144 17350 2208
rect 17414 2144 17430 2208
rect 17494 2144 17502 2208
rect 17182 1120 17502 2144
rect 17182 1056 17190 1120
rect 17254 1056 17270 1120
rect 17334 1056 17350 1120
rect 17414 1056 17430 1120
rect 17494 1056 17502 1120
rect 17182 496 17502 1056
rect 20540 31040 20860 31056
rect 20540 30976 20548 31040
rect 20612 30976 20628 31040
rect 20692 30976 20708 31040
rect 20772 30976 20788 31040
rect 20852 30976 20860 31040
rect 20540 29952 20860 30976
rect 20540 29888 20548 29952
rect 20612 29888 20628 29952
rect 20692 29888 20708 29952
rect 20772 29888 20788 29952
rect 20852 29888 20860 29952
rect 20540 28864 20860 29888
rect 20540 28800 20548 28864
rect 20612 28800 20628 28864
rect 20692 28800 20708 28864
rect 20772 28800 20788 28864
rect 20852 28800 20860 28864
rect 20540 27776 20860 28800
rect 20540 27712 20548 27776
rect 20612 27712 20628 27776
rect 20692 27712 20708 27776
rect 20772 27712 20788 27776
rect 20852 27712 20860 27776
rect 20540 26688 20860 27712
rect 20540 26624 20548 26688
rect 20612 26624 20628 26688
rect 20692 26624 20708 26688
rect 20772 26624 20788 26688
rect 20852 26624 20860 26688
rect 20540 25600 20860 26624
rect 20540 25536 20548 25600
rect 20612 25536 20628 25600
rect 20692 25536 20708 25600
rect 20772 25536 20788 25600
rect 20852 25536 20860 25600
rect 20540 24512 20860 25536
rect 20540 24448 20548 24512
rect 20612 24448 20628 24512
rect 20692 24448 20708 24512
rect 20772 24448 20788 24512
rect 20852 24448 20860 24512
rect 20540 23424 20860 24448
rect 20540 23360 20548 23424
rect 20612 23360 20628 23424
rect 20692 23360 20708 23424
rect 20772 23360 20788 23424
rect 20852 23360 20860 23424
rect 20540 22336 20860 23360
rect 20540 22272 20548 22336
rect 20612 22272 20628 22336
rect 20692 22272 20708 22336
rect 20772 22272 20788 22336
rect 20852 22272 20860 22336
rect 20540 21248 20860 22272
rect 20540 21184 20548 21248
rect 20612 21184 20628 21248
rect 20692 21184 20708 21248
rect 20772 21184 20788 21248
rect 20852 21184 20860 21248
rect 20540 20160 20860 21184
rect 20540 20096 20548 20160
rect 20612 20096 20628 20160
rect 20692 20096 20708 20160
rect 20772 20096 20788 20160
rect 20852 20096 20860 20160
rect 20540 19072 20860 20096
rect 20540 19008 20548 19072
rect 20612 19008 20628 19072
rect 20692 19008 20708 19072
rect 20772 19008 20788 19072
rect 20852 19008 20860 19072
rect 20540 17984 20860 19008
rect 20540 17920 20548 17984
rect 20612 17920 20628 17984
rect 20692 17920 20708 17984
rect 20772 17920 20788 17984
rect 20852 17920 20860 17984
rect 20540 16896 20860 17920
rect 20540 16832 20548 16896
rect 20612 16832 20628 16896
rect 20692 16832 20708 16896
rect 20772 16832 20788 16896
rect 20852 16832 20860 16896
rect 20540 15808 20860 16832
rect 20540 15744 20548 15808
rect 20612 15744 20628 15808
rect 20692 15744 20708 15808
rect 20772 15744 20788 15808
rect 20852 15744 20860 15808
rect 20540 14720 20860 15744
rect 20540 14656 20548 14720
rect 20612 14656 20628 14720
rect 20692 14656 20708 14720
rect 20772 14656 20788 14720
rect 20852 14656 20860 14720
rect 20540 13632 20860 14656
rect 20540 13568 20548 13632
rect 20612 13568 20628 13632
rect 20692 13568 20708 13632
rect 20772 13568 20788 13632
rect 20852 13568 20860 13632
rect 20540 12544 20860 13568
rect 20540 12480 20548 12544
rect 20612 12480 20628 12544
rect 20692 12480 20708 12544
rect 20772 12480 20788 12544
rect 20852 12480 20860 12544
rect 20540 11456 20860 12480
rect 20540 11392 20548 11456
rect 20612 11392 20628 11456
rect 20692 11392 20708 11456
rect 20772 11392 20788 11456
rect 20852 11392 20860 11456
rect 20540 10368 20860 11392
rect 20540 10304 20548 10368
rect 20612 10304 20628 10368
rect 20692 10304 20708 10368
rect 20772 10304 20788 10368
rect 20852 10304 20860 10368
rect 20540 9280 20860 10304
rect 20540 9216 20548 9280
rect 20612 9216 20628 9280
rect 20692 9216 20708 9280
rect 20772 9216 20788 9280
rect 20852 9216 20860 9280
rect 20540 8192 20860 9216
rect 20540 8128 20548 8192
rect 20612 8128 20628 8192
rect 20692 8128 20708 8192
rect 20772 8128 20788 8192
rect 20852 8128 20860 8192
rect 20540 7104 20860 8128
rect 20540 7040 20548 7104
rect 20612 7040 20628 7104
rect 20692 7040 20708 7104
rect 20772 7040 20788 7104
rect 20852 7040 20860 7104
rect 20540 6016 20860 7040
rect 20540 5952 20548 6016
rect 20612 5952 20628 6016
rect 20692 5952 20708 6016
rect 20772 5952 20788 6016
rect 20852 5952 20860 6016
rect 20540 4928 20860 5952
rect 20540 4864 20548 4928
rect 20612 4864 20628 4928
rect 20692 4864 20708 4928
rect 20772 4864 20788 4928
rect 20852 4864 20860 4928
rect 20540 3840 20860 4864
rect 20540 3776 20548 3840
rect 20612 3776 20628 3840
rect 20692 3776 20708 3840
rect 20772 3776 20788 3840
rect 20852 3776 20860 3840
rect 20540 2752 20860 3776
rect 20540 2688 20548 2752
rect 20612 2688 20628 2752
rect 20692 2688 20708 2752
rect 20772 2688 20788 2752
rect 20852 2688 20860 2752
rect 20540 1664 20860 2688
rect 20540 1600 20548 1664
rect 20612 1600 20628 1664
rect 20692 1600 20708 1664
rect 20772 1600 20788 1664
rect 20852 1600 20860 1664
rect 20540 576 20860 1600
rect 20540 512 20548 576
rect 20612 512 20628 576
rect 20692 512 20708 576
rect 20772 512 20788 576
rect 20852 512 20860 576
rect 20540 496 20860 512
rect 23898 30496 24218 31056
rect 23898 30432 23906 30496
rect 23970 30432 23986 30496
rect 24050 30432 24066 30496
rect 24130 30432 24146 30496
rect 24210 30432 24218 30496
rect 23898 29408 24218 30432
rect 23898 29344 23906 29408
rect 23970 29344 23986 29408
rect 24050 29344 24066 29408
rect 24130 29344 24146 29408
rect 24210 29344 24218 29408
rect 23898 28320 24218 29344
rect 23898 28256 23906 28320
rect 23970 28256 23986 28320
rect 24050 28256 24066 28320
rect 24130 28256 24146 28320
rect 24210 28256 24218 28320
rect 23898 27232 24218 28256
rect 27256 31040 27576 31056
rect 27256 30976 27264 31040
rect 27328 30976 27344 31040
rect 27408 30976 27424 31040
rect 27488 30976 27504 31040
rect 27568 30976 27576 31040
rect 27256 29952 27576 30976
rect 27256 29888 27264 29952
rect 27328 29888 27344 29952
rect 27408 29888 27424 29952
rect 27488 29888 27504 29952
rect 27568 29888 27576 29952
rect 27256 28864 27576 29888
rect 27256 28800 27264 28864
rect 27328 28800 27344 28864
rect 27408 28800 27424 28864
rect 27488 28800 27504 28864
rect 27568 28800 27576 28864
rect 27256 27776 27576 28800
rect 27256 27712 27264 27776
rect 27328 27712 27344 27776
rect 27408 27712 27424 27776
rect 27488 27712 27504 27776
rect 27568 27712 27576 27776
rect 24899 27708 24965 27709
rect 24899 27644 24900 27708
rect 24964 27644 24965 27708
rect 24899 27643 24965 27644
rect 23898 27168 23906 27232
rect 23970 27168 23986 27232
rect 24050 27168 24066 27232
rect 24130 27168 24146 27232
rect 24210 27168 24218 27232
rect 23898 26144 24218 27168
rect 23898 26080 23906 26144
rect 23970 26080 23986 26144
rect 24050 26080 24066 26144
rect 24130 26080 24146 26144
rect 24210 26080 24218 26144
rect 23898 25056 24218 26080
rect 23898 24992 23906 25056
rect 23970 24992 23986 25056
rect 24050 24992 24066 25056
rect 24130 24992 24146 25056
rect 24210 24992 24218 25056
rect 23898 23968 24218 24992
rect 23898 23904 23906 23968
rect 23970 23904 23986 23968
rect 24050 23904 24066 23968
rect 24130 23904 24146 23968
rect 24210 23904 24218 23968
rect 23898 22880 24218 23904
rect 23898 22816 23906 22880
rect 23970 22816 23986 22880
rect 24050 22816 24066 22880
rect 24130 22816 24146 22880
rect 24210 22816 24218 22880
rect 23898 21792 24218 22816
rect 23898 21728 23906 21792
rect 23970 21728 23986 21792
rect 24050 21728 24066 21792
rect 24130 21728 24146 21792
rect 24210 21728 24218 21792
rect 23898 20704 24218 21728
rect 23898 20640 23906 20704
rect 23970 20640 23986 20704
rect 24050 20640 24066 20704
rect 24130 20640 24146 20704
rect 24210 20640 24218 20704
rect 23898 19616 24218 20640
rect 23898 19552 23906 19616
rect 23970 19552 23986 19616
rect 24050 19552 24066 19616
rect 24130 19552 24146 19616
rect 24210 19552 24218 19616
rect 23898 18528 24218 19552
rect 23898 18464 23906 18528
rect 23970 18464 23986 18528
rect 24050 18464 24066 18528
rect 24130 18464 24146 18528
rect 24210 18464 24218 18528
rect 23898 17440 24218 18464
rect 23898 17376 23906 17440
rect 23970 17376 23986 17440
rect 24050 17376 24066 17440
rect 24130 17376 24146 17440
rect 24210 17376 24218 17440
rect 23898 16352 24218 17376
rect 24902 17101 24962 27643
rect 27256 26688 27576 27712
rect 27256 26624 27264 26688
rect 27328 26624 27344 26688
rect 27408 26624 27424 26688
rect 27488 26624 27504 26688
rect 27568 26624 27576 26688
rect 27256 25600 27576 26624
rect 27256 25536 27264 25600
rect 27328 25536 27344 25600
rect 27408 25536 27424 25600
rect 27488 25536 27504 25600
rect 27568 25536 27576 25600
rect 27256 24512 27576 25536
rect 27256 24448 27264 24512
rect 27328 24448 27344 24512
rect 27408 24448 27424 24512
rect 27488 24448 27504 24512
rect 27568 24448 27576 24512
rect 27256 23424 27576 24448
rect 27256 23360 27264 23424
rect 27328 23360 27344 23424
rect 27408 23360 27424 23424
rect 27488 23360 27504 23424
rect 27568 23360 27576 23424
rect 27256 22336 27576 23360
rect 27256 22272 27264 22336
rect 27328 22272 27344 22336
rect 27408 22272 27424 22336
rect 27488 22272 27504 22336
rect 27568 22272 27576 22336
rect 27256 21248 27576 22272
rect 27256 21184 27264 21248
rect 27328 21184 27344 21248
rect 27408 21184 27424 21248
rect 27488 21184 27504 21248
rect 27568 21184 27576 21248
rect 27256 20160 27576 21184
rect 27256 20096 27264 20160
rect 27328 20096 27344 20160
rect 27408 20096 27424 20160
rect 27488 20096 27504 20160
rect 27568 20096 27576 20160
rect 27256 19072 27576 20096
rect 27256 19008 27264 19072
rect 27328 19008 27344 19072
rect 27408 19008 27424 19072
rect 27488 19008 27504 19072
rect 27568 19008 27576 19072
rect 27256 17984 27576 19008
rect 27256 17920 27264 17984
rect 27328 17920 27344 17984
rect 27408 17920 27424 17984
rect 27488 17920 27504 17984
rect 27568 17920 27576 17984
rect 24899 17100 24965 17101
rect 24899 17036 24900 17100
rect 24964 17036 24965 17100
rect 24899 17035 24965 17036
rect 23898 16288 23906 16352
rect 23970 16288 23986 16352
rect 24050 16288 24066 16352
rect 24130 16288 24146 16352
rect 24210 16288 24218 16352
rect 23898 15264 24218 16288
rect 23898 15200 23906 15264
rect 23970 15200 23986 15264
rect 24050 15200 24066 15264
rect 24130 15200 24146 15264
rect 24210 15200 24218 15264
rect 23898 14176 24218 15200
rect 23898 14112 23906 14176
rect 23970 14112 23986 14176
rect 24050 14112 24066 14176
rect 24130 14112 24146 14176
rect 24210 14112 24218 14176
rect 23898 13088 24218 14112
rect 23898 13024 23906 13088
rect 23970 13024 23986 13088
rect 24050 13024 24066 13088
rect 24130 13024 24146 13088
rect 24210 13024 24218 13088
rect 23898 12000 24218 13024
rect 23898 11936 23906 12000
rect 23970 11936 23986 12000
rect 24050 11936 24066 12000
rect 24130 11936 24146 12000
rect 24210 11936 24218 12000
rect 23898 10912 24218 11936
rect 23898 10848 23906 10912
rect 23970 10848 23986 10912
rect 24050 10848 24066 10912
rect 24130 10848 24146 10912
rect 24210 10848 24218 10912
rect 23898 9824 24218 10848
rect 23898 9760 23906 9824
rect 23970 9760 23986 9824
rect 24050 9760 24066 9824
rect 24130 9760 24146 9824
rect 24210 9760 24218 9824
rect 23898 8736 24218 9760
rect 23898 8672 23906 8736
rect 23970 8672 23986 8736
rect 24050 8672 24066 8736
rect 24130 8672 24146 8736
rect 24210 8672 24218 8736
rect 23898 7648 24218 8672
rect 23898 7584 23906 7648
rect 23970 7584 23986 7648
rect 24050 7584 24066 7648
rect 24130 7584 24146 7648
rect 24210 7584 24218 7648
rect 23898 6560 24218 7584
rect 23898 6496 23906 6560
rect 23970 6496 23986 6560
rect 24050 6496 24066 6560
rect 24130 6496 24146 6560
rect 24210 6496 24218 6560
rect 23898 5472 24218 6496
rect 23898 5408 23906 5472
rect 23970 5408 23986 5472
rect 24050 5408 24066 5472
rect 24130 5408 24146 5472
rect 24210 5408 24218 5472
rect 23898 4384 24218 5408
rect 23898 4320 23906 4384
rect 23970 4320 23986 4384
rect 24050 4320 24066 4384
rect 24130 4320 24146 4384
rect 24210 4320 24218 4384
rect 23898 3296 24218 4320
rect 23898 3232 23906 3296
rect 23970 3232 23986 3296
rect 24050 3232 24066 3296
rect 24130 3232 24146 3296
rect 24210 3232 24218 3296
rect 23898 2208 24218 3232
rect 23898 2144 23906 2208
rect 23970 2144 23986 2208
rect 24050 2144 24066 2208
rect 24130 2144 24146 2208
rect 24210 2144 24218 2208
rect 23898 1120 24218 2144
rect 23898 1056 23906 1120
rect 23970 1056 23986 1120
rect 24050 1056 24066 1120
rect 24130 1056 24146 1120
rect 24210 1056 24218 1120
rect 23898 496 24218 1056
rect 27256 16896 27576 17920
rect 27256 16832 27264 16896
rect 27328 16832 27344 16896
rect 27408 16832 27424 16896
rect 27488 16832 27504 16896
rect 27568 16832 27576 16896
rect 27256 15808 27576 16832
rect 27256 15744 27264 15808
rect 27328 15744 27344 15808
rect 27408 15744 27424 15808
rect 27488 15744 27504 15808
rect 27568 15744 27576 15808
rect 27256 14720 27576 15744
rect 27256 14656 27264 14720
rect 27328 14656 27344 14720
rect 27408 14656 27424 14720
rect 27488 14656 27504 14720
rect 27568 14656 27576 14720
rect 27256 13632 27576 14656
rect 27256 13568 27264 13632
rect 27328 13568 27344 13632
rect 27408 13568 27424 13632
rect 27488 13568 27504 13632
rect 27568 13568 27576 13632
rect 27256 12544 27576 13568
rect 27256 12480 27264 12544
rect 27328 12480 27344 12544
rect 27408 12480 27424 12544
rect 27488 12480 27504 12544
rect 27568 12480 27576 12544
rect 27256 11456 27576 12480
rect 27256 11392 27264 11456
rect 27328 11392 27344 11456
rect 27408 11392 27424 11456
rect 27488 11392 27504 11456
rect 27568 11392 27576 11456
rect 27256 10368 27576 11392
rect 27256 10304 27264 10368
rect 27328 10304 27344 10368
rect 27408 10304 27424 10368
rect 27488 10304 27504 10368
rect 27568 10304 27576 10368
rect 27256 9280 27576 10304
rect 27256 9216 27264 9280
rect 27328 9216 27344 9280
rect 27408 9216 27424 9280
rect 27488 9216 27504 9280
rect 27568 9216 27576 9280
rect 27256 8192 27576 9216
rect 27256 8128 27264 8192
rect 27328 8128 27344 8192
rect 27408 8128 27424 8192
rect 27488 8128 27504 8192
rect 27568 8128 27576 8192
rect 27256 7104 27576 8128
rect 27256 7040 27264 7104
rect 27328 7040 27344 7104
rect 27408 7040 27424 7104
rect 27488 7040 27504 7104
rect 27568 7040 27576 7104
rect 27256 6016 27576 7040
rect 27256 5952 27264 6016
rect 27328 5952 27344 6016
rect 27408 5952 27424 6016
rect 27488 5952 27504 6016
rect 27568 5952 27576 6016
rect 27256 4928 27576 5952
rect 27256 4864 27264 4928
rect 27328 4864 27344 4928
rect 27408 4864 27424 4928
rect 27488 4864 27504 4928
rect 27568 4864 27576 4928
rect 27256 3840 27576 4864
rect 27256 3776 27264 3840
rect 27328 3776 27344 3840
rect 27408 3776 27424 3840
rect 27488 3776 27504 3840
rect 27568 3776 27576 3840
rect 27256 2752 27576 3776
rect 27256 2688 27264 2752
rect 27328 2688 27344 2752
rect 27408 2688 27424 2752
rect 27488 2688 27504 2752
rect 27568 2688 27576 2752
rect 27256 1664 27576 2688
rect 27256 1600 27264 1664
rect 27328 1600 27344 1664
rect 27408 1600 27424 1664
rect 27488 1600 27504 1664
rect 27568 1600 27576 1664
rect 27256 576 27576 1600
rect 27256 512 27264 576
rect 27328 512 27344 576
rect 27408 512 27424 576
rect 27488 512 27504 576
rect 27568 512 27576 576
rect 27256 496 27576 512
use sky130_fd_sc_hd__and4b_1  _1068_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7176 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__nand4b_1  _1069_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7728 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _1070_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6900 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_4  _1071_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4876 0 1 17952
box -38 -48 1418 592
use sky130_fd_sc_hd__buf_2  _1072_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3496 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1073_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4784 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1074_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5244 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1075_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5244 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1076_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5060 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1077_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4600 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1078_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3864 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1079_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5152 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1080_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4876 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1081_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3496 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1082_
timestamp 1704896540
transform 1 0 3772 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1083_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2208 0 -1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1084_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2852 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1085_
timestamp 1704896540
transform -1 0 2944 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1086_
timestamp 1704896540
transform 1 0 1196 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1087_
timestamp 1704896540
transform -1 0 3772 0 -1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1088_
timestamp 1704896540
transform 1 0 2668 0 1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1089_
timestamp 1704896540
transform 1 0 2668 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1090_
timestamp 1704896540
transform -1 0 3588 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1091_
timestamp 1704896540
transform 1 0 1656 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1092_
timestamp 1704896540
transform -1 0 3220 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1093_
timestamp 1704896540
transform 1 0 2116 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1094_
timestamp 1704896540
transform 1 0 1012 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1095_
timestamp 1704896540
transform -1 0 3680 0 1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1096_
timestamp 1704896540
transform 1 0 2208 0 -1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1097_
timestamp 1704896540
transform -1 0 2944 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1098_
timestamp 1704896540
transform 1 0 1012 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1099_
timestamp 1704896540
transform 1 0 2208 0 1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1100_
timestamp 1704896540
transform 1 0 2208 0 1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1101_
timestamp 1704896540
transform -1 0 3036 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1102_
timestamp 1704896540
transform 1 0 1380 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1103_
timestamp 1704896540
transform 1 0 2668 0 1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1104_
timestamp 1704896540
transform 1 0 3036 0 -1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1105_
timestamp 1704896540
transform 1 0 3220 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1106_
timestamp 1704896540
transform 1 0 3588 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1107_
timestamp 1704896540
transform 1 0 4508 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1108_
timestamp 1704896540
transform 1 0 4508 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1109_
timestamp 1704896540
transform -1 0 5796 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1110_
timestamp 1704896540
transform 1 0 4876 0 -1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1111_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5612 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1112_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5244 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1113_
timestamp 1704896540
transform -1 0 5796 0 1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1114_
timestamp 1704896540
transform 1 0 5796 0 1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1115_
timestamp 1704896540
transform 1 0 4692 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1116_
timestamp 1704896540
transform -1 0 5520 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1117_
timestamp 1704896540
transform -1 0 4600 0 -1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1118_
timestamp 1704896540
transform -1 0 4876 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1119_
timestamp 1704896540
transform -1 0 4140 0 -1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1120_
timestamp 1704896540
transform 1 0 2484 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1121_
timestamp 1704896540
transform -1 0 4048 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1122_
timestamp 1704896540
transform 1 0 2760 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1123_
timestamp 1704896540
transform -1 0 4508 0 -1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1124_
timestamp 1704896540
transform 1 0 2208 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1125_
timestamp 1704896540
transform -1 0 4416 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1126_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3680 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1127_
timestamp 1704896540
transform -1 0 4692 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1128_
timestamp 1704896540
transform 1 0 3496 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1129_
timestamp 1704896540
transform 1 0 3680 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1130_
timestamp 1704896540
transform 1 0 4508 0 -1 29920
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1131_
timestamp 1704896540
transform 1 0 4232 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1132_
timestamp 1704896540
transform 1 0 4784 0 1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1133_
timestamp 1704896540
transform -1 0 5520 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1134_
timestamp 1704896540
transform 1 0 4968 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1135_
timestamp 1704896540
transform 1 0 5796 0 -1 29920
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1136_
timestamp 1704896540
transform -1 0 6164 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1137_
timestamp 1704896540
transform -1 0 5704 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1138_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4416 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _1139_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8096 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _1140_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8280 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1141_
timestamp 1704896540
transform 1 0 9016 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1142_
timestamp 1704896540
transform 1 0 8464 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1143_
timestamp 1704896540
transform 1 0 8372 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1144_
timestamp 1704896540
transform -1 0 9016 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1145_
timestamp 1704896540
transform -1 0 9200 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1146_
timestamp 1704896540
transform 1 0 7636 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1147_
timestamp 1704896540
transform 1 0 8004 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1148_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7452 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1149_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8004 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1150_
timestamp 1704896540
transform -1 0 10396 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1151_
timestamp 1704896540
transform -1 0 9292 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1152_
timestamp 1704896540
transform 1 0 9016 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1153_
timestamp 1704896540
transform 1 0 9476 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1154_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9568 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1155_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10304 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nor2b_2  _1156_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 17020 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__nor2b_1  _1157_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 20424 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1158_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 21896 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1159_
timestamp 1704896540
transform -1 0 21068 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1160_
timestamp 1704896540
transform -1 0 23184 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1161_
timestamp 1704896540
transform 1 0 20884 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1162_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 13064 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_2  _1163_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11960 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1164_
timestamp 1704896540
transform -1 0 12512 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1165_
timestamp 1704896540
transform -1 0 11868 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1166_
timestamp 1704896540
transform -1 0 11868 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1167_
timestamp 1704896540
transform -1 0 12420 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1168_
timestamp 1704896540
transform -1 0 12328 0 1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1169_
timestamp 1704896540
transform -1 0 11592 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1170_
timestamp 1704896540
transform -1 0 13248 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1171_
timestamp 1704896540
transform -1 0 13340 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1172_
timestamp 1704896540
transform -1 0 9384 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1173_
timestamp 1704896540
transform 1 0 8648 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1174_
timestamp 1704896540
transform 1 0 8648 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1175_
timestamp 1704896540
transform -1 0 9384 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1176_
timestamp 1704896540
transform -1 0 7728 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1177_
timestamp 1704896540
transform 1 0 7728 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1178_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8556 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1179_
timestamp 1704896540
transform 1 0 8464 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1180_
timestamp 1704896540
transform 1 0 8924 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1181_
timestamp 1704896540
transform -1 0 9660 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1182_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8188 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1183_
timestamp 1704896540
transform -1 0 8004 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1184_
timestamp 1704896540
transform -1 0 8280 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1185_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7728 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1186_
timestamp 1704896540
transform 1 0 8372 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1187_
timestamp 1704896540
transform -1 0 8924 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1188_
timestamp 1704896540
transform -1 0 7912 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1189_
timestamp 1704896540
transform 1 0 7176 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1190_
timestamp 1704896540
transform -1 0 6440 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1191_
timestamp 1704896540
transform 1 0 6532 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1192_
timestamp 1704896540
transform 1 0 6440 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1193_
timestamp 1704896540
transform -1 0 7176 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1194_
timestamp 1704896540
transform -1 0 7084 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1195_
timestamp 1704896540
transform 1 0 6348 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1196_
timestamp 1704896540
transform -1 0 7544 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1197_
timestamp 1704896540
transform -1 0 4232 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1198_
timestamp 1704896540
transform -1 0 4692 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1199_
timestamp 1704896540
transform -1 0 5152 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1200_
timestamp 1704896540
transform -1 0 2852 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1201_
timestamp 1704896540
transform 1 0 2852 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1202_
timestamp 1704896540
transform 1 0 3404 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1203_
timestamp 1704896540
transform 1 0 4048 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1204_
timestamp 1704896540
transform 1 0 4232 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1205_
timestamp 1704896540
transform -1 0 5612 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1206_
timestamp 1704896540
transform -1 0 5520 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1207_
timestamp 1704896540
transform 1 0 3496 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1208_
timestamp 1704896540
transform -1 0 3496 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1209_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3220 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1210_
timestamp 1704896540
transform -1 0 2208 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1211_
timestamp 1704896540
transform 1 0 2208 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1212_
timestamp 1704896540
transform -1 0 2852 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _1213_
timestamp 1704896540
transform 1 0 1380 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1214_
timestamp 1704896540
transform 1 0 1380 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1215_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2024 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _1216_
timestamp 1704896540
transform 1 0 1932 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _1217_
timestamp 1704896540
transform 1 0 828 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1218_
timestamp 1704896540
transform 1 0 2024 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1219_
timestamp 1704896540
transform -1 0 3220 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1220_
timestamp 1704896540
transform -1 0 1932 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1221_
timestamp 1704896540
transform -1 0 18400 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1222_
timestamp 1704896540
transform 1 0 18308 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1223_
timestamp 1704896540
transform -1 0 18124 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1224_
timestamp 1704896540
transform 1 0 17480 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1225_
timestamp 1704896540
transform -1 0 17572 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1226_
timestamp 1704896540
transform 1 0 17572 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1227_
timestamp 1704896540
transform 1 0 18032 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1228_
timestamp 1704896540
transform 1 0 17756 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1229_
timestamp 1704896540
transform 1 0 18676 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1230_
timestamp 1704896540
transform -1 0 19412 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1231_
timestamp 1704896540
transform -1 0 18216 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1232_
timestamp 1704896540
transform -1 0 18400 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1233_
timestamp 1704896540
transform -1 0 18676 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1234_
timestamp 1704896540
transform 1 0 17940 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1235_
timestamp 1704896540
transform 1 0 17940 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1236_
timestamp 1704896540
transform 1 0 18860 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1237_
timestamp 1704896540
transform -1 0 19596 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1238_
timestamp 1704896540
transform 1 0 17572 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1239_
timestamp 1704896540
transform -1 0 16836 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1240_
timestamp 1704896540
transform -1 0 16836 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1241_
timestamp 1704896540
transform -1 0 17756 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1242_
timestamp 1704896540
transform 1 0 16560 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1243_
timestamp 1704896540
transform 1 0 17204 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1244_
timestamp 1704896540
transform -1 0 17664 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1245_
timestamp 1704896540
transform 1 0 16008 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1246_
timestamp 1704896540
transform 1 0 15456 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1247_
timestamp 1704896540
transform 1 0 14076 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1248_
timestamp 1704896540
transform 1 0 14904 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1249_
timestamp 1704896540
transform -1 0 13892 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1250_
timestamp 1704896540
transform -1 0 12972 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1251_
timestamp 1704896540
transform 1 0 14628 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1252_
timestamp 1704896540
transform -1 0 15456 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1253_
timestamp 1704896540
transform 1 0 15272 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1254_
timestamp 1704896540
transform 1 0 15916 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1255_
timestamp 1704896540
transform -1 0 16468 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1256_
timestamp 1704896540
transform 1 0 14720 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1257_
timestamp 1704896540
transform -1 0 14720 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1258_
timestamp 1704896540
transform 1 0 14444 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1259_
timestamp 1704896540
transform -1 0 12420 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1260_
timestamp 1704896540
transform -1 0 11592 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1261_
timestamp 1704896540
transform 1 0 11960 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _1262_
timestamp 1704896540
transform 1 0 11500 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1263_
timestamp 1704896540
transform 1 0 12512 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1264_
timestamp 1704896540
transform 1 0 10948 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1265_
timestamp 1704896540
transform -1 0 11960 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__a21boi_1  _1266_
timestamp 1704896540
transform 1 0 10028 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1267_
timestamp 1704896540
transform -1 0 12144 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1268_
timestamp 1704896540
transform -1 0 10488 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1269_
timestamp 1704896540
transform 1 0 9844 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _1270_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11132 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _1271_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10764 0 1 9248
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _1272_
timestamp 1704896540
transform 1 0 14536 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1273_
timestamp 1704896540
transform 1 0 7636 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_4  _1274_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 16192 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__a211o_2  _1275_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 13800 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _1276_
timestamp 1704896540
transform 1 0 10948 0 -1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _1277_
timestamp 1704896540
transform -1 0 14628 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_2  _1278_
timestamp 1704896540
transform 1 0 13708 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1279_
timestamp 1704896540
transform -1 0 3220 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _1280_
timestamp 1704896540
transform 1 0 10672 0 1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _1281_
timestamp 1704896540
transform -1 0 15180 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_2  _1282_
timestamp 1704896540
transform 1 0 13892 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1283_
timestamp 1704896540
transform -1 0 2852 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _1284_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10948 0 -1 9248
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _1285_
timestamp 1704896540
transform -1 0 14904 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_2  _1286_
timestamp 1704896540
transform 1 0 13708 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1287_
timestamp 1704896540
transform -1 0 2484 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_4  _1288_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 15548 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_1  _1289_
timestamp 1704896540
transform 1 0 3496 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1290_
timestamp 1704896540
transform 1 0 4232 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1291_
timestamp 1704896540
transform -1 0 5336 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1292_
timestamp 1704896540
transform 1 0 5612 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1293_
timestamp 1704896540
transform 1 0 4140 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1294_
timestamp 1704896540
transform 1 0 4784 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1295_
timestamp 1704896540
transform 1 0 4048 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1296_
timestamp 1704896540
transform -1 0 6532 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1297_
timestamp 1704896540
transform 1 0 2944 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1298_
timestamp 1704896540
transform 1 0 2668 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1299_
timestamp 1704896540
transform -1 0 2760 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1300_
timestamp 1704896540
transform 1 0 5796 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1301_
timestamp 1704896540
transform 1 0 3220 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1302_
timestamp 1704896540
transform 1 0 4692 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1303_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5152 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1304_
timestamp 1704896540
transform -1 0 5888 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1305_
timestamp 1704896540
transform 1 0 6624 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1306_
timestamp 1704896540
transform -1 0 7360 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1307_
timestamp 1704896540
transform -1 0 6992 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1308_
timestamp 1704896540
transform -1 0 6992 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1309_
timestamp 1704896540
transform -1 0 6716 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _1310_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3312 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1311_
timestamp 1704896540
transform -1 0 4600 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1312_
timestamp 1704896540
transform -1 0 5704 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1313_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6072 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1314_
timestamp 1704896540
transform -1 0 6992 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1315_
timestamp 1704896540
transform 1 0 2024 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1316_
timestamp 1704896540
transform 1 0 3404 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1317_
timestamp 1704896540
transform 1 0 6164 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1318_
timestamp 1704896540
transform 1 0 6072 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1319_
timestamp 1704896540
transform -1 0 6624 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1320_
timestamp 1704896540
transform -1 0 3496 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1321_
timestamp 1704896540
transform -1 0 5612 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1322_
timestamp 1704896540
transform -1 0 6256 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1323_
timestamp 1704896540
transform -1 0 5980 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1324_
timestamp 1704896540
transform 1 0 4968 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1325_
timestamp 1704896540
transform 1 0 4692 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1326_
timestamp 1704896540
transform -1 0 5152 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1327_
timestamp 1704896540
transform 1 0 2116 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1328_
timestamp 1704896540
transform 1 0 2668 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1329_
timestamp 1704896540
transform -1 0 4600 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1330_
timestamp 1704896540
transform -1 0 4876 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1331_
timestamp 1704896540
transform -1 0 4232 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1332_
timestamp 1704896540
transform 1 0 3496 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1333_
timestamp 1704896540
transform -1 0 3680 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1334_
timestamp 1704896540
transform -1 0 2208 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1335_
timestamp 1704896540
transform 1 0 1656 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_4  _1336_
timestamp 1704896540
transform -1 0 18952 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_1  _1337_
timestamp 1704896540
transform -1 0 13616 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_2  _1338_
timestamp 1704896540
transform 1 0 11868 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1339_
timestamp 1704896540
transform -1 0 13432 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_2  _1340_
timestamp 1704896540
transform 1 0 12604 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1341_
timestamp 1704896540
transform -1 0 11960 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1342_
timestamp 1704896540
transform 1 0 13156 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_2  _1343_
timestamp 1704896540
transform -1 0 13708 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1344_
timestamp 1704896540
transform -1 0 11408 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1345_
timestamp 1704896540
transform -1 0 12696 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1346_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12052 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1347_
timestamp 1704896540
transform -1 0 10856 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_2  _1348_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12420 0 1 8160
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1349_
timestamp 1704896540
transform 1 0 12236 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1350_
timestamp 1704896540
transform 1 0 12880 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1351_
timestamp 1704896540
transform -1 0 14168 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1352_
timestamp 1704896540
transform 1 0 15548 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1353_
timestamp 1704896540
transform 1 0 12696 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1354_
timestamp 1704896540
transform 1 0 13524 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1355_
timestamp 1704896540
transform 1 0 12512 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1356_
timestamp 1704896540
transform -1 0 14812 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1357_
timestamp 1704896540
transform -1 0 11960 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1358_
timestamp 1704896540
transform -1 0 11316 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1359_
timestamp 1704896540
transform -1 0 11040 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1360_
timestamp 1704896540
transform 1 0 14904 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1361_
timestamp 1704896540
transform 1 0 11684 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1362_
timestamp 1704896540
transform 1 0 13248 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1363_
timestamp 1704896540
transform 1 0 13708 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1364_
timestamp 1704896540
transform -1 0 14996 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1365_
timestamp 1704896540
transform 1 0 16100 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1366_
timestamp 1704896540
transform -1 0 16192 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1367_
timestamp 1704896540
transform 1 0 13156 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1368_
timestamp 1704896540
transform 1 0 12788 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1369_
timestamp 1704896540
transform 1 0 14260 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _1370_
timestamp 1704896540
transform -1 0 11684 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1371_
timestamp 1704896540
transform 1 0 12880 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1372_
timestamp 1704896540
transform -1 0 14076 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1373_
timestamp 1704896540
transform 1 0 14996 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1374_
timestamp 1704896540
transform -1 0 15548 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1375_
timestamp 1704896540
transform 1 0 10580 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1376_
timestamp 1704896540
transform 1 0 11500 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1377_
timestamp 1704896540
transform -1 0 14812 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1378_
timestamp 1704896540
transform 1 0 15180 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1379_
timestamp 1704896540
transform -1 0 15824 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1380_
timestamp 1704896540
transform -1 0 12236 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1381_
timestamp 1704896540
transform 1 0 14260 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1382_
timestamp 1704896540
transform 1 0 14720 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1383_
timestamp 1704896540
transform -1 0 15548 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1384_
timestamp 1704896540
transform -1 0 13892 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1385_
timestamp 1704896540
transform 1 0 13800 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1386_
timestamp 1704896540
transform -1 0 14444 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1387_
timestamp 1704896540
transform -1 0 12788 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1388_
timestamp 1704896540
transform -1 0 12788 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1389_
timestamp 1704896540
transform 1 0 12788 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1390_
timestamp 1704896540
transform -1 0 12788 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1391_
timestamp 1704896540
transform -1 0 12696 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1392_
timestamp 1704896540
transform 1 0 11960 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1393_
timestamp 1704896540
transform -1 0 11960 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1394_
timestamp 1704896540
transform -1 0 10764 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1395_
timestamp 1704896540
transform 1 0 10212 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_4  _1396_
timestamp 1704896540
transform -1 0 20516 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_1  _1397_
timestamp 1704896540
transform -1 0 19228 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_2  _1398_
timestamp 1704896540
transform -1 0 19320 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1399_
timestamp 1704896540
transform 1 0 18676 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_2  _1400_
timestamp 1704896540
transform 1 0 18216 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1401_
timestamp 1704896540
transform 1 0 19596 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1402_
timestamp 1704896540
transform -1 0 20332 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_2  _1403_
timestamp 1704896540
transform 1 0 19320 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1404_
timestamp 1704896540
transform -1 0 20516 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1405_
timestamp 1704896540
transform 1 0 18308 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1406_
timestamp 1704896540
transform -1 0 19688 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1407_
timestamp 1704896540
transform -1 0 19596 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_2  _1408_
timestamp 1704896540
transform -1 0 19872 0 1 7072
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1409_
timestamp 1704896540
transform 1 0 20516 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1410_
timestamp 1704896540
transform 1 0 21252 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1411_
timestamp 1704896540
transform -1 0 22540 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1412_
timestamp 1704896540
transform 1 0 22632 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1413_
timestamp 1704896540
transform 1 0 21160 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1414_
timestamp 1704896540
transform 1 0 22172 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1415_
timestamp 1704896540
transform 1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1416_
timestamp 1704896540
transform 1 0 22080 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1417_
timestamp 1704896540
transform -1 0 19964 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1418_
timestamp 1704896540
transform 1 0 19504 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1419_
timestamp 1704896540
transform -1 0 19872 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1420_
timestamp 1704896540
transform 1 0 22816 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1421_
timestamp 1704896540
transform 1 0 20056 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1422_
timestamp 1704896540
transform 1 0 21712 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1423_
timestamp 1704896540
transform 1 0 21988 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1424_
timestamp 1704896540
transform -1 0 23000 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1425_
timestamp 1704896540
transform 1 0 23092 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1426_
timestamp 1704896540
transform -1 0 24196 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1427_
timestamp 1704896540
transform -1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1428_
timestamp 1704896540
transform 1 0 20332 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1429_
timestamp 1704896540
transform -1 0 22816 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _1430_
timestamp 1704896540
transform -1 0 21528 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1431_
timestamp 1704896540
transform 1 0 21528 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1432_
timestamp 1704896540
transform -1 0 22356 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1433_
timestamp 1704896540
transform 1 0 23000 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1434_
timestamp 1704896540
transform -1 0 23920 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1435_
timestamp 1704896540
transform 1 0 19872 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1436_
timestamp 1704896540
transform -1 0 21160 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1437_
timestamp 1704896540
transform 1 0 22264 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1438_
timestamp 1704896540
transform 1 0 23000 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1439_
timestamp 1704896540
transform -1 0 24012 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1440_
timestamp 1704896540
transform -1 0 21068 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1441_
timestamp 1704896540
transform -1 0 22632 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1442_
timestamp 1704896540
transform 1 0 22724 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1443_
timestamp 1704896540
transform -1 0 23460 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1444_
timestamp 1704896540
transform 1 0 21988 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1445_
timestamp 1704896540
transform 1 0 22080 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1446_
timestamp 1704896540
transform 1 0 22816 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1447_
timestamp 1704896540
transform -1 0 21160 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1448_
timestamp 1704896540
transform 1 0 21252 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1449_
timestamp 1704896540
transform 1 0 21252 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1450_
timestamp 1704896540
transform -1 0 21068 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1451_
timestamp 1704896540
transform -1 0 21068 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1452_
timestamp 1704896540
transform -1 0 20516 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1453_
timestamp 1704896540
transform 1 0 20516 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1454_
timestamp 1704896540
transform 1 0 19872 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1455_
timestamp 1704896540
transform 1 0 19044 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_2  _1456_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12420 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__nand3b_2  _1457_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 13524 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1458_
timestamp 1704896540
transform -1 0 14720 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1459_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 14444 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1460_
timestamp 1704896540
transform 1 0 10396 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1461_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 20608 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1462_
timestamp 1704896540
transform 1 0 15180 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1463_
timestamp 1704896540
transform 1 0 15640 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1464_
timestamp 1704896540
transform 1 0 16928 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1465_
timestamp 1704896540
transform 1 0 17112 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1466_
timestamp 1704896540
transform 1 0 20516 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1467_
timestamp 1704896540
transform -1 0 19596 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1468_
timestamp 1704896540
transform -1 0 16652 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1469_
timestamp 1704896540
transform -1 0 17848 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1470_
timestamp 1704896540
transform 1 0 19872 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1471_
timestamp 1704896540
transform 1 0 17572 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  _1472_
timestamp 1704896540
transform 1 0 18676 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1473_
timestamp 1704896540
transform -1 0 18308 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1474_
timestamp 1704896540
transform 1 0 17020 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1475_
timestamp 1704896540
transform -1 0 18492 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1476_
timestamp 1704896540
transform 1 0 13064 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1477_
timestamp 1704896540
transform -1 0 20332 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__nand3b_4  _1478_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 14996 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_4  _1479_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 16744 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1480_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 19872 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1481_
timestamp 1704896540
transform 1 0 20332 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1482_
timestamp 1704896540
transform -1 0 18768 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1483_
timestamp 1704896540
transform 1 0 17756 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1484_
timestamp 1704896540
transform -1 0 17296 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1485_
timestamp 1704896540
transform -1 0 21160 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1486_
timestamp 1704896540
transform 1 0 20608 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1487_
timestamp 1704896540
transform 1 0 20424 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1488_
timestamp 1704896540
transform -1 0 18584 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1489_
timestamp 1704896540
transform 1 0 17296 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1490_
timestamp 1704896540
transform -1 0 17204 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1491_
timestamp 1704896540
transform 1 0 21252 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _1492_
timestamp 1704896540
transform 1 0 16376 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1493_
timestamp 1704896540
transform 1 0 21252 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1494_
timestamp 1704896540
transform 1 0 20516 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1495_
timestamp 1704896540
transform -1 0 20056 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1496_
timestamp 1704896540
transform 1 0 19044 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1497_
timestamp 1704896540
transform -1 0 19320 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1498_
timestamp 1704896540
transform -1 0 20792 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1499_
timestamp 1704896540
transform -1 0 19872 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1500_
timestamp 1704896540
transform 1 0 19412 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1501_
timestamp 1704896540
transform 1 0 20700 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1502_
timestamp 1704896540
transform 1 0 21252 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1503_
timestamp 1704896540
transform -1 0 20976 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1504_
timestamp 1704896540
transform 1 0 14260 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1505_
timestamp 1704896540
transform 1 0 14352 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1506_
timestamp 1704896540
transform 1 0 15364 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1507_
timestamp 1704896540
transform 1 0 16100 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1508_
timestamp 1704896540
transform 1 0 14812 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1509_
timestamp 1704896540
transform -1 0 13892 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1510_
timestamp 1704896540
transform -1 0 18584 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1511_
timestamp 1704896540
transform 1 0 17480 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1512_
timestamp 1704896540
transform 1 0 17204 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1513_
timestamp 1704896540
transform -1 0 18584 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1514_
timestamp 1704896540
transform 1 0 17572 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1515_
timestamp 1704896540
transform -1 0 17756 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1516_
timestamp 1704896540
transform -1 0 16836 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1517_
timestamp 1704896540
transform -1 0 15732 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1518_
timestamp 1704896540
transform 1 0 14628 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1519_
timestamp 1704896540
transform 1 0 14260 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1520_
timestamp 1704896540
transform -1 0 16928 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1521_
timestamp 1704896540
transform 1 0 16100 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1522_
timestamp 1704896540
transform -1 0 15732 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1523_
timestamp 1704896540
transform -1 0 18952 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1524_
timestamp 1704896540
transform 1 0 17480 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1525_
timestamp 1704896540
transform 1 0 17572 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_2  _1526_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 15364 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1527_
timestamp 1704896540
transform -1 0 13984 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1528_
timestamp 1704896540
transform 1 0 12512 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1529_
timestamp 1704896540
transform 1 0 11868 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1530_
timestamp 1704896540
transform -1 0 11684 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1531_
timestamp 1704896540
transform 1 0 9568 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1532_
timestamp 1704896540
transform 1 0 13340 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1533_
timestamp 1704896540
transform -1 0 11684 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1534_
timestamp 1704896540
transform -1 0 19964 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1535_
timestamp 1704896540
transform -1 0 19688 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1536_
timestamp 1704896540
transform 1 0 21252 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1537_
timestamp 1704896540
transform -1 0 20516 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1538_
timestamp 1704896540
transform 1 0 21252 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1539_
timestamp 1704896540
transform 1 0 21160 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1540_
timestamp 1704896540
transform 1 0 11960 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1541_
timestamp 1704896540
transform 1 0 26220 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1542_
timestamp 1704896540
transform -1 0 26220 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1543_
timestamp 1704896540
transform -1 0 25760 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1544_
timestamp 1704896540
transform 1 0 25024 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1545_
timestamp 1704896540
transform -1 0 25668 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1546_
timestamp 1704896540
transform 1 0 25024 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1547_
timestamp 1704896540
transform 1 0 26404 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1548_
timestamp 1704896540
transform 1 0 25116 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1549_
timestamp 1704896540
transform 1 0 26404 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1550_
timestamp 1704896540
transform 1 0 26864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1551_
timestamp 1704896540
transform -1 0 11040 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1552_
timestamp 1704896540
transform -1 0 26220 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1553_
timestamp 1704896540
transform -1 0 25760 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1554_
timestamp 1704896540
transform 1 0 25760 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1555_
timestamp 1704896540
transform -1 0 27048 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1556_
timestamp 1704896540
transform -1 0 26496 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1557_
timestamp 1704896540
transform 1 0 23920 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1558_
timestamp 1704896540
transform -1 0 24656 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1559_
timestamp 1704896540
transform 1 0 13524 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1560_
timestamp 1704896540
transform 1 0 25392 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1561_
timestamp 1704896540
transform -1 0 24288 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1562_
timestamp 1704896540
transform -1 0 25760 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1563_
timestamp 1704896540
transform 1 0 24748 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1564_
timestamp 1704896540
transform 1 0 24840 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1565_
timestamp 1704896540
transform 1 0 25392 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1566_
timestamp 1704896540
transform 1 0 26404 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1567_
timestamp 1704896540
transform 1 0 24288 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1568_
timestamp 1704896540
transform 1 0 23460 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1569_
timestamp 1704896540
transform 1 0 23460 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1570_
timestamp 1704896540
transform -1 0 24472 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1571_
timestamp 1704896540
transform -1 0 23276 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1572_
timestamp 1704896540
transform 1 0 22540 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1573_
timestamp 1704896540
transform 1 0 22540 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1574_
timestamp 1704896540
transform 1 0 23828 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1575_
timestamp 1704896540
transform 1 0 23828 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1576_
timestamp 1704896540
transform 1 0 24380 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1577_
timestamp 1704896540
transform -1 0 24932 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1578_
timestamp 1704896540
transform 1 0 23092 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1579_
timestamp 1704896540
transform 1 0 22908 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1580_
timestamp 1704896540
transform 1 0 22448 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1581_
timestamp 1704896540
transform 1 0 21804 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1582_
timestamp 1704896540
transform 1 0 22080 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1583_
timestamp 1704896540
transform -1 0 21896 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1584_
timestamp 1704896540
transform 1 0 21896 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _1585_
timestamp 1704896540
transform 1 0 20608 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1586_
timestamp 1704896540
transform 1 0 21252 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1587_
timestamp 1704896540
transform 1 0 20516 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1588_
timestamp 1704896540
transform -1 0 22264 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a21boi_1  _1589_
timestamp 1704896540
transform -1 0 22356 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1590_
timestamp 1704896540
transform -1 0 21804 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1591_
timestamp 1704896540
transform 1 0 20608 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1592_
timestamp 1704896540
transform 1 0 5796 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1593_
timestamp 1704896540
transform 1 0 20332 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1594_
timestamp 1704896540
transform -1 0 12604 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1595_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 16376 0 1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _1596_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 14076 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1597_
timestamp 1704896540
transform 1 0 15180 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1598_
timestamp 1704896540
transform 1 0 14904 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1599_
timestamp 1704896540
transform -1 0 15640 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1600_
timestamp 1704896540
transform 1 0 12604 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1601_
timestamp 1704896540
transform 1 0 12052 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1602_
timestamp 1704896540
transform 1 0 12512 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1603_
timestamp 1704896540
transform 1 0 16100 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1604_
timestamp 1704896540
transform 1 0 15364 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1605_
timestamp 1704896540
transform 1 0 16100 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1606_
timestamp 1704896540
transform 1 0 14168 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1607_
timestamp 1704896540
transform 1 0 13708 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1608_
timestamp 1704896540
transform 1 0 13984 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1609_
timestamp 1704896540
transform 1 0 13064 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1610_
timestamp 1704896540
transform -1 0 14076 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1611_
timestamp 1704896540
transform 1 0 1012 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1612_
timestamp 1704896540
transform 1 0 1196 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1613_
timestamp 1704896540
transform 1 0 1380 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1614_
timestamp 1704896540
transform -1 0 1380 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1615_
timestamp 1704896540
transform 1 0 3220 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1616_
timestamp 1704896540
transform 1 0 3312 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1617_
timestamp 1704896540
transform 1 0 2484 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1618_
timestamp 1704896540
transform -1 0 2760 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1619_
timestamp 1704896540
transform -1 0 2392 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1620_
timestamp 1704896540
transform -1 0 3036 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1621_
timestamp 1704896540
transform -1 0 2852 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1622_
timestamp 1704896540
transform 1 0 1380 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1623_
timestamp 1704896540
transform 1 0 1380 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1624_
timestamp 1704896540
transform -1 0 3036 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1625_
timestamp 1704896540
transform -1 0 3864 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1626_
timestamp 1704896540
transform 1 0 3956 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1627_
timestamp 1704896540
transform 1 0 4416 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1628_
timestamp 1704896540
transform 1 0 2484 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1629_
timestamp 1704896540
transform 1 0 2484 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1630_
timestamp 1704896540
transform -1 0 9292 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1631_
timestamp 1704896540
transform 1 0 8280 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1632_
timestamp 1704896540
transform 1 0 7820 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1633_
timestamp 1704896540
transform 1 0 8464 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1634_
timestamp 1704896540
transform -1 0 10396 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1635_
timestamp 1704896540
transform 1 0 9384 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1636_
timestamp 1704896540
transform 1 0 11500 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1637_
timestamp 1704896540
transform 1 0 11684 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1638_
timestamp 1704896540
transform 1 0 13432 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1639_
timestamp 1704896540
transform 1 0 14076 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1640_
timestamp 1704896540
transform -1 0 10120 0 -1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_2  _1641_
timestamp 1704896540
transform 1 0 9016 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1642_
timestamp 1704896540
transform -1 0 8648 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1643_
timestamp 1704896540
transform -1 0 9292 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1644_
timestamp 1704896540
transform -1 0 9476 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1645_
timestamp 1704896540
transform -1 0 10304 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1646_
timestamp 1704896540
transform 1 0 8280 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1647_
timestamp 1704896540
transform 1 0 10028 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1648_
timestamp 1704896540
transform 1 0 9476 0 -1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1649_
timestamp 1704896540
transform -1 0 9292 0 1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1650_
timestamp 1704896540
transform -1 0 18308 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _1651_
timestamp 1704896540
transform -1 0 15364 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1652_
timestamp 1704896540
transform 1 0 16652 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1653_
timestamp 1704896540
transform 1 0 17388 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1654_
timestamp 1704896540
transform 1 0 17388 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1655_
timestamp 1704896540
transform 1 0 19504 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1656_
timestamp 1704896540
transform 1 0 19320 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1657_
timestamp 1704896540
transform 1 0 19044 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1658_
timestamp 1704896540
transform 1 0 18676 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1659_
timestamp 1704896540
transform 1 0 19136 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1660_
timestamp 1704896540
transform 1 0 17940 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1661_
timestamp 1704896540
transform -1 0 18676 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1662_
timestamp 1704896540
transform 1 0 17020 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1663_
timestamp 1704896540
transform -1 0 16744 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1664_
timestamp 1704896540
transform 1 0 19412 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1665_
timestamp 1704896540
transform -1 0 20792 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1666_
timestamp 1704896540
transform 1 0 20516 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1667_
timestamp 1704896540
transform -1 0 14720 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1668_
timestamp 1704896540
transform -1 0 10856 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1669_
timestamp 1704896540
transform 1 0 9936 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1670_
timestamp 1704896540
transform 1 0 10948 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1671_
timestamp 1704896540
transform 1 0 8648 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1672_
timestamp 1704896540
transform -1 0 9936 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1673_
timestamp 1704896540
transform -1 0 9384 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1674_
timestamp 1704896540
transform 1 0 10120 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1675_
timestamp 1704896540
transform 1 0 8464 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1676_
timestamp 1704896540
transform -1 0 10488 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1677_
timestamp 1704896540
transform -1 0 12328 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1678_
timestamp 1704896540
transform -1 0 9292 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1679_
timestamp 1704896540
transform -1 0 13156 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1680_
timestamp 1704896540
transform -1 0 13984 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1681_
timestamp 1704896540
transform -1 0 12696 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1682_
timestamp 1704896540
transform 1 0 12236 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1683_
timestamp 1704896540
transform 1 0 12972 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1684_
timestamp 1704896540
transform 1 0 13892 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1685_
timestamp 1704896540
transform 1 0 12696 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1686_
timestamp 1704896540
transform -1 0 12788 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1687_
timestamp 1704896540
transform -1 0 12512 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1688_
timestamp 1704896540
transform 1 0 11960 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1689_
timestamp 1704896540
transform 1 0 13524 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1690_
timestamp 1704896540
transform 1 0 13524 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1691_
timestamp 1704896540
transform 1 0 12788 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1692_
timestamp 1704896540
transform -1 0 13892 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1693_
timestamp 1704896540
transform 1 0 12512 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1694_
timestamp 1704896540
transform -1 0 11684 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1695_
timestamp 1704896540
transform -1 0 18032 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1696_
timestamp 1704896540
transform 1 0 16652 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1697_
timestamp 1704896540
transform -1 0 17664 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1698_
timestamp 1704896540
transform -1 0 17204 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1699_
timestamp 1704896540
transform -1 0 19320 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1700_
timestamp 1704896540
transform -1 0 18952 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _1701_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 18032 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1702_
timestamp 1704896540
transform -1 0 19412 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1703_
timestamp 1704896540
transform -1 0 19044 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1704_
timestamp 1704896540
transform 1 0 17204 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__nor3b_1  _1705_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 16376 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1706_
timestamp 1704896540
transform 1 0 13340 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1707_
timestamp 1704896540
transform 1 0 13156 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1708_
timestamp 1704896540
transform -1 0 14444 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1709_
timestamp 1704896540
transform 1 0 13156 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1710_
timestamp 1704896540
transform 1 0 14260 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1711_
timestamp 1704896540
transform 1 0 14720 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1712_
timestamp 1704896540
transform 1 0 14812 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1713_
timestamp 1704896540
transform -1 0 15824 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1714_
timestamp 1704896540
transform 1 0 13892 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1715_
timestamp 1704896540
transform 1 0 13708 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1716_
timestamp 1704896540
transform 1 0 14352 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1717_
timestamp 1704896540
transform -1 0 15732 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1718_
timestamp 1704896540
transform 1 0 15732 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _1719_
timestamp 1704896540
transform 1 0 15456 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1720_
timestamp 1704896540
transform -1 0 15548 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1721_
timestamp 1704896540
transform -1 0 15548 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1722_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 14628 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1723_
timestamp 1704896540
transform 1 0 13524 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _1724_
timestamp 1704896540
transform -1 0 15180 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1725_
timestamp 1704896540
transform 1 0 15548 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1726_
timestamp 1704896540
transform 1 0 15088 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1727_
timestamp 1704896540
transform -1 0 16284 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1728_
timestamp 1704896540
transform 1 0 15180 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1729_
timestamp 1704896540
transform 1 0 15272 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1730_
timestamp 1704896540
transform -1 0 17664 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1731_
timestamp 1704896540
transform -1 0 16468 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1732_
timestamp 1704896540
transform 1 0 15548 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1733_
timestamp 1704896540
transform 1 0 14168 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_1  _1734_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 15548 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1735_
timestamp 1704896540
transform 1 0 15364 0 -1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1736_
timestamp 1704896540
transform 1 0 3864 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _1737_
timestamp 1704896540
transform -1 0 5888 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1738_
timestamp 1704896540
transform 1 0 3864 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1739_
timestamp 1704896540
transform 1 0 4784 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_1  _1740_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5152 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1741_
timestamp 1704896540
transform 1 0 5152 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1742_
timestamp 1704896540
transform 1 0 15824 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1743_
timestamp 1704896540
transform -1 0 16100 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1744_
timestamp 1704896540
transform 1 0 15732 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1745_
timestamp 1704896540
transform -1 0 4416 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1746_
timestamp 1704896540
transform -1 0 20700 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1747_
timestamp 1704896540
transform 1 0 15548 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1748_
timestamp 1704896540
transform 1 0 16284 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1749_
timestamp 1704896540
transform 1 0 16928 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1750_
timestamp 1704896540
transform -1 0 16928 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1751_
timestamp 1704896540
transform -1 0 14352 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1752_
timestamp 1704896540
transform 1 0 13616 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1753_
timestamp 1704896540
transform 1 0 13524 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1754_
timestamp 1704896540
transform 1 0 14168 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1755_
timestamp 1704896540
transform -1 0 12788 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1756_
timestamp 1704896540
transform -1 0 14536 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1757_
timestamp 1704896540
transform -1 0 13064 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1758_
timestamp 1704896540
transform -1 0 13708 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1759_
timestamp 1704896540
transform 1 0 12880 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1760_
timestamp 1704896540
transform 1 0 13708 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1761_
timestamp 1704896540
transform -1 0 15456 0 1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1762_
timestamp 1704896540
transform 1 0 14536 0 1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1763_
timestamp 1704896540
transform 1 0 14536 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1764_
timestamp 1704896540
transform -1 0 15732 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1765_
timestamp 1704896540
transform 1 0 14444 0 -1 29920
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1766_
timestamp 1704896540
transform 1 0 14168 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1767_
timestamp 1704896540
transform 1 0 14904 0 -1 29920
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1768_
timestamp 1704896540
transform 1 0 15088 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1769_
timestamp 1704896540
transform 1 0 15548 0 -1 29920
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1770_
timestamp 1704896540
transform 1 0 14904 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1771_
timestamp 1704896540
transform -1 0 17388 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1772_
timestamp 1704896540
transform -1 0 17204 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1773_
timestamp 1704896540
transform 1 0 16100 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1774_
timestamp 1704896540
transform 1 0 17388 0 1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1775_
timestamp 1704896540
transform 1 0 16744 0 1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1776_
timestamp 1704896540
transform -1 0 18308 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1777_
timestamp 1704896540
transform 1 0 16284 0 -1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1778_
timestamp 1704896540
transform 1 0 17480 0 -1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1779_
timestamp 1704896540
transform 1 0 16836 0 -1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1780_
timestamp 1704896540
transform -1 0 18952 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1781_
timestamp 1704896540
transform 1 0 16560 0 -1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1782_
timestamp 1704896540
transform 1 0 18216 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1783_
timestamp 1704896540
transform -1 0 17112 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1784_
timestamp 1704896540
transform 1 0 17296 0 1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1785_
timestamp 1704896540
transform 1 0 17020 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1786_
timestamp 1704896540
transform 1 0 17756 0 1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1787_
timestamp 1704896540
transform -1 0 19228 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1788_
timestamp 1704896540
transform -1 0 18584 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1789_
timestamp 1704896540
transform 1 0 17848 0 1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1790_
timestamp 1704896540
transform -1 0 18952 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1791_
timestamp 1704896540
transform 1 0 17756 0 -1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1792_
timestamp 1704896540
transform -1 0 18952 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1793_
timestamp 1704896540
transform 1 0 17940 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1794_
timestamp 1704896540
transform 1 0 25852 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1795_
timestamp 1704896540
transform -1 0 23644 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1796_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 22632 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1797_
timestamp 1704896540
transform -1 0 23736 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1798_
timestamp 1704896540
transform -1 0 23644 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1799_
timestamp 1704896540
transform -1 0 23000 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1800_
timestamp 1704896540
transform 1 0 23828 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1801_
timestamp 1704896540
transform 1 0 23184 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1802_
timestamp 1704896540
transform 1 0 24012 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1803_
timestamp 1704896540
transform 1 0 25208 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1804_
timestamp 1704896540
transform 1 0 23828 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _1805_
timestamp 1704896540
transform -1 0 25208 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1806_
timestamp 1704896540
transform 1 0 22172 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1807_
timestamp 1704896540
transform -1 0 24104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _1808_
timestamp 1704896540
transform -1 0 23092 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1809_
timestamp 1704896540
transform 1 0 22080 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1810_
timestamp 1704896540
transform -1 0 23552 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1811_
timestamp 1704896540
transform -1 0 24104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1812_
timestamp 1704896540
transform -1 0 25208 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1813_
timestamp 1704896540
transform 1 0 22172 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1814_
timestamp 1704896540
transform -1 0 23552 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_1  _1815_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 23644 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1816_
timestamp 1704896540
transform 1 0 23000 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1817_
timestamp 1704896540
transform -1 0 23276 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1818_
timestamp 1704896540
transform -1 0 23000 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1819_
timestamp 1704896540
transform -1 0 22632 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1820_
timestamp 1704896540
transform -1 0 24656 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1821_
timestamp 1704896540
transform 1 0 21988 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1822_
timestamp 1704896540
transform -1 0 23276 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1823_
timestamp 1704896540
transform 1 0 22632 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1824_
timestamp 1704896540
transform 1 0 22080 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1825_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 23092 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _1826_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 23000 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1827_
timestamp 1704896540
transform 1 0 23368 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _1828_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 22448 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1829_
timestamp 1704896540
transform -1 0 24104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1830_
timestamp 1704896540
transform 1 0 22724 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1831_
timestamp 1704896540
transform 1 0 19504 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1832_
timestamp 1704896540
transform 1 0 19964 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1833_
timestamp 1704896540
transform 1 0 23644 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1834_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 24012 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1835_
timestamp 1704896540
transform 1 0 24472 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1836_
timestamp 1704896540
transform 1 0 25116 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1837_
timestamp 1704896540
transform 1 0 23276 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1838_
timestamp 1704896540
transform 1 0 23828 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1839_
timestamp 1704896540
transform 1 0 23276 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1840_
timestamp 1704896540
transform 1 0 23460 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1841_
timestamp 1704896540
transform 1 0 24380 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1842_
timestamp 1704896540
transform 1 0 24104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1843_
timestamp 1704896540
transform 1 0 25024 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1844_
timestamp 1704896540
transform -1 0 25944 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1845_
timestamp 1704896540
transform -1 0 24196 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1846_
timestamp 1704896540
transform 1 0 24748 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1847_
timestamp 1704896540
transform 1 0 25208 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1848_
timestamp 1704896540
transform -1 0 25944 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1849_
timestamp 1704896540
transform 1 0 24748 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1850_
timestamp 1704896540
transform 1 0 24012 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1851_
timestamp 1704896540
transform 1 0 24196 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1852_
timestamp 1704896540
transform -1 0 25852 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1853_
timestamp 1704896540
transform -1 0 24748 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1854_
timestamp 1704896540
transform -1 0 25484 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1855_
timestamp 1704896540
transform 1 0 24288 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1856_
timestamp 1704896540
transform -1 0 25576 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1857_
timestamp 1704896540
transform 1 0 24380 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1858_
timestamp 1704896540
transform 1 0 24380 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1859_
timestamp 1704896540
transform 1 0 24656 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1860_
timestamp 1704896540
transform -1 0 25668 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1861_
timestamp 1704896540
transform -1 0 24380 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1862_
timestamp 1704896540
transform 1 0 25116 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1863_
timestamp 1704896540
transform 1 0 25576 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1864_
timestamp 1704896540
transform -1 0 26312 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1865_
timestamp 1704896540
transform -1 0 24932 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1866_
timestamp 1704896540
transform -1 0 24104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1867_
timestamp 1704896540
transform 1 0 24932 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1868_
timestamp 1704896540
transform 1 0 26404 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1869_
timestamp 1704896540
transform -1 0 24748 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1870_
timestamp 1704896540
transform -1 0 25300 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1871_
timestamp 1704896540
transform 1 0 24104 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1872_
timestamp 1704896540
transform -1 0 26680 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1873_
timestamp 1704896540
transform -1 0 25116 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1874_
timestamp 1704896540
transform -1 0 24840 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_1  _1875_
timestamp 1704896540
transform 1 0 23460 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1876_
timestamp 1704896540
transform -1 0 24748 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1877_
timestamp 1704896540
transform 1 0 23644 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1878_
timestamp 1704896540
transform -1 0 26312 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1879_
timestamp 1704896540
transform 1 0 23920 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1880_
timestamp 1704896540
transform -1 0 24932 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1881_
timestamp 1704896540
transform 1 0 23460 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _1882_
timestamp 1704896540
transform -1 0 24564 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1883_
timestamp 1704896540
transform 1 0 24564 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1884_
timestamp 1704896540
transform -1 0 24288 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1885_
timestamp 1704896540
transform -1 0 25300 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__nor3b_1  _1886_
timestamp 1704896540
transform 1 0 24564 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1887_
timestamp 1704896540
transform 1 0 23000 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1888_
timestamp 1704896540
transform 1 0 23184 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1889_
timestamp 1704896540
transform 1 0 22356 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1890_
timestamp 1704896540
transform 1 0 23828 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1891_
timestamp 1704896540
transform 1 0 21988 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1892_
timestamp 1704896540
transform 1 0 22540 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1893_
timestamp 1704896540
transform 1 0 21620 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1894_
timestamp 1704896540
transform -1 0 23644 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1895_
timestamp 1704896540
transform 1 0 22356 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1896_
timestamp 1704896540
transform -1 0 23736 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1897_
timestamp 1704896540
transform 1 0 23736 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1898_
timestamp 1704896540
transform -1 0 24564 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1899_
timestamp 1704896540
transform -1 0 25024 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _1900_
timestamp 1704896540
transform 1 0 24288 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1901_
timestamp 1704896540
transform 1 0 25576 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1902_
timestamp 1704896540
transform -1 0 25576 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1903_
timestamp 1704896540
transform 1 0 23460 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1904_
timestamp 1704896540
transform 1 0 23368 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _1905_
timestamp 1704896540
transform 1 0 22724 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1906_
timestamp 1704896540
transform 1 0 24472 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1907_
timestamp 1704896540
transform -1 0 24472 0 1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1908_
timestamp 1704896540
transform -1 0 25024 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1909_
timestamp 1704896540
transform 1 0 23828 0 1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1910_
timestamp 1704896540
transform 1 0 23828 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1911_
timestamp 1704896540
transform 1 0 24840 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1912_
timestamp 1704896540
transform -1 0 24104 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1913_
timestamp 1704896540
transform 1 0 23460 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1914_
timestamp 1704896540
transform 1 0 22540 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_1  _1915_
timestamp 1704896540
transform -1 0 23460 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1916_
timestamp 1704896540
transform -1 0 24840 0 1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1917_
timestamp 1704896540
transform 1 0 23828 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1918_
timestamp 1704896540
transform -1 0 21896 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1919_
timestamp 1704896540
transform -1 0 21160 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1920_
timestamp 1704896540
transform 1 0 21252 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1921_
timestamp 1704896540
transform 1 0 23828 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1922_
timestamp 1704896540
transform -1 0 24564 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1923_
timestamp 1704896540
transform -1 0 22080 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1924_
timestamp 1704896540
transform 1 0 21712 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1925_
timestamp 1704896540
transform 1 0 21712 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1926_
timestamp 1704896540
transform -1 0 21712 0 -1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1927_
timestamp 1704896540
transform 1 0 20700 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1928_
timestamp 1704896540
transform 1 0 23000 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1929_
timestamp 1704896540
transform -1 0 21436 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1930_
timestamp 1704896540
transform 1 0 21988 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1931_
timestamp 1704896540
transform -1 0 22264 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1932_
timestamp 1704896540
transform 1 0 21436 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1933_
timestamp 1704896540
transform -1 0 22356 0 1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1934_
timestamp 1704896540
transform 1 0 21436 0 1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1935_
timestamp 1704896540
transform 1 0 22356 0 1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1936_
timestamp 1704896540
transform 1 0 22356 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1937_
timestamp 1704896540
transform 1 0 22908 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1938_
timestamp 1704896540
transform 1 0 24564 0 1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1939_
timestamp 1704896540
transform 1 0 25300 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1940_
timestamp 1704896540
transform -1 0 25300 0 -1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1941_
timestamp 1704896540
transform -1 0 24840 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1942_
timestamp 1704896540
transform -1 0 25668 0 -1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1943_
timestamp 1704896540
transform -1 0 25944 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1944_
timestamp 1704896540
transform 1 0 25024 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1945_
timestamp 1704896540
transform -1 0 26128 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1946_
timestamp 1704896540
transform 1 0 24564 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1947_
timestamp 1704896540
transform -1 0 25024 0 1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1948_
timestamp 1704896540
transform 1 0 24932 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1949_
timestamp 1704896540
transform 1 0 26036 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1950_
timestamp 1704896540
transform -1 0 26036 0 -1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1951_
timestamp 1704896540
transform 1 0 26404 0 -1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1952_
timestamp 1704896540
transform 1 0 25024 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1953_
timestamp 1704896540
transform 1 0 26864 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1954_
timestamp 1704896540
transform 1 0 24932 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1955_
timestamp 1704896540
transform -1 0 25668 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1956_
timestamp 1704896540
transform -1 0 25576 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1957_
timestamp 1704896540
transform 1 0 26404 0 -1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1958_
timestamp 1704896540
transform 1 0 25944 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1959_
timestamp 1704896540
transform -1 0 26036 0 -1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1960_
timestamp 1704896540
transform -1 0 25668 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1961_
timestamp 1704896540
transform 1 0 26864 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1962_
timestamp 1704896540
transform -1 0 26864 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1963_
timestamp 1704896540
transform 1 0 26864 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1964_
timestamp 1704896540
transform 1 0 26404 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1965_
timestamp 1704896540
transform 1 0 26864 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1966_
timestamp 1704896540
transform 1 0 25668 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1967_
timestamp 1704896540
transform 1 0 16192 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1968_
timestamp 1704896540
transform -1 0 16652 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1969_
timestamp 1704896540
transform 1 0 16100 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1970_
timestamp 1704896540
transform -1 0 16284 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1971_
timestamp 1704896540
transform -1 0 15640 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1972_
timestamp 1704896540
transform 1 0 14904 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1973_
timestamp 1704896540
transform 1 0 14720 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1974_
timestamp 1704896540
transform 1 0 15548 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1975_
timestamp 1704896540
transform 1 0 15824 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1976_
timestamp 1704896540
transform -1 0 15548 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1977_
timestamp 1704896540
transform 1 0 14628 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1978_
timestamp 1704896540
transform 1 0 15180 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1979_
timestamp 1704896540
transform 1 0 14076 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1980_
timestamp 1704896540
transform 1 0 14628 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1981_
timestamp 1704896540
transform 1 0 14536 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1982_
timestamp 1704896540
transform 1 0 14352 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nor2b_2  _1983_
timestamp 1704896540
transform 1 0 11684 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1984_
timestamp 1704896540
transform 1 0 4968 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1985_
timestamp 1704896540
transform 1 0 5428 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1986_
timestamp 1704896540
transform -1 0 10948 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1987_
timestamp 1704896540
transform -1 0 11224 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1988_
timestamp 1704896540
transform 1 0 12512 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1989_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10948 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1990_
timestamp 1704896540
transform 1 0 8924 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1991_
timestamp 1704896540
transform -1 0 9476 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1992_
timestamp 1704896540
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1993_
timestamp 1704896540
transform 1 0 9936 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1994_
timestamp 1704896540
transform -1 0 10672 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__nor2b_2  _1995_
timestamp 1704896540
transform 1 0 6900 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1996_
timestamp 1704896540
transform 1 0 5888 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1997_
timestamp 1704896540
transform 1 0 6440 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1998_
timestamp 1704896540
transform 1 0 8464 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1999_
timestamp 1704896540
transform -1 0 8924 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2000_
timestamp 1704896540
transform 1 0 9016 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2001_
timestamp 1704896540
transform 1 0 10304 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _2002_
timestamp 1704896540
transform -1 0 8464 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2003_
timestamp 1704896540
transform 1 0 8372 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _2004_
timestamp 1704896540
transform -1 0 7728 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _2005_
timestamp 1704896540
transform 1 0 6808 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2006_
timestamp 1704896540
transform 1 0 7636 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2007_
timestamp 1704896540
transform 1 0 7912 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _2008_
timestamp 1704896540
transform 1 0 9108 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2009_
timestamp 1704896540
transform 1 0 10488 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2010_
timestamp 1704896540
transform -1 0 8372 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _2011_
timestamp 1704896540
transform 1 0 7728 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2012_
timestamp 1704896540
transform -1 0 5704 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2013_
timestamp 1704896540
transform 1 0 6348 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2014_
timestamp 1704896540
transform 1 0 6624 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_1  _2015_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6348 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _2016_
timestamp 1704896540
transform 1 0 6808 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _2017_
timestamp 1704896540
transform -1 0 4600 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _2018_
timestamp 1704896540
transform -1 0 6348 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _2019_
timestamp 1704896540
transform -1 0 3404 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2020_
timestamp 1704896540
transform -1 0 7544 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2021_
timestamp 1704896540
transform -1 0 6348 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2022_
timestamp 1704896540
transform -1 0 7636 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2023_
timestamp 1704896540
transform -1 0 5704 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2024_
timestamp 1704896540
transform 1 0 4140 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2025_
timestamp 1704896540
transform 1 0 4600 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2026_
timestamp 1704896540
transform 1 0 3312 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2027_
timestamp 1704896540
transform 1 0 3956 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2028_
timestamp 1704896540
transform 1 0 7544 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2029_
timestamp 1704896540
transform 1 0 6348 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2030_
timestamp 1704896540
transform -1 0 7544 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2031_
timestamp 1704896540
transform 1 0 4876 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2032_
timestamp 1704896540
transform -1 0 3864 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2033_
timestamp 1704896540
transform -1 0 4140 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2034_
timestamp 1704896540
transform -1 0 3680 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _2035_
timestamp 1704896540
transform -1 0 2668 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _2036_
timestamp 1704896540
transform -1 0 2668 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2037_
timestamp 1704896540
transform -1 0 3036 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2038_
timestamp 1704896540
transform -1 0 3128 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2039_
timestamp 1704896540
transform -1 0 1472 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2040_
timestamp 1704896540
transform 1 0 1472 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2041_
timestamp 1704896540
transform 1 0 1012 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2042_
timestamp 1704896540
transform -1 0 2208 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2043_
timestamp 1704896540
transform 1 0 1196 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2044_
timestamp 1704896540
transform -1 0 3036 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2045_
timestamp 1704896540
transform -1 0 3680 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2046_
timestamp 1704896540
transform 1 0 920 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2047_
timestamp 1704896540
transform 1 0 1012 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2048_
timestamp 1704896540
transform 1 0 1748 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2049_
timestamp 1704896540
transform 1 0 1012 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2050_
timestamp 1704896540
transform -1 0 3312 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2051_
timestamp 1704896540
transform 1 0 6256 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2052_
timestamp 1704896540
transform -1 0 3956 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _2053_
timestamp 1704896540
transform 1 0 2944 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2054_
timestamp 1704896540
transform 1 0 3404 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2055_
timestamp 1704896540
transform 1 0 5796 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2056_
timestamp 1704896540
transform 1 0 6624 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _2057_
timestamp 1704896540
transform 1 0 3956 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2058_
timestamp 1704896540
transform -1 0 5428 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _2059_
timestamp 1704896540
transform 1 0 7084 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2060_
timestamp 1704896540
transform -1 0 7084 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _2061_
timestamp 1704896540
transform -1 0 19780 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_2  _2062_
timestamp 1704896540
transform -1 0 19688 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2063_
timestamp 1704896540
transform -1 0 20608 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2064_
timestamp 1704896540
transform -1 0 21068 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2065_
timestamp 1704896540
transform -1 0 20332 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2066_
timestamp 1704896540
transform 1 0 17940 0 1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2067_
timestamp 1704896540
transform -1 0 23368 0 1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2068_
timestamp 1704896540
transform 1 0 18952 0 1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2069_
timestamp 1704896540
transform -1 0 19872 0 -1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2070_
timestamp 1704896540
transform -1 0 23736 0 -1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2071_
timestamp 1704896540
transform -1 0 10304 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2072_
timestamp 1704896540
transform 1 0 8096 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2073_
timestamp 1704896540
transform 1 0 9200 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_1  _2074_
timestamp 1704896540
transform 1 0 6072 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _2075_
timestamp 1704896540
transform -1 0 9936 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _2076_
timestamp 1704896540
transform 1 0 9016 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2077_
timestamp 1704896540
transform 1 0 9292 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2078_
timestamp 1704896540
transform -1 0 10580 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2079_
timestamp 1704896540
transform 1 0 10580 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _2080_
timestamp 1704896540
transform -1 0 7084 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _2081_
timestamp 1704896540
transform 1 0 5796 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _2082_
timestamp 1704896540
transform 1 0 5152 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2083_
timestamp 1704896540
transform -1 0 6716 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _2084_
timestamp 1704896540
transform 1 0 5796 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _2085_
timestamp 1704896540
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _2086_
timestamp 1704896540
transform -1 0 7912 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _2087_
timestamp 1704896540
transform -1 0 8188 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _2088_
timestamp 1704896540
transform 1 0 6624 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2089_
timestamp 1704896540
transform 1 0 6900 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2090_
timestamp 1704896540
transform -1 0 8004 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2091_
timestamp 1704896540
transform 1 0 5796 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2092_
timestamp 1704896540
transform -1 0 7084 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _2093_
timestamp 1704896540
transform -1 0 6992 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2094_
timestamp 1704896540
transform 1 0 4876 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _2095_
timestamp 1704896540
transform 1 0 6992 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _2096_
timestamp 1704896540
transform -1 0 7452 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2097_
timestamp 1704896540
transform -1 0 8280 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _2098_
timestamp 1704896540
transform 1 0 7452 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2099_
timestamp 1704896540
transform -1 0 8464 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _2100_
timestamp 1704896540
transform -1 0 7728 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2101_
timestamp 1704896540
transform 1 0 6808 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2102_
timestamp 1704896540
transform 1 0 7728 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2103_
timestamp 1704896540
transform -1 0 7820 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _2104_
timestamp 1704896540
transform 1 0 5980 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2105_
timestamp 1704896540
transform -1 0 8648 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2106_
timestamp 1704896540
transform -1 0 8740 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _2107_
timestamp 1704896540
transform 1 0 7636 0 1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2108_
timestamp 1704896540
transform -1 0 9752 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _2109_
timestamp 1704896540
transform -1 0 8188 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__a221oi_2  _2110_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7268 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _2111_
timestamp 1704896540
transform -1 0 8648 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _2112_
timestamp 1704896540
transform -1 0 6992 0 1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2113_
timestamp 1704896540
transform -1 0 7820 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  _2114_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6808 0 -1 29920
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2115_
timestamp 1704896540
transform -1 0 8096 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2116_
timestamp 1704896540
transform 1 0 6072 0 -1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2117_
timestamp 1704896540
transform -1 0 10580 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2118_
timestamp 1704896540
transform -1 0 8188 0 1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2119_
timestamp 1704896540
transform -1 0 8740 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2120_
timestamp 1704896540
transform -1 0 8832 0 1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _2121_
timestamp 1704896540
transform 1 0 7452 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _2122_
timestamp 1704896540
transform -1 0 8096 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2123_
timestamp 1704896540
transform -1 0 8648 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _2124_
timestamp 1704896540
transform -1 0 7820 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _2125_
timestamp 1704896540
transform 1 0 6532 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _2126_
timestamp 1704896540
transform 1 0 7268 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2127_
timestamp 1704896540
transform -1 0 7544 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _2128_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6716 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2129_
timestamp 1704896540
transform -1 0 7544 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _2130_
timestamp 1704896540
transform 1 0 6992 0 1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2131_
timestamp 1704896540
transform 1 0 6624 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _2132_
timestamp 1704896540
transform -1 0 8004 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2133_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10948 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2134_
timestamp 1704896540
transform -1 0 17572 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2135_
timestamp 1704896540
transform -1 0 18124 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2136_
timestamp 1704896540
transform 1 0 17940 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2137_
timestamp 1704896540
transform 1 0 17940 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2138_
timestamp 1704896540
transform 1 0 18952 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2139_
timestamp 1704896540
transform 1 0 17296 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2140_
timestamp 1704896540
transform 1 0 20332 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2141_
timestamp 1704896540
transform 1 0 17204 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2142_
timestamp 1704896540
transform 1 0 20424 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2143_
timestamp 1704896540
transform 1 0 18860 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2144_
timestamp 1704896540
transform 1 0 18860 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2145_
timestamp 1704896540
transform -1 0 22356 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2146_
timestamp 1704896540
transform 1 0 13892 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2147_
timestamp 1704896540
transform 1 0 17020 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2148_
timestamp 1704896540
transform 1 0 17572 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2149_
timestamp 1704896540
transform 1 0 13800 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2150_
timestamp 1704896540
transform 1 0 15732 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2151_
timestamp 1704896540
transform 1 0 17020 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2152_
timestamp 1704896540
transform -1 0 12512 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2153_
timestamp 1704896540
transform 1 0 10304 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2154_
timestamp 1704896540
transform -1 0 13340 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2155_
timestamp 1704896540
transform -1 0 13432 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2156_
timestamp 1704896540
transform -1 0 12420 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2157_
timestamp 1704896540
transform 1 0 21896 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2158_
timestamp 1704896540
transform 1 0 19780 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2159_
timestamp 1704896540
transform 1 0 21804 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2160_
timestamp 1704896540
transform 1 0 21896 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2161_
timestamp 1704896540
transform 1 0 24472 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2162_
timestamp 1704896540
transform -1 0 27140 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2163_
timestamp 1704896540
transform 1 0 24196 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2164_
timestamp 1704896540
transform -1 0 26312 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2165_
timestamp 1704896540
transform 1 0 22264 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2166_
timestamp 1704896540
transform -1 0 26036 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2167_
timestamp 1704896540
transform 1 0 19688 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2168_
timestamp 1704896540
transform -1 0 22724 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2169_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2392 0 -1 31008
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2170_
timestamp 1704896540
transform -1 0 16284 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2171_
timestamp 1704896540
transform 1 0 11776 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2172_
timestamp 1704896540
transform 1 0 15824 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2173_
timestamp 1704896540
transform 1 0 13708 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2174_
timestamp 1704896540
transform 1 0 11592 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2175_
timestamp 1704896540
transform 1 0 828 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2176_
timestamp 1704896540
transform 1 0 828 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2177_
timestamp 1704896540
transform 1 0 3588 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2178_
timestamp 1704896540
transform 1 0 2392 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2179_
timestamp 1704896540
transform 1 0 828 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2180_
timestamp 1704896540
transform -1 0 4692 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2181_
timestamp 1704896540
transform 1 0 1012 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2182_
timestamp 1704896540
transform 1 0 6716 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2183_
timestamp 1704896540
transform 1 0 6808 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2184_
timestamp 1704896540
transform 1 0 9016 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2185_
timestamp 1704896540
transform -1 0 10856 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2186_
timestamp 1704896540
transform 1 0 7912 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2187_
timestamp 1704896540
transform 1 0 8648 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2188_
timestamp 1704896540
transform -1 0 10396 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2189_
timestamp 1704896540
transform 1 0 9476 0 1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2190_
timestamp 1704896540
transform 1 0 8648 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2191_
timestamp 1704896540
transform 1 0 10948 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2192_
timestamp 1704896540
transform -1 0 11592 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2193_
timestamp 1704896540
transform -1 0 10028 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2194_
timestamp 1704896540
transform 1 0 17112 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2195_
timestamp 1704896540
transform 1 0 18952 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2196_
timestamp 1704896540
transform 1 0 17664 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2197_
timestamp 1704896540
transform 1 0 16744 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2198_
timestamp 1704896540
transform -1 0 20700 0 1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2199_
timestamp 1704896540
transform -1 0 9384 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2200_
timestamp 1704896540
transform -1 0 10856 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2201_
timestamp 1704896540
transform 1 0 8648 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2202_
timestamp 1704896540
transform -1 0 11500 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2203_
timestamp 1704896540
transform -1 0 9568 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2204_
timestamp 1704896540
transform 1 0 9936 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2205_
timestamp 1704896540
transform -1 0 10856 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2206_
timestamp 1704896540
transform -1 0 9844 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2207_
timestamp 1704896540
transform 1 0 11224 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2208_
timestamp 1704896540
transform 1 0 12420 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2209_
timestamp 1704896540
transform 1 0 11040 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2210_
timestamp 1704896540
transform 1 0 12512 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2211_
timestamp 1704896540
transform 1 0 11868 0 -1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2212_
timestamp 1704896540
transform -1 0 17572 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2213_
timestamp 1704896540
transform -1 0 16008 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2214_
timestamp 1704896540
transform -1 0 14536 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2215_
timestamp 1704896540
transform 1 0 11684 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2216_
timestamp 1704896540
transform -1 0 16652 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2217_
timestamp 1704896540
transform 1 0 13800 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2218_
timestamp 1704896540
transform -1 0 18492 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2219_
timestamp 1704896540
transform -1 0 18952 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2220_
timestamp 1704896540
transform -1 0 19412 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2221_
timestamp 1704896540
transform 1 0 17112 0 1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2222_
timestamp 1704896540
transform -1 0 19688 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2223_
timestamp 1704896540
transform -1 0 19872 0 -1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2224_
timestamp 1704896540
transform 1 0 18676 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2225_
timestamp 1704896540
transform -1 0 20240 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2226_
timestamp 1704896540
transform 1 0 25668 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2227_
timestamp 1704896540
transform 1 0 22908 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2228_
timestamp 1704896540
transform -1 0 26864 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2229_
timestamp 1704896540
transform 1 0 25668 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2230_
timestamp 1704896540
transform 1 0 25484 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2231_
timestamp 1704896540
transform -1 0 26864 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2232_
timestamp 1704896540
transform -1 0 27048 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2233_
timestamp 1704896540
transform -1 0 27048 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2234_
timestamp 1704896540
transform -1 0 26312 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2235_
timestamp 1704896540
transform -1 0 26956 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2236_
timestamp 1704896540
transform 1 0 24840 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2237_
timestamp 1704896540
transform 1 0 23644 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2238_
timestamp 1704896540
transform -1 0 21068 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2239_
timestamp 1704896540
transform 1 0 21896 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2240_
timestamp 1704896540
transform 1 0 20240 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2241_
timestamp 1704896540
transform 1 0 21252 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2242_
timestamp 1704896540
transform 1 0 22264 0 1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2243_
timestamp 1704896540
transform -1 0 26772 0 1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2244_
timestamp 1704896540
transform -1 0 27140 0 1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2245_
timestamp 1704896540
transform -1 0 26312 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2246_
timestamp 1704896540
transform -1 0 27140 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2247_
timestamp 1704896540
transform 1 0 25576 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2248_
timestamp 1704896540
transform 1 0 25668 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2249_
timestamp 1704896540
transform -1 0 27140 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2250_
timestamp 1704896540
transform -1 0 26312 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2251_
timestamp 1704896540
transform -1 0 17296 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2252_
timestamp 1704896540
transform 1 0 14444 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2253_
timestamp 1704896540
transform -1 0 17572 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2254_
timestamp 1704896540
transform 1 0 13708 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2255_
timestamp 1704896540
transform 1 0 13984 0 -1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2256_
timestamp 1704896540
transform 1 0 4600 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2257_
timestamp 1704896540
transform 1 0 6164 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2258_
timestamp 1704896540
transform -1 0 10304 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2259_
timestamp 1704896540
transform 1 0 6348 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2260_
timestamp 1704896540
transform -1 0 10488 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2261_
timestamp 1704896540
transform 1 0 8372 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2262_
timestamp 1704896540
transform 1 0 5980 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2263_
timestamp 1704896540
transform 1 0 5888 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2264_
timestamp 1704896540
transform -1 0 7636 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2265_
timestamp 1704896540
transform 1 0 5336 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2266_
timestamp 1704896540
transform 1 0 3496 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2267_
timestamp 1704896540
transform 1 0 5980 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2268_
timestamp 1704896540
transform 1 0 4508 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2269_
timestamp 1704896540
transform 1 0 3864 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2270_
timestamp 1704896540
transform 1 0 2116 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2271_
timestamp 1704896540
transform 1 0 2668 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2272_
timestamp 1704896540
transform 1 0 828 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2273_
timestamp 1704896540
transform -1 0 3128 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2274_
timestamp 1704896540
transform -1 0 2300 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2275_
timestamp 1704896540
transform 1 0 828 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2276_
timestamp 1704896540
transform 1 0 1656 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2277_
timestamp 1704896540
transform -1 0 4692 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2278_
timestamp 1704896540
transform 1 0 3220 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2279_
timestamp 1704896540
transform -1 0 6256 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2280_
timestamp 1704896540
transform 1 0 19688 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2281_
timestamp 1704896540
transform 1 0 20148 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2282_
timestamp 1704896540
transform 1 0 19504 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2283_
timestamp 1704896540
transform 1 0 19504 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2284_
timestamp 1704896540
transform 1 0 21252 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2285_
timestamp 1704896540
transform 1 0 19412 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2286_
timestamp 1704896540
transform 1 0 19320 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2287_
timestamp 1704896540
transform -1 0 22724 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2288_
timestamp 1704896540
transform 1 0 9936 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2289_
timestamp 1704896540
transform 1 0 5520 0 1 20128
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2290_
timestamp 1704896540
transform 1 0 3680 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2291_
timestamp 1704896540
transform 1 0 3404 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2292_
timestamp 1704896540
transform 1 0 828 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2293_
timestamp 1704896540
transform 1 0 3220 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2294_
timestamp 1704896540
transform 1 0 828 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2295_
timestamp 1704896540
transform 1 0 828 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2296_
timestamp 1704896540
transform 1 0 920 0 -1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2297_
timestamp 1704896540
transform 1 0 3220 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2298_
timestamp 1704896540
transform 1 0 4968 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2299_
timestamp 1704896540
transform 1 0 5796 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2300_
timestamp 1704896540
transform 1 0 2208 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2301_
timestamp 1704896540
transform 1 0 1840 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2302_
timestamp 1704896540
transform 1 0 3312 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2303_
timestamp 1704896540
transform 1 0 5796 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2304_
timestamp 1704896540
transform 1 0 6164 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2305_
timestamp 1704896540
transform 1 0 3956 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2306_
timestamp 1704896540
transform 1 0 6808 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2307_
timestamp 1704896540
transform 1 0 7176 0 -1 10336
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2308_
timestamp 1704896540
transform 1 0 6716 0 1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2309_
timestamp 1704896540
transform 1 0 9200 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2310_
timestamp 1704896540
transform -1 0 10856 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2311_
timestamp 1704896540
transform 1 0 21252 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2312_
timestamp 1704896540
transform 1 0 21436 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2313_
timestamp 1704896540
transform 1 0 21068 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2314_
timestamp 1704896540
transform 1 0 21252 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _2315__61 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8648 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2315_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8004 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2316__62
timestamp 1704896540
transform -1 0 8188 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2316_
timestamp 1704896540
transform 1 0 6808 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_2  _2317_
timestamp 1704896540
transform 1 0 7084 0 1 544
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2317__63
timestamp 1704896540
transform 1 0 6532 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2318_
timestamp 1704896540
transform 1 0 6716 0 1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2318__64
timestamp 1704896540
transform -1 0 7268 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2319__65
timestamp 1704896540
transform -1 0 6532 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2319_
timestamp 1704896540
transform 1 0 5888 0 1 544
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_2  _2320_
timestamp 1704896540
transform 1 0 5520 0 1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2320__66
timestamp 1704896540
transform -1 0 6072 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2321__67
timestamp 1704896540
transform -1 0 5520 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2321_
timestamp 1704896540
transform 1 0 4508 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_2  _2322_
timestamp 1704896540
transform 1 0 4416 0 1 544
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2322__68
timestamp 1704896540
transform 1 0 3772 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2323_
timestamp 1704896540
transform 1 0 4048 0 1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2323__69
timestamp 1704896540
transform -1 0 4324 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2324__70
timestamp 1704896540
transform -1 0 3496 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2324_
timestamp 1704896540
transform 1 0 3312 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_2  _2325_
timestamp 1704896540
transform 1 0 3220 0 1 544
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2325__71
timestamp 1704896540
transform 1 0 2852 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2326__72
timestamp 1704896540
transform -1 0 2484 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2326_
timestamp 1704896540
transform 1 0 2116 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_2  _2327_
timestamp 1704896540
transform 1 0 1840 0 1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2327__73
timestamp 1704896540
transform 1 0 1564 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2328_
timestamp 1704896540
transform 1 0 920 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2328__74
timestamp 1704896540
transform -1 0 1564 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2329__75
timestamp 1704896540
transform -1 0 1196 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2329_
timestamp 1704896540
transform 1 0 920 0 1 544
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_1  _2330_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7176 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2330__76
timestamp 1704896540
transform -1 0 7728 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2331__77
timestamp 1704896540
transform -1 0 7360 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _2331_
timestamp 1704896540
transform 1 0 6992 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2332__78
timestamp 1704896540
transform -1 0 7176 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _2332_
timestamp 1704896540
transform 1 0 6624 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _2333_
timestamp 1704896540
transform 1 0 5796 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2333__79
timestamp 1704896540
transform 1 0 5612 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _2334_
timestamp 1704896540
transform -1 0 5612 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2334__80
timestamp 1704896540
transform 1 0 4600 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _2335_
timestamp 1704896540
transform 1 0 2668 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2335__81
timestamp 1704896540
transform -1 0 2944 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2336__82
timestamp 1704896540
transform -1 0 1564 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _2336_
timestamp 1704896540
transform 1 0 1196 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2337__83
timestamp 1704896540
transform 1 0 920 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _2337_
timestamp 1704896540
transform 1 0 1196 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_2  _2338_
timestamp 1704896540
transform 1 0 17296 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2338__38
timestamp 1704896540
transform 1 0 16652 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2339__39
timestamp 1704896540
transform -1 0 16652 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2339_
timestamp 1704896540
transform 1 0 16192 0 1 544
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2340__40
timestamp 1704896540
transform 1 0 15548 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2340_
timestamp 1704896540
transform 1 0 16100 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_2  _2341_
timestamp 1704896540
transform 1 0 15180 0 1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2341__41
timestamp 1704896540
transform 1 0 14904 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2342_
timestamp 1704896540
transform 1 0 14628 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2342__42
timestamp 1704896540
transform -1 0 14904 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2343_
timestamp 1704896540
transform 1 0 14076 0 1 544
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2343__43
timestamp 1704896540
transform -1 0 14444 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2344_
timestamp 1704896540
transform 1 0 13432 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2344__44
timestamp 1704896540
transform -1 0 13800 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2345_
timestamp 1704896540
transform 1 0 12236 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2345__45
timestamp 1704896540
transform -1 0 13156 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2346_
timestamp 1704896540
transform 1 0 12236 0 1 544
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2346__46
timestamp 1704896540
transform -1 0 13432 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2347_
timestamp 1704896540
transform 1 0 11684 0 1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2347__47
timestamp 1704896540
transform -1 0 11960 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2348__48
timestamp 1704896540
transform -1 0 11500 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2348_
timestamp 1704896540
transform 1 0 11040 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2349__49
timestamp 1704896540
transform -1 0 10856 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2349_
timestamp 1704896540
transform 1 0 10488 0 1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_2  _2350_
timestamp 1704896540
transform -1 0 10488 0 1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2350__50
timestamp 1704896540
transform 1 0 10120 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2351__51
timestamp 1704896540
transform 1 0 9292 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2351_
timestamp 1704896540
transform 1 0 9568 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_2  _2352_
timestamp 1704896540
transform 1 0 9200 0 1 544
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2352__52
timestamp 1704896540
transform 1 0 9016 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2353__53
timestamp 1704896540
transform -1 0 16468 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _2353_
timestamp 1704896540
transform 1 0 16192 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2354__54
timestamp 1704896540
transform 1 0 15824 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _2354_
timestamp 1704896540
transform 1 0 16100 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _2355_
timestamp 1704896540
transform 1 0 16284 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2355__55
timestamp 1704896540
transform 1 0 15732 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2356__56
timestamp 1704896540
transform -1 0 15916 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _2356_
timestamp 1704896540
transform 1 0 15548 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _2357_
timestamp 1704896540
transform 1 0 14168 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2357__57
timestamp 1704896540
transform -1 0 14444 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2358__58
timestamp 1704896540
transform -1 0 13248 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _2358_
timestamp 1704896540
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2359__59
timestamp 1704896540
transform 1 0 11592 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _2359_
timestamp 1704896540
transform -1 0 12328 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _2360_
timestamp 1704896540
transform -1 0 10856 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2360__60
timestamp 1704896540
transform 1 0 10580 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2361_
timestamp 1704896540
transform 1 0 24564 0 1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2361__15
timestamp 1704896540
transform -1 0 25576 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2362__16
timestamp 1704896540
transform -1 0 25300 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2362_
timestamp 1704896540
transform 1 0 24840 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2363__17
timestamp 1704896540
transform -1 0 24104 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2363_
timestamp 1704896540
transform 1 0 23828 0 1 544
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_2  _2364_
timestamp 1704896540
transform 1 0 23276 0 -1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2364__18
timestamp 1704896540
transform -1 0 23644 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2365__19
timestamp 1704896540
transform 1 0 23000 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2365_
timestamp 1704896540
transform 1 0 23644 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2366__20
timestamp 1704896540
transform -1 0 23000 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2366_
timestamp 1704896540
transform 1 0 22356 0 1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_2  _2367_
timestamp 1704896540
transform 1 0 22448 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2367__21
timestamp 1704896540
transform -1 0 22724 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2368__22
timestamp 1704896540
transform -1 0 22172 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2368_
timestamp 1704896540
transform 1 0 21252 0 1 544
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2369__23
timestamp 1704896540
transform -1 0 21896 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2369_
timestamp 1704896540
transform 1 0 21252 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_2  _2370_
timestamp 1704896540
transform 1 0 20148 0 1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2370__24
timestamp 1704896540
transform -1 0 21620 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2371__25
timestamp 1704896540
transform 1 0 20884 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2371_
timestamp 1704896540
transform -1 0 21068 0 1 544
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_2  _2372_
timestamp 1704896540
transform 1 0 18952 0 1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2372__26
timestamp 1704896540
transform 1 0 18676 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2373_
timestamp 1704896540
transform 1 0 19688 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2373__27
timestamp 1704896540
transform 1 0 18308 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2374_
timestamp 1704896540
transform 1 0 18676 0 1 544
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2374__28
timestamp 1704896540
transform 1 0 18032 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_2  _2375_
timestamp 1704896540
transform -1 0 19688 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2375__29
timestamp 1704896540
transform 1 0 17664 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2376_
timestamp 1704896540
transform 1 0 11408 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2377_
timestamp 1704896540
transform 1 0 11408 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2378_
timestamp 1704896540
transform 1 0 10120 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2379_
timestamp 1704896540
transform 1 0 11592 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2380_
timestamp 1704896540
transform 1 0 10948 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2381_
timestamp 1704896540
transform 1 0 10948 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2382_
timestamp 1704896540
transform 1 0 12788 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2383_
timestamp 1704896540
transform 1 0 12788 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__dlxtn_1  _2384_
timestamp 1704896540
transform 1 0 23920 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2384__30
timestamp 1704896540
transform -1 0 24472 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2385__31
timestamp 1704896540
transform -1 0 24380 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _2385_
timestamp 1704896540
transform 1 0 23920 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2386__32
timestamp 1704896540
transform -1 0 24840 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _2386_
timestamp 1704896540
transform 1 0 24012 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _2387_
timestamp 1704896540
transform 1 0 23460 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2387__33
timestamp 1704896540
transform -1 0 24104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2388__34
timestamp 1704896540
transform -1 0 22816 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _2388_
timestamp 1704896540
transform 1 0 22540 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2389__35
timestamp 1704896540
transform -1 0 21896 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _2389_
timestamp 1704896540
transform 1 0 21620 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2390__36
timestamp 1704896540
transform 1 0 20792 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _2390_
timestamp 1704896540
transform 1 0 21436 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2391__37
timestamp 1704896540
transform 1 0 19780 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _2391_
timestamp 1704896540
transform 1 0 20332 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _2392_
timestamp 1704896540
transform 1 0 4508 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2393_
timestamp 1704896540
transform -1 0 10028 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2394_
timestamp 1704896540
transform -1 0 10580 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2395_
timestamp 1704896540
transform -1 0 9384 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2396_
timestamp 1704896540
transform 1 0 5244 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2397_
timestamp 1704896540
transform 1 0 3220 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2398_
timestamp 1704896540
transform -1 0 5704 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2399_
timestamp 1704896540
transform 1 0 828 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2400_
timestamp 1704896540
transform -1 0 2300 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2401_
timestamp 1704896540
transform 1 0 1932 0 -1 29920
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2402_
timestamp 1704896540
transform 1 0 16836 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2403_
timestamp 1704896540
transform -1 0 19688 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2404_
timestamp 1704896540
transform -1 0 20332 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2405_
timestamp 1704896540
transform -1 0 19044 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2406_
timestamp 1704896540
transform 1 0 12972 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2407_
timestamp 1704896540
transform -1 0 17572 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2408_
timestamp 1704896540
transform -1 0 12512 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2409_
timestamp 1704896540
transform -1 0 10580 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2410_
timestamp 1704896540
transform 1 0 1564 0 1 29920
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 16192 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1704896540
transform -1 0 10212 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1704896540
transform 1 0 18676 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_0_clk
timestamp 1704896540
transform 1 0 4048 0 1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_1_clk
timestamp 1704896540
transform 1 0 9016 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_2_clk
timestamp 1704896540
transform 1 0 11132 0 1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_3_clk
timestamp 1704896540
transform 1 0 5888 0 1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_4_clk
timestamp 1704896540
transform -1 0 3588 0 -1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_5_clk
timestamp 1704896540
transform 1 0 3220 0 1 27744
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_6_clk
timestamp 1704896540
transform -1 0 11132 0 1 28832
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_7_clk
timestamp 1704896540
transform 1 0 11592 0 1 26656
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_8_clk
timestamp 1704896540
transform -1 0 12604 0 1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_9_clk
timestamp 1704896540
transform -1 0 17940 0 -1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_10_clk
timestamp 1704896540
transform -1 0 21620 0 1 27744
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_11_clk
timestamp 1704896540
transform 1 0 25300 0 1 26656
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_12_clk
timestamp 1704896540
transform 1 0 25300 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_13_clk
timestamp 1704896540
transform 1 0 22908 0 -1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_14_clk
timestamp 1704896540
transform 1 0 18768 0 1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_15_clk
timestamp 1704896540
transform 1 0 19596 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_16_clk
timestamp 1704896540
transform 1 0 25300 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_17_clk
timestamp 1704896540
transform 1 0 24564 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_18_clk
timestamp 1704896540
transform -1 0 20516 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_19_clk
timestamp 1704896540
transform 1 0 12696 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_20_clk
timestamp 1704896540
transform -1 0 11592 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_21_clk
timestamp 1704896540
transform 1 0 3588 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 828 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_17
timestamp 1704896540
transform 1 0 2116 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2484 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 1704896540
transform 1 0 5612 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_57
timestamp 1704896540
transform 1 0 5796 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_88 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8648 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_107 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10396 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_113 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10948 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_119
timestamp 1704896540
transform 1 0 11500 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_124
timestamp 1704896540
transform 1 0 11960 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_144
timestamp 1704896540
transform 1 0 13800 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_160
timestamp 1704896540
transform 1 0 15272 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_166
timestamp 1704896540
transform 1 0 15824 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_169
timestamp 1704896540
transform 1 0 16100 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_183
timestamp 1704896540
transform 1 0 17388 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_189
timestamp 1704896540
transform 1 0 17940 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_223
timestamp 1704896540
transform 1 0 21068 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_247
timestamp 1704896540
transform 1 0 23276 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_251
timestamp 1704896540
transform 1 0 23644 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_272 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 25576 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_281
timestamp 1704896540
transform 1 0 26404 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_3
timestamp 1704896540
transform 1 0 828 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_60
timestamp 1704896540
transform 1 0 6072 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_94
timestamp 1704896540
transform 1 0 9200 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1704896540
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_113
timestamp 1704896540
transform 1 0 10948 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_166
timestamp 1704896540
transform 1 0 15824 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_277
timestamp 1704896540
transform 1 0 26036 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_281
timestamp 1704896540
transform 1 0 26404 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_3
timestamp 1704896540
transform 1 0 828 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_7
timestamp 1704896540
transform 1 0 1196 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1704896540
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1704896540
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_85
timestamp 1704896540
transform 1 0 8372 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_91
timestamp 1704896540
transform 1 0 8924 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_141
timestamp 1704896540
transform 1 0 13524 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_147
timestamp 1704896540
transform 1 0 14076 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_151
timestamp 1704896540
transform 1 0 14444 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_178
timestamp 1704896540
transform 1 0 16928 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_187
timestamp 1704896540
transform 1 0 17756 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1704896540
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_235
timestamp 1704896540
transform 1 0 22172 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_250
timestamp 1704896540
transform 1 0 23552 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_256
timestamp 1704896540
transform 1 0 24104 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_260
timestamp 1704896540
transform 1 0 24472 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_274 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 25760 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_286
timestamp 1704896540
transform 1 0 26864 0 1 1632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1704896540
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_15
timestamp 1704896540
transform 1 0 1932 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_24
timestamp 1704896540
transform 1 0 2760 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_30
timestamp 1704896540
transform 1 0 3312 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_34
timestamp 1704896540
transform 1 0 3680 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_47
timestamp 1704896540
transform 1 0 4876 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_51
timestamp 1704896540
transform 1 0 5244 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1704896540
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_65
timestamp 1704896540
transform 1 0 6532 0 -1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_73
timestamp 1704896540
transform 1 0 7268 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_85
timestamp 1704896540
transform 1 0 8372 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_96
timestamp 1704896540
transform 1 0 9384 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_107
timestamp 1704896540
transform 1 0 10396 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1704896540
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_113
timestamp 1704896540
transform 1 0 10948 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_127
timestamp 1704896540
transform 1 0 12236 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_136
timestamp 1704896540
transform 1 0 13064 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_145
timestamp 1704896540
transform 1 0 13892 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_155
timestamp 1704896540
transform 1 0 14812 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1704896540
transform 1 0 15364 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1704896540
transform 1 0 15916 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_169
timestamp 1704896540
transform 1 0 16100 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_173
timestamp 1704896540
transform 1 0 16468 0 -1 2720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_198
timestamp 1704896540
transform 1 0 18768 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_210
timestamp 1704896540
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1704896540
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_228
timestamp 1704896540
transform 1 0 21528 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_240
timestamp 1704896540
transform 1 0 22632 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_276
timestamp 1704896540
transform 1 0 25944 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_281
timestamp 1704896540
transform 1 0 26404 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_3
timestamp 1704896540
transform 1 0 828 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_11
timestamp 1704896540
transform 1 0 1564 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_21
timestamp 1704896540
transform 1 0 2484 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_26
timestamp 1704896540
transform 1 0 2944 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_29
timestamp 1704896540
transform 1 0 3220 0 1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_36
timestamp 1704896540
transform 1 0 3864 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_48
timestamp 1704896540
transform 1 0 4968 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_54
timestamp 1704896540
transform 1 0 5520 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_60
timestamp 1704896540
transform 1 0 6072 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_70
timestamp 1704896540
transform 1 0 6992 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_85
timestamp 1704896540
transform 1 0 8372 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_103
timestamp 1704896540
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_117
timestamp 1704896540
transform 1 0 11316 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_124
timestamp 1704896540
transform 1 0 11960 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_136
timestamp 1704896540
transform 1 0 13064 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_141
timestamp 1704896540
transform 1 0 13524 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_155
timestamp 1704896540
transform 1 0 14812 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_165
timestamp 1704896540
transform 1 0 15732 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_182
timestamp 1704896540
transform 1 0 17296 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_194
timestamp 1704896540
transform 1 0 18400 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_197
timestamp 1704896540
transform 1 0 18676 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_213
timestamp 1704896540
transform 1 0 20148 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_218
timestamp 1704896540
transform 1 0 20608 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_224
timestamp 1704896540
transform 1 0 21160 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_232
timestamp 1704896540
transform 1 0 21896 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_242
timestamp 1704896540
transform 1 0 22816 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1704896540
transform 1 0 23644 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_253
timestamp 1704896540
transform 1 0 23828 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_282
timestamp 1704896540
transform 1 0 26496 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_288
timestamp 1704896540
transform 1 0 27048 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1704896540
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_15
timestamp 1704896540
transform 1 0 1932 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_23
timestamp 1704896540
transform 1 0 2668 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_29
timestamp 1704896540
transform 1 0 3220 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_35
timestamp 1704896540
transform 1 0 3772 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_44
timestamp 1704896540
transform 1 0 4600 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_57
timestamp 1704896540
transform 1 0 5796 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_74
timestamp 1704896540
transform 1 0 7360 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_78
timestamp 1704896540
transform 1 0 7728 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_86
timestamp 1704896540
transform 1 0 8464 0 -1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_96
timestamp 1704896540
transform 1 0 9384 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_108
timestamp 1704896540
transform 1 0 10488 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_113
timestamp 1704896540
transform 1 0 10948 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_132
timestamp 1704896540
transform 1 0 12696 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_140
timestamp 1704896540
transform 1 0 13432 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_147
timestamp 1704896540
transform 1 0 14076 0 -1 3808
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_174
timestamp 1704896540
transform 1 0 16560 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_186
timestamp 1704896540
transform 1 0 17664 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_191
timestamp 1704896540
transform 1 0 18124 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_203
timestamp 1704896540
transform 1 0 19228 0 -1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_209
timestamp 1704896540
transform 1 0 19780 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_221
timestamp 1704896540
transform 1 0 20884 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_225
timestamp 1704896540
transform 1 0 21252 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_232
timestamp 1704896540
transform 1 0 21896 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_239
timestamp 1704896540
transform 1 0 22540 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_250
timestamp 1704896540
transform 1 0 23552 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_260
timestamp 1704896540
transform 1 0 24472 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_268
timestamp 1704896540
transform 1 0 25208 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1704896540
transform 1 0 25668 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1704896540
transform 1 0 26220 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_281
timestamp 1704896540
transform 1 0 26404 0 -1 3808
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1704896540
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_15
timestamp 1704896540
transform 1 0 1932 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_19
timestamp 1704896540
transform 1 0 2300 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_25
timestamp 1704896540
transform 1 0 2852 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_45
timestamp 1704896540
transform 1 0 4692 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_58
timestamp 1704896540
transform 1 0 5888 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_66
timestamp 1704896540
transform 1 0 6624 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_82
timestamp 1704896540
transform 1 0 8096 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_85
timestamp 1704896540
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_92
timestamp 1704896540
transform 1 0 9016 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_112
timestamp 1704896540
transform 1 0 10856 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_120
timestamp 1704896540
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_124
timestamp 1704896540
transform 1 0 11960 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_132
timestamp 1704896540
transform 1 0 12696 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1704896540
transform 1 0 13340 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_144
timestamp 1704896540
transform 1 0 13800 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_148
timestamp 1704896540
transform 1 0 14168 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_181
timestamp 1704896540
transform 1 0 17204 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1704896540
transform 1 0 18492 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_205
timestamp 1704896540
transform 1 0 19412 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_211
timestamp 1704896540
transform 1 0 19964 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_237
timestamp 1704896540
transform 1 0 22356 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_250
timestamp 1704896540
transform 1 0 23552 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_253
timestamp 1704896540
transform 1 0 23828 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_271
timestamp 1704896540
transform 1 0 25484 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_3
timestamp 1704896540
transform 1 0 828 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_19
timestamp 1704896540
transform 1 0 2300 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_23
timestamp 1704896540
transform 1 0 2668 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_35
timestamp 1704896540
transform 1 0 3772 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_53
timestamp 1704896540
transform 1 0 5428 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_62
timestamp 1704896540
transform 1 0 6256 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_70
timestamp 1704896540
transform 1 0 6992 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_74
timestamp 1704896540
transform 1 0 7360 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_99
timestamp 1704896540
transform 1 0 9660 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_118
timestamp 1704896540
transform 1 0 11408 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_130
timestamp 1704896540
transform 1 0 12512 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_146
timestamp 1704896540
transform 1 0 13984 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_151
timestamp 1704896540
transform 1 0 14444 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_159
timestamp 1704896540
transform 1 0 15180 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_169
timestamp 1704896540
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_183
timestamp 1704896540
transform 1 0 17388 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_208
timestamp 1704896540
transform 1 0 19688 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_213
timestamp 1704896540
transform 1 0 20148 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_221
timestamp 1704896540
transform 1 0 20884 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_230
timestamp 1704896540
transform 1 0 21712 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_239
timestamp 1704896540
transform 1 0 22540 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_243
timestamp 1704896540
transform 1 0 22908 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_250
timestamp 1704896540
transform 1 0 23552 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1704896540
transform 1 0 26220 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_3
timestamp 1704896540
transform 1 0 828 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_19
timestamp 1704896540
transform 1 0 2300 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_26
timestamp 1704896540
transform 1 0 2944 0 1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1704896540
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_41
timestamp 1704896540
transform 1 0 4324 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_50
timestamp 1704896540
transform 1 0 5152 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_59
timestamp 1704896540
transform 1 0 5980 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_78
timestamp 1704896540
transform 1 0 7728 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_85
timestamp 1704896540
transform 1 0 8372 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_90
timestamp 1704896540
transform 1 0 8832 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_102
timestamp 1704896540
transform 1 0 9936 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_112
timestamp 1704896540
transform 1 0 10856 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_128
timestamp 1704896540
transform 1 0 12328 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_133
timestamp 1704896540
transform 1 0 12788 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_138
timestamp 1704896540
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_141
timestamp 1704896540
transform 1 0 13524 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_147
timestamp 1704896540
transform 1 0 14076 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_175
timestamp 1704896540
transform 1 0 16652 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_187
timestamp 1704896540
transform 1 0 17756 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1704896540
transform 1 0 18492 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_197
timestamp 1704896540
transform 1 0 18676 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_205
timestamp 1704896540
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_223
timestamp 1704896540
transform 1 0 21068 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_238
timestamp 1704896540
transform 1 0 22448 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_246
timestamp 1704896540
transform 1 0 23184 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_253
timestamp 1704896540
transform 1 0 23828 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_259
timestamp 1704896540
transform 1 0 24380 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_286
timestamp 1704896540
transform 1 0 26864 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_3
timestamp 1704896540
transform 1 0 828 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_7
timestamp 1704896540
transform 1 0 1196 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_11
timestamp 1704896540
transform 1 0 1564 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_35
timestamp 1704896540
transform 1 0 3772 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1704896540
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_72
timestamp 1704896540
transform 1 0 7176 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_84
timestamp 1704896540
transform 1 0 8280 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_92
timestamp 1704896540
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_109
timestamp 1704896540
transform 1 0 10580 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_123
timestamp 1704896540
transform 1 0 11868 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_133
timestamp 1704896540
transform 1 0 12788 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_147
timestamp 1704896540
transform 1 0 14076 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_151
timestamp 1704896540
transform 1 0 14444 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_155
timestamp 1704896540
transform 1 0 14812 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_159
timestamp 1704896540
transform 1 0 15180 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_163
timestamp 1704896540
transform 1 0 15548 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1704896540
transform 1 0 15916 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_169
timestamp 1704896540
transform 1 0 16100 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_173
timestamp 1704896540
transform 1 0 16468 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_177
timestamp 1704896540
transform 1 0 16836 0 -1 5984
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_197
timestamp 1704896540
transform 1 0 18676 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_209
timestamp 1704896540
transform 1 0 19780 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_217
timestamp 1704896540
transform 1 0 20516 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1704896540
transform 1 0 21068 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1704896540
transform 1 0 21252 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_237
timestamp 1704896540
transform 1 0 22356 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_245
timestamp 1704896540
transform 1 0 23092 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_264
timestamp 1704896540
transform 1 0 24840 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_276
timestamp 1704896540
transform 1 0 25944 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_281
timestamp 1704896540
transform 1 0 26404 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_3
timestamp 1704896540
transform 1 0 828 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_21
timestamp 1704896540
transform 1 0 2484 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_26
timestamp 1704896540
transform 1 0 2944 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_29
timestamp 1704896540
transform 1 0 3220 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_38
timestamp 1704896540
transform 1 0 4048 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_47
timestamp 1704896540
transform 1 0 4876 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_58
timestamp 1704896540
transform 1 0 5888 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_64
timestamp 1704896540
transform 1 0 6440 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_68
timestamp 1704896540
transform 1 0 6808 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_92
timestamp 1704896540
transform 1 0 9016 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_129
timestamp 1704896540
transform 1 0 12420 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_137
timestamp 1704896540
transform 1 0 13156 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_145
timestamp 1704896540
transform 1 0 13892 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_167
timestamp 1704896540
transform 1 0 15916 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_187
timestamp 1704896540
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_197
timestamp 1704896540
transform 1 0 18676 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1704896540
transform 1 0 23644 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_256
timestamp 1704896540
transform 1 0 24104 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_273
timestamp 1704896540
transform 1 0 25668 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_288
timestamp 1704896540
transform 1 0 27048 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_25
timestamp 1704896540
transform 1 0 2852 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_57
timestamp 1704896540
transform 1 0 5796 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_76
timestamp 1704896540
transform 1 0 7544 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_96
timestamp 1704896540
transform 1 0 9384 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_108
timestamp 1704896540
transform 1 0 10488 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_113
timestamp 1704896540
transform 1 0 10948 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_130
timestamp 1704896540
transform 1 0 12512 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_162
timestamp 1704896540
transform 1 0 15456 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_169
timestamp 1704896540
transform 1 0 16100 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_173
timestamp 1704896540
transform 1 0 16468 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_177
timestamp 1704896540
transform 1 0 16836 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_195
timestamp 1704896540
transform 1 0 18492 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_207
timestamp 1704896540
transform 1 0 19596 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_212
timestamp 1704896540
transform 1 0 20056 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_228
timestamp 1704896540
transform 1 0 21528 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_241
timestamp 1704896540
transform 1 0 22724 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_253
timestamp 1704896540
transform 1 0 23828 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_262
timestamp 1704896540
transform 1 0 24656 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_270
timestamp 1704896540
transform 1 0 25392 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_277
timestamp 1704896540
transform 1 0 26036 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_281
timestamp 1704896540
transform 1 0 26404 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_3
timestamp 1704896540
transform 1 0 828 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_22
timestamp 1704896540
transform 1 0 2576 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_36
timestamp 1704896540
transform 1 0 3864 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_45
timestamp 1704896540
transform 1 0 4692 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_54
timestamp 1704896540
transform 1 0 5520 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_62
timestamp 1704896540
transform 1 0 6256 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_72
timestamp 1704896540
transform 1 0 7176 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_85
timestamp 1704896540
transform 1 0 8372 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_91
timestamp 1704896540
transform 1 0 8924 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_99
timestamp 1704896540
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_109
timestamp 1704896540
transform 1 0 10580 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_113
timestamp 1704896540
transform 1 0 10948 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_136
timestamp 1704896540
transform 1 0 13064 0 1 7072
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1704896540
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1704896540
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_165
timestamp 1704896540
transform 1 0 15732 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_172
timestamp 1704896540
transform 1 0 16376 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_180
timestamp 1704896540
transform 1 0 17112 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_186
timestamp 1704896540
transform 1 0 17664 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_194
timestamp 1704896540
transform 1 0 18400 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_197
timestamp 1704896540
transform 1 0 18676 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_210
timestamp 1704896540
transform 1 0 19872 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_222
timestamp 1704896540
transform 1 0 20976 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_228
timestamp 1704896540
transform 1 0 21528 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_232
timestamp 1704896540
transform 1 0 21896 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_253
timestamp 1704896540
transform 1 0 23828 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_261
timestamp 1704896540
transform 1 0 24564 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_274
timestamp 1704896540
transform 1 0 25760 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_286
timestamp 1704896540
transform 1 0 26864 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1704896540
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_15
timestamp 1704896540
transform 1 0 1932 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_34
timestamp 1704896540
transform 1 0 3680 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1704896540
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_57
timestamp 1704896540
transform 1 0 5796 0 -1 8160
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_71
timestamp 1704896540
transform 1 0 7084 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_83
timestamp 1704896540
transform 1 0 8188 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_95
timestamp 1704896540
transform 1 0 9292 0 -1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_100
timestamp 1704896540
transform 1 0 9752 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_113
timestamp 1704896540
transform 1 0 10948 0 -1 8160
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_132
timestamp 1704896540
transform 1 0 12696 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_144
timestamp 1704896540
transform 1 0 13800 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1704896540
transform 1 0 15916 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_237
timestamp 1704896540
transform 1 0 22356 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_247
timestamp 1704896540
transform 1 0 23276 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_254
timestamp 1704896540
transform 1 0 23920 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_284
timestamp 1704896540
transform 1 0 26680 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_288
timestamp 1704896540
transform 1 0 27048 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1704896540
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_45
timestamp 1704896540
transform 1 0 4692 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_85
timestamp 1704896540
transform 1 0 8372 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_93
timestamp 1704896540
transform 1 0 9108 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_123
timestamp 1704896540
transform 1 0 11868 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1704896540
transform 1 0 13340 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_141
timestamp 1704896540
transform 1 0 13524 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_163
timestamp 1704896540
transform 1 0 15548 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_169
timestamp 1704896540
transform 1 0 16100 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_173
timestamp 1704896540
transform 1 0 16468 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_181
timestamp 1704896540
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_186
timestamp 1704896540
transform 1 0 17664 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_192
timestamp 1704896540
transform 1 0 18216 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_217
timestamp 1704896540
transform 1 0 20516 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_224
timestamp 1704896540
transform 1 0 21160 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_236
timestamp 1704896540
transform 1 0 22264 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_242
timestamp 1704896540
transform 1 0 22816 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_247
timestamp 1704896540
transform 1 0 23276 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_260
timestamp 1704896540
transform 1 0 24472 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_269
timestamp 1704896540
transform 1 0 25300 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_275
timestamp 1704896540
transform 1 0 25852 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_287
timestamp 1704896540
transform 1 0 26956 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_3
timestamp 1704896540
transform 1 0 828 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_29
timestamp 1704896540
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_52
timestamp 1704896540
transform 1 0 5336 0 -1 9248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1704896540
transform 1 0 5796 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_69
timestamp 1704896540
transform 1 0 6900 0 -1 9248
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_99
timestamp 1704896540
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1704896540
transform 1 0 10764 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_151
timestamp 1704896540
transform 1 0 14444 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_159
timestamp 1704896540
transform 1 0 15180 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1704896540
transform 1 0 15916 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_169
timestamp 1704896540
transform 1 0 16100 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_175
timestamp 1704896540
transform 1 0 16652 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_179
timestamp 1704896540
transform 1 0 17020 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_215
timestamp 1704896540
transform 1 0 20332 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 1704896540
transform 1 0 21068 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_225
timestamp 1704896540
transform 1 0 21252 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_237
timestamp 1704896540
transform 1 0 22356 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_253
timestamp 1704896540
transform 1 0 23828 0 -1 9248
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_264
timestamp 1704896540
transform 1 0 24840 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_276
timestamp 1704896540
transform 1 0 25944 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_281
timestamp 1704896540
transform 1 0 26404 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_19
timestamp 1704896540
transform 1 0 2300 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_29
timestamp 1704896540
transform 1 0 3220 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_75
timestamp 1704896540
transform 1 0 7452 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_85
timestamp 1704896540
transform 1 0 8372 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_107
timestamp 1704896540
transform 1 0 10396 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_124
timestamp 1704896540
transform 1 0 11960 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_128
timestamp 1704896540
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_132
timestamp 1704896540
transform 1 0 12696 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_136
timestamp 1704896540
transform 1 0 13064 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_141
timestamp 1704896540
transform 1 0 13524 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_152
timestamp 1704896540
transform 1 0 14536 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_165
timestamp 1704896540
transform 1 0 15732 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_182
timestamp 1704896540
transform 1 0 17296 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_186
timestamp 1704896540
transform 1 0 17664 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_193
timestamp 1704896540
transform 1 0 18308 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_197
timestamp 1704896540
transform 1 0 18676 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_216
timestamp 1704896540
transform 1 0 20424 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_224
timestamp 1704896540
transform 1 0 21160 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_231
timestamp 1704896540
transform 1 0 21804 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_246
timestamp 1704896540
transform 1 0 23184 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_260
timestamp 1704896540
transform 1 0 24472 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_277
timestamp 1704896540
transform 1 0 26036 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_3
timestamp 1704896540
transform 1 0 828 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_15
timestamp 1704896540
transform 1 0 1932 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_53
timestamp 1704896540
transform 1 0 5428 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_63
timestamp 1704896540
transform 1 0 6348 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_94
timestamp 1704896540
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_126
timestamp 1704896540
transform 1 0 12144 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_130
timestamp 1704896540
transform 1 0 12512 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_142
timestamp 1704896540
transform 1 0 13616 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 1704896540
transform 1 0 15916 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_178
timestamp 1704896540
transform 1 0 16928 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_182
timestamp 1704896540
transform 1 0 17296 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_200
timestamp 1704896540
transform 1 0 18952 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_213
timestamp 1704896540
transform 1 0 20148 0 -1 10336
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_241
timestamp 1704896540
transform 1 0 22724 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_253
timestamp 1704896540
transform 1 0 23828 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_261
timestamp 1704896540
transform 1 0 24564 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_265
timestamp 1704896540
transform 1 0 24932 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_277
timestamp 1704896540
transform 1 0 26036 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_281
timestamp 1704896540
transform 1 0 26404 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_3
timestamp 1704896540
transform 1 0 828 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_18
timestamp 1704896540
transform 1 0 2208 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_29
timestamp 1704896540
transform 1 0 3220 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_85
timestamp 1704896540
transform 1 0 8372 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_93
timestamp 1704896540
transform 1 0 9108 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_114
timestamp 1704896540
transform 1 0 11040 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_122
timestamp 1704896540
transform 1 0 11776 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_131
timestamp 1704896540
transform 1 0 12604 0 1 10336
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1704896540
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_153
timestamp 1704896540
transform 1 0 14628 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_157
timestamp 1704896540
transform 1 0 14996 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_164
timestamp 1704896540
transform 1 0 15640 0 1 10336
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_171
timestamp 1704896540
transform 1 0 16284 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_183
timestamp 1704896540
transform 1 0 17388 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 1704896540
transform 1 0 18492 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_203
timestamp 1704896540
transform 1 0 19228 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_211
timestamp 1704896540
transform 1 0 19964 0 1 10336
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_237
timestamp 1704896540
transform 1 0 22356 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_249
timestamp 1704896540
transform 1 0 23460 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_253
timestamp 1704896540
transform 1 0 23828 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_261
timestamp 1704896540
transform 1 0 24564 0 1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_267
timestamp 1704896540
transform 1 0 25116 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_279
timestamp 1704896540
transform 1 0 26220 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_287
timestamp 1704896540
transform 1 0 26956 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_52
timestamp 1704896540
transform 1 0 5336 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_57
timestamp 1704896540
transform 1 0 5796 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_77
timestamp 1704896540
transform 1 0 7636 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_106
timestamp 1704896540
transform 1 0 10304 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_113
timestamp 1704896540
transform 1 0 10948 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_121
timestamp 1704896540
transform 1 0 11684 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_145
timestamp 1704896540
transform 1 0 13892 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_158
timestamp 1704896540
transform 1 0 15088 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_166
timestamp 1704896540
transform 1 0 15824 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_169
timestamp 1704896540
transform 1 0 16100 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_197
timestamp 1704896540
transform 1 0 18676 0 -1 11424
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_210
timestamp 1704896540
transform 1 0 19872 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_222
timestamp 1704896540
transform 1 0 20976 0 -1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_225
timestamp 1704896540
transform 1 0 21252 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_237
timestamp 1704896540
transform 1 0 22356 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_244
timestamp 1704896540
transform 1 0 23000 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_278
timestamp 1704896540
transform 1 0 26128 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_281
timestamp 1704896540
transform 1 0 26404 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_3
timestamp 1704896540
transform 1 0 828 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_26
timestamp 1704896540
transform 1 0 2944 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_29
timestamp 1704896540
transform 1 0 3220 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_101
timestamp 1704896540
transform 1 0 9844 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1704896540
transform 1 0 13340 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_141
timestamp 1704896540
transform 1 0 13524 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_168
timestamp 1704896540
transform 1 0 16008 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_176
timestamp 1704896540
transform 1 0 16744 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_188
timestamp 1704896540
transform 1 0 17848 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_192
timestamp 1704896540
transform 1 0 18216 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_219
timestamp 1704896540
transform 1 0 20700 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_239
timestamp 1704896540
transform 1 0 22540 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_3
timestamp 1704896540
transform 1 0 828 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_57
timestamp 1704896540
transform 1 0 5796 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_80
timestamp 1704896540
transform 1 0 7912 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_91
timestamp 1704896540
transform 1 0 8924 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_99
timestamp 1704896540
transform 1 0 9660 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_113
timestamp 1704896540
transform 1 0 10948 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_130
timestamp 1704896540
transform 1 0 12512 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_155
timestamp 1704896540
transform 1 0 14812 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_159
timestamp 1704896540
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_185
timestamp 1704896540
transform 1 0 17572 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_220
timestamp 1704896540
transform 1 0 20792 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_263
timestamp 1704896540
transform 1 0 24748 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_284
timestamp 1704896540
transform 1 0 26680 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_288
timestamp 1704896540
transform 1 0 27048 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_3
timestamp 1704896540
transform 1 0 828 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_53
timestamp 1704896540
transform 1 0 5428 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_82
timestamp 1704896540
transform 1 0 8096 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_85
timestamp 1704896540
transform 1 0 8372 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_93
timestamp 1704896540
transform 1 0 9108 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_106
timestamp 1704896540
transform 1 0 10304 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_118
timestamp 1704896540
transform 1 0 11408 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_127
timestamp 1704896540
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_136
timestamp 1704896540
transform 1 0 13064 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_150
timestamp 1704896540
transform 1 0 14352 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_161
timestamp 1704896540
transform 1 0 15364 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_165
timestamp 1704896540
transform 1 0 15732 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_175
timestamp 1704896540
transform 1 0 16652 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_187
timestamp 1704896540
transform 1 0 17756 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_220
timestamp 1704896540
transform 1 0 20792 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_228
timestamp 1704896540
transform 1 0 21528 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 1704896540
transform 1 0 23644 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_287
timestamp 1704896540
transform 1 0 26956 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_53
timestamp 1704896540
transform 1 0 5428 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_57
timestamp 1704896540
transform 1 0 5796 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_89
timestamp 1704896540
transform 1 0 8740 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_95
timestamp 1704896540
transform 1 0 9292 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_163
timestamp 1704896540
transform 1 0 15548 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1704896540
transform 1 0 15916 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_178
timestamp 1704896540
transform 1 0 16928 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_195
timestamp 1704896540
transform 1 0 18492 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_214
timestamp 1704896540
transform 1 0 20240 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1704896540
transform 1 0 21068 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_263
timestamp 1704896540
transform 1 0 24748 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_281
timestamp 1704896540
transform 1 0 26404 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_3
timestamp 1704896540
transform 1 0 828 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_26
timestamp 1704896540
transform 1 0 2944 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_45
timestamp 1704896540
transform 1 0 4692 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_75
timestamp 1704896540
transform 1 0 7452 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1704896540
transform 1 0 8188 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_85
timestamp 1704896540
transform 1 0 8372 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_91
timestamp 1704896540
transform 1 0 8924 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_112
timestamp 1704896540
transform 1 0 10856 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_137
timestamp 1704896540
transform 1 0 13156 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_146
timestamp 1704896540
transform 1 0 13984 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_158
timestamp 1704896540
transform 1 0 15088 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_193
timestamp 1704896540
transform 1 0 18308 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_197
timestamp 1704896540
transform 1 0 18676 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_205
timestamp 1704896540
transform 1 0 19412 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 1704896540
transform 1 0 23644 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_271
timestamp 1704896540
transform 1 0 25484 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_288
timestamp 1704896540
transform 1 0 27048 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_19
timestamp 1704896540
transform 1 0 2300 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_46
timestamp 1704896540
transform 1 0 4784 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_57
timestamp 1704896540
transform 1 0 5796 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_66
timestamp 1704896540
transform 1 0 6624 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_83
timestamp 1704896540
transform 1 0 8188 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_95
timestamp 1704896540
transform 1 0 9292 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_110
timestamp 1704896540
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_121
timestamp 1704896540
transform 1 0 11684 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_132
timestamp 1704896540
transform 1 0 12696 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_140
timestamp 1704896540
transform 1 0 13432 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 1704896540
transform 1 0 15364 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1704896540
transform 1 0 15916 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_169
timestamp 1704896540
transform 1 0 16100 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_178
timestamp 1704896540
transform 1 0 16928 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_200
timestamp 1704896540
transform 1 0 18952 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_221
timestamp 1704896540
transform 1 0 20884 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_249
timestamp 1704896540
transform 1 0 23460 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_257
timestamp 1704896540
transform 1 0 24196 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_284
timestamp 1704896540
transform 1 0 26680 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_288
timestamp 1704896540
transform 1 0 27048 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_3
timestamp 1704896540
transform 1 0 828 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_37
timestamp 1704896540
transform 1 0 3956 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_85
timestamp 1704896540
transform 1 0 8372 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_116
timestamp 1704896540
transform 1 0 11224 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_120
timestamp 1704896540
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_128
timestamp 1704896540
transform 1 0 12328 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_147
timestamp 1704896540
transform 1 0 14076 0 1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_170
timestamp 1704896540
transform 1 0 16192 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_182
timestamp 1704896540
transform 1 0 17296 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_194
timestamp 1704896540
transform 1 0 18400 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_197
timestamp 1704896540
transform 1 0 18676 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_223
timestamp 1704896540
transform 1 0 21068 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_232
timestamp 1704896540
transform 1 0 21896 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_250
timestamp 1704896540
transform 1 0 23552 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_288
timestamp 1704896540
transform 1 0 27048 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_3
timestamp 1704896540
transform 1 0 828 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_12
timestamp 1704896540
transform 1 0 1656 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_77
timestamp 1704896540
transform 1 0 7636 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1704896540
transform 1 0 10764 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_154
timestamp 1704896540
transform 1 0 14720 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_164
timestamp 1704896540
transform 1 0 15640 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_217
timestamp 1704896540
transform 1 0 20516 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_233
timestamp 1704896540
transform 1 0 21988 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_256
timestamp 1704896540
transform 1 0 24104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_264
timestamp 1704896540
transform 1 0 24840 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_273
timestamp 1704896540
transform 1 0 25668 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 1704896540
transform 1 0 26220 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_281
timestamp 1704896540
transform 1 0 26404 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_3
timestamp 1704896540
transform 1 0 828 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_11
timestamp 1704896540
transform 1 0 1564 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1704896540
transform 1 0 3036 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_34
timestamp 1704896540
transform 1 0 3680 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_42
timestamp 1704896540
transform 1 0 4416 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1704896540
transform 1 0 8188 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_105
timestamp 1704896540
transform 1 0 10212 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_121
timestamp 1704896540
transform 1 0 11684 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_130
timestamp 1704896540
transform 1 0 12512 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_138
timestamp 1704896540
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_141
timestamp 1704896540
transform 1 0 13524 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_152
timestamp 1704896540
transform 1 0 14536 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_177
timestamp 1704896540
transform 1 0 16836 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_183
timestamp 1704896540
transform 1 0 17388 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_187
timestamp 1704896540
transform 1 0 17756 0 1 15776
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_224
timestamp 1704896540
transform 1 0 21160 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_236
timestamp 1704896540
transform 1 0 22264 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_248
timestamp 1704896540
transform 1 0 23368 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_253
timestamp 1704896540
transform 1 0 23828 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_259
timestamp 1704896540
transform 1 0 24380 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_267
timestamp 1704896540
transform 1 0 25116 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_286
timestamp 1704896540
transform 1 0 26864 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_3
timestamp 1704896540
transform 1 0 828 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_27
timestamp 1704896540
transform 1 0 3036 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_45
timestamp 1704896540
transform 1 0 4692 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_53
timestamp 1704896540
transform 1 0 5428 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_57
timestamp 1704896540
transform 1 0 5796 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_65
timestamp 1704896540
transform 1 0 6532 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_76
timestamp 1704896540
transform 1 0 7544 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_98
timestamp 1704896540
transform 1 0 9568 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_109
timestamp 1704896540
transform 1 0 10580 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_129
timestamp 1704896540
transform 1 0 12420 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_135
timestamp 1704896540
transform 1 0 12972 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_140
timestamp 1704896540
transform 1 0 13432 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_165
timestamp 1704896540
transform 1 0 15732 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_177
timestamp 1704896540
transform 1 0 16836 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_200
timestamp 1704896540
transform 1 0 18952 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_210
timestamp 1704896540
transform 1 0 19872 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_216
timestamp 1704896540
transform 1 0 20424 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_220
timestamp 1704896540
transform 1 0 20792 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_234
timestamp 1704896540
transform 1 0 22080 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_249
timestamp 1704896540
transform 1 0 23460 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_268
timestamp 1704896540
transform 1 0 25208 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_275
timestamp 1704896540
transform 1 0 25852 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 1704896540
transform 1 0 26220 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_281
timestamp 1704896540
transform 1 0 26404 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_3
timestamp 1704896540
transform 1 0 828 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_15
timestamp 1704896540
transform 1 0 1932 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_21
timestamp 1704896540
transform 1 0 2484 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1704896540
transform 1 0 3036 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_66
timestamp 1704896540
transform 1 0 6624 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_71
timestamp 1704896540
transform 1 0 7084 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_77
timestamp 1704896540
transform 1 0 7636 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_149
timestamp 1704896540
transform 1 0 14260 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_193
timestamp 1704896540
transform 1 0 18308 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_197
timestamp 1704896540
transform 1 0 18676 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_215
timestamp 1704896540
transform 1 0 20332 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_232
timestamp 1704896540
transform 1 0 21896 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_236
timestamp 1704896540
transform 1 0 22264 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_250
timestamp 1704896540
transform 1 0 23552 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_287
timestamp 1704896540
transform 1 0 26956 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_27
timestamp 1704896540
transform 1 0 3036 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_45
timestamp 1704896540
transform 1 0 4692 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_57
timestamp 1704896540
transform 1 0 5796 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_79
timestamp 1704896540
transform 1 0 7820 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_98
timestamp 1704896540
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_108
timestamp 1704896540
transform 1 0 10488 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_113
timestamp 1704896540
transform 1 0 10948 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_154
timestamp 1704896540
transform 1 0 14720 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_169
timestamp 1704896540
transform 1 0 16100 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_188
timestamp 1704896540
transform 1 0 17848 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_192
timestamp 1704896540
transform 1 0 18216 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_198
timestamp 1704896540
transform 1 0 18768 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_204
timestamp 1704896540
transform 1 0 19320 0 -1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_212
timestamp 1704896540
transform 1 0 20056 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_230
timestamp 1704896540
transform 1 0 21712 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_234
timestamp 1704896540
transform 1 0 22080 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_242
timestamp 1704896540
transform 1 0 22816 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_247
timestamp 1704896540
transform 1 0 23276 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_253
timestamp 1704896540
transform 1 0 23828 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_262
timestamp 1704896540
transform 1 0 24656 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_276
timestamp 1704896540
transform 1 0 25944 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_281
timestamp 1704896540
transform 1 0 26404 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_3
timestamp 1704896540
transform 1 0 828 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_15
timestamp 1704896540
transform 1 0 1932 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1704896540
transform 1 0 3036 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_29
timestamp 1704896540
transform 1 0 3220 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_39
timestamp 1704896540
transform 1 0 4140 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_62
timestamp 1704896540
transform 1 0 6256 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_67
timestamp 1704896540
transform 1 0 6716 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_78
timestamp 1704896540
transform 1 0 7728 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_85
timestamp 1704896540
transform 1 0 8372 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_105
timestamp 1704896540
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_135
timestamp 1704896540
transform 1 0 12972 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1704896540
transform 1 0 13340 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_141
timestamp 1704896540
transform 1 0 13524 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_168
timestamp 1704896540
transform 1 0 16008 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_185
timestamp 1704896540
transform 1 0 17572 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_197
timestamp 1704896540
transform 1 0 18676 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_210
timestamp 1704896540
transform 1 0 19872 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_214
timestamp 1704896540
transform 1 0 20240 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_231
timestamp 1704896540
transform 1 0 21804 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_262
timestamp 1704896540
transform 1 0 24656 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_270
timestamp 1704896540
transform 1 0 25392 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_3
timestamp 1704896540
transform 1 0 828 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_11
timestamp 1704896540
transform 1 0 1564 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_36
timestamp 1704896540
transform 1 0 3864 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_57
timestamp 1704896540
transform 1 0 5796 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_77
timestamp 1704896540
transform 1 0 7636 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_109
timestamp 1704896540
transform 1 0 10580 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_113
timestamp 1704896540
transform 1 0 10948 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_133
timestamp 1704896540
transform 1 0 12788 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_141
timestamp 1704896540
transform 1 0 13524 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_157
timestamp 1704896540
transform 1 0 14996 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_165
timestamp 1704896540
transform 1 0 15732 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_178
timestamp 1704896540
transform 1 0 16928 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_198
timestamp 1704896540
transform 1 0 18768 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_225
timestamp 1704896540
transform 1 0 21252 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_231
timestamp 1704896540
transform 1 0 21804 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_240
timestamp 1704896540
transform 1 0 22632 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_276
timestamp 1704896540
transform 1 0 25944 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_281
timestamp 1704896540
transform 1 0 26404 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_19
timestamp 1704896540
transform 1 0 2300 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_25
timestamp 1704896540
transform 1 0 2852 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_29
timestamp 1704896540
transform 1 0 3220 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_78
timestamp 1704896540
transform 1 0 7728 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_97
timestamp 1704896540
transform 1 0 9476 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_113
timestamp 1704896540
transform 1 0 10948 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_136
timestamp 1704896540
transform 1 0 13064 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_146
timestamp 1704896540
transform 1 0 13984 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_197
timestamp 1704896540
transform 1 0 18676 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_227
timestamp 1704896540
transform 1 0 21436 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_233
timestamp 1704896540
transform 1 0 21988 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_240
timestamp 1704896540
transform 1 0 22632 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_259
timestamp 1704896540
transform 1 0 24380 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_286
timestamp 1704896540
transform 1 0 26864 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_3
timestamp 1704896540
transform 1 0 828 0 -1 20128
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_10
timestamp 1704896540
transform 1 0 1472 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_22
timestamp 1704896540
transform 1 0 2576 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_34
timestamp 1704896540
transform 1 0 3680 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_44
timestamp 1704896540
transform 1 0 4600 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_53
timestamp 1704896540
transform 1 0 5428 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_57
timestamp 1704896540
transform 1 0 5796 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_65
timestamp 1704896540
transform 1 0 6532 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_83
timestamp 1704896540
transform 1 0 8188 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_87
timestamp 1704896540
transform 1 0 8556 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_113
timestamp 1704896540
transform 1 0 10948 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_129
timestamp 1704896540
transform 1 0 12420 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_140
timestamp 1704896540
transform 1 0 13432 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_157
timestamp 1704896540
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_172
timestamp 1704896540
transform 1 0 16376 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_197
timestamp 1704896540
transform 1 0 18676 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_218
timestamp 1704896540
transform 1 0 20608 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_234
timestamp 1704896540
transform 1 0 22080 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_238
timestamp 1704896540
transform 1 0 22448 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_242
timestamp 1704896540
transform 1 0 22816 0 -1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_263
timestamp 1704896540
transform 1 0 24748 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_275
timestamp 1704896540
transform 1 0 25852 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_279
timestamp 1704896540
transform 1 0 26220 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_19
timestamp 1704896540
transform 1 0 2300 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_50
timestamp 1704896540
transform 1 0 5152 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_71
timestamp 1704896540
transform 1 0 7084 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_80
timestamp 1704896540
transform 1 0 7912 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_93
timestamp 1704896540
transform 1 0 9108 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_104
timestamp 1704896540
transform 1 0 10120 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_138
timestamp 1704896540
transform 1 0 13248 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_171
timestamp 1704896540
transform 1 0 16284 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_192
timestamp 1704896540
transform 1 0 18216 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_197
timestamp 1704896540
transform 1 0 18676 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_220
timestamp 1704896540
transform 1 0 20792 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_237
timestamp 1704896540
transform 1 0 22356 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_253
timestamp 1704896540
transform 1 0 23828 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_265
timestamp 1704896540
transform 1 0 24932 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_3
timestamp 1704896540
transform 1 0 828 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1704896540
transform 1 0 5612 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_57
timestamp 1704896540
transform 1 0 5796 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_65
timestamp 1704896540
transform 1 0 6532 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_117
timestamp 1704896540
transform 1 0 11316 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_133
timestamp 1704896540
transform 1 0 12788 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_139
timestamp 1704896540
transform 1 0 13340 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_153
timestamp 1704896540
transform 1 0 14628 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_164
timestamp 1704896540
transform 1 0 15640 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_208
timestamp 1704896540
transform 1 0 19688 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_216
timestamp 1704896540
transform 1 0 20424 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_222
timestamp 1704896540
transform 1 0 20976 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_248
timestamp 1704896540
transform 1 0 23368 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_258
timestamp 1704896540
transform 1 0 24288 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_3
timestamp 1704896540
transform 1 0 828 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_24
timestamp 1704896540
transform 1 0 2760 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_29
timestamp 1704896540
transform 1 0 3220 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_41
timestamp 1704896540
transform 1 0 4324 0 1 21216
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_51
timestamp 1704896540
transform 1 0 5244 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_63
timestamp 1704896540
transform 1 0 6348 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_81
timestamp 1704896540
transform 1 0 8004 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_85
timestamp 1704896540
transform 1 0 8372 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_96
timestamp 1704896540
transform 1 0 9384 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_102
timestamp 1704896540
transform 1 0 9936 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_119
timestamp 1704896540
transform 1 0 11500 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_123
timestamp 1704896540
transform 1 0 11868 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_131
timestamp 1704896540
transform 1 0 12604 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_139
timestamp 1704896540
transform 1 0 13340 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_141
timestamp 1704896540
transform 1 0 13524 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_151
timestamp 1704896540
transform 1 0 14444 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_170
timestamp 1704896540
transform 1 0 16192 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_174
timestamp 1704896540
transform 1 0 16560 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_191
timestamp 1704896540
transform 1 0 18124 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_195
timestamp 1704896540
transform 1 0 18492 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_197
timestamp 1704896540
transform 1 0 18676 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_201
timestamp 1704896540
transform 1 0 19044 0 1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_211
timestamp 1704896540
transform 1 0 19964 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_223
timestamp 1704896540
transform 1 0 21068 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_247
timestamp 1704896540
transform 1 0 23276 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_267
timestamp 1704896540
transform 1 0 25116 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_3
timestamp 1704896540
transform 1 0 828 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_10
timestamp 1704896540
transform 1 0 1472 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_18
timestamp 1704896540
transform 1 0 2208 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_25
timestamp 1704896540
transform 1 0 2852 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_31
timestamp 1704896540
transform 1 0 3404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_39
timestamp 1704896540
transform 1 0 4140 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_47
timestamp 1704896540
transform 1 0 4876 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_67
timestamp 1704896540
transform 1 0 6716 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_81
timestamp 1704896540
transform 1 0 8004 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_87
timestamp 1704896540
transform 1 0 8556 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_113
timestamp 1704896540
transform 1 0 10948 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_117
timestamp 1704896540
transform 1 0 11316 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_134
timestamp 1704896540
transform 1 0 12880 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_181
timestamp 1704896540
transform 1 0 17204 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_185
timestamp 1704896540
transform 1 0 17572 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_193
timestamp 1704896540
transform 1 0 18308 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_209
timestamp 1704896540
transform 1 0 19780 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_217
timestamp 1704896540
transform 1 0 20516 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 1704896540
transform 1 0 21068 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_233
timestamp 1704896540
transform 1 0 21988 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_252
timestamp 1704896540
transform 1 0 23736 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_260
timestamp 1704896540
transform 1 0 24472 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_279
timestamp 1704896540
transform 1 0 26220 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_26
timestamp 1704896540
transform 1 0 2944 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_29
timestamp 1704896540
transform 1 0 3220 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_54
timestamp 1704896540
transform 1 0 5520 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_78
timestamp 1704896540
transform 1 0 7728 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_85
timestamp 1704896540
transform 1 0 8372 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_91
timestamp 1704896540
transform 1 0 8924 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_107
timestamp 1704896540
transform 1 0 10396 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_136
timestamp 1704896540
transform 1 0 13064 0 1 22304
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_150
timestamp 1704896540
transform 1 0 14352 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_162
timestamp 1704896540
transform 1 0 15456 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_170
timestamp 1704896540
transform 1 0 16192 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 1704896540
transform 1 0 18492 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_200
timestamp 1704896540
transform 1 0 18952 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_208
timestamp 1704896540
transform 1 0 19688 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_248
timestamp 1704896540
transform 1 0 23368 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_269
timestamp 1704896540
transform 1 0 25300 0 1 22304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1704896540
transform 1 0 828 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_15
timestamp 1704896540
transform 1 0 1932 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_38
timestamp 1704896540
transform 1 0 4048 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_42
timestamp 1704896540
transform 1 0 4416 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_50
timestamp 1704896540
transform 1 0 5152 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_63
timestamp 1704896540
transform 1 0 6348 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_67
timestamp 1704896540
transform 1 0 6716 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_76
timestamp 1704896540
transform 1 0 7544 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_98
timestamp 1704896540
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 1704896540
transform 1 0 10764 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_113
timestamp 1704896540
transform 1 0 10948 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_138
timestamp 1704896540
transform 1 0 13248 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_146
timestamp 1704896540
transform 1 0 13984 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_161
timestamp 1704896540
transform 1 0 15364 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_167
timestamp 1704896540
transform 1 0 15916 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_185
timestamp 1704896540
transform 1 0 17572 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_219
timestamp 1704896540
transform 1 0 20700 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 1704896540
transform 1 0 21068 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_248
timestamp 1704896540
transform 1 0 23368 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_261
timestamp 1704896540
transform 1 0 24564 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_19
timestamp 1704896540
transform 1 0 2300 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_29
timestamp 1704896540
transform 1 0 3220 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_33
timestamp 1704896540
transform 1 0 3588 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_41
timestamp 1704896540
transform 1 0 4324 0 1 23392
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_56
timestamp 1704896540
transform 1 0 5704 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_68
timestamp 1704896540
transform 1 0 6808 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_85
timestamp 1704896540
transform 1 0 8372 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_101
timestamp 1704896540
transform 1 0 9844 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_137
timestamp 1704896540
transform 1 0 13156 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_152
timestamp 1704896540
transform 1 0 14536 0 1 23392
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_166
timestamp 1704896540
transform 1 0 15824 0 1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_178
timestamp 1704896540
transform 1 0 16928 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_190
timestamp 1704896540
transform 1 0 18032 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_201
timestamp 1704896540
transform 1 0 19044 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_209
timestamp 1704896540
transform 1 0 19780 0 1 23392
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_218
timestamp 1704896540
transform 1 0 20608 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_230
timestamp 1704896540
transform 1 0 21712 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_234
timestamp 1704896540
transform 1 0 22080 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_246
timestamp 1704896540
transform 1 0 23184 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_253
timestamp 1704896540
transform 1 0 23828 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_267
timestamp 1704896540
transform 1 0 25116 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_3
timestamp 1704896540
transform 1 0 828 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_8
timestamp 1704896540
transform 1 0 1288 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_45
timestamp 1704896540
transform 1 0 4692 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_57
timestamp 1704896540
transform 1 0 5796 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_86
timestamp 1704896540
transform 1 0 8464 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_95
timestamp 1704896540
transform 1 0 9292 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_128
timestamp 1704896540
transform 1 0 12328 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_166
timestamp 1704896540
transform 1 0 15824 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_173
timestamp 1704896540
transform 1 0 16468 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_189
timestamp 1704896540
transform 1 0 17940 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_198
timestamp 1704896540
transform 1 0 18768 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_205
timestamp 1704896540
transform 1 0 19412 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_251
timestamp 1704896540
transform 1 0 23644 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_256
timestamp 1704896540
transform 1 0 24104 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_263
timestamp 1704896540
transform 1 0 24748 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_273
timestamp 1704896540
transform 1 0 25668 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_279
timestamp 1704896540
transform 1 0 26220 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_26
timestamp 1704896540
transform 1 0 2944 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_34
timestamp 1704896540
transform 1 0 3680 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_42
timestamp 1704896540
transform 1 0 4416 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_60
timestamp 1704896540
transform 1 0 6072 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_79
timestamp 1704896540
transform 1 0 7820 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1704896540
transform 1 0 8188 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_116
timestamp 1704896540
transform 1 0 11224 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_120
timestamp 1704896540
transform 1 0 11592 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_137
timestamp 1704896540
transform 1 0 13156 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_141
timestamp 1704896540
transform 1 0 13524 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_151
timestamp 1704896540
transform 1 0 14444 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_165
timestamp 1704896540
transform 1 0 15732 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_186
timestamp 1704896540
transform 1 0 17664 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_194
timestamp 1704896540
transform 1 0 18400 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_235
timestamp 1704896540
transform 1 0 22172 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_239
timestamp 1704896540
transform 1 0 22540 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_288
timestamp 1704896540
transform 1 0 27048 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_3
timestamp 1704896540
transform 1 0 828 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_8
timestamp 1704896540
transform 1 0 1288 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_16
timestamp 1704896540
transform 1 0 2024 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_23
timestamp 1704896540
transform 1 0 2668 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_36
timestamp 1704896540
transform 1 0 3864 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_42
timestamp 1704896540
transform 1 0 4416 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 1704896540
transform 1 0 5244 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1704896540
transform 1 0 5612 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_57
timestamp 1704896540
transform 1 0 5796 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_65
timestamp 1704896540
transform 1 0 6532 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_71
timestamp 1704896540
transform 1 0 7084 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_79
timestamp 1704896540
transform 1 0 7820 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_104
timestamp 1704896540
transform 1 0 10120 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_113
timestamp 1704896540
transform 1 0 10948 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_121
timestamp 1704896540
transform 1 0 11684 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_129
timestamp 1704896540
transform 1 0 12420 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_150
timestamp 1704896540
transform 1 0 14352 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_159
timestamp 1704896540
transform 1 0 15180 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_166
timestamp 1704896540
transform 1 0 15824 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_169
timestamp 1704896540
transform 1 0 16100 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_178
timestamp 1704896540
transform 1 0 16928 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_186
timestamp 1704896540
transform 1 0 17664 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_195
timestamp 1704896540
transform 1 0 18492 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_204
timestamp 1704896540
transform 1 0 19320 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_223
timestamp 1704896540
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_233
timestamp 1704896540
transform 1 0 21988 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_245
timestamp 1704896540
transform 1 0 23092 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_259
timestamp 1704896540
transform 1 0 24380 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_263
timestamp 1704896540
transform 1 0 24748 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_3
timestamp 1704896540
transform 1 0 828 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_12
timestamp 1704896540
transform 1 0 1656 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_45
timestamp 1704896540
transform 1 0 4692 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_82
timestamp 1704896540
transform 1 0 8096 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_136
timestamp 1704896540
transform 1 0 13064 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_149
timestamp 1704896540
transform 1 0 14260 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_157
timestamp 1704896540
transform 1 0 14996 0 1 25568
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_175
timestamp 1704896540
transform 1 0 16652 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_187
timestamp 1704896540
transform 1 0 17756 0 1 25568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_200
timestamp 1704896540
transform 1 0 18952 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_212
timestamp 1704896540
transform 1 0 20056 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_236
timestamp 1704896540
transform 1 0 22264 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_243
timestamp 1704896540
transform 1 0 22908 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_250
timestamp 1704896540
transform 1 0 23552 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_256
timestamp 1704896540
transform 1 0 24104 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_3
timestamp 1704896540
transform 1 0 828 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_32
timestamp 1704896540
transform 1 0 3496 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_36
timestamp 1704896540
transform 1 0 3864 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_44
timestamp 1704896540
transform 1 0 4600 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 1704896540
transform 1 0 5612 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_57
timestamp 1704896540
transform 1 0 5796 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_79
timestamp 1704896540
transform 1 0 7820 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 1704896540
transform 1 0 10764 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_113
timestamp 1704896540
transform 1 0 10948 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_138
timestamp 1704896540
transform 1 0 13248 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_151
timestamp 1704896540
transform 1 0 14444 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_159
timestamp 1704896540
transform 1 0 15180 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_167
timestamp 1704896540
transform 1 0 15916 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_169
timestamp 1704896540
transform 1 0 16100 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_177
timestamp 1704896540
transform 1 0 16836 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_182
timestamp 1704896540
transform 1 0 17296 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_186
timestamp 1704896540
transform 1 0 17664 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_192
timestamp 1704896540
transform 1 0 18216 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_210
timestamp 1704896540
transform 1 0 19872 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_218
timestamp 1704896540
transform 1 0 20608 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_222
timestamp 1704896540
transform 1 0 20976 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_234
timestamp 1704896540
transform 1 0 22080 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_243
timestamp 1704896540
transform 1 0 22908 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_259
timestamp 1704896540
transform 1 0 24380 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_281
timestamp 1704896540
transform 1 0 26404 0 -1 26656
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 1704896540
transform 1 0 828 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_15
timestamp 1704896540
transform 1 0 1932 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_23
timestamp 1704896540
transform 1 0 2668 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1704896540
transform 1 0 3036 0 1 26656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 1704896540
transform 1 0 3220 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_41
timestamp 1704896540
transform 1 0 4324 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_62
timestamp 1704896540
transform 1 0 6256 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_66
timestamp 1704896540
transform 1 0 6624 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_82
timestamp 1704896540
transform 1 0 8096 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_90
timestamp 1704896540
transform 1 0 8832 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_107
timestamp 1704896540
transform 1 0 10396 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_149
timestamp 1704896540
transform 1 0 14260 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_157
timestamp 1704896540
transform 1 0 14996 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_171
timestamp 1704896540
transform 1 0 16284 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_195
timestamp 1704896540
transform 1 0 18492 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_203
timestamp 1704896540
transform 1 0 19228 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_222
timestamp 1704896540
transform 1 0 20976 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_242
timestamp 1704896540
transform 1 0 22816 0 1 26656
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_253
timestamp 1704896540
transform 1 0 23828 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_265
timestamp 1704896540
transform 1 0 24932 0 1 26656
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 1704896540
transform 1 0 828 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_15
timestamp 1704896540
transform 1 0 1932 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_47
timestamp 1704896540
transform 1 0 4876 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_54
timestamp 1704896540
transform 1 0 5520 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_73
timestamp 1704896540
transform 1 0 7268 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_82
timestamp 1704896540
transform 1 0 8096 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_109
timestamp 1704896540
transform 1 0 10580 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_129
timestamp 1704896540
transform 1 0 12420 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_149
timestamp 1704896540
transform 1 0 14260 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_166
timestamp 1704896540
transform 1 0 15824 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_169
timestamp 1704896540
transform 1 0 16100 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_173
timestamp 1704896540
transform 1 0 16468 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_190
timestamp 1704896540
transform 1 0 18032 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_215
timestamp 1704896540
transform 1 0 20332 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_223
timestamp 1704896540
transform 1 0 21068 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_236
timestamp 1704896540
transform 1 0 22264 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_247
timestamp 1704896540
transform 1 0 23276 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_255
timestamp 1704896540
transform 1 0 24012 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_276
timestamp 1704896540
transform 1 0 25944 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_281
timestamp 1704896540
transform 1 0 26404 0 -1 27744
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1704896540
transform 1 0 828 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_15
timestamp 1704896540
transform 1 0 1932 0 1 27744
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_49
timestamp 1704896540
transform 1 0 5060 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_61
timestamp 1704896540
transform 1 0 6164 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_65
timestamp 1704896540
transform 1 0 6532 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_70
timestamp 1704896540
transform 1 0 6992 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_83
timestamp 1704896540
transform 1 0 8188 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_85
timestamp 1704896540
transform 1 0 8372 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_89
timestamp 1704896540
transform 1 0 8740 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_121
timestamp 1704896540
transform 1 0 11684 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_139
timestamp 1704896540
transform 1 0 13340 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_144
timestamp 1704896540
transform 1 0 13800 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_152
timestamp 1704896540
transform 1 0 14536 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_170
timestamp 1704896540
transform 1 0 16192 0 1 27744
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_197
timestamp 1704896540
transform 1 0 18676 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_260
timestamp 1704896540
transform 1 0 24472 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_3
timestamp 1704896540
transform 1 0 828 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_11
timestamp 1704896540
transform 1 0 1564 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_30
timestamp 1704896540
transform 1 0 3312 0 -1 28832
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_43
timestamp 1704896540
transform 1 0 4508 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 1704896540
transform 1 0 5612 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_79
timestamp 1704896540
transform 1 0 7820 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_129
timestamp 1704896540
transform 1 0 12420 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_166
timestamp 1704896540
transform 1 0 15824 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_169
timestamp 1704896540
transform 1 0 16100 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_176
timestamp 1704896540
transform 1 0 16744 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_205
timestamp 1704896540
transform 1 0 19412 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_222
timestamp 1704896540
transform 1 0 20976 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_241
timestamp 1704896540
transform 1 0 22724 0 -1 28832
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_246
timestamp 1704896540
transform 1 0 23184 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_258
timestamp 1704896540
transform 1 0 24288 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_278
timestamp 1704896540
transform 1 0 26128 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_281
timestamp 1704896540
transform 1 0 26404 0 -1 28832
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_3
timestamp 1704896540
transform 1 0 828 0 1 28832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_15
timestamp 1704896540
transform 1 0 1932 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 1704896540
transform 1 0 3036 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_29
timestamp 1704896540
transform 1 0 3220 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_33
timestamp 1704896540
transform 1 0 3588 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_37
timestamp 1704896540
transform 1 0 3956 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_45
timestamp 1704896540
transform 1 0 4692 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_54
timestamp 1704896540
transform 1 0 5520 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_62
timestamp 1704896540
transform 1 0 6256 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_85
timestamp 1704896540
transform 1 0 8372 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_115
timestamp 1704896540
transform 1 0 11132 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_136
timestamp 1704896540
transform 1 0 13064 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_147
timestamp 1704896540
transform 1 0 14076 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_155
timestamp 1704896540
transform 1 0 14812 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_159
timestamp 1704896540
transform 1 0 15180 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_168
timestamp 1704896540
transform 1 0 16008 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_188
timestamp 1704896540
transform 1 0 17848 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_207
timestamp 1704896540
transform 1 0 19596 0 1 28832
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_230
timestamp 1704896540
transform 1 0 21712 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_242
timestamp 1704896540
transform 1 0 22816 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_250
timestamp 1704896540
transform 1 0 23552 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_266
timestamp 1704896540
transform 1 0 25024 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_285
timestamp 1704896540
transform 1 0 26772 0 1 28832
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 1704896540
transform 1 0 828 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_39
timestamp 1704896540
transform 1 0 4140 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 1704896540
transform 1 0 5612 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_62
timestamp 1704896540
transform 1 0 6256 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_85
timestamp 1704896540
transform 1 0 8372 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_100
timestamp 1704896540
transform 1 0 9752 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_110
timestamp 1704896540
transform 1 0 10672 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_147
timestamp 1704896540
transform 1 0 14076 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_161
timestamp 1704896540
transform 1 0 15364 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_183
timestamp 1704896540
transform 1 0 17388 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_200
timestamp 1704896540
transform 1 0 18952 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_204
timestamp 1704896540
transform 1 0 19320 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_221
timestamp 1704896540
transform 1 0 20884 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_272
timestamp 1704896540
transform 1 0 25576 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_281
timestamp 1704896540
transform 1 0 26404 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_3
timestamp 1704896540
transform 1 0 828 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_29
timestamp 1704896540
transform 1 0 3220 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_83
timestamp 1704896540
transform 1 0 8188 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_85
timestamp 1704896540
transform 1 0 8372 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_103
timestamp 1704896540
transform 1 0 10028 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_139
timestamp 1704896540
transform 1 0 13340 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_141
timestamp 1704896540
transform 1 0 13524 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_163
timestamp 1704896540
transform 1 0 15548 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_178
timestamp 1704896540
transform 1 0 16928 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_195
timestamp 1704896540
transform 1 0 18492 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_197
timestamp 1704896540
transform 1 0 18676 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_203
timestamp 1704896540
transform 1 0 19228 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_224
timestamp 1704896540
transform 1 0 21160 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_251
timestamp 1704896540
transform 1 0 23644 0 1 29920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_266
timestamp 1704896540
transform 1 0 25024 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_278
timestamp 1704896540
transform 1 0 26128 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_286
timestamp 1704896540
transform 1 0 26864 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_20
timestamp 1704896540
transform 1 0 2392 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_29
timestamp 1704896540
transform 1 0 3220 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_33
timestamp 1704896540
transform 1 0 3588 0 -1 31008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_37
timestamp 1704896540
transform 1 0 3956 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_49
timestamp 1704896540
transform 1 0 5060 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_55
timestamp 1704896540
transform 1 0 5612 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_57
timestamp 1704896540
transform 1 0 5796 0 -1 31008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_61
timestamp 1704896540
transform 1 0 6164 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_73
timestamp 1704896540
transform 1 0 7268 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_77
timestamp 1704896540
transform 1 0 7636 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_83
timestamp 1704896540
transform 1 0 8188 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_88
timestamp 1704896540
transform 1 0 8648 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_93
timestamp 1704896540
transform 1 0 9108 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_131
timestamp 1704896540
transform 1 0 12604 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_139
timestamp 1704896540
transform 1 0 13340 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_153
timestamp 1704896540
transform 1 0 14628 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_161
timestamp 1704896540
transform 1 0 15364 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_167
timestamp 1704896540
transform 1 0 15916 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_169
timestamp 1704896540
transform 1 0 16100 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_173
timestamp 1704896540
transform 1 0 16468 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_177
timestamp 1704896540
transform 1 0 16836 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_181
timestamp 1704896540
transform 1 0 17204 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_185
timestamp 1704896540
transform 1 0 17572 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_193
timestamp 1704896540
transform 1 0 18308 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_197
timestamp 1704896540
transform 1 0 18676 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_222
timestamp 1704896540
transform 1 0 20976 0 -1 31008
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_257
timestamp 1704896540
transform 1 0 24196 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_269
timestamp 1704896540
transform 1 0 25300 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_277
timestamp 1704896540
transform 1 0 26036 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_281
timestamp 1704896540
transform 1 0 26404 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_285
timestamp 1704896540
transform 1 0 26772 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11132 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1704896540
transform -1 0 11132 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1704896540
transform 1 0 8372 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1704896540
transform -1 0 14260 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1704896540
transform -1 0 25668 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1704896540
transform -1 0 23000 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1704896540
transform 1 0 25116 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1704896540
transform -1 0 24748 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1704896540
transform -1 0 5888 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1704896540
transform -1 0 20148 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1704896540
transform -1 0 12420 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1704896540
transform -1 0 14260 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1704896540
transform -1 0 9844 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1704896540
transform 1 0 11224 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1704896540
transform -1 0 13248 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1704896540
transform -1 0 23736 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1704896540
transform 1 0 8924 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1704896540
transform -1 0 20424 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1704896540
transform 1 0 9384 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1704896540
transform -1 0 13064 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1704896540
transform -1 0 22540 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1704896540
transform -1 0 10212 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1704896540
transform 1 0 8372 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1704896540
transform -1 0 10856 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1704896540
transform 1 0 11132 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1704896540
transform -1 0 23000 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1704896540
transform -1 0 21988 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1704896540
transform -1 0 21988 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1704896540
transform -1 0 10856 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1704896540
transform -1 0 10396 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1704896540
transform -1 0 12604 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1704896540
transform -1 0 11684 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1704896540
transform -1 0 10764 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1704896540
transform -1 0 10028 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1704896540
transform -1 0 12696 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1704896540
transform -1 0 11960 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1704896540
transform -1 0 11684 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1704896540
transform 1 0 10488 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1704896540
transform 1 0 22356 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1704896540
transform -1 0 14260 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1704896540
transform -1 0 19320 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1704896540
transform -1 0 10856 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1704896540
transform 1 0 22724 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1704896540
transform -1 0 3956 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1704896540
transform -1 0 23644 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1704896540
transform 1 0 16468 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1704896540
transform -1 0 21436 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1704896540
transform -1 0 24564 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1704896540
transform 1 0 4968 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1704896540
transform -1 0 6624 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1704896540
transform -1 0 20700 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1704896540
transform -1 0 10304 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1704896540
transform 1 0 10304 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1704896540
transform -1 0 2484 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1704896540
transform -1 0 1748 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1704896540
transform -1 0 21988 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1704896540
transform -1 0 20976 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1704896540
transform 1 0 8740 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1704896540
transform 1 0 16836 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1704896540
transform -1 0 2944 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1704896540
transform -1 0 2208 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1704896540
transform -1 0 3956 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1704896540
transform 1 0 2208 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1704896540
transform -1 0 3220 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1704896540
transform 1 0 1748 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1704896540
transform -1 0 10120 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1704896540
transform -1 0 6624 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1704896540
transform 1 0 4600 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1704896540
transform 1 0 6348 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1704896540
transform -1 0 14996 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1704896540
transform -1 0 14260 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1704896540
transform 1 0 5612 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1704896540
transform 1 0 4140 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1704896540
transform -1 0 4232 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1704896540
transform -1 0 8188 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1704896540
transform -1 0 4784 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1704896540
transform 1 0 3312 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1704896540
transform 1 0 1472 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1704896540
transform -1 0 2944 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1704896540
transform -1 0 1656 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1704896540
transform -1 0 5428 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1704896540
transform -1 0 3128 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1704896540
transform -1 0 4508 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 1704896540
transform -1 0 7176 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1704896540
transform -1 0 21988 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 1704896540
transform -1 0 5428 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1704896540
transform 1 0 21620 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 1704896540
transform -1 0 7176 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 1704896540
transform -1 0 27140 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1704896540
transform -1 0 4140 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 1704896540
transform -1 0 3036 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 1704896540
transform -1 0 17756 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 1704896540
transform -1 0 8096 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 1704896540
transform -1 0 25484 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 1704896540
transform 1 0 19228 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 1704896540
transform -1 0 11684 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 1704896540
transform -1 0 16836 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 1704896540
transform -1 0 21804 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 1704896540
transform 1 0 21252 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 1704896540
transform -1 0 27140 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 1704896540
transform -1 0 9844 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 1704896540
transform -1 0 8464 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 1704896540
transform -1 0 1932 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 1704896540
transform 1 0 14812 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 1704896540
transform -1 0 23184 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 1704896540
transform -1 0 9016 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 1704896540
transform 1 0 10948 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 1704896540
transform -1 0 7636 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 1704896540
transform -1 0 11224 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1704896540
transform 1 0 8832 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1704896540
transform -1 0 11224 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1704896540
transform 1 0 7360 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1704896540
transform 1 0 5888 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 1704896540
transform -1 0 21620 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input6
timestamp 1704896540
transform 1 0 20792 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1704896540
transform 1 0 19872 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1704896540
transform -1 0 18032 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1704896540
transform -1 0 16468 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input10
timestamp 1704896540
transform 1 0 14720 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input11
timestamp 1704896540
transform 1 0 14260 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input12
timestamp 1704896540
transform 1 0 11960 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1704896540
transform -1 0 26772 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input14
timestamp 1704896540
transform 1 0 23828 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1704896540
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1704896540
transform -1 0 27416 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1704896540
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1704896540
transform -1 0 27416 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1704896540
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1704896540
transform -1 0 27416 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1704896540
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1704896540
transform -1 0 27416 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1704896540
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1704896540
transform -1 0 27416 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1704896540
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1704896540
transform -1 0 27416 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1704896540
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1704896540
transform -1 0 27416 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1704896540
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1704896540
transform -1 0 27416 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1704896540
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1704896540
transform -1 0 27416 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1704896540
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1704896540
transform -1 0 27416 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1704896540
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1704896540
transform -1 0 27416 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1704896540
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1704896540
transform -1 0 27416 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1704896540
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1704896540
transform -1 0 27416 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1704896540
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1704896540
transform -1 0 27416 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1704896540
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1704896540
transform -1 0 27416 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1704896540
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1704896540
transform -1 0 27416 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1704896540
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1704896540
transform -1 0 27416 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1704896540
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1704896540
transform -1 0 27416 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1704896540
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1704896540
transform -1 0 27416 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1704896540
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1704896540
transform -1 0 27416 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1704896540
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1704896540
transform -1 0 27416 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1704896540
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1704896540
transform -1 0 27416 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1704896540
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1704896540
transform -1 0 27416 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1704896540
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1704896540
transform -1 0 27416 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1704896540
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1704896540
transform -1 0 27416 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1704896540
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1704896540
transform -1 0 27416 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1704896540
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1704896540
transform -1 0 27416 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1704896540
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1704896540
transform -1 0 27416 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1704896540
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1704896540
transform -1 0 27416 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1704896540
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1704896540
transform -1 0 27416 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1704896540
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1704896540
transform -1 0 27416 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1704896540
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1704896540
transform -1 0 27416 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1704896540
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1704896540
transform -1 0 27416 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1704896540
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1704896540
transform -1 0 27416 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1704896540
transform 1 0 552 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1704896540
transform -1 0 27416 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1704896540
transform 1 0 552 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1704896540
transform -1 0 27416 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1704896540
transform 1 0 552 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1704896540
transform -1 0 27416 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1704896540
transform 1 0 552 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1704896540
transform -1 0 27416 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1704896540
transform 1 0 552 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1704896540
transform -1 0 27416 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1704896540
transform 1 0 552 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1704896540
transform -1 0 27416 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1704896540
transform 1 0 552 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1704896540
transform -1 0 27416 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1704896540
transform 1 0 552 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1704896540
transform -1 0 27416 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1704896540
transform 1 0 552 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1704896540
transform -1 0 27416 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1704896540
transform 1 0 552 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1704896540
transform -1 0 27416 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1704896540
transform 1 0 552 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1704896540
transform -1 0 27416 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1704896540
transform 1 0 552 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1704896540
transform -1 0 27416 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1704896540
transform 1 0 552 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1704896540
transform -1 0 27416 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1704896540
transform 1 0 552 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1704896540
transform -1 0 27416 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1704896540
transform 1 0 552 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1704896540
transform -1 0 27416 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1704896540
transform 1 0 552 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1704896540
transform -1 0 27416 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1704896540
transform 1 0 552 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1704896540
transform -1 0 27416 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1704896540
transform 1 0 552 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1704896540
transform -1 0 27416 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1704896540
transform 1 0 552 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1704896540
transform -1 0 27416 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1704896540
transform 1 0 552 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1704896540
transform -1 0 27416 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1704896540
transform 1 0 552 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1704896540
transform -1 0 27416 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1704896540
transform 1 0 552 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1704896540
transform -1 0 27416 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1704896540
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1704896540
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1704896540
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1704896540
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1704896540
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1704896540
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1704896540
transform 1 0 21160 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1704896540
transform 1 0 23736 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1704896540
transform 1 0 26312 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1704896540
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1704896540
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1704896540
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1704896540
transform 1 0 21160 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1704896540
transform 1 0 26312 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1704896540
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1704896540
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1704896540
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1704896540
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1704896540
transform 1 0 23736 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1704896540
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1704896540
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1704896540
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1704896540
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1704896540
transform 1 0 26312 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1704896540
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1704896540
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1704896540
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1704896540
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1704896540
transform 1 0 23736 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1704896540
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1704896540
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1704896540
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1704896540
transform 1 0 21160 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1704896540
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1704896540
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1704896540
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1704896540
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1704896540
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1704896540
transform 1 0 23736 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1704896540
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1704896540
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1704896540
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1704896540
transform 1 0 21160 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1704896540
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1704896540
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1704896540
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1704896540
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1704896540
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1704896540
transform 1 0 23736 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1704896540
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1704896540
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1704896540
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1704896540
transform 1 0 21160 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1704896540
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1704896540
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1704896540
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1704896540
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1704896540
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1704896540
transform 1 0 23736 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1704896540
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1704896540
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1704896540
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1704896540
transform 1 0 21160 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1704896540
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1704896540
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1704896540
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1704896540
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1704896540
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1704896540
transform 1 0 23736 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1704896540
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1704896540
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1704896540
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1704896540
transform 1 0 21160 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1704896540
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1704896540
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1704896540
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1704896540
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1704896540
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1704896540
transform 1 0 23736 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1704896540
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1704896540
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1704896540
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1704896540
transform 1 0 21160 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1704896540
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1704896540
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1704896540
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1704896540
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1704896540
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1704896540
transform 1 0 23736 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1704896540
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1704896540
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1704896540
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1704896540
transform 1 0 21160 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1704896540
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1704896540
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1704896540
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1704896540
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1704896540
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1704896540
transform 1 0 23736 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1704896540
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1704896540
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1704896540
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1704896540
transform 1 0 21160 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1704896540
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1704896540
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1704896540
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1704896540
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1704896540
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1704896540
transform 1 0 23736 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1704896540
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1704896540
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1704896540
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1704896540
transform 1 0 21160 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1704896540
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1704896540
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1704896540
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1704896540
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1704896540
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1704896540
transform 1 0 23736 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1704896540
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1704896540
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1704896540
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1704896540
transform 1 0 21160 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1704896540
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1704896540
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1704896540
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1704896540
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1704896540
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1704896540
transform 1 0 23736 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1704896540
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1704896540
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1704896540
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1704896540
transform 1 0 21160 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1704896540
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1704896540
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1704896540
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1704896540
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1704896540
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1704896540
transform 1 0 23736 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1704896540
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1704896540
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1704896540
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1704896540
transform 1 0 21160 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1704896540
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1704896540
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1704896540
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1704896540
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1704896540
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1704896540
transform 1 0 23736 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1704896540
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1704896540
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1704896540
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1704896540
transform 1 0 21160 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1704896540
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1704896540
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1704896540
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1704896540
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1704896540
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1704896540
transform 1 0 23736 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1704896540
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1704896540
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1704896540
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1704896540
transform 1 0 21160 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1704896540
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1704896540
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1704896540
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1704896540
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1704896540
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1704896540
transform 1 0 23736 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1704896540
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1704896540
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1704896540
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1704896540
transform 1 0 21160 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1704896540
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1704896540
transform 1 0 3128 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1704896540
transform 1 0 8280 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1704896540
transform 1 0 13432 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1704896540
transform 1 0 18584 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1704896540
transform 1 0 23736 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1704896540
transform 1 0 5704 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1704896540
transform 1 0 10856 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1704896540
transform 1 0 16008 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1704896540
transform 1 0 21160 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1704896540
transform 1 0 26312 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1704896540
transform 1 0 3128 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1704896540
transform 1 0 8280 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1704896540
transform 1 0 13432 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1704896540
transform 1 0 18584 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1704896540
transform 1 0 23736 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1704896540
transform 1 0 5704 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1704896540
transform 1 0 10856 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1704896540
transform 1 0 16008 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1704896540
transform 1 0 21160 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1704896540
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1704896540
transform 1 0 3128 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1704896540
transform 1 0 8280 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1704896540
transform 1 0 13432 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1704896540
transform 1 0 18584 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1704896540
transform 1 0 23736 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1704896540
transform 1 0 5704 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1704896540
transform 1 0 10856 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1704896540
transform 1 0 16008 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1704896540
transform 1 0 21160 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1704896540
transform 1 0 26312 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1704896540
transform 1 0 3128 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1704896540
transform 1 0 8280 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1704896540
transform 1 0 13432 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1704896540
transform 1 0 18584 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1704896540
transform 1 0 23736 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1704896540
transform 1 0 5704 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1704896540
transform 1 0 10856 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1704896540
transform 1 0 16008 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1704896540
transform 1 0 21160 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1704896540
transform 1 0 26312 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1704896540
transform 1 0 3128 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1704896540
transform 1 0 8280 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1704896540
transform 1 0 13432 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1704896540
transform 1 0 18584 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1704896540
transform 1 0 23736 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1704896540
transform 1 0 5704 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1704896540
transform 1 0 10856 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1704896540
transform 1 0 16008 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1704896540
transform 1 0 21160 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1704896540
transform 1 0 26312 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1704896540
transform 1 0 3128 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1704896540
transform 1 0 8280 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1704896540
transform 1 0 13432 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1704896540
transform 1 0 18584 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1704896540
transform 1 0 23736 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1704896540
transform 1 0 5704 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1704896540
transform 1 0 10856 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1704896540
transform 1 0 16008 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1704896540
transform 1 0 21160 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1704896540
transform 1 0 26312 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1704896540
transform 1 0 3128 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1704896540
transform 1 0 8280 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1704896540
transform 1 0 13432 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1704896540
transform 1 0 18584 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1704896540
transform 1 0 23736 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1704896540
transform 1 0 5704 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1704896540
transform 1 0 10856 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1704896540
transform 1 0 16008 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1704896540
transform 1 0 21160 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1704896540
transform 1 0 26312 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1704896540
transform 1 0 3128 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1704896540
transform 1 0 8280 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1704896540
transform 1 0 13432 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1704896540
transform 1 0 18584 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1704896540
transform 1 0 23736 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1704896540
transform 1 0 5704 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1704896540
transform 1 0 10856 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1704896540
transform 1 0 16008 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1704896540
transform 1 0 21160 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1704896540
transform 1 0 26312 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1704896540
transform 1 0 3128 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1704896540
transform 1 0 8280 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1704896540
transform 1 0 13432 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1704896540
transform 1 0 18584 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1704896540
transform 1 0 23736 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1704896540
transform 1 0 5704 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1704896540
transform 1 0 10856 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1704896540
transform 1 0 16008 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1704896540
transform 1 0 21160 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1704896540
transform 1 0 26312 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1704896540
transform 1 0 3128 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1704896540
transform 1 0 8280 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1704896540
transform 1 0 13432 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1704896540
transform 1 0 18584 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1704896540
transform 1 0 23736 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1704896540
transform 1 0 5704 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1704896540
transform 1 0 10856 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1704896540
transform 1 0 16008 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1704896540
transform 1 0 21160 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1704896540
transform 1 0 26312 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1704896540
transform 1 0 3128 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1704896540
transform 1 0 8280 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1704896540
transform 1 0 13432 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1704896540
transform 1 0 18584 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1704896540
transform 1 0 23736 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1704896540
transform 1 0 3128 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1704896540
transform 1 0 5704 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1704896540
transform 1 0 8280 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1704896540
transform 1 0 10856 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1704896540
transform 1 0 13432 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1704896540
transform 1 0 16008 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1704896540
transform 1 0 18584 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1704896540
transform 1 0 21160 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1704896540
transform 1 0 23736 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1704896540
transform 1 0 26312 0 -1 31008
box -38 -48 130 592
<< labels >>
rlabel metal2 s 14064 31008 14064 31008 4 VGND
rlabel metal1 s 13984 30464 13984 30464 4 VPWR
rlabel metal1 s 10534 14348 10534 14348 4 _0003_
rlabel metal1 s 17158 22746 17158 22746 4 _0004_
rlabel metal2 s 18170 20978 18170 20978 4 _0005_
rlabel metal1 s 18062 21046 18062 21046 4 _0006_
rlabel metal2 s 17894 22950 17894 22950 4 _0007_
rlabel metal1 s 19821 18802 19821 18802 4 _0008_
rlabel metal1 s 17516 18802 17516 18802 4 _0009_
rlabel metal1 s 20552 18190 20552 18190 4 _0010_
rlabel metal1 s 17326 19958 17326 19958 4 _0011_
rlabel metal1 s 20470 16762 20470 16762 4 _0012_
rlabel metal1 s 19223 17034 19223 17034 4 _0013_
rlabel metal1 s 19269 20298 19269 20298 4 _0014_
rlabel metal1 s 21486 20366 21486 20366 4 _0015_
rlabel metal1 s 14014 14518 14014 14518 4 _0016_
rlabel metal2 s 17337 13362 17337 13362 4 _0017_
rlabel metal1 s 17786 15606 17786 15606 4 _0018_
rlabel metal1 s 14214 16218 14214 16218 4 _0019_
rlabel metal1 s 15860 13838 15860 13838 4 _0020_
rlabel metal1 s 17475 16626 17475 16626 4 _0021_
rlabel metal2 s 12282 19125 12282 19125 4 _0022_
rlabel metal2 s 11086 20162 11086 20162 4 _0023_
rlabel metal1 s 12838 17714 12838 17714 4 _0024_
rlabel metal1 s 13309 17034 13309 17034 4 _0025_
rlabel metal2 s 11086 16422 11086 16422 4 _0026_
rlabel metal1 s 21965 22406 21965 22406 4 _0027_
rlabel metal2 s 19918 22338 19918 22338 4 _0028_
rlabel metal1 s 21850 20944 21850 20944 4 _0029_
rlabel metal2 s 21758 21216 21758 21216 4 _0030_
rlabel metal1 s 24927 2550 24927 2550 4 _0031_
rlabel metal1 s 26822 4046 26822 4046 4 _0032_
rlabel metal2 s 24513 6222 24513 6222 4 _0033_
rlabel metal1 s 26092 7922 26092 7922 4 _0034_
rlabel metal2 s 22581 7242 22581 7242 4 _0035_
rlabel metal1 s 25304 9486 25304 9486 4 _0036_
rlabel metal1 s 20649 7922 20649 7922 4 _0037_
rlabel metal2 s 22126 9860 22126 9860 4 _0038_
rlabel metal4 s 2093 30396 2093 30396 4 _0039_
rlabel metal2 s 15966 20298 15966 20298 4 _0040_
rlabel metal2 s 12374 20570 12374 20570 4 _0041_
rlabel metal2 s 16141 19278 16141 19278 4 _0042_
rlabel metal1 s 14122 17306 14122 17306 4 _0043_
rlabel metal1 s 13800 29274 13800 29274 4 _0044_
rlabel metal2 s 1145 19278 1145 19278 4 _0045_
rlabel metal1 s 1472 21590 1472 21590 4 _0046_
rlabel metal1 s 2714 21046 2714 21046 4 _0047_
rlabel metal2 s 2806 19006 2806 19006 4 _0048_
rlabel metal2 s 1426 17510 1426 17510 4 _0049_
rlabel metal1 s 4426 16626 4426 16626 4 _0050_
rlabel metal1 s 1697 16626 1697 16626 4 _0051_
rlabel metal1 s 7677 14450 7677 14450 4 _0052_
rlabel metal1 s 7539 14858 7539 14858 4 _0053_
rlabel metal2 s 9430 14722 9430 14722 4 _0054_
rlabel metal1 s 11147 13430 11147 13430 4 _0055_
rlabel metal1 s 8126 25398 8126 25398 4 _0056_
rlabel metal1 s 8862 25738 8862 25738 4 _0057_
rlabel metal1 s 9986 26826 9986 26826 4 _0058_
rlabel metal1 s 9752 27642 9752 27642 4 _0059_
rlabel metal1 s 8924 27642 8924 27642 4 _0060_
rlabel metal1 s 10932 29750 10932 29750 4 _0061_
rlabel metal1 s 11182 30090 11182 30090 4 _0062_
rlabel metal2 s 8694 29682 8694 29682 4 _0063_
rlabel metal2 s 17424 9078 17424 9078 4 _0064_
rlabel metal1 s 19172 9486 19172 9486 4 _0065_
rlabel metal2 s 17986 12070 17986 12070 4 _0066_
rlabel metal1 s 16866 11254 16866 11254 4 _0067_
rlabel metal1 s 20470 12886 20470 12886 4 _0068_
rlabel metal2 s 9246 20502 9246 20502 4 _0069_
rlabel metal1 s 9660 20026 9660 20026 4 _0070_
rlabel metal2 s 8786 21862 8786 21862 4 _0071_
rlabel metal2 s 11182 21454 11182 21454 4 _0072_
rlabel metal1 s 9158 23222 9158 23222 4 _0073_
rlabel metal1 s 10058 23562 10058 23562 4 _0074_
rlabel metal1 s 11147 24310 11147 24310 4 _0075_
rlabel metal2 s 8694 24514 8694 24514 4 _0076_
rlabel metal2 s 12282 13634 12282 13634 4 _0077_
rlabel metal2 s 12742 15300 12742 15300 4 _0078_
rlabel metal1 s 11403 12342 11403 12342 4 _0079_
rlabel metal2 s 12834 13158 12834 13158 4 _0080_
rlabel metal1 s 11898 11254 11898 11254 4 _0081_
rlabel metal1 s 16564 15606 16564 15606 4 _0082_
rlabel metal1 s 16422 21930 16422 21930 4 _0083_
rlabel metal2 s 14214 21862 14214 21862 4 _0084_
rlabel metal2 s 12926 24242 12926 24242 4 _0085_
rlabel metal1 s 16008 24854 16008 24854 4 _0086_
rlabel metal1 s 14347 30158 14347 30158 4 _0087_
rlabel metal2 s 18174 30158 18174 30158 4 _0088_
rlabel metal1 s 18450 29750 18450 29750 4 _0089_
rlabel metal1 s 19002 28662 19002 28662 4 _0090_
rlabel metal1 s 17234 27914 17234 27914 4 _0091_
rlabel metal1 s 19274 27098 19274 27098 4 _0092_
rlabel metal1 s 19228 26010 19228 26010 4 _0093_
rlabel metal1 s 18568 24650 18568 24650 4 _0094_
rlabel metal1 s 19964 12954 19964 12954 4 _0095_
rlabel metal1 s 25438 19482 25438 19482 4 _0096_
rlabel metal1 s 23363 18870 23363 18870 4 _0097_
rlabel metal2 s 25898 19074 25898 19074 4 _0098_
rlabel metal1 s 25944 17850 25944 17850 4 _0099_
rlabel metal2 s 25806 16898 25806 16898 4 _0100_
rlabel metal1 s 26408 16014 26408 16014 4 _0101_
rlabel metal1 s 26500 14926 26500 14926 4 _0102_
rlabel metal1 s 26500 13838 26500 13838 4 _0103_
rlabel metal1 s 26097 13430 26097 13430 4 _0104_
rlabel metal2 s 26638 12682 26638 12682 4 _0105_
rlabel metal2 s 24794 12036 24794 12036 4 _0106_
rlabel metal1 s 24150 12206 24150 12206 4 _0107_
rlabel metal1 s 20802 14926 20802 14926 4 _0108_
rlabel metal2 s 22218 23358 22218 23358 4 _0109_
rlabel metal1 s 20649 25738 20649 25738 4 _0110_
rlabel metal1 s 21620 28934 21620 28934 4 _0111_
rlabel metal1 s 22765 27914 22765 27914 4 _0112_
rlabel metal1 s 25622 28458 25622 28458 4 _0113_
rlabel metal1 s 26454 27914 26454 27914 4 _0114_
rlabel metal1 s 25994 25330 25994 25330 4 _0115_
rlabel metal1 s 26864 25466 26864 25466 4 _0116_
rlabel metal1 s 25698 24650 25698 24650 4 _0117_
rlabel metal2 s 25622 23154 25622 23154 4 _0118_
rlabel metal1 s 26864 22202 26864 22202 4 _0119_
rlabel metal1 s 25948 21046 25948 21046 4 _0120_
rlabel metal1 s 16886 9418 16886 9418 4 _0121_
rlabel metal2 s 14756 10166 14756 10166 4 _0122_
rlabel metal1 s 16380 12342 16380 12342 4 _0123_
rlabel metal1 s 14168 11322 14168 11322 4 _0124_
rlabel metal2 s 14301 13362 14301 13362 4 _0125_
rlabel metal1 s 5060 17850 5060 17850 4 _0126_
rlabel metal2 s 6481 18802 6481 18802 4 _0127_
rlabel metal1 s 10089 18870 10089 18870 4 _0128_
rlabel metal1 s 6762 17306 6762 17306 4 _0129_
rlabel metal1 s 10365 15606 10365 15606 4 _0130_
rlabel metal1 s 8510 16660 8510 16660 4 _0131_
rlabel metal1 s 6435 15946 6435 15946 4 _0132_
rlabel metal2 s 6302 13192 6302 13192 4 _0133_
rlabel metal1 s 6490 12342 6490 12342 4 _0134_
rlabel metal2 s 4646 11492 4646 11492 4 _0135_
rlabel metal1 s 3905 12342 3905 12342 4 _0136_
rlabel metal1 s 6343 9418 6343 9418 4 _0137_
rlabel metal1 s 4600 10642 4600 10642 4 _0138_
rlabel metal2 s 4181 9010 4181 9010 4 _0139_
rlabel metal2 s 2433 10098 2433 10098 4 _0140_
rlabel metal1 s 3036 9622 3036 9622 4 _0141_
rlabel metal1 s 1794 10642 1794 10642 4 _0142_
rlabel metal1 s 2208 12206 2208 12206 4 _0143_
rlabel metal1 s 2944 13498 2944 13498 4 _0144_
rlabel metal2 s 1145 14518 1145 14518 4 _0145_
rlabel metal1 s 1794 15606 1794 15606 4 _0146_
rlabel metal1 s 3312 14382 3312 14382 4 _0147_
rlabel metal1 s 3726 15130 3726 15130 4 _0148_
rlabel metal1 s 6578 14314 6578 14314 4 _0149_
rlabel metal2 s 20010 24038 20010 24038 4 _0150_
rlabel metal2 s 20465 24718 20465 24718 4 _0151_
rlabel metal2 s 19821 26894 19821 26894 4 _0152_
rlabel metal1 s 19724 28594 19724 28594 4 _0153_
rlabel metal1 s 22770 30056 22770 30056 4 _0154_
rlabel metal1 s 19642 29274 19642 29274 4 _0155_
rlabel metal1 s 19637 30158 19637 30158 4 _0156_
rlabel metal1 s 22596 29682 22596 29682 4 _0157_
rlabel metal1 s 10299 11594 10299 11594 4 _0158_
rlabel metal1 s 5596 20298 5596 20298 4 _0159_
rlabel metal1 s 3956 20026 3956 20026 4 _0160_
rlabel metal1 s 3721 22474 3721 22474 4 _0161_
rlabel metal2 s 1242 22338 1242 22338 4 _0162_
rlabel metal2 s 3542 24038 3542 24038 4 _0163_
rlabel metal2 s 1145 23630 1145 23630 4 _0164_
rlabel metal2 s 1145 24650 1145 24650 4 _0165_
rlabel metal1 s 1334 26010 1334 26010 4 _0166_
rlabel metal1 s 3583 25738 3583 25738 4 _0167_
rlabel metal1 s 5244 25466 5244 25466 4 _0168_
rlabel metal1 s 6016 27506 6016 27506 4 _0169_
rlabel metal2 s 2525 27574 2525 27574 4 _0170_
rlabel metal1 s 2208 28186 2208 28186 4 _0171_
rlabel metal2 s 3629 30090 3629 30090 4 _0172_
rlabel metal1 s 6016 28594 6016 28594 4 _0173_
rlabel metal1 s 6240 30090 6240 30090 4 _0174_
rlabel metal2 s 4273 18802 4273 18802 4 _0175_
rlabel metal1 s 8418 11254 8418 11254 4 _0176_
rlabel metal1 s 7769 10098 7769 10098 4 _0177_
rlabel metal1 s 7539 8330 7539 8330 4 _0178_
rlabel metal2 s 9522 8194 9522 8194 4 _0179_
rlabel metal1 s 10304 10642 10304 10642 4 _0180_
rlabel metal2 s 21569 13362 21569 13362 4 _0181_
rlabel metal1 s 20792 13498 20792 13498 4 _0182_
rlabel metal1 s 21983 11662 21983 11662 4 _0183_
rlabel metal2 s 21528 12308 21528 12308 4 _0184_
rlabel metal2 s 11914 23256 11914 23256 4 _0185_
rlabel metal1 s 11484 22134 11484 22134 4 _0186_
rlabel metal1 s 10851 25738 10851 25738 4 _0187_
rlabel metal1 s 11868 25466 11868 25466 4 _0188_
rlabel metal1 s 11495 28662 11495 28662 4 _0189_
rlabel metal1 s 11040 27098 11040 27098 4 _0190_
rlabel metal1 s 12788 26554 12788 26554 4 _0191_
rlabel metal2 s 12742 28390 12742 28390 4 _0192_
rlabel metal1 s 6532 14994 6532 14994 4 _0193_
rlabel metal1 s 9522 2618 9522 2618 4 _0194_
rlabel metal1 s 9986 4046 9986 4046 4 _0195_
rlabel metal1 s 8836 6834 8836 6834 4 _0196_
rlabel metal2 s 6394 8194 6394 8194 4 _0197_
rlabel metal1 s 3036 7786 3036 7786 4 _0198_
rlabel metal2 s 5386 6902 5386 6902 4 _0199_
rlabel metal1 s 1288 6426 1288 6426 4 _0200_
rlabel metal1 s 2024 8466 2024 8466 4 _0201_
rlabel metal2 s 1886 16157 1886 16157 4 _0202_
rlabel metal1 s 17250 2074 17250 2074 4 _0203_
rlabel metal2 s 19366 4454 19366 4454 4 _0204_
rlabel metal1 s 19784 6154 19784 6154 4 _0205_
rlabel metal1 s 18450 7922 18450 7922 4 _0206_
rlabel metal1 s 13274 6902 13274 6902 4 _0207_
rlabel metal1 s 17070 7922 17070 7922 4 _0208_
rlabel metal1 s 12389 7242 12389 7242 4 _0209_
rlabel metal1 s 10963 5814 10963 5814 4 _0210_
rlabel metal4 s 1909 29716 1909 29716 4 _0211_
rlabel metal1 s 7452 2822 7452 2822 4 _0212_
rlabel metal1 s 3588 782 3588 782 4 _0213_
rlabel metal1 s 2438 1428 2438 1428 4 _0214_
rlabel metal1 s 4232 2346 4232 2346 4 _0215_
rlabel metal1 s 1288 1394 1288 1394 4 _0216_
rlabel metal1 s 1242 748 1242 748 4 _0217_
rlabel metal2 s 7038 1394 7038 1394 4 _0218_
rlabel metal2 s 6302 2176 6302 2176 4 _0219_
rlabel metal1 s 6808 2346 6808 2346 4 _0220_
rlabel metal1 s 5842 2278 5842 2278 4 _0221_
rlabel metal1 s 5474 3536 5474 3536 4 _0222_
rlabel metal1 s 4922 2618 4922 2618 4 _0223_
rlabel metal1 s 4692 782 4692 782 4 _0224_
rlabel metal1 s 4600 1870 4600 1870 4 _0225_
rlabel metal1 s 3588 1394 3588 1394 4 _0226_
rlabel metal1 s 7452 2958 7452 2958 4 _0227_
rlabel metal1 s 7314 4012 7314 4012 4 _0228_
rlabel metal1 s 6946 5100 6946 5100 4 _0229_
rlabel metal1 s 6026 5338 6026 5338 4 _0230_
rlabel metal1 s 5198 5338 5198 5338 4 _0231_
rlabel metal2 s 2990 5542 2990 5542 4 _0232_
rlabel metal1 s 1518 5100 1518 5100 4 _0233_
rlabel metal1 s 3358 3910 3358 3910 4 _0234_
rlabel metal1 s 17342 1462 17342 1462 4 _0235_
rlabel metal1 s 11638 1394 11638 1394 4 _0236_
rlabel metal2 s 10856 1870 10856 1870 4 _0237_
rlabel metal2 s 15042 2278 15042 2278 4 _0238_
rlabel metal2 s 9982 1394 9982 1394 4 _0239_
rlabel metal3 s 15778 3587 15778 3587 4 _0240_
rlabel metal1 s 16238 714 16238 714 4 _0241_
rlabel metal1 s 16146 1394 16146 1394 4 _0242_
rlabel metal1 s 14904 2550 14904 2550 4 _0243_
rlabel metal1 s 14628 2278 14628 2278 4 _0244_
rlabel metal1 s 14812 3570 14812 3570 4 _0245_
rlabel metal2 s 13754 1615 13754 1615 4 _0246_
rlabel metal1 s 12604 1394 12604 1394 4 _0247_
rlabel metal1 s 12650 782 12650 782 4 _0248_
rlabel metal2 s 12006 2074 12006 2074 4 _0249_
rlabel metal1 s 16514 2924 16514 2924 4 _0250_
rlabel metal1 s 16422 4012 16422 4012 4 _0251_
rlabel metal1 s 16192 3910 16192 3910 4 _0252_
rlabel metal1 s 15870 5100 15870 5100 4 _0253_
rlabel metal1 s 14444 4794 14444 4794 4 _0254_
rlabel metal1 s 12834 5338 12834 5338 4 _0255_
rlabel metal1 s 12374 4726 12374 4726 4 _0256_
rlabel metal1 s 12880 4182 12880 4182 4 _0257_
rlabel metal1 s 23782 2822 23782 2822 4 _0258_
rlabel metal1 s 20562 782 20562 782 4 _0259_
rlabel metal1 s 19550 1870 19550 1870 4 _0260_
rlabel metal1 s 22862 2414 22862 2414 4 _0261_
rlabel metal2 s 19090 782 19090 782 4 _0262_
rlabel metal2 s 19458 1394 19458 1394 4 _0263_
rlabel metal1 s 22724 3570 22724 3570 4 _0264_
rlabel metal1 s 23874 782 23874 782 4 _0265_
rlabel metal1 s 22632 2550 22632 2550 4 _0266_
rlabel metal1 s 22678 2618 22678 2618 4 _0267_
rlabel metal1 s 22724 4046 22724 4046 4 _0268_
rlabel metal1 s 22448 1462 22448 1462 4 _0269_
rlabel metal2 s 21574 1530 21574 1530 4 _0270_
rlabel metal1 s 21574 1428 21574 1428 4 _0271_
rlabel metal2 s 20470 2074 20470 2074 4 _0272_
rlabel metal1 s 24288 2958 24288 2958 4 _0273_
rlabel metal1 s 24058 3706 24058 3706 4 _0274_
rlabel metal1 s 24150 4658 24150 4658 4 _0275_
rlabel metal1 s 23598 5746 23598 5746 4 _0276_
rlabel metal2 s 22862 6052 22862 6052 4 _0277_
rlabel metal1 s 21850 6834 21850 6834 4 _0278_
rlabel metal1 s 21758 6154 21758 6154 4 _0279_
rlabel metal1 s 20792 4522 20792 4522 4 _0280_
rlabel metal1 s 15410 24922 15410 24922 4 _0281_
rlabel metal2 s 15732 20604 15732 20604 4 _0282_
rlabel metal1 s 15640 15538 15640 15538 4 _0283_
rlabel metal1 s 20654 23188 20654 23188 4 _0284_
rlabel metal1 s 16422 21522 16422 21522 4 _0285_
rlabel metal1 s 16376 21658 16376 21658 4 _0286_
rlabel metal1 s 16882 26418 16882 26418 4 _0287_
rlabel metal1 s 13386 24038 13386 24038 4 _0288_
rlabel metal1 s 14490 23698 14490 23698 4 _0289_
rlabel metal1 s 13716 22406 13716 22406 4 _0290_
rlabel metal2 s 14352 21828 14352 21828 4 _0291_
rlabel metal1 s 12834 24208 12834 24208 4 _0292_
rlabel metal2 s 14490 24242 14490 24242 4 _0293_
rlabel metal1 s 13110 24310 13110 24310 4 _0294_
rlabel metal1 s 13110 23732 13110 23732 4 _0295_
rlabel metal1 s 14122 24344 14122 24344 4 _0296_
rlabel metal1 s 14812 25194 14812 25194 4 _0297_
rlabel metal2 s 14950 25160 14950 25160 4 _0298_
rlabel metal1 s 15364 24718 15364 24718 4 _0299_
rlabel metal1 s 14996 29478 14996 29478 4 _0300_
rlabel metal1 s 14774 29818 14774 29818 4 _0301_
rlabel metal2 s 15318 30294 15318 30294 4 _0302_
rlabel metal1 s 16246 28730 16246 28730 4 _0303_
rlabel metal1 s 15456 29002 15456 29002 4 _0304_
rlabel metal2 s 16790 30294 16790 30294 4 _0305_
rlabel metal1 s 16798 27574 16798 27574 4 _0306_
rlabel metal1 s 17158 29036 17158 29036 4 _0307_
rlabel metal1 s 17710 29274 17710 29274 4 _0308_
rlabel metal1 s 16790 28458 16790 28458 4 _0309_
rlabel metal1 s 17572 28662 17572 28662 4 _0310_
rlabel metal1 s 18078 28730 18078 28730 4 _0311_
rlabel metal1 s 17020 26894 17020 26894 4 _0312_
rlabel metal2 s 18354 27472 18354 27472 4 _0313_
rlabel metal1 s 17848 27098 17848 27098 4 _0314_
rlabel metal2 s 17994 26758 17994 26758 4 _0315_
rlabel metal1 s 18998 26928 18998 26928 4 _0316_
rlabel metal1 s 18492 26010 18492 26010 4 _0317_
rlabel metal1 s 18124 26010 18124 26010 4 _0318_
rlabel metal1 s 18367 26554 18367 26554 4 _0319_
rlabel metal1 s 18722 25772 18722 25772 4 _0320_
rlabel metal2 s 23598 11492 23598 11492 4 _0321_
rlabel metal1 s 23138 11186 23138 11186 4 _0322_
rlabel metal2 s 23414 12551 23414 12551 4 _0323_
rlabel metal2 s 23598 12551 23598 12551 4 _0324_
rlabel metal1 s 23184 12954 23184 12954 4 _0325_
rlabel metal1 s 23184 11050 23184 11050 4 _0326_
rlabel metal1 s 24840 13906 24840 13906 4 _0327_
rlabel metal1 s 24104 13906 24104 13906 4 _0328_
rlabel metal1 s 24426 13498 24426 13498 4 _0329_
rlabel metal1 s 24196 13838 24196 13838 4 _0330_
rlabel metal1 s 24242 13974 24242 13974 4 _0331_
rlabel metal1 s 23046 13396 23046 13396 4 _0332_
rlabel metal1 s 22494 19686 22494 19686 4 _0333_
rlabel metal1 s 24196 14926 24196 14926 4 _0334_
rlabel metal1 s 23184 15470 23184 15470 4 _0335_
rlabel metal1 s 23092 15538 23092 15538 4 _0336_
rlabel metal1 s 22862 14552 22862 14552 4 _0337_
rlabel metal1 s 23506 17204 23506 17204 4 _0338_
rlabel metal1 s 22678 17136 22678 17136 4 _0339_
rlabel metal1 s 22954 16728 22954 16728 4 _0340_
rlabel metal2 s 23138 16694 23138 16694 4 _0341_
rlabel metal1 s 22862 16456 22862 16456 4 _0342_
rlabel metal1 s 22862 14450 22862 14450 4 _0343_
rlabel metal2 s 23138 18666 23138 18666 4 _0344_
rlabel metal2 s 22862 18768 22862 18768 4 _0345_
rlabel metal2 s 22586 19108 22586 19108 4 _0346_
rlabel metal1 s 22954 18224 22954 18224 4 _0347_
rlabel metal1 s 22540 18394 22540 18394 4 _0348_
rlabel metal1 s 23184 17850 23184 17850 4 _0349_
rlabel metal1 s 22494 18326 22494 18326 4 _0350_
rlabel metal1 s 22402 16626 22402 16626 4 _0351_
rlabel metal1 s 22586 16660 22586 16660 4 _0352_
rlabel metal1 s 22540 14450 22540 14450 4 _0353_
rlabel metal1 s 23230 13498 23230 13498 4 _0354_
rlabel metal1 s 22724 13294 22724 13294 4 _0355_
rlabel metal2 s 23322 17901 23322 17901 4 _0356_
rlabel metal1 s 20470 12784 20470 12784 4 _0357_
rlabel metal1 s 19964 12750 19964 12750 4 _0358_
rlabel metal1 s 24748 16762 24748 16762 4 _0359_
rlabel metal1 s 24196 12954 24196 12954 4 _0360_
rlabel metal1 s 25116 19278 25116 19278 4 _0361_
rlabel metal1 s 23644 18394 23644 18394 4 _0362_
rlabel metal1 s 23706 19210 23706 19210 4 _0363_
rlabel metal2 s 23690 19924 23690 19924 4 _0364_
rlabel metal1 s 25024 18666 25024 18666 4 _0365_
rlabel metal1 s 24840 18394 24840 18394 4 _0366_
rlabel metal1 s 25668 18802 25668 18802 4 _0367_
rlabel metal1 s 24058 16660 24058 16660 4 _0368_
rlabel metal1 s 25254 17714 25254 17714 4 _0369_
rlabel metal1 s 25668 17714 25668 17714 4 _0370_
rlabel metal1 s 24794 17306 24794 17306 4 _0371_
rlabel metal1 s 24288 16762 24288 16762 4 _0372_
rlabel metal1 s 25530 16626 25530 16626 4 _0373_
rlabel metal1 s 24242 16558 24242 16558 4 _0374_
rlabel metal1 s 24702 16456 24702 16456 4 _0375_
rlabel metal1 s 25346 16660 25346 16660 4 _0376_
rlabel metal1 s 24840 15130 24840 15130 4 _0377_
rlabel metal1 s 25040 14858 25040 14858 4 _0378_
rlabel metal1 s 25254 15130 25254 15130 4 _0379_
rlabel metal1 s 25622 14246 25622 14246 4 _0380_
rlabel metal1 s 25392 14790 25392 14790 4 _0381_
rlabel metal1 s 26036 14450 26036 14450 4 _0382_
rlabel metal1 s 24840 13362 24840 13362 4 _0383_
rlabel metal1 s 25438 14518 25438 14518 4 _0384_
rlabel metal1 s 26634 14416 26634 14416 4 _0385_
rlabel metal1 s 24242 12886 24242 12886 4 _0386_
rlabel metal1 s 24748 12682 24748 12682 4 _0387_
rlabel metal1 s 25484 12954 25484 12954 4 _0388_
rlabel metal1 s 24334 11696 24334 11696 4 _0389_
rlabel metal1 s 23966 23188 23966 23188 4 _0390_
rlabel metal1 s 24104 23290 24104 23290 4 _0391_
rlabel metal1 s 24978 22508 24978 22508 4 _0392_
rlabel metal1 s 24656 23630 24656 23630 4 _0393_
rlabel metal1 s 25438 21930 25438 21930 4 _0394_
rlabel metal1 s 23736 21454 23736 21454 4 _0395_
rlabel metal1 s 24610 21658 24610 21658 4 _0396_
rlabel metal1 s 25116 21658 25116 21658 4 _0397_
rlabel metal1 s 24426 20842 24426 20842 4 _0398_
rlabel metal1 s 25254 23222 25254 23222 4 _0399_
rlabel metal1 s 24702 23834 24702 23834 4 _0400_
rlabel metal1 s 23644 26282 23644 26282 4 _0401_
rlabel metal2 s 23506 26146 23506 26146 4 _0402_
rlabel metal1 s 23138 26418 23138 26418 4 _0403_
rlabel metal1 s 24150 26010 24150 26010 4 _0404_
rlabel metal1 s 23230 24208 23230 24208 4 _0405_
rlabel metal1 s 23000 24378 23000 24378 4 _0406_
rlabel metal1 s 22724 24786 22724 24786 4 _0407_
rlabel metal1 s 24012 24174 24012 24174 4 _0408_
rlabel metal1 s 23092 26554 23092 26554 4 _0409_
rlabel metal2 s 23138 25500 23138 25500 4 _0410_
rlabel metal2 s 24334 26928 24334 26928 4 _0411_
rlabel metal1 s 24564 27574 24564 27574 4 _0412_
rlabel metal1 s 24886 29750 24886 29750 4 _0413_
rlabel metal1 s 24380 29818 24380 29818 4 _0414_
rlabel metal2 s 25714 28118 25714 28118 4 _0415_
rlabel metal1 s 24288 29546 24288 29546 4 _0416_
rlabel metal2 s 24242 29750 24242 29750 4 _0417_
rlabel metal1 s 23828 30090 23828 30090 4 _0418_
rlabel metal1 s 23828 29206 23828 29206 4 _0419_
rlabel metal1 s 24058 30192 24058 30192 4 _0420_
rlabel metal1 s 24058 27914 24058 27914 4 _0421_
rlabel metal1 s 24334 27948 24334 27948 4 _0422_
rlabel metal2 s 24426 28458 24426 28458 4 _0423_
rlabel metal1 s 23736 24242 23736 24242 4 _0424_
rlabel metal1 s 24978 22950 24978 22950 4 _0425_
rlabel metal1 s 24146 24378 24146 24378 4 _0426_
rlabel metal1 s 23184 24854 23184 24854 4 _0427_
rlabel metal2 s 23046 24922 23046 24922 4 _0428_
rlabel metal1 s 24502 24650 24502 24650 4 _0429_
rlabel metal1 s 24334 24582 24334 24582 4 _0430_
rlabel metal2 s 23690 16320 23690 16320 4 _0431_
rlabel metal1 s 21252 15130 21252 15130 4 _0432_
rlabel metal2 s 21850 23460 21850 23460 4 _0433_
rlabel metal1 s 24518 25738 24518 25738 4 _0434_
rlabel metal1 s 25714 22100 25714 22100 4 _0435_
rlabel metal1 s 21804 26554 21804 26554 4 _0436_
rlabel metal1 s 21666 26010 21666 26010 4 _0437_
rlabel metal1 s 21114 26418 21114 26418 4 _0438_
rlabel metal1 s 22198 27506 22198 27506 4 _0439_
rlabel metal2 s 22402 27438 22402 27438 4 _0440_
rlabel metal2 s 21850 27710 21850 27710 4 _0441_
rlabel metal2 s 21666 28628 21666 28628 4 _0442_
rlabel metal1 s 21774 26826 21774 26826 4 _0443_
rlabel metal1 s 22402 27336 22402 27336 4 _0444_
rlabel metal2 s 22770 27336 22770 27336 4 _0445_
rlabel metal1 s 23046 27642 23046 27642 4 _0446_
rlabel metal1 s 25024 28186 25024 28186 4 _0447_
rlabel metal1 s 25622 28390 25622 28390 4 _0448_
rlabel metal1 s 24748 28594 24748 28594 4 _0449_
rlabel metal1 s 25606 26486 25606 26486 4 _0450_
rlabel metal1 s 25622 27642 25622 27642 4 _0451_
rlabel metal1 s 25760 28186 25760 28186 4 _0452_
rlabel metal1 s 25070 26350 25070 26350 4 _0453_
rlabel metal1 s 24794 26010 24794 26010 4 _0454_
rlabel metal1 s 26266 26486 26266 26486 4 _0455_
rlabel metal1 s 25162 24786 25162 24786 4 _0456_
rlabel metal1 s 26174 25126 26174 25126 4 _0457_
rlabel metal1 s 26910 25330 26910 25330 4 _0458_
rlabel metal1 s 25990 24208 25990 24208 4 _0459_
rlabel metal1 s 25484 24378 25484 24378 4 _0460_
rlabel metal1 s 25806 22984 25806 22984 4 _0461_
rlabel metal1 s 26818 20944 26818 20944 4 _0462_
rlabel metal2 s 25438 22746 25438 22746 4 _0463_
rlabel metal1 s 27048 20978 27048 20978 4 _0464_
rlabel metal1 s 26542 21862 26542 21862 4 _0465_
rlabel metal1 s 26834 22134 26834 22134 4 _0466_
rlabel metal1 s 26956 21930 26956 21930 4 _0467_
rlabel metal2 s 16606 9656 16606 9656 4 _0468_
rlabel metal1 s 15686 9554 15686 9554 4 _0469_
rlabel metal1 s 16100 10234 16100 10234 4 _0470_
rlabel metal1 s 15272 9486 15272 9486 4 _0471_
rlabel metal2 s 14950 10132 14950 10132 4 _0472_
rlabel metal1 s 16100 12410 16100 12410 4 _0473_
rlabel metal1 s 15778 12410 15778 12410 4 _0474_
rlabel metal2 s 15042 11458 15042 11458 4 _0475_
rlabel metal2 s 14306 11390 14306 11390 4 _0476_
rlabel metal1 s 14996 12750 14996 12750 4 _0477_
rlabel metal2 s 14582 13396 14582 13396 4 _0478_
rlabel metal1 s 5152 17714 5152 17714 4 _0479_
rlabel metal1 s 5520 17714 5520 17714 4 _0480_
rlabel metal1 s 10258 17204 10258 17204 4 _0481_
rlabel metal2 s 10258 16626 10258 16626 4 _0482_
rlabel metal2 s 10442 18972 10442 18972 4 _0483_
rlabel metal2 s 9154 17663 9154 17663 4 _0484_
rlabel metal2 s 8970 17952 8970 17952 4 _0485_
rlabel metal1 s 9706 17782 9706 17782 4 _0486_
rlabel metal2 s 10440 17102 10440 17102 4 _0487_
rlabel metal1 s 10442 16762 10442 16762 4 _0488_
rlabel metal1 s 7038 16660 7038 16660 4 _0489_
rlabel metal1 s 6992 16762 6992 16762 4 _0490_
rlabel metal1 s 6440 18190 6440 18190 4 _0491_
rlabel metal1 s 9016 18938 9016 18938 4 _0492_
rlabel metal1 s 9016 17850 9016 17850 4 _0493_
rlabel metal1 s 10534 18768 10534 18768 4 _0494_
rlabel metal1 s 7774 18326 7774 18326 4 _0495_
rlabel metal1 s 7866 18394 7866 18394 4 _0496_
rlabel metal2 s 7038 17578 7038 17578 4 _0497_
rlabel metal1 s 8556 16422 8556 16422 4 _0498_
rlabel metal1 s 8326 16625 8326 16625 4 _0499_
rlabel metal1 s 10810 15538 10810 15538 4 _0500_
rlabel metal1 s 8142 17136 8142 17136 4 _0501_
rlabel metal1 s 6118 14824 6118 14824 4 _0502_
rlabel metal1 s 6808 15674 6808 15674 4 _0503_
rlabel metal1 s 2622 13396 2622 13396 4 _0504_
rlabel metal1 s 2484 9690 2484 9690 4 _0505_
rlabel metal1 s 1058 13736 1058 13736 4 _0506_
rlabel metal1 s 1426 11764 1426 11764 4 _0507_
rlabel metal1 s 5842 12818 5842 12818 4 _0508_
rlabel metal1 s 6992 11118 6992 11118 4 _0509_
rlabel metal1 s 5106 11152 5106 11152 4 _0510_
rlabel metal1 s 4048 9622 4048 9622 4 _0511_
rlabel metal2 s 6854 10676 6854 10676 4 _0512_
rlabel metal1 s 5382 10540 5382 10540 4 _0513_
rlabel metal1 s 3404 9146 3404 9146 4 _0514_
rlabel metal1 s 2714 8058 2714 8058 4 _0515_
rlabel metal1 s 1610 15504 1610 15504 4 _0516_
rlabel metal2 s 2622 9044 2622 9044 4 _0517_
rlabel metal1 s 2024 11662 2024 11662 4 _0518_
rlabel metal1 s 1564 10710 1564 10710 4 _0519_
rlabel metal1 s 2024 12954 2024 12954 4 _0520_
rlabel metal1 s 1426 15572 1426 15572 4 _0521_
rlabel metal1 s 2116 15946 2116 15946 4 _0522_
rlabel metal2 s 2806 14246 2806 14246 4 _0523_
rlabel metal1 s 5888 14042 5888 14042 4 _0524_
rlabel metal1 s 3818 12410 3818 12410 4 _0525_
rlabel metal1 s 4094 13226 4094 13226 4 _0526_
rlabel metal1 s 6486 10234 6486 10234 4 _0527_
rlabel metal1 s 5658 13158 5658 13158 4 _0528_
rlabel metal1 s 4508 13430 4508 13430 4 _0529_
rlabel metal1 s 5750 13498 5750 13498 4 _0530_
rlabel metal1 s 7038 13872 7038 13872 4 _0531_
rlabel metal2 s 19458 30940 19458 30940 4 _0532_
rlabel metal1 s 19642 30872 19642 30872 4 _0533_
rlabel metal2 s 10166 12512 10166 12512 4 _0534_
rlabel metal1 s 9154 12818 9154 12818 4 _0535_
rlabel metal2 s 9246 12517 9246 12517 4 _0536_
rlabel metal2 s 9016 17170 9016 17170 4 _0537_
rlabel metal1 s 8694 11628 8694 11628 4 _0538_
rlabel metal1 s 9614 11220 9614 11220 4 _0539_
rlabel metal1 s 9982 11322 9982 11322 4 _0540_
rlabel metal1 s 10672 12274 10672 12274 4 _0541_
rlabel metal1 s 6532 22202 6532 22202 4 _0542_
rlabel metal1 s 6256 22610 6256 22610 4 _0543_
rlabel metal1 s 6394 21998 6394 21998 4 _0544_
rlabel metal2 s 6762 21964 6762 21964 4 _0545_
rlabel metal2 s 6302 22338 6302 22338 4 _0546_
rlabel metal1 s 7176 22474 7176 22474 4 _0547_
rlabel metal2 s 7498 20995 7498 20995 4 _0548_
rlabel metal1 s 7636 20910 7636 20910 4 _0549_
rlabel metal1 s 7084 21114 7084 21114 4 _0550_
rlabel metal1 s 7360 21590 7360 21590 4 _0551_
rlabel metal1 s 7636 22202 7636 22202 4 _0552_
rlabel metal1 s 6348 24582 6348 24582 4 _0553_
rlabel metal1 s 6670 24922 6670 24922 4 _0554_
rlabel metal2 s 7590 24242 7590 24242 4 _0555_
rlabel metal1 s 7130 24276 7130 24276 4 _0556_
rlabel metal1 s 7406 24208 7406 24208 4 _0557_
rlabel metal1 s 7682 23562 7682 23562 4 _0558_
rlabel metal2 s 8142 24004 8142 24004 4 _0559_
rlabel metal1 s 7358 24038 7358 24038 4 _0560_
rlabel metal1 s 7314 23664 7314 23664 4 _0561_
rlabel metal1 s 7130 23120 7130 23120 4 _0562_
rlabel metal1 s 7222 23222 7222 23222 4 _0563_
rlabel metal1 s 7544 23494 7544 23494 4 _0564_
rlabel metal2 s 6210 24463 6210 24463 4 _0565_
rlabel metal1 s 7314 23154 7314 23154 4 _0566_
rlabel metal1 s 8326 29274 8326 29274 4 _0567_
rlabel metal1 s 8464 29682 8464 29682 4 _0568_
rlabel metal1 s 7314 28593 7314 28593 4 _0569_
rlabel metal2 s 7769 29682 7769 29682 4 _0570_
rlabel metal1 s 7498 29682 7498 29682 4 _0571_
rlabel metal1 s 7590 28696 7590 28696 4 _0572_
rlabel metal1 s 6946 29002 6946 29002 4 _0573_
rlabel metal2 s 6946 29478 6946 29478 4 _0574_
rlabel metal1 s 7314 28458 7314 28458 4 _0575_
rlabel metal1 s 6670 27948 6670 27948 4 _0576_
rlabel metal1 s 7222 26010 7222 26010 4 _0577_
rlabel metal1 s 6900 26282 6900 26282 4 _0578_
rlabel metal1 s 9200 27302 9200 27302 4 _0579_
rlabel metal2 s 7774 27404 7774 27404 4 _0580_
rlabel metal2 s 8602 27370 8602 27370 4 _0581_
rlabel metal1 s 8188 27098 8188 27098 4 _0582_
rlabel metal1 s 7268 26962 7268 26962 4 _0583_
rlabel metal1 s 7268 27030 7268 27030 4 _0584_
rlabel metal1 s 7590 25874 7590 25874 4 _0585_
rlabel metal1 s 7130 26826 7130 26826 4 _0586_
rlabel metal1 s 7268 26418 7268 26418 4 _0587_
rlabel metal1 s 7636 23222 7636 23222 4 _0588_
rlabel metal1 s 7452 21998 7452 21998 4 _0589_
rlabel metal2 s 6762 27540 6762 27540 4 _0590_
rlabel metal1 s 7452 28730 7452 28730 4 _0591_
rlabel metal1 s 6992 28050 6992 28050 4 _0592_
rlabel metal1 s 6946 22066 6946 22066 4 _0593_
rlabel metal1 s 7602 21046 7602 21046 4 _0594_
rlabel metal1 s 7682 22474 7682 22474 4 _0595_
rlabel metal2 s 7498 22304 7498 22304 4 _0596_
rlabel metal1 s 5658 18768 5658 18768 4 _0597_
rlabel metal1 s 3358 19278 3358 19278 4 _0598_
rlabel metal1 s 4508 19958 4508 19958 4 _0599_
rlabel metal1 s 5290 20298 5290 20298 4 _0600_
rlabel metal1 s 4646 19686 4646 19686 4 _0601_
rlabel metal1 s 4730 20026 4730 20026 4 _0602_
rlabel metal1 s 4140 19890 4140 19890 4 _0603_
rlabel metal2 s 3534 23290 3534 23290 4 _0604_
rlabel metal1 s 4416 21862 4416 21862 4 _0605_
rlabel metal2 s 4094 22474 4094 22474 4 _0606_
rlabel metal1 s 2668 23290 2668 23290 4 _0607_
rlabel metal1 s 2484 22202 2484 22202 4 _0608_
rlabel metal1 s 1610 22066 1610 22066 4 _0609_
rlabel metal1 s 3414 24684 3414 24684 4 _0610_
rlabel metal2 s 3082 23222 3082 23222 4 _0611_
rlabel metal1 s 3312 23290 3312 23290 4 _0612_
rlabel metal1 s 2162 24310 2162 24310 4 _0613_
rlabel metal1 s 2668 24038 2668 24038 4 _0614_
rlabel metal1 s 1242 24174 1242 24174 4 _0615_
rlabel metal2 s 2484 25806 2484 25806 4 _0616_
rlabel metal1 s 2576 24922 2576 24922 4 _0617_
rlabel metal1 s 2346 24820 2346 24820 4 _0618_
rlabel metal2 s 2990 26112 2990 26112 4 _0619_
rlabel metal2 s 2622 26486 2622 26486 4 _0620_
rlabel metal1 s 1610 25840 1610 25840 4 _0621_
rlabel metal1 s 3174 25330 3174 25330 4 _0622_
rlabel metal1 s 3542 25398 3542 25398 4 _0623_
rlabel metal1 s 3680 25466 3680 25466 4 _0624_
rlabel metal1 s 5290 23290 5290 23290 4 _0625_
rlabel metal1 s 5244 24650 5244 24650 4 _0626_
rlabel metal1 s 5106 26350 5106 26350 4 _0627_
rlabel metal1 s 5704 26418 5704 26418 4 _0628_
rlabel metal1 s 4738 25364 4738 25364 4 _0629_
rlabel metal1 s 3542 28526 3542 28526 4 _0630_
rlabel metal1 s 5934 27030 5934 27030 4 _0631_
rlabel metal2 s 5290 27302 5290 27302 4 _0632_
rlabel metal1 s 4048 27302 4048 27302 4 _0633_
rlabel metal1 s 4370 27438 4370 27438 4 _0634_
rlabel metal1 s 3312 27642 3312 27642 4 _0635_
rlabel metal1 s 4278 28424 4278 28424 4 _0636_
rlabel metal2 s 4262 28662 4262 28662 4 _0637_
rlabel metal1 s 2438 28016 2438 28016 4 _0638_
rlabel metal1 s 4094 29206 4094 29206 4 _0639_
rlabel metal1 s 4278 29716 4278 29716 4 _0640_
rlabel metal1 s 4370 29274 4370 29274 4 _0641_
rlabel metal1 s 3818 29818 3818 29818 4 _0642_
rlabel metal1 s 4968 29274 4968 29274 4 _0643_
rlabel metal1 s 4738 29614 4738 29614 4 _0644_
rlabel metal1 s 5244 29070 5244 29070 4 _0645_
rlabel metal1 s 5796 29682 5796 29682 4 _0646_
rlabel metal1 s 6072 29818 6072 29818 4 _0647_
rlabel metal1 s 5290 18938 5290 18938 4 _0648_
rlabel metal1 s 7958 12614 7958 12614 4 _0649_
rlabel metal1 s 9016 11186 9016 11186 4 _0650_
rlabel metal1 s 8970 11254 8970 11254 4 _0651_
rlabel metal1 s 8924 11322 8924 11322 4 _0652_
rlabel metal1 s 10166 8942 10166 8942 4 _0653_
rlabel metal1 s 8372 9418 8372 9418 4 _0654_
rlabel metal2 s 8234 10132 8234 10132 4 _0655_
rlabel metal1 s 7958 8942 7958 8942 4 _0656_
rlabel metal2 s 9982 9180 9982 9180 4 _0657_
rlabel metal1 s 9338 9146 9338 9146 4 _0658_
rlabel metal1 s 9706 7990 9706 7990 4 _0659_
rlabel metal1 s 9476 10506 9476 10506 4 _0660_
rlabel metal1 s 20516 14450 20516 14450 4 _0661_
rlabel metal1 s 21114 12648 21114 12648 4 _0662_
rlabel metal1 s 12650 22644 12650 22644 4 _0663_
rlabel metal1 s 13064 26486 13064 26486 4 _0664_
rlabel metal1 s 9016 2278 9016 2278 4 _0665_
rlabel metal2 s 8891 2618 8891 2618 4 _0666_
rlabel metal1 s 9108 2482 9108 2482 4 _0667_
rlabel metal1 s 8602 4658 8602 4658 4 _0668_
rlabel metal1 s 8418 4692 8418 4692 4 _0669_
rlabel metal1 s 9062 4250 9062 4250 4 _0670_
rlabel metal1 s 8978 4794 8978 4794 4 _0671_
rlabel metal1 s 9384 4658 9384 4658 4 _0672_
rlabel metal1 s 8418 6222 8418 6222 4 _0673_
rlabel metal1 s 7682 6290 7682 6290 4 _0674_
rlabel metal2 s 8142 6120 8142 6120 4 _0675_
rlabel metal1 s 8372 6290 8372 6290 4 _0676_
rlabel metal1 s 8786 6426 8786 6426 4 _0677_
rlabel metal1 s 8096 6834 8096 6834 4 _0678_
rlabel metal1 s 6992 6834 6992 6834 4 _0679_
rlabel metal1 s 6394 6766 6394 6766 4 _0680_
rlabel metal1 s 6716 6698 6716 6698 4 _0681_
rlabel metal1 s 6992 6970 6992 6970 4 _0682_
rlabel metal1 s 6762 7514 6762 7514 4 _0683_
rlabel metal1 s 6624 7922 6624 7922 4 _0684_
rlabel metal1 s 4094 7276 4094 7276 4 _0685_
rlabel metal1 s 4830 7922 4830 7922 4 _0686_
rlabel metal1 s 4830 7514 4830 7514 4 _0687_
rlabel metal2 s 4186 7242 4186 7242 4 _0688_
rlabel metal1 s 2714 7990 2714 7990 4 _0689_
rlabel metal2 s 3634 7650 3634 7650 4 _0690_
rlabel metal1 s 4324 7514 4324 7514 4 _0691_
rlabel metal1 s 5382 7956 5382 7956 4 _0692_
rlabel metal1 s 5244 7310 5244 7310 4 _0693_
rlabel metal1 s 3496 6834 3496 6834 4 _0694_
rlabel metal1 s 3588 6698 3588 6698 4 _0695_
rlabel metal1 s 2070 7242 2070 7242 4 _0696_
rlabel metal2 s 2162 6868 2162 6868 4 _0697_
rlabel metal2 s 2530 6834 2530 6834 4 _0698_
rlabel metal1 s 2116 6970 2116 6970 4 _0699_
rlabel metal1 s 1656 6222 1656 6222 4 _0700_
rlabel metal1 s 1886 8602 1886 8602 4 _0701_
rlabel metal2 s 2438 8330 2438 8330 4 _0702_
rlabel metal1 s 2208 8398 2208 8398 4 _0703_
rlabel metal1 s 1426 10132 1426 10132 4 _0704_
rlabel metal1 s 17848 3502 17848 3502 4 _0705_
rlabel metal1 s 18446 2414 18446 2414 4 _0706_
rlabel metal2 s 17710 2346 17710 2346 4 _0707_
rlabel metal1 s 17802 4250 17802 4250 4 _0708_
rlabel metal1 s 17940 3910 17940 3910 4 _0709_
rlabel metal1 s 18676 4250 18676 4250 4 _0710_
rlabel metal2 s 18078 3808 18078 3808 4 _0711_
rlabel metal1 s 19136 4046 19136 4046 4 _0712_
rlabel metal2 s 18078 5270 18078 5270 4 _0713_
rlabel metal2 s 17986 6256 17986 6256 4 _0714_
rlabel metal1 s 18400 5882 18400 5882 4 _0715_
rlabel metal1 s 18354 6290 18354 6290 4 _0716_
rlabel metal1 s 18814 6358 18814 6358 4 _0717_
rlabel metal1 s 19320 6834 19320 6834 4 _0718_
rlabel metal1 s 17204 6222 17204 6222 4 _0719_
rlabel metal1 s 17204 5814 17204 5814 4 _0720_
rlabel metal1 s 16238 6290 16238 6290 4 _0721_
rlabel metal1 s 17066 6290 17066 6290 4 _0722_
rlabel metal2 s 17066 6834 17066 6834 4 _0723_
rlabel metal2 s 17618 7956 17618 7956 4 _0724_
rlabel metal1 s 13846 6188 13846 6188 4 _0725_
rlabel metal1 s 15502 5746 15502 5746 4 _0726_
rlabel metal1 s 14950 5780 14950 5780 4 _0727_
rlabel metal1 s 13156 6222 13156 6222 4 _0728_
rlabel metal1 s 13294 6426 13294 6426 4 _0729_
rlabel metal1 s 15180 7718 15180 7718 4 _0730_
rlabel metal1 s 15272 6970 15272 6970 4 _0731_
rlabel metal1 s 16146 7344 16146 7344 4 _0732_
rlabel metal1 s 16284 7514 16284 7514 4 _0733_
rlabel metal1 s 14720 6154 14720 6154 4 _0734_
rlabel metal1 s 14950 6800 14950 6800 4 _0735_
rlabel metal1 s 13754 7310 13754 7310 4 _0736_
rlabel metal1 s 11960 6630 11960 6630 4 _0737_
rlabel metal1 s 11546 6766 11546 6766 4 _0738_
rlabel metal2 s 12926 7684 12926 7684 4 _0739_
rlabel metal1 s 12742 7412 12742 7412 4 _0740_
rlabel metal2 s 11546 5304 11546 5304 4 _0741_
rlabel metal2 s 10258 5984 10258 5984 4 _0742_
rlabel metal1 s 11086 5338 11086 5338 4 _0743_
rlabel metal1 s 10396 6970 10396 6970 4 _0744_
rlabel metal1 s 11362 11084 11362 11084 4 _0745_
rlabel metal1 s 14122 9452 14122 9452 4 _0746_
rlabel metal2 s 14398 10778 14398 10778 4 _0747_
rlabel metal1 s 14950 14960 14950 14960 4 _0748_
rlabel metal1 s 14398 9996 14398 9996 4 _0749_
rlabel metal2 s 14490 3536 14490 3536 4 _0750_
rlabel metal1 s 14030 10132 14030 10132 4 _0751_
rlabel metal2 s 14306 10540 14306 10540 4 _0752_
rlabel metal2 s 14674 4131 14674 4131 4 _0753_
rlabel metal2 s 2622 4318 2622 4318 4 _0754_
rlabel metal1 s 19642 8976 19642 8976 4 _0755_
rlabel metal1 s 14490 7956 14490 7956 4 _0756_
rlabel metal2 s 14214 6800 14214 6800 4 _0757_
rlabel metal2 s 2254 4046 2254 4046 4 _0758_
rlabel metal1 s 19458 7956 19458 7956 4 _0759_
rlabel metal1 s 14812 8806 14812 8806 4 _0760_
rlabel metal1 s 12466 6222 12466 6222 4 _0761_
rlabel metal1 s 2024 2958 2024 2958 4 _0762_
rlabel metal1 s 3542 4590 3542 4590 4 _0763_
rlabel metal1 s 5014 4046 5014 4046 4 _0764_
rlabel metal1 s 6394 3536 6394 3536 4 _0765_
rlabel metal1 s 4784 4658 4784 4658 4 _0766_
rlabel metal1 s 5152 2482 5152 2482 4 _0767_
rlabel metal2 s 4370 2499 4370 2499 4 _0768_
rlabel metal1 s 4922 3604 4922 3604 4 _0769_
rlabel metal1 s 2162 2890 2162 2890 4 _0770_
rlabel metal1 s 6348 2618 6348 2618 4 _0771_
rlabel metal1 s 5382 4080 5382 4080 4 _0772_
rlabel metal1 s 5152 4658 5152 4658 4 _0773_
rlabel metal1 s 6256 3910 6256 3910 4 _0774_
rlabel metal1 s 7084 3570 7084 3570 4 _0775_
rlabel metal1 s 6486 2924 6486 2924 4 _0776_
rlabel metal1 s 6716 2618 6716 2618 4 _0777_
rlabel metal1 s 4554 3604 4554 3604 4 _0778_
rlabel metal1 s 4922 3400 4922 3400 4 _0779_
rlabel metal1 s 5888 3570 5888 3570 4 _0780_
rlabel metal1 s 6670 3706 6670 3706 4 _0781_
rlabel metal1 s 3634 2448 3634 2448 4 _0782_
rlabel metal1 s 6486 4250 6486 4250 4 _0783_
rlabel metal1 s 5796 4794 5796 4794 4 _0784_
rlabel metal2 s 5106 4420 5106 4420 4 _0785_
rlabel metal1 s 2438 5134 2438 5134 4 _0786_
rlabel metal1 s 3634 1870 3634 1870 4 _0787_
rlabel metal1 s 13156 10098 13156 10098 4 _0788_
rlabel metal2 s 13478 10370 13478 10370 4 _0789_
rlabel metal1 s 12742 4760 12742 4760 4 _0790_
rlabel metal2 s 13294 10268 13294 10268 4 _0791_
rlabel metal1 s 12926 9894 12926 9894 4 _0792_
rlabel metal1 s 11362 4726 11362 4726 4 _0793_
rlabel metal1 s 12926 9010 12926 9010 4 _0794_
rlabel metal1 s 12558 5780 12558 5780 4 _0795_
rlabel metal1 s 10626 4080 10626 4080 4 _0796_
rlabel metal1 s 12512 8466 12512 8466 4 _0797_
rlabel metal2 s 12374 6732 12374 6732 4 _0798_
rlabel metal1 s 12282 4624 12282 4624 4 _0799_
rlabel metal1 s 12236 4522 12236 4522 4 _0800_
rlabel metal1 s 13938 4012 13938 4012 4 _0801_
rlabel metal1 s 15640 3502 15640 3502 4 _0802_
rlabel metal1 s 13340 4658 13340 4658 4 _0803_
rlabel metal1 s 14490 2516 14490 2516 4 _0804_
rlabel metal1 s 12972 2482 12972 2482 4 _0805_
rlabel metal1 s 11454 3910 11454 3910 4 _0806_
rlabel metal1 s 10718 2992 10718 2992 4 _0807_
rlabel metal1 s 15410 2618 15410 2618 4 _0808_
rlabel metal1 s 14444 3570 14444 3570 4 _0809_
rlabel metal1 s 13708 4658 13708 4658 4 _0810_
rlabel metal2 s 14950 4182 14950 4182 4 _0811_
rlabel metal1 s 15962 3060 15962 3060 4 _0812_
rlabel metal1 s 14490 2992 14490 2992 4 _0813_
rlabel metal2 s 12788 2482 12788 2482 4 _0814_
rlabel metal1 s 11592 2482 11592 2482 4 _0815_
rlabel metal2 s 13846 3247 13846 3247 4 _0816_
rlabel metal1 s 14536 3638 14536 3638 4 _0817_
rlabel metal1 s 15410 3706 15410 3706 4 _0818_
rlabel metal1 s 14030 2482 14030 2482 4 _0819_
rlabel metal1 s 15640 3162 15640 3162 4 _0820_
rlabel metal1 s 15226 4794 15226 4794 4 _0821_
rlabel metal2 s 14214 3910 14214 3910 4 _0822_
rlabel metal2 s 12742 5338 12742 5338 4 _0823_
rlabel metal2 s 12190 2621 12190 2621 4 _0824_
rlabel metal1 s 19918 8942 19918 8942 4 _0825_
rlabel metal1 s 18630 9044 18630 9044 4 _0826_
rlabel metal1 s 20102 6834 20102 6834 4 _0827_
rlabel metal1 s 18906 10132 18906 10132 4 _0828_
rlabel metal1 s 21482 6800 21482 6800 4 _0829_
rlabel metal1 s 20148 5066 20148 5066 4 _0830_
rlabel metal1 s 20010 8976 20010 8976 4 _0831_
rlabel metal1 s 20930 6800 20930 6800 4 _0832_
rlabel metal1 s 19918 4692 19918 4692 4 _0833_
rlabel metal1 s 19090 7990 19090 7990 4 _0834_
rlabel metal1 s 20746 6868 20746 6868 4 _0835_
rlabel metal1 s 19090 2924 19090 2924 4 _0836_
rlabel metal1 s 20976 5134 20976 5134 4 _0837_
rlabel metal1 s 21666 4556 21666 4556 4 _0838_
rlabel metal1 s 23322 3638 23322 3638 4 _0839_
rlabel metal1 s 22034 5168 22034 5168 4 _0840_
rlabel metal1 s 22264 2482 22264 2482 4 _0841_
rlabel metal1 s 21804 2482 21804 2482 4 _0842_
rlabel metal1 s 19780 3570 19780 3570 4 _0843_
rlabel metal1 s 19780 2958 19780 2958 4 _0844_
rlabel metal1 s 23184 2618 23184 2618 4 _0845_
rlabel metal1 s 20838 4080 20838 4080 4 _0846_
rlabel metal1 s 22030 4658 22030 4658 4 _0847_
rlabel metal2 s 22954 4692 22954 4692 4 _0848_
rlabel metal1 s 23966 3536 23966 3536 4 _0849_
rlabel metal2 s 21482 3230 21482 3230 4 _0850_
rlabel metal1 s 22586 2448 22586 2448 4 _0851_
rlabel metal1 s 21252 2482 21252 2482 4 _0852_
rlabel metal1 s 21850 4114 21850 4114 4 _0853_
rlabel metal1 s 22678 3978 22678 3978 4 _0854_
rlabel metal1 s 23598 3570 23598 3570 4 _0855_
rlabel metal1 s 20746 2550 20746 2550 4 _0856_
rlabel metal1 s 23644 4658 23644 4658 4 _0857_
rlabel metal1 s 23184 5338 23184 5338 4 _0858_
rlabel metal1 s 22770 3366 22770 3366 4 _0859_
rlabel metal1 s 21206 6834 21206 6834 4 _0860_
rlabel metal1 s 20470 4046 20470 4046 4 _0861_
rlabel metal2 s 13156 29478 13156 29478 4 _0862_
rlabel metal1 s 14030 17714 14030 17714 4 _0863_
rlabel metal1 s 14176 17578 14176 17578 4 _0864_
rlabel metal1 s 8540 14518 8540 14518 4 _0865_
rlabel metal1 s 21160 15674 21160 15674 4 _0866_
rlabel metal1 s 15640 18190 15640 18190 4 _0867_
rlabel metal1 s 12742 21454 12742 21454 4 _0868_
rlabel metal1 s 17848 22066 17848 22066 4 _0869_
rlabel metal1 s 16882 17306 16882 17306 4 _0870_
rlabel metal1 s 13984 14926 13984 14926 4 _0871_
rlabel metal1 s 16422 22032 16422 22032 4 _0872_
rlabel metal1 s 17756 20366 17756 20366 4 _0873_
rlabel metal1 s 17894 20400 17894 20400 4 _0874_
rlabel metal1 s 18906 12682 18906 12682 4 _0875_
rlabel metal1 s 15088 12682 15088 12682 4 _0876_
rlabel metal2 s 20102 18836 20102 18836 4 _0877_
rlabel metal1 s 19688 18122 19688 18122 4 _0878_
rlabel metal1 s 14858 19686 14858 19686 4 _0879_
rlabel metal1 s 20792 16558 20792 16558 4 _0880_
rlabel metal1 s 20010 18394 20010 18394 4 _0881_
rlabel metal1 s 18262 17850 18262 17850 4 _0882_
rlabel metal1 s 17434 18394 17434 18394 4 _0883_
rlabel metal1 s 20884 18938 20884 18938 4 _0884_
rlabel metal1 s 20562 18802 20562 18802 4 _0885_
rlabel metal1 s 17843 19210 17843 19210 4 _0886_
rlabel metal1 s 17158 19482 17158 19482 4 _0887_
rlabel metal2 s 21666 17136 21666 17136 4 _0888_
rlabel metal2 s 21574 28645 21574 28645 4 _0889_
rlabel metal1 s 21022 16626 21022 16626 4 _0890_
rlabel metal1 s 19550 16762 19550 16762 4 _0891_
rlabel metal2 s 19090 17238 19090 17238 4 _0892_
rlabel metal1 s 19504 20026 19504 20026 4 _0893_
rlabel metal1 s 19734 20026 19734 20026 4 _0894_
rlabel metal1 s 21390 19890 21390 19890 4 _0895_
rlabel metal1 s 21160 20026 21160 20026 4 _0896_
rlabel metal1 s 14720 14926 14720 14926 4 _0897_
rlabel metal1 s 14536 19482 14536 19482 4 _0898_
rlabel metal1 s 16054 16626 16054 16626 4 _0899_
rlabel metal1 s 16422 16762 16422 16762 4 _0900_
rlabel metal1 s 14260 14450 14260 14450 4 _0901_
rlabel metal1 s 18032 12954 18032 12954 4 _0902_
rlabel metal1 s 17480 13838 17480 13838 4 _0903_
rlabel metal2 s 17986 15402 17986 15402 4 _0904_
rlabel metal1 s 17710 15130 17710 15130 4 _0905_
rlabel metal1 s 16882 14348 16882 14348 4 _0906_
rlabel metal1 s 15180 16014 15180 16014 4 _0907_
rlabel metal1 s 14582 16014 14582 16014 4 _0908_
rlabel metal2 s 16514 13872 16514 13872 4 _0909_
rlabel metal1 s 15824 13498 15824 13498 4 _0910_
rlabel metal1 s 18216 16762 18216 16762 4 _0911_
rlabel metal1 s 17664 17306 17664 17306 4 _0912_
rlabel metal1 s 19918 21522 19918 21522 4 _0913_
rlabel metal2 s 11270 19618 11270 19618 4 _0914_
rlabel metal1 s 13524 17714 13524 17714 4 _0915_
rlabel metal1 s 21620 21454 21620 21454 4 _0916_
rlabel metal1 s 21436 20978 21436 20978 4 _0917_
rlabel metal2 s 18722 4624 18722 4624 4 _0918_
rlabel metal1 s 25944 3162 25944 3162 4 _0919_
rlabel metal1 s 25660 2822 25660 2822 4 _0920_
rlabel metal1 s 25300 2958 25300 2958 4 _0921_
rlabel metal1 s 25760 4658 25760 4658 4 _0922_
rlabel metal1 s 26036 4658 26036 4658 4 _0923_
rlabel metal1 s 26726 4454 26726 4454 4 _0924_
rlabel metal1 s 25852 4726 25852 4726 4 _0925_
rlabel metal1 s 26956 4658 26956 4658 4 _0926_
rlabel metal1 s 2070 21522 2070 21522 4 _0927_
rlabel metal1 s 26036 5678 26036 5678 4 _0928_
rlabel metal1 s 25760 5610 25760 5610 4 _0929_
rlabel metal1 s 25852 6630 25852 6630 4 _0930_
rlabel metal1 s 26450 6290 26450 6290 4 _0931_
rlabel metal1 s 25852 6426 25852 6426 4 _0932_
rlabel metal1 s 24380 6834 24380 6834 4 _0933_
rlabel metal1 s 14076 14858 14076 14858 4 _0934_
rlabel metal1 s 25254 7310 25254 7310 4 _0935_
rlabel metal1 s 24748 7718 24748 7718 4 _0936_
rlabel metal1 s 25024 7922 25024 7922 4 _0937_
rlabel metal1 s 25208 7378 25208 7378 4 _0938_
rlabel metal1 s 25484 7514 25484 7514 4 _0939_
rlabel metal1 s 26634 7990 26634 7990 4 _0940_
rlabel metal1 s 22724 8058 22724 8058 4 _0941_
rlabel metal1 s 24058 8058 24058 8058 4 _0942_
rlabel metal1 s 23874 8466 23874 8466 4 _0943_
rlabel metal2 s 22862 8398 22862 8398 4 _0944_
rlabel metal1 s 22770 7990 22770 7990 4 _0945_
rlabel metal1 s 23598 9350 23598 9350 4 _0946_
rlabel metal1 s 24150 8602 24150 8602 4 _0947_
rlabel metal1 s 24518 9010 24518 9010 4 _0948_
rlabel metal1 s 24748 9146 24748 9146 4 _0949_
rlabel metal2 s 22954 8347 22954 8347 4 _0950_
rlabel metal1 s 22954 8908 22954 8908 4 _0951_
rlabel metal2 s 22034 8602 22034 8602 4 _0952_
rlabel metal1 s 21896 8058 21896 8058 4 _0953_
rlabel metal1 s 21850 8432 21850 8432 4 _0954_
rlabel metal1 s 21528 8262 21528 8262 4 _0955_
rlabel metal1 s 1426 18156 1426 18156 4 _0956_
rlabel metal1 s 21482 7956 21482 7956 4 _0957_
rlabel metal2 s 21114 10234 21114 10234 4 _0958_
rlabel metal1 s 21390 9452 21390 9452 4 _0959_
rlabel metal2 s 22218 10030 22218 10030 4 _0960_
rlabel metal1 s 20792 9622 20792 9622 4 _0961_
rlabel metal1 s 20930 15980 20930 15980 4 _0962_
rlabel metal1 s 12880 30158 12880 30158 4 _0963_
rlabel metal1 s 14030 29784 14030 29784 4 _0964_
rlabel metal1 s 13064 19822 13064 19822 4 _0965_
rlabel metal2 s 15226 20502 15226 20502 4 _0966_
rlabel metal1 s 15364 20978 15364 20978 4 _0967_
rlabel metal2 s 12650 20468 12650 20468 4 _0968_
rlabel metal1 s 12604 20978 12604 20978 4 _0969_
rlabel metal1 s 15870 18938 15870 18938 4 _0970_
rlabel metal1 s 15916 19482 15916 19482 4 _0971_
rlabel metal1 s 14076 18802 14076 18802 4 _0972_
rlabel metal1 s 14260 17102 14260 17102 4 _0973_
rlabel metal1 s 13432 29070 13432 29070 4 _0974_
rlabel metal1 s 1472 18938 1472 18938 4 _0975_
rlabel metal1 s 1518 21386 1518 21386 4 _0976_
rlabel metal1 s 2438 20366 2438 20366 4 _0977_
rlabel metal1 s 3128 20570 3128 20570 4 _0978_
rlabel metal1 s 2944 20502 2944 20502 4 _0979_
rlabel metal1 s 2300 18938 2300 18938 4 _0980_
rlabel metal1 s 2852 18394 2852 18394 4 _0981_
rlabel metal1 s 1656 17102 1656 17102 4 _0982_
rlabel metal1 s 2944 16490 2944 16490 4 _0983_
rlabel metal1 s 4278 17034 4278 17034 4 _0984_
rlabel metal1 s 4600 17306 4600 17306 4 _0985_
rlabel metal2 s 2714 16422 2714 16422 4 _0986_
rlabel metal1 s 8510 14416 8510 14416 4 _0987_
rlabel metal2 s 8694 15130 8694 15130 4 _0988_
rlabel metal2 s 9614 14382 9614 14382 4 _0989_
rlabel metal2 s 11914 13158 11914 13158 4 _0990_
rlabel metal1 s 14122 21046 14122 21046 4 _0991_
rlabel metal1 s 15640 21046 15640 21046 4 _0992_
rlabel metal2 s 9706 24888 9706 24888 4 _0993_
rlabel metal2 s 8418 24582 8418 24582 4 _0994_
rlabel metal1 s 17848 9690 17848 9690 4 _0995_
rlabel metal1 s 14812 17510 14812 17510 4 _0996_
rlabel metal1 s 17296 11730 17296 11730 4 _0997_
rlabel metal2 s 17618 9690 17618 9690 4 _0998_
rlabel metal1 s 19826 10234 19826 10234 4 _0999_
rlabel metal1 s 19320 10098 19320 10098 4 _1000_
rlabel metal1 s 19320 11866 19320 11866 4 _1001_
rlabel metal1 s 18170 11730 18170 11730 4 _1002_
rlabel metal1 s 17848 11322 17848 11322 4 _1003_
rlabel metal1 s 16560 11186 16560 11186 4 _1004_
rlabel metal2 s 19826 11798 19826 11798 4 _1005_
rlabel metal2 s 20838 12750 20838 12750 4 _1006_
rlabel metal2 s 14122 19618 14122 19618 4 _1007_
rlabel metal1 s 10626 19788 10626 19788 4 _1008_
rlabel metal1 s 10718 20026 10718 20026 4 _1009_
rlabel metal1 s 9154 21488 9154 21488 4 _1010_
rlabel metal2 s 12190 14212 12190 14212 4 _1011_
rlabel metal1 s 14490 15538 14490 15538 4 _1012_
rlabel metal1 s 12466 13430 12466 13430 4 _1013_
rlabel metal1 s 13616 15130 13616 15130 4 _1014_
rlabel metal1 s 12926 14960 12926 14960 4 _1015_
rlabel metal1 s 12190 11730 12190 11730 4 _1016_
rlabel metal2 s 12466 12308 12466 12308 4 _1017_
rlabel metal1 s 14122 12750 14122 12750 4 _1018_
rlabel metal1 s 13294 12750 13294 12750 4 _1019_
rlabel metal1 s 13248 11322 13248 11322 4 _1020_
rlabel metal1 s 12489 11526 12489 11526 4 _1021_
rlabel metal1 s 17342 25330 17342 25330 4 _1022_
rlabel metal2 s 16698 24956 16698 24956 4 _1023_
rlabel metal2 s 17526 24531 17526 24531 4 _1024_
rlabel metal1 s 16606 24820 16606 24820 4 _1025_
rlabel metal1 s 18768 25398 18768 25398 4 _1026_
rlabel metal1 s 18722 23562 18722 23562 4 _1027_
rlabel metal1 s 17710 24276 17710 24276 4 _1028_
rlabel metal1 s 18722 24378 18722 24378 4 _1029_
rlabel metal1 s 17894 24208 17894 24208 4 _1030_
rlabel metal1 s 16974 24616 16974 24616 4 _1031_
rlabel metal2 s 16422 25126 16422 25126 4 _1032_
rlabel metal2 s 13754 25534 13754 25534 4 _1033_
rlabel metal2 s 13662 25636 13662 25636 4 _1034_
rlabel metal1 s 14122 25466 14122 25466 4 _1035_
rlabel metal1 s 14766 25840 14766 25840 4 _1036_
rlabel metal1 s 15088 23494 15088 23494 4 _1037_
rlabel metal2 s 15226 23902 15226 23902 4 _1038_
rlabel metal1 s 15548 23630 15548 23630 4 _1039_
rlabel metal1 s 15824 23834 15824 23834 4 _1040_
rlabel metal1 s 14260 24922 14260 24922 4 _1041_
rlabel metal1 s 14858 25262 14858 25262 4 _1042_
rlabel metal1 s 15272 26010 15272 26010 4 _1043_
rlabel metal1 s 15640 27846 15640 27846 4 _1044_
rlabel metal1 s 15962 28186 15962 28186 4 _1045_
rlabel metal1 s 15686 26826 15686 26826 4 _1046_
rlabel metal1 s 14950 27948 14950 27948 4 _1047_
rlabel metal1 s 14674 28050 14674 28050 4 _1048_
rlabel metal1 s 15502 27302 15502 27302 4 _1049_
rlabel metal1 s 14536 27506 14536 27506 4 _1050_
rlabel metal1 s 15180 27370 15180 27370 4 _1051_
rlabel metal1 s 15594 26894 15594 26894 4 _1052_
rlabel metal1 s 15502 26452 15502 26452 4 _1053_
rlabel metal1 s 15778 26486 15778 26486 4 _1054_
rlabel metal1 s 15870 26486 15870 26486 4 _1055_
rlabel metal1 s 16146 24276 16146 24276 4 _1056_
rlabel metal1 s 16882 24310 16882 24310 4 _1057_
rlabel metal2 s 16326 24378 16326 24378 4 _1058_
rlabel metal1 s 15272 24106 15272 24106 4 _1059_
rlabel metal1 s 14904 24378 14904 24378 4 _1060_
rlabel metal2 s 15502 24888 15502 24888 4 _1061_
rlabel metal1 s 16008 24922 16008 24922 4 _1062_
rlabel metal1 s 4784 21658 4784 21658 4 _1063_
rlabel metal2 s 5568 23630 5568 23630 4 _1064_
rlabel metal1 s 4876 17578 4876 17578 4 _1065_
rlabel metal2 s 5198 26792 5198 26792 4 _1066_
rlabel metal1 s 5244 23834 5244 23834 4 _1067_
rlabel metal1 s 13432 30294 13432 30294 4 active
rlabel metal1 s 8878 3536 8878 3536 4 amp_A.pwm_out\[0\]
rlabel metal1 s 7912 4590 7912 4590 4 amp_A.pwm_out\[1\]
rlabel metal1 s 7728 5746 7728 5746 4 amp_A.pwm_out\[2\]
rlabel metal1 s 6762 6256 6762 6256 4 amp_A.pwm_out\[3\]
rlabel metal1 s 4002 6868 4002 6868 4 amp_A.pwm_out\[4\]
rlabel metal1 s 3726 6834 3726 6834 4 amp_A.pwm_out\[5\]
rlabel metal1 s 2438 6188 2438 6188 4 amp_A.pwm_out\[6\]
rlabel metal1 s 1748 10098 1748 10098 4 amp_A.pwm_out\[7\]
rlabel metal1 s 18400 2482 18400 2482 4 amp_B.pwm_out\[0\]
rlabel metal1 s 17250 4046 17250 4046 4 amp_B.pwm_out\[1\]
rlabel metal2 s 18170 5134 18170 5134 4 amp_B.pwm_out\[2\]
rlabel metal2 s 16606 6290 16606 6290 4 amp_B.pwm_out\[3\]
rlabel metal1 s 15226 6154 15226 6154 4 amp_B.pwm_out\[4\]
rlabel metal2 s 15042 6273 15042 6273 4 amp_B.pwm_out\[5\]
rlabel metal1 s 11362 6800 11362 6800 4 amp_B.pwm_out\[6\]
rlabel metal1 s 11178 5644 11178 5644 4 amp_B.pwm_out\[7\]
rlabel metal1 s 25990 2992 25990 2992 4 amp_C.pwm_out\[0\]
rlabel metal1 s 25024 4046 25024 4046 4 amp_C.pwm_out\[1\]
rlabel metal1 s 25300 6834 25300 6834 4 amp_C.pwm_out\[2\]
rlabel metal1 s 25530 7276 25530 7276 4 amp_C.pwm_out\[3\]
rlabel metal1 s 23644 7922 23644 7922 4 amp_C.pwm_out\[4\]
rlabel metal2 s 23138 7548 23138 7548 4 amp_C.pwm_out\[5\]
rlabel metal1 s 22034 7956 22034 7956 4 amp_C.pwm_out\[6\]
rlabel metal2 s 21022 7888 21022 7888 4 amp_C.pwm_out\[7\]
rlabel metal1 s 15640 9350 15640 9350 4 amplitude_A\[0\]
rlabel metal1 s 15686 9894 15686 9894 4 amplitude_A\[1\]
rlabel metal1 s 15778 12206 15778 12206 4 amplitude_A\[2\]
rlabel metal1 s 14996 11186 14996 11186 4 amplitude_A\[3\]
rlabel metal2 s 12604 9486 12604 9486 4 amplitude_B\[0\]
rlabel metal1 s 13662 15334 13662 15334 4 amplitude_B\[1\]
rlabel metal1 s 12926 12070 12926 12070 4 amplitude_B\[2\]
rlabel metal1 s 13800 13158 13800 13158 4 amplitude_B\[3\]
rlabel metal1 s 18308 9146 18308 9146 4 amplitude_C\[0\]
rlabel metal1 s 20056 9690 20056 9690 4 amplitude_C\[1\]
rlabel metal1 s 18998 11662 18998 11662 4 amplitude_C\[2\]
rlabel metal1 s 18308 11186 18308 11186 4 amplitude_C\[3\]
rlabel metal1 s 8832 30770 8832 30770 4 bc1
rlabel metal1 s 10672 30770 10672 30770 4 bdir
rlabel metal2 s 9522 874 9522 874 4 channel_A_dac_ctrl[0]
rlabel metal2 s 4002 568 4002 568 4 channel_A_dac_ctrl[10]
rlabel metal2 s 3450 551 3450 551 4 channel_A_dac_ctrl[11]
rlabel metal2 s 2898 1112 2898 1112 4 channel_A_dac_ctrl[12]
rlabel metal2 s 2346 874 2346 874 4 channel_A_dac_ctrl[13]
rlabel metal2 s 1794 568 1794 568 4 channel_A_dac_ctrl[14]
rlabel metal2 s 8970 908 8970 908 4 channel_A_dac_ctrl[1]
rlabel metal2 s 8418 568 8418 568 4 channel_A_dac_ctrl[2]
rlabel metal2 s 7866 1112 7866 1112 4 channel_A_dac_ctrl[3]
rlabel metal2 s 7286 0 7342 400 4 channel_A_dac_ctrl[4]
port 14 nsew
rlabel metal2 s 6762 415 6762 415 4 channel_A_dac_ctrl[5]
rlabel metal2 s 6210 908 6210 908 4 channel_A_dac_ctrl[6]
rlabel metal2 s 5658 568 5658 568 4 channel_A_dac_ctrl[7]
rlabel metal2 s 5106 1112 5106 1112 4 channel_A_dac_ctrl[8]
rlabel metal2 s 4554 874 4554 874 4 channel_A_dac_ctrl[9]
rlabel metal1 s 3588 29478 3588 29478 4 channel_A_pwm_out
rlabel metal2 s 17802 874 17802 874 4 channel_B_dac_ctrl[0]
rlabel metal2 s 12282 874 12282 874 4 channel_B_dac_ctrl[10]
rlabel metal2 s 11730 619 11730 619 4 channel_B_dac_ctrl[11]
rlabel metal2 s 11178 1044 11178 1044 4 channel_B_dac_ctrl[12]
rlabel metal2 s 10626 415 10626 415 4 channel_B_dac_ctrl[13]
rlabel metal2 s 10074 568 10074 568 4 channel_B_dac_ctrl[14]
rlabel metal2 s 17250 568 17250 568 4 channel_B_dac_ctrl[1]
rlabel metal2 s 16698 874 16698 874 4 channel_B_dac_ctrl[2]
rlabel metal2 s 16146 619 16146 619 4 channel_B_dac_ctrl[3]
rlabel metal2 s 15594 874 15594 874 4 channel_B_dac_ctrl[4]
rlabel metal2 s 15042 568 15042 568 4 channel_B_dac_ctrl[5]
rlabel metal2 s 14490 874 14490 874 4 channel_B_dac_ctrl[6]
rlabel metal2 s 13910 0 13966 400 4 channel_B_dac_ctrl[7]
port 33 nsew
rlabel metal2 s 13386 568 13386 568 4 channel_B_dac_ctrl[8]
rlabel metal2 s 12834 1112 12834 1112 4 channel_B_dac_ctrl[9]
rlabel metal1 s 2944 30294 2944 30294 4 channel_B_pwm_out
rlabel metal2 s 26082 1112 26082 1112 4 channel_C_dac_ctrl[0]
rlabel metal2 s 20534 0 20590 400 4 channel_C_dac_ctrl[10]
port 38 nsew
rlabel metal2 s 20010 1112 20010 1112 4 channel_C_dac_ctrl[11]
rlabel metal2 s 19458 415 19458 415 4 channel_C_dac_ctrl[12]
rlabel metal2 s 18906 415 18906 415 4 channel_C_dac_ctrl[13]
rlabel metal2 s 18354 874 18354 874 4 channel_C_dac_ctrl[14]
rlabel metal2 s 25530 874 25530 874 4 channel_C_dac_ctrl[1]
rlabel metal2 s 24978 568 24978 568 4 channel_C_dac_ctrl[2]
rlabel metal2 s 24426 1418 24426 1418 4 channel_C_dac_ctrl[3]
rlabel metal2 s 23874 415 23874 415 4 channel_C_dac_ctrl[4]
rlabel metal2 s 23322 1112 23322 1112 4 channel_C_dac_ctrl[5]
rlabel metal2 s 22770 551 22770 551 4 channel_C_dac_ctrl[6]
rlabel metal2 s 22218 568 22218 568 4 channel_C_dac_ctrl[7]
rlabel metal2 s 21666 415 21666 415 4 channel_C_dac_ctrl[8]
rlabel metal2 s 21114 619 21114 619 4 channel_C_dac_ctrl[9]
rlabel metal1 s 1196 30906 1196 30906 4 channel_C_pwm_out
rlabel metal3 s 16146 17051 16146 17051 4 clk
rlabel metal1 s 1656 19142 1656 19142 4 clk_counter\[0\]
rlabel metal1 s 2300 21454 2300 21454 4 clk_counter\[1\]
rlabel metal1 s 3496 21454 3496 21454 4 clk_counter\[2\]
rlabel metal1 s 2346 18666 2346 18666 4 clk_counter\[3\]
rlabel metal1 s 3772 17646 3772 17646 4 clk_counter\[4\]
rlabel metal1 s 3358 17578 3358 17578 4 clk_counter\[5\]
rlabel metal1 s 2438 17034 2438 17034 4 clk_counter\[6\]
rlabel metal2 s 14858 16456 14858 16456 4 clknet_0_clk
rlabel metal1 s 11408 18190 11408 18190 4 clknet_1_0__leaf_clk
rlabel metal1 s 18446 19210 18446 19210 4 clknet_1_1__leaf_clk
rlabel metal1 s 1380 14994 1380 14994 4 clknet_leaf_0_clk
rlabel metal1 s 19642 27574 19642 27574 4 clknet_leaf_10_clk
rlabel metal1 s 26680 25806 26680 25806 4 clknet_leaf_11_clk
rlabel metal1 s 26542 19278 26542 19278 4 clknet_leaf_12_clk
rlabel metal1 s 21942 20842 21942 20842 4 clknet_leaf_13_clk
rlabel metal1 s 18952 20366 18952 20366 4 clknet_leaf_14_clk
rlabel metal1 s 17572 15470 17572 15470 4 clknet_leaf_15_clk
rlabel metal1 s 26956 14926 26956 14926 4 clknet_leaf_16_clk
rlabel metal1 s 24012 6290 24012 6290 4 clknet_leaf_17_clk
rlabel metal1 s 17250 2550 17250 2550 4 clknet_leaf_18_clk
rlabel metal1 s 14030 13396 14030 13396 4 clknet_leaf_19_clk
rlabel metal1 s 9062 14892 9062 14892 4 clknet_leaf_1_clk
rlabel metal1 s 8004 8398 8004 8398 4 clknet_leaf_20_clk
rlabel metal1 s 874 11050 874 11050 4 clknet_leaf_21_clk
rlabel metal1 s 10074 20434 10074 20434 4 clknet_leaf_2_clk
rlabel metal1 s 7866 19278 7866 19278 4 clknet_leaf_3_clk
rlabel metal2 s 874 18496 874 18496 4 clknet_leaf_4_clk
rlabel metal1 s 2438 24616 2438 24616 4 clknet_leaf_5_clk
rlabel metal1 s 7774 28526 7774 28526 4 clknet_leaf_6_clk
rlabel metal2 s 12834 29376 12834 29376 4 clknet_leaf_7_clk
rlabel metal1 s 11638 21454 11638 21454 4 clknet_leaf_8_clk
rlabel metal1 s 13524 18190 13524 18190 4 clknet_leaf_9_clk
rlabel metal1 s 7544 30770 7544 30770 4 clock_select[0]
rlabel metal1 s 5980 30770 5980 30770 4 clock_select[1]
rlabel metal1 s 21804 30770 21804 30770 4 data[0]
rlabel metal1 s 20654 30158 20654 30158 4 data[1]
rlabel metal1 s 20010 30736 20010 30736 4 data[2]
rlabel metal1 s 17756 30838 17756 30838 4 data[3]
rlabel metal1 s 16192 30770 16192 30770 4 data[4]
rlabel metal1 s 14720 30770 14720 30770 4 data[5]
rlabel metal1 s 13754 30770 13754 30770 4 data[6]
rlabel metal1 s 11868 30770 11868 30770 4 data[7]
rlabel metal1 s 26588 30770 26588 30770 4 ena
rlabel metal1 s 14168 9010 14168 9010 4 envelope_A
rlabel metal1 s 13018 10608 13018 10608 4 envelope_B
rlabel metal1 s 19642 11220 19642 11220 4 envelope_C
rlabel metal1 s 8326 15130 8326 15130 4 envelope_generator.alternate
rlabel metal1 s 11224 13294 11224 13294 4 envelope_generator.attack
rlabel metal1 s 10212 13498 10212 13498 4 envelope_generator.continue_
rlabel metal2 s 9522 9214 9522 9214 4 envelope_generator.envelope_counter\[0\]
rlabel metal1 s 10580 9690 10580 9690 4 envelope_generator.envelope_counter\[1\]
rlabel metal1 s 9246 9418 9246 9418 4 envelope_generator.envelope_counter\[2\]
rlabel metal1 s 10534 10574 10534 10574 4 envelope_generator.envelope_counter\[3\]
rlabel metal1 s 8648 14586 8648 14586 4 envelope_generator.hold
rlabel metal1 s 11224 11186 11224 11186 4 envelope_generator.invert_output
rlabel metal1 s 8096 20570 8096 20570 4 envelope_generator.period\[0\]
rlabel metal1 s 8924 27438 8924 27438 4 envelope_generator.period\[10\]
rlabel metal1 s 11224 28118 11224 28118 4 envelope_generator.period\[11\]
rlabel metal1 s 9338 28730 9338 28730 4 envelope_generator.period\[12\]
rlabel metal1 s 11040 29818 11040 29818 4 envelope_generator.period\[13\]
rlabel metal1 s 9890 30022 9890 30022 4 envelope_generator.period\[14\]
rlabel metal1 s 8694 30022 8694 30022 4 envelope_generator.period\[15\]
rlabel metal1 s 7452 19686 7452 19686 4 envelope_generator.period\[1\]
rlabel metal1 s 8096 21862 8096 21862 4 envelope_generator.period\[2\]
rlabel metal1 s 6532 21658 6532 21658 4 envelope_generator.period\[3\]
rlabel metal1 s 8234 23698 8234 23698 4 envelope_generator.period\[4\]
rlabel metal1 s 11454 24174 11454 24174 4 envelope_generator.period\[5\]
rlabel metal1 s 9890 24378 9890 24378 4 envelope_generator.period\[6\]
rlabel metal1 s 8740 24922 8740 24922 4 envelope_generator.period\[7\]
rlabel metal1 s 9614 25466 9614 25466 4 envelope_generator.period\[8\]
rlabel metal1 s 9384 25670 9384 25670 4 envelope_generator.period\[9\]
rlabel metal1 s 6118 17306 6118 17306 4 envelope_generator.signal_edge.previous_signal_state_0
rlabel metal1 s 5750 18598 5750 18598 4 envelope_generator.signal_edge.signal
rlabel metal1 s 9706 11764 9706 11764 4 envelope_generator.stop
rlabel metal1 s 5290 21114 5290 21114 4 envelope_generator.tone.counter\[0\]
rlabel metal1 s 7820 27506 7820 27506 4 envelope_generator.tone.counter\[10\]
rlabel metal2 s 8050 27744 8050 27744 4 envelope_generator.tone.counter\[11\]
rlabel metal2 s 6670 28900 6670 28900 4 envelope_generator.tone.counter\[12\]
rlabel metal1 s 4784 28934 4784 28934 4 envelope_generator.tone.counter\[13\]
rlabel metal1 s 4600 29682 4600 29682 4 envelope_generator.tone.counter\[14\]
rlabel metal1 s 7176 30022 7176 30022 4 envelope_generator.tone.counter\[15\]
rlabel metal1 s 6670 20842 6670 20842 4 envelope_generator.tone.counter\[1\]
rlabel metal1 s 5704 22066 5704 22066 4 envelope_generator.tone.counter\[2\]
rlabel metal2 s 2254 22916 2254 22916 4 envelope_generator.tone.counter\[3\]
rlabel metal1 s 8142 24242 8142 24242 4 envelope_generator.tone.counter\[4\]
rlabel metal1 s 4922 24276 4922 24276 4 envelope_generator.tone.counter\[5\]
rlabel metal1 s 2346 24922 2346 24922 4 envelope_generator.tone.counter\[6\]
rlabel metal2 s 2346 26554 2346 26554 4 envelope_generator.tone.counter\[7\]
rlabel metal2 s 3358 26078 3358 26078 4 envelope_generator.tone.counter\[8\]
rlabel metal1 s 6072 25670 6072 25670 4 envelope_generator.tone.counter\[9\]
rlabel metal1 s 15088 20230 15088 20230 4 latched_register\[0\]
rlabel metal1 s 13156 20230 13156 20230 4 latched_register\[1\]
rlabel metal1 s 16560 18938 16560 18938 4 latched_register\[2\]
rlabel metal1 s 14490 18938 14490 18938 4 latched_register\[3\]
rlabel metal2 s 12466 30226 12466 30226 4 net1
rlabel metal1 s 17480 17034 17480 17034 4 net10
rlabel metal1 s 9522 27642 9522 27642 4 net100
rlabel metal1 s 19504 25330 19504 25330 4 net101
rlabel metal1 s 9982 19890 9982 19890 4 net102
rlabel metal1 s 12328 29070 12328 29070 4 net103
rlabel metal1 s 20930 12784 20930 12784 4 net104
rlabel metal1 s 8326 17748 8326 17748 4 net105
rlabel metal2 s 9062 16898 9062 16898 4 net106
rlabel metal1 s 8326 27540 8326 27540 4 net107
rlabel metal1 s 13386 17748 13386 17748 4 net108
rlabel metal1 s 21850 14484 21850 14484 4 net109
rlabel metal1 s 19596 19890 19596 19890 4 net11
rlabel metal1 s 21160 25330 21160 25330 4 net110
rlabel metal1 s 20792 27506 20792 27506 4 net111
rlabel metal2 s 10166 22678 10166 22678 4 net112
rlabel metal1 s 9522 21454 9522 21454 4 net113
rlabel metal1 s 11868 26418 11868 26418 4 net114
rlabel metal1 s 10258 27574 10258 27574 4 net115
rlabel metal1 s 9660 26418 9660 26418 4 net116
rlabel metal1 s 8602 26384 8602 26384 4 net117
rlabel metal2 s 11546 27370 11546 27370 4 net118
rlabel metal1 s 10074 29580 10074 29580 4 net119
rlabel metal1 s 21482 19822 21482 19822 4 net12
rlabel metal1 s 10718 24378 10718 24378 4 net120
rlabel metal1 s 12282 24310 12282 24310 4 net121
rlabel metal1 s 23322 30192 23322 30192 4 net122
rlabel metal1 s 13202 26452 13202 26452 4 net123
rlabel metal1 s 18446 22066 18446 22066 4 net124
rlabel metal1 s 9522 30736 9522 30736 4 net125
rlabel metal1 s 23276 12410 23276 12410 4 net126
rlabel metal1 s 3128 16626 3128 16626 4 net127
rlabel metal1 s 21390 13362 21390 13362 4 net128
rlabel metal1 s 17802 22576 17802 22576 4 net129
rlabel metal1 s 20930 30124 20930 30124 4 net13
rlabel metal1 s 17986 29036 17986 29036 4 net130
rlabel metal1 s 21298 22644 21298 22644 4 net131
rlabel metal1 s 6440 13770 6440 13770 4 net132
rlabel metal2 s 5938 13838 5938 13838 4 net133
rlabel metal1 s 18998 29104 18998 29104 4 net134
rlabel metal1 s 9844 10778 9844 10778 4 net135
rlabel metal1 s 10687 10166 10687 10166 4 net136
rlabel metal1 s 1472 21318 1472 21318 4 net137
rlabel metal2 s 1145 20366 1145 20366 4 net138
rlabel metal1 s 20884 22066 20884 22066 4 net139
rlabel metal1 s 17664 17102 17664 17102 4 net14
rlabel metal1 s 19826 30804 19826 30804 4 net140
rlabel metal1 s 9338 29070 9338 29070 4 net141
rlabel metal1 s 17572 20366 17572 20366 4 net142
rlabel metal1 s 2530 11526 2530 11526 4 net143
rlabel metal1 s 1334 10778 1334 10778 4 net144
rlabel metal1 s 1886 12308 1886 12308 4 net145
rlabel metal2 s 2810 12682 2810 12682 4 net146
rlabel metal1 s 2070 16048 2070 16048 4 net147
rlabel metal1 s 2203 14926 2203 14926 4 net148
rlabel metal1 s 9338 24242 9338 24242 4 net149
rlabel metal2 s 25346 1394 25346 1394 4 net15
rlabel metal1 s 6670 11254 6670 11254 4 net150
rlabel metal1 s 5458 11594 5458 11594 4 net151
rlabel metal1 s 7176 12682 7176 12682 4 net152
rlabel metal1 s 13294 28016 13294 28016 4 net153
rlabel metal1 s 13018 23154 13018 23154 4 net154
rlabel metal1 s 7038 10710 7038 10710 4 net155
rlabel metal2 s 4825 9486 4825 9486 4 net156
rlabel metal1 s 3036 9486 3036 9486 4 net157
rlabel metal1 s 6486 15572 6486 15572 4 net158
rlabel metal1 s 3542 14450 3542 14450 4 net159
rlabel metal1 s 24978 986 24978 986 4 net16
rlabel metal2 s 4374 13838 4374 13838 4 net160
rlabel metal1 s 2714 13328 2714 13328 4 net161
rlabel metal1 s 2085 13430 2085 13430 4 net162
rlabel metal1 s 1104 15538 1104 15538 4 net163
rlabel metal1 s 3634 14960 3634 14960 4 net164
rlabel metal1 s 2392 10438 2392 10438 4 net165
rlabel metal1 s 3680 9690 3680 9690 4 net166
rlabel metal2 s 6486 9622 6486 9622 4 net167
rlabel metal1 s 20930 23630 20930 23630 4 net168
rlabel metal1 s 4278 12716 4278 12716 4 net169
rlabel metal1 s 23828 850 23828 850 4 net17
rlabel metal1 s 23690 30702 23690 30702 4 net170
rlabel metal1 s 5704 25330 5704 25330 4 net171
rlabel metal1 s 25254 24752 25254 24752 4 net172
rlabel metal1 s 3220 18190 3220 18190 4 net173
rlabel metal1 s 2070 17850 2070 17850 4 net174
rlabel metal1 s 17020 27506 17020 27506 4 net175
rlabel metal1 s 6026 12784 6026 12784 4 net176
rlabel metal2 s 24794 12517 24794 12517 4 net177
rlabel metal1 s 20148 12614 20148 12614 4 net178
rlabel metal1 s 10626 12750 10626 12750 4 net179
rlabel metal2 s 23322 2587 23322 2587 4 net18
rlabel metal1 s 16008 16014 16008 16014 4 net180
rlabel metal1 s 20746 10608 20746 10608 4 net181
rlabel metal1 s 21804 14926 21804 14926 4 net182
rlabel metal1 s 24702 19244 24702 19244 4 net183
rlabel metal1 s 8832 11866 8832 11866 4 net184
rlabel metal2 s 7774 11458 7774 11458 4 net185
rlabel metal1 s 1288 9146 1288 9146 4 net186
rlabel metal1 s 15640 21454 15640 21454 4 net187
rlabel metal2 s 22034 23375 22034 23375 4 net188
rlabel metal1 s 8050 15368 8050 15368 4 net189
rlabel metal1 s 23460 986 23460 986 4 net19
rlabel metal1 s 11592 12682 11592 12682 4 net190
rlabel metal1 s 6532 19890 6532 19890 4 net191
rlabel metal1 s 10166 14280 10166 14280 4 net192
rlabel metal1 s 12650 30770 12650 30770 4 net2
rlabel metal1 s 22678 986 22678 986 4 net20
rlabel metal2 s 22494 1156 22494 1156 4 net21
rlabel metal1 s 21298 918 21298 918 4 net22
rlabel metal1 s 21390 1394 21390 1394 4 net23
rlabel metal1 s 20194 2006 20194 2006 4 net24
rlabel metal1 s 21068 850 21068 850 4 net25
rlabel metal1 s 18952 1870 18952 1870 4 net26
rlabel metal1 s 19136 986 19136 986 4 net27
rlabel metal1 s 18492 850 18492 850 4 net28
rlabel metal2 s 17894 1088 17894 1088 4 net29
rlabel metal1 s 5842 30192 5842 30192 4 net3
rlabel metal1 s 23966 3094 23966 3094 4 net30
rlabel metal1 s 23874 4114 23874 4114 4 net31
rlabel metal1 s 24058 4522 24058 4522 4 net32
rlabel metal2 s 23506 5950 23506 5950 4 net33
rlabel metal1 s 22586 5814 22586 5814 4 net34
rlabel metal2 s 21666 7072 21666 7072 4 net35
rlabel metal1 s 21252 5746 21252 5746 4 net36
rlabel metal1 s 20378 6358 20378 6358 4 net37
rlabel metal2 s 17342 1632 17342 1632 4 net38
rlabel metal1 s 16330 782 16330 782 4 net39
rlabel metal1 s 5842 30362 5842 30362 4 net4
rlabel metal1 s 15962 986 15962 986 4 net40
rlabel metal1 s 15180 1870 15180 1870 4 net41
rlabel metal2 s 14674 1632 14674 1632 4 net42
rlabel metal1 s 14122 884 14122 884 4 net43
rlabel metal1 s 13524 986 13524 986 4 net44
rlabel metal1 s 12926 1428 12926 1428 4 net45
rlabel metal2 s 13202 1428 13202 1428 4 net46
rlabel metal2 s 11730 1428 11730 1428 4 net47
rlabel metal1 s 11178 986 11178 986 4 net48
rlabel metal1 s 10488 986 10488 986 4 net49
rlabel metal1 s 19366 18224 19366 18224 4 net5
rlabel metal1 s 10442 1972 10442 1972 4 net50
rlabel metal1 s 9568 1326 9568 1326 4 net51
rlabel metal2 s 9246 1360 9246 1360 4 net52
rlabel metal2 s 16238 2720 16238 2720 4 net53
rlabel metal1 s 16100 4046 16100 4046 4 net54
rlabel metal1 s 16146 4590 16146 4590 4 net55
rlabel metal2 s 15594 5338 15594 5338 4 net56
rlabel metal2 s 14214 5372 14214 5372 4 net57
rlabel metal2 s 13018 5508 13018 5508 4 net58
rlabel metal1 s 12190 5134 12190 5134 4 net59
rlabel metal1 s 18400 18190 18400 18190 4 net6
rlabel metal1 s 10810 4726 10810 4726 4 net60
rlabel metal1 s 8234 986 8234 986 4 net61
rlabel metal1 s 6854 1360 6854 1360 4 net62
rlabel metal1 s 6946 850 6946 850 4 net63
rlabel metal1 s 6762 2006 6762 2006 4 net64
rlabel metal1 s 5934 918 5934 918 4 net65
rlabel metal1 s 5796 1394 5796 1394 4 net66
rlabel metal1 s 4554 1428 4554 1428 4 net67
rlabel metal1 s 4324 850 4324 850 4 net68
rlabel metal1 s 4094 2006 4094 2006 4 net69
rlabel metal1 s 20424 19278 20424 19278 4 net7
rlabel metal2 s 3358 1598 3358 1598 4 net70
rlabel metal1 s 3174 782 3174 782 4 net71
rlabel metal1 s 2208 986 2208 986 4 net72
rlabel metal1 s 1840 1870 1840 1870 4 net73
rlabel metal1 s 1058 1394 1058 1394 4 net74
rlabel metal2 s 966 1360 966 1360 4 net75
rlabel metal1 s 7222 3094 7222 3094 4 net76
rlabel metal2 s 7038 4250 7038 4250 4 net77
rlabel metal1 s 6670 5270 6670 5270 4 net78
rlabel metal1 s 5842 5814 5842 5814 4 net79
rlabel metal1 s 17710 19278 17710 19278 4 net8
rlabel metal1 s 5566 5780 5566 5780 4 net80
rlabel metal1 s 2714 5814 2714 5814 4 net81
rlabel metal2 s 1242 5338 1242 5338 4 net82
rlabel metal1 s 1196 4658 1196 4658 4 net83
rlabel metal1 s 11868 19278 11868 19278 4 net84
rlabel metal1 s 9614 19210 9614 19210 4 net85
rlabel metal1 s 8694 19924 8694 19924 4 net86
rlabel metal2 s 13570 25568 13570 25568 4 net87
rlabel metal1 s 24932 22066 24932 22066 4 net88
rlabel metal1 s 21206 21488 21206 21488 4 net89
rlabel metal1 s 16330 30362 16330 30362 4 net9
rlabel metal1 s 25852 11186 25852 11186 4 net90
rlabel metal1 s 23858 11254 23858 11254 4 net91
rlabel metal2 s 5014 18462 5014 18462 4 net92
rlabel metal1 s 18446 22576 18446 22576 4 net93
rlabel metal1 s 11684 19890 11684 19890 4 net94
rlabel metal1 s 13432 30158 13432 30158 4 net95
rlabel metal1 s 8510 23664 8510 23664 4 net96
rlabel metal1 s 11776 16014 11776 16014 4 net97
rlabel metal1 s 11822 23120 11822 23120 4 net98
rlabel metal1 s 21298 21012 21298 21012 4 net99
rlabel metal1 s 15456 16626 15456 16626 4 noise_disable_A
rlabel metal1 s 16836 14450 16836 14450 4 noise_disable_B
rlabel metal1 s 19090 16626 19090 16626 4 noise_disable_C
rlabel metal1 s 7314 13294 7314 13294 4 noise_generator.lfsr\[0\]
rlabel metal1 s 1518 12614 1518 12614 4 noise_generator.lfsr\[10\]
rlabel metal1 s 1058 13158 1058 13158 4 noise_generator.lfsr\[11\]
rlabel metal1 s 2070 12682 2070 12682 4 noise_generator.lfsr\[12\]
rlabel metal1 s 3266 14790 3266 14790 4 noise_generator.lfsr\[13\]
rlabel metal1 s 1242 12206 1242 12206 4 noise_generator.lfsr\[14\]
rlabel metal1 s 2622 13872 2622 13872 4 noise_generator.lfsr\[15\]
rlabel metal2 s 4830 13600 4830 13600 4 noise_generator.lfsr\[16\]
rlabel metal1 s 6532 12070 6532 12070 4 noise_generator.lfsr\[1\]
rlabel metal2 s 6578 11356 6578 11356 4 noise_generator.lfsr\[2\]
rlabel metal1 s 5060 12750 5060 12750 4 noise_generator.lfsr\[3\]
rlabel metal1 s 6992 10098 6992 10098 4 noise_generator.lfsr\[4\]
rlabel metal2 s 5842 10438 5842 10438 4 noise_generator.lfsr\[5\]
rlabel metal1 s 6256 10030 6256 10030 4 noise_generator.lfsr\[6\]
rlabel metal1 s 4692 9894 4692 9894 4 noise_generator.lfsr\[7\]
rlabel metal1 s 5106 11050 5106 11050 4 noise_generator.lfsr\[8\]
rlabel metal1 s 2944 11730 2944 11730 4 noise_generator.lfsr\[9\]
rlabel metal1 s 11040 19278 11040 19278 4 noise_generator.period\[0\]
rlabel metal2 s 12558 19346 12558 19346 4 noise_generator.period\[1\]
rlabel metal1 s 10534 18258 10534 18258 4 noise_generator.period\[2\]
rlabel metal1 s 11592 17102 11592 17102 4 noise_generator.period\[3\]
rlabel metal1 s 10902 17136 10902 17136 4 noise_generator.period\[4\]
rlabel metal1 s 6256 14858 6256 14858 4 noise_generator.signal_edge.previous_signal_state_0
rlabel metal1 s 7728 16082 7728 16082 4 noise_generator.signal_edge.signal
rlabel metal2 s 7590 19380 7590 19380 4 noise_generator.tone.counter\[0\]
rlabel metal1 s 9706 18598 9706 18598 4 noise_generator.tone.counter\[1\]
rlabel metal1 s 8372 18666 8372 18666 4 noise_generator.tone.counter\[2\]
rlabel metal1 s 10258 16660 10258 16660 4 noise_generator.tone.counter\[3\]
rlabel metal2 s 10074 17646 10074 17646 4 noise_generator.tone.counter\[4\]
rlabel metal1 s 8648 3570 8648 3570 4 pwm_A.accumulator\[0\]
rlabel metal1 s 7958 4692 7958 4692 4 pwm_A.accumulator\[1\]
rlabel metal2 s 7958 6188 7958 6188 4 pwm_A.accumulator\[2\]
rlabel metal1 s 6532 6834 6532 6834 4 pwm_A.accumulator\[3\]
rlabel metal2 s 4186 8092 4186 8092 4 pwm_A.accumulator\[4\]
rlabel metal1 s 3910 6800 3910 6800 4 pwm_A.accumulator\[5\]
rlabel metal1 s 2254 6324 2254 6324 4 pwm_A.accumulator\[6\]
rlabel metal1 s 1334 9010 1334 9010 4 pwm_A.accumulator\[7\]
rlabel metal1 s 18308 2618 18308 2618 4 pwm_B.accumulator\[0\]
rlabel metal1 s 17802 4080 17802 4080 4 pwm_B.accumulator\[1\]
rlabel metal1 s 18768 5746 18768 5746 4 pwm_B.accumulator\[2\]
rlabel metal1 s 16836 6834 16836 6834 4 pwm_B.accumulator\[3\]
rlabel metal1 s 14122 6290 14122 6290 4 pwm_B.accumulator\[4\]
rlabel metal1 s 14950 7820 14950 7820 4 pwm_B.accumulator\[5\]
rlabel metal1 s 11546 6868 11546 6868 4 pwm_B.accumulator\[6\]
rlabel metal1 s 9844 6834 9844 6834 4 pwm_B.accumulator\[7\]
rlabel metal1 s 25990 2618 25990 2618 4 pwm_C.accumulator\[0\]
rlabel metal1 s 25484 4046 25484 4046 4 pwm_C.accumulator\[1\]
rlabel metal1 s 25668 6834 25668 6834 4 pwm_C.accumulator\[2\]
rlabel metal1 s 25116 7718 25116 7718 4 pwm_C.accumulator\[3\]
rlabel metal2 s 23506 8636 23506 8636 4 pwm_C.accumulator\[4\]
rlabel metal1 s 22862 9588 22862 9588 4 pwm_C.accumulator\[5\]
rlabel metal1 s 21850 7854 21850 7854 4 pwm_C.accumulator\[6\]
rlabel metal2 s 21298 10438 21298 10438 4 pwm_C.accumulator\[7\]
rlabel metal1 s 12098 14926 12098 14926 4 restart_envelope
rlabel metal1 s 23874 30804 23874 30804 4 rst_n
rlabel metal2 s 14766 24378 14766 24378 4 tone_A_generator.counter\[0\]
rlabel metal1 s 18538 25840 18538 25840 4 tone_A_generator.counter\[10\]
rlabel metal1 s 19918 24582 19918 24582 4 tone_A_generator.counter\[11\]
rlabel metal1 s 13478 21862 13478 21862 4 tone_A_generator.counter\[1\]
rlabel metal1 s 13938 24752 13938 24752 4 tone_A_generator.counter\[2\]
rlabel metal1 s 14766 24752 14766 24752 4 tone_A_generator.counter\[3\]
rlabel metal1 s 15870 28594 15870 28594 4 tone_A_generator.counter\[4\]
rlabel metal1 s 16468 29818 16468 29818 4 tone_A_generator.counter\[5\]
rlabel metal1 s 16330 28390 16330 28390 4 tone_A_generator.counter\[6\]
rlabel metal1 s 17848 28594 17848 28594 4 tone_A_generator.counter\[7\]
rlabel metal1 s 18262 27506 18262 27506 4 tone_A_generator.counter\[8\]
rlabel metal1 s 17250 26928 17250 26928 4 tone_A_generator.counter\[9\]
rlabel metal1 s 16192 15674 16192 15674 4 tone_A_generator.out
rlabel metal1 s 14122 23596 14122 23596 4 tone_A_generator.period\[0\]
rlabel metal1 s 19320 21114 19320 21114 4 tone_A_generator.period\[10\]
rlabel metal1 s 18814 24310 18814 24310 4 tone_A_generator.period\[11\]
rlabel metal1 s 12972 23086 12972 23086 4 tone_A_generator.period\[1\]
rlabel metal1 s 14352 26418 14352 26418 4 tone_A_generator.period\[2\]
rlabel metal1 s 13708 26214 13708 26214 4 tone_A_generator.period\[3\]
rlabel metal1 s 13018 29036 13018 29036 4 tone_A_generator.period\[4\]
rlabel metal2 s 12558 27676 12558 27676 4 tone_A_generator.period\[5\]
rlabel metal1 s 15092 27982 15092 27982 4 tone_A_generator.period\[6\]
rlabel metal1 s 15410 28424 15410 28424 4 tone_A_generator.period\[7\]
rlabel metal2 s 16974 24752 16974 24752 4 tone_A_generator.period\[8\]
rlabel metal1 s 16790 21318 16790 21318 4 tone_A_generator.period\[9\]
rlabel metal2 s 27094 20060 27094 20060 4 tone_B_generator.counter\[0\]
rlabel metal1 s 24472 11186 24472 11186 4 tone_B_generator.counter\[10\]
rlabel metal1 s 25162 11084 25162 11084 4 tone_B_generator.counter\[11\]
rlabel metal1 s 23644 19278 23644 19278 4 tone_B_generator.counter\[1\]
rlabel metal1 s 24656 18734 24656 18734 4 tone_B_generator.counter\[2\]
rlabel metal1 s 25024 17782 25024 17782 4 tone_B_generator.counter\[3\]
rlabel metal1 s 24794 16966 24794 16966 4 tone_B_generator.counter\[4\]
rlabel metal1 s 24794 17034 24794 17034 4 tone_B_generator.counter\[5\]
rlabel metal1 s 23598 15572 23598 15572 4 tone_B_generator.counter\[6\]
rlabel metal1 s 24886 14450 24886 14450 4 tone_B_generator.counter\[7\]
rlabel metal2 s 24886 13906 24886 13906 4 tone_B_generator.counter\[8\]
rlabel metal1 s 25300 12614 25300 12614 4 tone_B_generator.counter\[9\]
rlabel metal1 s 19228 14450 19228 14450 4 tone_B_generator.out
rlabel metal1 s 20332 18666 20332 18666 4 tone_B_generator.period\[0\]
rlabel metal1 s 22862 11764 22862 11764 4 tone_B_generator.period\[10\]
rlabel metal1 s 22586 12410 22586 12410 4 tone_B_generator.period\[11\]
rlabel metal2 s 18722 17884 18722 17884 4 tone_B_generator.period\[1\]
rlabel metal1 s 21436 18394 21436 18394 4 tone_B_generator.period\[2\]
rlabel metal1 s 18538 19380 18538 19380 4 tone_B_generator.period\[3\]
rlabel metal2 s 21850 17476 21850 17476 4 tone_B_generator.period\[4\]
rlabel metal1 s 20010 17612 20010 17612 4 tone_B_generator.period\[5\]
rlabel metal1 s 20746 20332 20746 20332 4 tone_B_generator.period\[6\]
rlabel metal1 s 20838 19822 20838 19822 4 tone_B_generator.period\[7\]
rlabel metal1 s 22770 13498 22770 13498 4 tone_B_generator.period\[8\]
rlabel metal1 s 23506 13940 23506 13940 4 tone_B_generator.period\[9\]
rlabel metal2 s 21896 26486 21896 26486 4 tone_C_generator.counter\[0\]
rlabel metal1 s 24840 21522 24840 21522 4 tone_C_generator.counter\[10\]
rlabel metal1 s 25254 21590 25254 21590 4 tone_C_generator.counter\[11\]
rlabel metal2 s 21666 24446 21666 24446 4 tone_C_generator.counter\[1\]
rlabel metal1 s 23046 27540 23046 27540 4 tone_C_generator.counter\[2\]
rlabel metal2 s 23414 27472 23414 27472 4 tone_C_generator.counter\[3\]
rlabel metal1 s 24702 30124 24702 30124 4 tone_C_generator.counter\[4\]
rlabel metal1 s 25208 27574 25208 27574 4 tone_C_generator.counter\[5\]
rlabel metal1 s 24564 27506 24564 27506 4 tone_C_generator.counter\[6\]
rlabel metal1 s 25254 29682 25254 29682 4 tone_C_generator.counter\[7\]
rlabel metal1 s 27002 24310 27002 24310 4 tone_C_generator.counter\[8\]
rlabel metal1 s 26266 23222 26266 23222 4 tone_C_generator.counter\[9\]
rlabel metal1 s 20792 15470 20792 15470 4 tone_C_generator.out
rlabel metal1 s 21850 24140 21850 24140 4 tone_C_generator.period\[0\]
rlabel metal1 s 23506 21488 23506 21488 4 tone_C_generator.period\[10\]
rlabel metal1 s 23138 21114 23138 21114 4 tone_C_generator.period\[11\]
rlabel metal2 s 22034 24446 22034 24446 4 tone_C_generator.period\[1\]
rlabel metal1 s 21758 27336 21758 27336 4 tone_C_generator.period\[2\]
rlabel metal1 s 21482 28390 21482 28390 4 tone_C_generator.period\[3\]
rlabel metal1 s 22586 30362 22586 30362 4 tone_C_generator.period\[4\]
rlabel metal1 s 20746 29478 20746 29478 4 tone_C_generator.period\[5\]
rlabel metal1 s 20792 30362 20792 30362 4 tone_C_generator.period\[6\]
rlabel metal1 s 25116 30158 25116 30158 4 tone_C_generator.period\[7\]
rlabel metal1 s 23644 23154 23644 23154 4 tone_C_generator.period\[8\]
rlabel metal1 s 21804 22066 21804 22066 4 tone_C_generator.period\[9\]
rlabel metal1 s 15594 14892 15594 14892 4 tone_disable_A
rlabel metal2 s 18446 13974 18446 13974 4 tone_disable_B
rlabel metal1 s 18676 15674 18676 15674 4 tone_disable_C
flabel metal4 s 27256 496 27576 31056 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 20540 496 20860 31056 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 13824 496 14144 31056 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 7108 496 7428 31056 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 23898 496 24218 31056 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 17182 496 17502 31056 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 10466 496 10786 31056 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 3750 496 4070 31056 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal2 s 8758 31600 8814 32000 0 FreeSans 280 90 0 0 bc1
port 3 nsew
flabel metal2 s 10230 31600 10286 32000 0 FreeSans 280 90 0 0 bdir
port 4 nsew
flabel metal2 s 9494 0 9550 400 0 FreeSans 280 90 0 0 channel_A_dac_ctrl[0]
port 5 nsew
flabel metal2 s 3974 0 4030 400 0 FreeSans 280 90 0 0 channel_A_dac_ctrl[10]
port 6 nsew
flabel metal2 s 3422 0 3478 400 0 FreeSans 280 90 0 0 channel_A_dac_ctrl[11]
port 7 nsew
flabel metal2 s 2870 0 2926 400 0 FreeSans 280 90 0 0 channel_A_dac_ctrl[12]
port 8 nsew
flabel metal2 s 2318 0 2374 400 0 FreeSans 280 90 0 0 channel_A_dac_ctrl[13]
port 9 nsew
flabel metal2 s 1766 0 1822 400 0 FreeSans 280 90 0 0 channel_A_dac_ctrl[14]
port 10 nsew
flabel metal2 s 8942 0 8998 400 0 FreeSans 280 90 0 0 channel_A_dac_ctrl[1]
port 11 nsew
flabel metal2 s 8390 0 8446 400 0 FreeSans 280 90 0 0 channel_A_dac_ctrl[2]
port 12 nsew
flabel metal2 s 7838 0 7894 400 0 FreeSans 280 90 0 0 channel_A_dac_ctrl[3]
port 13 nsew
flabel metal2 s 7314 200 7314 200 0 FreeSans 280 90 0 0 channel_A_dac_ctrl[4]
flabel metal2 s 6734 0 6790 400 0 FreeSans 280 90 0 0 channel_A_dac_ctrl[5]
port 15 nsew
flabel metal2 s 6182 0 6238 400 0 FreeSans 280 90 0 0 channel_A_dac_ctrl[6]
port 16 nsew
flabel metal2 s 5630 0 5686 400 0 FreeSans 280 90 0 0 channel_A_dac_ctrl[7]
port 17 nsew
flabel metal2 s 5078 0 5134 400 0 FreeSans 280 90 0 0 channel_A_dac_ctrl[8]
port 18 nsew
flabel metal2 s 4526 0 4582 400 0 FreeSans 280 90 0 0 channel_A_dac_ctrl[9]
port 19 nsew
flabel metal2 s 4342 31600 4398 32000 0 FreeSans 280 90 0 0 channel_A_pwm_out
port 20 nsew
flabel metal2 s 17774 0 17830 400 0 FreeSans 280 90 0 0 channel_B_dac_ctrl[0]
port 21 nsew
flabel metal2 s 12254 0 12310 400 0 FreeSans 280 90 0 0 channel_B_dac_ctrl[10]
port 22 nsew
flabel metal2 s 11702 0 11758 400 0 FreeSans 280 90 0 0 channel_B_dac_ctrl[11]
port 23 nsew
flabel metal2 s 11150 0 11206 400 0 FreeSans 280 90 0 0 channel_B_dac_ctrl[12]
port 24 nsew
flabel metal2 s 10598 0 10654 400 0 FreeSans 280 90 0 0 channel_B_dac_ctrl[13]
port 25 nsew
flabel metal2 s 10046 0 10102 400 0 FreeSans 280 90 0 0 channel_B_dac_ctrl[14]
port 26 nsew
flabel metal2 s 17222 0 17278 400 0 FreeSans 280 90 0 0 channel_B_dac_ctrl[1]
port 27 nsew
flabel metal2 s 16670 0 16726 400 0 FreeSans 280 90 0 0 channel_B_dac_ctrl[2]
port 28 nsew
flabel metal2 s 16118 0 16174 400 0 FreeSans 280 90 0 0 channel_B_dac_ctrl[3]
port 29 nsew
flabel metal2 s 15566 0 15622 400 0 FreeSans 280 90 0 0 channel_B_dac_ctrl[4]
port 30 nsew
flabel metal2 s 15014 0 15070 400 0 FreeSans 280 90 0 0 channel_B_dac_ctrl[5]
port 31 nsew
flabel metal2 s 14462 0 14518 400 0 FreeSans 280 90 0 0 channel_B_dac_ctrl[6]
port 32 nsew
flabel metal2 s 13938 200 13938 200 0 FreeSans 280 90 0 0 channel_B_dac_ctrl[7]
flabel metal2 s 13358 0 13414 400 0 FreeSans 280 90 0 0 channel_B_dac_ctrl[8]
port 34 nsew
flabel metal2 s 12806 0 12862 400 0 FreeSans 280 90 0 0 channel_B_dac_ctrl[9]
port 35 nsew
flabel metal2 s 2870 31600 2926 32000 0 FreeSans 280 90 0 0 channel_B_pwm_out
port 36 nsew
flabel metal2 s 26054 0 26110 400 0 FreeSans 280 90 0 0 channel_C_dac_ctrl[0]
port 37 nsew
flabel metal2 s 20562 200 20562 200 0 FreeSans 280 90 0 0 channel_C_dac_ctrl[10]
flabel metal2 s 19982 0 20038 400 0 FreeSans 280 90 0 0 channel_C_dac_ctrl[11]
port 39 nsew
flabel metal2 s 19430 0 19486 400 0 FreeSans 280 90 0 0 channel_C_dac_ctrl[12]
port 40 nsew
flabel metal2 s 18878 0 18934 400 0 FreeSans 280 90 0 0 channel_C_dac_ctrl[13]
port 41 nsew
flabel metal2 s 18326 0 18382 400 0 FreeSans 280 90 0 0 channel_C_dac_ctrl[14]
port 42 nsew
flabel metal2 s 25502 0 25558 400 0 FreeSans 280 90 0 0 channel_C_dac_ctrl[1]
port 43 nsew
flabel metal2 s 24950 0 25006 400 0 FreeSans 280 90 0 0 channel_C_dac_ctrl[2]
port 44 nsew
flabel metal2 s 24398 0 24454 400 0 FreeSans 280 90 0 0 channel_C_dac_ctrl[3]
port 45 nsew
flabel metal2 s 23846 0 23902 400 0 FreeSans 280 90 0 0 channel_C_dac_ctrl[4]
port 46 nsew
flabel metal2 s 23294 0 23350 400 0 FreeSans 280 90 0 0 channel_C_dac_ctrl[5]
port 47 nsew
flabel metal2 s 22742 0 22798 400 0 FreeSans 280 90 0 0 channel_C_dac_ctrl[6]
port 48 nsew
flabel metal2 s 22190 0 22246 400 0 FreeSans 280 90 0 0 channel_C_dac_ctrl[7]
port 49 nsew
flabel metal2 s 21638 0 21694 400 0 FreeSans 280 90 0 0 channel_C_dac_ctrl[8]
port 50 nsew
flabel metal2 s 21086 0 21142 400 0 FreeSans 280 90 0 0 channel_C_dac_ctrl[9]
port 51 nsew
flabel metal2 s 1398 31600 1454 32000 0 FreeSans 280 90 0 0 channel_C_pwm_out
port 52 nsew
flabel metal2 s 24950 31600 25006 32000 0 FreeSans 280 90 0 0 clk
port 53 nsew
flabel metal2 s 7286 31600 7342 32000 0 FreeSans 280 90 0 0 clock_select[0]
port 54 nsew
flabel metal2 s 5814 31600 5870 32000 0 FreeSans 280 90 0 0 clock_select[1]
port 55 nsew
flabel metal2 s 22006 31600 22062 32000 0 FreeSans 280 90 0 0 data[0]
port 56 nsew
flabel metal2 s 20534 31600 20590 32000 0 FreeSans 280 90 0 0 data[1]
port 57 nsew
flabel metal2 s 19062 31600 19118 32000 0 FreeSans 280 90 0 0 data[2]
port 58 nsew
flabel metal2 s 17590 31600 17646 32000 0 FreeSans 280 90 0 0 data[3]
port 59 nsew
flabel metal2 s 16118 31600 16174 32000 0 FreeSans 280 90 0 0 data[4]
port 60 nsew
flabel metal2 s 14646 31600 14702 32000 0 FreeSans 280 90 0 0 data[5]
port 61 nsew
flabel metal2 s 13174 31600 13230 32000 0 FreeSans 280 90 0 0 data[6]
port 62 nsew
flabel metal2 s 11702 31600 11758 32000 0 FreeSans 280 90 0 0 data[7]
port 63 nsew
flabel metal2 s 26422 31600 26478 32000 0 FreeSans 280 90 0 0 ena
port 64 nsew
flabel metal2 s 23478 31600 23534 32000 0 FreeSans 280 90 0 0 rst_n
port 65 nsew
<< properties >>
string FIXED_BBOX 0 0 28000 32000
string GDS_END 3773574
string GDS_FILE ../gds/ay8913.gds
string GDS_START 552086
<< end >>
